module  ep2c61a(
   sys_clk,
   rst_n,
   ofc3555,
   mg1aaad,
   jcd5569,
   jraab4b,
   vv55a5f,
   vkad2fe,
   lq697f3,
   kd4bf9b,
   jp5fcdc,
   lqfe6e7,
   thf373b,
   bn9b9df,
   aldceff,
   ofe77fc,
   ym3bfe4,
   jpd27c8,
   do93e46,
   mt9f233,
   hq99d4a,
   qgcea52,
   en75290,
   mt18edf,
   hbc76fc,
   ie3b7e7,
   sudbf39,
   fadf9c9,
   hbfce4b,
   mre725f,
   kf392fc,
   gbc97e4,
   cz4bf24,
   xj5f924,
   vvfc927,
   tue493f,
   mg249fa,
   ie24fd0,
   fp27e80,
   je3f407,
   ayfa03b,
`ifdef AER
   hod01d9,
   sj80ecb,
   ux765d,
   ie3b2ed,
   uvd9769 ,
   uicbb4d,
   jc5da68,
   iped342,
   lq69a15,
   fa4d0aa,
`endif
   ym1549d,
   zzaa4e9,
   ne5274e,
   je93a72,
   gq9d393,
   pfe9c99,
   mr4e4ce,
   ay72675,
   do933a9,
   wlb4393,
   uxa1c9c,
   vke4e4,
`ifdef AER
   zxece0b,
`endif
   me6705e,
   lf382f0,
   mec1786
   );
parameter twbc30 = 3'b111;
parameter uvc3724   = 2'b00;
parameter je1b925  = 2'b01;
parameter mrdc92b = 2'b10;
input                     sys_clk;
input                     rst_n;
input  [7:0]              ofc3555;
input  [7:0]              mg1aaad;
input  [7:0]              jcd5569;
input  [11:0]             jraab4b;
input  [11:0]             vv55a5f;
input  [11:0]             vkad2fe;
input  [6:0]              lq697f3;
input  [10:0]             kd4bf9b;
input  [6:0]              jp5fcdc;
input  [10:0]             lqfe6e7;
input  [6:0]              thf373b;
input  [10:0]             bn9b9df;
input                     aldceff;
input                     ofe77fc;
input                     ym3bfe4;
input                     jpd27c8;
input                     do93e46;
input                     mt9f233;
input                     hq99d4a;
input                     qgcea52;
input                     en75290;
input                     mt18edf;
input                     hbc76fc;
input                     ie3b7e7;
input                     sudbf39;
input                     fadf9c9;
input                     hbfce4b;
input                     mre725f;
input                     kf392fc;
input                     gbc97e4;
input                     cz4bf24;
input                     xj5f924;
input                     vvfc927;
input [7:0]                tue493f;
input [7:0]                mg249fa;
input [7:0]                ie24fd0;
input                     fp27e80;
input                     je3f407;
input                     ayfa03b;
`ifdef AER
input                     hod01d9;
input                     sj80ecb;
input                     ux765d;
input                     ie3b2ed;
input                     uvd9769;
input  [8:0]              uicbb4d;
input                     jc5da68;
input                     iped342;
input                     lq69a15;
input                     fa4d0aa;
`endif
output                    ym1549d;
output                    zzaa4e9;
output                    ne5274e;
output                    je93a72;
output                    gq9d393;
output                    pfe9c99;
output                    mr4e4ce;
output                    ay72675;
output                    do933a9;
output                    wlb4393;
output                    uxa1c9c;
output                    vke4e4;
output [23:0]             me6705e;
output [23:0]             lf382f0;
output [23:0]             mec1786;
`ifdef AER
output                    zxece0b;
`endif
reg                       ym1549d;
reg                       zzaa4e9;
reg                       ne5274e;
reg                       je93a72;
reg                       gq9d393;
reg                       pfe9c99;
reg                       mr4e4ce;
reg                       ay72675;
reg                       do933a9;
reg                       wlb4393;
reg                       uxa1c9c;
reg                       vke4e4;
reg                       zxece0b;
wire   [23:0]             me6705e;
wire   [23:0]             lf382f0;
wire   [23:0]             mec1786;
`ifdef CUMULATIVE_CREDIT_CHECK
reg  [7:0]                vvf37aa, rv9bd57, wwdeabf;
reg  [11:0]               kqf55f9,   dbaafc8,   xw57e47,   rvbf23b,   pff91df;
reg  [11:0]               vvc8efe,  vi477f7,  qi3bfbb,  bydfdd8,  zkfeec3;
reg  [11:0]               wjf761a, yzbb0d5, thd86ad, ofc356f, mg1ab7d;
`endif
reg  [11:0]               jcd5be9;
reg  [7:0]                doadf4a;
reg  [11:0]               uv6fa52;
reg  [7:0]                cm7d295;
reg  [11:0]               vve94a8;
reg  [7:0]                nr4a547;
reg                       jc52a3f;
reg                       ir951fb;
reg                       zma8fdd;
reg  [2:0]                ne47eea;
reg  [2:0]                ba3f752;
reg  [13:0]               psfba93;
reg  [13:0]               vvdd49a;
reg  [13:0]               cmea4d7;
reg  [6:0]                lq526b8;
reg  [11:0]               tw935c2;
reg  [6:0]                gd9ae12;
reg  [11:0]               pfd7095;
reg  [6:0]                zmb84ae;
reg  [11:0]               xjc2572;
reg  [7:0]                ir12b97;
reg  [11:0]               an95cbd;
reg  [7:0]                kfae5ec;
reg  [11:0]               ww72f64;
reg  [7:0]                sw97b20;
reg  [11:0]               babd901;
reg  [7:0]                rtec80b;
reg  [11:0]               dz6405e;
wire [7:0]                tw202f7;
wire [11:0]               ri17bb;
wire [7:0]                hqbdda;
wire [11:0]               kd5eed2;
reg                       uvf7695;
reg                       irbb4ad;
reg                       tuda56d;
reg                       ldd2b6a;
wire                      yz95b57;
wire                      twadabc;
wire                      qg6d5e2;
wire                      yx6af11;
wire                      jc5788d;
wire                      gqbc46b;
wire                      ale2358;
wire                      ri11ac4;
wire                      ou8d622;
wire                      pf6b110;
wire                      lq58886;
wire                      wwc4432;
wire                      xl22190;
wire                      sw10c86;
wire                      xy86430;
wire                      jr32183;
wire                      yz90c1f;
wire                      tw860fc;
wire [5:0]                ba307e3;
`ifdef CUMULATIVE_CREDIT_CHECK
`else
`endif
`ifdef AER
`endif
reg [7 : 0] hq83f1a;
reg [7 : 0] ec1f8d2;
reg [7 : 0] zxfc691;
reg [11 : 0] xje348e;
reg [11 : 0] sw1a476;
reg [11 : 0] dzd23b0;
reg [6 : 0] jr91d86;
reg [10 : 0] fp8ec36;
reg [6 : 0] tu761b6;
reg [10 : 0] bnb0db3;
reg [6 : 0] ls86d9f;
reg [10 : 0] mt36cfa;
reg qib67d4;
reg aab3ea1;
reg an9f508;
reg mefa844;
reg uid4220;
reg sja1101;
reg kf880d;
reg mr4406d;
reg tw2036c;
reg ri1b63;
reg mtdb1b;
reg ay6d8dd;
reg vi6c6e8;
reg lq63743;
reg ba1ba1a;
reg bldd0d3;
reg ale869f;
reg yk434fd;
reg ou1a7e9;
reg wjd3f48;
reg ir9fa45;
reg [7 : 0] enfd22d;
reg [7 : 0] lde916c;
reg [7 : 0] jc48b67;
reg fn45b3b;
reg vx2d9df;
reg ho6cefe;
reg [11 : 0] yk677f2;
reg [7 : 0] aa3bf90;
reg [11 : 0] dmdfc80;
reg [7 : 0] psfe403;
reg [11 : 0] yxf201b;
reg [7 : 0] oh900dd;
reg wl806ed;
reg xl376c;
reg hq1bb67;
reg [2 : 0] xjddb3b;
reg [2 : 0] qted9de;
reg [13 : 0] tu6cef4;
reg [13 : 0] qg677a2;
reg [13 : 0] ou3bd10;
reg [6 : 0] kqde880;
reg [11 : 0] tuf4401;
reg [6 : 0] vka200a;
reg [11 : 0] co10052;
reg [6 : 0] ep80291;
reg [11 : 0] hq148c;
reg [7 : 0] eca462;
reg [11 : 0] ps52311;
reg [7 : 0] bn9188a;
reg [11 : 0] ri8c456;
reg [7 : 0] kq622b2;
reg [11 : 0] tw11590;
reg [7 : 0] kf8ac83;
reg [11 : 0] go5641c;
reg [7 : 0] fcb20e0;
reg [11 : 0] sj90703;
reg [7 : 0] ba8381d;
reg [11 : 0] lf1c0ea;
reg aye0757;
reg xl3ab9;
reg ep1d5ce;
reg wweae75;
reg tu573a9;
reg ecb9d4a;
reg mecea51;
reg yx75288;
reg iea9444;
reg nr4a221;
reg kd5110f;
reg ou8887d;
reg sh443e9;
reg ou21f4c;
reg ymfa60;
reg os7d300;
reg nre9800;
reg ui4c006;
reg kd60030;
reg wy185;
reg ukc28;
reg lf6141;
reg [5 : 0] pu30a0f;
reg [2047:0] necf6c2;
wire [93:0] ld7b613;
`ifdef AER
`endif
`ifdef AER
`endif
`ifdef CUMULATIVE_CREDIT_CHECK
`endif
`ifdef CUMULATIVE_CREDIT_CHECK
`else
`endif
`ifdef AER
`endif
localparam qgdb09f = 94,nrd84f8 = 32'hfdffca8b;
localparam [31:0] thc27c7 = nrd84f8;
localparam mt9f1ff = nrd84f8 & 4'hf;
localparam [11:0] fnc7fe5 = 'h7ff;
wire  [(1 << mt9f1ff)  -1:0] suff972;
reg    [qgdb09f-1:0] cme5c87;
reg [mt9f1ff-1:0] qg721c0 [0:1];
reg [mt9f1ff-1:0] ym8700c;
reg rv38061;
integer jcc030e;
integer vk1872;
`ifdef AER
`endif
`ifdef AER
`endif
`ifdef CUMULATIVE_CREDIT_CHECK
`endif
`ifdef CUMULATIVE_CREDIT_CHECK
`else
`endif
`ifdef AER
`endif
`ifdef AER
`endif
`ifdef AER
`endif
`ifdef CUMULATIVE_CREDIT_CHECK
`endif
assign me6705e   = {2'b00, aa3bf90, 2'b00, yk677f2};
assign lf382f0  = {2'b00, psfe403, 2'b00, dmdfc80};
assign mec1786 = {2'b00, oh900dd, 2'b00, yxf201b};
assign ale2358   = (hq83f1a == 0);
assign ri11ac4   = (xje348e == 0);
assign ou8d622  = (ec1f8d2 == 0);
assign pf6b110  = (sw1a476 == 0);
assign lq58886 = (zxfc691 == 0);
assign wwc4432 = (dzd23b0 == 0);
assign yx6af11 = yk434fd | fn45b3b;
assign jc5788d = ou1a7e9 | vx2d9df;
assign gqbc46b = bldd0d3 | ho6cefe;
assign ba307e3 = (vx2d9df) ? (lde916c + 1'b1) : lde916c;
`ifdef CUMULATIVE_CREDIT_CHECK
always @(posedge sys_clk or negedge rst_n) begin   if (rst_n == 1'b0) begin      kqf55f9            <= 12'd0;      dbaafc8            <= 12'd0;      xw57e47            <= 12'd0;      rvbf23b         <= 12'd0;      pff91df   <= 12'd0;      vvc8efe           <= 12'd0;      vi477f7           <= 12'd0;      qi3bfbb           <= 12'd0;      bydfdd8        <= 12'd0;      zkfeec3  <= 12'd0;      wjf761a          <= 12'd0;      yzbb0d5          <= 12'd0;      thd86ad          <= 12'd0;      ofc356f       <= 12'd0;      mg1ab7d <= 12'd0;      vvf37aa            <= 8'd0;      rv9bd57           <= 8'd0;      wwdeabf          <= 8'd0;   end   else begin                  if(qib67d4) begin            dbaafc8  <= 12'd0;         xw57e47  <= 12'd0;      end      else begin                  dbaafc8 <= (ale869f) ? (dbaafc8 + enfd22d) : dbaafc8;
                  xw57e47  <= (mefa844) ? kqf55f9 : xw57e47;       end                  rvbf23b       <= dbaafc8 - xw57e47;                  pff91df <= kqf55f9 - xw57e47;                  if(rvbf23b <= 12'd2047)                      kqf55f9 <= dbaafc8;      else if(pff91df <= 12'd2047)           kqf55f9 <= xw57e47 + 12'd2047;            if(qib67d4) begin            vi477f7  <= 12'd0;         qi3bfbb  <= 12'd0;      end      else begin         case({ou1a7e9, vx2d9df})            2'b01   : vi477f7  <= vi477f7 + 1'b1;            2'b10,            2'b11   : vi477f7  <= vi477f7 + pu30a0f;            default : vi477f7  <= vi477f7;         endcase         qi3bfbb  <= (uid4220) ? vvc8efe : qi3bfbb;      end      bydfdd8       <= vi477f7 - qi3bfbb;      zkfeec3 <= vvc8efe - qi3bfbb;      if(bydfdd8 <= 12'd2047)         vvc8efe <= vi477f7;      else if(zkfeec3 <= 12'd2047)         vvc8efe <= qi3bfbb + 12'd2047;            if(qib67d4) begin            yzbb0d5  <= 12'd0;         thd86ad  <= 12'd0;      end      else begin         yzbb0d5  <= (ir9fa45) ? (yzbb0d5 + jc48b67) : yzbb0d5;         thd86ad  <= (sja1101) ? wjf761a : thd86ad;      end      ofc356f       <= yzbb0d5 - thd86ad;      mg1ab7d <= wjf761a - thd86ad;      if(ofc356f <= 12'd2047)         wjf761a <= yzbb0d5;      else if(mg1ab7d <= 12'd2047)         wjf761a <= thd86ad + 12'd2047;                  if(qib67d4) begin            vvf37aa   <= 8'd0;         rv9bd57  <= 8'd0;         wwdeabf <= 8'd0;      end      else begin         vvf37aa   <= (bldd0d3) ? (vvf37aa + 1'b1) : vvf37aa;         rv9bd57  <= (yk434fd) ? (rv9bd57 + 1'b1) : rv9bd57;         wwdeabf <= (wjd3f48) ? (wwdeabf + 1'b1) : wwdeabf;      end   end
end
always @(posedge sys_clk or negedge rst_n) begin   if (rst_n == 1'b0) begin      doadf4a    <= 8'd0;      cm7d295   <= 8'd0;      nr4a547  <= 8'd0;      jcd5be9   <= 12'd0;      uv6fa52  <= 12'd0;      vve94a8 <= 12'd0;   end   else begin            doadf4a     <= (!kd5110f) ? (hq83f1a + vvf37aa) : hq83f1a;      jcd5be9    <= (!ou8887d) ? (xje348e + kqf55f9) : xje348e;            cm7d295    <= (!sh443e9) ? (ec1f8d2 + rv9bd57) : ec1f8d2;      uv6fa52   <= (!ou21f4c) ? (sw1a476 + vvc8efe) : sw1a476;            nr4a547   <= (!ymfa60) ? (zxfc691 + wwdeabf) : zxfc691;      vve94a8  <= (!os7d300) ? (dzd23b0 + wjf761a) : dzd23b0;   end
end
`else
always @(posedge sys_clk or negedge rst_n) begin   if (rst_n == 1'b0) begin         doadf4a    <= 8'd0;         cm7d295   <= 8'd0;         nr4a547  <= 8'd0;         jcd5be9   <= 12'd0;         uv6fa52  <= 12'd0;         vve94a8 <= 12'd0;   end   else begin      if(qib67d4) begin            doadf4a    <= hq83f1a;         cm7d295   <= ec1f8d2;         nr4a547  <= zxfc691;         jcd5be9   <= xje348e;         uv6fa52  <= sw1a476;         vve94a8 <= dzd23b0;      end      else begin                  if (!kd5110f && bldd0d3 && ho6cefe)            doadf4a <= (aa3bf90 + 2) ;         else if (!kd5110f && nr4a221)            doadf4a <= (aa3bf90 + 1) ;         jcd5be9   <= (!ou8887d && ale869f) ? (yk677f2 + enfd22d) : yk677f2;                  if (!sh443e9 && yk434fd && fn45b3b)            cm7d295 <= (psfe403 + 2) ;         else if (!sh443e9 && yx75288)            cm7d295 <= (psfe403 + 1) ;         if (!ou21f4c) begin            case({ou1a7e9, vx2d9df})               2'b01   : uv6fa52  <= dmdfc80 + 1'b1;               2'b10,               2'b11   : uv6fa52  <= dmdfc80 + pu30a0f;               default : uv6fa52  <= dmdfc80;            endcase         end                  nr4a547  <= (!ymfa60 && wjd3f48) ? (oh900dd + 1) : oh900dd;         vve94a8 <= (!os7d300 && ir9fa45) ? (yxf201b + jc48b67) : yxf201b;      end   end
end
`endif
`ifdef AER
assign tw202f7   = aa3bf90   - eca462;
assign ri17bb   = yk677f2  - ps52311;
assign hqbdda  = psfe403  - bn9188a;
assign kd5eed2  = dmdfc80 - ri8c456;
always @(posedge sys_clk or negedge rst_n) begin   if (rst_n == 1'b0) begin      ir12b97        <= 8'd0;      an95cbd       <= 12'd0;      kfae5ec       <= 8'd0;      ww72f64      <= 12'd0;      sw97b20   <= 8'd0;      babd901  <= 12'd0;      rtec80b  <= 8'd0;      dz6405e <= 12'd0;            uvf7695     <= 1'b0;      irbb4ad     <= 1'b0;      tuda56d    <= 1'b0;      ldd2b6a    <= 1'b0;      zxece0b        <= 1'b0;   end   else begin            if(hod01d9) begin            sw97b20   <= (!kd5110f  && sj80ecb)  ? eca462   : kq622b2;         babd901  <= (!ou8887d  && ux765d)  ? ps52311  : tw11590;         rtec80b  <= (!sh443e9 && ie3b2ed) ? bn9188a  : kf8ac83;         dz6405e <= (!ou21f4c && uvd9769) ? ri8c456 : go5641c;      end                  uvf7695  <= (fcb20e0  >= 'd128)  ? 1'b1 : 1'b0;      irbb4ad  <= (sj90703  >= 'd2048) ? 1'b1 : 1'b0;      tuda56d <= (ba8381d >= 'd128)  ? 1'b1 : 1'b0;      ldd2b6a <= (lf1c0ea >= 'd2048) ? 1'b1 : 1'b0;      zxece0b     <= aye0757 | xl3ab9 | ep1d5ce | wweae75;            if(qib67d4)          ir12b97      <= 8'd0;      else if(!kd5110f && hod01d9) begin            if(sj80ecb)            ir12b97      <= eca462 + 1;         else if(aye0757 || xl3ab9 || jc5da68)            ir12b97      <= kq622b2;      end      if(qib67d4)          an95cbd     <= 12'd0;      else if(!ou8887d && hod01d9) begin            if(ux765d)            an95cbd     <= ps52311 + uicbb4d;         else if(aye0757 || xl3ab9 || iped342)            an95cbd     <= tw11590;      end      if(qib67d4)          kfae5ec     <= 8'd0;      else if(!sh443e9 && hod01d9) begin            if(ie3b2ed)            kfae5ec     <= bn9188a + 1;         else if(ep1d5ce || wweae75 || lq69a15)            kfae5ec     <= kf8ac83;      end      if(qib67d4)          ww72f64     <= 12'd0;      else if(!ou21f4c && hod01d9) begin            if(uvd9769)            ww72f64    <= ri8c456 + uicbb4d;         else if(ep1d5ce || wweae75 || fa4d0aa)            ww72f64    <= go5641c;      end   end
end
`endif
always @(posedge sys_clk or negedge rst_n) begin   if (rst_n == 1'b0) begin      jc52a3f      <= 1'b0;      ir951fb     <= 1'b0;      zma8fdd    <= 1'b0;      wlb4393   <= 1'b0;      uxa1c9c  <= 1'b0;      vke4e4 <= 1'b0;   end   else begin                        jc52a3f    <= mefa844 | wlb4393 | qib67d4 | !an9f508;      ir951fb   <= uid4220 | uxa1c9c | qib67d4 | !an9f508;      zma8fdd  <= sja1101 | vke4e4 | qib67d4 | !an9f508;            wlb4393   <= ((hq83f1a == 0)   && (xje348e == 0))   ? 1'b1 : 1'b0;      uxa1c9c  <= ((ec1f8d2 == 0)  && (sw1a476 == 0))  ? 1'b1 : 1'b0;      vke4e4 <= ((zxfc691 == 0) && (dzd23b0 == 0)) ? 1'b1 : 1'b0;   end
end
assign yz95b57   = kf880d | wl806ed;
assign twadabc  = mr4406d | xl376c;
assign qg6d5e2 = tw2036c | hq1bb67;
always @(posedge sys_clk or negedge rst_n) begin   if (rst_n == 1'b0) begin      ne47eea    <= 0;      ba3f752  <= 0;      ym1549d       <= 1'b0;      zzaa4e9      <= 1'b0;      ne5274e     <= 1'b0;   end   else begin                                    if(ym1549d) begin         if(tu573a9)            ym1549d  <= 1'b0;      end      else         ym1549d   <= (ri1b63 & nr4a221) | (mtdb1b & ale869f);                              if(zzaa4e9) begin         if(ecb9d4a)            zzaa4e9  <= 1'b0;      end      else         zzaa4e9  <= (ay6d8dd & yx75288) | (vi6c6e8 & iea9444) ;      if(ne5274e) begin         if(mecea51)            ne5274e  <= 1'b0;      end      else         ne5274e <= (lq63743 & wjd3f48) | (ba1ba1a & ir9fa45);                           end
end
assign xl22190   = (kqde880 == (jr91d86 - 1)) ? 1'b1 : 1'b0;
assign xy86430  = (vka200a == (tu761b6 - 1)) ? 1'b1 : 1'b0;
assign yz90c1f = (ep80291 == (ls86d9f - 1)) ? 1'b1 : 1'b0;
assign sw10c86   = (tuf4401 >= fp8ec36) ? 1'b1 : 1'b0;
assign jr32183  = (co10052 >= bnb0db3) ? 1'b1 : 1'b0;
assign tw860fc = (hq148c >= mt36cfa) ? 1'b1 : 1'b0;
always @(posedge sys_clk or negedge rst_n) begin   if (rst_n == 1'b0) begin      lq526b8    <= 0;      tw935c2    <= 0;      gd9ae12   <= 0;      pfd7095   <= 0;      zmb84ae  <= 0;      xjc2572  <= 0;      psfba93           <= 0;      vvdd49a          <= 0;      cmea4d7         <= 0;      je93a72      <= 1'b0;      gq9d393     <= 1'b0;      pfe9c99    <= 1'b0;   end   else begin                              if(ri1b63 || wl806ed || (nre9800 && nr4a221))         lq526b8  <= 0;      else         lq526b8  <= (nr4a221) ? (kqde880 + 1) : kqde880;
      if(mtdb1b || wl806ed || ui4c006)         tw935c2  <= 0;      else if (ale869f)         tw935c2  <= tuf4401 + enfd22d;            if(ay6d8dd || xl376c || (kd60030 && yx75288))         gd9ae12  <= 0;      else         gd9ae12  <= (yx75288) ? (vka200a + 1) : vka200a;
      if(vi6c6e8 || xl376c || wy185)         pfd7095  <= 0;      else if (ou1a7e9)         pfd7095  <= co10052 + lde916c;
            if(lq63743 || hq1bb67 || (ukc28 && wjd3f48))         zmb84ae  <= 0;      else        zmb84ae  <= (wjd3f48) ? (ep80291 + 1) : ep80291;
      if(ba1ba1a || hq1bb67 || lf6141)         xjc2572  <= 0;      else if (ir9fa45)         xjc2572  <= hq148c + jc48b67;            if(je93a72) begin         if(tu573a9)            je93a72  <= 1'b0;      end      else         je93a72   <= (nr4a221 && nre9800) | (ui4c006) |                         (!wl806ed && aab3ea1);      if(gq9d393) begin         if(ecb9d4a)            gq9d393  <= 1'b0;      end      else         gq9d393  <= (yx75288 && kd60030) | (wy185) |                         (!xl376c && aab3ea1);      if(pfe9c99) begin         if(mecea51)            pfe9c99  <= 1'b0;      end      else         pfe9c99 <= (wjd3f48 && ukc28) | (lf6141) |                         (!hq1bb67 && aab3ea1);   end
end
always @(posedge sys_clk or negedge rst_n) begin   if (rst_n == 1'b0) begin                  mr4e4ce       <= 1'b0;      ay72675      <= 1'b0;      do933a9     <= 1'b0;   end   else begin                  if(mr4e4ce) begin         if(tu573a9)            mr4e4ce  <= 1'b0;      end      else         mr4e4ce   <=  !wl806ed && (nr4a221 | ale869f);               if(ay72675) begin         if(ecb9d4a)            ay72675  <= 1'b0;      end      else         ay72675   <=  !xl376c && ((yx75288) | (iea9444));      if(do933a9) begin         if(mecea51)            do933a9  <= 1'b0;      end      else         do933a9 <=  !hq1bb67 && (wjd3f48 | ir9fa45);            end
end
always@* begin hq83f1a<={ofc3555>>1,ld7b613[0]};ec1f8d2<={mg1aaad>>1,ld7b613[1]};zxfc691<={jcd5569>>1,ld7b613[2]};xje348e<={jraab4b>>1,ld7b613[3]};sw1a476<={vv55a5f>>1,ld7b613[4]};dzd23b0<={vkad2fe>>1,ld7b613[5]};jr91d86<={lq697f3>>1,ld7b613[6]};fp8ec36<={kd4bf9b>>1,ld7b613[7]};tu761b6<={jp5fcdc>>1,ld7b613[8]};bnb0db3<={lqfe6e7>>1,ld7b613[9]};ls86d9f<={thf373b>>1,ld7b613[10]};mt36cfa<={bn9b9df>>1,ld7b613[11]};qib67d4<=ld7b613[12];aab3ea1<=ld7b613[13];an9f508<=ld7b613[14];mefa844<=ld7b613[15];uid4220<=ld7b613[16];sja1101<=ld7b613[17];kf880d<=ld7b613[18];mr4406d<=ld7b613[19];tw2036c<=ld7b613[20];ri1b63<=ld7b613[21];mtdb1b<=ld7b613[22];ay6d8dd<=ld7b613[23];vi6c6e8<=ld7b613[24];lq63743<=ld7b613[25];ba1ba1a<=ld7b613[26];bldd0d3<=ld7b613[27];ale869f<=ld7b613[28];yk434fd<=ld7b613[29];ou1a7e9<=ld7b613[30];wjd3f48<=ld7b613[31];ir9fa45<=ld7b613[32];enfd22d<={tue493f>>1,ld7b613[33]};lde916c<={mg249fa>>1,ld7b613[34]};jc48b67<={ie24fd0>>1,ld7b613[35]};fn45b3b<=ld7b613[36];vx2d9df<=ld7b613[37];ho6cefe<=ld7b613[38];yk677f2<={jcd5be9>>1,ld7b613[39]};aa3bf90<={doadf4a>>1,ld7b613[40]};dmdfc80<={uv6fa52>>1,ld7b613[41]};psfe403<={cm7d295>>1,ld7b613[42]};yxf201b<={vve94a8>>1,ld7b613[43]};oh900dd<={nr4a547>>1,ld7b613[44]};wl806ed<=ld7b613[45];xl376c<=ld7b613[46];hq1bb67<=ld7b613[47];xjddb3b<={ne47eea>>1,ld7b613[48]};qted9de<={ba3f752>>1,ld7b613[49]};tu6cef4<={psfba93>>1,ld7b613[50]};qg677a2<={vvdd49a>>1,ld7b613[51]};ou3bd10<={cmea4d7>>1,ld7b613[52]};kqde880<={lq526b8>>1,ld7b613[53]};tuf4401<={tw935c2>>1,ld7b613[54]};vka200a<={gd9ae12>>1,ld7b613[55]};co10052<={pfd7095>>1,ld7b613[56]};ep80291<={zmb84ae>>1,ld7b613[57]};hq148c<={xjc2572>>1,ld7b613[58]};eca462<={ir12b97>>1,ld7b613[59]};ps52311<={an95cbd>>1,ld7b613[60]};bn9188a<={kfae5ec>>1,ld7b613[61]};ri8c456<={ww72f64>>1,ld7b613[62]};kq622b2<={sw97b20>>1,ld7b613[63]};tw11590<={babd901>>1,ld7b613[64]};kf8ac83<={rtec80b>>1,ld7b613[65]};go5641c<={dz6405e>>1,ld7b613[66]};fcb20e0<={tw202f7>>1,ld7b613[67]};sj90703<={ri17bb>>1,ld7b613[68]};ba8381d<={hqbdda>>1,ld7b613[69]};lf1c0ea<={kd5eed2>>1,ld7b613[70]};aye0757<=ld7b613[71];xl3ab9<=ld7b613[72];ep1d5ce<=ld7b613[73];wweae75<=ld7b613[74];tu573a9<=ld7b613[75];ecb9d4a<=ld7b613[76];mecea51<=ld7b613[77];yx75288<=ld7b613[78];iea9444<=ld7b613[79];nr4a221<=ld7b613[80];kd5110f<=ld7b613[81];ou8887d<=ld7b613[82];sh443e9<=ld7b613[83];ou21f4c<=ld7b613[84];ymfa60<=ld7b613[85];os7d300<=ld7b613[86];nre9800<=ld7b613[87];ui4c006<=ld7b613[88];kd60030<=ld7b613[89];wy185<=ld7b613[90];ukc28<=ld7b613[91];lf6141<=ld7b613[92];pu30a0f<={ba307e3>>1,ld7b613[93]};end
always@* begin necf6c2[2047]<=mg1aaad[0];necf6c2[2046]<=jcd5569[0];necf6c2[2044]<=jraab4b[0];necf6c2[2040]<=vv55a5f[0];necf6c2[2032]<=vkad2fe[0];necf6c2[2028]<=tw860fc;necf6c2[2017]<=lq697f3[0];necf6c2[2008]<=ba307e3[0];necf6c2[1988]<=yz95b57;necf6c2[1987]<=kd4bf9b[0];necf6c2[1928]<=twadabc;necf6c2[1926]<=jp5fcdc[0];necf6c2[1809]<=qg6d5e2;necf6c2[1805]<=ie24fd0[0];necf6c2[1804]<=lqfe6e7[0];necf6c2[1803]<=ie3b7e7;necf6c2[1761]<=vvfc927;necf6c2[1748]<=kfae5ec[0];necf6c2[1727]<=xl22190;necf6c2[1696]<=babd901[0];necf6c2[1668]<=cm7d295[0];necf6c2[1571]<=yx6af11;necf6c2[1562]<=fp27e80;necf6c2[1560]<=thf373b[0];necf6c2[1558]<=sudbf39;necf6c2[1550]<=do93e46;necf6c2[1531]<=jr32183;necf6c2[1475]<=tue493f[0];necf6c2[1464]<=cz4bf24;necf6c2[1448]<=ww72f64[0];necf6c2[1406]<=sw10c86;necf6c2[1345]<=rtec80b[0];necf6c2[1288]<=vve94a8[0];necf6c2[1287]<=tw202f7[0];necf6c2[1242]<=xjc2572[0];necf6c2[1131]<=ou8d622;necf6c2[1094]<=jc5788d;necf6c2[1076]<=je3f407;necf6c2[1072]<=bn9b9df[0];necf6c2[1069]<=fadf9c9;necf6c2[1056]<=jc52a3f;necf6c2[1055]<=hqbdda[0];necf6c2[1052]<=mt9f233;necf6c2[1028]<=psfba93[0];necf6c2[1023]<=ofc3555[0];necf6c2[1014]<=yz90c1f;necf6c2[994]<=ldd2b6a;necf6c2[902]<=mg249fa[0];necf6c2[901]<=hbc76fc;necf6c2[880]<=xj5f924;necf6c2[874]<=an95cbd[0];necf6c2[863]<=wwc4432;necf6c2[848]<=sw97b20[0];necf6c2[834]<=uv6fa52[0];necf6c2[775]<=jpd27c8;necf6c2[765]<=xy86430;necf6c2[732]<=gbc97e4;necf6c2[643]<=dz6405e[0];necf6c2[621]<=zmb84ae[0];necf6c2[565]<=ri11ac4;necf6c2[528]<=nr4a547[0];necf6c2[527]<=ri17bb[0];necf6c2[514]<=ba3f752[0];necf6c2[497]<=tuda56d;necf6c2[450]<=mt18edf;necf6c2[437]<=ir12b97[0];necf6c2[431]<=lq58886;necf6c2[417]<=doadf4a[0];necf6c2[387]<=ym3bfe4;necf6c2[366]<=kf392fc;necf6c2[310]<=pfd7095[0];necf6c2[282]<=ale2358;necf6c2[257]<=ne47eea[0];necf6c2[248]<=irbb4ad;necf6c2[225]<=en75290;necf6c2[215]<=pf6b110;necf6c2[208]<=jcd5be9[0];necf6c2[193]<=ofe77fc;necf6c2[183]<=mre725f;necf6c2[155]<=gd9ae12[0];necf6c2[141]<=gqbc46b;necf6c2[128]<=zma8fdd;necf6c2[124]<=uvf7695;necf6c2[112]<=qgcea52;necf6c2[104]<=ayfa03b;necf6c2[96]<=aldceff;necf6c2[91]<=hbfce4b;necf6c2[77]<=tw935c2[0];necf6c2[64]<=ir951fb;necf6c2[62]<=kd5eed2[0];necf6c2[56]<=hq99d4a;necf6c2[38]<=lq526b8[0];necf6c2[19]<=cmea4d7[0];necf6c2[9]<=vvdd49a[0];end         assign suff972 = necf6c2,ld7b613 = cme5c87;   initial begin   jcc030e = $fopen(".fred");   $fdisplay( jcc030e, "%3h\n%3h", (thc27c7 >> 4) & fnc7fe5, (thc27c7 >> (mt9f1ff+4)) & fnc7fe5 );   $fclose(jcc030e);   $readmemh(".fred", qg721c0);   end   always @ (suff972) begin   ym8700c = qg721c0[1];       for (vk1872=0; vk1872<qgdb09f; vk1872=vk1872+1) begin           cme5c87[vk1872] = suff972[ym8700c];       rv38061  = ^(ym8700c & qg721c0[0]);       ym8700c =  {ym8700c, rv38061};       end   end
endmodule