module or1200_monitor2;
	wire [31:0] r0;
	wire [31:0] r1;
	wire [31:0] r2;
	wire [31:0] r3;
	wire [31:0] r4;
	wire [31:0] r5;
	wire [31:0] r6;
	wire [31:0] r7;
	wire [31:0] r8;
	wire [31:0] r9;
	wire [31:0] r10;
	wire [31:0] r11;
	wire [31:0] r12;
	wire [31:0] r13;
	wire [31:0] r14;
	wire [31:0] r15;
	wire [31:0] r16;
	wire [31:0] r17;
	wire [31:0] r18;
	wire [31:0] r19;
	wire [31:0] r20;
	wire [31:0] r21;
	wire [31:0] r22;
	wire [31:0] r23;
	wire [31:0] r24;
	wire [31:0] r25;
	wire [31:0] r26;
	wire [31:0] r27;
	wire [31:0] r28;
	wire [31:0] r29;
	wire [31:0] r30;
	wire [31:0] r31;
	assign r0 = `OR1200_TOP.or1200_cpu.or1200_rf.rf_a.mem[32*0+31:32*0];
	assign r1 = `OR1200_TOP.or1200_cpu.or1200_rf.rf_a.mem[32*1+31:32*1];
	assign r2 = `OR1200_TOP.or1200_cpu.or1200_rf.rf_a.mem[32*2+31:32*2];
	assign r3 = `OR1200_TOP.or1200_cpu.or1200_rf.rf_a.mem[32*3+31:32*3];
	assign r4 = `OR1200_TOP.or1200_cpu.or1200_rf.rf_a.mem[32*4+31:32*4];
	assign r5 = `OR1200_TOP.or1200_cpu.or1200_rf.rf_a.mem[32*5+31:32*5];
	assign r6 = `OR1200_TOP.or1200_cpu.or1200_rf.rf_a.mem[32*6+31:32*6];
	assign r7 = `OR1200_TOP.or1200_cpu.or1200_rf.rf_a.mem[32*7+31:32*7];
	assign r8 = `OR1200_TOP.or1200_cpu.or1200_rf.rf_a.mem[32*8+31:32*8];
	assign r9 = `OR1200_TOP.or1200_cpu.or1200_rf.rf_a.mem[32*9+31:32*9];
	assign r10 = `OR1200_TOP.or1200_cpu.or1200_rf.rf_a.mem[32*10+31:32*10];
	assign r11 = `OR1200_TOP.or1200_cpu.or1200_rf.rf_a.mem[32*11+31:32*11];
	assign r12 = `OR1200_TOP.or1200_cpu.or1200_rf.rf_a.mem[32*12+31:32*12];
	assign r13 = `OR1200_TOP.or1200_cpu.or1200_rf.rf_a.mem[32*13+31:32*13];
	assign r14 = `OR1200_TOP.or1200_cpu.or1200_rf.rf_a.mem[32*14+31:32*14];
	assign r15 = `OR1200_TOP.or1200_cpu.or1200_rf.rf_a.mem[32*15+31:32*15];
	assign r16 = `OR1200_TOP.or1200_cpu.or1200_rf.rf_a.mem[32*16+31:32*16];
	assign r17 = `OR1200_TOP.or1200_cpu.or1200_rf.rf_a.mem[32*17+31:32*17];
	assign r18 = `OR1200_TOP.or1200_cpu.or1200_rf.rf_a.mem[32*18+31:32*18];
	assign r19 = `OR1200_TOP.or1200_cpu.or1200_rf.rf_a.mem[32*19+31:32*19];
	assign r20 = `OR1200_TOP.or1200_cpu.or1200_rf.rf_a.mem[32*20+31:32*20];
	assign r21 = `OR1200_TOP.or1200_cpu.or1200_rf.rf_a.mem[32*21+31:32*21];
	assign r22 = `OR1200_TOP.or1200_cpu.or1200_rf.rf_a.mem[32*22+31:32*22];
	assign r23 = `OR1200_TOP.or1200_cpu.or1200_rf.rf_a.mem[32*23+31:32*23];
	assign r24 = `OR1200_TOP.or1200_cpu.or1200_rf.rf_a.mem[32*24+31:32*24];
	assign r25 = `OR1200_TOP.or1200_cpu.or1200_rf.rf_a.mem[32*25+31:32*25];
	assign r26 = `OR1200_TOP.or1200_cpu.or1200_rf.rf_a.mem[32*26+31:32*26];
	assign r27 = `OR1200_TOP.or1200_cpu.or1200_rf.rf_a.mem[32*27+31:32*27];
	assign r28 = `OR1200_TOP.or1200_cpu.or1200_rf.rf_a.mem[32*28+31:32*28];
	assign r29 = `OR1200_TOP.or1200_cpu.or1200_rf.rf_a.mem[32*29+31:32*29];
	assign r30 = `OR1200_TOP.or1200_cpu.or1200_rf.rf_a.mem[32*30+31:32*30];
	assign r31 = `OR1200_TOP.or1200_cpu.or1200_rf.rf_a.mem[32*31+31:32*31];
endmodule