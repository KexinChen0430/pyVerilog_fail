module SCB_P4_v1_20_0 (
    sclk,
    interrupt,
    clock);
    output      sclk;
    output      interrupt;
    input       clock;
          wire  Net_427;
          wire  Net_416;
          wire  Net_245;
          wire  Net_676;
          wire  Net_452;
          wire  Net_459;
          wire  Net_496;
          wire  Net_660;
          wire  Net_656;
          wire  Net_687;
          wire  Net_703;
          wire  Net_682;
          wire  Net_422;
          wire  Net_379;
          wire  Net_555;
          wire  Net_387;
          wire  uncfg_rx_irq;
          wire  Net_458;
          wire  Net_596;
          wire  Net_252;
          wire  Net_547;
          wire  rx_irq;
          wire [3:0] ss;
          wire  Net_467;
          wire  Net_655;
          wire  Net_663;
          wire  Net_581;
          wire  Net_474;
          wire  Net_651;
          wire  Net_580;
          wire  Net_654;
          wire  Net_653;
          wire  Net_652;
          wire  Net_284;
	cy_clock_v1_0
		#(.id("38321056-ba6d-401c-98e7-a21e84ee201e/81fcee8a-3b8b-4be1-9a5f-a5e2e619a938"),
		  .source_clock_id(""),
		  .divisor(0),
		  .period("156250000"),
		  .is_direct(0),
		  .is_digital(0))
		SCBCLK
		 (.clock_out(Net_284));
    ZeroTerminal ZeroTerminal_5 (
        .z(Net_459));
	// select_s_VM (cy_virtualmux_v1_0)
	assign Net_652 = Net_459;
    ZeroTerminal ZeroTerminal_4 (
        .z(Net_452));
    ZeroTerminal ZeroTerminal_3 (
        .z(Net_676));
    ZeroTerminal ZeroTerminal_2 (
        .z(Net_245));
    ZeroTerminal ZeroTerminal_1 (
        .z(Net_416));
	// rx_VM (cy_virtualmux_v1_0)
	assign Net_654 = Net_452;
	// rx_wake_VM (cy_virtualmux_v1_0)
	assign Net_682 = uncfg_rx_irq;
	// clock_VM (cy_virtualmux_v1_0)
	assign Net_655 = Net_284;
	// sclk_s_VM (cy_virtualmux_v1_0)
	assign Net_653 = Net_416;
	// mosi_s_VM (cy_virtualmux_v1_0)
	assign Net_651 = Net_676;
	// miso_m_VM (cy_virtualmux_v1_0)
	assign Net_663 = Net_245;
	wire [0:0] tmpOE__sda_net;
	wire [0:0] tmpFB_0__sda_net;
	wire [0:0] tmpINTERRUPT_0__sda_net;
	electrical [0:0] tmpSIOVREF__sda_net;
	cy_psoc3_pins_v1_10
		#(.id("38321056-ba6d-401c-98e7-a21e84ee201e/5382e105-1382-4a2e-b9f4-3bb2feba71e0"),
		  .drive_mode(3'b100),
		  .ibuf_enabled(1'b1),
		  .init_dr_st(1'b1),
		  .input_clk_en(0),
		  .input_sync(1'b0),
		  .input_sync_mode(1'b0),
		  .intr_mode(2'b00),
		  .invert_in_clock(0),
		  .invert_in_clock_en(0),
		  .invert_in_reset(0),
		  .invert_out_clock(0),
		  .invert_out_clock_en(0),
		  .invert_out_reset(0),
		  .io_voltage(""),
		  .layout_mode("CONTIGUOUS"),
		  .oe_conn(1'b0),
		  .oe_reset(0),
		  .oe_sync(1'b0),
		  .output_clk_en(0),
		  .output_clock_mode(1'b0),
		  .output_conn(1'b0),
		  .output_mode(1'b0),
		  .output_reset(0),
		  .output_sync(1'b0),
		  .pa_in_clock(-1),
		  .pa_in_clock_en(-1),
		  .pa_in_reset(-1),
		  .pa_out_clock(-1),
		  .pa_out_clock_en(-1),
		  .pa_out_reset(-1),
		  .pin_aliases(""),
		  .pin_mode("B"),
		  .por_state(4),
		  .sio_group_cnt(0),
		  .sio_hyst(1'b0),
		  .sio_ibuf(""),
		  .sio_info(2'b00),
		  .sio_obuf(""),
		  .sio_refsel(""),
		  .sio_vtrip(""),
		  .slew_rate(1'b0),
		  .spanning(0),
		  .use_annotation(1'b0),
		  .vtrip(2'b00),
		  .width(1))
		sda
		 (.oe(tmpOE__sda_net),
		  .y({1'b0}),
		  .fb({tmpFB_0__sda_net[0:0]}),
		  .io({Net_581}),
		  .siovref(tmpSIOVREF__sda_net),
		  .interrupt({tmpINTERRUPT_0__sda_net[0:0]}),
		  .in_clock({1'b0}),
		  .in_clock_en({1'b1}),
		  .in_reset({1'b0}),
		  .out_clock({1'b0}),
		  .out_clock_en({1'b1}),
		  .out_reset({1'b0}));
	assign tmpOE__sda_net = (`CYDEV_CHIP_MEMBER_USED == `CYDEV_CHIP_MEMBER_3A && `CYDEV_CHIP_REVISION_USED < `CYDEV_CHIP_REVISION_3A_ES3) ? ~{1'b1} : {1'b1};
	wire [0:0] tmpOE__scl_net;
	wire [0:0] tmpFB_0__scl_net;
	wire [0:0] tmpINTERRUPT_0__scl_net;
	electrical [0:0] tmpSIOVREF__scl_net;
	cy_psoc3_pins_v1_10
		#(.id("38321056-ba6d-401c-98e7-a21e84ee201e/22863ebe-a37b-476f-b252-6e49a8c00b12"),
		  .drive_mode(3'b100),
		  .ibuf_enabled(1'b1),
		  .init_dr_st(1'b1),
		  .input_clk_en(0),
		  .input_sync(1'b0),
		  .input_sync_mode(1'b0),
		  .intr_mode(2'b00),
		  .invert_in_clock(0),
		  .invert_in_clock_en(0),
		  .invert_in_reset(0),
		  .invert_out_clock(0),
		  .invert_out_clock_en(0),
		  .invert_out_reset(0),
		  .io_voltage(""),
		  .layout_mode("CONTIGUOUS"),
		  .oe_conn(1'b0),
		  .oe_reset(0),
		  .oe_sync(1'b0),
		  .output_clk_en(0),
		  .output_clock_mode(1'b0),
		  .output_conn(1'b0),
		  .output_mode(1'b0),
		  .output_reset(0),
		  .output_sync(1'b0),
		  .pa_in_clock(-1),
		  .pa_in_clock_en(-1),
		  .pa_in_reset(-1),
		  .pa_out_clock(-1),
		  .pa_out_clock_en(-1),
		  .pa_out_reset(-1),
		  .pin_aliases(""),
		  .pin_mode("B"),
		  .por_state(4),
		  .sio_group_cnt(0),
		  .sio_hyst(1'b0),
		  .sio_ibuf(""),
		  .sio_info(2'b00),
		  .sio_obuf(""),
		  .sio_refsel(""),
		  .sio_vtrip(""),
		  .slew_rate(1'b0),
		  .spanning(0),
		  .use_annotation(1'b0),
		  .vtrip(2'b00),
		  .width(1))
		scl
		 (.oe(tmpOE__scl_net),
		  .y({1'b0}),
		  .fb({tmpFB_0__scl_net[0:0]}),
		  .io({Net_580}),
		  .siovref(tmpSIOVREF__scl_net),
		  .interrupt({tmpINTERRUPT_0__scl_net[0:0]}),
		  .in_clock({1'b0}),
		  .in_clock_en({1'b1}),
		  .in_reset({1'b0}),
		  .out_clock({1'b0}),
		  .out_clock_en({1'b1}),
		  .out_reset({1'b0}));
	assign tmpOE__scl_net = (`CYDEV_CHIP_MEMBER_USED == `CYDEV_CHIP_MEMBER_3A && `CYDEV_CHIP_REVISION_USED < `CYDEV_CHIP_REVISION_3A_ES3) ? ~{1'b1} : {1'b1};
    ZeroTerminal ZeroTerminal_7 (
        .z(Net_427));
    assign sclk = Net_284 | Net_427;
	cy_isr_v1_0
		#(.int_type(2'b10))
		SCB_IRQ
		 (.int_signal(interrupt));
    cy_m0s8_scb_v1_0 SCB (
        .rx(Net_654),
        .miso_m(Net_663),
        .clock(Net_655),
        .select_m(ss[3:0]),
        .sclk_m(Net_687),
        .mosi_s(Net_651),
        .select_s(Net_652),
        .sclk_s(Net_653),
        .mosi_m(Net_660),
        .scl(Net_580),
        .sda(Net_581),
        .tx(Net_656),
        .miso_s(Net_703),
        .interrupt(interrupt));
    defparam SCB.scb_mode = 0;
endmodule