module outputs
  wire [127 : 0] wmemiM_MData;
  wire [35 : 0] wmemiM_MAddr;
  wire [31 : 0] wci_s_0_SData,
		wci_s_1_SData,
		wci_s_2_SData,
		wci_s_3_SData,
		wci_s_4_SData,
		wci_s_5_SData,
		wci_s_6_SData,
		wci_s_7_SData,
		wmiM0_MData,
		wmiM0_MFlag,
		wmiM1_MData,
		wmiM1_MFlag,
		wsi_m_dac_MData;
  wire [15 : 0] wmemiM_MDataByteEn;
  wire [13 : 0] wmiM0_MAddr, wmiM1_MAddr;
  wire [11 : 0] wmemiM_MBurstLength,
		wmiM0_MBurstLength,
		wmiM1_MBurstLength,
		wsi_m_dac_MBurstLength;
  wire [7 : 0] wsi_m_dac_MReqInfo;
  wire [3 : 0] wmiM0_MDataByteEn, wmiM1_MDataByteEn, wsi_m_dac_MByteEn;
  wire [2 : 0] wmemiM_MCmd, wmiM0_MCmd, wmiM1_MCmd, wsi_m_dac_MCmd;
  wire [1 : 0] wci_s_0_SFlag,
	       wci_s_0_SResp,
	       wci_s_1_SFlag,
	       wci_s_1_SResp,
	       wci_s_2_SFlag,
	       wci_s_2_SResp,
	       wci_s_3_SFlag,
	       wci_s_3_SResp,
	       wci_s_4_SFlag,
	       wci_s_4_SResp,
	       wci_s_5_SFlag,
	       wci_s_5_SResp,
	       wci_s_6_SFlag,
	       wci_s_6_SResp,
	       wci_s_7_SFlag,
	       wci_s_7_SResp;
  wire wci_s_0_SThreadBusy,
       wci_s_1_SThreadBusy,
       wci_s_2_SThreadBusy,
       wci_s_3_SThreadBusy,
       wci_s_4_SThreadBusy,
       wci_s_5_SThreadBusy,
       wci_s_6_SThreadBusy,
       wci_s_7_SThreadBusy,
       wmemiM_MDataLast,
       wmemiM_MDataValid,
       wmemiM_MReqLast,
       wmemiM_MReset_n,
       wmiM0_MAddrSpace,
       wmiM0_MDataLast,
       wmiM0_MDataValid,
       wmiM0_MReqInfo,
       wmiM0_MReqLast,
       wmiM0_MReset_n,
       wmiM1_MAddrSpace,
       wmiM1_MDataLast,
       wmiM1_MDataValid,
       wmiM1_MReqInfo,
       wmiM1_MReqLast,
       wmiM1_MReset_n,
       wsi_m_dac_MBurstPrecise,
       wsi_m_dac_MReqLast,
       wsi_m_dac_MReset_n,
       wsi_s_adc_SReset_n,
       wsi_s_adc_SThreadBusy;
  // Instantiate the wip-compliant app
  ocpi_app #(.hasDebugLogic(hasDebugLogic)) app(
				      .wci0_MReset_n(RST_N_rst_2),
				      .wci1_MReset_n(RST_N_rst_3),
				      .wci2_MReset_n(RST_N_rst_4),
				      .wci_Clk(CLK),
				      .wci0_MAddr(wci_s_2_MAddr),
				      .wci0_MAddrSpace(wci_s_2_MAddrSpace),
				      .wci0_MByteEn(wci_s_2_MByteEn),
				      .wci0_MCmd(wci_s_2_MCmd),
				      .wci0_MData(wci_s_2_MData),
				      .wci0_MFlag(wci_s_2_MFlag),
				      .wci1_MAddr(wci_s_3_MAddr),
				      .wci1_MAddrSpace(wci_s_3_MAddrSpace),
				      .wci1_MByteEn(wci_s_3_MByteEn),
				      .wci1_MCmd(wci_s_3_MCmd),
				      .wci1_MData(wci_s_3_MData),
				      .wci1_MFlag(wci_s_3_MFlag),
				      .wci2_MAddr(wci_s_4_MAddr),
				      .wci2_MAddrSpace(wci_s_4_MAddrSpace),
				      .wci2_MByteEn(wci_s_4_MByteEn),
				      .wci2_MCmd(wci_s_4_MCmd),
				      .wci2_MData(wci_s_4_MData),
				      .wci2_MFlag(wci_s_4_MFlag),
`ifdef NOTHERE
				      .wmemi0_SData(wmemiM_SData),
				      .wmemi0_SResp(wmemiM_SResp),
`endif
				      .FC_SData(wmiM0_SData),
				      .FC_SFlag(wmiM0_SFlag),
				      .FC_SResp(wmiM0_SResp),
				      .FP_SData(wmiM1_SData),
				      .FP_SFlag(wmiM1_SFlag),
				      .FP_SResp(wmiM1_SResp),
`ifdef NOTHERE
				      .adc_MBurstLength(wsi_s_adc_MBurstLength),
				      .adc_MByteEn(wsi_s_adc_MByteEn),
				      .adc_MCmd(wsi_s_adc_MCmd),
				      .adc_MData(wsi_s_adc_MData),
				      .adc_MReqInfo(wsi_s_adc_MReqInfo),
`endif
				      .FC_SThreadBusy(wmiM0_SThreadBusy),
				      .FC_SDataThreadBusy(wmiM0_SDataThreadBusy),
				      .FC_SRespLast(wmiM0_SRespLast),
				      .FC_SReset_n(wmiM0_SReset_n),
				      .FP_SThreadBusy(wmiM1_SThreadBusy),
				      .FP_SDataThreadBusy(wmiM1_SDataThreadBusy),
				      .FP_SRespLast(wmiM1_SRespLast),
				      .FP_SReset_n(wmiM1_SReset_n),
`ifdef NOTHERE
				      .wmemi0_SRespLast(wmemiM_SRespLast),
				      .wmemi0_SCmdAccept(wmemiM_SCmdAccept),
				      .wmemi0_SDataAccept(wmemiM_SDataAccept),
				      .adc_MReqLast(wsi_s_adc_MReqLast),
				      .adc_MBurstPrecise(wsi_s_adc_MBurstPrecise),
				      .adc_MReset_n(wsi_s_adc_MReset_n),
				      .dac_SThreadBusy(wsi_m_dac_SThreadBusy),
				      .dac_SReset_n(wsi_m_dac_SReset_n),
`endif
				      .wci0_SResp(wci_s_2_SResp),
				      .wci0_SData(wci_s_2_SData),
				      .wci0_SThreadBusy(wci_s_2_SThreadBusy),
				      .wci0_SFlag(wci_s_2_SFlag),
				      .wci1_SResp(wci_s_3_SResp),
				      .wci1_SData(wci_s_3_SData),
				      .wci1_SThreadBusy(wci_s_3_SThreadBusy),
				      .wci1_SFlag(wci_s_3_SFlag),
				      .wci2_SResp(wci_s_4_SResp),
				      .wci2_SData(wci_s_4_SData),
				      .wci2_SThreadBusy(wci_s_4_SThreadBusy),
				      .wci2_SFlag(wci_s_4_SFlag),
				      .FC_MCmd(wmiM0_MCmd),
				      .FC_MReqLast(wmiM0_MReqLast),
				      .FC_MReqInfo(wmiM0_MReqInfo),
				      .FC_MAddrSpace(wmiM0_MAddrSpace),
				      .FC_MAddr(wmiM0_MAddr),
				      .FC_MBurstLength(wmiM0_MBurstLength),
				      .FC_MDataValid(wmiM0_MDataValid),
				      .FC_MDataLast(wmiM0_MDataLast),
				      .FC_MData(wmiM0_MData),
				      .FC_MDataByteEn(wmiM0_MDataByteEn),
				      .FC_MFlag(wmiM0_MFlag),
				      .FC_MReset_n(wmiM0_MReset_n),
				      .FP_MCmd(wmiM1_MCmd),
				      .FP_MReqLast(wmiM1_MReqLast),
				      .FP_MReqInfo(wmiM1_MReqInfo),
				      .FP_MAddrSpace(wmiM1_MAddrSpace),
				      .FP_MAddr(wmiM1_MAddr),
				      .FP_MBurstLength(wmiM1_MBurstLength),
				      .FP_MDataValid(wmiM1_MDataValid),
				      .FP_MDataLast(wmiM1_MDataLast),
				      .FP_MData(wmiM1_MData),
				      .FP_MDataByteEn(wmiM1_MDataByteEn),
				      .FP_MFlag(wmiM1_MFlag),
				      .FP_MReset_n(wmiM1_MReset_n)
`ifdef NOTTHERE
				      .wmemi0_MCmd(wmemiM_MCmd),
				      .wmemi0_MReqLast(wmemiM_MReqLast),
				      .wmemi0_MAddr(wmemiM_MAddr),
				      .wmemi0_MBurstLength(wmemiM_MBurstLength),
				      .wmemi0_MDataValid(wmemiM_MDataValid),
				      .wmemi0_MDataLast(wmemiM_MDataLast),
				      .wmemi0_MData(wmemiM_MData),
				      .wmemi0_MDataByteEn(wmemiM_MDataByteEn),
				      .wmemi0_MReset_n(wmemiM_MReset_n)
`endif
);
//				      .adc_SThreadBusy(wsi_s_adc_SThreadBusy),
//				      .adc_SReset_n(wsi_s_adc_SReset_n),
//				      .dac_MCmd(wsi_m_dac_MCmd),
//				      .dac_MReqLast(wsi_m_dac_MReqLast),
//				      .dac_MBurstPrecise(wsi_m_dac_MBurstPrecise),
//				      .dac_MBurstLength(wsi_m_dac_MBurstLength),
//				      .dac_MData(wsi_m_dac_MData),
//				      .dac_MByteEn(wsi_m_dac_MByteEn),
//				      .dac_MReqInfo(wsi_m_dac_MReqInfo),
//				      .dac_MReset_n(wsi_m_dac_MReset_n));
endmodule