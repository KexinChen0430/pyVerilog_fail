module reset logic
	module_reset <= (tens_digit == 4'h6);
end
endmodule