module emFile_v1_20_7 ;
          wire  Net_31;
          wire  Net_30;
          wire  Net_29;
          wire  Net_28;
          wire  Net_27;
          wire  Net_26;
          wire  Net_24;
          wire  Net_23;
          wire  Net_21;
          wire  Net_20;
          wire  Net_18;
          wire  Net_17;
          wire  Net_14;
          wire  Net_13;
          wire  Net_12;
          wire  Net_11;
          wire  Net_9;
          wire  Net_8;
          wire  Net_6;
          wire  Net_5;
          wire  Net_4;
          wire  Net_3;
          wire  Net_2;
          wire  Net_1;
          wire  Net_58;
          wire  Net_57;
          wire  Net_55;
          wire  Net_54;
          wire  Net_43;
          wire  Net_42;
          wire  Net_40;
          wire  Net_39;
          wire  Net_83;
          wire  Net_81;
          wire  Net_80;
          wire  Net_66;
          wire  Net_19;
          wire  Net_16;
          wire  Net_22;
          wire  Net_10;
    SPI_Master_v2_40_6 SPI0 (
        .mosi(Net_10),
        .sclk(Net_22),
        .ss(Net_1),
        .miso(Net_16),
        .clock(Net_19),
        .reset(Net_2),
        .rx_interrupt(Net_3),
        .sdat(Net_4),
        .tx_interrupt(Net_5));
    defparam SPI0.BidirectMode = 0;
    defparam SPI0.HighSpeedMode = 1;
    defparam SPI0.NumberOfDataBits = 8;
    defparam SPI0.ShiftDir = 0;
	wire [0:0] tmpOE__mosi0_net;
	wire [0:0] tmpFB_0__mosi0_net;
	wire [0:0] tmpIO_0__mosi0_net;
	wire [0:0] tmpINTERRUPT_0__mosi0_net;
	electrical [0:0] tmpSIOVREF__mosi0_net;
	cy_psoc3_pins_v1_10
		#(.id("62946763-63ac-47e7-8754-b206ba7765cc/ed092b9b-d398-4703-be89-cebf998501f6"),
		  .drive_mode(3'b110),
		  .ibuf_enabled(1'b1),
		  .init_dr_st(1'b0),
		  .input_clk_en(0),
		  .input_sync(1'b1),
		  .input_sync_mode(1'b0),
		  .intr_mode(2'b00),
		  .invert_in_clock(0),
		  .invert_in_clock_en(0),
		  .invert_in_reset(0),
		  .invert_out_clock(0),
		  .invert_out_clock_en(0),
		  .invert_out_reset(0),
		  .io_voltage(""),
		  .layout_mode("CONTIGUOUS"),
		  .oe_conn(1'b0),
		  .oe_reset(0),
		  .oe_sync(1'b0),
		  .output_clk_en(0),
		  .output_clock_mode(1'b0),
		  .output_conn(1'b1),
		  .output_mode(1'b0),
		  .output_reset(0),
		  .output_sync(1'b0),
		  .pa_in_clock(-1),
		  .pa_in_clock_en(-1),
		  .pa_in_reset(-1),
		  .pa_out_clock(-1),
		  .pa_out_clock_en(-1),
		  .pa_out_reset(-1),
		  .pin_aliases(""),
		  .pin_mode("O"),
		  .por_state(4),
		  .sio_group_cnt(0),
		  .sio_hyst(1'b0),
		  .sio_ibuf(""),
		  .sio_info(2'b00),
		  .sio_obuf(""),
		  .sio_refsel(""),
		  .sio_vtrip(""),
		  .slew_rate(1'b0),
		  .spanning(0),
		  .use_annotation(1'b0),
		  .vtrip(2'b10),
		  .width(1))
		mosi0
		 (.oe(tmpOE__mosi0_net),
		  .y({Net_10}),
		  .fb({tmpFB_0__mosi0_net[0:0]}),
		  .io({tmpIO_0__mosi0_net[0:0]}),
		  .siovref(tmpSIOVREF__mosi0_net),
		  .interrupt({tmpINTERRUPT_0__mosi0_net[0:0]}),
		  .in_clock({1'b0}),
		  .in_clock_en({1'b1}),
		  .in_reset({1'b0}),
		  .out_clock({1'b0}),
		  .out_clock_en({1'b1}),
		  .out_reset({1'b0}));
	assign tmpOE__mosi0_net = (`CYDEV_CHIP_MEMBER_USED == `CYDEV_CHIP_MEMBER_3A && `CYDEV_CHIP_REVISION_USED < `CYDEV_CHIP_REVISION_3A_ES3) ? ~{1'b1} : {1'b1};
	cy_clock_v1_0
		#(.id("62946763-63ac-47e7-8754-b206ba7765cc/5ed615c6-e1f0-40ed-8816-f906ef67d531"),
		  .source_clock_id("61737EF6-3B74-48f9-8B91-F7473A442AE7"),
		  .divisor(1),
		  .period("0"),
		  .is_direct(0),
		  .is_digital(1))
		Clock_1
		 (.clock_out(Net_19));
	wire [0:0] tmpOE__miso0_net;
	wire [0:0] tmpIO_0__miso0_net;
	wire [0:0] tmpINTERRUPT_0__miso0_net;
	electrical [0:0] tmpSIOVREF__miso0_net;
	cy_psoc3_pins_v1_10
		#(.id("62946763-63ac-47e7-8754-b206ba7765cc/1425177d-0d0e-4468-8bcc-e638e5509a9b"),
		  .drive_mode(3'b001),
		  .ibuf_enabled(1'b1),
		  .init_dr_st(1'b0),
		  .input_clk_en(0),
		  .input_sync(1'b0),
		  .input_sync_mode(1'b0),
		  .intr_mode(2'b00),
		  .invert_in_clock(0),
		  .invert_in_clock_en(0),
		  .invert_in_reset(0),
		  .invert_out_clock(0),
		  .invert_out_clock_en(0),
		  .invert_out_reset(0),
		  .io_voltage(""),
		  .layout_mode("CONTIGUOUS"),
		  .oe_conn(1'b0),
		  .oe_reset(0),
		  .oe_sync(1'b0),
		  .output_clk_en(0),
		  .output_clock_mode(1'b0),
		  .output_conn(1'b0),
		  .output_mode(1'b0),
		  .output_reset(0),
		  .output_sync(1'b0),
		  .pa_in_clock(-1),
		  .pa_in_clock_en(-1),
		  .pa_in_reset(-1),
		  .pa_out_clock(-1),
		  .pa_out_clock_en(-1),
		  .pa_out_reset(-1),
		  .pin_aliases(""),
		  .pin_mode("I"),
		  .por_state(4),
		  .sio_group_cnt(0),
		  .sio_hyst(1'b0),
		  .sio_ibuf(""),
		  .sio_info(2'b00),
		  .sio_obuf(""),
		  .sio_refsel(""),
		  .sio_vtrip(""),
		  .slew_rate(1'b0),
		  .spanning(0),
		  .use_annotation(1'b0),
		  .vtrip(2'b00),
		  .width(1))
		miso0
		 (.oe(tmpOE__miso0_net),
		  .y({1'b0}),
		  .fb({Net_16}),
		  .io({tmpIO_0__miso0_net[0:0]}),
		  .siovref(tmpSIOVREF__miso0_net),
		  .interrupt({tmpINTERRUPT_0__miso0_net[0:0]}),
		  .in_clock({1'b0}),
		  .in_clock_en({1'b1}),
		  .in_reset({1'b0}),
		  .out_clock({1'b0}),
		  .out_clock_en({1'b1}),
		  .out_reset({1'b0}));
	assign tmpOE__miso0_net = (`CYDEV_CHIP_MEMBER_USED == `CYDEV_CHIP_MEMBER_3A && `CYDEV_CHIP_REVISION_USED < `CYDEV_CHIP_REVISION_3A_ES3) ? ~{1'b1} : {1'b1};
    ZeroTerminal ZeroTerminal_1 (
        .z(Net_2));
	wire [0:0] tmpOE__sclk0_net;
	wire [0:0] tmpFB_0__sclk0_net;
	wire [0:0] tmpIO_0__sclk0_net;
	wire [0:0] tmpINTERRUPT_0__sclk0_net;
	electrical [0:0] tmpSIOVREF__sclk0_net;
	cy_psoc3_pins_v1_10
		#(.id("62946763-63ac-47e7-8754-b206ba7765cc/ae249072-87dc-41aa-9405-888517aefa28"),
		  .drive_mode(3'b110),
		  .ibuf_enabled(1'b1),
		  .init_dr_st(1'b0),
		  .input_clk_en(0),
		  .input_sync(1'b1),
		  .input_sync_mode(1'b0),
		  .intr_mode(2'b00),
		  .invert_in_clock(0),
		  .invert_in_clock_en(0),
		  .invert_in_reset(0),
		  .invert_out_clock(0),
		  .invert_out_clock_en(0),
		  .invert_out_reset(0),
		  .io_voltage(""),
		  .layout_mode("CONTIGUOUS"),
		  .oe_conn(1'b0),
		  .oe_reset(0),
		  .oe_sync(1'b0),
		  .output_clk_en(0),
		  .output_clock_mode(1'b0),
		  .output_conn(1'b1),
		  .output_mode(1'b0),
		  .output_reset(0),
		  .output_sync(1'b0),
		  .pa_in_clock(-1),
		  .pa_in_clock_en(-1),
		  .pa_in_reset(-1),
		  .pa_out_clock(-1),
		  .pa_out_clock_en(-1),
		  .pa_out_reset(-1),
		  .pin_aliases(""),
		  .pin_mode("O"),
		  .por_state(4),
		  .sio_group_cnt(0),
		  .sio_hyst(1'b0),
		  .sio_ibuf(""),
		  .sio_info(2'b00),
		  .sio_obuf(""),
		  .sio_refsel(""),
		  .sio_vtrip(""),
		  .slew_rate(1'b0),
		  .spanning(0),
		  .use_annotation(1'b0),
		  .vtrip(2'b10),
		  .width(1))
		sclk0
		 (.oe(tmpOE__sclk0_net),
		  .y({Net_22}),
		  .fb({tmpFB_0__sclk0_net[0:0]}),
		  .io({tmpIO_0__sclk0_net[0:0]}),
		  .siovref(tmpSIOVREF__sclk0_net),
		  .interrupt({tmpINTERRUPT_0__sclk0_net[0:0]}),
		  .in_clock({1'b0}),
		  .in_clock_en({1'b1}),
		  .in_reset({1'b0}),
		  .out_clock({1'b0}),
		  .out_clock_en({1'b1}),
		  .out_reset({1'b0}));
	assign tmpOE__sclk0_net = (`CYDEV_CHIP_MEMBER_USED == `CYDEV_CHIP_MEMBER_3A && `CYDEV_CHIP_REVISION_USED < `CYDEV_CHIP_REVISION_3A_ES3) ? ~{1'b1} : {1'b1};
	wire [0:0] tmpOE__SPI0_CS_net;
	wire [0:0] tmpFB_0__SPI0_CS_net;
	wire [0:0] tmpIO_0__SPI0_CS_net;
	wire [0:0] tmpINTERRUPT_0__SPI0_CS_net;
	electrical [0:0] tmpSIOVREF__SPI0_CS_net;
	cy_psoc3_pins_v1_10
		#(.id("62946763-63ac-47e7-8754-b206ba7765cc/6df85302-e45f-45fb-97de-4bdf3128e07b"),
		  .drive_mode(3'b110),
		  .ibuf_enabled(1'b1),
		  .init_dr_st(1'b0),
		  .input_clk_en(0),
		  .input_sync(1'b1),
		  .input_sync_mode(1'b0),
		  .intr_mode(2'b00),
		  .invert_in_clock(0),
		  .invert_in_clock_en(0),
		  .invert_in_reset(0),
		  .invert_out_clock(0),
		  .invert_out_clock_en(0),
		  .invert_out_reset(0),
		  .io_voltage(""),
		  .layout_mode("CONTIGUOUS"),
		  .oe_conn(1'b0),
		  .oe_reset(0),
		  .oe_sync(1'b0),
		  .output_clk_en(0),
		  .output_clock_mode(1'b0),
		  .output_conn(1'b0),
		  .output_mode(1'b0),
		  .output_reset(0),
		  .output_sync(1'b0),
		  .pa_in_clock(-1),
		  .pa_in_clock_en(-1),
		  .pa_in_reset(-1),
		  .pa_out_clock(-1),
		  .pa_out_clock_en(-1),
		  .pa_out_reset(-1),
		  .pin_aliases(""),
		  .pin_mode("O"),
		  .por_state(4),
		  .sio_group_cnt(0),
		  .sio_hyst(1'b0),
		  .sio_ibuf(""),
		  .sio_info(2'b00),
		  .sio_obuf(""),
		  .sio_refsel(""),
		  .sio_vtrip(""),
		  .slew_rate(1'b0),
		  .spanning(0),
		  .use_annotation(1'b0),
		  .vtrip(2'b10),
		  .width(1))
		SPI0_CS
		 (.oe(tmpOE__SPI0_CS_net),
		  .y({1'b0}),
		  .fb({tmpFB_0__SPI0_CS_net[0:0]}),
		  .io({tmpIO_0__SPI0_CS_net[0:0]}),
		  .siovref(tmpSIOVREF__SPI0_CS_net),
		  .interrupt({tmpINTERRUPT_0__SPI0_CS_net[0:0]}),
		  .in_clock({1'b0}),
		  .in_clock_en({1'b1}),
		  .in_reset({1'b0}),
		  .out_clock({1'b0}),
		  .out_clock_en({1'b1}),
		  .out_reset({1'b0}));
	assign tmpOE__SPI0_CS_net = (`CYDEV_CHIP_MEMBER_USED == `CYDEV_CHIP_MEMBER_3A && `CYDEV_CHIP_REVISION_USED < `CYDEV_CHIP_REVISION_3A_ES3) ? ~{1'b1} : {1'b1};
endmodule