module sky130_fd_sc_hs__a31o (
    //# {{data|Data Signals}}
    input  A1,
    input  A2,
    input  A3,
    input  B1,
    output X
);
    // Voltage supply signals
    supply1 VPWR;
    supply0 VGND;
endmodule