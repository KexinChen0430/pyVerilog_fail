module to generate a "tone".
// Port Map
//   clock : circuit synchronous clock
//   reset : circult reset
//   note  : digital signal for the note
//   nv    : note valid strobe
input clock;
input reset;
output signed [14:0] note;
reg signed [14:0] note;
output nv;
reg nv;
reg [13:0] noteidx = 0;
reg [10:0] sample_rate_cnt = 1;
always @(posedge clock, negedge reset) begin: M_MUSICBOX_RTL
    if (reset == 0) begin
        sample_rate_cnt <= 1;
        note <= 0;
        noteidx <= 0;
        nv <= 0;
    end
    else begin
        if ((sample_rate_cnt == 1042)) begin
            sample_rate_cnt <= 1;
            case (noteidx)
                0: note <= 0;
                1: note <= 5378;
                2: note <= 9626;
                3: note <= 11911;
                4: note <= 11910;
                5: note <= 9889;
                6: note <= 6627;
                7: note <= 3203;
                8: note <= 697;
                9: note <= (-101);
                10: note <= 1098;
                11: note <= 3995;
                12: note <= 7791;
                13: note <= 11395;
                14: note <= 13722;
                15: note <= 13985;
                16: note <= 11910;
                17: note <= 7815;
                18: note <= 2531;
                19: note <= (-2814);
                20: note <= (-7094);
                21: note <= (-9474);
                22: note <= (-9626);
                23: note <= (-7815);
                24: note <= (-4815);
                25: note <= (-1697);
                26: note <= 467;
                27: note <= 893;
                28: note <= (-697);
                29: note <= (-3995);
                30: note <= (-8192);
                31: note <= (-12187);
                32: note <= (-14886);
                33: note <= (-15491);
                34: note <= (-13722);
                35: note <= (-9889);
                36: note <= (-4815);
                37: note <= 377;
                38: note <= 4563;
                39: note <= 6910;
                40: note <= 7094;
                41: note <= 5378;
                42: note <= 2531;
                43: note <= (-377);
                44: note <= (-2279);
                45: note <= (-2399);
                46: note <= (-467);
                47: note <= 3203;
                48: note <= 7791;
                49: note <= 12187;
                50: note <= 15286;
                51: note <= 16283;
                52: note <= 14886;
                53: note <= 11395;
                54: note <= 6627;
                55: note <= 1697;
                56: note <= (-2279);
                57: note <= (-4473);
                58: note <= (-4563);
                59: note <= (-2814);
                60: note <= 0;
                61: note <= 2814;
                62: note <= 4563;
                63: note <= 4473;
                64: note <= 2279;
                65: note <= (-1697);
                66: note <= (-6627);
                67: note <= (-11395);
                68: note <= (-14886);
                69: note <= (-16283);
                70: note <= (-15286);
                71: note <= (-12187);
                72: note <= (-7791);
                73: note <= (-3203);
                74: note <= 467;
                75: note <= 2399;
                76: note <= 2279;
                77: note <= 377;
                78: note <= (-2531);
                79: note <= (-5378);
                80: note <= (-7094);
                81: note <= (-6910);
                82: note <= (-4563);
                83: note <= (-377);
                84: note <= 4815;
                85: note <= 9889;
                86: note <= 13722;
                87: note <= 15491;
                88: note <= 14886;
                89: note <= 12187;
                90: note <= 8192;
                91: note <= 3995;
                92: note <= 697;
                93: note <= (-893);
                94: note <= (-467);
                95: note <= 1697;
                96: note <= 4815;
                97: note <= 7815;
                98: note <= 9626;
                99: note <= 9474;
                100: note <= 7094;
                101: note <= 2814;
                102: note <= (-2531);
                103: note <= (-7815);
                104: note <= (-11910);
                105: note <= (-13985);
                106: note <= (-13722);
                107: note <= (-11395);
                108: note <= (-7791);
                109: note <= (-3995);
                110: note <= (-1098);
                111: note <= 101;
                112: note <= (-697);
                113: note <= (-3203);
                114: note <= (-6627);
                115: note <= (-9889);
                116: note <= (-11910);
                117: note <= (-11911);
                118: note <= (-9626);
                119: note <= (-5378);
                120: note <= 0;
                121: note <= 5378;
                122: note <= 9626;
                123: note <= 11911;
                124: note <= 11910;
                125: note <= 9889;
                126: note <= 6627;
                127: note <= 3203;
                128: note <= 697;
                129: note <= (-101);
                130: note <= 1098;
                131: note <= 3995;
                132: note <= 7791;
                133: note <= 11395;
                134: note <= 13722;
                135: note <= 13985;
                136: note <= 11910;
                137: note <= 7815;
                138: note <= 2531;
                139: note <= (-2814);
                140: note <= (-7094);
                141: note <= (-9474);
                142: note <= (-9626);
                143: note <= (-7815);
                144: note <= (-4815);
                145: note <= (-1697);
                146: note <= 467;
                147: note <= 893;
                148: note <= (-697);
                149: note <= (-3995);
                150: note <= (-8192);
                151: note <= (-12187);
                152: note <= (-14886);
                153: note <= (-15491);
                154: note <= (-13722);
                155: note <= (-9889);
                156: note <= (-4815);
                157: note <= 377;
                158: note <= 4563;
                159: note <= 6910;
                160: note <= 7094;
                161: note <= 5378;
                162: note <= 2531;
                163: note <= (-377);
                164: note <= (-2279);
                165: note <= (-2399);
                166: note <= (-467);
                167: note <= 3203;
                168: note <= 7791;
                169: note <= 12187;
                170: note <= 15286;
                171: note <= 16283;
                172: note <= 14886;
                173: note <= 11395;
                174: note <= 6627;
                175: note <= 1697;
                176: note <= (-2279);
                177: note <= (-4473);
                178: note <= (-4563);
                179: note <= (-2814);
                180: note <= 0;
                181: note <= 2814;
                182: note <= 4563;
                183: note <= 4473;
                184: note <= 2279;
                185: note <= (-1697);
                186: note <= (-6627);
                187: note <= (-11395);
                188: note <= (-14886);
                189: note <= (-16283);
                190: note <= (-15286);
                191: note <= (-12187);
                192: note <= (-7791);
                193: note <= (-3203);
                194: note <= 467;
                195: note <= 2399;
                196: note <= 2279;
                197: note <= 377;
                198: note <= (-2531);
                199: note <= (-5378);
                200: note <= (-7094);
                201: note <= (-6910);
                202: note <= (-4563);
                203: note <= (-377);
                204: note <= 4815;
                205: note <= 9889;
                206: note <= 13722;
                207: note <= 15491;
                208: note <= 14886;
                209: note <= 12187;
                210: note <= 8192;
                211: note <= 3995;
                212: note <= 697;
                213: note <= (-893);
                214: note <= (-467);
                215: note <= 1697;
                216: note <= 4815;
                217: note <= 7815;
                218: note <= 9626;
                219: note <= 9474;
                220: note <= 7094;
                221: note <= 2814;
                222: note <= (-2531);
                223: note <= (-7815);
                224: note <= (-11910);
                225: note <= (-13985);
                226: note <= (-13722);
                227: note <= (-11395);
                228: note <= (-7791);
                229: note <= (-3995);
                230: note <= (-1098);
                231: note <= 101;
                232: note <= (-697);
                233: note <= (-3203);
                234: note <= (-6627);
                235: note <= (-9889);
                236: note <= (-11910);
                237: note <= (-11911);
                238: note <= (-9626);
                239: note <= (-5378);
                240: note <= 0;
                241: note <= 5378;
                242: note <= 9626;
                243: note <= 11911;
                244: note <= 11910;
                245: note <= 9889;
                246: note <= 6627;
                247: note <= 3203;
                248: note <= 697;
                249: note <= (-101);
                250: note <= 1098;
                251: note <= 3995;
                252: note <= 7791;
                253: note <= 11395;
                254: note <= 13722;
                255: note <= 13985;
                256: note <= 11910;
                257: note <= 7815;
                258: note <= 2531;
                259: note <= (-2814);
                260: note <= (-7094);
                261: note <= (-9474);
                262: note <= (-9626);
                263: note <= (-7815);
                264: note <= (-4815);
                265: note <= (-1697);
                266: note <= 467;
                267: note <= 893;
                268: note <= (-697);
                269: note <= (-3995);
                270: note <= (-8192);
                271: note <= (-12187);
                272: note <= (-14886);
                273: note <= (-15491);
                274: note <= (-13722);
                275: note <= (-9889);
                276: note <= (-4815);
                277: note <= 377;
                278: note <= 4563;
                279: note <= 6910;
                280: note <= 7094;
                281: note <= 5378;
                282: note <= 2531;
                283: note <= (-377);
                284: note <= (-2279);
                285: note <= (-2399);
                286: note <= (-467);
                287: note <= 3203;
                288: note <= 7791;
                289: note <= 12187;
                290: note <= 15286;
                291: note <= 16283;
                292: note <= 14886;
                293: note <= 11395;
                294: note <= 6627;
                295: note <= 1697;
                296: note <= (-2279);
                297: note <= (-4473);
                298: note <= (-4563);
                299: note <= (-2814);
                300: note <= 0;
                301: note <= 2814;
                302: note <= 4563;
                303: note <= 4473;
                304: note <= 2279;
                305: note <= (-1697);
                306: note <= (-6627);
                307: note <= (-11395);
                308: note <= (-14886);
                309: note <= (-16283);
                310: note <= (-15286);
                311: note <= (-12187);
                312: note <= (-7791);
                313: note <= (-3203);
                314: note <= 467;
                315: note <= 2399;
                316: note <= 2279;
                317: note <= 377;
                318: note <= (-2531);
                319: note <= (-5378);
                320: note <= (-7094);
                321: note <= (-6910);
                322: note <= (-4563);
                323: note <= (-377);
                324: note <= 4815;
                325: note <= 9889;
                326: note <= 13722;
                327: note <= 15491;
                328: note <= 14886;
                329: note <= 12187;
                330: note <= 8192;
                331: note <= 3995;
                332: note <= 697;
                333: note <= (-893);
                334: note <= (-467);
                335: note <= 1697;
                336: note <= 4815;
                337: note <= 7815;
                338: note <= 9626;
                339: note <= 9474;
                340: note <= 7094;
                341: note <= 2814;
                342: note <= (-2531);
                343: note <= (-7815);
                344: note <= (-11910);
                345: note <= (-13985);
                346: note <= (-13722);
                347: note <= (-11395);
                348: note <= (-7791);
                349: note <= (-3995);
                350: note <= (-1098);
                351: note <= 101;
                352: note <= (-697);
                353: note <= (-3203);
                354: note <= (-6627);
                355: note <= (-9889);
                356: note <= (-11910);
                357: note <= (-11911);
                358: note <= (-9626);
                359: note <= (-5378);
                360: note <= 0;
                361: note <= 5378;
                362: note <= 9626;
                363: note <= 11911;
                364: note <= 11910;
                365: note <= 9889;
                366: note <= 6627;
                367: note <= 3203;
                368: note <= 697;
                369: note <= (-101);
                370: note <= 1098;
                371: note <= 3995;
                372: note <= 7791;
                373: note <= 11395;
                374: note <= 13722;
                375: note <= 13985;
                376: note <= 11910;
                377: note <= 7815;
                378: note <= 2531;
                379: note <= (-2814);
                380: note <= (-7094);
                381: note <= (-9474);
                382: note <= (-9626);
                383: note <= (-7815);
                384: note <= (-4815);
                385: note <= (-1697);
                386: note <= 467;
                387: note <= 893;
                388: note <= (-697);
                389: note <= (-3995);
                390: note <= (-8192);
                391: note <= (-12187);
                392: note <= (-14886);
                393: note <= (-15491);
                394: note <= (-13722);
                395: note <= (-9889);
                396: note <= (-4815);
                397: note <= 377;
                398: note <= 4563;
                399: note <= 6910;
                400: note <= 7094;
                401: note <= 5378;
                402: note <= 2531;
                403: note <= (-377);
                404: note <= (-2279);
                405: note <= (-2399);
                406: note <= (-467);
                407: note <= 3203;
                408: note <= 7791;
                409: note <= 12187;
                410: note <= 15286;
                411: note <= 16283;
                412: note <= 14886;
                413: note <= 11395;
                414: note <= 6627;
                415: note <= 1697;
                416: note <= (-2279);
                417: note <= (-4473);
                418: note <= (-4563);
                419: note <= (-2814);
                420: note <= 0;
                421: note <= 2814;
                422: note <= 4563;
                423: note <= 4473;
                424: note <= 2279;
                425: note <= (-1697);
                426: note <= (-6627);
                427: note <= (-11395);
                428: note <= (-14886);
                429: note <= (-16283);
                430: note <= (-15286);
                431: note <= (-12187);
                432: note <= (-7791);
                433: note <= (-3203);
                434: note <= 467;
                435: note <= 2399;
                436: note <= 2279;
                437: note <= 377;
                438: note <= (-2531);
                439: note <= (-5378);
                440: note <= (-7094);
                441: note <= (-6910);
                442: note <= (-4563);
                443: note <= (-377);
                444: note <= 4815;
                445: note <= 9889;
                446: note <= 13722;
                447: note <= 15491;
                448: note <= 14886;
                449: note <= 12187;
                450: note <= 8192;
                451: note <= 3995;
                452: note <= 697;
                453: note <= (-893);
                454: note <= (-467);
                455: note <= 1697;
                456: note <= 4815;
                457: note <= 7815;
                458: note <= 9626;
                459: note <= 9474;
                460: note <= 7094;
                461: note <= 2814;
                462: note <= (-2531);
                463: note <= (-7815);
                464: note <= (-11910);
                465: note <= (-13985);
                466: note <= (-13722);
                467: note <= (-11395);
                468: note <= (-7791);
                469: note <= (-3995);
                470: note <= (-1098);
                471: note <= 101;
                472: note <= (-697);
                473: note <= (-3203);
                474: note <= (-6627);
                475: note <= (-9889);
                476: note <= (-11910);
                477: note <= (-11911);
                478: note <= (-9626);
                479: note <= (-5378);
                480: note <= 0;
                481: note <= 5378;
                482: note <= 9626;
                483: note <= 11911;
                484: note <= 11910;
                485: note <= 9889;
                486: note <= 6627;
                487: note <= 3203;
                488: note <= 697;
                489: note <= (-101);
                490: note <= 1098;
                491: note <= 3995;
                492: note <= 7791;
                493: note <= 11395;
                494: note <= 13722;
                495: note <= 13985;
                496: note <= 11910;
                497: note <= 7815;
                498: note <= 2531;
                499: note <= (-2814);
                500: note <= (-7094);
                501: note <= (-9474);
                502: note <= (-9626);
                503: note <= (-7815);
                504: note <= (-4815);
                505: note <= (-1697);
                506: note <= 467;
                507: note <= 893;
                508: note <= (-697);
                509: note <= (-3995);
                510: note <= (-8192);
                511: note <= (-12187);
                512: note <= (-14886);
                513: note <= (-15491);
                514: note <= (-13722);
                515: note <= (-9889);
                516: note <= (-4815);
                517: note <= 377;
                518: note <= 4563;
                519: note <= 6910;
                520: note <= 7094;
                521: note <= 5378;
                522: note <= 2531;
                523: note <= (-377);
                524: note <= (-2279);
                525: note <= (-2399);
                526: note <= (-467);
                527: note <= 3203;
                528: note <= 7791;
                529: note <= 12187;
                530: note <= 15286;
                531: note <= 16283;
                532: note <= 14886;
                533: note <= 11395;
                534: note <= 6627;
                535: note <= 1697;
                536: note <= (-2279);
                537: note <= (-4473);
                538: note <= (-4563);
                539: note <= (-2814);
                540: note <= 0;
                541: note <= 2814;
                542: note <= 4563;
                543: note <= 4473;
                544: note <= 2279;
                545: note <= (-1697);
                546: note <= (-6627);
                547: note <= (-11395);
                548: note <= (-14886);
                549: note <= (-16283);
                550: note <= (-15286);
                551: note <= (-12187);
                552: note <= (-7791);
                553: note <= (-3203);
                554: note <= 467;
                555: note <= 2399;
                556: note <= 2279;
                557: note <= 377;
                558: note <= (-2531);
                559: note <= (-5378);
                560: note <= (-7094);
                561: note <= (-6910);
                562: note <= (-4563);
                563: note <= (-377);
                564: note <= 4815;
                565: note <= 9889;
                566: note <= 13722;
                567: note <= 15491;
                568: note <= 14886;
                569: note <= 12187;
                570: note <= 8192;
                571: note <= 3995;
                572: note <= 697;
                573: note <= (-893);
                574: note <= (-467);
                575: note <= 1697;
                576: note <= 4815;
                577: note <= 7815;
                578: note <= 9626;
                579: note <= 9474;
                580: note <= 7094;
                581: note <= 2814;
                582: note <= (-2531);
                583: note <= (-7815);
                584: note <= (-11910);
                585: note <= (-13985);
                586: note <= (-13722);
                587: note <= (-11395);
                588: note <= (-7791);
                589: note <= (-3995);
                590: note <= (-1098);
                591: note <= 101;
                592: note <= (-697);
                593: note <= (-3203);
                594: note <= (-6627);
                595: note <= (-9889);
                596: note <= (-11910);
                597: note <= (-11911);
                598: note <= (-9626);
                599: note <= (-5378);
                600: note <= 0;
                601: note <= 5378;
                602: note <= 9626;
                603: note <= 11911;
                604: note <= 11910;
                605: note <= 9889;
                606: note <= 6627;
                607: note <= 3203;
                608: note <= 697;
                609: note <= (-101);
                610: note <= 1098;
                611: note <= 3995;
                612: note <= 7791;
                613: note <= 11395;
                614: note <= 13722;
                615: note <= 13985;
                616: note <= 11910;
                617: note <= 7815;
                618: note <= 2531;
                619: note <= (-2814);
                620: note <= (-7094);
                621: note <= (-9474);
                622: note <= (-9626);
                623: note <= (-7815);
                624: note <= (-4815);
                625: note <= (-1697);
                626: note <= 467;
                627: note <= 893;
                628: note <= (-697);
                629: note <= (-3995);
                630: note <= (-8192);
                631: note <= (-12187);
                632: note <= (-14886);
                633: note <= (-15491);
                634: note <= (-13722);
                635: note <= (-9889);
                636: note <= (-4815);
                637: note <= 377;
                638: note <= 4563;
                639: note <= 6910;
                640: note <= 7094;
                641: note <= 5378;
                642: note <= 2531;
                643: note <= (-377);
                644: note <= (-2279);
                645: note <= (-2399);
                646: note <= (-467);
                647: note <= 3203;
                648: note <= 7791;
                649: note <= 12187;
                650: note <= 15286;
                651: note <= 16283;
                652: note <= 14886;
                653: note <= 11395;
                654: note <= 6627;
                655: note <= 1697;
                656: note <= (-2279);
                657: note <= (-4473);
                658: note <= (-4563);
                659: note <= (-2814);
                660: note <= 0;
                661: note <= 2814;
                662: note <= 4563;
                663: note <= 4473;
                664: note <= 2279;
                665: note <= (-1697);
                666: note <= (-6627);
                667: note <= (-11395);
                668: note <= (-14886);
                669: note <= (-16283);
                670: note <= (-15286);
                671: note <= (-12187);
                672: note <= (-7791);
                673: note <= (-3203);
                674: note <= 467;
                675: note <= 2399;
                676: note <= 2279;
                677: note <= 377;
                678: note <= (-2531);
                679: note <= (-5378);
                680: note <= (-7094);
                681: note <= (-6910);
                682: note <= (-4563);
                683: note <= (-377);
                684: note <= 4815;
                685: note <= 9889;
                686: note <= 13722;
                687: note <= 15491;
                688: note <= 14886;
                689: note <= 12187;
                690: note <= 8192;
                691: note <= 3995;
                692: note <= 697;
                693: note <= (-893);
                694: note <= (-467);
                695: note <= 1697;
                696: note <= 4815;
                697: note <= 7815;
                698: note <= 9626;
                699: note <= 9474;
                700: note <= 7094;
                701: note <= 2814;
                702: note <= (-2531);
                703: note <= (-7815);
                704: note <= (-11910);
                705: note <= (-13985);
                706: note <= (-13722);
                707: note <= (-11395);
                708: note <= (-7791);
                709: note <= (-3995);
                710: note <= (-1098);
                711: note <= 101;
                712: note <= (-697);
                713: note <= (-3203);
                714: note <= (-6627);
                715: note <= (-9889);
                716: note <= (-11910);
                717: note <= (-11911);
                718: note <= (-9626);
                719: note <= (-5378);
                720: note <= 0;
                721: note <= 5378;
                722: note <= 9626;
                723: note <= 11911;
                724: note <= 11910;
                725: note <= 9889;
                726: note <= 6627;
                727: note <= 3203;
                728: note <= 697;
                729: note <= (-101);
                730: note <= 1098;
                731: note <= 3995;
                732: note <= 7791;
                733: note <= 11395;
                734: note <= 13722;
                735: note <= 13985;
                736: note <= 11910;
                737: note <= 7815;
                738: note <= 2531;
                739: note <= (-2814);
                740: note <= (-7094);
                741: note <= (-9474);
                742: note <= (-9626);
                743: note <= (-7815);
                744: note <= (-4815);
                745: note <= (-1697);
                746: note <= 467;
                747: note <= 893;
                748: note <= (-697);
                749: note <= (-3995);
                750: note <= (-8192);
                751: note <= (-12187);
                752: note <= (-14886);
                753: note <= (-15491);
                754: note <= (-13722);
                755: note <= (-9889);
                756: note <= (-4815);
                757: note <= 377;
                758: note <= 4563;
                759: note <= 6910;
                760: note <= 7094;
                761: note <= 5378;
                762: note <= 2531;
                763: note <= (-377);
                764: note <= (-2279);
                765: note <= (-2399);
                766: note <= (-467);
                767: note <= 3203;
                768: note <= 7791;
                769: note <= 12187;
                770: note <= 15286;
                771: note <= 16283;
                772: note <= 14886;
                773: note <= 11395;
                774: note <= 6627;
                775: note <= 1697;
                776: note <= (-2279);
                777: note <= (-4473);
                778: note <= (-4563);
                779: note <= (-2814);
                780: note <= 0;
                781: note <= 2814;
                782: note <= 4563;
                783: note <= 4473;
                784: note <= 2279;
                785: note <= (-1697);
                786: note <= (-6627);
                787: note <= (-11395);
                788: note <= (-14886);
                789: note <= (-16283);
                790: note <= (-15286);
                791: note <= (-12187);
                792: note <= (-7791);
                793: note <= (-3203);
                794: note <= 467;
                795: note <= 2399;
                796: note <= 2279;
                797: note <= 377;
                798: note <= (-2531);
                799: note <= (-5378);
                800: note <= (-7094);
                801: note <= (-6910);
                802: note <= (-4563);
                803: note <= (-377);
                804: note <= 4815;
                805: note <= 9889;
                806: note <= 13722;
                807: note <= 15491;
                808: note <= 14886;
                809: note <= 12187;
                810: note <= 8192;
                811: note <= 3995;
                812: note <= 697;
                813: note <= (-893);
                814: note <= (-467);
                815: note <= 1697;
                816: note <= 4815;
                817: note <= 7815;
                818: note <= 9626;
                819: note <= 9474;
                820: note <= 7094;
                821: note <= 2814;
                822: note <= (-2531);
                823: note <= (-7815);
                824: note <= (-11910);
                825: note <= (-13985);
                826: note <= (-13722);
                827: note <= (-11395);
                828: note <= (-7791);
                829: note <= (-3995);
                830: note <= (-1098);
                831: note <= 101;
                832: note <= (-697);
                833: note <= (-3203);
                834: note <= (-6627);
                835: note <= (-9889);
                836: note <= (-11910);
                837: note <= (-11911);
                838: note <= (-9626);
                839: note <= (-5378);
                840: note <= 0;
                841: note <= 5378;
                842: note <= 9626;
                843: note <= 11911;
                844: note <= 11910;
                845: note <= 9889;
                846: note <= 6627;
                847: note <= 3203;
                848: note <= 697;
                849: note <= (-101);
                850: note <= 1098;
                851: note <= 3995;
                852: note <= 7791;
                853: note <= 11395;
                854: note <= 13722;
                855: note <= 13985;
                856: note <= 11910;
                857: note <= 7815;
                858: note <= 2531;
                859: note <= (-2814);
                860: note <= (-7094);
                861: note <= (-9474);
                862: note <= (-9626);
                863: note <= (-7815);
                864: note <= (-4815);
                865: note <= (-1697);
                866: note <= 467;
                867: note <= 893;
                868: note <= (-697);
                869: note <= (-3995);
                870: note <= (-8192);
                871: note <= (-12187);
                872: note <= (-14886);
                873: note <= (-15491);
                874: note <= (-13722);
                875: note <= (-9889);
                876: note <= (-4815);
                877: note <= 377;
                878: note <= 4563;
                879: note <= 6910;
                880: note <= 7094;
                881: note <= 5378;
                882: note <= 2531;
                883: note <= (-377);
                884: note <= (-2279);
                885: note <= (-2399);
                886: note <= (-467);
                887: note <= 3203;
                888: note <= 7791;
                889: note <= 12187;
                890: note <= 15286;
                891: note <= 16283;
                892: note <= 14886;
                893: note <= 11395;
                894: note <= 6627;
                895: note <= 1697;
                896: note <= (-2279);
                897: note <= (-4473);
                898: note <= (-4563);
                899: note <= (-2814);
                900: note <= 0;
                901: note <= 2814;
                902: note <= 4563;
                903: note <= 4473;
                904: note <= 2279;
                905: note <= (-1697);
                906: note <= (-6627);
                907: note <= (-11395);
                908: note <= (-14886);
                909: note <= (-16283);
                910: note <= (-15286);
                911: note <= (-12187);
                912: note <= (-7791);
                913: note <= (-3203);
                914: note <= 467;
                915: note <= 2399;
                916: note <= 2279;
                917: note <= 377;
                918: note <= (-2531);
                919: note <= (-5378);
                920: note <= (-7094);
                921: note <= (-6910);
                922: note <= (-4563);
                923: note <= (-377);
                924: note <= 4815;
                925: note <= 9889;
                926: note <= 13722;
                927: note <= 15491;
                928: note <= 14886;
                929: note <= 12187;
                930: note <= 8192;
                931: note <= 3995;
                932: note <= 697;
                933: note <= (-893);
                934: note <= (-467);
                935: note <= 1697;
                936: note <= 4815;
                937: note <= 7815;
                938: note <= 9626;
                939: note <= 9474;
                940: note <= 7094;
                941: note <= 2814;
                942: note <= (-2531);
                943: note <= (-7815);
                944: note <= (-11910);
                945: note <= (-13985);
                946: note <= (-13722);
                947: note <= (-11395);
                948: note <= (-7791);
                949: note <= (-3995);
                950: note <= (-1098);
                951: note <= 101;
                952: note <= (-697);
                953: note <= (-3203);
                954: note <= (-6627);
                955: note <= (-9889);
                956: note <= (-11910);
                957: note <= (-11911);
                958: note <= (-9626);
                959: note <= (-5378);
                960: note <= 0;
                961: note <= 5378;
                962: note <= 9626;
                963: note <= 11911;
                964: note <= 11910;
                965: note <= 9889;
                966: note <= 6627;
                967: note <= 3203;
                968: note <= 697;
                969: note <= (-101);
                970: note <= 1098;
                971: note <= 3995;
                972: note <= 7791;
                973: note <= 11395;
                974: note <= 13722;
                975: note <= 13985;
                976: note <= 11910;
                977: note <= 7815;
                978: note <= 2531;
                979: note <= (-2814);
                980: note <= (-7094);
                981: note <= (-9474);
                982: note <= (-9626);
                983: note <= (-7815);
                984: note <= (-4815);
                985: note <= (-1697);
                986: note <= 467;
                987: note <= 893;
                988: note <= (-697);
                989: note <= (-3995);
                990: note <= (-8192);
                991: note <= (-12187);
                992: note <= (-14886);
                993: note <= (-15491);
                994: note <= (-13722);
                995: note <= (-9889);
                996: note <= (-4815);
                997: note <= 377;
                998: note <= 4563;
                999: note <= 6910;
                1000: note <= 7094;
                1001: note <= 5378;
                1002: note <= 2531;
                1003: note <= (-377);
                1004: note <= (-2279);
                1005: note <= (-2399);
                1006: note <= (-467);
                1007: note <= 3203;
                1008: note <= 7791;
                1009: note <= 12187;
                1010: note <= 15286;
                1011: note <= 16283;
                1012: note <= 14886;
                1013: note <= 11395;
                1014: note <= 6627;
                1015: note <= 1697;
                1016: note <= (-2279);
                1017: note <= (-4473);
                1018: note <= (-4563);
                1019: note <= (-2814);
                1020: note <= 0;
                1021: note <= 2814;
                1022: note <= 4563;
                1023: note <= 4473;
                1024: note <= 2279;
                1025: note <= (-1697);
                1026: note <= (-6627);
                1027: note <= (-11395);
                1028: note <= (-14886);
                1029: note <= (-16283);
                1030: note <= (-15286);
                1031: note <= (-12187);
                1032: note <= (-7791);
                1033: note <= (-3203);
                1034: note <= 467;
                1035: note <= 2399;
                1036: note <= 2279;
                1037: note <= 377;
                1038: note <= (-2531);
                1039: note <= (-5378);
                1040: note <= (-7094);
                1041: note <= (-6910);
                1042: note <= (-4563);
                1043: note <= (-377);
                1044: note <= 4815;
                1045: note <= 9889;
                1046: note <= 13722;
                1047: note <= 15491;
                1048: note <= 14886;
                1049: note <= 12187;
                1050: note <= 8192;
                1051: note <= 3995;
                1052: note <= 697;
                1053: note <= (-893);
                1054: note <= (-467);
                1055: note <= 1697;
                1056: note <= 4815;
                1057: note <= 7815;
                1058: note <= 9626;
                1059: note <= 9474;
                1060: note <= 7094;
                1061: note <= 2814;
                1062: note <= (-2531);
                1063: note <= (-7815);
                1064: note <= (-11910);
                1065: note <= (-13985);
                1066: note <= (-13722);
                1067: note <= (-11395);
                1068: note <= (-7791);
                1069: note <= (-3995);
                1070: note <= (-1098);
                1071: note <= 101;
                1072: note <= (-697);
                1073: note <= (-3203);
                1074: note <= (-6627);
                1075: note <= (-9889);
                1076: note <= (-11910);
                1077: note <= (-11911);
                1078: note <= (-9626);
                1079: note <= (-5378);
                1080: note <= 0;
                1081: note <= 5378;
                1082: note <= 9626;
                1083: note <= 11911;
                1084: note <= 11910;
                1085: note <= 9889;
                1086: note <= 6627;
                1087: note <= 3203;
                1088: note <= 697;
                1089: note <= (-101);
                1090: note <= 1098;
                1091: note <= 3995;
                1092: note <= 7791;
                1093: note <= 11395;
                1094: note <= 13722;
                1095: note <= 13985;
                1096: note <= 11910;
                1097: note <= 7815;
                1098: note <= 2531;
                1099: note <= (-2814);
                1100: note <= (-7094);
                1101: note <= (-9474);
                1102: note <= (-9626);
                1103: note <= (-7815);
                1104: note <= (-4815);
                1105: note <= (-1697);
                1106: note <= 467;
                1107: note <= 893;
                1108: note <= (-697);
                1109: note <= (-3995);
                1110: note <= (-8192);
                1111: note <= (-12187);
                1112: note <= (-14886);
                1113: note <= (-15491);
                1114: note <= (-13722);
                1115: note <= (-9889);
                1116: note <= (-4815);
                1117: note <= 377;
                1118: note <= 4563;
                1119: note <= 6910;
                1120: note <= 7094;
                1121: note <= 5378;
                1122: note <= 2531;
                1123: note <= (-377);
                1124: note <= (-2279);
                1125: note <= (-2399);
                1126: note <= (-467);
                1127: note <= 3203;
                1128: note <= 7791;
                1129: note <= 12187;
                1130: note <= 15286;
                1131: note <= 16283;
                1132: note <= 14886;
                1133: note <= 11395;
                1134: note <= 6627;
                1135: note <= 1697;
                1136: note <= (-2279);
                1137: note <= (-4473);
                1138: note <= (-4563);
                1139: note <= (-2814);
                1140: note <= 0;
                1141: note <= 2814;
                1142: note <= 4563;
                1143: note <= 4473;
                1144: note <= 2279;
                1145: note <= (-1697);
                1146: note <= (-6627);
                1147: note <= (-11395);
                1148: note <= (-14886);
                1149: note <= (-16283);
                1150: note <= (-15286);
                1151: note <= (-12187);
                1152: note <= (-7791);
                1153: note <= (-3203);
                1154: note <= 467;
                1155: note <= 2399;
                1156: note <= 2279;
                1157: note <= 377;
                1158: note <= (-2531);
                1159: note <= (-5378);
                1160: note <= (-7094);
                1161: note <= (-6910);
                1162: note <= (-4563);
                1163: note <= (-377);
                1164: note <= 4815;
                1165: note <= 9889;
                1166: note <= 13722;
                1167: note <= 15491;
                1168: note <= 14886;
                1169: note <= 12187;
                1170: note <= 8192;
                1171: note <= 3995;
                1172: note <= 697;
                1173: note <= (-893);
                1174: note <= (-467);
                1175: note <= 1697;
                1176: note <= 4815;
                1177: note <= 7815;
                1178: note <= 9626;
                1179: note <= 9474;
                1180: note <= 7094;
                1181: note <= 2814;
                1182: note <= (-2531);
                1183: note <= (-7815);
                1184: note <= (-11910);
                1185: note <= (-13985);
                1186: note <= (-13722);
                1187: note <= (-11395);
                1188: note <= (-7791);
                1189: note <= (-3995);
                1190: note <= (-1098);
                1191: note <= 101;
                1192: note <= (-697);
                1193: note <= (-3203);
                1194: note <= (-6627);
                1195: note <= (-9889);
                1196: note <= (-11910);
                1197: note <= (-11911);
                1198: note <= (-9626);
                1199: note <= (-5378);
                1200: note <= 0;
                1201: note <= 5378;
                1202: note <= 9626;
                1203: note <= 11911;
                1204: note <= 11910;
                1205: note <= 9889;
                1206: note <= 6627;
                1207: note <= 3203;
                1208: note <= 697;
                1209: note <= (-101);
                1210: note <= 1098;
                1211: note <= 3995;
                1212: note <= 7791;
                1213: note <= 11395;
                1214: note <= 13722;
                1215: note <= 13985;
                1216: note <= 11910;
                1217: note <= 7815;
                1218: note <= 2531;
                1219: note <= (-2814);
                1220: note <= (-7094);
                1221: note <= (-9474);
                1222: note <= (-9626);
                1223: note <= (-7815);
                1224: note <= (-4815);
                1225: note <= (-1697);
                1226: note <= 467;
                1227: note <= 893;
                1228: note <= (-697);
                1229: note <= (-3995);
                1230: note <= (-8192);
                1231: note <= (-12187);
                1232: note <= (-14886);
                1233: note <= (-15491);
                1234: note <= (-13722);
                1235: note <= (-9889);
                1236: note <= (-4815);
                1237: note <= 377;
                1238: note <= 4563;
                1239: note <= 6910;
                1240: note <= 7094;
                1241: note <= 5378;
                1242: note <= 2531;
                1243: note <= (-377);
                1244: note <= (-2279);
                1245: note <= (-2399);
                1246: note <= (-467);
                1247: note <= 3203;
                1248: note <= 7791;
                1249: note <= 12187;
                1250: note <= 15286;
                1251: note <= 16283;
                1252: note <= 14886;
                1253: note <= 11395;
                1254: note <= 6627;
                1255: note <= 1697;
                1256: note <= (-2279);
                1257: note <= (-4473);
                1258: note <= (-4563);
                1259: note <= (-2814);
                1260: note <= 0;
                1261: note <= 2814;
                1262: note <= 4563;
                1263: note <= 4473;
                1264: note <= 2279;
                1265: note <= (-1697);
                1266: note <= (-6627);
                1267: note <= (-11395);
                1268: note <= (-14886);
                1269: note <= (-16283);
                1270: note <= (-15286);
                1271: note <= (-12187);
                1272: note <= (-7791);
                1273: note <= (-3203);
                1274: note <= 467;
                1275: note <= 2399;
                1276: note <= 2279;
                1277: note <= 377;
                1278: note <= (-2531);
                1279: note <= (-5378);
                1280: note <= (-7094);
                1281: note <= (-6910);
                1282: note <= (-4563);
                1283: note <= (-377);
                1284: note <= 4815;
                1285: note <= 9889;
                1286: note <= 13722;
                1287: note <= 15491;
                1288: note <= 14886;
                1289: note <= 12187;
                1290: note <= 8192;
                1291: note <= 3995;
                1292: note <= 697;
                1293: note <= (-893);
                1294: note <= (-467);
                1295: note <= 1697;
                1296: note <= 4815;
                1297: note <= 7815;
                1298: note <= 9626;
                1299: note <= 9474;
                1300: note <= 7094;
                1301: note <= 2814;
                1302: note <= (-2531);
                1303: note <= (-7815);
                1304: note <= (-11910);
                1305: note <= (-13985);
                1306: note <= (-13722);
                1307: note <= (-11395);
                1308: note <= (-7791);
                1309: note <= (-3995);
                1310: note <= (-1098);
                1311: note <= 101;
                1312: note <= (-697);
                1313: note <= (-3203);
                1314: note <= (-6627);
                1315: note <= (-9889);
                1316: note <= (-11910);
                1317: note <= (-11911);
                1318: note <= (-9626);
                1319: note <= (-5378);
                1320: note <= 0;
                1321: note <= 5378;
                1322: note <= 9626;
                1323: note <= 11911;
                1324: note <= 11910;
                1325: note <= 9889;
                1326: note <= 6627;
                1327: note <= 3203;
                1328: note <= 697;
                1329: note <= (-101);
                1330: note <= 1098;
                1331: note <= 3995;
                1332: note <= 7791;
                1333: note <= 11395;
                1334: note <= 13722;
                1335: note <= 13985;
                1336: note <= 11910;
                1337: note <= 7815;
                1338: note <= 2531;
                1339: note <= (-2814);
                1340: note <= (-7094);
                1341: note <= (-9474);
                1342: note <= (-9626);
                1343: note <= (-7815);
                1344: note <= (-4815);
                1345: note <= (-1697);
                1346: note <= 467;
                1347: note <= 893;
                1348: note <= (-697);
                1349: note <= (-3995);
                1350: note <= (-8192);
                1351: note <= (-12187);
                1352: note <= (-14886);
                1353: note <= (-15491);
                1354: note <= (-13722);
                1355: note <= (-9889);
                1356: note <= (-4815);
                1357: note <= 377;
                1358: note <= 4563;
                1359: note <= 6910;
                1360: note <= 7094;
                1361: note <= 5378;
                1362: note <= 2531;
                1363: note <= (-377);
                1364: note <= (-2279);
                1365: note <= (-2399);
                1366: note <= (-467);
                1367: note <= 3203;
                1368: note <= 7791;
                1369: note <= 12187;
                1370: note <= 15286;
                1371: note <= 16283;
                1372: note <= 14886;
                1373: note <= 11395;
                1374: note <= 6627;
                1375: note <= 1697;
                1376: note <= (-2279);
                1377: note <= (-4473);
                1378: note <= (-4563);
                1379: note <= (-2814);
                1380: note <= 0;
                1381: note <= 2814;
                1382: note <= 4563;
                1383: note <= 4473;
                1384: note <= 2279;
                1385: note <= (-1697);
                1386: note <= (-6627);
                1387: note <= (-11395);
                1388: note <= (-14886);
                1389: note <= (-16283);
                1390: note <= (-15286);
                1391: note <= (-12187);
                1392: note <= (-7791);
                1393: note <= (-3203);
                1394: note <= 467;
                1395: note <= 2399;
                1396: note <= 2279;
                1397: note <= 377;
                1398: note <= (-2531);
                1399: note <= (-5378);
                1400: note <= (-7094);
                1401: note <= (-6910);
                1402: note <= (-4563);
                1403: note <= (-377);
                1404: note <= 4815;
                1405: note <= 9889;
                1406: note <= 13722;
                1407: note <= 15491;
                1408: note <= 14886;
                1409: note <= 12187;
                1410: note <= 8192;
                1411: note <= 3995;
                1412: note <= 697;
                1413: note <= (-893);
                1414: note <= (-467);
                1415: note <= 1697;
                1416: note <= 4815;
                1417: note <= 7815;
                1418: note <= 9626;
                1419: note <= 9474;
                1420: note <= 7094;
                1421: note <= 2814;
                1422: note <= (-2531);
                1423: note <= (-7815);
                1424: note <= (-11910);
                1425: note <= (-13985);
                1426: note <= (-13722);
                1427: note <= (-11395);
                1428: note <= (-7791);
                1429: note <= (-3995);
                1430: note <= (-1098);
                1431: note <= 101;
                1432: note <= (-697);
                1433: note <= (-3203);
                1434: note <= (-6627);
                1435: note <= (-9889);
                1436: note <= (-11910);
                1437: note <= (-11911);
                1438: note <= (-9626);
                1439: note <= (-5378);
                1440: note <= 0;
                1441: note <= 5378;
                1442: note <= 9626;
                1443: note <= 11911;
                1444: note <= 11910;
                1445: note <= 9889;
                1446: note <= 6627;
                1447: note <= 3203;
                1448: note <= 697;
                1449: note <= (-101);
                1450: note <= 1098;
                1451: note <= 3995;
                1452: note <= 7791;
                1453: note <= 11395;
                1454: note <= 13722;
                1455: note <= 13985;
                1456: note <= 11910;
                1457: note <= 7815;
                1458: note <= 2531;
                1459: note <= (-2814);
                1460: note <= (-7094);
                1461: note <= (-9474);
                1462: note <= (-9626);
                1463: note <= (-7815);
                1464: note <= (-4815);
                1465: note <= (-1697);
                1466: note <= 467;
                1467: note <= 893;
                1468: note <= (-697);
                1469: note <= (-3995);
                1470: note <= (-8192);
                1471: note <= (-12187);
                1472: note <= (-14886);
                1473: note <= (-15491);
                1474: note <= (-13722);
                1475: note <= (-9889);
                1476: note <= (-4815);
                1477: note <= 377;
                1478: note <= 4563;
                1479: note <= 6910;
                1480: note <= 7094;
                1481: note <= 5378;
                1482: note <= 2531;
                1483: note <= (-377);
                1484: note <= (-2279);
                1485: note <= (-2399);
                1486: note <= (-467);
                1487: note <= 3203;
                1488: note <= 7791;
                1489: note <= 12187;
                1490: note <= 15286;
                1491: note <= 16283;
                1492: note <= 14886;
                1493: note <= 11395;
                1494: note <= 6627;
                1495: note <= 1697;
                1496: note <= (-2279);
                1497: note <= (-4473);
                1498: note <= (-4563);
                1499: note <= (-2814);
                1500: note <= 0;
                1501: note <= 2814;
                1502: note <= 4563;
                1503: note <= 4473;
                1504: note <= 2279;
                1505: note <= (-1697);
                1506: note <= (-6627);
                1507: note <= (-11395);
                1508: note <= (-14886);
                1509: note <= (-16283);
                1510: note <= (-15286);
                1511: note <= (-12187);
                1512: note <= (-7791);
                1513: note <= (-3203);
                1514: note <= 467;
                1515: note <= 2399;
                1516: note <= 2279;
                1517: note <= 377;
                1518: note <= (-2531);
                1519: note <= (-5378);
                1520: note <= (-7094);
                1521: note <= (-6910);
                1522: note <= (-4563);
                1523: note <= (-377);
                1524: note <= 4815;
                1525: note <= 9889;
                1526: note <= 13722;
                1527: note <= 15491;
                1528: note <= 14886;
                1529: note <= 12187;
                1530: note <= 8192;
                1531: note <= 3995;
                1532: note <= 697;
                1533: note <= (-893);
                1534: note <= (-467);
                1535: note <= 1697;
                1536: note <= 4815;
                1537: note <= 7815;
                1538: note <= 9626;
                1539: note <= 9474;
                1540: note <= 7094;
                1541: note <= 2814;
                1542: note <= (-2531);
                1543: note <= (-7815);
                1544: note <= (-11910);
                1545: note <= (-13985);
                1546: note <= (-13722);
                1547: note <= (-11395);
                1548: note <= (-7791);
                1549: note <= (-3995);
                1550: note <= (-1098);
                1551: note <= 101;
                1552: note <= (-697);
                1553: note <= (-3203);
                1554: note <= (-6627);
                1555: note <= (-9889);
                1556: note <= (-11910);
                1557: note <= (-11911);
                1558: note <= (-9626);
                1559: note <= (-5378);
                1560: note <= 0;
                1561: note <= 5378;
                1562: note <= 9626;
                1563: note <= 11911;
                1564: note <= 11910;
                1565: note <= 9889;
                1566: note <= 6627;
                1567: note <= 3203;
                1568: note <= 697;
                1569: note <= (-101);
                1570: note <= 1098;
                1571: note <= 3995;
                1572: note <= 7791;
                1573: note <= 11395;
                1574: note <= 13722;
                1575: note <= 13985;
                1576: note <= 11910;
                1577: note <= 7815;
                1578: note <= 2531;
                1579: note <= (-2814);
                1580: note <= (-7094);
                1581: note <= (-9474);
                1582: note <= (-9626);
                1583: note <= (-7815);
                1584: note <= (-4815);
                1585: note <= (-1697);
                1586: note <= 467;
                1587: note <= 893;
                1588: note <= (-697);
                1589: note <= (-3995);
                1590: note <= (-8192);
                1591: note <= (-12187);
                1592: note <= (-14886);
                1593: note <= (-15491);
                1594: note <= (-13722);
                1595: note <= (-9889);
                1596: note <= (-4815);
                1597: note <= 377;
                1598: note <= 4563;
                1599: note <= 6910;
                1600: note <= 7094;
                1601: note <= 5378;
                1602: note <= 2531;
                1603: note <= (-377);
                1604: note <= (-2279);
                1605: note <= (-2399);
                1606: note <= (-467);
                1607: note <= 3203;
                1608: note <= 7791;
                1609: note <= 12187;
                1610: note <= 15286;
                1611: note <= 16283;
                1612: note <= 14886;
                1613: note <= 11395;
                1614: note <= 6627;
                1615: note <= 1697;
                1616: note <= (-2279);
                1617: note <= (-4473);
                1618: note <= (-4563);
                1619: note <= (-2814);
                1620: note <= 0;
                1621: note <= 2814;
                1622: note <= 4563;
                1623: note <= 4473;
                1624: note <= 2279;
                1625: note <= (-1697);
                1626: note <= (-6627);
                1627: note <= (-11395);
                1628: note <= (-14886);
                1629: note <= (-16283);
                1630: note <= (-15286);
                1631: note <= (-12187);
                1632: note <= (-7791);
                1633: note <= (-3203);
                1634: note <= 467;
                1635: note <= 2399;
                1636: note <= 2279;
                1637: note <= 377;
                1638: note <= (-2531);
                1639: note <= (-5378);
                1640: note <= (-7094);
                1641: note <= (-6910);
                1642: note <= (-4563);
                1643: note <= (-377);
                1644: note <= 4815;
                1645: note <= 9889;
                1646: note <= 13722;
                1647: note <= 15491;
                1648: note <= 14886;
                1649: note <= 12187;
                1650: note <= 8192;
                1651: note <= 3995;
                1652: note <= 697;
                1653: note <= (-893);
                1654: note <= (-467);
                1655: note <= 1697;
                1656: note <= 4815;
                1657: note <= 7815;
                1658: note <= 9626;
                1659: note <= 9474;
                1660: note <= 7094;
                1661: note <= 2814;
                1662: note <= (-2531);
                1663: note <= (-7815);
                1664: note <= (-11910);
                1665: note <= (-13985);
                1666: note <= (-13722);
                1667: note <= (-11395);
                1668: note <= (-7791);
                1669: note <= (-3995);
                1670: note <= (-1098);
                1671: note <= 101;
                1672: note <= (-697);
                1673: note <= (-3203);
                1674: note <= (-6627);
                1675: note <= (-9889);
                1676: note <= (-11910);
                1677: note <= (-11911);
                1678: note <= (-9626);
                1679: note <= (-5378);
                1680: note <= 0;
                1681: note <= 5378;
                1682: note <= 9626;
                1683: note <= 11911;
                1684: note <= 11910;
                1685: note <= 9889;
                1686: note <= 6627;
                1687: note <= 3203;
                1688: note <= 697;
                1689: note <= (-101);
                1690: note <= 1098;
                1691: note <= 3995;
                1692: note <= 7791;
                1693: note <= 11395;
                1694: note <= 13722;
                1695: note <= 13985;
                1696: note <= 11910;
                1697: note <= 7815;
                1698: note <= 2531;
                1699: note <= (-2814);
                1700: note <= (-7094);
                1701: note <= (-9474);
                1702: note <= (-9626);
                1703: note <= (-7815);
                1704: note <= (-4815);
                1705: note <= (-1697);
                1706: note <= 467;
                1707: note <= 893;
                1708: note <= (-697);
                1709: note <= (-3995);
                1710: note <= (-8192);
                1711: note <= (-12187);
                1712: note <= (-14886);
                1713: note <= (-15491);
                1714: note <= (-13722);
                1715: note <= (-9889);
                1716: note <= (-4815);
                1717: note <= 377;
                1718: note <= 4563;
                1719: note <= 6910;
                1720: note <= 7094;
                1721: note <= 5378;
                1722: note <= 2531;
                1723: note <= (-377);
                1724: note <= (-2279);
                1725: note <= (-2399);
                1726: note <= (-467);
                1727: note <= 3203;
                1728: note <= 7791;
                1729: note <= 12187;
                1730: note <= 15286;
                1731: note <= 16283;
                1732: note <= 14886;
                1733: note <= 11395;
                1734: note <= 6627;
                1735: note <= 1697;
                1736: note <= (-2279);
                1737: note <= (-4473);
                1738: note <= (-4563);
                1739: note <= (-2814);
                1740: note <= 0;
                1741: note <= 2814;
                1742: note <= 4563;
                1743: note <= 4473;
                1744: note <= 2279;
                1745: note <= (-1697);
                1746: note <= (-6627);
                1747: note <= (-11395);
                1748: note <= (-14886);
                1749: note <= (-16283);
                1750: note <= (-15286);
                1751: note <= (-12187);
                1752: note <= (-7791);
                1753: note <= (-3203);
                1754: note <= 467;
                1755: note <= 2399;
                1756: note <= 2279;
                1757: note <= 377;
                1758: note <= (-2531);
                1759: note <= (-5378);
                1760: note <= (-7094);
                1761: note <= (-6910);
                1762: note <= (-4563);
                1763: note <= (-377);
                1764: note <= 4815;
                1765: note <= 9889;
                1766: note <= 13722;
                1767: note <= 15491;
                1768: note <= 14886;
                1769: note <= 12187;
                1770: note <= 8192;
                1771: note <= 3995;
                1772: note <= 697;
                1773: note <= (-893);
                1774: note <= (-467);
                1775: note <= 1697;
                1776: note <= 4815;
                1777: note <= 7815;
                1778: note <= 9626;
                1779: note <= 9474;
                1780: note <= 7094;
                1781: note <= 2814;
                1782: note <= (-2531);
                1783: note <= (-7815);
                1784: note <= (-11910);
                1785: note <= (-13985);
                1786: note <= (-13722);
                1787: note <= (-11395);
                1788: note <= (-7791);
                1789: note <= (-3995);
                1790: note <= (-1098);
                1791: note <= 101;
                1792: note <= (-697);
                1793: note <= (-3203);
                1794: note <= (-6627);
                1795: note <= (-9889);
                1796: note <= (-11910);
                1797: note <= (-11911);
                1798: note <= (-9626);
                1799: note <= (-5378);
                1800: note <= 0;
                1801: note <= 5378;
                1802: note <= 9626;
                1803: note <= 11911;
                1804: note <= 11910;
                1805: note <= 9889;
                1806: note <= 6627;
                1807: note <= 3203;
                1808: note <= 697;
                1809: note <= (-101);
                1810: note <= 1098;
                1811: note <= 3995;
                1812: note <= 7791;
                1813: note <= 11395;
                1814: note <= 13722;
                1815: note <= 13985;
                1816: note <= 11910;
                1817: note <= 7815;
                1818: note <= 2531;
                1819: note <= (-2814);
                1820: note <= (-7094);
                1821: note <= (-9474);
                1822: note <= (-9626);
                1823: note <= (-7815);
                1824: note <= (-4815);
                1825: note <= (-1697);
                1826: note <= 467;
                1827: note <= 893;
                1828: note <= (-697);
                1829: note <= (-3995);
                1830: note <= (-8192);
                1831: note <= (-12187);
                1832: note <= (-14886);
                1833: note <= (-15491);
                1834: note <= (-13722);
                1835: note <= (-9889);
                1836: note <= (-4815);
                1837: note <= 377;
                1838: note <= 4563;
                1839: note <= 6910;
                1840: note <= 7094;
                1841: note <= 5378;
                1842: note <= 2531;
                1843: note <= (-377);
                1844: note <= (-2279);
                1845: note <= (-2399);
                1846: note <= (-467);
                1847: note <= 3203;
                1848: note <= 7791;
                1849: note <= 12187;
                1850: note <= 15286;
                1851: note <= 16283;
                1852: note <= 14886;
                1853: note <= 11395;
                1854: note <= 6627;
                1855: note <= 1697;
                1856: note <= (-2279);
                1857: note <= (-4473);
                1858: note <= (-4563);
                1859: note <= (-2814);
                1860: note <= 0;
                1861: note <= 2814;
                1862: note <= 4563;
                1863: note <= 4473;
                1864: note <= 2279;
                1865: note <= (-1697);
                1866: note <= (-6627);
                1867: note <= (-11395);
                1868: note <= (-14886);
                1869: note <= (-16283);
                1870: note <= (-15286);
                1871: note <= (-12187);
                1872: note <= (-7791);
                1873: note <= (-3203);
                1874: note <= 467;
                1875: note <= 2399;
                1876: note <= 2279;
                1877: note <= 377;
                1878: note <= (-2531);
                1879: note <= (-5378);
                1880: note <= (-7094);
                1881: note <= (-6910);
                1882: note <= (-4563);
                1883: note <= (-377);
                1884: note <= 4815;
                1885: note <= 9889;
                1886: note <= 13722;
                1887: note <= 15491;
                1888: note <= 14886;
                1889: note <= 12187;
                1890: note <= 8192;
                1891: note <= 3995;
                1892: note <= 697;
                1893: note <= (-893);
                1894: note <= (-467);
                1895: note <= 1697;
                1896: note <= 4815;
                1897: note <= 7815;
                1898: note <= 9626;
                1899: note <= 9474;
                1900: note <= 7094;
                1901: note <= 2814;
                1902: note <= (-2531);
                1903: note <= (-7815);
                1904: note <= (-11910);
                1905: note <= (-13985);
                1906: note <= (-13722);
                1907: note <= (-11395);
                1908: note <= (-7791);
                1909: note <= (-3995);
                1910: note <= (-1098);
                1911: note <= 101;
                1912: note <= (-697);
                1913: note <= (-3203);
                1914: note <= (-6627);
                1915: note <= (-9889);
                1916: note <= (-11910);
                1917: note <= (-11911);
                1918: note <= (-9626);
                1919: note <= (-5378);
                1920: note <= 0;
                1921: note <= 5378;
                1922: note <= 9626;
                1923: note <= 11911;
                1924: note <= 11910;
                1925: note <= 9889;
                1926: note <= 6627;
                1927: note <= 3203;
                1928: note <= 697;
                1929: note <= (-101);
                1930: note <= 1098;
                1931: note <= 3995;
                1932: note <= 7791;
                1933: note <= 11395;
                1934: note <= 13722;
                1935: note <= 13985;
                1936: note <= 11910;
                1937: note <= 7815;
                1938: note <= 2531;
                1939: note <= (-2814);
                1940: note <= (-7094);
                1941: note <= (-9474);
                1942: note <= (-9626);
                1943: note <= (-7815);
                1944: note <= (-4815);
                1945: note <= (-1697);
                1946: note <= 467;
                1947: note <= 893;
                1948: note <= (-697);
                1949: note <= (-3995);
                1950: note <= (-8192);
                1951: note <= (-12187);
                1952: note <= (-14886);
                1953: note <= (-15491);
                1954: note <= (-13722);
                1955: note <= (-9889);
                1956: note <= (-4815);
                1957: note <= 377;
                1958: note <= 4563;
                1959: note <= 6910;
                1960: note <= 7094;
                1961: note <= 5378;
                1962: note <= 2531;
                1963: note <= (-377);
                1964: note <= (-2279);
                1965: note <= (-2399);
                1966: note <= (-467);
                1967: note <= 3203;
                1968: note <= 7791;
                1969: note <= 12187;
                1970: note <= 15286;
                1971: note <= 16283;
                1972: note <= 14886;
                1973: note <= 11395;
                1974: note <= 6627;
                1975: note <= 1697;
                1976: note <= (-2279);
                1977: note <= (-4473);
                1978: note <= (-4563);
                1979: note <= (-2814);
                1980: note <= 0;
                1981: note <= 2814;
                1982: note <= 4563;
                1983: note <= 4473;
                1984: note <= 2279;
                1985: note <= (-1697);
                1986: note <= (-6627);
                1987: note <= (-11395);
                1988: note <= (-14886);
                1989: note <= (-16283);
                1990: note <= (-15286);
                1991: note <= (-12187);
                1992: note <= (-7791);
                1993: note <= (-3203);
                1994: note <= 467;
                1995: note <= 2399;
                1996: note <= 2279;
                1997: note <= 377;
                1998: note <= (-2531);
                1999: note <= (-5378);
                2000: note <= (-7094);
                2001: note <= (-6910);
                2002: note <= (-4563);
                2003: note <= (-377);
                2004: note <= 4815;
                2005: note <= 9889;
                2006: note <= 13722;
                2007: note <= 15491;
                2008: note <= 14886;
                2009: note <= 12187;
                2010: note <= 8192;
                2011: note <= 3995;
                2012: note <= 697;
                2013: note <= (-893);
                2014: note <= (-467);
                2015: note <= 1697;
                2016: note <= 4815;
                2017: note <= 7815;
                2018: note <= 9626;
                2019: note <= 9474;
                2020: note <= 7094;
                2021: note <= 2814;
                2022: note <= (-2531);
                2023: note <= (-7815);
                2024: note <= (-11910);
                2025: note <= (-13985);
                2026: note <= (-13722);
                2027: note <= (-11395);
                2028: note <= (-7791);
                2029: note <= (-3995);
                2030: note <= (-1098);
                2031: note <= 101;
                2032: note <= (-697);
                2033: note <= (-3203);
                2034: note <= (-6627);
                2035: note <= (-9889);
                2036: note <= (-11910);
                2037: note <= (-11911);
                2038: note <= (-9626);
                2039: note <= (-5378);
                2040: note <= 0;
                2041: note <= 5378;
                2042: note <= 9626;
                2043: note <= 11911;
                2044: note <= 11910;
                2045: note <= 9889;
                2046: note <= 6627;
                2047: note <= 3203;
                2048: note <= 697;
                2049: note <= (-101);
                2050: note <= 1098;
                2051: note <= 3995;
                2052: note <= 7791;
                2053: note <= 11395;
                2054: note <= 13722;
                2055: note <= 13985;
                2056: note <= 11910;
                2057: note <= 7815;
                2058: note <= 2531;
                2059: note <= (-2814);
                2060: note <= (-7094);
                2061: note <= (-9474);
                2062: note <= (-9626);
                2063: note <= (-7815);
                2064: note <= (-4815);
                2065: note <= (-1697);
                2066: note <= 467;
                2067: note <= 893;
                2068: note <= (-697);
                2069: note <= (-3995);
                2070: note <= (-8192);
                2071: note <= (-12187);
                2072: note <= (-14886);
                2073: note <= (-15491);
                2074: note <= (-13722);
                2075: note <= (-9889);
                2076: note <= (-4815);
                2077: note <= 377;
                2078: note <= 4563;
                2079: note <= 6910;
                2080: note <= 7094;
                2081: note <= 5378;
                2082: note <= 2531;
                2083: note <= (-377);
                2084: note <= (-2279);
                2085: note <= (-2399);
                2086: note <= (-467);
                2087: note <= 3203;
                2088: note <= 7791;
                2089: note <= 12187;
                2090: note <= 15286;
                2091: note <= 16283;
                2092: note <= 14886;
                2093: note <= 11395;
                2094: note <= 6627;
                2095: note <= 1697;
                2096: note <= (-2279);
                2097: note <= (-4473);
                2098: note <= (-4563);
                2099: note <= (-2814);
                2100: note <= 0;
                2101: note <= 2814;
                2102: note <= 4563;
                2103: note <= 4473;
                2104: note <= 2279;
                2105: note <= (-1697);
                2106: note <= (-6627);
                2107: note <= (-11395);
                2108: note <= (-14886);
                2109: note <= (-16283);
                2110: note <= (-15286);
                2111: note <= (-12187);
                2112: note <= (-7791);
                2113: note <= (-3203);
                2114: note <= 467;
                2115: note <= 2399;
                2116: note <= 2279;
                2117: note <= 377;
                2118: note <= (-2531);
                2119: note <= (-5378);
                2120: note <= (-7094);
                2121: note <= (-6910);
                2122: note <= (-4563);
                2123: note <= (-377);
                2124: note <= 4815;
                2125: note <= 9889;
                2126: note <= 13722;
                2127: note <= 15491;
                2128: note <= 14886;
                2129: note <= 12187;
                2130: note <= 8192;
                2131: note <= 3995;
                2132: note <= 697;
                2133: note <= (-893);
                2134: note <= (-467);
                2135: note <= 1697;
                2136: note <= 4815;
                2137: note <= 7815;
                2138: note <= 9626;
                2139: note <= 9474;
                2140: note <= 7094;
                2141: note <= 2814;
                2142: note <= (-2531);
                2143: note <= (-7815);
                2144: note <= (-11910);
                2145: note <= (-13985);
                2146: note <= (-13722);
                2147: note <= (-11395);
                2148: note <= (-7791);
                2149: note <= (-3995);
                2150: note <= (-1098);
                2151: note <= 101;
                2152: note <= (-697);
                2153: note <= (-3203);
                2154: note <= (-6627);
                2155: note <= (-9889);
                2156: note <= (-11910);
                2157: note <= (-11911);
                2158: note <= (-9626);
                2159: note <= (-5378);
                2160: note <= 0;
                2161: note <= 5378;
                2162: note <= 9626;
                2163: note <= 11911;
                2164: note <= 11910;
                2165: note <= 9889;
                2166: note <= 6627;
                2167: note <= 3203;
                2168: note <= 697;
                2169: note <= (-101);
                2170: note <= 1098;
                2171: note <= 3995;
                2172: note <= 7791;
                2173: note <= 11395;
                2174: note <= 13722;
                2175: note <= 13985;
                2176: note <= 11910;
                2177: note <= 7815;
                2178: note <= 2531;
                2179: note <= (-2814);
                2180: note <= (-7094);
                2181: note <= (-9474);
                2182: note <= (-9626);
                2183: note <= (-7815);
                2184: note <= (-4815);
                2185: note <= (-1697);
                2186: note <= 467;
                2187: note <= 893;
                2188: note <= (-697);
                2189: note <= (-3995);
                2190: note <= (-8192);
                2191: note <= (-12187);
                2192: note <= (-14886);
                2193: note <= (-15491);
                2194: note <= (-13722);
                2195: note <= (-9889);
                2196: note <= (-4815);
                2197: note <= 377;
                2198: note <= 4563;
                2199: note <= 6910;
                2200: note <= 7094;
                2201: note <= 5378;
                2202: note <= 2531;
                2203: note <= (-377);
                2204: note <= (-2279);
                2205: note <= (-2399);
                2206: note <= (-467);
                2207: note <= 3203;
                2208: note <= 7791;
                2209: note <= 12187;
                2210: note <= 15286;
                2211: note <= 16283;
                2212: note <= 14886;
                2213: note <= 11395;
                2214: note <= 6627;
                2215: note <= 1697;
                2216: note <= (-2279);
                2217: note <= (-4473);
                2218: note <= (-4563);
                2219: note <= (-2814);
                2220: note <= 0;
                2221: note <= 2814;
                2222: note <= 4563;
                2223: note <= 4473;
                2224: note <= 2279;
                2225: note <= (-1697);
                2226: note <= (-6627);
                2227: note <= (-11395);
                2228: note <= (-14886);
                2229: note <= (-16283);
                2230: note <= (-15286);
                2231: note <= (-12187);
                2232: note <= (-7791);
                2233: note <= (-3203);
                2234: note <= 467;
                2235: note <= 2399;
                2236: note <= 2279;
                2237: note <= 377;
                2238: note <= (-2531);
                2239: note <= (-5378);
                2240: note <= (-7094);
                2241: note <= (-6910);
                2242: note <= (-4563);
                2243: note <= (-377);
                2244: note <= 4815;
                2245: note <= 9889;
                2246: note <= 13722;
                2247: note <= 15491;
                2248: note <= 14886;
                2249: note <= 12187;
                2250: note <= 8192;
                2251: note <= 3995;
                2252: note <= 697;
                2253: note <= (-893);
                2254: note <= (-467);
                2255: note <= 1697;
                2256: note <= 4815;
                2257: note <= 7815;
                2258: note <= 9626;
                2259: note <= 9474;
                2260: note <= 7094;
                2261: note <= 2814;
                2262: note <= (-2531);
                2263: note <= (-7815);
                2264: note <= (-11910);
                2265: note <= (-13985);
                2266: note <= (-13722);
                2267: note <= (-11395);
                2268: note <= (-7791);
                2269: note <= (-3995);
                2270: note <= (-1098);
                2271: note <= 101;
                2272: note <= (-697);
                2273: note <= (-3203);
                2274: note <= (-6627);
                2275: note <= (-9889);
                2276: note <= (-11910);
                2277: note <= (-11911);
                2278: note <= (-9626);
                2279: note <= (-5378);
                2280: note <= 0;
                2281: note <= 5378;
                2282: note <= 9626;
                2283: note <= 11911;
                2284: note <= 11910;
                2285: note <= 9889;
                2286: note <= 6627;
                2287: note <= 3203;
                2288: note <= 697;
                2289: note <= (-101);
                2290: note <= 1098;
                2291: note <= 3995;
                2292: note <= 7791;
                2293: note <= 11395;
                2294: note <= 13722;
                2295: note <= 13985;
                2296: note <= 11910;
                2297: note <= 7815;
                2298: note <= 2531;
                2299: note <= (-2814);
                2300: note <= (-7094);
                2301: note <= (-9474);
                2302: note <= (-9626);
                2303: note <= (-7815);
                2304: note <= (-4815);
                2305: note <= (-1697);
                2306: note <= 467;
                2307: note <= 893;
                2308: note <= (-697);
                2309: note <= (-3995);
                2310: note <= (-8192);
                2311: note <= (-12187);
                2312: note <= (-14886);
                2313: note <= (-15491);
                2314: note <= (-13722);
                2315: note <= (-9889);
                2316: note <= (-4815);
                2317: note <= 377;
                2318: note <= 4563;
                2319: note <= 6910;
                2320: note <= 7094;
                2321: note <= 5378;
                2322: note <= 2531;
                2323: note <= (-377);
                2324: note <= (-2279);
                2325: note <= (-2399);
                2326: note <= (-467);
                2327: note <= 3203;
                2328: note <= 7791;
                2329: note <= 12187;
                2330: note <= 15286;
                2331: note <= 16283;
                2332: note <= 14886;
                2333: note <= 11395;
                2334: note <= 6627;
                2335: note <= 1697;
                2336: note <= (-2279);
                2337: note <= (-4473);
                2338: note <= (-4563);
                2339: note <= (-2814);
                2340: note <= 0;
                2341: note <= 2814;
                2342: note <= 4563;
                2343: note <= 4473;
                2344: note <= 2279;
                2345: note <= (-1697);
                2346: note <= (-6627);
                2347: note <= (-11395);
                2348: note <= (-14886);
                2349: note <= (-16283);
                2350: note <= (-15286);
                2351: note <= (-12187);
                2352: note <= (-7791);
                2353: note <= (-3203);
                2354: note <= 467;
                2355: note <= 2399;
                2356: note <= 2279;
                2357: note <= 377;
                2358: note <= (-2531);
                2359: note <= (-5378);
                2360: note <= (-7094);
                2361: note <= (-6910);
                2362: note <= (-4563);
                2363: note <= (-377);
                2364: note <= 4815;
                2365: note <= 9889;
                2366: note <= 13722;
                2367: note <= 15491;
                2368: note <= 14886;
                2369: note <= 12187;
                2370: note <= 8192;
                2371: note <= 3995;
                2372: note <= 697;
                2373: note <= (-893);
                2374: note <= (-467);
                2375: note <= 1697;
                2376: note <= 4815;
                2377: note <= 7815;
                2378: note <= 9626;
                2379: note <= 9474;
                2380: note <= 7094;
                2381: note <= 2814;
                2382: note <= (-2531);
                2383: note <= (-7815);
                2384: note <= (-11910);
                2385: note <= (-13985);
                2386: note <= (-13722);
                2387: note <= (-11395);
                2388: note <= (-7791);
                2389: note <= (-3995);
                2390: note <= (-1098);
                2391: note <= 101;
                2392: note <= (-697);
                2393: note <= (-3203);
                2394: note <= (-6627);
                2395: note <= (-9889);
                2396: note <= (-11910);
                2397: note <= (-11911);
                2398: note <= (-9626);
                2399: note <= (-5378);
                2400: note <= 0;
                2401: note <= 5378;
                2402: note <= 9626;
                2403: note <= 11911;
                2404: note <= 11910;
                2405: note <= 9889;
                2406: note <= 6627;
                2407: note <= 3203;
                2408: note <= 697;
                2409: note <= (-101);
                2410: note <= 1098;
                2411: note <= 3995;
                2412: note <= 7791;
                2413: note <= 11395;
                2414: note <= 13722;
                2415: note <= 13985;
                2416: note <= 11910;
                2417: note <= 7815;
                2418: note <= 2531;
                2419: note <= (-2814);
                2420: note <= (-7094);
                2421: note <= (-9474);
                2422: note <= (-9626);
                2423: note <= (-7815);
                2424: note <= (-4815);
                2425: note <= (-1697);
                2426: note <= 467;
                2427: note <= 893;
                2428: note <= (-697);
                2429: note <= (-3995);
                2430: note <= (-8192);
                2431: note <= (-12187);
                2432: note <= (-14886);
                2433: note <= (-15491);
                2434: note <= (-13722);
                2435: note <= (-9889);
                2436: note <= (-4815);
                2437: note <= 377;
                2438: note <= 4563;
                2439: note <= 6910;
                2440: note <= 7094;
                2441: note <= 5378;
                2442: note <= 2531;
                2443: note <= (-377);
                2444: note <= (-2279);
                2445: note <= (-2399);
                2446: note <= (-467);
                2447: note <= 3203;
                2448: note <= 7791;
                2449: note <= 12187;
                2450: note <= 15286;
                2451: note <= 16283;
                2452: note <= 14886;
                2453: note <= 11395;
                2454: note <= 6627;
                2455: note <= 1697;
                2456: note <= (-2279);
                2457: note <= (-4473);
                2458: note <= (-4563);
                2459: note <= (-2814);
                2460: note <= 0;
                2461: note <= 2814;
                2462: note <= 4563;
                2463: note <= 4473;
                2464: note <= 2279;
                2465: note <= (-1697);
                2466: note <= (-6627);
                2467: note <= (-11395);
                2468: note <= (-14886);
                2469: note <= (-16283);
                2470: note <= (-15286);
                2471: note <= (-12187);
                2472: note <= (-7791);
                2473: note <= (-3203);
                2474: note <= 467;
                2475: note <= 2399;
                2476: note <= 2279;
                2477: note <= 377;
                2478: note <= (-2531);
                2479: note <= (-5378);
                2480: note <= (-7094);
                2481: note <= (-6910);
                2482: note <= (-4563);
                2483: note <= (-377);
                2484: note <= 4815;
                2485: note <= 9889;
                2486: note <= 13722;
                2487: note <= 15491;
                2488: note <= 14886;
                2489: note <= 12187;
                2490: note <= 8192;
                2491: note <= 3995;
                2492: note <= 697;
                2493: note <= (-893);
                2494: note <= (-467);
                2495: note <= 1697;
                2496: note <= 4815;
                2497: note <= 7815;
                2498: note <= 9626;
                2499: note <= 9474;
                2500: note <= 7094;
                2501: note <= 2814;
                2502: note <= (-2531);
                2503: note <= (-7815);
                2504: note <= (-11910);
                2505: note <= (-13985);
                2506: note <= (-13722);
                2507: note <= (-11395);
                2508: note <= (-7791);
                2509: note <= (-3995);
                2510: note <= (-1098);
                2511: note <= 101;
                2512: note <= (-697);
                2513: note <= (-3203);
                2514: note <= (-6627);
                2515: note <= (-9889);
                2516: note <= (-11910);
                2517: note <= (-11911);
                2518: note <= (-9626);
                2519: note <= (-5378);
                2520: note <= 0;
                2521: note <= 5378;
                2522: note <= 9626;
                2523: note <= 11911;
                2524: note <= 11910;
                2525: note <= 9889;
                2526: note <= 6627;
                2527: note <= 3203;
                2528: note <= 697;
                2529: note <= (-101);
                2530: note <= 1098;
                2531: note <= 3995;
                2532: note <= 7791;
                2533: note <= 11395;
                2534: note <= 13722;
                2535: note <= 13985;
                2536: note <= 11910;
                2537: note <= 7815;
                2538: note <= 2531;
                2539: note <= (-2814);
                2540: note <= (-7094);
                2541: note <= (-9474);
                2542: note <= (-9626);
                2543: note <= (-7815);
                2544: note <= (-4815);
                2545: note <= (-1697);
                2546: note <= 467;
                2547: note <= 893;
                2548: note <= (-697);
                2549: note <= (-3995);
                2550: note <= (-8192);
                2551: note <= (-12187);
                2552: note <= (-14886);
                2553: note <= (-15491);
                2554: note <= (-13722);
                2555: note <= (-9889);
                2556: note <= (-4815);
                2557: note <= 377;
                2558: note <= 4563;
                2559: note <= 6910;
                2560: note <= 7094;
                2561: note <= 5378;
                2562: note <= 2531;
                2563: note <= (-377);
                2564: note <= (-2279);
                2565: note <= (-2399);
                2566: note <= (-467);
                2567: note <= 3203;
                2568: note <= 7791;
                2569: note <= 12187;
                2570: note <= 15286;
                2571: note <= 16283;
                2572: note <= 14886;
                2573: note <= 11395;
                2574: note <= 6627;
                2575: note <= 1697;
                2576: note <= (-2279);
                2577: note <= (-4473);
                2578: note <= (-4563);
                2579: note <= (-2814);
                2580: note <= 0;
                2581: note <= 2814;
                2582: note <= 4563;
                2583: note <= 4473;
                2584: note <= 2279;
                2585: note <= (-1697);
                2586: note <= (-6627);
                2587: note <= (-11395);
                2588: note <= (-14886);
                2589: note <= (-16283);
                2590: note <= (-15286);
                2591: note <= (-12187);
                2592: note <= (-7791);
                2593: note <= (-3203);
                2594: note <= 467;
                2595: note <= 2399;
                2596: note <= 2279;
                2597: note <= 377;
                2598: note <= (-2531);
                2599: note <= (-5378);
                2600: note <= (-7094);
                2601: note <= (-6910);
                2602: note <= (-4563);
                2603: note <= (-377);
                2604: note <= 4815;
                2605: note <= 9889;
                2606: note <= 13722;
                2607: note <= 15491;
                2608: note <= 14886;
                2609: note <= 12187;
                2610: note <= 8192;
                2611: note <= 3995;
                2612: note <= 697;
                2613: note <= (-893);
                2614: note <= (-467);
                2615: note <= 1697;
                2616: note <= 4815;
                2617: note <= 7815;
                2618: note <= 9626;
                2619: note <= 9474;
                2620: note <= 7094;
                2621: note <= 2814;
                2622: note <= (-2531);
                2623: note <= (-7815);
                2624: note <= (-11910);
                2625: note <= (-13985);
                2626: note <= (-13722);
                2627: note <= (-11395);
                2628: note <= (-7791);
                2629: note <= (-3995);
                2630: note <= (-1098);
                2631: note <= 101;
                2632: note <= (-697);
                2633: note <= (-3203);
                2634: note <= (-6627);
                2635: note <= (-9889);
                2636: note <= (-11910);
                2637: note <= (-11911);
                2638: note <= (-9626);
                2639: note <= (-5378);
                2640: note <= 0;
                2641: note <= 5378;
                2642: note <= 9626;
                2643: note <= 11911;
                2644: note <= 11910;
                2645: note <= 9889;
                2646: note <= 6627;
                2647: note <= 3203;
                2648: note <= 697;
                2649: note <= (-101);
                2650: note <= 1098;
                2651: note <= 3995;
                2652: note <= 7791;
                2653: note <= 11395;
                2654: note <= 13722;
                2655: note <= 13985;
                2656: note <= 11910;
                2657: note <= 7815;
                2658: note <= 2531;
                2659: note <= (-2814);
                2660: note <= (-7094);
                2661: note <= (-9474);
                2662: note <= (-9626);
                2663: note <= (-7815);
                2664: note <= (-4815);
                2665: note <= (-1697);
                2666: note <= 467;
                2667: note <= 893;
                2668: note <= (-697);
                2669: note <= (-3995);
                2670: note <= (-8192);
                2671: note <= (-12187);
                2672: note <= (-14886);
                2673: note <= (-15491);
                2674: note <= (-13722);
                2675: note <= (-9889);
                2676: note <= (-4815);
                2677: note <= 377;
                2678: note <= 4563;
                2679: note <= 6910;
                2680: note <= 7094;
                2681: note <= 5378;
                2682: note <= 2531;
                2683: note <= (-377);
                2684: note <= (-2279);
                2685: note <= (-2399);
                2686: note <= (-467);
                2687: note <= 3203;
                2688: note <= 7791;
                2689: note <= 12187;
                2690: note <= 15286;
                2691: note <= 16283;
                2692: note <= 14886;
                2693: note <= 11395;
                2694: note <= 6627;
                2695: note <= 1697;
                2696: note <= (-2279);
                2697: note <= (-4473);
                2698: note <= (-4563);
                2699: note <= (-2814);
                2700: note <= 0;
                2701: note <= 2814;
                2702: note <= 4563;
                2703: note <= 4473;
                2704: note <= 2279;
                2705: note <= (-1697);
                2706: note <= (-6627);
                2707: note <= (-11395);
                2708: note <= (-14886);
                2709: note <= (-16283);
                2710: note <= (-15286);
                2711: note <= (-12187);
                2712: note <= (-7791);
                2713: note <= (-3203);
                2714: note <= 467;
                2715: note <= 2399;
                2716: note <= 2279;
                2717: note <= 377;
                2718: note <= (-2531);
                2719: note <= (-5378);
                2720: note <= (-7094);
                2721: note <= (-6910);
                2722: note <= (-4563);
                2723: note <= (-377);
                2724: note <= 4815;
                2725: note <= 9889;
                2726: note <= 13722;
                2727: note <= 15491;
                2728: note <= 14886;
                2729: note <= 12187;
                2730: note <= 8192;
                2731: note <= 3995;
                2732: note <= 697;
                2733: note <= (-893);
                2734: note <= (-467);
                2735: note <= 1697;
                2736: note <= 4815;
                2737: note <= 7815;
                2738: note <= 9626;
                2739: note <= 9474;
                2740: note <= 7094;
                2741: note <= 2814;
                2742: note <= (-2531);
                2743: note <= (-7815);
                2744: note <= (-11910);
                2745: note <= (-13985);
                2746: note <= (-13722);
                2747: note <= (-11395);
                2748: note <= (-7791);
                2749: note <= (-3995);
                2750: note <= (-1098);
                2751: note <= 101;
                2752: note <= (-697);
                2753: note <= (-3203);
                2754: note <= (-6627);
                2755: note <= (-9889);
                2756: note <= (-11910);
                2757: note <= (-11911);
                2758: note <= (-9626);
                2759: note <= (-5378);
                2760: note <= 0;
                2761: note <= 5378;
                2762: note <= 9626;
                2763: note <= 11911;
                2764: note <= 11910;
                2765: note <= 9889;
                2766: note <= 6627;
                2767: note <= 3203;
                2768: note <= 697;
                2769: note <= (-101);
                2770: note <= 1098;
                2771: note <= 3995;
                2772: note <= 7791;
                2773: note <= 11395;
                2774: note <= 13722;
                2775: note <= 13985;
                2776: note <= 11910;
                2777: note <= 7815;
                2778: note <= 2531;
                2779: note <= (-2814);
                2780: note <= (-7094);
                2781: note <= (-9474);
                2782: note <= (-9626);
                2783: note <= (-7815);
                2784: note <= (-4815);
                2785: note <= (-1697);
                2786: note <= 467;
                2787: note <= 893;
                2788: note <= (-697);
                2789: note <= (-3995);
                2790: note <= (-8192);
                2791: note <= (-12187);
                2792: note <= (-14886);
                2793: note <= (-15491);
                2794: note <= (-13722);
                2795: note <= (-9889);
                2796: note <= (-4815);
                2797: note <= 377;
                2798: note <= 4563;
                2799: note <= 6910;
                2800: note <= 7094;
                2801: note <= 5378;
                2802: note <= 2531;
                2803: note <= (-377);
                2804: note <= (-2279);
                2805: note <= (-2399);
                2806: note <= (-467);
                2807: note <= 3203;
                2808: note <= 7791;
                2809: note <= 12187;
                2810: note <= 15286;
                2811: note <= 16283;
                2812: note <= 14886;
                2813: note <= 11395;
                2814: note <= 6627;
                2815: note <= 1697;
                2816: note <= (-2279);
                2817: note <= (-4473);
                2818: note <= (-4563);
                2819: note <= (-2814);
                2820: note <= 0;
                2821: note <= 2814;
                2822: note <= 4563;
                2823: note <= 4473;
                2824: note <= 2279;
                2825: note <= (-1697);
                2826: note <= (-6627);
                2827: note <= (-11395);
                2828: note <= (-14886);
                2829: note <= (-16283);
                2830: note <= (-15286);
                2831: note <= (-12187);
                2832: note <= (-7791);
                2833: note <= (-3203);
                2834: note <= 467;
                2835: note <= 2399;
                2836: note <= 2279;
                2837: note <= 377;
                2838: note <= (-2531);
                2839: note <= (-5378);
                2840: note <= (-7094);
                2841: note <= (-6910);
                2842: note <= (-4563);
                2843: note <= (-377);
                2844: note <= 4815;
                2845: note <= 9889;
                2846: note <= 13722;
                2847: note <= 15491;
                2848: note <= 14886;
                2849: note <= 12187;
                2850: note <= 8192;
                2851: note <= 3995;
                2852: note <= 697;
                2853: note <= (-893);
                2854: note <= (-467);
                2855: note <= 1697;
                2856: note <= 4815;
                2857: note <= 7815;
                2858: note <= 9626;
                2859: note <= 9474;
                2860: note <= 7094;
                2861: note <= 2814;
                2862: note <= (-2531);
                2863: note <= (-7815);
                2864: note <= (-11910);
                2865: note <= (-13985);
                2866: note <= (-13722);
                2867: note <= (-11395);
                2868: note <= (-7791);
                2869: note <= (-3995);
                2870: note <= (-1098);
                2871: note <= 101;
                2872: note <= (-697);
                2873: note <= (-3203);
                2874: note <= (-6627);
                2875: note <= (-9889);
                2876: note <= (-11910);
                2877: note <= (-11911);
                2878: note <= (-9626);
                2879: note <= (-5378);
                2880: note <= 0;
                2881: note <= 5378;
                2882: note <= 9626;
                2883: note <= 11911;
                2884: note <= 11910;
                2885: note <= 9889;
                2886: note <= 6627;
                2887: note <= 3203;
                2888: note <= 697;
                2889: note <= (-101);
                2890: note <= 1098;
                2891: note <= 3995;
                2892: note <= 7791;
                2893: note <= 11395;
                2894: note <= 13722;
                2895: note <= 13985;
                2896: note <= 11910;
                2897: note <= 7815;
                2898: note <= 2531;
                2899: note <= (-2814);
                2900: note <= (-7094);
                2901: note <= (-9474);
                2902: note <= (-9626);
                2903: note <= (-7815);
                2904: note <= (-4815);
                2905: note <= (-1697);
                2906: note <= 467;
                2907: note <= 893;
                2908: note <= (-697);
                2909: note <= (-3995);
                2910: note <= (-8192);
                2911: note <= (-12187);
                2912: note <= (-14886);
                2913: note <= (-15491);
                2914: note <= (-13722);
                2915: note <= (-9889);
                2916: note <= (-4815);
                2917: note <= 377;
                2918: note <= 4563;
                2919: note <= 6910;
                2920: note <= 7094;
                2921: note <= 5378;
                2922: note <= 2531;
                2923: note <= (-377);
                2924: note <= (-2279);
                2925: note <= (-2399);
                2926: note <= (-467);
                2927: note <= 3203;
                2928: note <= 7791;
                2929: note <= 12187;
                2930: note <= 15286;
                2931: note <= 16283;
                2932: note <= 14886;
                2933: note <= 11395;
                2934: note <= 6627;
                2935: note <= 1697;
                2936: note <= (-2279);
                2937: note <= (-4473);
                2938: note <= (-4563);
                2939: note <= (-2814);
                2940: note <= 0;
                2941: note <= 2814;
                2942: note <= 4563;
                2943: note <= 4473;
                2944: note <= 2279;
                2945: note <= (-1697);
                2946: note <= (-6627);
                2947: note <= (-11395);
                2948: note <= (-14886);
                2949: note <= (-16283);
                2950: note <= (-15286);
                2951: note <= (-12187);
                2952: note <= (-7791);
                2953: note <= (-3203);
                2954: note <= 467;
                2955: note <= 2399;
                2956: note <= 2279;
                2957: note <= 377;
                2958: note <= (-2531);
                2959: note <= (-5378);
                2960: note <= (-7094);
                2961: note <= (-6910);
                2962: note <= (-4563);
                2963: note <= (-377);
                2964: note <= 4815;
                2965: note <= 9889;
                2966: note <= 13722;
                2967: note <= 15491;
                2968: note <= 14886;
                2969: note <= 12187;
                2970: note <= 8192;
                2971: note <= 3995;
                2972: note <= 697;
                2973: note <= (-893);
                2974: note <= (-467);
                2975: note <= 1697;
                2976: note <= 4815;
                2977: note <= 7815;
                2978: note <= 9626;
                2979: note <= 9474;
                2980: note <= 7094;
                2981: note <= 2814;
                2982: note <= (-2531);
                2983: note <= (-7815);
                2984: note <= (-11910);
                2985: note <= (-13985);
                2986: note <= (-13722);
                2987: note <= (-11395);
                2988: note <= (-7791);
                2989: note <= (-3995);
                2990: note <= (-1098);
                2991: note <= 101;
                2992: note <= (-697);
                2993: note <= (-3203);
                2994: note <= (-6627);
                2995: note <= (-9889);
                2996: note <= (-11910);
                2997: note <= (-11911);
                2998: note <= (-9626);
                2999: note <= (-5378);
                3000: note <= 0;
                3001: note <= 5378;
                3002: note <= 9626;
                3003: note <= 11911;
                3004: note <= 11910;
                3005: note <= 9889;
                3006: note <= 6627;
                3007: note <= 3203;
                3008: note <= 697;
                3009: note <= (-101);
                3010: note <= 1098;
                3011: note <= 3995;
                3012: note <= 7791;
                3013: note <= 11395;
                3014: note <= 13722;
                3015: note <= 13985;
                3016: note <= 11910;
                3017: note <= 7815;
                3018: note <= 2531;
                3019: note <= (-2814);
                3020: note <= (-7094);
                3021: note <= (-9474);
                3022: note <= (-9626);
                3023: note <= (-7815);
                3024: note <= (-4815);
                3025: note <= (-1697);
                3026: note <= 467;
                3027: note <= 893;
                3028: note <= (-697);
                3029: note <= (-3995);
                3030: note <= (-8192);
                3031: note <= (-12187);
                3032: note <= (-14886);
                3033: note <= (-15491);
                3034: note <= (-13722);
                3035: note <= (-9889);
                3036: note <= (-4815);
                3037: note <= 377;
                3038: note <= 4563;
                3039: note <= 6910;
                3040: note <= 7094;
                3041: note <= 5378;
                3042: note <= 2531;
                3043: note <= (-377);
                3044: note <= (-2279);
                3045: note <= (-2399);
                3046: note <= (-467);
                3047: note <= 3203;
                3048: note <= 7791;
                3049: note <= 12187;
                3050: note <= 15286;
                3051: note <= 16283;
                3052: note <= 14886;
                3053: note <= 11395;
                3054: note <= 6627;
                3055: note <= 1697;
                3056: note <= (-2279);
                3057: note <= (-4473);
                3058: note <= (-4563);
                3059: note <= (-2814);
                3060: note <= 0;
                3061: note <= 2814;
                3062: note <= 4563;
                3063: note <= 4473;
                3064: note <= 2279;
                3065: note <= (-1697);
                3066: note <= (-6627);
                3067: note <= (-11395);
                3068: note <= (-14886);
                3069: note <= (-16283);
                3070: note <= (-15286);
                3071: note <= (-12187);
                3072: note <= (-7791);
                3073: note <= (-3203);
                3074: note <= 467;
                3075: note <= 2399;
                3076: note <= 2279;
                3077: note <= 377;
                3078: note <= (-2531);
                3079: note <= (-5378);
                3080: note <= (-7094);
                3081: note <= (-6910);
                3082: note <= (-4563);
                3083: note <= (-377);
                3084: note <= 4815;
                3085: note <= 9889;
                3086: note <= 13722;
                3087: note <= 15491;
                3088: note <= 14886;
                3089: note <= 12187;
                3090: note <= 8192;
                3091: note <= 3995;
                3092: note <= 697;
                3093: note <= (-893);
                3094: note <= (-467);
                3095: note <= 1697;
                3096: note <= 4815;
                3097: note <= 7815;
                3098: note <= 9626;
                3099: note <= 9474;
                3100: note <= 7094;
                3101: note <= 2814;
                3102: note <= (-2531);
                3103: note <= (-7815);
                3104: note <= (-11910);
                3105: note <= (-13985);
                3106: note <= (-13722);
                3107: note <= (-11395);
                3108: note <= (-7791);
                3109: note <= (-3995);
                3110: note <= (-1098);
                3111: note <= 101;
                3112: note <= (-697);
                3113: note <= (-3203);
                3114: note <= (-6627);
                3115: note <= (-9889);
                3116: note <= (-11910);
                3117: note <= (-11911);
                3118: note <= (-9626);
                3119: note <= (-5378);
                3120: note <= 0;
                3121: note <= 5378;
                3122: note <= 9626;
                3123: note <= 11911;
                3124: note <= 11910;
                3125: note <= 9889;
                3126: note <= 6627;
                3127: note <= 3203;
                3128: note <= 697;
                3129: note <= (-101);
                3130: note <= 1098;
                3131: note <= 3995;
                3132: note <= 7791;
                3133: note <= 11395;
                3134: note <= 13722;
                3135: note <= 13985;
                3136: note <= 11910;
                3137: note <= 7815;
                3138: note <= 2531;
                3139: note <= (-2814);
                3140: note <= (-7094);
                3141: note <= (-9474);
                3142: note <= (-9626);
                3143: note <= (-7815);
                3144: note <= (-4815);
                3145: note <= (-1697);
                3146: note <= 467;
                3147: note <= 893;
                3148: note <= (-697);
                3149: note <= (-3995);
                3150: note <= (-8192);
                3151: note <= (-12187);
                3152: note <= (-14886);
                3153: note <= (-15491);
                3154: note <= (-13722);
                3155: note <= (-9889);
                3156: note <= (-4815);
                3157: note <= 377;
                3158: note <= 4563;
                3159: note <= 6910;
                3160: note <= 7094;
                3161: note <= 5378;
                3162: note <= 2531;
                3163: note <= (-377);
                3164: note <= (-2279);
                3165: note <= (-2399);
                3166: note <= (-467);
                3167: note <= 3203;
                3168: note <= 7791;
                3169: note <= 12187;
                3170: note <= 15286;
                3171: note <= 16283;
                3172: note <= 14886;
                3173: note <= 11395;
                3174: note <= 6627;
                3175: note <= 1697;
                3176: note <= (-2279);
                3177: note <= (-4473);
                3178: note <= (-4563);
                3179: note <= (-2814);
                3180: note <= 0;
                3181: note <= 2814;
                3182: note <= 4563;
                3183: note <= 4473;
                3184: note <= 2279;
                3185: note <= (-1697);
                3186: note <= (-6627);
                3187: note <= (-11395);
                3188: note <= (-14886);
                3189: note <= (-16283);
                3190: note <= (-15286);
                3191: note <= (-12187);
                3192: note <= (-7791);
                3193: note <= (-3203);
                3194: note <= 467;
                3195: note <= 2399;
                3196: note <= 2279;
                3197: note <= 377;
                3198: note <= (-2531);
                3199: note <= (-5378);
                3200: note <= (-7094);
                3201: note <= (-6910);
                3202: note <= (-4563);
                3203: note <= (-377);
                3204: note <= 4815;
                3205: note <= 9889;
                3206: note <= 13722;
                3207: note <= 15491;
                3208: note <= 14886;
                3209: note <= 12187;
                3210: note <= 8192;
                3211: note <= 3995;
                3212: note <= 697;
                3213: note <= (-893);
                3214: note <= (-467);
                3215: note <= 1697;
                3216: note <= 4815;
                3217: note <= 7815;
                3218: note <= 9626;
                3219: note <= 9474;
                3220: note <= 7094;
                3221: note <= 2814;
                3222: note <= (-2531);
                3223: note <= (-7815);
                3224: note <= (-11910);
                3225: note <= (-13985);
                3226: note <= (-13722);
                3227: note <= (-11395);
                3228: note <= (-7791);
                3229: note <= (-3995);
                3230: note <= (-1098);
                3231: note <= 101;
                3232: note <= (-697);
                3233: note <= (-3203);
                3234: note <= (-6627);
                3235: note <= (-9889);
                3236: note <= (-11910);
                3237: note <= (-11911);
                3238: note <= (-9626);
                3239: note <= (-5378);
                3240: note <= 0;
                3241: note <= 5378;
                3242: note <= 9626;
                3243: note <= 11911;
                3244: note <= 11910;
                3245: note <= 9889;
                3246: note <= 6627;
                3247: note <= 3203;
                3248: note <= 697;
                3249: note <= (-101);
                3250: note <= 1098;
                3251: note <= 3995;
                3252: note <= 7791;
                3253: note <= 11395;
                3254: note <= 13722;
                3255: note <= 13985;
                3256: note <= 11910;
                3257: note <= 7815;
                3258: note <= 2531;
                3259: note <= (-2814);
                3260: note <= (-7094);
                3261: note <= (-9474);
                3262: note <= (-9626);
                3263: note <= (-7815);
                3264: note <= (-4815);
                3265: note <= (-1697);
                3266: note <= 467;
                3267: note <= 893;
                3268: note <= (-697);
                3269: note <= (-3995);
                3270: note <= (-8192);
                3271: note <= (-12187);
                3272: note <= (-14886);
                3273: note <= (-15491);
                3274: note <= (-13722);
                3275: note <= (-9889);
                3276: note <= (-4815);
                3277: note <= 377;
                3278: note <= 4563;
                3279: note <= 6910;
                3280: note <= 7094;
                3281: note <= 5378;
                3282: note <= 2531;
                3283: note <= (-377);
                3284: note <= (-2279);
                3285: note <= (-2399);
                3286: note <= (-467);
                3287: note <= 3203;
                3288: note <= 7791;
                3289: note <= 12187;
                3290: note <= 15286;
                3291: note <= 16283;
                3292: note <= 14886;
                3293: note <= 11395;
                3294: note <= 6627;
                3295: note <= 1697;
                3296: note <= (-2279);
                3297: note <= (-4473);
                3298: note <= (-4563);
                3299: note <= (-2814);
                3300: note <= 0;
                3301: note <= 2814;
                3302: note <= 4563;
                3303: note <= 4473;
                3304: note <= 2279;
                3305: note <= (-1697);
                3306: note <= (-6627);
                3307: note <= (-11395);
                3308: note <= (-14886);
                3309: note <= (-16283);
                3310: note <= (-15286);
                3311: note <= (-12187);
                3312: note <= (-7791);
                3313: note <= (-3203);
                3314: note <= 467;
                3315: note <= 2399;
                3316: note <= 2279;
                3317: note <= 377;
                3318: note <= (-2531);
                3319: note <= (-5378);
                3320: note <= (-7094);
                3321: note <= (-6910);
                3322: note <= (-4563);
                3323: note <= (-377);
                3324: note <= 4815;
                3325: note <= 9889;
                3326: note <= 13722;
                3327: note <= 15491;
                3328: note <= 14886;
                3329: note <= 12187;
                3330: note <= 8192;
                3331: note <= 3995;
                3332: note <= 697;
                3333: note <= (-893);
                3334: note <= (-467);
                3335: note <= 1697;
                3336: note <= 4815;
                3337: note <= 7815;
                3338: note <= 9626;
                3339: note <= 9474;
                3340: note <= 7094;
                3341: note <= 2814;
                3342: note <= (-2531);
                3343: note <= (-7815);
                3344: note <= (-11910);
                3345: note <= (-13985);
                3346: note <= (-13722);
                3347: note <= (-11395);
                3348: note <= (-7791);
                3349: note <= (-3995);
                3350: note <= (-1098);
                3351: note <= 101;
                3352: note <= (-697);
                3353: note <= (-3203);
                3354: note <= (-6627);
                3355: note <= (-9889);
                3356: note <= (-11910);
                3357: note <= (-11911);
                3358: note <= (-9626);
                3359: note <= (-5378);
                3360: note <= 0;
                3361: note <= 5378;
                3362: note <= 9626;
                3363: note <= 11911;
                3364: note <= 11910;
                3365: note <= 9889;
                3366: note <= 6627;
                3367: note <= 3203;
                3368: note <= 697;
                3369: note <= (-101);
                3370: note <= 1098;
                3371: note <= 3995;
                3372: note <= 7791;
                3373: note <= 11395;
                3374: note <= 13722;
                3375: note <= 13985;
                3376: note <= 11910;
                3377: note <= 7815;
                3378: note <= 2531;
                3379: note <= (-2814);
                3380: note <= (-7094);
                3381: note <= (-9474);
                3382: note <= (-9626);
                3383: note <= (-7815);
                3384: note <= (-4815);
                3385: note <= (-1697);
                3386: note <= 467;
                3387: note <= 893;
                3388: note <= (-697);
                3389: note <= (-3995);
                3390: note <= (-8192);
                3391: note <= (-12187);
                3392: note <= (-14886);
                3393: note <= (-15491);
                3394: note <= (-13722);
                3395: note <= (-9889);
                3396: note <= (-4815);
                3397: note <= 377;
                3398: note <= 4563;
                3399: note <= 6910;
                3400: note <= 7094;
                3401: note <= 5378;
                3402: note <= 2531;
                3403: note <= (-377);
                3404: note <= (-2279);
                3405: note <= (-2399);
                3406: note <= (-467);
                3407: note <= 3203;
                3408: note <= 7791;
                3409: note <= 12187;
                3410: note <= 15286;
                3411: note <= 16283;
                3412: note <= 14886;
                3413: note <= 11395;
                3414: note <= 6627;
                3415: note <= 1697;
                3416: note <= (-2279);
                3417: note <= (-4473);
                3418: note <= (-4563);
                3419: note <= (-2814);
                3420: note <= 0;
                3421: note <= 2814;
                3422: note <= 4563;
                3423: note <= 4473;
                3424: note <= 2279;
                3425: note <= (-1697);
                3426: note <= (-6627);
                3427: note <= (-11395);
                3428: note <= (-14886);
                3429: note <= (-16283);
                3430: note <= (-15286);
                3431: note <= (-12187);
                3432: note <= (-7791);
                3433: note <= (-3203);
                3434: note <= 467;
                3435: note <= 2399;
                3436: note <= 2279;
                3437: note <= 377;
                3438: note <= (-2531);
                3439: note <= (-5378);
                3440: note <= (-7094);
                3441: note <= (-6910);
                3442: note <= (-4563);
                3443: note <= (-377);
                3444: note <= 4815;
                3445: note <= 9889;
                3446: note <= 13722;
                3447: note <= 15491;
                3448: note <= 14886;
                3449: note <= 12187;
                3450: note <= 8192;
                3451: note <= 3995;
                3452: note <= 697;
                3453: note <= (-893);
                3454: note <= (-467);
                3455: note <= 1697;
                3456: note <= 4815;
                3457: note <= 7815;
                3458: note <= 9626;
                3459: note <= 9474;
                3460: note <= 7094;
                3461: note <= 2814;
                3462: note <= (-2531);
                3463: note <= (-7815);
                3464: note <= (-11910);
                3465: note <= (-13985);
                3466: note <= (-13722);
                3467: note <= (-11395);
                3468: note <= (-7791);
                3469: note <= (-3995);
                3470: note <= (-1098);
                3471: note <= 101;
                3472: note <= (-697);
                3473: note <= (-3203);
                3474: note <= (-6627);
                3475: note <= (-9889);
                3476: note <= (-11910);
                3477: note <= (-11911);
                3478: note <= (-9626);
                3479: note <= (-5378);
                3480: note <= 0;
                3481: note <= 5378;
                3482: note <= 9626;
                3483: note <= 11911;
                3484: note <= 11910;
                3485: note <= 9889;
                3486: note <= 6627;
                3487: note <= 3203;
                3488: note <= 697;
                3489: note <= (-101);
                3490: note <= 1098;
                3491: note <= 3995;
                3492: note <= 7791;
                3493: note <= 11395;
                3494: note <= 13722;
                3495: note <= 13985;
                3496: note <= 11910;
                3497: note <= 7815;
                3498: note <= 2531;
                3499: note <= (-2814);
                3500: note <= (-7094);
                3501: note <= (-9474);
                3502: note <= (-9626);
                3503: note <= (-7815);
                3504: note <= (-4815);
                3505: note <= (-1697);
                3506: note <= 467;
                3507: note <= 893;
                3508: note <= (-697);
                3509: note <= (-3995);
                3510: note <= (-8192);
                3511: note <= (-12187);
                3512: note <= (-14886);
                3513: note <= (-15491);
                3514: note <= (-13722);
                3515: note <= (-9889);
                3516: note <= (-4815);
                3517: note <= 377;
                3518: note <= 4563;
                3519: note <= 6910;
                3520: note <= 7094;
                3521: note <= 5378;
                3522: note <= 2531;
                3523: note <= (-377);
                3524: note <= (-2279);
                3525: note <= (-2399);
                3526: note <= (-467);
                3527: note <= 3203;
                3528: note <= 7791;
                3529: note <= 12187;
                3530: note <= 15286;
                3531: note <= 16283;
                3532: note <= 14886;
                3533: note <= 11395;
                3534: note <= 6627;
                3535: note <= 1697;
                3536: note <= (-2279);
                3537: note <= (-4473);
                3538: note <= (-4563);
                3539: note <= (-2814);
                3540: note <= 0;
                3541: note <= 2814;
                3542: note <= 4563;
                3543: note <= 4473;
                3544: note <= 2279;
                3545: note <= (-1697);
                3546: note <= (-6627);
                3547: note <= (-11395);
                3548: note <= (-14886);
                3549: note <= (-16283);
                3550: note <= (-15286);
                3551: note <= (-12187);
                3552: note <= (-7791);
                3553: note <= (-3203);
                3554: note <= 467;
                3555: note <= 2399;
                3556: note <= 2279;
                3557: note <= 377;
                3558: note <= (-2531);
                3559: note <= (-5378);
                3560: note <= (-7094);
                3561: note <= (-6910);
                3562: note <= (-4563);
                3563: note <= (-377);
                3564: note <= 4815;
                3565: note <= 9889;
                3566: note <= 13722;
                3567: note <= 15491;
                3568: note <= 14886;
                3569: note <= 12187;
                3570: note <= 8192;
                3571: note <= 3995;
                3572: note <= 697;
                3573: note <= (-893);
                3574: note <= (-467);
                3575: note <= 1697;
                3576: note <= 4815;
                3577: note <= 7815;
                3578: note <= 9626;
                3579: note <= 9474;
                3580: note <= 7094;
                3581: note <= 2814;
                3582: note <= (-2531);
                3583: note <= (-7815);
                3584: note <= (-11910);
                3585: note <= (-13985);
                3586: note <= (-13722);
                3587: note <= (-11395);
                3588: note <= (-7791);
                3589: note <= (-3995);
                3590: note <= (-1098);
                3591: note <= 101;
                3592: note <= (-697);
                3593: note <= (-3203);
                3594: note <= (-6627);
                3595: note <= (-9889);
                3596: note <= (-11910);
                3597: note <= (-11911);
                3598: note <= (-9626);
                3599: note <= (-5378);
                3600: note <= 0;
                3601: note <= 5378;
                3602: note <= 9626;
                3603: note <= 11911;
                3604: note <= 11910;
                3605: note <= 9889;
                3606: note <= 6627;
                3607: note <= 3203;
                3608: note <= 697;
                3609: note <= (-101);
                3610: note <= 1098;
                3611: note <= 3995;
                3612: note <= 7791;
                3613: note <= 11395;
                3614: note <= 13722;
                3615: note <= 13985;
                3616: note <= 11910;
                3617: note <= 7815;
                3618: note <= 2531;
                3619: note <= (-2814);
                3620: note <= (-7094);
                3621: note <= (-9474);
                3622: note <= (-9626);
                3623: note <= (-7815);
                3624: note <= (-4815);
                3625: note <= (-1697);
                3626: note <= 467;
                3627: note <= 893;
                3628: note <= (-697);
                3629: note <= (-3995);
                3630: note <= (-8192);
                3631: note <= (-12187);
                3632: note <= (-14886);
                3633: note <= (-15491);
                3634: note <= (-13722);
                3635: note <= (-9889);
                3636: note <= (-4815);
                3637: note <= 377;
                3638: note <= 4563;
                3639: note <= 6910;
                3640: note <= 7094;
                3641: note <= 5378;
                3642: note <= 2531;
                3643: note <= (-377);
                3644: note <= (-2279);
                3645: note <= (-2399);
                3646: note <= (-467);
                3647: note <= 3203;
                3648: note <= 7791;
                3649: note <= 12187;
                3650: note <= 15286;
                3651: note <= 16283;
                3652: note <= 14886;
                3653: note <= 11395;
                3654: note <= 6627;
                3655: note <= 1697;
                3656: note <= (-2279);
                3657: note <= (-4473);
                3658: note <= (-4563);
                3659: note <= (-2814);
                3660: note <= 0;
                3661: note <= 2814;
                3662: note <= 4563;
                3663: note <= 4473;
                3664: note <= 2279;
                3665: note <= (-1697);
                3666: note <= (-6627);
                3667: note <= (-11395);
                3668: note <= (-14886);
                3669: note <= (-16283);
                3670: note <= (-15286);
                3671: note <= (-12187);
                3672: note <= (-7791);
                3673: note <= (-3203);
                3674: note <= 467;
                3675: note <= 2399;
                3676: note <= 2279;
                3677: note <= 377;
                3678: note <= (-2531);
                3679: note <= (-5378);
                3680: note <= (-7094);
                3681: note <= (-6910);
                3682: note <= (-4563);
                3683: note <= (-377);
                3684: note <= 4815;
                3685: note <= 9889;
                3686: note <= 13722;
                3687: note <= 15491;
                3688: note <= 14886;
                3689: note <= 12187;
                3690: note <= 8192;
                3691: note <= 3995;
                3692: note <= 697;
                3693: note <= (-893);
                3694: note <= (-467);
                3695: note <= 1697;
                3696: note <= 4815;
                3697: note <= 7815;
                3698: note <= 9626;
                3699: note <= 9474;
                3700: note <= 7094;
                3701: note <= 2814;
                3702: note <= (-2531);
                3703: note <= (-7815);
                3704: note <= (-11910);
                3705: note <= (-13985);
                3706: note <= (-13722);
                3707: note <= (-11395);
                3708: note <= (-7791);
                3709: note <= (-3995);
                3710: note <= (-1098);
                3711: note <= 101;
                3712: note <= (-697);
                3713: note <= (-3203);
                3714: note <= (-6627);
                3715: note <= (-9889);
                3716: note <= (-11910);
                3717: note <= (-11911);
                3718: note <= (-9626);
                3719: note <= (-5378);
                3720: note <= 0;
                3721: note <= 5378;
                3722: note <= 9626;
                3723: note <= 11911;
                3724: note <= 11910;
                3725: note <= 9889;
                3726: note <= 6627;
                3727: note <= 3203;
                3728: note <= 697;
                3729: note <= (-101);
                3730: note <= 1098;
                3731: note <= 3995;
                3732: note <= 7791;
                3733: note <= 11395;
                3734: note <= 13722;
                3735: note <= 13985;
                3736: note <= 11910;
                3737: note <= 7815;
                3738: note <= 2531;
                3739: note <= (-2814);
                3740: note <= (-7094);
                3741: note <= (-9474);
                3742: note <= (-9626);
                3743: note <= (-7815);
                3744: note <= (-4815);
                3745: note <= (-1697);
                3746: note <= 467;
                3747: note <= 893;
                3748: note <= (-697);
                3749: note <= (-3995);
                3750: note <= (-8192);
                3751: note <= (-12187);
                3752: note <= (-14886);
                3753: note <= (-15491);
                3754: note <= (-13722);
                3755: note <= (-9889);
                3756: note <= (-4815);
                3757: note <= 377;
                3758: note <= 4563;
                3759: note <= 6910;
                3760: note <= 7094;
                3761: note <= 5378;
                3762: note <= 2531;
                3763: note <= (-377);
                3764: note <= (-2279);
                3765: note <= (-2399);
                3766: note <= (-467);
                3767: note <= 3203;
                3768: note <= 7791;
                3769: note <= 12187;
                3770: note <= 15286;
                3771: note <= 16283;
                3772: note <= 14886;
                3773: note <= 11395;
                3774: note <= 6627;
                3775: note <= 1697;
                3776: note <= (-2279);
                3777: note <= (-4473);
                3778: note <= (-4563);
                3779: note <= (-2814);
                3780: note <= 0;
                3781: note <= 2814;
                3782: note <= 4563;
                3783: note <= 4473;
                3784: note <= 2279;
                3785: note <= (-1697);
                3786: note <= (-6627);
                3787: note <= (-11395);
                3788: note <= (-14886);
                3789: note <= (-16283);
                3790: note <= (-15286);
                3791: note <= (-12187);
                3792: note <= (-7791);
                3793: note <= (-3203);
                3794: note <= 467;
                3795: note <= 2399;
                3796: note <= 2279;
                3797: note <= 377;
                3798: note <= (-2531);
                3799: note <= (-5378);
                3800: note <= (-7094);
                3801: note <= (-6910);
                3802: note <= (-4563);
                3803: note <= (-377);
                3804: note <= 4815;
                3805: note <= 9889;
                3806: note <= 13722;
                3807: note <= 15491;
                3808: note <= 14886;
                3809: note <= 12187;
                3810: note <= 8192;
                3811: note <= 3995;
                3812: note <= 697;
                3813: note <= (-893);
                3814: note <= (-467);
                3815: note <= 1697;
                3816: note <= 4815;
                3817: note <= 7815;
                3818: note <= 9626;
                3819: note <= 9474;
                3820: note <= 7094;
                3821: note <= 2814;
                3822: note <= (-2531);
                3823: note <= (-7815);
                3824: note <= (-11910);
                3825: note <= (-13985);
                3826: note <= (-13722);
                3827: note <= (-11395);
                3828: note <= (-7791);
                3829: note <= (-3995);
                3830: note <= (-1098);
                3831: note <= 101;
                3832: note <= (-697);
                3833: note <= (-3203);
                3834: note <= (-6627);
                3835: note <= (-9889);
                3836: note <= (-11910);
                3837: note <= (-11911);
                3838: note <= (-9626);
                3839: note <= (-5378);
                3840: note <= 0;
                3841: note <= 5378;
                3842: note <= 9626;
                3843: note <= 11911;
                3844: note <= 11910;
                3845: note <= 9889;
                3846: note <= 6627;
                3847: note <= 3203;
                3848: note <= 697;
                3849: note <= (-101);
                3850: note <= 1098;
                3851: note <= 3995;
                3852: note <= 7791;
                3853: note <= 11395;
                3854: note <= 13722;
                3855: note <= 13985;
                3856: note <= 11910;
                3857: note <= 7815;
                3858: note <= 2531;
                3859: note <= (-2814);
                3860: note <= (-7094);
                3861: note <= (-9474);
                3862: note <= (-9626);
                3863: note <= (-7815);
                3864: note <= (-4815);
                3865: note <= (-1697);
                3866: note <= 467;
                3867: note <= 893;
                3868: note <= (-697);
                3869: note <= (-3995);
                3870: note <= (-8192);
                3871: note <= (-12187);
                3872: note <= (-14886);
                3873: note <= (-15491);
                3874: note <= (-13722);
                3875: note <= (-9889);
                3876: note <= (-4815);
                3877: note <= 377;
                3878: note <= 4563;
                3879: note <= 6910;
                3880: note <= 7094;
                3881: note <= 5378;
                3882: note <= 2531;
                3883: note <= (-377);
                3884: note <= (-2279);
                3885: note <= (-2399);
                3886: note <= (-467);
                3887: note <= 3203;
                3888: note <= 7791;
                3889: note <= 12187;
                3890: note <= 15286;
                3891: note <= 16283;
                3892: note <= 14886;
                3893: note <= 11395;
                3894: note <= 6627;
                3895: note <= 1697;
                3896: note <= (-2279);
                3897: note <= (-4473);
                3898: note <= (-4563);
                3899: note <= (-2814);
                3900: note <= 0;
                3901: note <= 2814;
                3902: note <= 4563;
                3903: note <= 4473;
                3904: note <= 2279;
                3905: note <= (-1697);
                3906: note <= (-6627);
                3907: note <= (-11395);
                3908: note <= (-14886);
                3909: note <= (-16283);
                3910: note <= (-15286);
                3911: note <= (-12187);
                3912: note <= (-7791);
                3913: note <= (-3203);
                3914: note <= 467;
                3915: note <= 2399;
                3916: note <= 2279;
                3917: note <= 377;
                3918: note <= (-2531);
                3919: note <= (-5378);
                3920: note <= (-7094);
                3921: note <= (-6910);
                3922: note <= (-4563);
                3923: note <= (-377);
                3924: note <= 4815;
                3925: note <= 9889;
                3926: note <= 13722;
                3927: note <= 15491;
                3928: note <= 14886;
                3929: note <= 12187;
                3930: note <= 8192;
                3931: note <= 3995;
                3932: note <= 697;
                3933: note <= (-893);
                3934: note <= (-467);
                3935: note <= 1697;
                3936: note <= 4815;
                3937: note <= 7815;
                3938: note <= 9626;
                3939: note <= 9474;
                3940: note <= 7094;
                3941: note <= 2814;
                3942: note <= (-2531);
                3943: note <= (-7815);
                3944: note <= (-11910);
                3945: note <= (-13985);
                3946: note <= (-13722);
                3947: note <= (-11395);
                3948: note <= (-7791);
                3949: note <= (-3995);
                3950: note <= (-1098);
                3951: note <= 101;
                3952: note <= (-697);
                3953: note <= (-3203);
                3954: note <= (-6627);
                3955: note <= (-9889);
                3956: note <= (-11910);
                3957: note <= (-11911);
                3958: note <= (-9626);
                3959: note <= (-5378);
                3960: note <= 0;
                3961: note <= 5378;
                3962: note <= 9626;
                3963: note <= 11911;
                3964: note <= 11910;
                3965: note <= 9889;
                3966: note <= 6627;
                3967: note <= 3203;
                3968: note <= 697;
                3969: note <= (-101);
                3970: note <= 1098;
                3971: note <= 3995;
                3972: note <= 7791;
                3973: note <= 11395;
                3974: note <= 13722;
                3975: note <= 13985;
                3976: note <= 11910;
                3977: note <= 7815;
                3978: note <= 2531;
                3979: note <= (-2814);
                3980: note <= (-7094);
                3981: note <= (-9474);
                3982: note <= (-9626);
                3983: note <= (-7815);
                3984: note <= (-4815);
                3985: note <= (-1697);
                3986: note <= 467;
                3987: note <= 893;
                3988: note <= (-697);
                3989: note <= (-3995);
                3990: note <= (-8192);
                3991: note <= (-12187);
                3992: note <= (-14886);
                3993: note <= (-15491);
                3994: note <= (-13722);
                3995: note <= (-9889);
                3996: note <= (-4815);
                3997: note <= 377;
                3998: note <= 4563;
                3999: note <= 6910;
                4000: note <= 7094;
                4001: note <= 5378;
                4002: note <= 2531;
                4003: note <= (-377);
                4004: note <= (-2279);
                4005: note <= (-2399);
                4006: note <= (-467);
                4007: note <= 3203;
                4008: note <= 7791;
                4009: note <= 12187;
                4010: note <= 15286;
                4011: note <= 16283;
                4012: note <= 14886;
                4013: note <= 11395;
                4014: note <= 6627;
                4015: note <= 1697;
                4016: note <= (-2279);
                4017: note <= (-4473);
                4018: note <= (-4563);
                4019: note <= (-2814);
                4020: note <= 0;
                4021: note <= 2814;
                4022: note <= 4563;
                4023: note <= 4473;
                4024: note <= 2279;
                4025: note <= (-1697);
                4026: note <= (-6627);
                4027: note <= (-11395);
                4028: note <= (-14886);
                4029: note <= (-16283);
                4030: note <= (-15286);
                4031: note <= (-12187);
                4032: note <= (-7791);
                4033: note <= (-3203);
                4034: note <= 467;
                4035: note <= 2399;
                4036: note <= 2279;
                4037: note <= 377;
                4038: note <= (-2531);
                4039: note <= (-5378);
                4040: note <= (-7094);
                4041: note <= (-6910);
                4042: note <= (-4563);
                4043: note <= (-377);
                4044: note <= 4815;
                4045: note <= 9889;
                4046: note <= 13722;
                4047: note <= 15491;
                4048: note <= 14886;
                4049: note <= 12187;
                4050: note <= 8192;
                4051: note <= 3995;
                4052: note <= 697;
                4053: note <= (-893);
                4054: note <= (-467);
                4055: note <= 1697;
                4056: note <= 4815;
                4057: note <= 7815;
                4058: note <= 9626;
                4059: note <= 9474;
                4060: note <= 7094;
                4061: note <= 2814;
                4062: note <= (-2531);
                4063: note <= (-7815);
                4064: note <= (-11910);
                4065: note <= (-13985);
                4066: note <= (-13722);
                4067: note <= (-11395);
                4068: note <= (-7791);
                4069: note <= (-3995);
                4070: note <= (-1098);
                4071: note <= 101;
                4072: note <= (-697);
                4073: note <= (-3203);
                4074: note <= (-6627);
                4075: note <= (-9889);
                4076: note <= (-11910);
                4077: note <= (-11911);
                4078: note <= (-9626);
                4079: note <= (-5378);
                4080: note <= 0;
                4081: note <= 5378;
                4082: note <= 9626;
                4083: note <= 11911;
                4084: note <= 11910;
                4085: note <= 9889;
                4086: note <= 6627;
                4087: note <= 3203;
                4088: note <= 697;
                4089: note <= (-101);
                4090: note <= 1098;
                4091: note <= 3995;
                4092: note <= 7791;
                4093: note <= 11395;
                4094: note <= 13722;
                4095: note <= 13985;
                4096: note <= 11910;
                4097: note <= 7815;
                4098: note <= 2531;
                4099: note <= (-2814);
                4100: note <= (-7094);
                4101: note <= (-9474);
                4102: note <= (-9626);
                4103: note <= (-7815);
                4104: note <= (-4815);
                4105: note <= (-1697);
                4106: note <= 467;
                4107: note <= 893;
                4108: note <= (-697);
                4109: note <= (-3995);
                4110: note <= (-8192);
                4111: note <= (-12187);
                4112: note <= (-14886);
                4113: note <= (-15491);
                4114: note <= (-13722);
                4115: note <= (-9889);
                4116: note <= (-4815);
                4117: note <= 377;
                4118: note <= 4563;
                4119: note <= 6910;
                4120: note <= 7094;
                4121: note <= 5378;
                4122: note <= 2531;
                4123: note <= (-377);
                4124: note <= (-2279);
                4125: note <= (-2399);
                4126: note <= (-467);
                4127: note <= 3203;
                4128: note <= 7791;
                4129: note <= 12187;
                4130: note <= 15286;
                4131: note <= 16283;
                4132: note <= 14886;
                4133: note <= 11395;
                4134: note <= 6627;
                4135: note <= 1697;
                4136: note <= (-2279);
                4137: note <= (-4473);
                4138: note <= (-4563);
                4139: note <= (-2814);
                4140: note <= 0;
                4141: note <= 2814;
                4142: note <= 4563;
                4143: note <= 4473;
                4144: note <= 2279;
                4145: note <= (-1697);
                4146: note <= (-6627);
                4147: note <= (-11395);
                4148: note <= (-14886);
                4149: note <= (-16283);
                4150: note <= (-15286);
                4151: note <= (-12187);
                4152: note <= (-7791);
                4153: note <= (-3203);
                4154: note <= 467;
                4155: note <= 2399;
                4156: note <= 2279;
                4157: note <= 377;
                4158: note <= (-2531);
                4159: note <= (-5378);
                4160: note <= (-7094);
                4161: note <= (-6910);
                4162: note <= (-4563);
                4163: note <= (-377);
                4164: note <= 4815;
                4165: note <= 9889;
                4166: note <= 13722;
                4167: note <= 15491;
                4168: note <= 14886;
                4169: note <= 12187;
                4170: note <= 8192;
                4171: note <= 3995;
                4172: note <= 697;
                4173: note <= (-893);
                4174: note <= (-467);
                4175: note <= 1697;
                4176: note <= 4815;
                4177: note <= 7815;
                4178: note <= 9626;
                4179: note <= 9474;
                4180: note <= 7094;
                4181: note <= 2814;
                4182: note <= (-2531);
                4183: note <= (-7815);
                4184: note <= (-11910);
                4185: note <= (-13985);
                4186: note <= (-13722);
                4187: note <= (-11395);
                4188: note <= (-7791);
                4189: note <= (-3995);
                4190: note <= (-1098);
                4191: note <= 101;
                4192: note <= (-697);
                4193: note <= (-3203);
                4194: note <= (-6627);
                4195: note <= (-9889);
                4196: note <= (-11910);
                4197: note <= (-11911);
                4198: note <= (-9626);
                4199: note <= (-5378);
                4200: note <= 0;
                4201: note <= 5378;
                4202: note <= 9626;
                4203: note <= 11911;
                4204: note <= 11910;
                4205: note <= 9889;
                4206: note <= 6627;
                4207: note <= 3203;
                4208: note <= 697;
                4209: note <= (-101);
                4210: note <= 1098;
                4211: note <= 3995;
                4212: note <= 7791;
                4213: note <= 11395;
                4214: note <= 13722;
                4215: note <= 13985;
                4216: note <= 11910;
                4217: note <= 7815;
                4218: note <= 2531;
                4219: note <= (-2814);
                4220: note <= (-7094);
                4221: note <= (-9474);
                4222: note <= (-9626);
                4223: note <= (-7815);
                4224: note <= (-4815);
                4225: note <= (-1697);
                4226: note <= 467;
                4227: note <= 893;
                4228: note <= (-697);
                4229: note <= (-3995);
                4230: note <= (-8192);
                4231: note <= (-12187);
                4232: note <= (-14886);
                4233: note <= (-15491);
                4234: note <= (-13722);
                4235: note <= (-9889);
                4236: note <= (-4815);
                4237: note <= 377;
                4238: note <= 4563;
                4239: note <= 6910;
                4240: note <= 7094;
                4241: note <= 5378;
                4242: note <= 2531;
                4243: note <= (-377);
                4244: note <= (-2279);
                4245: note <= (-2399);
                4246: note <= (-467);
                4247: note <= 3203;
                4248: note <= 7791;
                4249: note <= 12187;
                4250: note <= 15286;
                4251: note <= 16283;
                4252: note <= 14886;
                4253: note <= 11395;
                4254: note <= 6627;
                4255: note <= 1697;
                4256: note <= (-2279);
                4257: note <= (-4473);
                4258: note <= (-4563);
                4259: note <= (-2814);
                4260: note <= 0;
                4261: note <= 2814;
                4262: note <= 4563;
                4263: note <= 4473;
                4264: note <= 2279;
                4265: note <= (-1697);
                4266: note <= (-6627);
                4267: note <= (-11395);
                4268: note <= (-14886);
                4269: note <= (-16283);
                4270: note <= (-15286);
                4271: note <= (-12187);
                4272: note <= (-7791);
                4273: note <= (-3203);
                4274: note <= 467;
                4275: note <= 2399;
                4276: note <= 2279;
                4277: note <= 377;
                4278: note <= (-2531);
                4279: note <= (-5378);
                4280: note <= (-7094);
                4281: note <= (-6910);
                4282: note <= (-4563);
                4283: note <= (-377);
                4284: note <= 4815;
                4285: note <= 9889;
                4286: note <= 13722;
                4287: note <= 15491;
                4288: note <= 14886;
                4289: note <= 12187;
                4290: note <= 8192;
                4291: note <= 3995;
                4292: note <= 697;
                4293: note <= (-893);
                4294: note <= (-467);
                4295: note <= 1697;
                4296: note <= 4815;
                4297: note <= 7815;
                4298: note <= 9626;
                4299: note <= 9474;
                4300: note <= 7094;
                4301: note <= 2814;
                4302: note <= (-2531);
                4303: note <= (-7815);
                4304: note <= (-11910);
                4305: note <= (-13985);
                4306: note <= (-13722);
                4307: note <= (-11395);
                4308: note <= (-7791);
                4309: note <= (-3995);
                4310: note <= (-1098);
                4311: note <= 101;
                4312: note <= (-697);
                4313: note <= (-3203);
                4314: note <= (-6627);
                4315: note <= (-9889);
                4316: note <= (-11910);
                4317: note <= (-11911);
                4318: note <= (-9626);
                4319: note <= (-5378);
                4320: note <= 0;
                4321: note <= 5378;
                4322: note <= 9626;
                4323: note <= 11911;
                4324: note <= 11910;
                4325: note <= 9889;
                4326: note <= 6627;
                4327: note <= 3203;
                4328: note <= 697;
                4329: note <= (-101);
                4330: note <= 1098;
                4331: note <= 3995;
                4332: note <= 7791;
                4333: note <= 11395;
                4334: note <= 13722;
                4335: note <= 13985;
                4336: note <= 11910;
                4337: note <= 7815;
                4338: note <= 2531;
                4339: note <= (-2814);
                4340: note <= (-7094);
                4341: note <= (-9474);
                4342: note <= (-9626);
                4343: note <= (-7815);
                4344: note <= (-4815);
                4345: note <= (-1697);
                4346: note <= 467;
                4347: note <= 893;
                4348: note <= (-697);
                4349: note <= (-3995);
                4350: note <= (-8192);
                4351: note <= (-12187);
                4352: note <= (-14886);
                4353: note <= (-15491);
                4354: note <= (-13722);
                4355: note <= (-9889);
                4356: note <= (-4815);
                4357: note <= 377;
                4358: note <= 4563;
                4359: note <= 6910;
                4360: note <= 7094;
                4361: note <= 5378;
                4362: note <= 2531;
                4363: note <= (-377);
                4364: note <= (-2279);
                4365: note <= (-2399);
                4366: note <= (-467);
                4367: note <= 3203;
                4368: note <= 7791;
                4369: note <= 12187;
                4370: note <= 15286;
                4371: note <= 16283;
                4372: note <= 14886;
                4373: note <= 11395;
                4374: note <= 6627;
                4375: note <= 1697;
                4376: note <= (-2279);
                4377: note <= (-4473);
                4378: note <= (-4563);
                4379: note <= (-2814);
                4380: note <= 0;
                4381: note <= 2814;
                4382: note <= 4563;
                4383: note <= 4473;
                4384: note <= 2279;
                4385: note <= (-1697);
                4386: note <= (-6627);
                4387: note <= (-11395);
                4388: note <= (-14886);
                4389: note <= (-16283);
                4390: note <= (-15286);
                4391: note <= (-12187);
                4392: note <= (-7791);
                4393: note <= (-3203);
                4394: note <= 467;
                4395: note <= 2399;
                4396: note <= 2279;
                4397: note <= 377;
                4398: note <= (-2531);
                4399: note <= (-5378);
                4400: note <= (-7094);
                4401: note <= (-6910);
                4402: note <= (-4563);
                4403: note <= (-377);
                4404: note <= 4815;
                4405: note <= 9889;
                4406: note <= 13722;
                4407: note <= 15491;
                4408: note <= 14886;
                4409: note <= 12187;
                4410: note <= 8192;
                4411: note <= 3995;
                4412: note <= 697;
                4413: note <= (-893);
                4414: note <= (-467);
                4415: note <= 1697;
                4416: note <= 4815;
                4417: note <= 7815;
                4418: note <= 9626;
                4419: note <= 9474;
                4420: note <= 7094;
                4421: note <= 2814;
                4422: note <= (-2531);
                4423: note <= (-7815);
                4424: note <= (-11910);
                4425: note <= (-13985);
                4426: note <= (-13722);
                4427: note <= (-11395);
                4428: note <= (-7791);
                4429: note <= (-3995);
                4430: note <= (-1098);
                4431: note <= 101;
                4432: note <= (-697);
                4433: note <= (-3203);
                4434: note <= (-6627);
                4435: note <= (-9889);
                4436: note <= (-11910);
                4437: note <= (-11911);
                4438: note <= (-9626);
                4439: note <= (-5378);
                4440: note <= 0;
                4441: note <= 5378;
                4442: note <= 9626;
                4443: note <= 11911;
                4444: note <= 11910;
                4445: note <= 9889;
                4446: note <= 6627;
                4447: note <= 3203;
                4448: note <= 697;
                4449: note <= (-101);
                4450: note <= 1098;
                4451: note <= 3995;
                4452: note <= 7791;
                4453: note <= 11395;
                4454: note <= 13722;
                4455: note <= 13985;
                4456: note <= 11910;
                4457: note <= 7815;
                4458: note <= 2531;
                4459: note <= (-2814);
                4460: note <= (-7094);
                4461: note <= (-9474);
                4462: note <= (-9626);
                4463: note <= (-7815);
                4464: note <= (-4815);
                4465: note <= (-1697);
                4466: note <= 467;
                4467: note <= 893;
                4468: note <= (-697);
                4469: note <= (-3995);
                4470: note <= (-8192);
                4471: note <= (-12187);
                4472: note <= (-14886);
                4473: note <= (-15491);
                4474: note <= (-13722);
                4475: note <= (-9889);
                4476: note <= (-4815);
                4477: note <= 377;
                4478: note <= 4563;
                4479: note <= 6910;
                4480: note <= 7094;
                4481: note <= 5378;
                4482: note <= 2531;
                4483: note <= (-377);
                4484: note <= (-2279);
                4485: note <= (-2399);
                4486: note <= (-467);
                4487: note <= 3203;
                4488: note <= 7791;
                4489: note <= 12187;
                4490: note <= 15286;
                4491: note <= 16283;
                4492: note <= 14886;
                4493: note <= 11395;
                4494: note <= 6627;
                4495: note <= 1697;
                4496: note <= (-2279);
                4497: note <= (-4473);
                4498: note <= (-4563);
                4499: note <= (-2814);
                4500: note <= 0;
                4501: note <= 2814;
                4502: note <= 4563;
                4503: note <= 4473;
                4504: note <= 2279;
                4505: note <= (-1697);
                4506: note <= (-6627);
                4507: note <= (-11395);
                4508: note <= (-14886);
                4509: note <= (-16283);
                4510: note <= (-15286);
                4511: note <= (-12187);
                4512: note <= (-7791);
                4513: note <= (-3203);
                4514: note <= 467;
                4515: note <= 2399;
                4516: note <= 2279;
                4517: note <= 377;
                4518: note <= (-2531);
                4519: note <= (-5378);
                4520: note <= (-7094);
                4521: note <= (-6910);
                4522: note <= (-4563);
                4523: note <= (-377);
                4524: note <= 4815;
                4525: note <= 9889;
                4526: note <= 13722;
                4527: note <= 15491;
                4528: note <= 14886;
                4529: note <= 12187;
                4530: note <= 8192;
                4531: note <= 3995;
                4532: note <= 697;
                4533: note <= (-893);
                4534: note <= (-467);
                4535: note <= 1697;
                4536: note <= 4815;
                4537: note <= 7815;
                4538: note <= 9626;
                4539: note <= 9474;
                4540: note <= 7094;
                4541: note <= 2814;
                4542: note <= (-2531);
                4543: note <= (-7815);
                4544: note <= (-11910);
                4545: note <= (-13985);
                4546: note <= (-13722);
                4547: note <= (-11395);
                4548: note <= (-7791);
                4549: note <= (-3995);
                4550: note <= (-1098);
                4551: note <= 101;
                4552: note <= (-697);
                4553: note <= (-3203);
                4554: note <= (-6627);
                4555: note <= (-9889);
                4556: note <= (-11910);
                4557: note <= (-11911);
                4558: note <= (-9626);
                4559: note <= (-5378);
                4560: note <= 0;
                4561: note <= 5378;
                4562: note <= 9626;
                4563: note <= 11911;
                4564: note <= 11910;
                4565: note <= 9889;
                4566: note <= 6627;
                4567: note <= 3203;
                4568: note <= 697;
                4569: note <= (-101);
                4570: note <= 1098;
                4571: note <= 3995;
                4572: note <= 7791;
                4573: note <= 11395;
                4574: note <= 13722;
                4575: note <= 13985;
                4576: note <= 11910;
                4577: note <= 7815;
                4578: note <= 2531;
                4579: note <= (-2814);
                4580: note <= (-7094);
                4581: note <= (-9474);
                4582: note <= (-9626);
                4583: note <= (-7815);
                4584: note <= (-4815);
                4585: note <= (-1697);
                4586: note <= 467;
                4587: note <= 893;
                4588: note <= (-697);
                4589: note <= (-3995);
                4590: note <= (-8192);
                4591: note <= (-12187);
                4592: note <= (-14886);
                4593: note <= (-15491);
                4594: note <= (-13722);
                4595: note <= (-9889);
                4596: note <= (-4815);
                4597: note <= 377;
                4598: note <= 4563;
                4599: note <= 6910;
                4600: note <= 7094;
                4601: note <= 5378;
                4602: note <= 2531;
                4603: note <= (-377);
                4604: note <= (-2279);
                4605: note <= (-2399);
                4606: note <= (-467);
                4607: note <= 3203;
                4608: note <= 7791;
                4609: note <= 12187;
                4610: note <= 15286;
                4611: note <= 16283;
                4612: note <= 14886;
                4613: note <= 11395;
                4614: note <= 6627;
                4615: note <= 1697;
                4616: note <= (-2279);
                4617: note <= (-4473);
                4618: note <= (-4563);
                4619: note <= (-2814);
                4620: note <= 0;
                4621: note <= 2814;
                4622: note <= 4563;
                4623: note <= 4473;
                4624: note <= 2279;
                4625: note <= (-1697);
                4626: note <= (-6627);
                4627: note <= (-11395);
                4628: note <= (-14886);
                4629: note <= (-16283);
                4630: note <= (-15286);
                4631: note <= (-12187);
                4632: note <= (-7791);
                4633: note <= (-3203);
                4634: note <= 467;
                4635: note <= 2399;
                4636: note <= 2279;
                4637: note <= 377;
                4638: note <= (-2531);
                4639: note <= (-5378);
                4640: note <= (-7094);
                4641: note <= (-6910);
                4642: note <= (-4563);
                4643: note <= (-377);
                4644: note <= 4815;
                4645: note <= 9889;
                4646: note <= 13722;
                4647: note <= 15491;
                4648: note <= 14886;
                4649: note <= 12187;
                4650: note <= 8192;
                4651: note <= 3995;
                4652: note <= 697;
                4653: note <= (-893);
                4654: note <= (-467);
                4655: note <= 1697;
                4656: note <= 4815;
                4657: note <= 7815;
                4658: note <= 9626;
                4659: note <= 9474;
                4660: note <= 7094;
                4661: note <= 2814;
                4662: note <= (-2531);
                4663: note <= (-7815);
                4664: note <= (-11910);
                4665: note <= (-13985);
                4666: note <= (-13722);
                4667: note <= (-11395);
                4668: note <= (-7791);
                4669: note <= (-3995);
                4670: note <= (-1098);
                4671: note <= 101;
                4672: note <= (-697);
                4673: note <= (-3203);
                4674: note <= (-6627);
                4675: note <= (-9889);
                4676: note <= (-11910);
                4677: note <= (-11911);
                4678: note <= (-9626);
                4679: note <= (-5378);
                4680: note <= 0;
                4681: note <= 5378;
                4682: note <= 9626;
                4683: note <= 11911;
                4684: note <= 11910;
                4685: note <= 9889;
                4686: note <= 6627;
                4687: note <= 3203;
                4688: note <= 697;
                4689: note <= (-101);
                4690: note <= 1098;
                4691: note <= 3995;
                4692: note <= 7791;
                4693: note <= 11395;
                4694: note <= 13722;
                4695: note <= 13985;
                4696: note <= 11910;
                4697: note <= 7815;
                4698: note <= 2531;
                4699: note <= (-2814);
                4700: note <= (-7094);
                4701: note <= (-9474);
                4702: note <= (-9626);
                4703: note <= (-7815);
                4704: note <= (-4815);
                4705: note <= (-1697);
                4706: note <= 467;
                4707: note <= 893;
                4708: note <= (-697);
                4709: note <= (-3995);
                4710: note <= (-8192);
                4711: note <= (-12187);
                4712: note <= (-14886);
                4713: note <= (-15491);
                4714: note <= (-13722);
                4715: note <= (-9889);
                4716: note <= (-4815);
                4717: note <= 377;
                4718: note <= 4563;
                4719: note <= 6910;
                4720: note <= 7094;
                4721: note <= 5378;
                4722: note <= 2531;
                4723: note <= (-377);
                4724: note <= (-2279);
                4725: note <= (-2399);
                4726: note <= (-467);
                4727: note <= 3203;
                4728: note <= 7791;
                4729: note <= 12187;
                4730: note <= 15286;
                4731: note <= 16283;
                4732: note <= 14886;
                4733: note <= 11395;
                4734: note <= 6627;
                4735: note <= 1697;
                4736: note <= (-2279);
                4737: note <= (-4473);
                4738: note <= (-4563);
                4739: note <= (-2814);
                4740: note <= 0;
                4741: note <= 2814;
                4742: note <= 4563;
                4743: note <= 4473;
                4744: note <= 2279;
                4745: note <= (-1697);
                4746: note <= (-6627);
                4747: note <= (-11395);
                4748: note <= (-14886);
                4749: note <= (-16283);
                4750: note <= (-15286);
                4751: note <= (-12187);
                4752: note <= (-7791);
                4753: note <= (-3203);
                4754: note <= 467;
                4755: note <= 2399;
                4756: note <= 2279;
                4757: note <= 377;
                4758: note <= (-2531);
                4759: note <= (-5378);
                4760: note <= (-7094);
                4761: note <= (-6910);
                4762: note <= (-4563);
                4763: note <= (-377);
                4764: note <= 4815;
                4765: note <= 9889;
                4766: note <= 13722;
                4767: note <= 15491;
                4768: note <= 14886;
                4769: note <= 12187;
                4770: note <= 8192;
                4771: note <= 3995;
                4772: note <= 697;
                4773: note <= (-893);
                4774: note <= (-467);
                4775: note <= 1697;
                4776: note <= 4815;
                4777: note <= 7815;
                4778: note <= 9626;
                4779: note <= 9474;
                4780: note <= 7094;
                4781: note <= 2814;
                4782: note <= (-2531);
                4783: note <= (-7815);
                4784: note <= (-11910);
                4785: note <= (-13985);
                4786: note <= (-13722);
                4787: note <= (-11395);
                4788: note <= (-7791);
                4789: note <= (-3995);
                4790: note <= (-1098);
                4791: note <= 101;
                4792: note <= (-697);
                4793: note <= (-3203);
                4794: note <= (-6627);
                4795: note <= (-9889);
                4796: note <= (-11910);
                4797: note <= (-11911);
                4798: note <= (-9626);
                4799: note <= (-5378);
                4800: note <= 0;
                4801: note <= 5378;
                4802: note <= 9626;
                4803: note <= 11911;
                4804: note <= 11910;
                4805: note <= 9889;
                4806: note <= 6627;
                4807: note <= 3203;
                4808: note <= 697;
                4809: note <= (-101);
                4810: note <= 1098;
                4811: note <= 3995;
                4812: note <= 7791;
                4813: note <= 11395;
                4814: note <= 13722;
                4815: note <= 13985;
                4816: note <= 11910;
                4817: note <= 7815;
                4818: note <= 2531;
                4819: note <= (-2814);
                4820: note <= (-7094);
                4821: note <= (-9474);
                4822: note <= (-9626);
                4823: note <= (-7815);
                4824: note <= (-4815);
                4825: note <= (-1697);
                4826: note <= 467;
                4827: note <= 893;
                4828: note <= (-697);
                4829: note <= (-3995);
                4830: note <= (-8192);
                4831: note <= (-12187);
                4832: note <= (-14886);
                4833: note <= (-15491);
                4834: note <= (-13722);
                4835: note <= (-9889);
                4836: note <= (-4815);
                4837: note <= 377;
                4838: note <= 4563;
                4839: note <= 6910;
                4840: note <= 7094;
                4841: note <= 5378;
                4842: note <= 2531;
                4843: note <= (-377);
                4844: note <= (-2279);
                4845: note <= (-2399);
                4846: note <= (-467);
                4847: note <= 3203;
                4848: note <= 7791;
                4849: note <= 12187;
                4850: note <= 15286;
                4851: note <= 16283;
                4852: note <= 14886;
                4853: note <= 11395;
                4854: note <= 6627;
                4855: note <= 1697;
                4856: note <= (-2279);
                4857: note <= (-4473);
                4858: note <= (-4563);
                4859: note <= (-2814);
                4860: note <= 0;
                4861: note <= 2814;
                4862: note <= 4563;
                4863: note <= 4473;
                4864: note <= 2279;
                4865: note <= (-1697);
                4866: note <= (-6627);
                4867: note <= (-11395);
                4868: note <= (-14886);
                4869: note <= (-16283);
                4870: note <= (-15286);
                4871: note <= (-12187);
                4872: note <= (-7791);
                4873: note <= (-3203);
                4874: note <= 467;
                4875: note <= 2399;
                4876: note <= 2279;
                4877: note <= 377;
                4878: note <= (-2531);
                4879: note <= (-5378);
                4880: note <= (-7094);
                4881: note <= (-6910);
                4882: note <= (-4563);
                4883: note <= (-377);
                4884: note <= 4815;
                4885: note <= 9889;
                4886: note <= 13722;
                4887: note <= 15491;
                4888: note <= 14886;
                4889: note <= 12187;
                4890: note <= 8192;
                4891: note <= 3995;
                4892: note <= 697;
                4893: note <= (-893);
                4894: note <= (-467);
                4895: note <= 1697;
                4896: note <= 4815;
                4897: note <= 7815;
                4898: note <= 9626;
                4899: note <= 9474;
                4900: note <= 7094;
                4901: note <= 2814;
                4902: note <= (-2531);
                4903: note <= (-7815);
                4904: note <= (-11910);
                4905: note <= (-13985);
                4906: note <= (-13722);
                4907: note <= (-11395);
                4908: note <= (-7791);
                4909: note <= (-3995);
                4910: note <= (-1098);
                4911: note <= 101;
                4912: note <= (-697);
                4913: note <= (-3203);
                4914: note <= (-6627);
                4915: note <= (-9889);
                4916: note <= (-11910);
                4917: note <= (-11911);
                4918: note <= (-9626);
                4919: note <= (-5378);
                4920: note <= 0;
                4921: note <= 5378;
                4922: note <= 9626;
                4923: note <= 11911;
                4924: note <= 11910;
                4925: note <= 9889;
                4926: note <= 6627;
                4927: note <= 3203;
                4928: note <= 697;
                4929: note <= (-101);
                4930: note <= 1098;
                4931: note <= 3995;
                4932: note <= 7791;
                4933: note <= 11395;
                4934: note <= 13722;
                4935: note <= 13985;
                4936: note <= 11910;
                4937: note <= 7815;
                4938: note <= 2531;
                4939: note <= (-2814);
                4940: note <= (-7094);
                4941: note <= (-9474);
                4942: note <= (-9626);
                4943: note <= (-7815);
                4944: note <= (-4815);
                4945: note <= (-1697);
                4946: note <= 467;
                4947: note <= 893;
                4948: note <= (-697);
                4949: note <= (-3995);
                4950: note <= (-8192);
                4951: note <= (-12187);
                4952: note <= (-14886);
                4953: note <= (-15491);
                4954: note <= (-13722);
                4955: note <= (-9889);
                4956: note <= (-4815);
                4957: note <= 377;
                4958: note <= 4563;
                4959: note <= 6910;
                4960: note <= 7094;
                4961: note <= 5378;
                4962: note <= 2531;
                4963: note <= (-377);
                4964: note <= (-2279);
                4965: note <= (-2399);
                4966: note <= (-467);
                4967: note <= 3203;
                4968: note <= 7791;
                4969: note <= 12187;
                4970: note <= 15286;
                4971: note <= 16283;
                4972: note <= 14886;
                4973: note <= 11395;
                4974: note <= 6627;
                4975: note <= 1697;
                4976: note <= (-2279);
                4977: note <= (-4473);
                4978: note <= (-4563);
                4979: note <= (-2814);
                4980: note <= 0;
                4981: note <= 2814;
                4982: note <= 4563;
                4983: note <= 4473;
                4984: note <= 2279;
                4985: note <= (-1697);
                4986: note <= (-6627);
                4987: note <= (-11395);
                4988: note <= (-14886);
                4989: note <= (-16283);
                4990: note <= (-15286);
                4991: note <= (-12187);
                4992: note <= (-7791);
                4993: note <= (-3203);
                4994: note <= 467;
                4995: note <= 2399;
                4996: note <= 2279;
                4997: note <= 377;
                4998: note <= (-2531);
                4999: note <= (-5378);
                5000: note <= (-7094);
                5001: note <= (-6910);
                5002: note <= (-4563);
                5003: note <= (-377);
                5004: note <= 4815;
                5005: note <= 9889;
                5006: note <= 13722;
                5007: note <= 15491;
                5008: note <= 14886;
                5009: note <= 12187;
                5010: note <= 8192;
                5011: note <= 3995;
                5012: note <= 697;
                5013: note <= (-893);
                5014: note <= (-467);
                5015: note <= 1697;
                5016: note <= 4815;
                5017: note <= 7815;
                5018: note <= 9626;
                5019: note <= 9474;
                5020: note <= 7094;
                5021: note <= 2814;
                5022: note <= (-2531);
                5023: note <= (-7815);
                5024: note <= (-11910);
                5025: note <= (-13985);
                5026: note <= (-13722);
                5027: note <= (-11395);
                5028: note <= (-7791);
                5029: note <= (-3995);
                5030: note <= (-1098);
                5031: note <= 101;
                5032: note <= (-697);
                5033: note <= (-3203);
                5034: note <= (-6627);
                5035: note <= (-9889);
                5036: note <= (-11910);
                5037: note <= (-11911);
                5038: note <= (-9626);
                5039: note <= (-5378);
                5040: note <= 0;
                5041: note <= 5378;
                5042: note <= 9626;
                5043: note <= 11911;
                5044: note <= 11910;
                5045: note <= 9889;
                5046: note <= 6627;
                5047: note <= 3203;
                5048: note <= 697;
                5049: note <= (-101);
                5050: note <= 1098;
                5051: note <= 3995;
                5052: note <= 7791;
                5053: note <= 11395;
                5054: note <= 13722;
                5055: note <= 13985;
                5056: note <= 11910;
                5057: note <= 7815;
                5058: note <= 2531;
                5059: note <= (-2814);
                5060: note <= (-7094);
                5061: note <= (-9474);
                5062: note <= (-9626);
                5063: note <= (-7815);
                5064: note <= (-4815);
                5065: note <= (-1697);
                5066: note <= 467;
                5067: note <= 893;
                5068: note <= (-697);
                5069: note <= (-3995);
                5070: note <= (-8192);
                5071: note <= (-12187);
                5072: note <= (-14886);
                5073: note <= (-15491);
                5074: note <= (-13722);
                5075: note <= (-9889);
                5076: note <= (-4815);
                5077: note <= 377;
                5078: note <= 4563;
                5079: note <= 6910;
                5080: note <= 7094;
                5081: note <= 5378;
                5082: note <= 2531;
                5083: note <= (-377);
                5084: note <= (-2279);
                5085: note <= (-2399);
                5086: note <= (-467);
                5087: note <= 3203;
                5088: note <= 7791;
                5089: note <= 12187;
                5090: note <= 15286;
                5091: note <= 16283;
                5092: note <= 14886;
                5093: note <= 11395;
                5094: note <= 6627;
                5095: note <= 1697;
                5096: note <= (-2279);
                5097: note <= (-4473);
                5098: note <= (-4563);
                5099: note <= (-2814);
                5100: note <= 0;
                5101: note <= 2814;
                5102: note <= 4563;
                5103: note <= 4473;
                5104: note <= 2279;
                5105: note <= (-1697);
                5106: note <= (-6627);
                5107: note <= (-11395);
                5108: note <= (-14886);
                5109: note <= (-16283);
                5110: note <= (-15286);
                5111: note <= (-12187);
                5112: note <= (-7791);
                5113: note <= (-3203);
                5114: note <= 467;
                5115: note <= 2399;
                5116: note <= 2279;
                5117: note <= 377;
                5118: note <= (-2531);
                5119: note <= (-5378);
                5120: note <= (-7094);
                5121: note <= (-6910);
                5122: note <= (-4563);
                5123: note <= (-377);
                5124: note <= 4815;
                5125: note <= 9889;
                5126: note <= 13722;
                5127: note <= 15491;
                5128: note <= 14886;
                5129: note <= 12187;
                5130: note <= 8192;
                5131: note <= 3995;
                5132: note <= 697;
                5133: note <= (-893);
                5134: note <= (-467);
                5135: note <= 1697;
                5136: note <= 4815;
                5137: note <= 7815;
                5138: note <= 9626;
                5139: note <= 9474;
                5140: note <= 7094;
                5141: note <= 2814;
                5142: note <= (-2531);
                5143: note <= (-7815);
                5144: note <= (-11910);
                5145: note <= (-13985);
                5146: note <= (-13722);
                5147: note <= (-11395);
                5148: note <= (-7791);
                5149: note <= (-3995);
                5150: note <= (-1098);
                5151: note <= 101;
                5152: note <= (-697);
                5153: note <= (-3203);
                5154: note <= (-6627);
                5155: note <= (-9889);
                5156: note <= (-11910);
                5157: note <= (-11911);
                5158: note <= (-9626);
                5159: note <= (-5378);
                5160: note <= 0;
                5161: note <= 5378;
                5162: note <= 9626;
                5163: note <= 11911;
                5164: note <= 11910;
                5165: note <= 9889;
                5166: note <= 6627;
                5167: note <= 3203;
                5168: note <= 697;
                5169: note <= (-101);
                5170: note <= 1098;
                5171: note <= 3995;
                5172: note <= 7791;
                5173: note <= 11395;
                5174: note <= 13722;
                5175: note <= 13985;
                5176: note <= 11910;
                5177: note <= 7815;
                5178: note <= 2531;
                5179: note <= (-2814);
                5180: note <= (-7094);
                5181: note <= (-9474);
                5182: note <= (-9626);
                5183: note <= (-7815);
                5184: note <= (-4815);
                5185: note <= (-1697);
                5186: note <= 467;
                5187: note <= 893;
                5188: note <= (-697);
                5189: note <= (-3995);
                5190: note <= (-8192);
                5191: note <= (-12187);
                5192: note <= (-14886);
                5193: note <= (-15491);
                5194: note <= (-13722);
                5195: note <= (-9889);
                5196: note <= (-4815);
                5197: note <= 377;
                5198: note <= 4563;
                5199: note <= 6910;
                5200: note <= 7094;
                5201: note <= 5378;
                5202: note <= 2531;
                5203: note <= (-377);
                5204: note <= (-2279);
                5205: note <= (-2399);
                5206: note <= (-467);
                5207: note <= 3203;
                5208: note <= 7791;
                5209: note <= 12187;
                5210: note <= 15286;
                5211: note <= 16283;
                5212: note <= 14886;
                5213: note <= 11395;
                5214: note <= 6627;
                5215: note <= 1697;
                5216: note <= (-2279);
                5217: note <= (-4473);
                5218: note <= (-4563);
                5219: note <= (-2814);
                5220: note <= 0;
                5221: note <= 2814;
                5222: note <= 4563;
                5223: note <= 4473;
                5224: note <= 2279;
                5225: note <= (-1697);
                5226: note <= (-6627);
                5227: note <= (-11395);
                5228: note <= (-14886);
                5229: note <= (-16283);
                5230: note <= (-15286);
                5231: note <= (-12187);
                5232: note <= (-7791);
                5233: note <= (-3203);
                5234: note <= 467;
                5235: note <= 2399;
                5236: note <= 2279;
                5237: note <= 377;
                5238: note <= (-2531);
                5239: note <= (-5378);
                5240: note <= (-7094);
                5241: note <= (-6910);
                5242: note <= (-4563);
                5243: note <= (-377);
                5244: note <= 4815;
                5245: note <= 9889;
                5246: note <= 13722;
                5247: note <= 15491;
                5248: note <= 14886;
                5249: note <= 12187;
                5250: note <= 8192;
                5251: note <= 3995;
                5252: note <= 697;
                5253: note <= (-893);
                5254: note <= (-467);
                5255: note <= 1697;
                5256: note <= 4815;
                5257: note <= 7815;
                5258: note <= 9626;
                5259: note <= 9474;
                5260: note <= 7094;
                5261: note <= 2814;
                5262: note <= (-2531);
                5263: note <= (-7815);
                5264: note <= (-11910);
                5265: note <= (-13985);
                5266: note <= (-13722);
                5267: note <= (-11395);
                5268: note <= (-7791);
                5269: note <= (-3995);
                5270: note <= (-1098);
                5271: note <= 101;
                5272: note <= (-697);
                5273: note <= (-3203);
                5274: note <= (-6627);
                5275: note <= (-9889);
                5276: note <= (-11910);
                5277: note <= (-11911);
                5278: note <= (-9626);
                5279: note <= (-5378);
                5280: note <= 0;
                5281: note <= 5378;
                5282: note <= 9626;
                5283: note <= 11911;
                5284: note <= 11910;
                5285: note <= 9889;
                5286: note <= 6627;
                5287: note <= 3203;
                5288: note <= 697;
                5289: note <= (-101);
                5290: note <= 1098;
                5291: note <= 3995;
                5292: note <= 7791;
                5293: note <= 11395;
                5294: note <= 13722;
                5295: note <= 13985;
                5296: note <= 11910;
                5297: note <= 7815;
                5298: note <= 2531;
                5299: note <= (-2814);
                5300: note <= (-7094);
                5301: note <= (-9474);
                5302: note <= (-9626);
                5303: note <= (-7815);
                5304: note <= (-4815);
                5305: note <= (-1697);
                5306: note <= 467;
                5307: note <= 893;
                5308: note <= (-697);
                5309: note <= (-3995);
                5310: note <= (-8192);
                5311: note <= (-12187);
                5312: note <= (-14886);
                5313: note <= (-15491);
                5314: note <= (-13722);
                5315: note <= (-9889);
                5316: note <= (-4815);
                5317: note <= 377;
                5318: note <= 4563;
                5319: note <= 6910;
                5320: note <= 7094;
                5321: note <= 5378;
                5322: note <= 2531;
                5323: note <= (-377);
                5324: note <= (-2279);
                5325: note <= (-2399);
                5326: note <= (-467);
                5327: note <= 3203;
                5328: note <= 7791;
                5329: note <= 12187;
                5330: note <= 15286;
                5331: note <= 16283;
                5332: note <= 14886;
                5333: note <= 11395;
                5334: note <= 6627;
                5335: note <= 1697;
                5336: note <= (-2279);
                5337: note <= (-4473);
                5338: note <= (-4563);
                5339: note <= (-2814);
                5340: note <= 0;
                5341: note <= 2814;
                5342: note <= 4563;
                5343: note <= 4473;
                5344: note <= 2279;
                5345: note <= (-1697);
                5346: note <= (-6627);
                5347: note <= (-11395);
                5348: note <= (-14886);
                5349: note <= (-16283);
                5350: note <= (-15286);
                5351: note <= (-12187);
                5352: note <= (-7791);
                5353: note <= (-3203);
                5354: note <= 467;
                5355: note <= 2399;
                5356: note <= 2279;
                5357: note <= 377;
                5358: note <= (-2531);
                5359: note <= (-5378);
                5360: note <= (-7094);
                5361: note <= (-6910);
                5362: note <= (-4563);
                5363: note <= (-377);
                5364: note <= 4815;
                5365: note <= 9889;
                5366: note <= 13722;
                5367: note <= 15491;
                5368: note <= 14886;
                5369: note <= 12187;
                5370: note <= 8192;
                5371: note <= 3995;
                5372: note <= 697;
                5373: note <= (-893);
                5374: note <= (-467);
                5375: note <= 1697;
                5376: note <= 4815;
                5377: note <= 7815;
                5378: note <= 9626;
                5379: note <= 9474;
                5380: note <= 7094;
                5381: note <= 2814;
                5382: note <= (-2531);
                5383: note <= (-7815);
                5384: note <= (-11910);
                5385: note <= (-13985);
                5386: note <= (-13722);
                5387: note <= (-11395);
                5388: note <= (-7791);
                5389: note <= (-3995);
                5390: note <= (-1098);
                5391: note <= 101;
                5392: note <= (-697);
                5393: note <= (-3203);
                5394: note <= (-6627);
                5395: note <= (-9889);
                5396: note <= (-11910);
                5397: note <= (-11911);
                5398: note <= (-9626);
                5399: note <= (-5378);
                5400: note <= 0;
                5401: note <= 5378;
                5402: note <= 9626;
                5403: note <= 11911;
                5404: note <= 11910;
                5405: note <= 9889;
                5406: note <= 6627;
                5407: note <= 3203;
                5408: note <= 697;
                5409: note <= (-101);
                5410: note <= 1098;
                5411: note <= 3995;
                5412: note <= 7791;
                5413: note <= 11395;
                5414: note <= 13722;
                5415: note <= 13985;
                5416: note <= 11910;
                5417: note <= 7815;
                5418: note <= 2531;
                5419: note <= (-2814);
                5420: note <= (-7094);
                5421: note <= (-9474);
                5422: note <= (-9626);
                5423: note <= (-7815);
                5424: note <= (-4815);
                5425: note <= (-1697);
                5426: note <= 467;
                5427: note <= 893;
                5428: note <= (-697);
                5429: note <= (-3995);
                5430: note <= (-8192);
                5431: note <= (-12187);
                5432: note <= (-14886);
                5433: note <= (-15491);
                5434: note <= (-13722);
                5435: note <= (-9889);
                5436: note <= (-4815);
                5437: note <= 377;
                5438: note <= 4563;
                5439: note <= 6910;
                5440: note <= 7094;
                5441: note <= 5378;
                5442: note <= 2531;
                5443: note <= (-377);
                5444: note <= (-2279);
                5445: note <= (-2399);
                5446: note <= (-467);
                5447: note <= 3203;
                5448: note <= 7791;
                5449: note <= 12187;
                5450: note <= 15286;
                5451: note <= 16283;
                5452: note <= 14886;
                5453: note <= 11395;
                5454: note <= 6627;
                5455: note <= 1697;
                5456: note <= (-2279);
                5457: note <= (-4473);
                5458: note <= (-4563);
                5459: note <= (-2814);
                5460: note <= 0;
                5461: note <= 2814;
                5462: note <= 4563;
                5463: note <= 4473;
                5464: note <= 2279;
                5465: note <= (-1697);
                5466: note <= (-6627);
                5467: note <= (-11395);
                5468: note <= (-14886);
                5469: note <= (-16283);
                5470: note <= (-15286);
                5471: note <= (-12187);
                5472: note <= (-7791);
                5473: note <= (-3203);
                5474: note <= 467;
                5475: note <= 2399;
                5476: note <= 2279;
                5477: note <= 377;
                5478: note <= (-2531);
                5479: note <= (-5378);
                5480: note <= (-7094);
                5481: note <= (-6910);
                5482: note <= (-4563);
                5483: note <= (-377);
                5484: note <= 4815;
                5485: note <= 9889;
                5486: note <= 13722;
                5487: note <= 15491;
                5488: note <= 14886;
                5489: note <= 12187;
                5490: note <= 8192;
                5491: note <= 3995;
                5492: note <= 697;
                5493: note <= (-893);
                5494: note <= (-467);
                5495: note <= 1697;
                5496: note <= 4815;
                5497: note <= 7815;
                5498: note <= 9626;
                5499: note <= 9474;
                5500: note <= 7094;
                5501: note <= 2814;
                5502: note <= (-2531);
                5503: note <= (-7815);
                5504: note <= (-11910);
                5505: note <= (-13985);
                5506: note <= (-13722);
                5507: note <= (-11395);
                5508: note <= (-7791);
                5509: note <= (-3995);
                5510: note <= (-1098);
                5511: note <= 101;
                5512: note <= (-697);
                5513: note <= (-3203);
                5514: note <= (-6627);
                5515: note <= (-9889);
                5516: note <= (-11910);
                5517: note <= (-11911);
                5518: note <= (-9626);
                5519: note <= (-5378);
                5520: note <= 0;
                5521: note <= 5378;
                5522: note <= 9626;
                5523: note <= 11911;
                5524: note <= 11910;
                5525: note <= 9889;
                5526: note <= 6627;
                5527: note <= 3203;
                5528: note <= 697;
                5529: note <= (-101);
                5530: note <= 1098;
                5531: note <= 3995;
                5532: note <= 7791;
                5533: note <= 11395;
                5534: note <= 13722;
                5535: note <= 13985;
                5536: note <= 11910;
                5537: note <= 7815;
                5538: note <= 2531;
                5539: note <= (-2814);
                5540: note <= (-7094);
                5541: note <= (-9474);
                5542: note <= (-9626);
                5543: note <= (-7815);
                5544: note <= (-4815);
                5545: note <= (-1697);
                5546: note <= 467;
                5547: note <= 893;
                5548: note <= (-697);
                5549: note <= (-3995);
                5550: note <= (-8192);
                5551: note <= (-12187);
                5552: note <= (-14886);
                5553: note <= (-15491);
                5554: note <= (-13722);
                5555: note <= (-9889);
                5556: note <= (-4815);
                5557: note <= 377;
                5558: note <= 4563;
                5559: note <= 6910;
                5560: note <= 7094;
                5561: note <= 5378;
                5562: note <= 2531;
                5563: note <= (-377);
                5564: note <= (-2279);
                5565: note <= (-2399);
                5566: note <= (-467);
                5567: note <= 3203;
                5568: note <= 7791;
                5569: note <= 12187;
                5570: note <= 15286;
                5571: note <= 16283;
                5572: note <= 14886;
                5573: note <= 11395;
                5574: note <= 6627;
                5575: note <= 1697;
                5576: note <= (-2279);
                5577: note <= (-4473);
                5578: note <= (-4563);
                5579: note <= (-2814);
                5580: note <= 0;
                5581: note <= 2814;
                5582: note <= 4563;
                5583: note <= 4473;
                5584: note <= 2279;
                5585: note <= (-1697);
                5586: note <= (-6627);
                5587: note <= (-11395);
                5588: note <= (-14886);
                5589: note <= (-16283);
                5590: note <= (-15286);
                5591: note <= (-12187);
                5592: note <= (-7791);
                5593: note <= (-3203);
                5594: note <= 467;
                5595: note <= 2399;
                5596: note <= 2279;
                5597: note <= 377;
                5598: note <= (-2531);
                5599: note <= (-5378);
                5600: note <= (-7094);
                5601: note <= (-6910);
                5602: note <= (-4563);
                5603: note <= (-377);
                5604: note <= 4815;
                5605: note <= 9889;
                5606: note <= 13722;
                5607: note <= 15491;
                5608: note <= 14886;
                5609: note <= 12187;
                5610: note <= 8192;
                5611: note <= 3995;
                5612: note <= 697;
                5613: note <= (-893);
                5614: note <= (-467);
                5615: note <= 1697;
                5616: note <= 4815;
                5617: note <= 7815;
                5618: note <= 9626;
                5619: note <= 9474;
                5620: note <= 7094;
                5621: note <= 2814;
                5622: note <= (-2531);
                5623: note <= (-7815);
                5624: note <= (-11910);
                5625: note <= (-13985);
                5626: note <= (-13722);
                5627: note <= (-11395);
                5628: note <= (-7791);
                5629: note <= (-3995);
                5630: note <= (-1098);
                5631: note <= 101;
                5632: note <= (-697);
                5633: note <= (-3203);
                5634: note <= (-6627);
                5635: note <= (-9889);
                5636: note <= (-11910);
                5637: note <= (-11911);
                5638: note <= (-9626);
                5639: note <= (-5378);
                5640: note <= 0;
                5641: note <= 5378;
                5642: note <= 9626;
                5643: note <= 11911;
                5644: note <= 11910;
                5645: note <= 9889;
                5646: note <= 6627;
                5647: note <= 3203;
                5648: note <= 697;
                5649: note <= (-101);
                5650: note <= 1098;
                5651: note <= 3995;
                5652: note <= 7791;
                5653: note <= 11395;
                5654: note <= 13722;
                5655: note <= 13985;
                5656: note <= 11910;
                5657: note <= 7815;
                5658: note <= 2531;
                5659: note <= (-2814);
                5660: note <= (-7094);
                5661: note <= (-9474);
                5662: note <= (-9626);
                5663: note <= (-7815);
                5664: note <= (-4815);
                5665: note <= (-1697);
                5666: note <= 467;
                5667: note <= 893;
                5668: note <= (-697);
                5669: note <= (-3995);
                5670: note <= (-8192);
                5671: note <= (-12187);
                5672: note <= (-14886);
                5673: note <= (-15491);
                5674: note <= (-13722);
                5675: note <= (-9889);
                5676: note <= (-4815);
                5677: note <= 377;
                5678: note <= 4563;
                5679: note <= 6910;
                5680: note <= 7094;
                5681: note <= 5378;
                5682: note <= 2531;
                5683: note <= (-377);
                5684: note <= (-2279);
                5685: note <= (-2399);
                5686: note <= (-467);
                5687: note <= 3203;
                5688: note <= 7791;
                5689: note <= 12187;
                5690: note <= 15286;
                5691: note <= 16283;
                5692: note <= 14886;
                5693: note <= 11395;
                5694: note <= 6627;
                5695: note <= 1697;
                5696: note <= (-2279);
                5697: note <= (-4473);
                5698: note <= (-4563);
                5699: note <= (-2814);
                5700: note <= 0;
                5701: note <= 2814;
                5702: note <= 4563;
                5703: note <= 4473;
                5704: note <= 2279;
                5705: note <= (-1697);
                5706: note <= (-6627);
                5707: note <= (-11395);
                5708: note <= (-14886);
                5709: note <= (-16283);
                5710: note <= (-15286);
                5711: note <= (-12187);
                5712: note <= (-7791);
                5713: note <= (-3203);
                5714: note <= 467;
                5715: note <= 2399;
                5716: note <= 2279;
                5717: note <= 377;
                5718: note <= (-2531);
                5719: note <= (-5378);
                5720: note <= (-7094);
                5721: note <= (-6910);
                5722: note <= (-4563);
                5723: note <= (-377);
                5724: note <= 4815;
                5725: note <= 9889;
                5726: note <= 13722;
                5727: note <= 15491;
                5728: note <= 14886;
                5729: note <= 12187;
                5730: note <= 8192;
                5731: note <= 3995;
                5732: note <= 697;
                5733: note <= (-893);
                5734: note <= (-467);
                5735: note <= 1697;
                5736: note <= 4815;
                5737: note <= 7815;
                5738: note <= 9626;
                5739: note <= 9474;
                5740: note <= 7094;
                5741: note <= 2814;
                5742: note <= (-2531);
                5743: note <= (-7815);
                5744: note <= (-11910);
                5745: note <= (-13985);
                5746: note <= (-13722);
                5747: note <= (-11395);
                5748: note <= (-7791);
                5749: note <= (-3995);
                5750: note <= (-1098);
                5751: note <= 101;
                5752: note <= (-697);
                5753: note <= (-3203);
                5754: note <= (-6627);
                5755: note <= (-9889);
                5756: note <= (-11910);
                5757: note <= (-11911);
                5758: note <= (-9626);
                5759: note <= (-5378);
                5760: note <= 0;
                5761: note <= 5378;
                5762: note <= 9626;
                5763: note <= 11911;
                5764: note <= 11910;
                5765: note <= 9889;
                5766: note <= 6627;
                5767: note <= 3203;
                5768: note <= 697;
                5769: note <= (-101);
                5770: note <= 1098;
                5771: note <= 3995;
                5772: note <= 7791;
                5773: note <= 11395;
                5774: note <= 13722;
                5775: note <= 13985;
                5776: note <= 11910;
                5777: note <= 7815;
                5778: note <= 2531;
                5779: note <= (-2814);
                5780: note <= (-7094);
                5781: note <= (-9474);
                5782: note <= (-9626);
                5783: note <= (-7815);
                5784: note <= (-4815);
                5785: note <= (-1697);
                5786: note <= 467;
                5787: note <= 893;
                5788: note <= (-697);
                5789: note <= (-3995);
                5790: note <= (-8192);
                5791: note <= (-12187);
                5792: note <= (-14886);
                5793: note <= (-15491);
                5794: note <= (-13722);
                5795: note <= (-9889);
                5796: note <= (-4815);
                5797: note <= 377;
                5798: note <= 4563;
                5799: note <= 6910;
                5800: note <= 7094;
                5801: note <= 5378;
                5802: note <= 2531;
                5803: note <= (-377);
                5804: note <= (-2279);
                5805: note <= (-2399);
                5806: note <= (-467);
                5807: note <= 3203;
                5808: note <= 7791;
                5809: note <= 12187;
                5810: note <= 15286;
                5811: note <= 16283;
                5812: note <= 14886;
                5813: note <= 11395;
                5814: note <= 6627;
                5815: note <= 1697;
                5816: note <= (-2279);
                5817: note <= (-4473);
                5818: note <= (-4563);
                5819: note <= (-2814);
                5820: note <= 0;
                5821: note <= 2814;
                5822: note <= 4563;
                5823: note <= 4473;
                5824: note <= 2279;
                5825: note <= (-1697);
                5826: note <= (-6627);
                5827: note <= (-11395);
                5828: note <= (-14886);
                5829: note <= (-16283);
                5830: note <= (-15286);
                5831: note <= (-12187);
                5832: note <= (-7791);
                5833: note <= (-3203);
                5834: note <= 467;
                5835: note <= 2399;
                5836: note <= 2279;
                5837: note <= 377;
                5838: note <= (-2531);
                5839: note <= (-5378);
                5840: note <= (-7094);
                5841: note <= (-6910);
                5842: note <= (-4563);
                5843: note <= (-377);
                5844: note <= 4815;
                5845: note <= 9889;
                5846: note <= 13722;
                5847: note <= 15491;
                5848: note <= 14886;
                5849: note <= 12187;
                5850: note <= 8192;
                5851: note <= 3995;
                5852: note <= 697;
                5853: note <= (-893);
                5854: note <= (-467);
                5855: note <= 1697;
                5856: note <= 4815;
                5857: note <= 7815;
                5858: note <= 9626;
                5859: note <= 9474;
                5860: note <= 7094;
                5861: note <= 2814;
                5862: note <= (-2531);
                5863: note <= (-7815);
                5864: note <= (-11910);
                5865: note <= (-13985);
                5866: note <= (-13722);
                5867: note <= (-11395);
                5868: note <= (-7791);
                5869: note <= (-3995);
                5870: note <= (-1098);
                5871: note <= 101;
                5872: note <= (-697);
                5873: note <= (-3203);
                5874: note <= (-6627);
                5875: note <= (-9889);
                5876: note <= (-11910);
                5877: note <= (-11911);
                5878: note <= (-9626);
                5879: note <= (-5378);
                5880: note <= 0;
                5881: note <= 5378;
                5882: note <= 9626;
                5883: note <= 11911;
                5884: note <= 11910;
                5885: note <= 9889;
                5886: note <= 6627;
                5887: note <= 3203;
                5888: note <= 697;
                5889: note <= (-101);
                5890: note <= 1098;
                5891: note <= 3995;
                5892: note <= 7791;
                5893: note <= 11395;
                5894: note <= 13722;
                5895: note <= 13985;
                5896: note <= 11910;
                5897: note <= 7815;
                5898: note <= 2531;
                5899: note <= (-2814);
                5900: note <= (-7094);
                5901: note <= (-9474);
                5902: note <= (-9626);
                5903: note <= (-7815);
                5904: note <= (-4815);
                5905: note <= (-1697);
                5906: note <= 467;
                5907: note <= 893;
                5908: note <= (-697);
                5909: note <= (-3995);
                5910: note <= (-8192);
                5911: note <= (-12187);
                5912: note <= (-14886);
                5913: note <= (-15491);
                5914: note <= (-13722);
                5915: note <= (-9889);
                5916: note <= (-4815);
                5917: note <= 377;
                5918: note <= 4563;
                5919: note <= 6910;
                5920: note <= 7094;
                5921: note <= 5378;
                5922: note <= 2531;
                5923: note <= (-377);
                5924: note <= (-2279);
                5925: note <= (-2399);
                5926: note <= (-467);
                5927: note <= 3203;
                5928: note <= 7791;
                5929: note <= 12187;
                5930: note <= 15286;
                5931: note <= 16283;
                5932: note <= 14886;
                5933: note <= 11395;
                5934: note <= 6627;
                5935: note <= 1697;
                5936: note <= (-2279);
                5937: note <= (-4473);
                5938: note <= (-4563);
                5939: note <= (-2814);
                5940: note <= 0;
                5941: note <= 2814;
                5942: note <= 4563;
                5943: note <= 4473;
                5944: note <= 2279;
                5945: note <= (-1697);
                5946: note <= (-6627);
                5947: note <= (-11395);
                5948: note <= (-14886);
                5949: note <= (-16283);
                5950: note <= (-15286);
                5951: note <= (-12187);
                5952: note <= (-7791);
                5953: note <= (-3203);
                5954: note <= 467;
                5955: note <= 2399;
                5956: note <= 2279;
                5957: note <= 377;
                5958: note <= (-2531);
                5959: note <= (-5378);
                5960: note <= (-7094);
                5961: note <= (-6910);
                5962: note <= (-4563);
                5963: note <= (-377);
                5964: note <= 4815;
                5965: note <= 9889;
                5966: note <= 13722;
                5967: note <= 15491;
                5968: note <= 14886;
                5969: note <= 12187;
                5970: note <= 8192;
                5971: note <= 3995;
                5972: note <= 697;
                5973: note <= (-893);
                5974: note <= (-467);
                5975: note <= 1697;
                5976: note <= 4815;
                5977: note <= 7815;
                5978: note <= 9626;
                5979: note <= 9474;
                5980: note <= 7094;
                5981: note <= 2814;
                5982: note <= (-2531);
                5983: note <= (-7815);
                5984: note <= (-11910);
                5985: note <= (-13985);
                5986: note <= (-13722);
                5987: note <= (-11395);
                5988: note <= (-7791);
                5989: note <= (-3995);
                5990: note <= (-1098);
                5991: note <= 101;
                5992: note <= (-697);
                5993: note <= (-3203);
                5994: note <= (-6627);
                5995: note <= (-9889);
                5996: note <= (-11910);
                5997: note <= (-11911);
                5998: note <= (-9626);
                5999: note <= (-5378);
                6000: note <= 0;
                6001: note <= 5378;
                6002: note <= 9626;
                6003: note <= 11911;
                6004: note <= 11910;
                6005: note <= 9889;
                6006: note <= 6627;
                6007: note <= 3203;
                6008: note <= 697;
                6009: note <= (-101);
                6010: note <= 1098;
                6011: note <= 3995;
                6012: note <= 7791;
                6013: note <= 11395;
                6014: note <= 13722;
                6015: note <= 13985;
                6016: note <= 11910;
                6017: note <= 7815;
                6018: note <= 2531;
                6019: note <= (-2814);
                6020: note <= (-7094);
                6021: note <= (-9474);
                6022: note <= (-9626);
                6023: note <= (-7815);
                6024: note <= (-4815);
                6025: note <= (-1697);
                6026: note <= 467;
                6027: note <= 893;
                6028: note <= (-697);
                6029: note <= (-3995);
                6030: note <= (-8192);
                6031: note <= (-12187);
                6032: note <= (-14886);
                6033: note <= (-15491);
                6034: note <= (-13722);
                6035: note <= (-9889);
                6036: note <= (-4815);
                6037: note <= 377;
                6038: note <= 4563;
                6039: note <= 6910;
                6040: note <= 7094;
                6041: note <= 5378;
                6042: note <= 2531;
                6043: note <= (-377);
                6044: note <= (-2279);
                6045: note <= (-2399);
                6046: note <= (-467);
                6047: note <= 3203;
                6048: note <= 7791;
                6049: note <= 12187;
                6050: note <= 15286;
                6051: note <= 16283;
                6052: note <= 14886;
                6053: note <= 11395;
                6054: note <= 6627;
                6055: note <= 1697;
                6056: note <= (-2279);
                6057: note <= (-4473);
                6058: note <= (-4563);
                6059: note <= (-2814);
                6060: note <= 0;
                6061: note <= 2814;
                6062: note <= 4563;
                6063: note <= 4473;
                6064: note <= 2279;
                6065: note <= (-1697);
                6066: note <= (-6627);
                6067: note <= (-11395);
                6068: note <= (-14886);
                6069: note <= (-16283);
                6070: note <= (-15286);
                6071: note <= (-12187);
                6072: note <= (-7791);
                6073: note <= (-3203);
                6074: note <= 467;
                6075: note <= 2399;
                6076: note <= 2279;
                6077: note <= 377;
                6078: note <= (-2531);
                6079: note <= (-5378);
                6080: note <= (-7094);
                6081: note <= (-6910);
                6082: note <= (-4563);
                6083: note <= (-377);
                6084: note <= 4815;
                6085: note <= 9889;
                6086: note <= 13722;
                6087: note <= 15491;
                6088: note <= 14886;
                6089: note <= 12187;
                6090: note <= 8192;
                6091: note <= 3995;
                6092: note <= 697;
                6093: note <= (-893);
                6094: note <= (-467);
                6095: note <= 1697;
                6096: note <= 4815;
                6097: note <= 7815;
                6098: note <= 9626;
                6099: note <= 9474;
                6100: note <= 7094;
                6101: note <= 2814;
                6102: note <= (-2531);
                6103: note <= (-7815);
                6104: note <= (-11910);
                6105: note <= (-13985);
                6106: note <= (-13722);
                6107: note <= (-11395);
                6108: note <= (-7791);
                6109: note <= (-3995);
                6110: note <= (-1098);
                6111: note <= 101;
                6112: note <= (-697);
                6113: note <= (-3203);
                6114: note <= (-6627);
                6115: note <= (-9889);
                6116: note <= (-11910);
                6117: note <= (-11911);
                6118: note <= (-9626);
                6119: note <= (-5378);
                6120: note <= 0;
                6121: note <= 5378;
                6122: note <= 9626;
                6123: note <= 11911;
                6124: note <= 11910;
                6125: note <= 9889;
                6126: note <= 6627;
                6127: note <= 3203;
                6128: note <= 697;
                6129: note <= (-101);
                6130: note <= 1098;
                6131: note <= 3995;
                6132: note <= 7791;
                6133: note <= 11395;
                6134: note <= 13722;
                6135: note <= 13985;
                6136: note <= 11910;
                6137: note <= 7815;
                6138: note <= 2531;
                6139: note <= (-2814);
                6140: note <= (-7094);
                6141: note <= (-9474);
                6142: note <= (-9626);
                6143: note <= (-7815);
                6144: note <= (-4815);
                6145: note <= (-1697);
                6146: note <= 467;
                6147: note <= 893;
                6148: note <= (-697);
                6149: note <= (-3995);
                6150: note <= (-8192);
                6151: note <= (-12187);
                6152: note <= (-14886);
                6153: note <= (-15491);
                6154: note <= (-13722);
                6155: note <= (-9889);
                6156: note <= (-4815);
                6157: note <= 377;
                6158: note <= 4563;
                6159: note <= 6910;
                6160: note <= 7094;
                6161: note <= 5378;
                6162: note <= 2531;
                6163: note <= (-377);
                6164: note <= (-2279);
                6165: note <= (-2399);
                6166: note <= (-467);
                6167: note <= 3203;
                6168: note <= 7791;
                6169: note <= 12187;
                6170: note <= 15286;
                6171: note <= 16283;
                6172: note <= 14886;
                6173: note <= 11395;
                6174: note <= 6627;
                6175: note <= 1697;
                6176: note <= (-2279);
                6177: note <= (-4473);
                6178: note <= (-4563);
                6179: note <= (-2814);
                6180: note <= 0;
                6181: note <= 2814;
                6182: note <= 4563;
                6183: note <= 4473;
                6184: note <= 2279;
                6185: note <= (-1697);
                6186: note <= (-6627);
                6187: note <= (-11395);
                6188: note <= (-14886);
                6189: note <= (-16283);
                6190: note <= (-15286);
                6191: note <= (-12187);
                6192: note <= (-7791);
                6193: note <= (-3203);
                6194: note <= 467;
                6195: note <= 2399;
                6196: note <= 2279;
                6197: note <= 377;
                6198: note <= (-2531);
                6199: note <= (-5378);
                6200: note <= (-7094);
                6201: note <= (-6910);
                6202: note <= (-4563);
                6203: note <= (-377);
                6204: note <= 4815;
                6205: note <= 9889;
                6206: note <= 13722;
                6207: note <= 15491;
                6208: note <= 14886;
                6209: note <= 12187;
                6210: note <= 8192;
                6211: note <= 3995;
                6212: note <= 697;
                6213: note <= (-893);
                6214: note <= (-467);
                6215: note <= 1697;
                6216: note <= 4815;
                6217: note <= 7815;
                6218: note <= 9626;
                6219: note <= 9474;
                6220: note <= 7094;
                6221: note <= 2814;
                6222: note <= (-2531);
                6223: note <= (-7815);
                6224: note <= (-11910);
                6225: note <= (-13985);
                6226: note <= (-13722);
                6227: note <= (-11395);
                6228: note <= (-7791);
                6229: note <= (-3995);
                6230: note <= (-1098);
                6231: note <= 101;
                6232: note <= (-697);
                6233: note <= (-3203);
                6234: note <= (-6627);
                6235: note <= (-9889);
                6236: note <= (-11910);
                6237: note <= (-11911);
                6238: note <= (-9626);
                6239: note <= (-5378);
                6240: note <= 0;
                6241: note <= 5378;
                6242: note <= 9626;
                6243: note <= 11911;
                6244: note <= 11910;
                6245: note <= 9889;
                6246: note <= 6627;
                6247: note <= 3203;
                6248: note <= 697;
                6249: note <= (-101);
                6250: note <= 1098;
                6251: note <= 3995;
                6252: note <= 7791;
                6253: note <= 11395;
                6254: note <= 13722;
                6255: note <= 13985;
                6256: note <= 11910;
                6257: note <= 7815;
                6258: note <= 2531;
                6259: note <= (-2814);
                6260: note <= (-7094);
                6261: note <= (-9474);
                6262: note <= (-9626);
                6263: note <= (-7815);
                6264: note <= (-4815);
                6265: note <= (-1697);
                6266: note <= 467;
                6267: note <= 893;
                6268: note <= (-697);
                6269: note <= (-3995);
                6270: note <= (-8192);
                6271: note <= (-12187);
                6272: note <= (-14886);
                6273: note <= (-15491);
                6274: note <= (-13722);
                6275: note <= (-9889);
                6276: note <= (-4815);
                6277: note <= 377;
                6278: note <= 4563;
                6279: note <= 6910;
                6280: note <= 7094;
                6281: note <= 5378;
                6282: note <= 2531;
                6283: note <= (-377);
                6284: note <= (-2279);
                6285: note <= (-2399);
                6286: note <= (-467);
                6287: note <= 3203;
                6288: note <= 7791;
                6289: note <= 12187;
                6290: note <= 15286;
                6291: note <= 16283;
                6292: note <= 14886;
                6293: note <= 11395;
                6294: note <= 6627;
                6295: note <= 1697;
                6296: note <= (-2279);
                6297: note <= (-4473);
                6298: note <= (-4563);
                6299: note <= (-2814);
                6300: note <= 0;
                6301: note <= 2814;
                6302: note <= 4563;
                6303: note <= 4473;
                6304: note <= 2279;
                6305: note <= (-1697);
                6306: note <= (-6627);
                6307: note <= (-11395);
                6308: note <= (-14886);
                6309: note <= (-16283);
                6310: note <= (-15286);
                6311: note <= (-12187);
                6312: note <= (-7791);
                6313: note <= (-3203);
                6314: note <= 467;
                6315: note <= 2399;
                6316: note <= 2279;
                6317: note <= 377;
                6318: note <= (-2531);
                6319: note <= (-5378);
                6320: note <= (-7094);
                6321: note <= (-6910);
                6322: note <= (-4563);
                6323: note <= (-377);
                6324: note <= 4815;
                6325: note <= 9889;
                6326: note <= 13722;
                6327: note <= 15491;
                6328: note <= 14886;
                6329: note <= 12187;
                6330: note <= 8192;
                6331: note <= 3995;
                6332: note <= 697;
                6333: note <= (-893);
                6334: note <= (-467);
                6335: note <= 1697;
                6336: note <= 4815;
                6337: note <= 7815;
                6338: note <= 9626;
                6339: note <= 9474;
                6340: note <= 7094;
                6341: note <= 2814;
                6342: note <= (-2531);
                6343: note <= (-7815);
                6344: note <= (-11910);
                6345: note <= (-13985);
                6346: note <= (-13722);
                6347: note <= (-11395);
                6348: note <= (-7791);
                6349: note <= (-3995);
                6350: note <= (-1098);
                6351: note <= 101;
                6352: note <= (-697);
                6353: note <= (-3203);
                6354: note <= (-6627);
                6355: note <= (-9889);
                6356: note <= (-11910);
                6357: note <= (-11911);
                6358: note <= (-9626);
                6359: note <= (-5378);
                6360: note <= 0;
                6361: note <= 5378;
                6362: note <= 9626;
                6363: note <= 11911;
                6364: note <= 11910;
                6365: note <= 9889;
                6366: note <= 6627;
                6367: note <= 3203;
                6368: note <= 697;
                6369: note <= (-101);
                6370: note <= 1098;
                6371: note <= 3995;
                6372: note <= 7791;
                6373: note <= 11395;
                6374: note <= 13722;
                6375: note <= 13985;
                6376: note <= 11910;
                6377: note <= 7815;
                6378: note <= 2531;
                6379: note <= (-2814);
                6380: note <= (-7094);
                6381: note <= (-9474);
                6382: note <= (-9626);
                6383: note <= (-7815);
                6384: note <= (-4815);
                6385: note <= (-1697);
                6386: note <= 467;
                6387: note <= 893;
                6388: note <= (-697);
                6389: note <= (-3995);
                6390: note <= (-8192);
                6391: note <= (-12187);
                6392: note <= (-14886);
                6393: note <= (-15491);
                6394: note <= (-13722);
                6395: note <= (-9889);
                6396: note <= (-4815);
                6397: note <= 377;
                6398: note <= 4563;
                6399: note <= 6910;
                6400: note <= 7094;
                6401: note <= 5378;
                6402: note <= 2531;
                6403: note <= (-377);
                6404: note <= (-2279);
                6405: note <= (-2399);
                6406: note <= (-467);
                6407: note <= 3203;
                6408: note <= 7791;
                6409: note <= 12187;
                6410: note <= 15286;
                6411: note <= 16283;
                6412: note <= 14886;
                6413: note <= 11395;
                6414: note <= 6627;
                6415: note <= 1697;
                6416: note <= (-2279);
                6417: note <= (-4473);
                6418: note <= (-4563);
                6419: note <= (-2814);
                6420: note <= 0;
                6421: note <= 2814;
                6422: note <= 4563;
                6423: note <= 4473;
                6424: note <= 2279;
                6425: note <= (-1697);
                6426: note <= (-6627);
                6427: note <= (-11395);
                6428: note <= (-14886);
                6429: note <= (-16283);
                6430: note <= (-15286);
                6431: note <= (-12187);
                6432: note <= (-7791);
                6433: note <= (-3203);
                6434: note <= 467;
                6435: note <= 2399;
                6436: note <= 2279;
                6437: note <= 377;
                6438: note <= (-2531);
                6439: note <= (-5378);
                6440: note <= (-7094);
                6441: note <= (-6910);
                6442: note <= (-4563);
                6443: note <= (-377);
                6444: note <= 4815;
                6445: note <= 9889;
                6446: note <= 13722;
                6447: note <= 15491;
                6448: note <= 14886;
                6449: note <= 12187;
                6450: note <= 8192;
                6451: note <= 3995;
                6452: note <= 697;
                6453: note <= (-893);
                6454: note <= (-467);
                6455: note <= 1697;
                6456: note <= 4815;
                6457: note <= 7815;
                6458: note <= 9626;
                6459: note <= 9474;
                6460: note <= 7094;
                6461: note <= 2814;
                6462: note <= (-2531);
                6463: note <= (-7815);
                6464: note <= (-11910);
                6465: note <= (-13985);
                6466: note <= (-13722);
                6467: note <= (-11395);
                6468: note <= (-7791);
                6469: note <= (-3995);
                6470: note <= (-1098);
                6471: note <= 101;
                6472: note <= (-697);
                6473: note <= (-3203);
                6474: note <= (-6627);
                6475: note <= (-9889);
                6476: note <= (-11910);
                6477: note <= (-11911);
                6478: note <= (-9626);
                6479: note <= (-5378);
                6480: note <= 0;
                6481: note <= 5378;
                6482: note <= 9626;
                6483: note <= 11911;
                6484: note <= 11910;
                6485: note <= 9889;
                6486: note <= 6627;
                6487: note <= 3203;
                6488: note <= 697;
                6489: note <= (-101);
                6490: note <= 1098;
                6491: note <= 3995;
                6492: note <= 7791;
                6493: note <= 11395;
                6494: note <= 13722;
                6495: note <= 13985;
                6496: note <= 11910;
                6497: note <= 7815;
                6498: note <= 2531;
                6499: note <= (-2814);
                6500: note <= (-7094);
                6501: note <= (-9474);
                6502: note <= (-9626);
                6503: note <= (-7815);
                6504: note <= (-4815);
                6505: note <= (-1697);
                6506: note <= 467;
                6507: note <= 893;
                6508: note <= (-697);
                6509: note <= (-3995);
                6510: note <= (-8192);
                6511: note <= (-12187);
                6512: note <= (-14886);
                6513: note <= (-15491);
                6514: note <= (-13722);
                6515: note <= (-9889);
                6516: note <= (-4815);
                6517: note <= 377;
                6518: note <= 4563;
                6519: note <= 6910;
                6520: note <= 7094;
                6521: note <= 5378;
                6522: note <= 2531;
                6523: note <= (-377);
                6524: note <= (-2279);
                6525: note <= (-2399);
                6526: note <= (-467);
                6527: note <= 3203;
                6528: note <= 7791;
                6529: note <= 12187;
                6530: note <= 15286;
                6531: note <= 16283;
                6532: note <= 14886;
                6533: note <= 11395;
                6534: note <= 6627;
                6535: note <= 1697;
                6536: note <= (-2279);
                6537: note <= (-4473);
                6538: note <= (-4563);
                6539: note <= (-2814);
                6540: note <= 0;
                6541: note <= 2814;
                6542: note <= 4563;
                6543: note <= 4473;
                6544: note <= 2279;
                6545: note <= (-1697);
                6546: note <= (-6627);
                6547: note <= (-11395);
                6548: note <= (-14886);
                6549: note <= (-16283);
                6550: note <= (-15286);
                6551: note <= (-12187);
                6552: note <= (-7791);
                6553: note <= (-3203);
                6554: note <= 467;
                6555: note <= 2399;
                6556: note <= 2279;
                6557: note <= 377;
                6558: note <= (-2531);
                6559: note <= (-5378);
                6560: note <= (-7094);
                6561: note <= (-6910);
                6562: note <= (-4563);
                6563: note <= (-377);
                6564: note <= 4815;
                6565: note <= 9889;
                6566: note <= 13722;
                6567: note <= 15491;
                6568: note <= 14886;
                6569: note <= 12187;
                6570: note <= 8192;
                6571: note <= 3995;
                6572: note <= 697;
                6573: note <= (-893);
                6574: note <= (-467);
                6575: note <= 1697;
                6576: note <= 4815;
                6577: note <= 7815;
                6578: note <= 9626;
                6579: note <= 9474;
                6580: note <= 7094;
                6581: note <= 2814;
                6582: note <= (-2531);
                6583: note <= (-7815);
                6584: note <= (-11910);
                6585: note <= (-13985);
                6586: note <= (-13722);
                6587: note <= (-11395);
                6588: note <= (-7791);
                6589: note <= (-3995);
                6590: note <= (-1098);
                6591: note <= 101;
                6592: note <= (-697);
                6593: note <= (-3203);
                6594: note <= (-6627);
                6595: note <= (-9889);
                6596: note <= (-11910);
                6597: note <= (-11911);
                6598: note <= (-9626);
                6599: note <= (-5378);
                6600: note <= 0;
                6601: note <= 5378;
                6602: note <= 9626;
                6603: note <= 11911;
                6604: note <= 11910;
                6605: note <= 9889;
                6606: note <= 6627;
                6607: note <= 3203;
                6608: note <= 697;
                6609: note <= (-101);
                6610: note <= 1098;
                6611: note <= 3995;
                6612: note <= 7791;
                6613: note <= 11395;
                6614: note <= 13722;
                6615: note <= 13985;
                6616: note <= 11910;
                6617: note <= 7815;
                6618: note <= 2531;
                6619: note <= (-2814);
                6620: note <= (-7094);
                6621: note <= (-9474);
                6622: note <= (-9626);
                6623: note <= (-7815);
                6624: note <= (-4815);
                6625: note <= (-1697);
                6626: note <= 467;
                6627: note <= 893;
                6628: note <= (-697);
                6629: note <= (-3995);
                6630: note <= (-8192);
                6631: note <= (-12187);
                6632: note <= (-14886);
                6633: note <= (-15491);
                6634: note <= (-13722);
                6635: note <= (-9889);
                6636: note <= (-4815);
                6637: note <= 377;
                6638: note <= 4563;
                6639: note <= 6910;
                6640: note <= 7094;
                6641: note <= 5378;
                6642: note <= 2531;
                6643: note <= (-377);
                6644: note <= (-2279);
                6645: note <= (-2399);
                6646: note <= (-467);
                6647: note <= 3203;
                6648: note <= 7791;
                6649: note <= 12187;
                6650: note <= 15286;
                6651: note <= 16283;
                6652: note <= 14886;
                6653: note <= 11395;
                6654: note <= 6627;
                6655: note <= 1697;
                6656: note <= (-2279);
                6657: note <= (-4473);
                6658: note <= (-4563);
                6659: note <= (-2814);
                6660: note <= 0;
                6661: note <= 2814;
                6662: note <= 4563;
                6663: note <= 4473;
                6664: note <= 2279;
                6665: note <= (-1697);
                6666: note <= (-6627);
                6667: note <= (-11395);
                6668: note <= (-14886);
                6669: note <= (-16283);
                6670: note <= (-15286);
                6671: note <= (-12187);
                6672: note <= (-7791);
                6673: note <= (-3203);
                6674: note <= 467;
                6675: note <= 2399;
                6676: note <= 2279;
                6677: note <= 377;
                6678: note <= (-2531);
                6679: note <= (-5378);
                6680: note <= (-7094);
                6681: note <= (-6910);
                6682: note <= (-4563);
                6683: note <= (-377);
                6684: note <= 4815;
                6685: note <= 9889;
                6686: note <= 13722;
                6687: note <= 15491;
                6688: note <= 14886;
                6689: note <= 12187;
                6690: note <= 8192;
                6691: note <= 3995;
                6692: note <= 697;
                6693: note <= (-893);
                6694: note <= (-467);
                6695: note <= 1697;
                6696: note <= 4815;
                6697: note <= 7815;
                6698: note <= 9626;
                6699: note <= 9474;
                6700: note <= 7094;
                6701: note <= 2814;
                6702: note <= (-2531);
                6703: note <= (-7815);
                6704: note <= (-11910);
                6705: note <= (-13985);
                6706: note <= (-13722);
                6707: note <= (-11395);
                6708: note <= (-7791);
                6709: note <= (-3995);
                6710: note <= (-1098);
                6711: note <= 101;
                6712: note <= (-697);
                6713: note <= (-3203);
                6714: note <= (-6627);
                6715: note <= (-9889);
                6716: note <= (-11910);
                6717: note <= (-11911);
                6718: note <= (-9626);
                6719: note <= (-5378);
                6720: note <= 0;
                6721: note <= 5378;
                6722: note <= 9626;
                6723: note <= 11911;
                6724: note <= 11910;
                6725: note <= 9889;
                6726: note <= 6627;
                6727: note <= 3203;
                6728: note <= 697;
                6729: note <= (-101);
                6730: note <= 1098;
                6731: note <= 3995;
                6732: note <= 7791;
                6733: note <= 11395;
                6734: note <= 13722;
                6735: note <= 13985;
                6736: note <= 11910;
                6737: note <= 7815;
                6738: note <= 2531;
                6739: note <= (-2814);
                6740: note <= (-7094);
                6741: note <= (-9474);
                6742: note <= (-9626);
                6743: note <= (-7815);
                6744: note <= (-4815);
                6745: note <= (-1697);
                6746: note <= 467;
                6747: note <= 893;
                6748: note <= (-697);
                6749: note <= (-3995);
                6750: note <= (-8192);
                6751: note <= (-12187);
                6752: note <= (-14886);
                6753: note <= (-15491);
                6754: note <= (-13722);
                6755: note <= (-9889);
                6756: note <= (-4815);
                6757: note <= 377;
                6758: note <= 4563;
                6759: note <= 6910;
                6760: note <= 7094;
                6761: note <= 5378;
                6762: note <= 2531;
                6763: note <= (-377);
                6764: note <= (-2279);
                6765: note <= (-2399);
                6766: note <= (-467);
                6767: note <= 3203;
                6768: note <= 7791;
                6769: note <= 12187;
                6770: note <= 15286;
                6771: note <= 16283;
                6772: note <= 14886;
                6773: note <= 11395;
                6774: note <= 6627;
                6775: note <= 1697;
                6776: note <= (-2279);
                6777: note <= (-4473);
                6778: note <= (-4563);
                6779: note <= (-2814);
                6780: note <= 0;
                6781: note <= 2814;
                6782: note <= 4563;
                6783: note <= 4473;
                6784: note <= 2279;
                6785: note <= (-1697);
                6786: note <= (-6627);
                6787: note <= (-11395);
                6788: note <= (-14886);
                6789: note <= (-16283);
                6790: note <= (-15286);
                6791: note <= (-12187);
                6792: note <= (-7791);
                6793: note <= (-3203);
                6794: note <= 467;
                6795: note <= 2399;
                6796: note <= 2279;
                6797: note <= 377;
                6798: note <= (-2531);
                6799: note <= (-5378);
                6800: note <= (-7094);
                6801: note <= (-6910);
                6802: note <= (-4563);
                6803: note <= (-377);
                6804: note <= 4815;
                6805: note <= 9889;
                6806: note <= 13722;
                6807: note <= 15491;
                6808: note <= 14886;
                6809: note <= 12187;
                6810: note <= 8192;
                6811: note <= 3995;
                6812: note <= 697;
                6813: note <= (-893);
                6814: note <= (-467);
                6815: note <= 1697;
                6816: note <= 4815;
                6817: note <= 7815;
                6818: note <= 9626;
                6819: note <= 9474;
                6820: note <= 7094;
                6821: note <= 2814;
                6822: note <= (-2531);
                6823: note <= (-7815);
                6824: note <= (-11910);
                6825: note <= (-13985);
                6826: note <= (-13722);
                6827: note <= (-11395);
                6828: note <= (-7791);
                6829: note <= (-3995);
                6830: note <= (-1098);
                6831: note <= 101;
                6832: note <= (-697);
                6833: note <= (-3203);
                6834: note <= (-6627);
                6835: note <= (-9889);
                6836: note <= (-11910);
                6837: note <= (-11911);
                6838: note <= (-9626);
                6839: note <= (-5378);
                6840: note <= 0;
                6841: note <= 5378;
                6842: note <= 9626;
                6843: note <= 11911;
                6844: note <= 11910;
                6845: note <= 9889;
                6846: note <= 6627;
                6847: note <= 3203;
                6848: note <= 697;
                6849: note <= (-101);
                6850: note <= 1098;
                6851: note <= 3995;
                6852: note <= 7791;
                6853: note <= 11395;
                6854: note <= 13722;
                6855: note <= 13985;
                6856: note <= 11910;
                6857: note <= 7815;
                6858: note <= 2531;
                6859: note <= (-2814);
                6860: note <= (-7094);
                6861: note <= (-9474);
                6862: note <= (-9626);
                6863: note <= (-7815);
                6864: note <= (-4815);
                6865: note <= (-1697);
                6866: note <= 467;
                6867: note <= 893;
                6868: note <= (-697);
                6869: note <= (-3995);
                6870: note <= (-8192);
                6871: note <= (-12187);
                6872: note <= (-14886);
                6873: note <= (-15491);
                6874: note <= (-13722);
                6875: note <= (-9889);
                6876: note <= (-4815);
                6877: note <= 377;
                6878: note <= 4563;
                6879: note <= 6910;
                6880: note <= 7094;
                6881: note <= 5378;
                6882: note <= 2531;
                6883: note <= (-377);
                6884: note <= (-2279);
                6885: note <= (-2399);
                6886: note <= (-467);
                6887: note <= 3203;
                6888: note <= 7791;
                6889: note <= 12187;
                6890: note <= 15286;
                6891: note <= 16283;
                6892: note <= 14886;
                6893: note <= 11395;
                6894: note <= 6627;
                6895: note <= 1697;
                6896: note <= (-2279);
                6897: note <= (-4473);
                6898: note <= (-4563);
                6899: note <= (-2814);
                6900: note <= 0;
                6901: note <= 2814;
                6902: note <= 4563;
                6903: note <= 4473;
                6904: note <= 2279;
                6905: note <= (-1697);
                6906: note <= (-6627);
                6907: note <= (-11395);
                6908: note <= (-14886);
                6909: note <= (-16283);
                6910: note <= (-15286);
                6911: note <= (-12187);
                6912: note <= (-7791);
                6913: note <= (-3203);
                6914: note <= 467;
                6915: note <= 2399;
                6916: note <= 2279;
                6917: note <= 377;
                6918: note <= (-2531);
                6919: note <= (-5378);
                6920: note <= (-7094);
                6921: note <= (-6910);
                6922: note <= (-4563);
                6923: note <= (-377);
                6924: note <= 4815;
                6925: note <= 9889;
                6926: note <= 13722;
                6927: note <= 15491;
                6928: note <= 14886;
                6929: note <= 12187;
                6930: note <= 8192;
                6931: note <= 3995;
                6932: note <= 697;
                6933: note <= (-893);
                6934: note <= (-467);
                6935: note <= 1697;
                6936: note <= 4815;
                6937: note <= 7815;
                6938: note <= 9626;
                6939: note <= 9474;
                6940: note <= 7094;
                6941: note <= 2814;
                6942: note <= (-2531);
                6943: note <= (-7815);
                6944: note <= (-11910);
                6945: note <= (-13985);
                6946: note <= (-13722);
                6947: note <= (-11395);
                6948: note <= (-7791);
                6949: note <= (-3995);
                6950: note <= (-1098);
                6951: note <= 101;
                6952: note <= (-697);
                6953: note <= (-3203);
                6954: note <= (-6627);
                6955: note <= (-9889);
                6956: note <= (-11910);
                6957: note <= (-11911);
                6958: note <= (-9626);
                6959: note <= (-5378);
                6960: note <= 0;
                6961: note <= 5378;
                6962: note <= 9626;
                6963: note <= 11911;
                6964: note <= 11910;
                6965: note <= 9889;
                6966: note <= 6627;
                6967: note <= 3203;
                6968: note <= 697;
                6969: note <= (-101);
                6970: note <= 1098;
                6971: note <= 3995;
                6972: note <= 7791;
                6973: note <= 11395;
                6974: note <= 13722;
                6975: note <= 13985;
                6976: note <= 11910;
                6977: note <= 7815;
                6978: note <= 2531;
                6979: note <= (-2814);
                6980: note <= (-7094);
                6981: note <= (-9474);
                6982: note <= (-9626);
                6983: note <= (-7815);
                6984: note <= (-4815);
                6985: note <= (-1697);
                6986: note <= 467;
                6987: note <= 893;
                6988: note <= (-697);
                6989: note <= (-3995);
                6990: note <= (-8192);
                6991: note <= (-12187);
                6992: note <= (-14886);
                6993: note <= (-15491);
                6994: note <= (-13722);
                6995: note <= (-9889);
                6996: note <= (-4815);
                6997: note <= 377;
                6998: note <= 4563;
                6999: note <= 6910;
                7000: note <= 7094;
                7001: note <= 5378;
                7002: note <= 2531;
                7003: note <= (-377);
                7004: note <= (-2279);
                7005: note <= (-2399);
                7006: note <= (-467);
                7007: note <= 3203;
                7008: note <= 7791;
                7009: note <= 12187;
                7010: note <= 15286;
                7011: note <= 16283;
                7012: note <= 14886;
                7013: note <= 11395;
                7014: note <= 6627;
                7015: note <= 1697;
                7016: note <= (-2279);
                7017: note <= (-4473);
                7018: note <= (-4563);
                7019: note <= (-2814);
                7020: note <= 0;
                7021: note <= 2814;
                7022: note <= 4563;
                7023: note <= 4473;
                7024: note <= 2279;
                7025: note <= (-1697);
                7026: note <= (-6627);
                7027: note <= (-11395);
                7028: note <= (-14886);
                7029: note <= (-16283);
                7030: note <= (-15286);
                7031: note <= (-12187);
                7032: note <= (-7791);
                7033: note <= (-3203);
                7034: note <= 467;
                7035: note <= 2399;
                7036: note <= 2279;
                7037: note <= 377;
                7038: note <= (-2531);
                7039: note <= (-5378);
                7040: note <= (-7094);
                7041: note <= (-6910);
                7042: note <= (-4563);
                7043: note <= (-377);
                7044: note <= 4815;
                7045: note <= 9889;
                7046: note <= 13722;
                7047: note <= 15491;
                7048: note <= 14886;
                7049: note <= 12187;
                7050: note <= 8192;
                7051: note <= 3995;
                7052: note <= 697;
                7053: note <= (-893);
                7054: note <= (-467);
                7055: note <= 1697;
                7056: note <= 4815;
                7057: note <= 7815;
                7058: note <= 9626;
                7059: note <= 9474;
                7060: note <= 7094;
                7061: note <= 2814;
                7062: note <= (-2531);
                7063: note <= (-7815);
                7064: note <= (-11910);
                7065: note <= (-13985);
                7066: note <= (-13722);
                7067: note <= (-11395);
                7068: note <= (-7791);
                7069: note <= (-3995);
                7070: note <= (-1098);
                7071: note <= 101;
                7072: note <= (-697);
                7073: note <= (-3203);
                7074: note <= (-6627);
                7075: note <= (-9889);
                7076: note <= (-11910);
                7077: note <= (-11911);
                7078: note <= (-9626);
                7079: note <= (-5378);
                7080: note <= 0;
                7081: note <= 5378;
                7082: note <= 9626;
                7083: note <= 11911;
                7084: note <= 11910;
                7085: note <= 9889;
                7086: note <= 6627;
                7087: note <= 3203;
                7088: note <= 697;
                7089: note <= (-101);
                7090: note <= 1098;
                7091: note <= 3995;
                7092: note <= 7791;
                7093: note <= 11395;
                7094: note <= 13722;
                7095: note <= 13985;
                7096: note <= 11910;
                7097: note <= 7815;
                7098: note <= 2531;
                7099: note <= (-2814);
                7100: note <= (-7094);
                7101: note <= (-9474);
                7102: note <= (-9626);
                7103: note <= (-7815);
                7104: note <= (-4815);
                7105: note <= (-1697);
                7106: note <= 467;
                7107: note <= 893;
                7108: note <= (-697);
                7109: note <= (-3995);
                7110: note <= (-8192);
                7111: note <= (-12187);
                7112: note <= (-14886);
                7113: note <= (-15491);
                7114: note <= (-13722);
                7115: note <= (-9889);
                7116: note <= (-4815);
                7117: note <= 377;
                7118: note <= 4563;
                7119: note <= 6910;
                7120: note <= 7094;
                7121: note <= 5378;
                7122: note <= 2531;
                7123: note <= (-377);
                7124: note <= (-2279);
                7125: note <= (-2399);
                7126: note <= (-467);
                7127: note <= 3203;
                7128: note <= 7791;
                7129: note <= 12187;
                7130: note <= 15286;
                7131: note <= 16283;
                7132: note <= 14886;
                7133: note <= 11395;
                7134: note <= 6627;
                7135: note <= 1697;
                7136: note <= (-2279);
                7137: note <= (-4473);
                7138: note <= (-4563);
                7139: note <= (-2814);
                7140: note <= 0;
                7141: note <= 2814;
                7142: note <= 4563;
                7143: note <= 4473;
                7144: note <= 2279;
                7145: note <= (-1697);
                7146: note <= (-6627);
                7147: note <= (-11395);
                7148: note <= (-14886);
                7149: note <= (-16283);
                7150: note <= (-15286);
                7151: note <= (-12187);
                7152: note <= (-7791);
                7153: note <= (-3203);
                7154: note <= 467;
                7155: note <= 2399;
                7156: note <= 2279;
                7157: note <= 377;
                7158: note <= (-2531);
                7159: note <= (-5378);
                7160: note <= (-7094);
                7161: note <= (-6910);
                7162: note <= (-4563);
                7163: note <= (-377);
                7164: note <= 4815;
                7165: note <= 9889;
                7166: note <= 13722;
                7167: note <= 15491;
                7168: note <= 14886;
                7169: note <= 12187;
                7170: note <= 8192;
                7171: note <= 3995;
                7172: note <= 697;
                7173: note <= (-893);
                7174: note <= (-467);
                7175: note <= 1697;
                7176: note <= 4815;
                7177: note <= 7815;
                7178: note <= 9626;
                7179: note <= 9474;
                7180: note <= 7094;
                7181: note <= 2814;
                7182: note <= (-2531);
                7183: note <= (-7815);
                7184: note <= (-11910);
                7185: note <= (-13985);
                7186: note <= (-13722);
                7187: note <= (-11395);
                7188: note <= (-7791);
                7189: note <= (-3995);
                7190: note <= (-1098);
                7191: note <= 101;
                7192: note <= (-697);
                7193: note <= (-3203);
                7194: note <= (-6627);
                7195: note <= (-9889);
                7196: note <= (-11910);
                7197: note <= (-11911);
                7198: note <= (-9626);
                7199: note <= (-5378);
                7200: note <= 0;
                7201: note <= 5378;
                7202: note <= 9626;
                7203: note <= 11911;
                7204: note <= 11910;
                7205: note <= 9889;
                7206: note <= 6627;
                7207: note <= 3203;
                7208: note <= 697;
                7209: note <= (-101);
                7210: note <= 1098;
                7211: note <= 3995;
                7212: note <= 7791;
                7213: note <= 11395;
                7214: note <= 13722;
                7215: note <= 13985;
                7216: note <= 11910;
                7217: note <= 7815;
                7218: note <= 2531;
                7219: note <= (-2814);
                7220: note <= (-7094);
                7221: note <= (-9474);
                7222: note <= (-9626);
                7223: note <= (-7815);
                7224: note <= (-4815);
                7225: note <= (-1697);
                7226: note <= 467;
                7227: note <= 893;
                7228: note <= (-697);
                7229: note <= (-3995);
                7230: note <= (-8192);
                7231: note <= (-12187);
                7232: note <= (-14886);
                7233: note <= (-15491);
                7234: note <= (-13722);
                7235: note <= (-9889);
                7236: note <= (-4815);
                7237: note <= 377;
                7238: note <= 4563;
                7239: note <= 6910;
                7240: note <= 7094;
                7241: note <= 5378;
                7242: note <= 2531;
                7243: note <= (-377);
                7244: note <= (-2279);
                7245: note <= (-2399);
                7246: note <= (-467);
                7247: note <= 3203;
                7248: note <= 7791;
                7249: note <= 12187;
                7250: note <= 15286;
                7251: note <= 16283;
                7252: note <= 14886;
                7253: note <= 11395;
                7254: note <= 6627;
                7255: note <= 1697;
                7256: note <= (-2279);
                7257: note <= (-4473);
                7258: note <= (-4563);
                7259: note <= (-2814);
                7260: note <= 0;
                7261: note <= 2814;
                7262: note <= 4563;
                7263: note <= 4473;
                7264: note <= 2279;
                7265: note <= (-1697);
                7266: note <= (-6627);
                7267: note <= (-11395);
                7268: note <= (-14886);
                7269: note <= (-16283);
                7270: note <= (-15286);
                7271: note <= (-12187);
                7272: note <= (-7791);
                7273: note <= (-3203);
                7274: note <= 467;
                7275: note <= 2399;
                7276: note <= 2279;
                7277: note <= 377;
                7278: note <= (-2531);
                7279: note <= (-5378);
                7280: note <= (-7094);
                7281: note <= (-6910);
                7282: note <= (-4563);
                7283: note <= (-377);
                7284: note <= 4815;
                7285: note <= 9889;
                7286: note <= 13722;
                7287: note <= 15491;
                7288: note <= 14886;
                7289: note <= 12187;
                7290: note <= 8192;
                7291: note <= 3995;
                7292: note <= 697;
                7293: note <= (-893);
                7294: note <= (-467);
                7295: note <= 1697;
                7296: note <= 4815;
                7297: note <= 7815;
                7298: note <= 9626;
                7299: note <= 9474;
                7300: note <= 7094;
                7301: note <= 2814;
                7302: note <= (-2531);
                7303: note <= (-7815);
                7304: note <= (-11910);
                7305: note <= (-13985);
                7306: note <= (-13722);
                7307: note <= (-11395);
                7308: note <= (-7791);
                7309: note <= (-3995);
                7310: note <= (-1098);
                7311: note <= 101;
                7312: note <= (-697);
                7313: note <= (-3203);
                7314: note <= (-6627);
                7315: note <= (-9889);
                7316: note <= (-11910);
                7317: note <= (-11911);
                7318: note <= (-9626);
                7319: note <= (-5378);
                7320: note <= 0;
                7321: note <= 5378;
                7322: note <= 9626;
                7323: note <= 11911;
                7324: note <= 11910;
                7325: note <= 9889;
                7326: note <= 6627;
                7327: note <= 3203;
                7328: note <= 697;
                7329: note <= (-101);
                7330: note <= 1098;
                7331: note <= 3995;
                7332: note <= 7791;
                7333: note <= 11395;
                7334: note <= 13722;
                7335: note <= 13985;
                7336: note <= 11910;
                7337: note <= 7815;
                7338: note <= 2531;
                7339: note <= (-2814);
                7340: note <= (-7094);
                7341: note <= (-9474);
                7342: note <= (-9626);
                7343: note <= (-7815);
                7344: note <= (-4815);
                7345: note <= (-1697);
                7346: note <= 467;
                7347: note <= 893;
                7348: note <= (-697);
                7349: note <= (-3995);
                7350: note <= (-8192);
                7351: note <= (-12187);
                7352: note <= (-14886);
                7353: note <= (-15491);
                7354: note <= (-13722);
                7355: note <= (-9889);
                7356: note <= (-4815);
                7357: note <= 377;
                7358: note <= 4563;
                7359: note <= 6910;
                7360: note <= 7094;
                7361: note <= 5378;
                7362: note <= 2531;
                7363: note <= (-377);
                7364: note <= (-2279);
                7365: note <= (-2399);
                7366: note <= (-467);
                7367: note <= 3203;
                7368: note <= 7791;
                7369: note <= 12187;
                7370: note <= 15286;
                7371: note <= 16283;
                7372: note <= 14886;
                7373: note <= 11395;
                7374: note <= 6627;
                7375: note <= 1697;
                7376: note <= (-2279);
                7377: note <= (-4473);
                7378: note <= (-4563);
                7379: note <= (-2814);
                7380: note <= 0;
                7381: note <= 2814;
                7382: note <= 4563;
                7383: note <= 4473;
                7384: note <= 2279;
                7385: note <= (-1697);
                7386: note <= (-6627);
                7387: note <= (-11395);
                7388: note <= (-14886);
                7389: note <= (-16283);
                7390: note <= (-15286);
                7391: note <= (-12187);
                7392: note <= (-7791);
                7393: note <= (-3203);
                7394: note <= 467;
                7395: note <= 2399;
                7396: note <= 2279;
                7397: note <= 377;
                7398: note <= (-2531);
                7399: note <= (-5378);
                7400: note <= (-7094);
                7401: note <= (-6910);
                7402: note <= (-4563);
                7403: note <= (-377);
                7404: note <= 4815;
                7405: note <= 9889;
                7406: note <= 13722;
                7407: note <= 15491;
                7408: note <= 14886;
                7409: note <= 12187;
                7410: note <= 8192;
                7411: note <= 3995;
                7412: note <= 697;
                7413: note <= (-893);
                7414: note <= (-467);
                7415: note <= 1697;
                7416: note <= 4815;
                7417: note <= 7815;
                7418: note <= 9626;
                7419: note <= 9474;
                7420: note <= 7094;
                7421: note <= 2814;
                7422: note <= (-2531);
                7423: note <= (-7815);
                7424: note <= (-11910);
                7425: note <= (-13985);
                7426: note <= (-13722);
                7427: note <= (-11395);
                7428: note <= (-7791);
                7429: note <= (-3995);
                7430: note <= (-1098);
                7431: note <= 101;
                7432: note <= (-697);
                7433: note <= (-3203);
                7434: note <= (-6627);
                7435: note <= (-9889);
                7436: note <= (-11910);
                7437: note <= (-11911);
                7438: note <= (-9626);
                7439: note <= (-5378);
                7440: note <= 0;
                7441: note <= 5378;
                7442: note <= 9626;
                7443: note <= 11911;
                7444: note <= 11910;
                7445: note <= 9889;
                7446: note <= 6627;
                7447: note <= 3203;
                7448: note <= 697;
                7449: note <= (-101);
                7450: note <= 1098;
                7451: note <= 3995;
                7452: note <= 7791;
                7453: note <= 11395;
                7454: note <= 13722;
                7455: note <= 13985;
                7456: note <= 11910;
                7457: note <= 7815;
                7458: note <= 2531;
                7459: note <= (-2814);
                7460: note <= (-7094);
                7461: note <= (-9474);
                7462: note <= (-9626);
                7463: note <= (-7815);
                7464: note <= (-4815);
                7465: note <= (-1697);
                7466: note <= 467;
                7467: note <= 893;
                7468: note <= (-697);
                7469: note <= (-3995);
                7470: note <= (-8192);
                7471: note <= (-12187);
                7472: note <= (-14886);
                7473: note <= (-15491);
                7474: note <= (-13722);
                7475: note <= (-9889);
                7476: note <= (-4815);
                7477: note <= 377;
                7478: note <= 4563;
                7479: note <= 6910;
                7480: note <= 7094;
                7481: note <= 5378;
                7482: note <= 2531;
                7483: note <= (-377);
                7484: note <= (-2279);
                7485: note <= (-2399);
                7486: note <= (-467);
                7487: note <= 3203;
                7488: note <= 7791;
                7489: note <= 12187;
                7490: note <= 15286;
                7491: note <= 16283;
                7492: note <= 14886;
                7493: note <= 11395;
                7494: note <= 6627;
                7495: note <= 1697;
                7496: note <= (-2279);
                7497: note <= (-4473);
                7498: note <= (-4563);
                7499: note <= (-2814);
                7500: note <= 0;
                7501: note <= 2814;
                7502: note <= 4563;
                7503: note <= 4473;
                7504: note <= 2279;
                7505: note <= (-1697);
                7506: note <= (-6627);
                7507: note <= (-11395);
                7508: note <= (-14886);
                7509: note <= (-16283);
                7510: note <= (-15286);
                7511: note <= (-12187);
                7512: note <= (-7791);
                7513: note <= (-3203);
                7514: note <= 467;
                7515: note <= 2399;
                7516: note <= 2279;
                7517: note <= 377;
                7518: note <= (-2531);
                7519: note <= (-5378);
                7520: note <= (-7094);
                7521: note <= (-6910);
                7522: note <= (-4563);
                7523: note <= (-377);
                7524: note <= 4815;
                7525: note <= 9889;
                7526: note <= 13722;
                7527: note <= 15491;
                7528: note <= 14886;
                7529: note <= 12187;
                7530: note <= 8192;
                7531: note <= 3995;
                7532: note <= 697;
                7533: note <= (-893);
                7534: note <= (-467);
                7535: note <= 1697;
                7536: note <= 4815;
                7537: note <= 7815;
                7538: note <= 9626;
                7539: note <= 9474;
                7540: note <= 7094;
                7541: note <= 2814;
                7542: note <= (-2531);
                7543: note <= (-7815);
                7544: note <= (-11910);
                7545: note <= (-13985);
                7546: note <= (-13722);
                7547: note <= (-11395);
                7548: note <= (-7791);
                7549: note <= (-3995);
                7550: note <= (-1098);
                7551: note <= 101;
                7552: note <= (-697);
                7553: note <= (-3203);
                7554: note <= (-6627);
                7555: note <= (-9889);
                7556: note <= (-11910);
                7557: note <= (-11911);
                7558: note <= (-9626);
                7559: note <= (-5378);
                7560: note <= 0;
                7561: note <= 5378;
                7562: note <= 9626;
                7563: note <= 11911;
                7564: note <= 11910;
                7565: note <= 9889;
                7566: note <= 6627;
                7567: note <= 3203;
                7568: note <= 697;
                7569: note <= (-101);
                7570: note <= 1098;
                7571: note <= 3995;
                7572: note <= 7791;
                7573: note <= 11395;
                7574: note <= 13722;
                7575: note <= 13985;
                7576: note <= 11910;
                7577: note <= 7815;
                7578: note <= 2531;
                7579: note <= (-2814);
                7580: note <= (-7094);
                7581: note <= (-9474);
                7582: note <= (-9626);
                7583: note <= (-7815);
                7584: note <= (-4815);
                7585: note <= (-1697);
                7586: note <= 467;
                7587: note <= 893;
                7588: note <= (-697);
                7589: note <= (-3995);
                7590: note <= (-8192);
                7591: note <= (-12187);
                7592: note <= (-14886);
                7593: note <= (-15491);
                7594: note <= (-13722);
                7595: note <= (-9889);
                7596: note <= (-4815);
                7597: note <= 377;
                7598: note <= 4563;
                7599: note <= 6910;
                7600: note <= 7094;
                7601: note <= 5378;
                7602: note <= 2531;
                7603: note <= (-377);
                7604: note <= (-2279);
                7605: note <= (-2399);
                7606: note <= (-467);
                7607: note <= 3203;
                7608: note <= 7791;
                7609: note <= 12187;
                7610: note <= 15286;
                7611: note <= 16283;
                7612: note <= 14886;
                7613: note <= 11395;
                7614: note <= 6627;
                7615: note <= 1697;
                7616: note <= (-2279);
                7617: note <= (-4473);
                7618: note <= (-4563);
                7619: note <= (-2814);
                7620: note <= 0;
                7621: note <= 2814;
                7622: note <= 4563;
                7623: note <= 4473;
                7624: note <= 2279;
                7625: note <= (-1697);
                7626: note <= (-6627);
                7627: note <= (-11395);
                7628: note <= (-14886);
                7629: note <= (-16283);
                7630: note <= (-15286);
                7631: note <= (-12187);
                7632: note <= (-7791);
                7633: note <= (-3203);
                7634: note <= 467;
                7635: note <= 2399;
                7636: note <= 2279;
                7637: note <= 377;
                7638: note <= (-2531);
                7639: note <= (-5378);
                7640: note <= (-7094);
                7641: note <= (-6910);
                7642: note <= (-4563);
                7643: note <= (-377);
                7644: note <= 4815;
                7645: note <= 9889;
                7646: note <= 13722;
                7647: note <= 15491;
                7648: note <= 14886;
                7649: note <= 12187;
                7650: note <= 8192;
                7651: note <= 3995;
                7652: note <= 697;
                7653: note <= (-893);
                7654: note <= (-467);
                7655: note <= 1697;
                7656: note <= 4815;
                7657: note <= 7815;
                7658: note <= 9626;
                7659: note <= 9474;
                7660: note <= 7094;
                7661: note <= 2814;
                7662: note <= (-2531);
                7663: note <= (-7815);
                7664: note <= (-11910);
                7665: note <= (-13985);
                7666: note <= (-13722);
                7667: note <= (-11395);
                7668: note <= (-7791);
                7669: note <= (-3995);
                7670: note <= (-1098);
                7671: note <= 101;
                7672: note <= (-697);
                7673: note <= (-3203);
                7674: note <= (-6627);
                7675: note <= (-9889);
                7676: note <= (-11910);
                7677: note <= (-11911);
                7678: note <= (-9626);
                7679: note <= (-5378);
                7680: note <= 0;
                7681: note <= 5378;
                7682: note <= 9626;
                7683: note <= 11911;
                7684: note <= 11910;
                7685: note <= 9889;
                7686: note <= 6627;
                7687: note <= 3203;
                7688: note <= 697;
                7689: note <= (-101);
                7690: note <= 1098;
                7691: note <= 3995;
                7692: note <= 7791;
                7693: note <= 11395;
                7694: note <= 13722;
                7695: note <= 13985;
                7696: note <= 11910;
                7697: note <= 7815;
                7698: note <= 2531;
                7699: note <= (-2814);
                7700: note <= (-7094);
                7701: note <= (-9474);
                7702: note <= (-9626);
                7703: note <= (-7815);
                7704: note <= (-4815);
                7705: note <= (-1697);
                7706: note <= 467;
                7707: note <= 893;
                7708: note <= (-697);
                7709: note <= (-3995);
                7710: note <= (-8192);
                7711: note <= (-12187);
                7712: note <= (-14886);
                7713: note <= (-15491);
                7714: note <= (-13722);
                7715: note <= (-9889);
                7716: note <= (-4815);
                7717: note <= 377;
                7718: note <= 4563;
                7719: note <= 6910;
                7720: note <= 7094;
                7721: note <= 5378;
                7722: note <= 2531;
                7723: note <= (-377);
                7724: note <= (-2279);
                7725: note <= (-2399);
                7726: note <= (-467);
                7727: note <= 3203;
                7728: note <= 7791;
                7729: note <= 12187;
                7730: note <= 15286;
                7731: note <= 16283;
                7732: note <= 14886;
                7733: note <= 11395;
                7734: note <= 6627;
                7735: note <= 1697;
                7736: note <= (-2279);
                7737: note <= (-4473);
                7738: note <= (-4563);
                7739: note <= (-2814);
                7740: note <= 0;
                7741: note <= 2814;
                7742: note <= 4563;
                7743: note <= 4473;
                7744: note <= 2279;
                7745: note <= (-1697);
                7746: note <= (-6627);
                7747: note <= (-11395);
                7748: note <= (-14886);
                7749: note <= (-16283);
                7750: note <= (-15286);
                7751: note <= (-12187);
                7752: note <= (-7791);
                7753: note <= (-3203);
                7754: note <= 467;
                7755: note <= 2399;
                7756: note <= 2279;
                7757: note <= 377;
                7758: note <= (-2531);
                7759: note <= (-5378);
                7760: note <= (-7094);
                7761: note <= (-6910);
                7762: note <= (-4563);
                7763: note <= (-377);
                7764: note <= 4815;
                7765: note <= 9889;
                7766: note <= 13722;
                7767: note <= 15491;
                7768: note <= 14886;
                7769: note <= 12187;
                7770: note <= 8192;
                7771: note <= 3995;
                7772: note <= 697;
                7773: note <= (-893);
                7774: note <= (-467);
                7775: note <= 1697;
                7776: note <= 4815;
                7777: note <= 7815;
                7778: note <= 9626;
                7779: note <= 9474;
                7780: note <= 7094;
                7781: note <= 2814;
                7782: note <= (-2531);
                7783: note <= (-7815);
                7784: note <= (-11910);
                7785: note <= (-13985);
                7786: note <= (-13722);
                7787: note <= (-11395);
                7788: note <= (-7791);
                7789: note <= (-3995);
                7790: note <= (-1098);
                7791: note <= 101;
                7792: note <= (-697);
                7793: note <= (-3203);
                7794: note <= (-6627);
                7795: note <= (-9889);
                7796: note <= (-11910);
                7797: note <= (-11911);
                7798: note <= (-9626);
                7799: note <= (-5378);
                7800: note <= 0;
                7801: note <= 5378;
                7802: note <= 9626;
                7803: note <= 11911;
                7804: note <= 11910;
                7805: note <= 9889;
                7806: note <= 6627;
                7807: note <= 3203;
                7808: note <= 697;
                7809: note <= (-101);
                7810: note <= 1098;
                7811: note <= 3995;
                7812: note <= 7791;
                7813: note <= 11395;
                7814: note <= 13722;
                7815: note <= 13985;
                7816: note <= 11910;
                7817: note <= 7815;
                7818: note <= 2531;
                7819: note <= (-2814);
                7820: note <= (-7094);
                7821: note <= (-9474);
                7822: note <= (-9626);
                7823: note <= (-7815);
                7824: note <= (-4815);
                7825: note <= (-1697);
                7826: note <= 467;
                7827: note <= 893;
                7828: note <= (-697);
                7829: note <= (-3995);
                7830: note <= (-8192);
                7831: note <= (-12187);
                7832: note <= (-14886);
                7833: note <= (-15491);
                7834: note <= (-13722);
                7835: note <= (-9889);
                7836: note <= (-4815);
                7837: note <= 377;
                7838: note <= 4563;
                7839: note <= 6910;
                7840: note <= 7094;
                7841: note <= 5378;
                7842: note <= 2531;
                7843: note <= (-377);
                7844: note <= (-2279);
                7845: note <= (-2399);
                7846: note <= (-467);
                7847: note <= 3203;
                7848: note <= 7791;
                7849: note <= 12187;
                7850: note <= 15286;
                7851: note <= 16283;
                7852: note <= 14886;
                7853: note <= 11395;
                7854: note <= 6627;
                7855: note <= 1697;
                7856: note <= (-2279);
                7857: note <= (-4473);
                7858: note <= (-4563);
                7859: note <= (-2814);
                7860: note <= 0;
                7861: note <= 2814;
                7862: note <= 4563;
                7863: note <= 4473;
                7864: note <= 2279;
                7865: note <= (-1697);
                7866: note <= (-6627);
                7867: note <= (-11395);
                7868: note <= (-14886);
                7869: note <= (-16283);
                7870: note <= (-15286);
                7871: note <= (-12187);
                7872: note <= (-7791);
                7873: note <= (-3203);
                7874: note <= 467;
                7875: note <= 2399;
                7876: note <= 2279;
                7877: note <= 377;
                7878: note <= (-2531);
                7879: note <= (-5378);
                7880: note <= (-7094);
                7881: note <= (-6910);
                7882: note <= (-4563);
                7883: note <= (-377);
                7884: note <= 4815;
                7885: note <= 9889;
                7886: note <= 13722;
                7887: note <= 15491;
                7888: note <= 14886;
                7889: note <= 12187;
                7890: note <= 8192;
                7891: note <= 3995;
                7892: note <= 697;
                7893: note <= (-893);
                7894: note <= (-467);
                7895: note <= 1697;
                7896: note <= 4815;
                7897: note <= 7815;
                7898: note <= 9626;
                7899: note <= 9474;
                7900: note <= 7094;
                7901: note <= 2814;
                7902: note <= (-2531);
                7903: note <= (-7815);
                7904: note <= (-11910);
                7905: note <= (-13985);
                7906: note <= (-13722);
                7907: note <= (-11395);
                7908: note <= (-7791);
                7909: note <= (-3995);
                7910: note <= (-1098);
                7911: note <= 101;
                7912: note <= (-697);
                7913: note <= (-3203);
                7914: note <= (-6627);
                7915: note <= (-9889);
                7916: note <= (-11910);
                7917: note <= (-11911);
                7918: note <= (-9626);
                7919: note <= (-5378);
                7920: note <= 0;
                7921: note <= 5378;
                7922: note <= 9626;
                7923: note <= 11911;
                7924: note <= 11910;
                7925: note <= 9889;
                7926: note <= 6627;
                7927: note <= 3203;
                7928: note <= 697;
                7929: note <= (-101);
                7930: note <= 1098;
                7931: note <= 3995;
                7932: note <= 7791;
                7933: note <= 11395;
                7934: note <= 13722;
                7935: note <= 13985;
                7936: note <= 11910;
                7937: note <= 7815;
                7938: note <= 2531;
                7939: note <= (-2814);
                7940: note <= (-7094);
                7941: note <= (-9474);
                7942: note <= (-9626);
                7943: note <= (-7815);
                7944: note <= (-4815);
                7945: note <= (-1697);
                7946: note <= 467;
                7947: note <= 893;
                7948: note <= (-697);
                7949: note <= (-3995);
                7950: note <= (-8192);
                7951: note <= (-12187);
                7952: note <= (-14886);
                7953: note <= (-15491);
                7954: note <= (-13722);
                7955: note <= (-9889);
                7956: note <= (-4815);
                7957: note <= 377;
                7958: note <= 4563;
                7959: note <= 6910;
                7960: note <= 7094;
                7961: note <= 5378;
                7962: note <= 2531;
                7963: note <= (-377);
                7964: note <= (-2279);
                7965: note <= (-2399);
                7966: note <= (-467);
                7967: note <= 3203;
                7968: note <= 7791;
                7969: note <= 12187;
                7970: note <= 15286;
                7971: note <= 16283;
                7972: note <= 14886;
                7973: note <= 11395;
                7974: note <= 6627;
                7975: note <= 1697;
                7976: note <= (-2279);
                7977: note <= (-4473);
                7978: note <= (-4563);
                7979: note <= (-2814);
                7980: note <= 0;
                7981: note <= 2814;
                7982: note <= 4563;
                7983: note <= 4473;
                7984: note <= 2279;
                7985: note <= (-1697);
                7986: note <= (-6627);
                7987: note <= (-11395);
                7988: note <= (-14886);
                7989: note <= (-16283);
                7990: note <= (-15286);
                7991: note <= (-12187);
                7992: note <= (-7791);
                7993: note <= (-3203);
                7994: note <= 467;
                7995: note <= 2399;
                7996: note <= 2279;
                7997: note <= 377;
                7998: note <= (-2531);
                7999: note <= (-5378);
                8000: note <= (-7094);
                8001: note <= (-6910);
                8002: note <= (-4563);
                8003: note <= (-377);
                8004: note <= 4815;
                8005: note <= 9889;
                8006: note <= 13722;
                8007: note <= 15491;
                8008: note <= 14886;
                8009: note <= 12187;
                8010: note <= 8192;
                8011: note <= 3995;
                8012: note <= 697;
                8013: note <= (-893);
                8014: note <= (-467);
                8015: note <= 1697;
                8016: note <= 4815;
                8017: note <= 7815;
                8018: note <= 9626;
                8019: note <= 9474;
                8020: note <= 7094;
                8021: note <= 2814;
                8022: note <= (-2531);
                8023: note <= (-7815);
                8024: note <= (-11910);
                8025: note <= (-13985);
                8026: note <= (-13722);
                8027: note <= (-11395);
                8028: note <= (-7791);
                8029: note <= (-3995);
                8030: note <= (-1098);
                8031: note <= 101;
                8032: note <= (-697);
                8033: note <= (-3203);
                8034: note <= (-6627);
                8035: note <= (-9889);
                8036: note <= (-11910);
                8037: note <= (-11911);
                8038: note <= (-9626);
                8039: note <= (-5378);
                8040: note <= 0;
                8041: note <= 5378;
                8042: note <= 9626;
                8043: note <= 11911;
                8044: note <= 11910;
                8045: note <= 9889;
                8046: note <= 6627;
                8047: note <= 3203;
                8048: note <= 697;
                8049: note <= (-101);
                8050: note <= 1098;
                8051: note <= 3995;
                8052: note <= 7791;
                8053: note <= 11395;
                8054: note <= 13722;
                8055: note <= 13985;
                8056: note <= 11910;
                8057: note <= 7815;
                8058: note <= 2531;
                8059: note <= (-2814);
                8060: note <= (-7094);
                8061: note <= (-9474);
                8062: note <= (-9626);
                8063: note <= (-7815);
                8064: note <= (-4815);
                8065: note <= (-1697);
                8066: note <= 467;
                8067: note <= 893;
                8068: note <= (-697);
                8069: note <= (-3995);
                8070: note <= (-8192);
                8071: note <= (-12187);
                8072: note <= (-14886);
                8073: note <= (-15491);
                8074: note <= (-13722);
                8075: note <= (-9889);
                8076: note <= (-4815);
                8077: note <= 377;
                8078: note <= 4563;
                8079: note <= 6910;
                8080: note <= 7094;
                8081: note <= 5378;
                8082: note <= 2531;
                8083: note <= (-377);
                8084: note <= (-2279);
                8085: note <= (-2399);
                8086: note <= (-467);
                8087: note <= 3203;
                8088: note <= 7791;
                8089: note <= 12187;
                8090: note <= 15286;
                8091: note <= 16283;
                8092: note <= 14886;
                8093: note <= 11395;
                8094: note <= 6627;
                8095: note <= 1697;
                8096: note <= (-2279);
                8097: note <= (-4473);
                8098: note <= (-4563);
                8099: note <= (-2814);
                8100: note <= 0;
                8101: note <= 2814;
                8102: note <= 4563;
                8103: note <= 4473;
                8104: note <= 2279;
                8105: note <= (-1697);
                8106: note <= (-6627);
                8107: note <= (-11395);
                8108: note <= (-14886);
                8109: note <= (-16283);
                8110: note <= (-15286);
                8111: note <= (-12187);
                8112: note <= (-7791);
                8113: note <= (-3203);
                8114: note <= 467;
                8115: note <= 2399;
                8116: note <= 2279;
                8117: note <= 377;
                8118: note <= (-2531);
                8119: note <= (-5378);
                8120: note <= (-7094);
                8121: note <= (-6910);
                8122: note <= (-4563);
                8123: note <= (-377);
                8124: note <= 4815;
                8125: note <= 9889;
                8126: note <= 13722;
                8127: note <= 15491;
                8128: note <= 14886;
                8129: note <= 12187;
                8130: note <= 8192;
                8131: note <= 3995;
                8132: note <= 697;
                8133: note <= (-893);
                8134: note <= (-467);
                8135: note <= 1697;
                8136: note <= 4815;
                8137: note <= 7815;
                8138: note <= 9626;
                8139: note <= 9474;
                8140: note <= 7094;
                8141: note <= 2814;
                8142: note <= (-2531);
                8143: note <= (-7815);
                8144: note <= (-11910);
                8145: note <= (-13985);
                8146: note <= (-13722);
                8147: note <= (-11395);
                8148: note <= (-7791);
                8149: note <= (-3995);
                8150: note <= (-1098);
                8151: note <= 101;
                8152: note <= (-697);
                8153: note <= (-3203);
                8154: note <= (-6627);
                8155: note <= (-9889);
                8156: note <= (-11910);
                8157: note <= (-11911);
                8158: note <= (-9626);
                8159: note <= (-5378);
                8160: note <= 0;
                8161: note <= 5378;
                8162: note <= 9626;
                8163: note <= 11911;
                8164: note <= 11910;
                8165: note <= 9889;
                8166: note <= 6627;
                8167: note <= 3203;
                8168: note <= 697;
                8169: note <= (-101);
                8170: note <= 1098;
                8171: note <= 3995;
                8172: note <= 7791;
                8173: note <= 11395;
                8174: note <= 13722;
                8175: note <= 13985;
                8176: note <= 11910;
                8177: note <= 7815;
                8178: note <= 2531;
                8179: note <= (-2814);
                8180: note <= (-7094);
                8181: note <= (-9474);
                8182: note <= (-9626);
                8183: note <= (-7815);
                8184: note <= (-4815);
                8185: note <= (-1697);
                8186: note <= 467;
                8187: note <= 893;
                8188: note <= (-697);
                8189: note <= (-3995);
                8190: note <= (-8192);
                8191: note <= (-12187);
                8192: note <= (-14886);
                8193: note <= (-15491);
                8194: note <= (-13722);
                8195: note <= (-9889);
                8196: note <= (-4815);
                8197: note <= 377;
                8198: note <= 4563;
                8199: note <= 6910;
                8200: note <= 7094;
                8201: note <= 5378;
                8202: note <= 2531;
                8203: note <= (-377);
                8204: note <= (-2279);
                8205: note <= (-2399);
                8206: note <= (-467);
                8207: note <= 3203;
                8208: note <= 7791;
                8209: note <= 12187;
                8210: note <= 15286;
                8211: note <= 16283;
                8212: note <= 14886;
                8213: note <= 11395;
                8214: note <= 6627;
                8215: note <= 1697;
                8216: note <= (-2279);
                8217: note <= (-4473);
                8218: note <= (-4563);
                8219: note <= (-2814);
                8220: note <= 0;
                8221: note <= 2814;
                8222: note <= 4563;
                8223: note <= 4473;
                8224: note <= 2279;
                8225: note <= (-1697);
                8226: note <= (-6627);
                8227: note <= (-11395);
                8228: note <= (-14886);
                8229: note <= (-16283);
                8230: note <= (-15286);
                8231: note <= (-12187);
                8232: note <= (-7791);
                8233: note <= (-3203);
                8234: note <= 467;
                8235: note <= 2399;
                8236: note <= 2279;
                8237: note <= 377;
                8238: note <= (-2531);
                8239: note <= (-5378);
                8240: note <= (-7094);
                8241: note <= (-6910);
                8242: note <= (-4563);
                8243: note <= (-377);
                8244: note <= 4815;
                8245: note <= 9889;
                8246: note <= 13722;
                8247: note <= 15491;
                8248: note <= 14886;
                8249: note <= 12187;
                8250: note <= 8192;
                8251: note <= 3995;
                8252: note <= 697;
                8253: note <= (-893);
                8254: note <= (-467);
                8255: note <= 1697;
                8256: note <= 4815;
                8257: note <= 7815;
                8258: note <= 9626;
                8259: note <= 9474;
                8260: note <= 7094;
                8261: note <= 2814;
                8262: note <= (-2531);
                8263: note <= (-7815);
                8264: note <= (-11910);
                8265: note <= (-13985);
                8266: note <= (-13722);
                8267: note <= (-11395);
                8268: note <= (-7791);
                8269: note <= (-3995);
                8270: note <= (-1098);
                8271: note <= 101;
                8272: note <= (-697);
                8273: note <= (-3203);
                8274: note <= (-6627);
                8275: note <= (-9889);
                8276: note <= (-11910);
                8277: note <= (-11911);
                8278: note <= (-9626);
                8279: note <= (-5378);
                8280: note <= 0;
                8281: note <= 5378;
                8282: note <= 9626;
                8283: note <= 11911;
                8284: note <= 11910;
                8285: note <= 9889;
                8286: note <= 6627;
                8287: note <= 3203;
                8288: note <= 697;
                8289: note <= (-101);
                8290: note <= 1098;
                8291: note <= 3995;
                8292: note <= 7791;
                8293: note <= 11395;
                8294: note <= 13722;
                8295: note <= 13985;
                8296: note <= 11910;
                8297: note <= 7815;
                8298: note <= 2531;
                8299: note <= (-2814);
                8300: note <= (-7094);
                8301: note <= (-9474);
                8302: note <= (-9626);
                8303: note <= (-7815);
                8304: note <= (-4815);
                8305: note <= (-1697);
                8306: note <= 467;
                8307: note <= 893;
                8308: note <= (-697);
                8309: note <= (-3995);
                8310: note <= (-8192);
                8311: note <= (-12187);
                8312: note <= (-14886);
                8313: note <= (-15491);
                8314: note <= (-13722);
                8315: note <= (-9889);
                8316: note <= (-4815);
                8317: note <= 377;
                8318: note <= 4563;
                8319: note <= 6910;
                8320: note <= 7094;
                8321: note <= 5378;
                8322: note <= 2531;
                8323: note <= (-377);
                8324: note <= (-2279);
                8325: note <= (-2399);
                8326: note <= (-467);
                8327: note <= 3203;
                8328: note <= 7791;
                8329: note <= 12187;
                8330: note <= 15286;
                8331: note <= 16283;
                8332: note <= 14886;
                8333: note <= 11395;
                8334: note <= 6627;
                8335: note <= 1697;
                8336: note <= (-2279);
                8337: note <= (-4473);
                8338: note <= (-4563);
                8339: note <= (-2814);
                8340: note <= 0;
                8341: note <= 2814;
                8342: note <= 4563;
                8343: note <= 4473;
                8344: note <= 2279;
                8345: note <= (-1697);
                8346: note <= (-6627);
                8347: note <= (-11395);
                8348: note <= (-14886);
                8349: note <= (-16283);
                8350: note <= (-15286);
                8351: note <= (-12187);
                8352: note <= (-7791);
                8353: note <= (-3203);
                8354: note <= 467;
                8355: note <= 2399;
                8356: note <= 2279;
                8357: note <= 377;
                8358: note <= (-2531);
                8359: note <= (-5378);
                8360: note <= (-7094);
                8361: note <= (-6910);
                8362: note <= (-4563);
                8363: note <= (-377);
                8364: note <= 4815;
                8365: note <= 9889;
                8366: note <= 13722;
                8367: note <= 15491;
                8368: note <= 14886;
                8369: note <= 12187;
                8370: note <= 8192;
                8371: note <= 3995;
                8372: note <= 697;
                8373: note <= (-893);
                8374: note <= (-467);
                8375: note <= 1697;
                8376: note <= 4815;
                8377: note <= 7815;
                8378: note <= 9626;
                8379: note <= 9474;
                8380: note <= 7094;
                8381: note <= 2814;
                8382: note <= (-2531);
                8383: note <= (-7815);
                8384: note <= (-11910);
                8385: note <= (-13985);
                8386: note <= (-13722);
                8387: note <= (-11395);
                8388: note <= (-7791);
                8389: note <= (-3995);
                8390: note <= (-1098);
                8391: note <= 101;
                8392: note <= (-697);
                8393: note <= (-3203);
                8394: note <= (-6627);
                8395: note <= (-9889);
                8396: note <= (-11910);
                8397: note <= (-11911);
                8398: note <= (-9626);
                8399: note <= (-5378);
                8400: note <= 0;
                8401: note <= 5378;
                8402: note <= 9626;
                8403: note <= 11911;
                8404: note <= 11910;
                8405: note <= 9889;
                8406: note <= 6627;
                8407: note <= 3203;
                8408: note <= 697;
                8409: note <= (-101);
                8410: note <= 1098;
                8411: note <= 3995;
                8412: note <= 7791;
                8413: note <= 11395;
                8414: note <= 13722;
                8415: note <= 13985;
                8416: note <= 11910;
                8417: note <= 7815;
                8418: note <= 2531;
                8419: note <= (-2814);
                8420: note <= (-7094);
                8421: note <= (-9474);
                8422: note <= (-9626);
                8423: note <= (-7815);
                8424: note <= (-4815);
                8425: note <= (-1697);
                8426: note <= 467;
                8427: note <= 893;
                8428: note <= (-697);
                8429: note <= (-3995);
                8430: note <= (-8192);
                8431: note <= (-12187);
                8432: note <= (-14886);
                8433: note <= (-15491);
                8434: note <= (-13722);
                8435: note <= (-9889);
                8436: note <= (-4815);
                8437: note <= 377;
                8438: note <= 4563;
                8439: note <= 6910;
                8440: note <= 7094;
                8441: note <= 5378;
                8442: note <= 2531;
                8443: note <= (-377);
                8444: note <= (-2279);
                8445: note <= (-2399);
                8446: note <= (-467);
                8447: note <= 3203;
                8448: note <= 7791;
                8449: note <= 12187;
                8450: note <= 15286;
                8451: note <= 16283;
                8452: note <= 14886;
                8453: note <= 11395;
                8454: note <= 6627;
                8455: note <= 1697;
                8456: note <= (-2279);
                8457: note <= (-4473);
                8458: note <= (-4563);
                8459: note <= (-2814);
                8460: note <= 0;
                8461: note <= 2814;
                8462: note <= 4563;
                8463: note <= 4473;
                8464: note <= 2279;
                8465: note <= (-1697);
                8466: note <= (-6627);
                8467: note <= (-11395);
                8468: note <= (-14886);
                8469: note <= (-16283);
                8470: note <= (-15286);
                8471: note <= (-12187);
                8472: note <= (-7791);
                8473: note <= (-3203);
                8474: note <= 467;
                8475: note <= 2399;
                8476: note <= 2279;
                8477: note <= 377;
                8478: note <= (-2531);
                8479: note <= (-5378);
                8480: note <= (-7094);
                8481: note <= (-6910);
                8482: note <= (-4563);
                8483: note <= (-377);
                8484: note <= 4815;
                8485: note <= 9889;
                8486: note <= 13722;
                8487: note <= 15491;
                8488: note <= 14886;
                8489: note <= 12187;
                8490: note <= 8192;
                8491: note <= 3995;
                8492: note <= 697;
                8493: note <= (-893);
                8494: note <= (-467);
                8495: note <= 1697;
                8496: note <= 4815;
                8497: note <= 7815;
                8498: note <= 9626;
                8499: note <= 9474;
                8500: note <= 7094;
                8501: note <= 2814;
                8502: note <= (-2531);
                8503: note <= (-7815);
                8504: note <= (-11910);
                8505: note <= (-13985);
                8506: note <= (-13722);
                8507: note <= (-11395);
                8508: note <= (-7791);
                8509: note <= (-3995);
                8510: note <= (-1098);
                8511: note <= 101;
                8512: note <= (-697);
                8513: note <= (-3203);
                8514: note <= (-6627);
                8515: note <= (-9889);
                8516: note <= (-11910);
                8517: note <= (-11911);
                8518: note <= (-9626);
                8519: note <= (-5378);
                8520: note <= 0;
                8521: note <= 5378;
                8522: note <= 9626;
                8523: note <= 11911;
                8524: note <= 11910;
                8525: note <= 9889;
                8526: note <= 6627;
                8527: note <= 3203;
                8528: note <= 697;
                8529: note <= (-101);
                8530: note <= 1098;
                8531: note <= 3995;
                8532: note <= 7791;
                8533: note <= 11395;
                8534: note <= 13722;
                8535: note <= 13985;
                8536: note <= 11910;
                8537: note <= 7815;
                8538: note <= 2531;
                8539: note <= (-2814);
                8540: note <= (-7094);
                8541: note <= (-9474);
                8542: note <= (-9626);
                8543: note <= (-7815);
                8544: note <= (-4815);
                8545: note <= (-1697);
                8546: note <= 467;
                8547: note <= 893;
                8548: note <= (-697);
                8549: note <= (-3995);
                8550: note <= (-8192);
                8551: note <= (-12187);
                8552: note <= (-14886);
                8553: note <= (-15491);
                8554: note <= (-13722);
                8555: note <= (-9889);
                8556: note <= (-4815);
                8557: note <= 377;
                8558: note <= 4563;
                8559: note <= 6910;
                8560: note <= 7094;
                8561: note <= 5378;
                8562: note <= 2531;
                8563: note <= (-377);
                8564: note <= (-2279);
                8565: note <= (-2399);
                8566: note <= (-467);
                8567: note <= 3203;
                8568: note <= 7791;
                8569: note <= 12187;
                8570: note <= 15286;
                8571: note <= 16283;
                8572: note <= 14886;
                8573: note <= 11395;
                8574: note <= 6627;
                8575: note <= 1697;
                8576: note <= (-2279);
                8577: note <= (-4473);
                8578: note <= (-4563);
                8579: note <= (-2814);
                8580: note <= 0;
                8581: note <= 2814;
                8582: note <= 4563;
                8583: note <= 4473;
                8584: note <= 2279;
                8585: note <= (-1697);
                8586: note <= (-6627);
                8587: note <= (-11395);
                8588: note <= (-14886);
                8589: note <= (-16283);
                8590: note <= (-15286);
                8591: note <= (-12187);
                8592: note <= (-7791);
                8593: note <= (-3203);
                8594: note <= 467;
                8595: note <= 2399;
                8596: note <= 2279;
                8597: note <= 377;
                8598: note <= (-2531);
                8599: note <= (-5378);
                8600: note <= (-7094);
                8601: note <= (-6910);
                8602: note <= (-4563);
                8603: note <= (-377);
                8604: note <= 4815;
                8605: note <= 9889;
                8606: note <= 13722;
                8607: note <= 15491;
                8608: note <= 14886;
                8609: note <= 12187;
                8610: note <= 8192;
                8611: note <= 3995;
                8612: note <= 697;
                8613: note <= (-893);
                8614: note <= (-467);
                8615: note <= 1697;
                8616: note <= 4815;
                8617: note <= 7815;
                8618: note <= 9626;
                8619: note <= 9474;
                8620: note <= 7094;
                8621: note <= 2814;
                8622: note <= (-2531);
                8623: note <= (-7815);
                8624: note <= (-11910);
                8625: note <= (-13985);
                8626: note <= (-13722);
                8627: note <= (-11395);
                8628: note <= (-7791);
                8629: note <= (-3995);
                8630: note <= (-1098);
                8631: note <= 101;
                8632: note <= (-697);
                8633: note <= (-3203);
                8634: note <= (-6627);
                8635: note <= (-9889);
                8636: note <= (-11910);
                8637: note <= (-11911);
                8638: note <= (-9626);
                8639: note <= (-5378);
                8640: note <= 0;
                8641: note <= 5378;
                8642: note <= 9626;
                8643: note <= 11911;
                8644: note <= 11910;
                8645: note <= 9889;
                8646: note <= 6627;
                8647: note <= 3203;
                8648: note <= 697;
                8649: note <= (-101);
                8650: note <= 1098;
                8651: note <= 3995;
                8652: note <= 7791;
                8653: note <= 11395;
                8654: note <= 13722;
                8655: note <= 13985;
                8656: note <= 11910;
                8657: note <= 7815;
                8658: note <= 2531;
                8659: note <= (-2814);
                8660: note <= (-7094);
                8661: note <= (-9474);
                8662: note <= (-9626);
                8663: note <= (-7815);
                8664: note <= (-4815);
                8665: note <= (-1697);
                8666: note <= 467;
                8667: note <= 893;
                8668: note <= (-697);
                8669: note <= (-3995);
                8670: note <= (-8192);
                8671: note <= (-12187);
                8672: note <= (-14886);
                8673: note <= (-15491);
                8674: note <= (-13722);
                8675: note <= (-9889);
                8676: note <= (-4815);
                8677: note <= 377;
                8678: note <= 4563;
                8679: note <= 6910;
                8680: note <= 7094;
                8681: note <= 5378;
                8682: note <= 2531;
                8683: note <= (-377);
                8684: note <= (-2279);
                8685: note <= (-2399);
                8686: note <= (-467);
                8687: note <= 3203;
                8688: note <= 7791;
                8689: note <= 12187;
                8690: note <= 15286;
                8691: note <= 16283;
                8692: note <= 14886;
                8693: note <= 11395;
                8694: note <= 6627;
                8695: note <= 1697;
                8696: note <= (-2279);
                8697: note <= (-4473);
                8698: note <= (-4563);
                8699: note <= (-2814);
                8700: note <= 0;
                8701: note <= 2814;
                8702: note <= 4563;
                8703: note <= 4473;
                8704: note <= 2279;
                8705: note <= (-1697);
                8706: note <= (-6627);
                8707: note <= (-11395);
                8708: note <= (-14886);
                8709: note <= (-16283);
                8710: note <= (-15286);
                8711: note <= (-12187);
                8712: note <= (-7791);
                8713: note <= (-3203);
                8714: note <= 467;
                8715: note <= 2399;
                8716: note <= 2279;
                8717: note <= 377;
                8718: note <= (-2531);
                8719: note <= (-5378);
                8720: note <= (-7094);
                8721: note <= (-6910);
                8722: note <= (-4563);
                8723: note <= (-377);
                8724: note <= 4815;
                8725: note <= 9889;
                8726: note <= 13722;
                8727: note <= 15491;
                8728: note <= 14886;
                8729: note <= 12187;
                8730: note <= 8192;
                8731: note <= 3995;
                8732: note <= 697;
                8733: note <= (-893);
                8734: note <= (-467);
                8735: note <= 1697;
                8736: note <= 4815;
                8737: note <= 7815;
                8738: note <= 9626;
                8739: note <= 9474;
                8740: note <= 7094;
                8741: note <= 2814;
                8742: note <= (-2531);
                8743: note <= (-7815);
                8744: note <= (-11910);
                8745: note <= (-13985);
                8746: note <= (-13722);
                8747: note <= (-11395);
                8748: note <= (-7791);
                8749: note <= (-3995);
                8750: note <= (-1098);
                8751: note <= 101;
                8752: note <= (-697);
                8753: note <= (-3203);
                8754: note <= (-6627);
                8755: note <= (-9889);
                8756: note <= (-11910);
                8757: note <= (-11911);
                8758: note <= (-9626);
                8759: note <= (-5378);
                8760: note <= 0;
                8761: note <= 5378;
                8762: note <= 9626;
                8763: note <= 11911;
                8764: note <= 11910;
                8765: note <= 9889;
                8766: note <= 6627;
                8767: note <= 3203;
                8768: note <= 697;
                8769: note <= (-101);
                8770: note <= 1098;
                8771: note <= 3995;
                8772: note <= 7791;
                8773: note <= 11395;
                8774: note <= 13722;
                8775: note <= 13985;
                8776: note <= 11910;
                8777: note <= 7815;
                8778: note <= 2531;
                8779: note <= (-2814);
                8780: note <= (-7094);
                8781: note <= (-9474);
                8782: note <= (-9626);
                8783: note <= (-7815);
                8784: note <= (-4815);
                8785: note <= (-1697);
                8786: note <= 467;
                8787: note <= 893;
                8788: note <= (-697);
                8789: note <= (-3995);
                8790: note <= (-8192);
                8791: note <= (-12187);
                8792: note <= (-14886);
                8793: note <= (-15491);
                8794: note <= (-13722);
                8795: note <= (-9889);
                8796: note <= (-4815);
                8797: note <= 377;
                8798: note <= 4563;
                8799: note <= 6910;
                8800: note <= 7094;
                8801: note <= 5378;
                8802: note <= 2531;
                8803: note <= (-377);
                8804: note <= (-2279);
                8805: note <= (-2399);
                8806: note <= (-467);
                8807: note <= 3203;
                8808: note <= 7791;
                8809: note <= 12187;
                8810: note <= 15286;
                8811: note <= 16283;
                8812: note <= 14886;
                8813: note <= 11395;
                8814: note <= 6627;
                8815: note <= 1697;
                8816: note <= (-2279);
                8817: note <= (-4473);
                8818: note <= (-4563);
                8819: note <= (-2814);
                8820: note <= 0;
                8821: note <= 2814;
                8822: note <= 4563;
                8823: note <= 4473;
                8824: note <= 2279;
                8825: note <= (-1697);
                8826: note <= (-6627);
                8827: note <= (-11395);
                8828: note <= (-14886);
                8829: note <= (-16283);
                8830: note <= (-15286);
                8831: note <= (-12187);
                8832: note <= (-7791);
                8833: note <= (-3203);
                8834: note <= 467;
                8835: note <= 2399;
                8836: note <= 2279;
                8837: note <= 377;
                8838: note <= (-2531);
                8839: note <= (-5378);
                8840: note <= (-7094);
                8841: note <= (-6910);
                8842: note <= (-4563);
                8843: note <= (-377);
                8844: note <= 4815;
                8845: note <= 9889;
                8846: note <= 13722;
                8847: note <= 15491;
                8848: note <= 14886;
                8849: note <= 12187;
                8850: note <= 8192;
                8851: note <= 3995;
                8852: note <= 697;
                8853: note <= (-893);
                8854: note <= (-467);
                8855: note <= 1697;
                8856: note <= 4815;
                8857: note <= 7815;
                8858: note <= 9626;
                8859: note <= 9474;
                8860: note <= 7094;
                8861: note <= 2814;
                8862: note <= (-2531);
                8863: note <= (-7815);
                8864: note <= (-11910);
                8865: note <= (-13985);
                8866: note <= (-13722);
                8867: note <= (-11395);
                8868: note <= (-7791);
                8869: note <= (-3995);
                8870: note <= (-1098);
                8871: note <= 101;
                8872: note <= (-697);
                8873: note <= (-3203);
                8874: note <= (-6627);
                8875: note <= (-9889);
                8876: note <= (-11910);
                8877: note <= (-11911);
                8878: note <= (-9626);
                8879: note <= (-5378);
                8880: note <= 0;
                8881: note <= 5378;
                8882: note <= 9626;
                8883: note <= 11911;
                8884: note <= 11910;
                8885: note <= 9889;
                8886: note <= 6627;
                8887: note <= 3203;
                8888: note <= 697;
                8889: note <= (-101);
                8890: note <= 1098;
                8891: note <= 3995;
                8892: note <= 7791;
                8893: note <= 11395;
                8894: note <= 13722;
                8895: note <= 13985;
                8896: note <= 11910;
                8897: note <= 7815;
                8898: note <= 2531;
                8899: note <= (-2814);
                8900: note <= (-7094);
                8901: note <= (-9474);
                8902: note <= (-9626);
                8903: note <= (-7815);
                8904: note <= (-4815);
                8905: note <= (-1697);
                8906: note <= 467;
                8907: note <= 893;
                8908: note <= (-697);
                8909: note <= (-3995);
                8910: note <= (-8192);
                8911: note <= (-12187);
                8912: note <= (-14886);
                8913: note <= (-15491);
                8914: note <= (-13722);
                8915: note <= (-9889);
                8916: note <= (-4815);
                8917: note <= 377;
                8918: note <= 4563;
                8919: note <= 6910;
                8920: note <= 7094;
                8921: note <= 5378;
                8922: note <= 2531;
                8923: note <= (-377);
                8924: note <= (-2279);
                8925: note <= (-2399);
                8926: note <= (-467);
                8927: note <= 3203;
                8928: note <= 7791;
                8929: note <= 12187;
                8930: note <= 15286;
                8931: note <= 16283;
                8932: note <= 14886;
                8933: note <= 11395;
                8934: note <= 6627;
                8935: note <= 1697;
                8936: note <= (-2279);
                8937: note <= (-4473);
                8938: note <= (-4563);
                8939: note <= (-2814);
                8940: note <= 0;
                8941: note <= 2814;
                8942: note <= 4563;
                8943: note <= 4473;
                8944: note <= 2279;
                8945: note <= (-1697);
                8946: note <= (-6627);
                8947: note <= (-11395);
                8948: note <= (-14886);
                8949: note <= (-16283);
                8950: note <= (-15286);
                8951: note <= (-12187);
                8952: note <= (-7791);
                8953: note <= (-3203);
                8954: note <= 467;
                8955: note <= 2399;
                8956: note <= 2279;
                8957: note <= 377;
                8958: note <= (-2531);
                8959: note <= (-5378);
                8960: note <= (-7094);
                8961: note <= (-6910);
                8962: note <= (-4563);
                8963: note <= (-377);
                8964: note <= 4815;
                8965: note <= 9889;
                8966: note <= 13722;
                8967: note <= 15491;
                8968: note <= 14886;
                8969: note <= 12187;
                8970: note <= 8192;
                8971: note <= 3995;
                8972: note <= 697;
                8973: note <= (-893);
                8974: note <= (-467);
                8975: note <= 1697;
                8976: note <= 4815;
                8977: note <= 7815;
                8978: note <= 9626;
                8979: note <= 9474;
                8980: note <= 7094;
                8981: note <= 2814;
                8982: note <= (-2531);
                8983: note <= (-7815);
                8984: note <= (-11910);
                8985: note <= (-13985);
                8986: note <= (-13722);
                8987: note <= (-11395);
                8988: note <= (-7791);
                8989: note <= (-3995);
                8990: note <= (-1098);
                8991: note <= 101;
                8992: note <= (-697);
                8993: note <= (-3203);
                8994: note <= (-6627);
                8995: note <= (-9889);
                8996: note <= (-11910);
                8997: note <= (-11911);
                8998: note <= (-9626);
                8999: note <= (-5378);
                9000: note <= 0;
                9001: note <= 5378;
                9002: note <= 9626;
                9003: note <= 11911;
                9004: note <= 11910;
                9005: note <= 9889;
                9006: note <= 6627;
                9007: note <= 3203;
                9008: note <= 697;
                9009: note <= (-101);
                9010: note <= 1098;
                9011: note <= 3995;
                9012: note <= 7791;
                9013: note <= 11395;
                9014: note <= 13722;
                9015: note <= 13985;
                9016: note <= 11910;
                9017: note <= 7815;
                9018: note <= 2531;
                9019: note <= (-2814);
                9020: note <= (-7094);
                9021: note <= (-9474);
                9022: note <= (-9626);
                9023: note <= (-7815);
                9024: note <= (-4815);
                9025: note <= (-1697);
                9026: note <= 467;
                9027: note <= 893;
                9028: note <= (-697);
                9029: note <= (-3995);
                9030: note <= (-8192);
                9031: note <= (-12187);
                9032: note <= (-14886);
                9033: note <= (-15491);
                9034: note <= (-13722);
                9035: note <= (-9889);
                9036: note <= (-4815);
                9037: note <= 377;
                9038: note <= 4563;
                9039: note <= 6910;
                9040: note <= 7094;
                9041: note <= 5378;
                9042: note <= 2531;
                9043: note <= (-377);
                9044: note <= (-2279);
                9045: note <= (-2399);
                9046: note <= (-467);
                9047: note <= 3203;
                9048: note <= 7791;
                9049: note <= 12187;
                9050: note <= 15286;
                9051: note <= 16283;
                9052: note <= 14886;
                9053: note <= 11395;
                9054: note <= 6627;
                9055: note <= 1697;
                9056: note <= (-2279);
                9057: note <= (-4473);
                9058: note <= (-4563);
                9059: note <= (-2814);
                9060: note <= 0;
                9061: note <= 2814;
                9062: note <= 4563;
                9063: note <= 4473;
                9064: note <= 2279;
                9065: note <= (-1697);
                9066: note <= (-6627);
                9067: note <= (-11395);
                9068: note <= (-14886);
                9069: note <= (-16283);
                9070: note <= (-15286);
                9071: note <= (-12187);
                9072: note <= (-7791);
                9073: note <= (-3203);
                9074: note <= 467;
                9075: note <= 2399;
                9076: note <= 2279;
                9077: note <= 377;
                9078: note <= (-2531);
                9079: note <= (-5378);
                9080: note <= (-7094);
                9081: note <= (-6910);
                9082: note <= (-4563);
                9083: note <= (-377);
                9084: note <= 4815;
                9085: note <= 9889;
                9086: note <= 13722;
                9087: note <= 15491;
                9088: note <= 14886;
                9089: note <= 12187;
                9090: note <= 8192;
                9091: note <= 3995;
                9092: note <= 697;
                9093: note <= (-893);
                9094: note <= (-467);
                9095: note <= 1697;
                9096: note <= 4815;
                9097: note <= 7815;
                9098: note <= 9626;
                9099: note <= 9474;
                9100: note <= 7094;
                9101: note <= 2814;
                9102: note <= (-2531);
                9103: note <= (-7815);
                9104: note <= (-11910);
                9105: note <= (-13985);
                9106: note <= (-13722);
                9107: note <= (-11395);
                9108: note <= (-7791);
                9109: note <= (-3995);
                9110: note <= (-1098);
                9111: note <= 101;
                9112: note <= (-697);
                9113: note <= (-3203);
                9114: note <= (-6627);
                9115: note <= (-9889);
                9116: note <= (-11910);
                9117: note <= (-11911);
                9118: note <= (-9626);
                9119: note <= (-5378);
                9120: note <= 0;
                9121: note <= 5378;
                9122: note <= 9626;
                9123: note <= 11911;
                9124: note <= 11910;
                9125: note <= 9889;
                9126: note <= 6627;
                9127: note <= 3203;
                9128: note <= 697;
                9129: note <= (-101);
                9130: note <= 1098;
                9131: note <= 3995;
                9132: note <= 7791;
                9133: note <= 11395;
                9134: note <= 13722;
                9135: note <= 13985;
                9136: note <= 11910;
                9137: note <= 7815;
                9138: note <= 2531;
                9139: note <= (-2814);
                9140: note <= (-7094);
                9141: note <= (-9474);
                9142: note <= (-9626);
                9143: note <= (-7815);
                9144: note <= (-4815);
                9145: note <= (-1697);
                9146: note <= 467;
                9147: note <= 893;
                9148: note <= (-697);
                9149: note <= (-3995);
                9150: note <= (-8192);
                9151: note <= (-12187);
                9152: note <= (-14886);
                9153: note <= (-15491);
                9154: note <= (-13722);
                9155: note <= (-9889);
                9156: note <= (-4815);
                9157: note <= 377;
                9158: note <= 4563;
                9159: note <= 6910;
                9160: note <= 7094;
                9161: note <= 5378;
                9162: note <= 2531;
                9163: note <= (-377);
                9164: note <= (-2279);
                9165: note <= (-2399);
                9166: note <= (-467);
                9167: note <= 3203;
                9168: note <= 7791;
                9169: note <= 12187;
                9170: note <= 15286;
                9171: note <= 16283;
                9172: note <= 14886;
                9173: note <= 11395;
                9174: note <= 6627;
                9175: note <= 1697;
                9176: note <= (-2279);
                9177: note <= (-4473);
                9178: note <= (-4563);
                9179: note <= (-2814);
                9180: note <= 0;
                9181: note <= 2814;
                9182: note <= 4563;
                9183: note <= 4473;
                9184: note <= 2279;
                9185: note <= (-1697);
                9186: note <= (-6627);
                9187: note <= (-11395);
                9188: note <= (-14886);
                9189: note <= (-16283);
                9190: note <= (-15286);
                9191: note <= (-12187);
                9192: note <= (-7791);
                9193: note <= (-3203);
                9194: note <= 467;
                9195: note <= 2399;
                9196: note <= 2279;
                9197: note <= 377;
                9198: note <= (-2531);
                9199: note <= (-5378);
                9200: note <= (-7094);
                9201: note <= (-6910);
                9202: note <= (-4563);
                9203: note <= (-377);
                9204: note <= 4815;
                9205: note <= 9889;
                9206: note <= 13722;
                9207: note <= 15491;
                9208: note <= 14886;
                9209: note <= 12187;
                9210: note <= 8192;
                9211: note <= 3995;
                9212: note <= 697;
                9213: note <= (-893);
                9214: note <= (-467);
                9215: note <= 1697;
                9216: note <= 4815;
                9217: note <= 7815;
                9218: note <= 9626;
                9219: note <= 9474;
                9220: note <= 7094;
                9221: note <= 2814;
                9222: note <= (-2531);
                9223: note <= (-7815);
                9224: note <= (-11910);
                9225: note <= (-13985);
                9226: note <= (-13722);
                9227: note <= (-11395);
                9228: note <= (-7791);
                9229: note <= (-3995);
                9230: note <= (-1098);
                9231: note <= 101;
                9232: note <= (-697);
                9233: note <= (-3203);
                9234: note <= (-6627);
                9235: note <= (-9889);
                9236: note <= (-11910);
                9237: note <= (-11911);
                9238: note <= (-9626);
                9239: note <= (-5378);
                9240: note <= 0;
                9241: note <= 5378;
                9242: note <= 9626;
                9243: note <= 11911;
                9244: note <= 11910;
                9245: note <= 9889;
                9246: note <= 6627;
                9247: note <= 3203;
                9248: note <= 697;
                9249: note <= (-101);
                9250: note <= 1098;
                9251: note <= 3995;
                9252: note <= 7791;
                9253: note <= 11395;
                9254: note <= 13722;
                9255: note <= 13985;
                9256: note <= 11910;
                9257: note <= 7815;
                9258: note <= 2531;
                9259: note <= (-2814);
                9260: note <= (-7094);
                9261: note <= (-9474);
                9262: note <= (-9626);
                9263: note <= (-7815);
                9264: note <= (-4815);
                9265: note <= (-1697);
                9266: note <= 467;
                9267: note <= 893;
                9268: note <= (-697);
                9269: note <= (-3995);
                9270: note <= (-8192);
                9271: note <= (-12187);
                9272: note <= (-14886);
                9273: note <= (-15491);
                9274: note <= (-13722);
                9275: note <= (-9889);
                9276: note <= (-4815);
                9277: note <= 377;
                9278: note <= 4563;
                9279: note <= 6910;
                9280: note <= 7094;
                9281: note <= 5378;
                9282: note <= 2531;
                9283: note <= (-377);
                9284: note <= (-2279);
                9285: note <= (-2399);
                9286: note <= (-467);
                9287: note <= 3203;
                9288: note <= 7791;
                9289: note <= 12187;
                9290: note <= 15286;
                9291: note <= 16283;
                9292: note <= 14886;
                9293: note <= 11395;
                9294: note <= 6627;
                9295: note <= 1697;
                9296: note <= (-2279);
                9297: note <= (-4473);
                9298: note <= (-4563);
                9299: note <= (-2814);
                9300: note <= 0;
                9301: note <= 2814;
                9302: note <= 4563;
                9303: note <= 4473;
                9304: note <= 2279;
                9305: note <= (-1697);
                9306: note <= (-6627);
                9307: note <= (-11395);
                9308: note <= (-14886);
                9309: note <= (-16283);
                9310: note <= (-15286);
                9311: note <= (-12187);
                9312: note <= (-7791);
                9313: note <= (-3203);
                9314: note <= 467;
                9315: note <= 2399;
                9316: note <= 2279;
                9317: note <= 377;
                9318: note <= (-2531);
                9319: note <= (-5378);
                9320: note <= (-7094);
                9321: note <= (-6910);
                9322: note <= (-4563);
                9323: note <= (-377);
                9324: note <= 4815;
                9325: note <= 9889;
                9326: note <= 13722;
                9327: note <= 15491;
                9328: note <= 14886;
                9329: note <= 12187;
                9330: note <= 8192;
                9331: note <= 3995;
                9332: note <= 697;
                9333: note <= (-893);
                9334: note <= (-467);
                9335: note <= 1697;
                9336: note <= 4815;
                9337: note <= 7815;
                9338: note <= 9626;
                9339: note <= 9474;
                9340: note <= 7094;
                9341: note <= 2814;
                9342: note <= (-2531);
                9343: note <= (-7815);
                9344: note <= (-11910);
                9345: note <= (-13985);
                9346: note <= (-13722);
                9347: note <= (-11395);
                9348: note <= (-7791);
                9349: note <= (-3995);
                9350: note <= (-1098);
                9351: note <= 101;
                9352: note <= (-697);
                9353: note <= (-3203);
                9354: note <= (-6627);
                9355: note <= (-9889);
                9356: note <= (-11910);
                9357: note <= (-11911);
                9358: note <= (-9626);
                9359: note <= (-5378);
                9360: note <= 0;
                9361: note <= 5378;
                9362: note <= 9626;
                9363: note <= 11911;
                9364: note <= 11910;
                9365: note <= 9889;
                9366: note <= 6627;
                9367: note <= 3203;
                9368: note <= 697;
                9369: note <= (-101);
                9370: note <= 1098;
                9371: note <= 3995;
                9372: note <= 7791;
                9373: note <= 11395;
                9374: note <= 13722;
                9375: note <= 13985;
                9376: note <= 11910;
                9377: note <= 7815;
                9378: note <= 2531;
                9379: note <= (-2814);
                9380: note <= (-7094);
                9381: note <= (-9474);
                9382: note <= (-9626);
                9383: note <= (-7815);
                9384: note <= (-4815);
                9385: note <= (-1697);
                9386: note <= 467;
                9387: note <= 893;
                9388: note <= (-697);
                9389: note <= (-3995);
                9390: note <= (-8192);
                9391: note <= (-12187);
                9392: note <= (-14886);
                9393: note <= (-15491);
                9394: note <= (-13722);
                9395: note <= (-9889);
                9396: note <= (-4815);
                9397: note <= 377;
                9398: note <= 4563;
                9399: note <= 6910;
                9400: note <= 7094;
                9401: note <= 5378;
                9402: note <= 2531;
                9403: note <= (-377);
                9404: note <= (-2279);
                9405: note <= (-2399);
                9406: note <= (-467);
                9407: note <= 3203;
                9408: note <= 7791;
                9409: note <= 12187;
                9410: note <= 15286;
                9411: note <= 16283;
                9412: note <= 14886;
                9413: note <= 11395;
                9414: note <= 6627;
                9415: note <= 1697;
                9416: note <= (-2279);
                9417: note <= (-4473);
                9418: note <= (-4563);
                9419: note <= (-2814);
                9420: note <= 0;
                9421: note <= 2814;
                9422: note <= 4563;
                9423: note <= 4473;
                9424: note <= 2279;
                9425: note <= (-1697);
                9426: note <= (-6627);
                9427: note <= (-11395);
                9428: note <= (-14886);
                9429: note <= (-16283);
                9430: note <= (-15286);
                9431: note <= (-12187);
                9432: note <= (-7791);
                9433: note <= (-3203);
                9434: note <= 467;
                9435: note <= 2399;
                9436: note <= 2279;
                9437: note <= 377;
                9438: note <= (-2531);
                9439: note <= (-5378);
                9440: note <= (-7094);
                9441: note <= (-6910);
                9442: note <= (-4563);
                9443: note <= (-377);
                9444: note <= 4815;
                9445: note <= 9889;
                9446: note <= 13722;
                9447: note <= 15491;
                9448: note <= 14886;
                9449: note <= 12187;
                9450: note <= 8192;
                9451: note <= 3995;
                9452: note <= 697;
                9453: note <= (-893);
                9454: note <= (-467);
                9455: note <= 1697;
                9456: note <= 4815;
                9457: note <= 7815;
                9458: note <= 9626;
                9459: note <= 9474;
                9460: note <= 7094;
                9461: note <= 2814;
                9462: note <= (-2531);
                9463: note <= (-7815);
                9464: note <= (-11910);
                9465: note <= (-13985);
                9466: note <= (-13722);
                9467: note <= (-11395);
                9468: note <= (-7791);
                9469: note <= (-3995);
                9470: note <= (-1098);
                9471: note <= 101;
                9472: note <= (-697);
                9473: note <= (-3203);
                9474: note <= (-6627);
                9475: note <= (-9889);
                9476: note <= (-11910);
                9477: note <= (-11911);
                9478: note <= (-9626);
                9479: note <= (-5378);
                9480: note <= 0;
                9481: note <= 5378;
                9482: note <= 9626;
                9483: note <= 11911;
                9484: note <= 11910;
                9485: note <= 9889;
                9486: note <= 6627;
                9487: note <= 3203;
                9488: note <= 697;
                9489: note <= (-101);
                9490: note <= 1098;
                9491: note <= 3995;
                9492: note <= 7791;
                9493: note <= 11395;
                9494: note <= 13722;
                9495: note <= 13985;
                9496: note <= 11910;
                9497: note <= 7815;
                9498: note <= 2531;
                9499: note <= (-2814);
                9500: note <= (-7094);
                9501: note <= (-9474);
                9502: note <= (-9626);
                9503: note <= (-7815);
                9504: note <= (-4815);
                9505: note <= (-1697);
                9506: note <= 467;
                9507: note <= 893;
                9508: note <= (-697);
                9509: note <= (-3995);
                9510: note <= (-8192);
                9511: note <= (-12187);
                9512: note <= (-14886);
                9513: note <= (-15491);
                9514: note <= (-13722);
                9515: note <= (-9889);
                9516: note <= (-4815);
                9517: note <= 377;
                9518: note <= 4563;
                9519: note <= 6910;
                9520: note <= 7094;
                9521: note <= 5378;
                9522: note <= 2531;
                9523: note <= (-377);
                9524: note <= (-2279);
                9525: note <= (-2399);
                9526: note <= (-467);
                9527: note <= 3203;
                9528: note <= 7791;
                9529: note <= 12187;
                9530: note <= 15286;
                9531: note <= 16283;
                9532: note <= 14886;
                9533: note <= 11395;
                9534: note <= 6627;
                9535: note <= 1697;
                9536: note <= (-2279);
                9537: note <= (-4473);
                9538: note <= (-4563);
                9539: note <= (-2814);
                9540: note <= 0;
                9541: note <= 2814;
                9542: note <= 4563;
                9543: note <= 4473;
                9544: note <= 2279;
                9545: note <= (-1697);
                9546: note <= (-6627);
                9547: note <= (-11395);
                9548: note <= (-14886);
                9549: note <= (-16283);
                9550: note <= (-15286);
                9551: note <= (-12187);
                9552: note <= (-7791);
                9553: note <= (-3203);
                9554: note <= 467;
                9555: note <= 2399;
                9556: note <= 2279;
                9557: note <= 377;
                9558: note <= (-2531);
                9559: note <= (-5378);
                9560: note <= (-7094);
                9561: note <= (-6910);
                9562: note <= (-4563);
                9563: note <= (-377);
                9564: note <= 4815;
                9565: note <= 9889;
                9566: note <= 13722;
                9567: note <= 15491;
                9568: note <= 14886;
                9569: note <= 12187;
                9570: note <= 8192;
                9571: note <= 3995;
                9572: note <= 697;
                9573: note <= (-893);
                9574: note <= (-467);
                9575: note <= 1697;
                9576: note <= 4815;
                9577: note <= 7815;
                9578: note <= 9626;
                9579: note <= 9474;
                9580: note <= 7094;
                9581: note <= 2814;
                9582: note <= (-2531);
                9583: note <= (-7815);
                9584: note <= (-11910);
                9585: note <= (-13985);
                9586: note <= (-13722);
                9587: note <= (-11395);
                9588: note <= (-7791);
                9589: note <= (-3995);
                9590: note <= (-1098);
                9591: note <= 101;
                9592: note <= (-697);
                9593: note <= (-3203);
                9594: note <= (-6627);
                9595: note <= (-9889);
                9596: note <= (-11910);
                9597: note <= (-11911);
                9598: note <= (-9626);
                9599: note <= (-5378);
                9600: note <= 0;
                9601: note <= 5378;
                9602: note <= 9626;
                9603: note <= 11911;
                9604: note <= 11910;
                9605: note <= 9889;
                9606: note <= 6627;
                9607: note <= 3203;
                9608: note <= 697;
                9609: note <= (-101);
                9610: note <= 1098;
                9611: note <= 3995;
                9612: note <= 7791;
                9613: note <= 11395;
                9614: note <= 13722;
                9615: note <= 13985;
                9616: note <= 11910;
                9617: note <= 7815;
                9618: note <= 2531;
                9619: note <= (-2814);
                9620: note <= (-7094);
                9621: note <= (-9474);
                9622: note <= (-9626);
                9623: note <= (-7815);
                9624: note <= (-4815);
                9625: note <= (-1697);
                9626: note <= 467;
                9627: note <= 893;
                9628: note <= (-697);
                9629: note <= (-3995);
                9630: note <= (-8192);
                9631: note <= (-12187);
                9632: note <= (-14886);
                9633: note <= (-15491);
                9634: note <= (-13722);
                9635: note <= (-9889);
                9636: note <= (-4815);
                9637: note <= 377;
                9638: note <= 4563;
                9639: note <= 6910;
                9640: note <= 7094;
                9641: note <= 5378;
                9642: note <= 2531;
                9643: note <= (-377);
                9644: note <= (-2279);
                9645: note <= (-2399);
                9646: note <= (-467);
                9647: note <= 3203;
                9648: note <= 7791;
                9649: note <= 12187;
                9650: note <= 15286;
                9651: note <= 16283;
                9652: note <= 14886;
                9653: note <= 11395;
                9654: note <= 6627;
                9655: note <= 1697;
                9656: note <= (-2279);
                9657: note <= (-4473);
                9658: note <= (-4563);
                9659: note <= (-2814);
                9660: note <= 0;
                9661: note <= 2814;
                9662: note <= 4563;
                9663: note <= 4473;
                9664: note <= 2279;
                9665: note <= (-1697);
                9666: note <= (-6627);
                9667: note <= (-11395);
                9668: note <= (-14886);
                9669: note <= (-16283);
                9670: note <= (-15286);
                9671: note <= (-12187);
                9672: note <= (-7791);
                9673: note <= (-3203);
                9674: note <= 467;
                9675: note <= 2399;
                9676: note <= 2279;
                9677: note <= 377;
                9678: note <= (-2531);
                9679: note <= (-5378);
                9680: note <= (-7094);
                9681: note <= (-6910);
                9682: note <= (-4563);
                9683: note <= (-377);
                9684: note <= 4815;
                9685: note <= 9889;
                9686: note <= 13722;
                9687: note <= 15491;
                9688: note <= 14886;
                9689: note <= 12187;
                9690: note <= 8192;
                9691: note <= 3995;
                9692: note <= 697;
                9693: note <= (-893);
                9694: note <= (-467);
                9695: note <= 1697;
                9696: note <= 4815;
                9697: note <= 7815;
                9698: note <= 9626;
                9699: note <= 9474;
                9700: note <= 7094;
                9701: note <= 2814;
                9702: note <= (-2531);
                9703: note <= (-7815);
                9704: note <= (-11910);
                9705: note <= (-13985);
                9706: note <= (-13722);
                9707: note <= (-11395);
                9708: note <= (-7791);
                9709: note <= (-3995);
                9710: note <= (-1098);
                9711: note <= 101;
                9712: note <= (-697);
                9713: note <= (-3203);
                9714: note <= (-6627);
                9715: note <= (-9889);
                9716: note <= (-11910);
                9717: note <= (-11911);
                9718: note <= (-9626);
                9719: note <= (-5378);
                9720: note <= 0;
                9721: note <= 5378;
                9722: note <= 9626;
                9723: note <= 11911;
                9724: note <= 11910;
                9725: note <= 9889;
                9726: note <= 6627;
                9727: note <= 3203;
                9728: note <= 697;
                9729: note <= (-101);
                9730: note <= 1098;
                9731: note <= 3995;
                9732: note <= 7791;
                9733: note <= 11395;
                9734: note <= 13722;
                9735: note <= 13985;
                9736: note <= 11910;
                9737: note <= 7815;
                9738: note <= 2531;
                9739: note <= (-2814);
                9740: note <= (-7094);
                9741: note <= (-9474);
                9742: note <= (-9626);
                9743: note <= (-7815);
                9744: note <= (-4815);
                9745: note <= (-1697);
                9746: note <= 467;
                9747: note <= 893;
                9748: note <= (-697);
                9749: note <= (-3995);
                9750: note <= (-8192);
                9751: note <= (-12187);
                9752: note <= (-14886);
                9753: note <= (-15491);
                9754: note <= (-13722);
                9755: note <= (-9889);
                9756: note <= (-4815);
                9757: note <= 377;
                9758: note <= 4563;
                9759: note <= 6910;
                9760: note <= 7094;
                9761: note <= 5378;
                9762: note <= 2531;
                9763: note <= (-377);
                9764: note <= (-2279);
                9765: note <= (-2399);
                9766: note <= (-467);
                9767: note <= 3203;
                9768: note <= 7791;
                9769: note <= 12187;
                9770: note <= 15286;
                9771: note <= 16283;
                9772: note <= 14886;
                9773: note <= 11395;
                9774: note <= 6627;
                9775: note <= 1697;
                9776: note <= (-2279);
                9777: note <= (-4473);
                9778: note <= (-4563);
                9779: note <= (-2814);
                9780: note <= 0;
                9781: note <= 2814;
                9782: note <= 4563;
                9783: note <= 4473;
                9784: note <= 2279;
                9785: note <= (-1697);
                9786: note <= (-6627);
                9787: note <= (-11395);
                9788: note <= (-14886);
                9789: note <= (-16283);
                9790: note <= (-15286);
                9791: note <= (-12187);
                9792: note <= (-7791);
                9793: note <= (-3203);
                9794: note <= 467;
                9795: note <= 2399;
                9796: note <= 2279;
                9797: note <= 377;
                9798: note <= (-2531);
                9799: note <= (-5378);
                9800: note <= (-7094);
                9801: note <= (-6910);
                9802: note <= (-4563);
                9803: note <= (-377);
                9804: note <= 4815;
                9805: note <= 9889;
                9806: note <= 13722;
                9807: note <= 15491;
                9808: note <= 14886;
                9809: note <= 12187;
                9810: note <= 8192;
                9811: note <= 3995;
                9812: note <= 697;
                9813: note <= (-893);
                9814: note <= (-467);
                9815: note <= 1697;
                9816: note <= 4815;
                9817: note <= 7815;
                9818: note <= 9626;
                9819: note <= 9474;
                9820: note <= 7094;
                9821: note <= 2814;
                9822: note <= (-2531);
                9823: note <= (-7815);
                9824: note <= (-11910);
                9825: note <= (-13985);
                9826: note <= (-13722);
                9827: note <= (-11395);
                9828: note <= (-7791);
                9829: note <= (-3995);
                9830: note <= (-1098);
                9831: note <= 101;
                9832: note <= (-697);
                9833: note <= (-3203);
                9834: note <= (-6627);
                9835: note <= (-9889);
                9836: note <= (-11910);
                9837: note <= (-11911);
                9838: note <= (-9626);
                9839: note <= (-5378);
                9840: note <= 0;
                9841: note <= 5378;
                9842: note <= 9626;
                9843: note <= 11911;
                9844: note <= 11910;
                9845: note <= 9889;
                9846: note <= 6627;
                9847: note <= 3203;
                9848: note <= 697;
                9849: note <= (-101);
                9850: note <= 1098;
                9851: note <= 3995;
                9852: note <= 7791;
                9853: note <= 11395;
                9854: note <= 13722;
                9855: note <= 13985;
                9856: note <= 11910;
                9857: note <= 7815;
                9858: note <= 2531;
                9859: note <= (-2814);
                9860: note <= (-7094);
                9861: note <= (-9474);
                9862: note <= (-9626);
                9863: note <= (-7815);
                9864: note <= (-4815);
                9865: note <= (-1697);
                9866: note <= 467;
                9867: note <= 893;
                9868: note <= (-697);
                9869: note <= (-3995);
                9870: note <= (-8192);
                9871: note <= (-12187);
                9872: note <= (-14886);
                9873: note <= (-15491);
                9874: note <= (-13722);
                9875: note <= (-9889);
                9876: note <= (-4815);
                9877: note <= 377;
                9878: note <= 4563;
                9879: note <= 6910;
                9880: note <= 7094;
                9881: note <= 5378;
                9882: note <= 2531;
                9883: note <= (-377);
                9884: note <= (-2279);
                9885: note <= (-2399);
                9886: note <= (-467);
                9887: note <= 3203;
                9888: note <= 7791;
                9889: note <= 12187;
                9890: note <= 15286;
                9891: note <= 16283;
                9892: note <= 14886;
                9893: note <= 11395;
                9894: note <= 6627;
                9895: note <= 1697;
                9896: note <= (-2279);
                9897: note <= (-4473);
                9898: note <= (-4563);
                9899: note <= (-2814);
                9900: note <= 0;
                9901: note <= 2814;
                9902: note <= 4563;
                9903: note <= 4473;
                9904: note <= 2279;
                9905: note <= (-1697);
                9906: note <= (-6627);
                9907: note <= (-11395);
                9908: note <= (-14886);
                9909: note <= (-16283);
                9910: note <= (-15286);
                9911: note <= (-12187);
                9912: note <= (-7791);
                9913: note <= (-3203);
                9914: note <= 467;
                9915: note <= 2399;
                9916: note <= 2279;
                9917: note <= 377;
                9918: note <= (-2531);
                9919: note <= (-5378);
                9920: note <= (-7094);
                9921: note <= (-6910);
                9922: note <= (-4563);
                9923: note <= (-377);
                9924: note <= 4815;
                9925: note <= 9889;
                9926: note <= 13722;
                9927: note <= 15491;
                9928: note <= 14886;
                9929: note <= 12187;
                9930: note <= 8192;
                9931: note <= 3995;
                9932: note <= 697;
                9933: note <= (-893);
                9934: note <= (-467);
                9935: note <= 1697;
                9936: note <= 4815;
                9937: note <= 7815;
                9938: note <= 9626;
                9939: note <= 9474;
                9940: note <= 7094;
                9941: note <= 2814;
                9942: note <= (-2531);
                9943: note <= (-7815);
                9944: note <= (-11910);
                9945: note <= (-13985);
                9946: note <= (-13722);
                9947: note <= (-11395);
                9948: note <= (-7791);
                9949: note <= (-3995);
                9950: note <= (-1098);
                9951: note <= 101;
                9952: note <= (-697);
                9953: note <= (-3203);
                9954: note <= (-6627);
                9955: note <= (-9889);
                9956: note <= (-11910);
                9957: note <= (-11911);
                9958: note <= (-9626);
                9959: note <= (-5378);
                9960: note <= 0;
                9961: note <= 5378;
                9962: note <= 9626;
                9963: note <= 11911;
                9964: note <= 11910;
                9965: note <= 9889;
                9966: note <= 6627;
                9967: note <= 3203;
                9968: note <= 697;
                9969: note <= (-101);
                9970: note <= 1098;
                9971: note <= 3995;
                9972: note <= 7791;
                9973: note <= 11395;
                9974: note <= 13722;
                9975: note <= 13985;
                9976: note <= 11910;
                9977: note <= 7815;
                9978: note <= 2531;
                9979: note <= (-2814);
                9980: note <= (-7094);
                9981: note <= (-9474);
                9982: note <= (-9626);
                9983: note <= (-7815);
                9984: note <= (-4815);
                9985: note <= (-1697);
                9986: note <= 467;
                9987: note <= 893;
                9988: note <= (-697);
                9989: note <= (-3995);
                9990: note <= (-8192);
                9991: note <= (-12187);
                9992: note <= (-14886);
                9993: note <= (-15491);
                9994: note <= (-13722);
                9995: note <= (-9889);
                9996: note <= (-4815);
                9997: note <= 377;
                9998: note <= 4563;
                9999: note <= 6910;
                10000: note <= 7094;
                10001: note <= 5378;
                10002: note <= 2531;
                10003: note <= (-377);
                10004: note <= (-2279);
                10005: note <= (-2399);
                10006: note <= (-467);
                10007: note <= 3203;
                10008: note <= 7791;
                10009: note <= 12187;
                10010: note <= 15286;
                10011: note <= 16283;
                10012: note <= 14886;
                10013: note <= 11395;
                10014: note <= 6627;
                10015: note <= 1697;
                10016: note <= (-2279);
                10017: note <= (-4473);
                10018: note <= (-4563);
                10019: note <= (-2814);
                10020: note <= 0;
                10021: note <= 2814;
                10022: note <= 4563;
                10023: note <= 4473;
                10024: note <= 2279;
                10025: note <= (-1697);
                10026: note <= (-6627);
                10027: note <= (-11395);
                10028: note <= (-14886);
                10029: note <= (-16283);
                10030: note <= (-15286);
                10031: note <= (-12187);
                10032: note <= (-7791);
                10033: note <= (-3203);
                10034: note <= 467;
                10035: note <= 2399;
                10036: note <= 2279;
                10037: note <= 377;
                10038: note <= (-2531);
                10039: note <= (-5378);
                10040: note <= (-7094);
                10041: note <= (-6910);
                10042: note <= (-4563);
                10043: note <= (-377);
                10044: note <= 4815;
                10045: note <= 9889;
                10046: note <= 13722;
                10047: note <= 15491;
                10048: note <= 14886;
                10049: note <= 12187;
                10050: note <= 8192;
                10051: note <= 3995;
                10052: note <= 697;
                10053: note <= (-893);
                10054: note <= (-467);
                10055: note <= 1697;
                10056: note <= 4815;
                10057: note <= 7815;
                10058: note <= 9626;
                10059: note <= 9474;
                10060: note <= 7094;
                10061: note <= 2814;
                10062: note <= (-2531);
                10063: note <= (-7815);
                10064: note <= (-11910);
                10065: note <= (-13985);
                10066: note <= (-13722);
                10067: note <= (-11395);
                10068: note <= (-7791);
                10069: note <= (-3995);
                10070: note <= (-1098);
                10071: note <= 101;
                10072: note <= (-697);
                10073: note <= (-3203);
                10074: note <= (-6627);
                10075: note <= (-9889);
                10076: note <= (-11910);
                10077: note <= (-11911);
                10078: note <= (-9626);
                10079: note <= (-5378);
                10080: note <= 0;
                10081: note <= 5378;
                10082: note <= 9626;
                10083: note <= 11911;
                10084: note <= 11910;
                10085: note <= 9889;
                10086: note <= 6627;
                10087: note <= 3203;
                10088: note <= 697;
                10089: note <= (-101);
                10090: note <= 1098;
                10091: note <= 3995;
                10092: note <= 7791;
                10093: note <= 11395;
                10094: note <= 13722;
                10095: note <= 13985;
                10096: note <= 11910;
                10097: note <= 7815;
                10098: note <= 2531;
                10099: note <= (-2814);
                10100: note <= (-7094);
                10101: note <= (-9474);
                10102: note <= (-9626);
                10103: note <= (-7815);
                10104: note <= (-4815);
                10105: note <= (-1697);
                10106: note <= 467;
                10107: note <= 893;
                10108: note <= (-697);
                10109: note <= (-3995);
                10110: note <= (-8192);
                10111: note <= (-12187);
                10112: note <= (-14886);
                10113: note <= (-15491);
                10114: note <= (-13722);
                10115: note <= (-9889);
                10116: note <= (-4815);
                10117: note <= 377;
                10118: note <= 4563;
                10119: note <= 6910;
                10120: note <= 7094;
                10121: note <= 5378;
                10122: note <= 2531;
                10123: note <= (-377);
                10124: note <= (-2279);
                10125: note <= (-2399);
                10126: note <= (-467);
                10127: note <= 3203;
                10128: note <= 7791;
                10129: note <= 12187;
                10130: note <= 15286;
                10131: note <= 16283;
                10132: note <= 14886;
                10133: note <= 11395;
                10134: note <= 6627;
                10135: note <= 1697;
                10136: note <= (-2279);
                10137: note <= (-4473);
                10138: note <= (-4563);
                10139: note <= (-2814);
                10140: note <= 0;
                10141: note <= 2814;
                10142: note <= 4563;
                10143: note <= 4473;
                10144: note <= 2279;
                10145: note <= (-1697);
                10146: note <= (-6627);
                10147: note <= (-11395);
                10148: note <= (-14886);
                10149: note <= (-16283);
                10150: note <= (-15286);
                10151: note <= (-12187);
                10152: note <= (-7791);
                10153: note <= (-3203);
                10154: note <= 467;
                10155: note <= 2399;
                10156: note <= 2279;
                10157: note <= 377;
                10158: note <= (-2531);
                10159: note <= (-5378);
                10160: note <= (-7094);
                10161: note <= (-6910);
                10162: note <= (-4563);
                10163: note <= (-377);
                10164: note <= 4815;
                10165: note <= 9889;
                10166: note <= 13722;
                10167: note <= 15491;
                10168: note <= 14886;
                10169: note <= 12187;
                10170: note <= 8192;
                10171: note <= 3995;
                10172: note <= 697;
                10173: note <= (-893);
                10174: note <= (-467);
                10175: note <= 1697;
                10176: note <= 4815;
                10177: note <= 7815;
                10178: note <= 9626;
                10179: note <= 9474;
                10180: note <= 7094;
                10181: note <= 2814;
                10182: note <= (-2531);
                10183: note <= (-7815);
                10184: note <= (-11910);
                10185: note <= (-13985);
                10186: note <= (-13722);
                10187: note <= (-11395);
                10188: note <= (-7791);
                10189: note <= (-3995);
                10190: note <= (-1098);
                10191: note <= 101;
                10192: note <= (-697);
                10193: note <= (-3203);
                10194: note <= (-6627);
                10195: note <= (-9889);
                10196: note <= (-11910);
                10197: note <= (-11911);
                10198: note <= (-9626);
                10199: note <= (-5378);
                10200: note <= 0;
                10201: note <= 5378;
                10202: note <= 9626;
                10203: note <= 11911;
                10204: note <= 11910;
                10205: note <= 9889;
                10206: note <= 6627;
                10207: note <= 3203;
                10208: note <= 697;
                10209: note <= (-101);
                10210: note <= 1098;
                10211: note <= 3995;
                10212: note <= 7791;
                10213: note <= 11395;
                10214: note <= 13722;
                10215: note <= 13985;
                10216: note <= 11910;
                10217: note <= 7815;
                10218: note <= 2531;
                10219: note <= (-2814);
                10220: note <= (-7094);
                10221: note <= (-9474);
                10222: note <= (-9626);
                10223: note <= (-7815);
                10224: note <= (-4815);
                10225: note <= (-1697);
                10226: note <= 467;
                10227: note <= 893;
                10228: note <= (-697);
                10229: note <= (-3995);
                10230: note <= (-8192);
                10231: note <= (-12187);
                10232: note <= (-14886);
                10233: note <= (-15491);
                10234: note <= (-13722);
                10235: note <= (-9889);
                10236: note <= (-4815);
                10237: note <= 377;
                10238: note <= 4563;
                10239: note <= 6910;
                10240: note <= 7094;
                10241: note <= 5378;
                10242: note <= 2531;
                10243: note <= (-377);
                10244: note <= (-2279);
                10245: note <= (-2399);
                10246: note <= (-467);
                10247: note <= 3203;
                10248: note <= 7791;
                10249: note <= 12187;
                10250: note <= 15286;
                10251: note <= 16283;
                10252: note <= 14886;
                10253: note <= 11395;
                10254: note <= 6627;
                10255: note <= 1697;
                10256: note <= (-2279);
                10257: note <= (-4473);
                10258: note <= (-4563);
                10259: note <= (-2814);
                10260: note <= 0;
                10261: note <= 2814;
                10262: note <= 4563;
                10263: note <= 4473;
                10264: note <= 2279;
                10265: note <= (-1697);
                10266: note <= (-6627);
                10267: note <= (-11395);
                10268: note <= (-14886);
                10269: note <= (-16283);
                10270: note <= (-15286);
                10271: note <= (-12187);
                10272: note <= (-7791);
                10273: note <= (-3203);
                10274: note <= 467;
                10275: note <= 2399;
                10276: note <= 2279;
                10277: note <= 377;
                10278: note <= (-2531);
                10279: note <= (-5378);
                10280: note <= (-7094);
                10281: note <= (-6910);
                10282: note <= (-4563);
                10283: note <= (-377);
                10284: note <= 4815;
                10285: note <= 9889;
                10286: note <= 13722;
                10287: note <= 15491;
                10288: note <= 14886;
                10289: note <= 12187;
                10290: note <= 8192;
                10291: note <= 3995;
                10292: note <= 697;
                10293: note <= (-893);
                10294: note <= (-467);
                10295: note <= 1697;
                10296: note <= 4815;
                10297: note <= 7815;
                10298: note <= 9626;
                10299: note <= 9474;
                10300: note <= 7094;
                10301: note <= 2814;
                10302: note <= (-2531);
                10303: note <= (-7815);
                10304: note <= (-11910);
                10305: note <= (-13985);
                10306: note <= (-13722);
                10307: note <= (-11395);
                10308: note <= (-7791);
                10309: note <= (-3995);
                10310: note <= (-1098);
                10311: note <= 101;
                10312: note <= (-697);
                10313: note <= (-3203);
                10314: note <= (-6627);
                10315: note <= (-9889);
                10316: note <= (-11910);
                10317: note <= (-11911);
                10318: note <= (-9626);
                10319: note <= (-5378);
                10320: note <= 0;
                10321: note <= 5378;
                10322: note <= 9626;
                10323: note <= 11911;
                10324: note <= 11910;
                10325: note <= 9889;
                10326: note <= 6627;
                10327: note <= 3203;
                10328: note <= 697;
                10329: note <= (-101);
                10330: note <= 1098;
                10331: note <= 3995;
                10332: note <= 7791;
                10333: note <= 11395;
                10334: note <= 13722;
                10335: note <= 13985;
                10336: note <= 11910;
                10337: note <= 7815;
                10338: note <= 2531;
                10339: note <= (-2814);
                10340: note <= (-7094);
                10341: note <= (-9474);
                10342: note <= (-9626);
                10343: note <= (-7815);
                10344: note <= (-4815);
                10345: note <= (-1697);
                10346: note <= 467;
                10347: note <= 893;
                10348: note <= (-697);
                10349: note <= (-3995);
                10350: note <= (-8192);
                10351: note <= (-12187);
                10352: note <= (-14886);
                10353: note <= (-15491);
                10354: note <= (-13722);
                10355: note <= (-9889);
                10356: note <= (-4815);
                10357: note <= 377;
                10358: note <= 4563;
                10359: note <= 6910;
                10360: note <= 7094;
                10361: note <= 5378;
                10362: note <= 2531;
                10363: note <= (-377);
                10364: note <= (-2279);
                10365: note <= (-2399);
                10366: note <= (-467);
                10367: note <= 3203;
                10368: note <= 7791;
                10369: note <= 12187;
                10370: note <= 15286;
                10371: note <= 16283;
                10372: note <= 14886;
                10373: note <= 11395;
                10374: note <= 6627;
                10375: note <= 1697;
                10376: note <= (-2279);
                10377: note <= (-4473);
                10378: note <= (-4563);
                10379: note <= (-2814);
                10380: note <= 0;
                10381: note <= 2814;
                10382: note <= 4563;
                10383: note <= 4473;
                10384: note <= 2279;
                10385: note <= (-1697);
                10386: note <= (-6627);
                10387: note <= (-11395);
                10388: note <= (-14886);
                10389: note <= (-16283);
                10390: note <= (-15286);
                10391: note <= (-12187);
                10392: note <= (-7791);
                10393: note <= (-3203);
                10394: note <= 467;
                10395: note <= 2399;
                10396: note <= 2279;
                10397: note <= 377;
                10398: note <= (-2531);
                10399: note <= (-5378);
                10400: note <= (-7094);
                10401: note <= (-6910);
                10402: note <= (-4563);
                10403: note <= (-377);
                10404: note <= 4815;
                10405: note <= 9889;
                10406: note <= 13722;
                10407: note <= 15491;
                10408: note <= 14886;
                10409: note <= 12187;
                10410: note <= 8192;
                10411: note <= 3995;
                10412: note <= 697;
                10413: note <= (-893);
                10414: note <= (-467);
                10415: note <= 1697;
                10416: note <= 4815;
                10417: note <= 7815;
                10418: note <= 9626;
                10419: note <= 9474;
                10420: note <= 7094;
                10421: note <= 2814;
                10422: note <= (-2531);
                10423: note <= (-7815);
                10424: note <= (-11910);
                10425: note <= (-13985);
                10426: note <= (-13722);
                10427: note <= (-11395);
                10428: note <= (-7791);
                10429: note <= (-3995);
                10430: note <= (-1098);
                10431: note <= 101;
                10432: note <= (-697);
                10433: note <= (-3203);
                10434: note <= (-6627);
                10435: note <= (-9889);
                10436: note <= (-11910);
                10437: note <= (-11911);
                10438: note <= (-9626);
                10439: note <= (-5378);
                10440: note <= 0;
                10441: note <= 5378;
                10442: note <= 9626;
                10443: note <= 11911;
                10444: note <= 11910;
                10445: note <= 9889;
                10446: note <= 6627;
                10447: note <= 3203;
                10448: note <= 697;
                10449: note <= (-101);
                10450: note <= 1098;
                10451: note <= 3995;
                10452: note <= 7791;
                10453: note <= 11395;
                10454: note <= 13722;
                10455: note <= 13985;
                10456: note <= 11910;
                10457: note <= 7815;
                10458: note <= 2531;
                10459: note <= (-2814);
                10460: note <= (-7094);
                10461: note <= (-9474);
                10462: note <= (-9626);
                10463: note <= (-7815);
                10464: note <= (-4815);
                10465: note <= (-1697);
                10466: note <= 467;
                10467: note <= 893;
                10468: note <= (-697);
                10469: note <= (-3995);
                10470: note <= (-8192);
                10471: note <= (-12187);
                10472: note <= (-14886);
                10473: note <= (-15491);
                10474: note <= (-13722);
                10475: note <= (-9889);
                10476: note <= (-4815);
                10477: note <= 377;
                10478: note <= 4563;
                10479: note <= 6910;
                10480: note <= 7094;
                10481: note <= 5378;
                10482: note <= 2531;
                10483: note <= (-377);
                10484: note <= (-2279);
                10485: note <= (-2399);
                10486: note <= (-467);
                10487: note <= 3203;
                10488: note <= 7791;
                10489: note <= 12187;
                10490: note <= 15286;
                10491: note <= 16283;
                10492: note <= 14886;
                10493: note <= 11395;
                10494: note <= 6627;
                10495: note <= 1697;
                10496: note <= (-2279);
                10497: note <= (-4473);
                10498: note <= (-4563);
                10499: note <= (-2814);
                10500: note <= 0;
                10501: note <= 2814;
                10502: note <= 4563;
                10503: note <= 4473;
                10504: note <= 2279;
                10505: note <= (-1697);
                10506: note <= (-6627);
                10507: note <= (-11395);
                10508: note <= (-14886);
                10509: note <= (-16283);
                10510: note <= (-15286);
                10511: note <= (-12187);
                10512: note <= (-7791);
                10513: note <= (-3203);
                10514: note <= 467;
                10515: note <= 2399;
                10516: note <= 2279;
                10517: note <= 377;
                10518: note <= (-2531);
                10519: note <= (-5378);
                10520: note <= (-7094);
                10521: note <= (-6910);
                10522: note <= (-4563);
                10523: note <= (-377);
                10524: note <= 4815;
                10525: note <= 9889;
                10526: note <= 13722;
                10527: note <= 15491;
                10528: note <= 14886;
                10529: note <= 12187;
                10530: note <= 8192;
                10531: note <= 3995;
                10532: note <= 697;
                10533: note <= (-893);
                10534: note <= (-467);
                10535: note <= 1697;
                10536: note <= 4815;
                10537: note <= 7815;
                10538: note <= 9626;
                10539: note <= 9474;
                10540: note <= 7094;
                10541: note <= 2814;
                10542: note <= (-2531);
                10543: note <= (-7815);
                10544: note <= (-11910);
                10545: note <= (-13985);
                10546: note <= (-13722);
                10547: note <= (-11395);
                10548: note <= (-7791);
                10549: note <= (-3995);
                10550: note <= (-1098);
                10551: note <= 101;
                10552: note <= (-697);
                10553: note <= (-3203);
                10554: note <= (-6627);
                10555: note <= (-9889);
                10556: note <= (-11910);
                10557: note <= (-11911);
                10558: note <= (-9626);
                10559: note <= (-5378);
                10560: note <= 0;
                10561: note <= 5378;
                10562: note <= 9626;
                10563: note <= 11911;
                10564: note <= 11910;
                10565: note <= 9889;
                10566: note <= 6627;
                10567: note <= 3203;
                10568: note <= 697;
                10569: note <= (-101);
                10570: note <= 1098;
                10571: note <= 3995;
                10572: note <= 7791;
                10573: note <= 11395;
                10574: note <= 13722;
                10575: note <= 13985;
                10576: note <= 11910;
                10577: note <= 7815;
                10578: note <= 2531;
                10579: note <= (-2814);
                10580: note <= (-7094);
                10581: note <= (-9474);
                10582: note <= (-9626);
                10583: note <= (-7815);
                10584: note <= (-4815);
                10585: note <= (-1697);
                10586: note <= 467;
                10587: note <= 893;
                10588: note <= (-697);
                10589: note <= (-3995);
                10590: note <= (-8192);
                10591: note <= (-12187);
                10592: note <= (-14886);
                10593: note <= (-15491);
                10594: note <= (-13722);
                10595: note <= (-9889);
                10596: note <= (-4815);
                10597: note <= 377;
                10598: note <= 4563;
                10599: note <= 6910;
                10600: note <= 7094;
                10601: note <= 5378;
                10602: note <= 2531;
                10603: note <= (-377);
                10604: note <= (-2279);
                10605: note <= (-2399);
                10606: note <= (-467);
                10607: note <= 3203;
                10608: note <= 7791;
                10609: note <= 12187;
                10610: note <= 15286;
                10611: note <= 16283;
                10612: note <= 14886;
                10613: note <= 11395;
                10614: note <= 6627;
                10615: note <= 1697;
                10616: note <= (-2279);
                10617: note <= (-4473);
                10618: note <= (-4563);
                10619: note <= (-2814);
                10620: note <= 0;
                10621: note <= 2814;
                10622: note <= 4563;
                10623: note <= 4473;
                10624: note <= 2279;
                10625: note <= (-1697);
                10626: note <= (-6627);
                10627: note <= (-11395);
                10628: note <= (-14886);
                10629: note <= (-16283);
                10630: note <= (-15286);
                10631: note <= (-12187);
                10632: note <= (-7791);
                10633: note <= (-3203);
                10634: note <= 467;
                10635: note <= 2399;
                10636: note <= 2279;
                10637: note <= 377;
                10638: note <= (-2531);
                10639: note <= (-5378);
                10640: note <= (-7094);
                10641: note <= (-6910);
                10642: note <= (-4563);
                10643: note <= (-377);
                10644: note <= 4815;
                10645: note <= 9889;
                10646: note <= 13722;
                10647: note <= 15491;
                10648: note <= 14886;
                10649: note <= 12187;
                10650: note <= 8192;
                10651: note <= 3995;
                10652: note <= 697;
                10653: note <= (-893);
                10654: note <= (-467);
                10655: note <= 1697;
                10656: note <= 4815;
                10657: note <= 7815;
                10658: note <= 9626;
                10659: note <= 9474;
                10660: note <= 7094;
                10661: note <= 2814;
                10662: note <= (-2531);
                10663: note <= (-7815);
                10664: note <= (-11910);
                10665: note <= (-13985);
                10666: note <= (-13722);
                10667: note <= (-11395);
                10668: note <= (-7791);
                10669: note <= (-3995);
                10670: note <= (-1098);
                10671: note <= 101;
                10672: note <= (-697);
                10673: note <= (-3203);
                10674: note <= (-6627);
                10675: note <= (-9889);
                10676: note <= (-11910);
                10677: note <= (-11911);
                10678: note <= (-9626);
                10679: note <= (-5378);
                10680: note <= 0;
                10681: note <= 5378;
                10682: note <= 9626;
                10683: note <= 11911;
                10684: note <= 11910;
                10685: note <= 9889;
                10686: note <= 6627;
                10687: note <= 3203;
                10688: note <= 697;
                10689: note <= (-101);
                10690: note <= 1098;
                10691: note <= 3995;
                10692: note <= 7791;
                10693: note <= 11395;
                10694: note <= 13722;
                10695: note <= 13985;
                10696: note <= 11910;
                10697: note <= 7815;
                10698: note <= 2531;
                10699: note <= (-2814);
                10700: note <= (-7094);
                10701: note <= (-9474);
                10702: note <= (-9626);
                10703: note <= (-7815);
                10704: note <= (-4815);
                10705: note <= (-1697);
                10706: note <= 467;
                10707: note <= 893;
                10708: note <= (-697);
                10709: note <= (-3995);
                10710: note <= (-8192);
                10711: note <= (-12187);
                10712: note <= (-14886);
                10713: note <= (-15491);
                10714: note <= (-13722);
                10715: note <= (-9889);
                10716: note <= (-4815);
                10717: note <= 377;
                10718: note <= 4563;
                10719: note <= 6910;
                10720: note <= 7094;
                10721: note <= 5378;
                10722: note <= 2531;
                10723: note <= (-377);
                10724: note <= (-2279);
                10725: note <= (-2399);
                10726: note <= (-467);
                10727: note <= 3203;
                10728: note <= 7791;
                10729: note <= 12187;
                10730: note <= 15286;
                10731: note <= 16283;
                10732: note <= 14886;
                10733: note <= 11395;
                10734: note <= 6627;
                10735: note <= 1697;
                10736: note <= (-2279);
                10737: note <= (-4473);
                10738: note <= (-4563);
                10739: note <= (-2814);
                10740: note <= 0;
                10741: note <= 2814;
                10742: note <= 4563;
                10743: note <= 4473;
                10744: note <= 2279;
                10745: note <= (-1697);
                10746: note <= (-6627);
                10747: note <= (-11395);
                10748: note <= (-14886);
                10749: note <= (-16283);
                10750: note <= (-15286);
                10751: note <= (-12187);
                10752: note <= (-7791);
                10753: note <= (-3203);
                10754: note <= 467;
                10755: note <= 2399;
                10756: note <= 2279;
                10757: note <= 377;
                10758: note <= (-2531);
                10759: note <= (-5378);
                10760: note <= (-7094);
                10761: note <= (-6910);
                10762: note <= (-4563);
                10763: note <= (-377);
                10764: note <= 4815;
                10765: note <= 9889;
                10766: note <= 13722;
                10767: note <= 15491;
                10768: note <= 14886;
                10769: note <= 12187;
                10770: note <= 8192;
                10771: note <= 3995;
                10772: note <= 697;
                10773: note <= (-893);
                10774: note <= (-467);
                10775: note <= 1697;
                10776: note <= 4815;
                10777: note <= 7815;
                10778: note <= 9626;
                10779: note <= 9474;
                10780: note <= 7094;
                10781: note <= 2814;
                10782: note <= (-2531);
                10783: note <= (-7815);
                10784: note <= (-11910);
                10785: note <= (-13985);
                10786: note <= (-13722);
                10787: note <= (-11395);
                10788: note <= (-7791);
                10789: note <= (-3995);
                10790: note <= (-1098);
                10791: note <= 101;
                10792: note <= (-697);
                10793: note <= (-3203);
                10794: note <= (-6627);
                10795: note <= (-9889);
                10796: note <= (-11910);
                10797: note <= (-11911);
                10798: note <= (-9626);
                10799: note <= (-5378);
                10800: note <= 0;
                10801: note <= 5378;
                10802: note <= 9626;
                10803: note <= 11911;
                10804: note <= 11910;
                10805: note <= 9889;
                10806: note <= 6627;
                10807: note <= 3203;
                10808: note <= 697;
                10809: note <= (-101);
                10810: note <= 1098;
                10811: note <= 3995;
                10812: note <= 7791;
                10813: note <= 11395;
                10814: note <= 13722;
                10815: note <= 13985;
                10816: note <= 11910;
                10817: note <= 7815;
                10818: note <= 2531;
                10819: note <= (-2814);
                10820: note <= (-7094);
                10821: note <= (-9474);
                10822: note <= (-9626);
                10823: note <= (-7815);
                10824: note <= (-4815);
                10825: note <= (-1697);
                10826: note <= 467;
                10827: note <= 893;
                10828: note <= (-697);
                10829: note <= (-3995);
                10830: note <= (-8192);
                10831: note <= (-12187);
                10832: note <= (-14886);
                10833: note <= (-15491);
                10834: note <= (-13722);
                10835: note <= (-9889);
                10836: note <= (-4815);
                10837: note <= 377;
                10838: note <= 4563;
                10839: note <= 6910;
                10840: note <= 7094;
                10841: note <= 5378;
                10842: note <= 2531;
                10843: note <= (-377);
                10844: note <= (-2279);
                10845: note <= (-2399);
                10846: note <= (-467);
                10847: note <= 3203;
                10848: note <= 7791;
                10849: note <= 12187;
                10850: note <= 15286;
                10851: note <= 16283;
                10852: note <= 14886;
                10853: note <= 11395;
                10854: note <= 6627;
                10855: note <= 1697;
                10856: note <= (-2279);
                10857: note <= (-4473);
                10858: note <= (-4563);
                10859: note <= (-2814);
                10860: note <= 0;
                10861: note <= 2814;
                10862: note <= 4563;
                10863: note <= 4473;
                10864: note <= 2279;
                10865: note <= (-1697);
                10866: note <= (-6627);
                10867: note <= (-11395);
                10868: note <= (-14886);
                10869: note <= (-16283);
                10870: note <= (-15286);
                10871: note <= (-12187);
                10872: note <= (-7791);
                10873: note <= (-3203);
                10874: note <= 467;
                10875: note <= 2399;
                10876: note <= 2279;
                10877: note <= 377;
                10878: note <= (-2531);
                10879: note <= (-5378);
                10880: note <= (-7094);
                10881: note <= (-6910);
                10882: note <= (-4563);
                10883: note <= (-377);
                10884: note <= 4815;
                10885: note <= 9889;
                10886: note <= 13722;
                10887: note <= 15491;
                10888: note <= 14886;
                10889: note <= 12187;
                10890: note <= 8192;
                10891: note <= 3995;
                10892: note <= 697;
                10893: note <= (-893);
                10894: note <= (-467);
                10895: note <= 1697;
                10896: note <= 4815;
                10897: note <= 7815;
                10898: note <= 9626;
                10899: note <= 9474;
                10900: note <= 7094;
                10901: note <= 2814;
                10902: note <= (-2531);
                10903: note <= (-7815);
                10904: note <= (-11910);
                10905: note <= (-13985);
                10906: note <= (-13722);
                10907: note <= (-11395);
                10908: note <= (-7791);
                10909: note <= (-3995);
                10910: note <= (-1098);
                10911: note <= 101;
                10912: note <= (-697);
                10913: note <= (-3203);
                10914: note <= (-6627);
                10915: note <= (-9889);
                10916: note <= (-11910);
                10917: note <= (-11911);
                10918: note <= (-9626);
                10919: note <= (-5378);
                10920: note <= 0;
                10921: note <= 5378;
                10922: note <= 9626;
                10923: note <= 11911;
                10924: note <= 11910;
                10925: note <= 9889;
                10926: note <= 6627;
                10927: note <= 3203;
                10928: note <= 697;
                10929: note <= (-101);
                10930: note <= 1098;
                10931: note <= 3995;
                10932: note <= 7791;
                10933: note <= 11395;
                10934: note <= 13722;
                10935: note <= 13985;
                10936: note <= 11910;
                10937: note <= 7815;
                10938: note <= 2531;
                10939: note <= (-2814);
                10940: note <= (-7094);
                10941: note <= (-9474);
                10942: note <= (-9626);
                10943: note <= (-7815);
                10944: note <= (-4815);
                10945: note <= (-1697);
                10946: note <= 467;
                10947: note <= 893;
                10948: note <= (-697);
                10949: note <= (-3995);
                10950: note <= (-8192);
                10951: note <= (-12187);
                10952: note <= (-14886);
                10953: note <= (-15491);
                10954: note <= (-13722);
                10955: note <= (-9889);
                10956: note <= (-4815);
                10957: note <= 377;
                10958: note <= 4563;
                10959: note <= 6910;
                10960: note <= 7094;
                10961: note <= 5378;
                10962: note <= 2531;
                10963: note <= (-377);
                10964: note <= (-2279);
                10965: note <= (-2399);
                10966: note <= (-467);
                10967: note <= 3203;
                10968: note <= 7791;
                10969: note <= 12187;
                10970: note <= 15286;
                10971: note <= 16283;
                10972: note <= 14886;
                10973: note <= 11395;
                10974: note <= 6627;
                10975: note <= 1697;
                10976: note <= (-2279);
                10977: note <= (-4473);
                10978: note <= (-4563);
                10979: note <= (-2814);
                10980: note <= 0;
                10981: note <= 2814;
                10982: note <= 4563;
                10983: note <= 4473;
                10984: note <= 2279;
                10985: note <= (-1697);
                10986: note <= (-6627);
                10987: note <= (-11395);
                10988: note <= (-14886);
                10989: note <= (-16283);
                10990: note <= (-15286);
                10991: note <= (-12187);
                10992: note <= (-7791);
                10993: note <= (-3203);
                10994: note <= 467;
                10995: note <= 2399;
                10996: note <= 2279;
                10997: note <= 377;
                10998: note <= (-2531);
                10999: note <= (-5378);
                11000: note <= (-7094);
                11001: note <= (-6910);
                11002: note <= (-4563);
                11003: note <= (-377);
                11004: note <= 4815;
                11005: note <= 9889;
                11006: note <= 13722;
                11007: note <= 15491;
                11008: note <= 14886;
                11009: note <= 12187;
                11010: note <= 8192;
                11011: note <= 3995;
                11012: note <= 697;
                11013: note <= (-893);
                11014: note <= (-467);
                11015: note <= 1697;
                11016: note <= 4815;
                11017: note <= 7815;
                11018: note <= 9626;
                11019: note <= 9474;
                11020: note <= 7094;
                11021: note <= 2814;
                11022: note <= (-2531);
                11023: note <= (-7815);
                11024: note <= (-11910);
                11025: note <= (-13985);
                11026: note <= (-13722);
                11027: note <= (-11395);
                11028: note <= (-7791);
                11029: note <= (-3995);
                11030: note <= (-1098);
                11031: note <= 101;
                11032: note <= (-697);
                11033: note <= (-3203);
                11034: note <= (-6627);
                11035: note <= (-9889);
                11036: note <= (-11910);
                11037: note <= (-11911);
                11038: note <= (-9626);
                11039: note <= (-5378);
                11040: note <= 0;
                11041: note <= 5378;
                11042: note <= 9626;
                11043: note <= 11911;
                11044: note <= 11910;
                11045: note <= 9889;
                11046: note <= 6627;
                11047: note <= 3203;
                11048: note <= 697;
                11049: note <= (-101);
                11050: note <= 1098;
                11051: note <= 3995;
                11052: note <= 7791;
                11053: note <= 11395;
                11054: note <= 13722;
                11055: note <= 13985;
                11056: note <= 11910;
                11057: note <= 7815;
                11058: note <= 2531;
                11059: note <= (-2814);
                11060: note <= (-7094);
                11061: note <= (-9474);
                11062: note <= (-9626);
                11063: note <= (-7815);
                11064: note <= (-4815);
                11065: note <= (-1697);
                11066: note <= 467;
                11067: note <= 893;
                11068: note <= (-697);
                11069: note <= (-3995);
                11070: note <= (-8192);
                11071: note <= (-12187);
                11072: note <= (-14886);
                11073: note <= (-15491);
                11074: note <= (-13722);
                11075: note <= (-9889);
                11076: note <= (-4815);
                11077: note <= 377;
                11078: note <= 4563;
                11079: note <= 6910;
                11080: note <= 7094;
                11081: note <= 5378;
                11082: note <= 2531;
                11083: note <= (-377);
                11084: note <= (-2279);
                11085: note <= (-2399);
                11086: note <= (-467);
                11087: note <= 3203;
                11088: note <= 7791;
                11089: note <= 12187;
                11090: note <= 15286;
                11091: note <= 16283;
                11092: note <= 14886;
                11093: note <= 11395;
                11094: note <= 6627;
                11095: note <= 1697;
                11096: note <= (-2279);
                11097: note <= (-4473);
                11098: note <= (-4563);
                11099: note <= (-2814);
                11100: note <= 0;
                11101: note <= 2814;
                11102: note <= 4563;
                11103: note <= 4473;
                11104: note <= 2279;
                11105: note <= (-1697);
                11106: note <= (-6627);
                11107: note <= (-11395);
                11108: note <= (-14886);
                11109: note <= (-16283);
                11110: note <= (-15286);
                11111: note <= (-12187);
                11112: note <= (-7791);
                11113: note <= (-3203);
                11114: note <= 467;
                11115: note <= 2399;
                11116: note <= 2279;
                11117: note <= 377;
                11118: note <= (-2531);
                11119: note <= (-5378);
                11120: note <= (-7094);
                11121: note <= (-6910);
                11122: note <= (-4563);
                11123: note <= (-377);
                11124: note <= 4815;
                11125: note <= 9889;
                11126: note <= 13722;
                11127: note <= 15491;
                11128: note <= 14886;
                11129: note <= 12187;
                11130: note <= 8192;
                11131: note <= 3995;
                11132: note <= 697;
                11133: note <= (-893);
                11134: note <= (-467);
                11135: note <= 1697;
                11136: note <= 4815;
                11137: note <= 7815;
                11138: note <= 9626;
                11139: note <= 9474;
                11140: note <= 7094;
                11141: note <= 2814;
                11142: note <= (-2531);
                11143: note <= (-7815);
                11144: note <= (-11910);
                11145: note <= (-13985);
                11146: note <= (-13722);
                11147: note <= (-11395);
                11148: note <= (-7791);
                11149: note <= (-3995);
                11150: note <= (-1098);
                11151: note <= 101;
                11152: note <= (-697);
                11153: note <= (-3203);
                11154: note <= (-6627);
                11155: note <= (-9889);
                11156: note <= (-11910);
                11157: note <= (-11911);
                11158: note <= (-9626);
                11159: note <= (-5378);
                11160: note <= 0;
                11161: note <= 5378;
                11162: note <= 9626;
                11163: note <= 11911;
                11164: note <= 11910;
                11165: note <= 9889;
                11166: note <= 6627;
                11167: note <= 3203;
                11168: note <= 697;
                11169: note <= (-101);
                11170: note <= 1098;
                11171: note <= 3995;
                11172: note <= 7791;
                11173: note <= 11395;
                11174: note <= 13722;
                11175: note <= 13985;
                11176: note <= 11910;
                11177: note <= 7815;
                11178: note <= 2531;
                11179: note <= (-2814);
                11180: note <= (-7094);
                11181: note <= (-9474);
                11182: note <= (-9626);
                11183: note <= (-7815);
                11184: note <= (-4815);
                11185: note <= (-1697);
                11186: note <= 467;
                11187: note <= 893;
                11188: note <= (-697);
                11189: note <= (-3995);
                11190: note <= (-8192);
                11191: note <= (-12187);
                11192: note <= (-14886);
                11193: note <= (-15491);
                11194: note <= (-13722);
                11195: note <= (-9889);
                11196: note <= (-4815);
                11197: note <= 377;
                11198: note <= 4563;
                11199: note <= 6910;
                11200: note <= 7094;
                11201: note <= 5378;
                11202: note <= 2531;
                11203: note <= (-377);
                11204: note <= (-2279);
                11205: note <= (-2399);
                11206: note <= (-467);
                11207: note <= 3203;
                11208: note <= 7791;
                11209: note <= 12187;
                11210: note <= 15286;
                11211: note <= 16283;
                11212: note <= 14886;
                11213: note <= 11395;
                11214: note <= 6627;
                11215: note <= 1697;
                11216: note <= (-2279);
                11217: note <= (-4473);
                11218: note <= (-4563);
                11219: note <= (-2814);
                11220: note <= 0;
                11221: note <= 2814;
                11222: note <= 4563;
                11223: note <= 4473;
                11224: note <= 2279;
                11225: note <= (-1697);
                11226: note <= (-6627);
                11227: note <= (-11395);
                11228: note <= (-14886);
                11229: note <= (-16283);
                11230: note <= (-15286);
                11231: note <= (-12187);
                11232: note <= (-7791);
                11233: note <= (-3203);
                11234: note <= 467;
                11235: note <= 2399;
                11236: note <= 2279;
                11237: note <= 377;
                11238: note <= (-2531);
                11239: note <= (-5378);
                11240: note <= (-7094);
                11241: note <= (-6910);
                11242: note <= (-4563);
                11243: note <= (-377);
                11244: note <= 4815;
                11245: note <= 9889;
                11246: note <= 13722;
                11247: note <= 15491;
                11248: note <= 14886;
                11249: note <= 12187;
                11250: note <= 8192;
                11251: note <= 3995;
                11252: note <= 697;
                11253: note <= (-893);
                11254: note <= (-467);
                11255: note <= 1697;
                11256: note <= 4815;
                11257: note <= 7815;
                11258: note <= 9626;
                11259: note <= 9474;
                11260: note <= 7094;
                11261: note <= 2814;
                11262: note <= (-2531);
                11263: note <= (-7815);
                11264: note <= (-11910);
                11265: note <= (-13985);
                11266: note <= (-13722);
                11267: note <= (-11395);
                11268: note <= (-7791);
                11269: note <= (-3995);
                11270: note <= (-1098);
                11271: note <= 101;
                11272: note <= (-697);
                11273: note <= (-3203);
                11274: note <= (-6627);
                11275: note <= (-9889);
                11276: note <= (-11910);
                11277: note <= (-11911);
                11278: note <= (-9626);
                11279: note <= (-5378);
                11280: note <= 0;
                11281: note <= 5378;
                11282: note <= 9626;
                11283: note <= 11911;
                11284: note <= 11910;
                11285: note <= 9889;
                11286: note <= 6627;
                11287: note <= 3203;
                11288: note <= 697;
                11289: note <= (-101);
                11290: note <= 1098;
                11291: note <= 3995;
                11292: note <= 7791;
                11293: note <= 11395;
                11294: note <= 13722;
                11295: note <= 13985;
                11296: note <= 11910;
                11297: note <= 7815;
                11298: note <= 2531;
                11299: note <= (-2814);
                11300: note <= (-7094);
                11301: note <= (-9474);
                11302: note <= (-9626);
                11303: note <= (-7815);
                11304: note <= (-4815);
                11305: note <= (-1697);
                11306: note <= 467;
                11307: note <= 893;
                11308: note <= (-697);
                11309: note <= (-3995);
                11310: note <= (-8192);
                11311: note <= (-12187);
                11312: note <= (-14886);
                11313: note <= (-15491);
                11314: note <= (-13722);
                11315: note <= (-9889);
                11316: note <= (-4815);
                11317: note <= 377;
                11318: note <= 4563;
                11319: note <= 6910;
                11320: note <= 7094;
                11321: note <= 5378;
                11322: note <= 2531;
                11323: note <= (-377);
                11324: note <= (-2279);
                11325: note <= (-2399);
                11326: note <= (-467);
                11327: note <= 3203;
                11328: note <= 7791;
                11329: note <= 12187;
                11330: note <= 15286;
                11331: note <= 16283;
                11332: note <= 14886;
                11333: note <= 11395;
                11334: note <= 6627;
                11335: note <= 1697;
                11336: note <= (-2279);
                11337: note <= (-4473);
                11338: note <= (-4563);
                11339: note <= (-2814);
                11340: note <= 0;
                11341: note <= 2814;
                11342: note <= 4563;
                11343: note <= 4473;
                11344: note <= 2279;
                11345: note <= (-1697);
                11346: note <= (-6627);
                11347: note <= (-11395);
                11348: note <= (-14886);
                11349: note <= (-16283);
                11350: note <= (-15286);
                11351: note <= (-12187);
                11352: note <= (-7791);
                11353: note <= (-3203);
                11354: note <= 467;
                11355: note <= 2399;
                11356: note <= 2279;
                11357: note <= 377;
                11358: note <= (-2531);
                11359: note <= (-5378);
                11360: note <= (-7094);
                11361: note <= (-6910);
                11362: note <= (-4563);
                11363: note <= (-377);
                11364: note <= 4815;
                11365: note <= 9889;
                11366: note <= 13722;
                11367: note <= 15491;
                11368: note <= 14886;
                11369: note <= 12187;
                11370: note <= 8192;
                11371: note <= 3995;
                11372: note <= 697;
                11373: note <= (-893);
                11374: note <= (-467);
                11375: note <= 1697;
                11376: note <= 4815;
                11377: note <= 7815;
                11378: note <= 9626;
                11379: note <= 9474;
                11380: note <= 7094;
                11381: note <= 2814;
                11382: note <= (-2531);
                11383: note <= (-7815);
                11384: note <= (-11910);
                11385: note <= (-13985);
                11386: note <= (-13722);
                11387: note <= (-11395);
                11388: note <= (-7791);
                11389: note <= (-3995);
                11390: note <= (-1098);
                11391: note <= 101;
                11392: note <= (-697);
                11393: note <= (-3203);
                11394: note <= (-6627);
                11395: note <= (-9889);
                11396: note <= (-11910);
                11397: note <= (-11911);
                11398: note <= (-9626);
                11399: note <= (-5378);
                11400: note <= 0;
                11401: note <= 5378;
                11402: note <= 9626;
                11403: note <= 11911;
                11404: note <= 11910;
                11405: note <= 9889;
                11406: note <= 6627;
                11407: note <= 3203;
                11408: note <= 697;
                11409: note <= (-101);
                11410: note <= 1098;
                11411: note <= 3995;
                11412: note <= 7791;
                11413: note <= 11395;
                11414: note <= 13722;
                11415: note <= 13985;
                11416: note <= 11910;
                11417: note <= 7815;
                11418: note <= 2531;
                11419: note <= (-2814);
                11420: note <= (-7094);
                11421: note <= (-9474);
                11422: note <= (-9626);
                11423: note <= (-7815);
                11424: note <= (-4815);
                11425: note <= (-1697);
                11426: note <= 467;
                11427: note <= 893;
                11428: note <= (-697);
                11429: note <= (-3995);
                11430: note <= (-8192);
                11431: note <= (-12187);
                11432: note <= (-14886);
                11433: note <= (-15491);
                11434: note <= (-13722);
                11435: note <= (-9889);
                11436: note <= (-4815);
                11437: note <= 377;
                11438: note <= 4563;
                11439: note <= 6910;
                11440: note <= 7094;
                11441: note <= 5378;
                11442: note <= 2531;
                11443: note <= (-377);
                11444: note <= (-2279);
                11445: note <= (-2399);
                11446: note <= (-467);
                11447: note <= 3203;
                11448: note <= 7791;
                11449: note <= 12187;
                11450: note <= 15286;
                11451: note <= 16283;
                11452: note <= 14886;
                11453: note <= 11395;
                11454: note <= 6627;
                11455: note <= 1697;
                11456: note <= (-2279);
                11457: note <= (-4473);
                11458: note <= (-4563);
                11459: note <= (-2814);
                11460: note <= 0;
                11461: note <= 2814;
                11462: note <= 4563;
                11463: note <= 4473;
                11464: note <= 2279;
                11465: note <= (-1697);
                11466: note <= (-6627);
                11467: note <= (-11395);
                11468: note <= (-14886);
                11469: note <= (-16283);
                11470: note <= (-15286);
                11471: note <= (-12187);
                11472: note <= (-7791);
                11473: note <= (-3203);
                11474: note <= 467;
                11475: note <= 2399;
                11476: note <= 2279;
                11477: note <= 377;
                11478: note <= (-2531);
                11479: note <= (-5378);
                11480: note <= (-7094);
                11481: note <= (-6910);
                11482: note <= (-4563);
                11483: note <= (-377);
                11484: note <= 4815;
                11485: note <= 9889;
                11486: note <= 13722;
                11487: note <= 15491;
                11488: note <= 14886;
                11489: note <= 12187;
                11490: note <= 8192;
                11491: note <= 3995;
                11492: note <= 697;
                11493: note <= (-893);
                11494: note <= (-467);
                11495: note <= 1697;
                11496: note <= 4815;
                11497: note <= 7815;
                11498: note <= 9626;
                11499: note <= 9474;
                11500: note <= 7094;
                11501: note <= 2814;
                11502: note <= (-2531);
                11503: note <= (-7815);
                11504: note <= (-11910);
                11505: note <= (-13985);
                11506: note <= (-13722);
                11507: note <= (-11395);
                11508: note <= (-7791);
                11509: note <= (-3995);
                11510: note <= (-1098);
                11511: note <= 101;
                11512: note <= (-697);
                11513: note <= (-3203);
                11514: note <= (-6627);
                11515: note <= (-9889);
                11516: note <= (-11910);
                11517: note <= (-11911);
                11518: note <= (-9626);
                11519: note <= (-5378);
                11520: note <= 0;
                11521: note <= 5378;
                11522: note <= 9626;
                11523: note <= 11911;
                11524: note <= 11910;
                11525: note <= 9889;
                11526: note <= 6627;
                11527: note <= 3203;
                11528: note <= 697;
                11529: note <= (-101);
                11530: note <= 1098;
                11531: note <= 3995;
                11532: note <= 7791;
                11533: note <= 11395;
                11534: note <= 13722;
                11535: note <= 13985;
                11536: note <= 11910;
                11537: note <= 7815;
                11538: note <= 2531;
                11539: note <= (-2814);
                11540: note <= (-7094);
                11541: note <= (-9474);
                11542: note <= (-9626);
                11543: note <= (-7815);
                11544: note <= (-4815);
                11545: note <= (-1697);
                11546: note <= 467;
                11547: note <= 893;
                11548: note <= (-697);
                11549: note <= (-3995);
                11550: note <= (-8192);
                11551: note <= (-12187);
                11552: note <= (-14886);
                11553: note <= (-15491);
                11554: note <= (-13722);
                11555: note <= (-9889);
                11556: note <= (-4815);
                11557: note <= 377;
                11558: note <= 4563;
                11559: note <= 6910;
                11560: note <= 7094;
                11561: note <= 5378;
                11562: note <= 2531;
                11563: note <= (-377);
                11564: note <= (-2279);
                11565: note <= (-2399);
                11566: note <= (-467);
                11567: note <= 3203;
                11568: note <= 7791;
                11569: note <= 12187;
                11570: note <= 15286;
                11571: note <= 16283;
                11572: note <= 14886;
                11573: note <= 11395;
                11574: note <= 6627;
                11575: note <= 1697;
                11576: note <= (-2279);
                11577: note <= (-4473);
                11578: note <= (-4563);
                11579: note <= (-2814);
                11580: note <= 0;
                11581: note <= 2814;
                11582: note <= 4563;
                11583: note <= 4473;
                11584: note <= 2279;
                11585: note <= (-1697);
                11586: note <= (-6627);
                11587: note <= (-11395);
                11588: note <= (-14886);
                11589: note <= (-16283);
                11590: note <= (-15286);
                11591: note <= (-12187);
                11592: note <= (-7791);
                11593: note <= (-3203);
                11594: note <= 467;
                11595: note <= 2399;
                11596: note <= 2279;
                11597: note <= 377;
                11598: note <= (-2531);
                11599: note <= (-5378);
                11600: note <= (-7094);
                11601: note <= (-6910);
                11602: note <= (-4563);
                11603: note <= (-377);
                11604: note <= 4815;
                11605: note <= 9889;
                11606: note <= 13722;
                11607: note <= 15491;
                11608: note <= 14886;
                11609: note <= 12187;
                11610: note <= 8192;
                11611: note <= 3995;
                11612: note <= 697;
                11613: note <= (-893);
                11614: note <= (-467);
                11615: note <= 1697;
                11616: note <= 4815;
                11617: note <= 7815;
                11618: note <= 9626;
                11619: note <= 9474;
                11620: note <= 7094;
                11621: note <= 2814;
                11622: note <= (-2531);
                11623: note <= (-7815);
                11624: note <= (-11910);
                11625: note <= (-13985);
                11626: note <= (-13722);
                11627: note <= (-11395);
                11628: note <= (-7791);
                11629: note <= (-3995);
                11630: note <= (-1098);
                11631: note <= 101;
                11632: note <= (-697);
                11633: note <= (-3203);
                11634: note <= (-6627);
                11635: note <= (-9889);
                11636: note <= (-11910);
                11637: note <= (-11911);
                11638: note <= (-9626);
                11639: note <= (-5378);
                11640: note <= 0;
                11641: note <= 5378;
                11642: note <= 9626;
                11643: note <= 11911;
                11644: note <= 11910;
                11645: note <= 9889;
                11646: note <= 6627;
                11647: note <= 3203;
                11648: note <= 697;
                11649: note <= (-101);
                11650: note <= 1098;
                11651: note <= 3995;
                11652: note <= 7791;
                11653: note <= 11395;
                11654: note <= 13722;
                11655: note <= 13985;
                11656: note <= 11910;
                11657: note <= 7815;
                11658: note <= 2531;
                11659: note <= (-2814);
                11660: note <= (-7094);
                11661: note <= (-9474);
                11662: note <= (-9626);
                11663: note <= (-7815);
                11664: note <= (-4815);
                11665: note <= (-1697);
                11666: note <= 467;
                11667: note <= 893;
                11668: note <= (-697);
                11669: note <= (-3995);
                11670: note <= (-8192);
                11671: note <= (-12187);
                11672: note <= (-14886);
                11673: note <= (-15491);
                11674: note <= (-13722);
                11675: note <= (-9889);
                11676: note <= (-4815);
                11677: note <= 377;
                11678: note <= 4563;
                11679: note <= 6910;
                11680: note <= 7094;
                11681: note <= 5378;
                11682: note <= 2531;
                11683: note <= (-377);
                11684: note <= (-2279);
                11685: note <= (-2399);
                11686: note <= (-467);
                11687: note <= 3203;
                11688: note <= 7791;
                11689: note <= 12187;
                11690: note <= 15286;
                11691: note <= 16283;
                11692: note <= 14886;
                11693: note <= 11395;
                11694: note <= 6627;
                11695: note <= 1697;
                11696: note <= (-2279);
                11697: note <= (-4473);
                11698: note <= (-4563);
                11699: note <= (-2814);
                11700: note <= 0;
                11701: note <= 2814;
                11702: note <= 4563;
                11703: note <= 4473;
                11704: note <= 2279;
                11705: note <= (-1697);
                11706: note <= (-6627);
                11707: note <= (-11395);
                11708: note <= (-14886);
                11709: note <= (-16283);
                11710: note <= (-15286);
                11711: note <= (-12187);
                11712: note <= (-7791);
                11713: note <= (-3203);
                11714: note <= 467;
                11715: note <= 2399;
                11716: note <= 2279;
                11717: note <= 377;
                11718: note <= (-2531);
                11719: note <= (-5378);
                11720: note <= (-7094);
                11721: note <= (-6910);
                11722: note <= (-4563);
                11723: note <= (-377);
                11724: note <= 4815;
                11725: note <= 9889;
                11726: note <= 13722;
                11727: note <= 15491;
                11728: note <= 14886;
                11729: note <= 12187;
                11730: note <= 8192;
                11731: note <= 3995;
                11732: note <= 697;
                11733: note <= (-893);
                11734: note <= (-467);
                11735: note <= 1697;
                11736: note <= 4815;
                11737: note <= 7815;
                11738: note <= 9626;
                11739: note <= 9474;
                11740: note <= 7094;
                11741: note <= 2814;
                11742: note <= (-2531);
                11743: note <= (-7815);
                11744: note <= (-11910);
                11745: note <= (-13985);
                11746: note <= (-13722);
                11747: note <= (-11395);
                11748: note <= (-7791);
                11749: note <= (-3995);
                11750: note <= (-1098);
                11751: note <= 101;
                11752: note <= (-697);
                11753: note <= (-3203);
                11754: note <= (-6627);
                11755: note <= (-9889);
                11756: note <= (-11910);
                11757: note <= (-11911);
                11758: note <= (-9626);
                11759: note <= (-5378);
                11760: note <= 0;
                11761: note <= 5378;
                11762: note <= 9626;
                11763: note <= 11911;
                11764: note <= 11910;
                11765: note <= 9889;
                11766: note <= 6627;
                11767: note <= 3203;
                11768: note <= 697;
                11769: note <= (-101);
                11770: note <= 1098;
                11771: note <= 3995;
                11772: note <= 7791;
                11773: note <= 11395;
                11774: note <= 13722;
                11775: note <= 13985;
                11776: note <= 11910;
                11777: note <= 7815;
                11778: note <= 2531;
                11779: note <= (-2814);
                11780: note <= (-7094);
                11781: note <= (-9474);
                11782: note <= (-9626);
                11783: note <= (-7815);
                11784: note <= (-4815);
                11785: note <= (-1697);
                11786: note <= 467;
                11787: note <= 893;
                11788: note <= (-697);
                11789: note <= (-3995);
                11790: note <= (-8192);
                11791: note <= (-12187);
                11792: note <= (-14886);
                11793: note <= (-15491);
                11794: note <= (-13722);
                11795: note <= (-9889);
                11796: note <= (-4815);
                11797: note <= 377;
                11798: note <= 4563;
                11799: note <= 6910;
                11800: note <= 7094;
                11801: note <= 5378;
                11802: note <= 2531;
                11803: note <= (-377);
                11804: note <= (-2279);
                11805: note <= (-2399);
                11806: note <= (-467);
                11807: note <= 3203;
                11808: note <= 7791;
                11809: note <= 12187;
                11810: note <= 15286;
                11811: note <= 16283;
                11812: note <= 14886;
                11813: note <= 11395;
                11814: note <= 6627;
                11815: note <= 1697;
                11816: note <= (-2279);
                11817: note <= (-4473);
                11818: note <= (-4563);
                11819: note <= (-2814);
                11820: note <= 0;
                11821: note <= 2814;
                11822: note <= 4563;
                11823: note <= 4473;
                11824: note <= 2279;
                11825: note <= (-1697);
                11826: note <= (-6627);
                11827: note <= (-11395);
                11828: note <= (-14886);
                11829: note <= (-16283);
                11830: note <= (-15286);
                11831: note <= (-12187);
                11832: note <= (-7791);
                11833: note <= (-3203);
                11834: note <= 467;
                11835: note <= 2399;
                11836: note <= 2279;
                11837: note <= 377;
                11838: note <= (-2531);
                11839: note <= (-5378);
                11840: note <= (-7094);
                11841: note <= (-6910);
                11842: note <= (-4563);
                11843: note <= (-377);
                11844: note <= 4815;
                11845: note <= 9889;
                11846: note <= 13722;
                11847: note <= 15491;
                11848: note <= 14886;
                11849: note <= 12187;
                11850: note <= 8192;
                11851: note <= 3995;
                11852: note <= 697;
                11853: note <= (-893);
                11854: note <= (-467);
                11855: note <= 1697;
                11856: note <= 4815;
                11857: note <= 7815;
                11858: note <= 9626;
                11859: note <= 9474;
                11860: note <= 7094;
                11861: note <= 2814;
                11862: note <= (-2531);
                11863: note <= (-7815);
                11864: note <= (-11910);
                11865: note <= (-13985);
                11866: note <= (-13722);
                11867: note <= (-11395);
                11868: note <= (-7791);
                11869: note <= (-3995);
                11870: note <= (-1098);
                11871: note <= 101;
                11872: note <= (-697);
                11873: note <= (-3203);
                11874: note <= (-6627);
                11875: note <= (-9889);
                11876: note <= (-11910);
                11877: note <= (-11911);
                11878: note <= (-9626);
                11879: note <= (-5378);
                11880: note <= 0;
                11881: note <= 5378;
                11882: note <= 9626;
                11883: note <= 11911;
                11884: note <= 11910;
                11885: note <= 9889;
                11886: note <= 6627;
                11887: note <= 3203;
                11888: note <= 697;
                11889: note <= (-101);
                11890: note <= 1098;
                11891: note <= 3995;
                11892: note <= 7791;
                11893: note <= 11395;
                11894: note <= 13722;
                11895: note <= 13985;
                11896: note <= 11910;
                11897: note <= 7815;
                11898: note <= 2531;
                11899: note <= (-2814);
                11900: note <= (-7094);
                11901: note <= (-9474);
                11902: note <= (-9626);
                11903: note <= (-7815);
                11904: note <= (-4815);
                11905: note <= (-1697);
                11906: note <= 467;
                11907: note <= 893;
                11908: note <= (-697);
                11909: note <= (-3995);
                11910: note <= (-8192);
                11911: note <= (-12187);
                11912: note <= (-14886);
                11913: note <= (-15491);
                11914: note <= (-13722);
                11915: note <= (-9889);
                11916: note <= (-4815);
                11917: note <= 377;
                11918: note <= 4563;
                11919: note <= 6910;
                11920: note <= 7094;
                11921: note <= 5378;
                11922: note <= 2531;
                11923: note <= (-377);
                11924: note <= (-2279);
                11925: note <= (-2399);
                11926: note <= (-467);
                11927: note <= 3203;
                11928: note <= 7791;
                11929: note <= 12187;
                11930: note <= 15286;
                11931: note <= 16283;
                11932: note <= 14886;
                11933: note <= 11395;
                11934: note <= 6627;
                11935: note <= 1697;
                11936: note <= (-2279);
                11937: note <= (-4473);
                11938: note <= (-4563);
                11939: note <= (-2814);
                11940: note <= 0;
                11941: note <= 2814;
                11942: note <= 4563;
                11943: note <= 4473;
                11944: note <= 2279;
                11945: note <= (-1697);
                11946: note <= (-6627);
                11947: note <= (-11395);
                11948: note <= (-14886);
                11949: note <= (-16283);
                11950: note <= (-15286);
                11951: note <= (-12187);
                11952: note <= (-7791);
                11953: note <= (-3203);
                11954: note <= 467;
                11955: note <= 2399;
                11956: note <= 2279;
                11957: note <= 377;
                11958: note <= (-2531);
                11959: note <= (-5378);
                11960: note <= (-7094);
                11961: note <= (-6910);
                11962: note <= (-4563);
                11963: note <= (-377);
                11964: note <= 4815;
                11965: note <= 9889;
                11966: note <= 13722;
                11967: note <= 15491;
                11968: note <= 14886;
                11969: note <= 12187;
                11970: note <= 8192;
                11971: note <= 3995;
                11972: note <= 697;
                11973: note <= (-893);
                11974: note <= (-467);
                11975: note <= 1697;
                11976: note <= 4815;
                11977: note <= 7815;
                11978: note <= 9626;
                11979: note <= 9474;
                11980: note <= 7094;
                11981: note <= 2814;
                11982: note <= (-2531);
                11983: note <= (-7815);
                11984: note <= (-11910);
                11985: note <= (-13985);
                11986: note <= (-13722);
                11987: note <= (-11395);
                11988: note <= (-7791);
                11989: note <= (-3995);
                11990: note <= (-1098);
                11991: note <= 101;
                11992: note <= (-697);
                11993: note <= (-3203);
                11994: note <= (-6627);
                11995: note <= (-9889);
                11996: note <= (-11910);
                11997: note <= (-11911);
                11998: note <= (-9626);
                default: note <= (-5378);
            endcase
            nv <= 1'b1;
            noteidx <= ($signed({1'b0, noteidx}) < (12000 - 1)) ? (noteidx + 1) : 0;
        end
        else begin
            sample_rate_cnt <= (sample_rate_cnt + 1);
            nv <= 1'b0;
        end
    end
end
endmodule