module header
    // Internal signals
		// Generated Signal List
		// End of Generated Signal List
    // %COMPILER_OPTS%
    //TODO: %VERI_CONSTANTS%
    // %VERI_CONCURS%
	// Generated Signal Assignments
    // Generated Instances
    // wiring ...
	// Generated Instances and Port Mappings
		// Generated Instance Port Map for inst_ba
		ent_ba inst_ba(
		);// End of Generated Instance Port Map for inst_ba
		// Generated Instance Port Map for inst_bb
		ent_bb inst_bb(
		);// End of Generated Instance Port Map for inst_bb
endmodule