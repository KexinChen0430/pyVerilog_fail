module alu_ctrl ( .OP({\OP[4] , \OP[3] , \OP[2] , \OP[1] , \OP[0] }), ALU_WORD
 );
  output [12:0] ALU_WORD;
  input \OP[4] , \OP[3] , \OP[2] , \OP[1] , \OP[0] ;
  wire   N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, N33,
         n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35;
  DLH_X1 \comp_sel_reg[2]  ( .G(N32), .D(N33), .Q(ALU_WORD[4]) );
  DLH_X1 \comp_sel_reg[1]  ( .G(N32), .D(N31), .Q(ALU_WORD[3]) );
  DLH_X1 \comp_sel_reg[0]  ( .G(N32), .D(N30), .Q(ALU_WORD[2]) );
  DLH_X1 sign_to_booth_reg ( .G(N20), .D(N21), .Q(ALU_WORD[0]) );
  DLH_X1 left_right_reg ( .G(N23), .D(N22), .Q(ALU_WORD[9]) );
  DLH_X1 logic_arith_reg ( .G(N23), .D(N24), .Q(ALU_WORD[8]) );
  DLH_X1 sign_to_adder_reg ( .G(N25), .D(N26), .Q(ALU_WORD[7]) );
  DLH_X1 \lu_ctrl_reg[1]  ( .G(N28), .D(N29), .Q(ALU_WORD[6]) );
  DLH_X1 \lu_ctrl_reg[0]  ( .G(N28), .D(N27), .Q(ALU_WORD[5]) );
  NAND3_X1 U53 ( .A1(n9), .A2(OP[1]), .A3(n28), .ZN(n30) );
  NAND3_X1 U54 ( .A1(n15), .A2(n35), .A3(n22), .ZN(n19) );
  NOR3_X1 U48 ( .A1(OP[2]), .A2(OP[0]), .A3(n22), .ZN(n10) );
  NAND2_X1 U47 ( .A1(OP[3]), .A2(n23), .ZN(n3) );
  NOR3_X1 U45 ( .A1(OP[2]), .A2(n35), .A3(n22), .ZN(n33) );
  NOR2_X1 U43 ( .A1(n3), .A2(n2), .ZN(n32) );
  NOR2_X1 U41 ( .A1(OP[0]), .A2(n15), .ZN(n28) );
  NAND2_X1 U40 ( .A1(n28), .A2(n22), .ZN(n1) );
  NOR2_X1 U39 ( .A1(n19), .A2(OP[3]), .ZN(n34) );
  NOR4_X1 U38 ( .A1(n15), .A2(n3), .A3(n35), .A4(n22), .ZN(n8) );
  AOI21_X1 U37 ( .B1(n34), .B2(OP[4]), .A(n8), .ZN(n18) );
  NAND2_X1 U36 ( .A1(n33), .A2(n26), .ZN(n6) );
  OAI211_X1 U35 ( .C1(n1), .C2(n16), .A(n18), .B(n6), .ZN(N30) );
  AOI211_X1 U34 ( .C1(n26), .C2(n10), .A(n32), .B(N30), .ZN(n29) );
  NAND2_X1 U33 ( .A1(OP[0]), .A2(n22), .ZN(n27) );
  NOR2_X1 U32 ( .A1(n3), .A2(n27), .ZN(n31) );
  NAND2_X1 U31 ( .A1(OP[2]), .A2(n31), .ZN(n4) );
  NOR2_X1 U29 ( .A1(OP[2]), .A2(n27), .ZN(n24) );
  NAND2_X1 U28 ( .A1(n26), .A2(n24), .ZN(n7) );
  NAND4_X1 U27 ( .A1(n29), .A2(n4), .A3(n30), .A4(n7), .ZN(N32) );
  AOI211_X1 U26 ( .C1(OP[0]), .C2(OP[1]), .A(OP[2]), .B(n3), .ZN(N28) );
  NAND2_X1 U25 ( .A1(OP[1]), .A2(n28), .ZN(n17) );
  OAI21_X1 U24 ( .B1(n27), .B2(n15), .A(n17), .ZN(n25) );
  NAND2_X1 U23 ( .A1(n25), .A2(n26), .ZN(n20) );
  NOR3_X1 U18 ( .A1(OP[2]), .A2(n22), .A3(n13), .ZN(N22) );
  OAI21_X1 U16 ( .B1(n11), .B2(n13), .A(n21), .ZN(N23) );
  OAI21_X1 U14 ( .B1(n19), .B2(n13), .A(n20), .ZN(ALU_WORD[12]) );
  NOR2_X1 U6 ( .A1(n3), .A2(n11), .ZN(N27) );
  NAND2_X1 U8 ( .A1(OP[2]), .A2(OP[1]), .ZN(n12) );
  OAI21_X1 U7 ( .B1(n12), .B2(n13), .A(n14), .ZN(N26) );
  NOR2_X1 U11 ( .A1(n2), .A2(n13), .ZN(N24) );
  OAI211_X1 U12 ( .C1(n16), .C2(n17), .A(n18), .B(n4), .ZN(N21) );
  NAND4_X1 U3 ( .A1(n4), .A2(n5), .A3(n6), .A4(n7), .ZN(N31) );
  AOI21_X1 U2 ( .B1(n1), .B2(n2), .A(n3), .ZN(N33) );
  OAI21_X1 U9 ( .B1(n15), .B2(n13), .A(n14), .ZN(N25) );
  NAND2_X1 U19 ( .A1(n23), .A2(n16), .ZN(n13) );
  NOR2_X1 U50 ( .A1(n23), .A2(n16), .ZN(n26) );
  INV_X1 U52 ( .A(OP[4]), .ZN(n23) );
  INV_X1 U51 ( .A(OP[3]), .ZN(n16) );
  INV_X1 U49 ( .A(OP[1]), .ZN(n22) );
  INV_X1 U46 ( .A(OP[0]), .ZN(n35) );
  INV_X1 U44 ( .A(n33), .ZN(n2) );
  INV_X1 U42 ( .A(OP[2]), .ZN(n15) );
  INV_X1 U30 ( .A(n3), .ZN(n9) );
  INV_X1 U22 ( .A(n20), .ZN(ALU_WORD[1]) );
  OR3_X1 U21 ( .A1(N32), .A2(N28), .A3(ALU_WORD[1]), .ZN(ALU_WORD[10]) );
  INV_X1 U20 ( .A(n24), .ZN(n11) );
  INV_X1 U17 ( .A(N22), .ZN(n21) );
  OR2_X1 U15 ( .A1(N32), .A2(N23), .ZN(ALU_WORD[11]) );
  AND2_X1 U5 ( .A1(n9), .A2(n10), .ZN(N29) );
  INV_X1 U10 ( .A(N32), .ZN(n14) );
  INV_X1 U4 ( .A(n8), .ZN(n5) );
  OR2_X1 U13 ( .A1(N32), .A2(ALU_WORD[12]), .ZN(N20) );
endmodule