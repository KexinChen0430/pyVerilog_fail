module to control the memory
	// MC0 even request port signals
	assign mc0_req_ld_e         = r_mc0_req_ld_e;
	assign mc0_req_st_e			= r_mc0_req_st_e;
	assign mc0_req_size_e		= r_mc0_req_size_e;
	assign mc0_req_vadr_e		= r_mc0_req_vadr_e;
	assign mc0_req_wrd_rdctl_e	= r_mc0_req_wrd_rdctl_e;
	assign mc0_req_flush_e		= r_mc0_req_flush_e;
	// MC0 even response port signals
	assign mc0_rsp_stall_e		= r_mc0_rsp_stall_e;
	// MC0 odd request port signals
	assign mc0_req_ld_o			= r_mc0_req_ld_o;
	assign mc0_req_st_o			= r_mc0_req_st_o;
	assign mc0_req_size_o		= r_mc0_req_size_o;
	assign mc0_req_vadr_o		= r_mc0_req_vadr_o;
	assign mc0_req_wrd_rdctl_o	= r_mc0_req_wrd_rdctl_o;
	assign mc0_req_flush_o		= r_mc0_req_flush_o;
	// MC0 odd response port signals
	assign mc0_rsp_stall_o		= r_mc0_rsp_stall_o;
	// MC1 even request port signals
	assign mc1_req_ld_e			= r_mc1_req_ld_e;
	assign mc1_req_st_e			= r_mc1_req_st_e;
	assign mc1_req_size_e		= r_mc1_req_size_e;
	assign mc1_req_vadr_e		= r_mc1_req_vadr_e;
	assign mc1_req_wrd_rdctl_e	= r_mc1_req_wrd_rdctl_e;
	assign mc1_req_flush_e		= r_mc1_req_flush_e;
	// MC1 even response port signals
	assign mc1_rsp_stall_e		= r_mc1_rsp_stall_e;
	// MC1 odd request port signals
	assign mc1_req_ld_o			= r_mc1_req_ld_o;
	assign mc1_req_st_o			= r_mc1_req_st_o;
	assign mc1_req_size_o		= r_mc1_req_size_o;
	assign mc1_req_vadr_o		= r_mc1_req_vadr_o;
	assign mc1_req_wrd_rdctl_o	= r_mc1_req_wrd_rdctl_o;
	assign mc1_req_flush_o		= r_mc1_req_flush_o;
	// MC1 odd response port signals
	assign mc1_rsp_stall_o		= r_mc1_rsp_stall_o;
	// MC2 even request port signals
	assign mc2_req_ld_e			= r_mc2_req_ld_e;
	assign mc2_req_st_e			= r_mc2_req_st_e;
	assign mc2_req_size_e		= r_mc2_req_size_e;
	assign mc2_req_vadr_e		= r_mc2_req_vadr_e;
	assign mc2_req_wrd_rdctl_e	= r_mc2_req_wrd_rdctl_e;
	assign mc2_req_flush_e		= r_mc2_req_flush_e;
	// MC2 even response port signals
	assign mc2_rsp_stall_e		= r_mc2_rsp_stall_e;
	// MC2 odd request port signals
	assign mc2_req_ld_o			= r_mc2_req_ld_o;
	assign mc2_req_st_o			= r_mc2_req_st_o;
	assign mc2_req_size_o		= r_mc2_req_size_o;
	assign mc2_req_vadr_o		= r_mc2_req_vadr_o;
	assign mc2_req_wrd_rdctl_o	= r_mc2_req_wrd_rdctl_o;
	assign mc2_req_flush_o		= r_mc2_req_flush_o;
	// MC2 odd response port signals
	assign mc2_rsp_stall_o		= r_mc2_rsp_stall_o;
	// MC3 even request port signals
	assign mc3_req_ld_e			= r_mc3_req_ld_e;
	assign mc3_req_st_e			= r_mc3_req_st_e;
	assign mc3_req_size_e		= r_mc3_req_size_e;
	assign mc3_req_vadr_e		= r_mc3_req_vadr_e;
	assign mc3_req_wrd_rdctl_e	= r_mc3_req_wrd_rdctl_e;
	assign mc3_req_flush_e		= r_mc3_req_flush_e;
	// MC3 even response port signals
	assign mc3_rsp_stall_e		= r_mc3_rsp_stall_e;
	// MC3 odd request port signals
	assign mc3_req_ld_o			= r_mc3_req_ld_o;
	assign mc3_req_st_o			= r_mc3_req_st_o;
	assign mc3_req_size_o		= r_mc3_req_size_o;
	assign mc3_req_vadr_o		= r_mc3_req_vadr_o;
	assign mc3_req_wrd_rdctl_o	= r_mc3_req_wrd_rdctl_o;
	assign mc3_req_flush_o		= r_mc3_req_flush_o;
	// MC3 odd response port signals
	assign mc3_rsp_stall_o		= r_mc3_rsp_stall_o;
	// MC4 even request port signals
	assign mc4_req_ld_e			= r_mc4_req_ld_e;
	assign mc4_req_st_e			= r_mc4_req_st_e;
	assign mc4_req_size_e		= r_mc4_req_size_e;
	assign mc4_req_vadr_e		= r_mc4_req_vadr_e;
	assign mc4_req_wrd_rdctl_e	= r_mc4_req_wrd_rdctl_e;
	assign mc4_req_flush_e		= r_mc4_req_flush_e;
	// MC4 even response port signals
	assign mc4_rsp_stall_e		= r_mc4_rsp_stall_e;
	// MC4 odd request port signals
	assign mc4_req_ld_o			= r_mc4_req_ld_o;
	assign mc4_req_st_o			= r_mc4_req_st_o;
	assign mc4_req_size_o		= r_mc4_req_size_o;
	assign mc4_req_vadr_o		= r_mc4_req_vadr_o;
	assign mc4_req_wrd_rdctl_o	= r_mc4_req_wrd_rdctl_o;
	assign mc4_req_flush_o		= r_mc4_req_flush_o;
	// MC4 odd response port signals
	assign mc4_rsp_stall_o		= r_mc4_rsp_stall_o;
	// MC5 even request port signals
	assign mc5_req_ld_e			= r_mc5_req_ld_e;
	assign mc5_req_st_e			= r_mc5_req_st_e;
	assign mc5_req_size_e		= r_mc5_req_size_e;
	assign mc5_req_vadr_e		= r_mc5_req_vadr_e;
	assign mc5_req_wrd_rdctl_e	= r_mc5_req_wrd_rdctl_e;
	assign mc5_req_flush_e		= r_mc5_req_flush_e;
	// MC5 even response port signals
	assign mc5_rsp_stall_e		= r_mc5_rsp_stall_e;
	// MC5 odd request port signals
	assign mc5_req_ld_o			= r_mc5_req_ld_o;
	assign mc5_req_st_o			= r_mc5_req_st_o;
	assign mc5_req_size_o		= r_mc5_req_size_o;
	assign mc5_req_vadr_o		= r_mc5_req_vadr_o;
	assign mc5_req_wrd_rdctl_o	= r_mc5_req_wrd_rdctl_o;
	assign mc5_req_flush_o		= r_mc5_req_flush_o;
	// MC5 odd response port signals
	assign mc5_rsp_stall_o		= r_mc5_rsp_stall_o;
	// MC6 even request port signals
	assign mc6_req_ld_e			= r_mc6_req_ld_e;
	assign mc6_req_st_e			= r_mc6_req_st_e;
	assign mc6_req_size_e		= r_mc6_req_size_e;
	assign mc6_req_vadr_e		= r_mc6_req_vadr_e;
	assign mc6_req_wrd_rdctl_e	= r_mc6_req_wrd_rdctl_e;
	assign mc6_req_flush_e		= r_mc6_req_flush_e;
	// MC6 even response port signals
	assign mc6_rsp_stall_e		= r_mc6_rsp_stall_e;
	// MC6 odd request port signals
	assign mc6_req_ld_o			= r_mc6_req_ld_o;
	assign mc6_req_st_o			= r_mc6_req_st_o;
	assign mc6_req_size_o		= r_mc6_req_size_o;
	assign mc6_req_vadr_o		= r_mc6_req_vadr_o;
	assign mc6_req_wrd_rdctl_o	= r_mc6_req_wrd_rdctl_o;
	assign mc6_req_flush_o		= r_mc6_req_flush_o;
	// MC6 odd response port signals
	assign mc6_rsp_stall_o		= r_mc6_rsp_stall_o;
	// MC7 even request port signals
	assign mc7_req_ld_e			= r_mc7_req_ld_e;
	assign mc7_req_st_e			= r_mc7_req_st_e;
	assign mc7_req_size_e		= r_mc7_req_size_e;
	assign mc7_req_vadr_e		= r_mc7_req_vadr_e;
	assign mc7_req_wrd_rdctl_e	= r_mc7_req_wrd_rdctl_e;
	assign mc7_req_flush_e		= r_mc7_req_flush_e;
	// MC7 even response port signals
	assign mc7_rsp_stall_e		= r_mc7_rsp_stall_e;
	// MC7 odd request port signals
	assign mc7_req_ld_o			= r_mc7_req_ld_o;
	assign mc7_req_st_o			= r_mc7_req_st_o;
	assign mc7_req_size_o		= r_mc7_req_size_o;
	assign mc7_req_vadr_o		= r_mc7_req_vadr_o;
	assign mc7_req_wrd_rdctl_o	= r_mc7_req_wrd_rdctl_o;
	assign mc7_req_flush_o		= r_mc7_req_flush_o;
	// MC7 odd response port signals
	assign mc7_rsp_stall_o		= r_mc7_rsp_stall_o;
	/* ---------- debug & synopsys off blocks  ---------- */
	// synopsys translate_off
	// Parameters: 1-Severity: Don't Stop, 2-start check only after negedge of reset
	//assert_never #(1, 2, "***ERROR ASSERT: unimplemented instruction cracked") a0 (.clk(clk), .reset_n(~reset), .test_expr(r_unimplemented_inst));
	// synopsys translate_on
endmodule