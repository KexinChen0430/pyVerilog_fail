module header
	// Internal signals
	// Generated Signal List
	// End of Generated Signal List
	// %COMPILER_OPTS%
	// Generated Signal Assignments
	// Generated Instances and Port Mappings
		// Generated Instance Port Map for inst_eaa
		inst_eaa_e inst_eaa (
		);
		// End of Generated Instance Port Map for inst_eaa
		// Generated Instance Port Map for inst_eab
		inst_eab_e inst_eab (
		);
		// End of Generated Instance Port Map for inst_eab
		// Generated Instance Port Map for inst_eac
		inst_eac_e inst_eac (
		);
		// End of Generated Instance Port Map for inst_eac
		// Generated Instance Port Map for inst_ead
		inst_ead_e inst_ead (
		);
		// End of Generated Instance Port Map for inst_ead
endmodule