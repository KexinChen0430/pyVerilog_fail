module pcc2_cfg;
  generate
   `simple_svfcov_clk(a, b, c, d);
  endgenerate
endmodule