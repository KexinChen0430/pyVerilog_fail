module DSP_M_DATA #(
`ifdef XIL_TIMING
  parameter LOC = "UNPLACED",
`endif
  parameter [0:0] IS_CLK_INVERTED = 1'b0,
  parameter [0:0] IS_RSTM_INVERTED = 1'b0,
  parameter integer MREG = 1
)(
  output [44:0] U_DATA,
  output [44:0] V_DATA,
  input CEM,
  input CLK,
  input RSTM,
  input [44:0] U,
  input [44:0] V
);
// define constants
  localparam MODULE_NAME = "DSP_M_DATA";
  reg trig_attr;
// include dynamic registers - XILINX test only
`ifdef XIL_DR
  `include "DSP_M_DATA_dr.v"
`else
  reg [0:0] IS_CLK_INVERTED_REG = IS_CLK_INVERTED;
  reg [0:0] IS_RSTM_INVERTED_REG = IS_RSTM_INVERTED;
  reg [31:0] MREG_REG = MREG;
`endif
`ifdef XIL_XECLIB
  wire MREG_BIN;
`else
  reg MREG_BIN;
`endif
`ifdef XIL_XECLIB
  reg glblGSR = 1'b0;
`else
  tri0 glblGSR = glbl.GSR;
`endif
  wire CEM_in;
  wire CLK_in;
  wire RSTM_in;
  wire [44:0] U_in;
  wire [44:0] V_in;
`ifdef XIL_TIMING
  wire CEM_delay;
  wire CLK_delay;
  wire RSTM_delay;
  wire [44:0] U_delay;
  wire [44:0] V_delay;
`endif
`ifdef XIL_TIMING
// bus inputs with only partial timing checks
  assign U_delay[44] = U[44];
  assign V_delay[1] = V[1];
  assign V_delay[2] = V[2];
  assign V_delay[3] = V[3];
  assign V_delay[44] = V[44];
`endif
`ifdef XIL_TIMING
  assign CEM_in = (CEM !== 1'bz) && CEM_delay; // rv 0
  assign CLK_in = (CLK !== 1'bz) && (CLK_delay ^ IS_CLK_INVERTED_REG); // rv 0
  assign RSTM_in = (RSTM !== 1'bz) && (RSTM_delay ^ IS_RSTM_INVERTED_REG); // rv 0
  assign U_in = U_delay;
  assign V_in = V_delay;
`else
  assign CEM_in = (CEM !== 1'bz) && CEM; // rv 0
  assign CLK_in = (CLK !== 1'bz) && (CLK ^ IS_CLK_INVERTED_REG); // rv 0
  assign RSTM_in = (RSTM !== 1'bz) && (RSTM ^ IS_RSTM_INVERTED_REG); // rv 0
  assign U_in = U;
  assign V_in = V;
`endif
`ifndef XIL_XECLIB
  reg attr_test;
  reg attr_err;
initial begin
  trig_attr = 1'b0;
`ifdef XIL_ATTR_TEST
  attr_test = 1'b1;
`else
  attr_test = 1'b0;
`endif
  attr_err = 1'b0;
  #1;
  trig_attr = ~trig_attr;
end
`endif
`ifdef XIL_XECLIB
  assign MREG_BIN = MREG_REG[0];
`else
always @(trig_attr) begin
#1;
  MREG_BIN = MREG_REG[0];
end
`endif
`ifndef XIL_TIMING
  initial begin
    $display("Error: [Unisim %s-100] SIMPRIM primitive is not intended for direct instantiation in RTL or functional netlists. This primitive is only available in the SIMPRIM library for implemented netlists, please ensure you are pointing to the correct library. Instance %m", MODULE_NAME);
    #1 $finish;
  end
`endif
`ifndef XIL_XECLIB
  always @(trig_attr) begin
  #1;
    if ((attr_test == 1'b1) ||
        ((MREG_REG != 1) &&
         (MREG_REG != 0))) begin
      $display("Error: [Unisim %s-103] MREG attribute is set to %d.  Legal values for this attribute are 1 or 0. Instance: %m", MODULE_NAME, MREG_REG);
      attr_err = 1'b1;
    end
    if (attr_err == 1'b1) #1 $finish;
  end
`endif
`ifdef XIL_TIMING
  reg notifier;
`endif
// begin behavioral model
  localparam M_WIDTH   = 45;
  reg [M_WIDTH-1:0] U_DATA_reg;
  reg [M_WIDTH-1:0] V_DATA_reg;
// initialize regs
`ifndef XIL_XECLIB
initial begin
  U_DATA_reg = {1'b0, {M_WIDTH-1{1'b0}}};
  V_DATA_reg = {1'b0, {M_WIDTH-1{1'b0}}};
end
`endif
   always @(posedge CLK_in) begin
      if  (RSTM_in || (MREG_BIN == 1'b0) || glblGSR) begin
         U_DATA_reg <= {1'b0, {M_WIDTH-1{1'b0}}};
         V_DATA_reg <= {1'b0, {M_WIDTH-1{1'b0}}};
      end else if (CEM_in)  begin
         U_DATA_reg <= U_in;
         V_DATA_reg <= V_in;
      end
   end
   assign U_DATA = (MREG_BIN == 1'b1) ? U_DATA_reg    : U_in;
   assign V_DATA = (MREG_BIN == 1'b1) ? V_DATA_reg    : V_in;
// end behavioral model
`ifndef XIL_XECLIB
`ifdef XIL_TIMING
  wire clk_en_n;
  wire clk_en_p;
  assign clk_en_n = IS_CLK_INVERTED_REG;
  assign clk_en_p = ~IS_CLK_INVERTED_REG;
`endif
  specify
    (CLK => U_DATA[0]) = (0:0:0, 0:0:0);
    (CLK => U_DATA[10]) = (0:0:0, 0:0:0);
    (CLK => U_DATA[11]) = (0:0:0, 0:0:0);
    (CLK => U_DATA[12]) = (0:0:0, 0:0:0);
    (CLK => U_DATA[13]) = (0:0:0, 0:0:0);
    (CLK => U_DATA[14]) = (0:0:0, 0:0:0);
    (CLK => U_DATA[15]) = (0:0:0, 0:0:0);
    (CLK => U_DATA[16]) = (0:0:0, 0:0:0);
    (CLK => U_DATA[17]) = (0:0:0, 0:0:0);
    (CLK => U_DATA[18]) = (0:0:0, 0:0:0);
    (CLK => U_DATA[19]) = (0:0:0, 0:0:0);
    (CLK => U_DATA[1]) = (0:0:0, 0:0:0);
    (CLK => U_DATA[20]) = (0:0:0, 0:0:0);
    (CLK => U_DATA[21]) = (0:0:0, 0:0:0);
    (CLK => U_DATA[22]) = (0:0:0, 0:0:0);
    (CLK => U_DATA[23]) = (0:0:0, 0:0:0);
    (CLK => U_DATA[24]) = (0:0:0, 0:0:0);
    (CLK => U_DATA[25]) = (0:0:0, 0:0:0);
    (CLK => U_DATA[26]) = (0:0:0, 0:0:0);
    (CLK => U_DATA[27]) = (0:0:0, 0:0:0);
    (CLK => U_DATA[28]) = (0:0:0, 0:0:0);
    (CLK => U_DATA[29]) = (0:0:0, 0:0:0);
    (CLK => U_DATA[2]) = (0:0:0, 0:0:0);
    (CLK => U_DATA[30]) = (0:0:0, 0:0:0);
    (CLK => U_DATA[31]) = (0:0:0, 0:0:0);
    (CLK => U_DATA[32]) = (0:0:0, 0:0:0);
    (CLK => U_DATA[33]) = (0:0:0, 0:0:0);
    (CLK => U_DATA[34]) = (0:0:0, 0:0:0);
    (CLK => U_DATA[35]) = (0:0:0, 0:0:0);
    (CLK => U_DATA[36]) = (0:0:0, 0:0:0);
    (CLK => U_DATA[37]) = (0:0:0, 0:0:0);
    (CLK => U_DATA[38]) = (0:0:0, 0:0:0);
    (CLK => U_DATA[39]) = (0:0:0, 0:0:0);
    (CLK => U_DATA[3]) = (0:0:0, 0:0:0);
    (CLK => U_DATA[40]) = (0:0:0, 0:0:0);
    (CLK => U_DATA[41]) = (0:0:0, 0:0:0);
    (CLK => U_DATA[42]) = (0:0:0, 0:0:0);
    (CLK => U_DATA[43]) = (0:0:0, 0:0:0);
    (CLK => U_DATA[44]) = (0:0:0, 0:0:0);
    (CLK => U_DATA[4]) = (0:0:0, 0:0:0);
    (CLK => U_DATA[5]) = (0:0:0, 0:0:0);
    (CLK => U_DATA[6]) = (0:0:0, 0:0:0);
    (CLK => U_DATA[7]) = (0:0:0, 0:0:0);
    (CLK => U_DATA[8]) = (0:0:0, 0:0:0);
    (CLK => U_DATA[9]) = (0:0:0, 0:0:0);
    (CLK => V_DATA[0]) = (0:0:0, 0:0:0);
    (CLK => V_DATA[10]) = (0:0:0, 0:0:0);
    (CLK => V_DATA[11]) = (0:0:0, 0:0:0);
    (CLK => V_DATA[12]) = (0:0:0, 0:0:0);
    (CLK => V_DATA[13]) = (0:0:0, 0:0:0);
    (CLK => V_DATA[14]) = (0:0:0, 0:0:0);
    (CLK => V_DATA[15]) = (0:0:0, 0:0:0);
    (CLK => V_DATA[16]) = (0:0:0, 0:0:0);
    (CLK => V_DATA[17]) = (0:0:0, 0:0:0);
    (CLK => V_DATA[18]) = (0:0:0, 0:0:0);
    (CLK => V_DATA[19]) = (0:0:0, 0:0:0);
    (CLK => V_DATA[1]) = (0:0:0, 0:0:0);
    (CLK => V_DATA[20]) = (0:0:0, 0:0:0);
    (CLK => V_DATA[21]) = (0:0:0, 0:0:0);
    (CLK => V_DATA[22]) = (0:0:0, 0:0:0);
    (CLK => V_DATA[23]) = (0:0:0, 0:0:0);
    (CLK => V_DATA[24]) = (0:0:0, 0:0:0);
    (CLK => V_DATA[25]) = (0:0:0, 0:0:0);
    (CLK => V_DATA[26]) = (0:0:0, 0:0:0);
    (CLK => V_DATA[27]) = (0:0:0, 0:0:0);
    (CLK => V_DATA[28]) = (0:0:0, 0:0:0);
    (CLK => V_DATA[29]) = (0:0:0, 0:0:0);
    (CLK => V_DATA[2]) = (0:0:0, 0:0:0);
    (CLK => V_DATA[30]) = (0:0:0, 0:0:0);
    (CLK => V_DATA[31]) = (0:0:0, 0:0:0);
    (CLK => V_DATA[32]) = (0:0:0, 0:0:0);
    (CLK => V_DATA[33]) = (0:0:0, 0:0:0);
    (CLK => V_DATA[34]) = (0:0:0, 0:0:0);
    (CLK => V_DATA[35]) = (0:0:0, 0:0:0);
    (CLK => V_DATA[36]) = (0:0:0, 0:0:0);
    (CLK => V_DATA[37]) = (0:0:0, 0:0:0);
    (CLK => V_DATA[38]) = (0:0:0, 0:0:0);
    (CLK => V_DATA[39]) = (0:0:0, 0:0:0);
    (CLK => V_DATA[3]) = (0:0:0, 0:0:0);
    (CLK => V_DATA[40]) = (0:0:0, 0:0:0);
    (CLK => V_DATA[41]) = (0:0:0, 0:0:0);
    (CLK => V_DATA[42]) = (0:0:0, 0:0:0);
    (CLK => V_DATA[43]) = (0:0:0, 0:0:0);
    (CLK => V_DATA[44]) = (0:0:0, 0:0:0);
    (CLK => V_DATA[4]) = (0:0:0, 0:0:0);
    (CLK => V_DATA[5]) = (0:0:0, 0:0:0);
    (CLK => V_DATA[6]) = (0:0:0, 0:0:0);
    (CLK => V_DATA[7]) = (0:0:0, 0:0:0);
    (CLK => V_DATA[8]) = (0:0:0, 0:0:0);
    (CLK => V_DATA[9]) = (0:0:0, 0:0:0);
    (U[0] => U_DATA[0]) = (0:0:0, 0:0:0);
    (U[10] => U_DATA[10]) = (0:0:0, 0:0:0);
    (U[11] => U_DATA[11]) = (0:0:0, 0:0:0);
    (U[12] => U_DATA[12]) = (0:0:0, 0:0:0);
    (U[13] => U_DATA[13]) = (0:0:0, 0:0:0);
    (U[14] => U_DATA[14]) = (0:0:0, 0:0:0);
    (U[15] => U_DATA[15]) = (0:0:0, 0:0:0);
    (U[16] => U_DATA[16]) = (0:0:0, 0:0:0);
    (U[17] => U_DATA[17]) = (0:0:0, 0:0:0);
    (U[18] => U_DATA[18]) = (0:0:0, 0:0:0);
    (U[19] => U_DATA[19]) = (0:0:0, 0:0:0);
    (U[1] => U_DATA[1]) = (0:0:0, 0:0:0);
    (U[20] => U_DATA[20]) = (0:0:0, 0:0:0);
    (U[21] => U_DATA[21]) = (0:0:0, 0:0:0);
    (U[22] => U_DATA[22]) = (0:0:0, 0:0:0);
    (U[23] => U_DATA[23]) = (0:0:0, 0:0:0);
    (U[24] => U_DATA[24]) = (0:0:0, 0:0:0);
    (U[25] => U_DATA[25]) = (0:0:0, 0:0:0);
    (U[26] => U_DATA[26]) = (0:0:0, 0:0:0);
    (U[27] => U_DATA[27]) = (0:0:0, 0:0:0);
    (U[28] => U_DATA[28]) = (0:0:0, 0:0:0);
    (U[29] => U_DATA[29]) = (0:0:0, 0:0:0);
    (U[2] => U_DATA[2]) = (0:0:0, 0:0:0);
    (U[30] => U_DATA[30]) = (0:0:0, 0:0:0);
    (U[31] => U_DATA[31]) = (0:0:0, 0:0:0);
    (U[32] => U_DATA[32]) = (0:0:0, 0:0:0);
    (U[33] => U_DATA[33]) = (0:0:0, 0:0:0);
    (U[34] => U_DATA[34]) = (0:0:0, 0:0:0);
    (U[35] => U_DATA[35]) = (0:0:0, 0:0:0);
    (U[36] => U_DATA[36]) = (0:0:0, 0:0:0);
    (U[37] => U_DATA[37]) = (0:0:0, 0:0:0);
    (U[38] => U_DATA[38]) = (0:0:0, 0:0:0);
    (U[39] => U_DATA[39]) = (0:0:0, 0:0:0);
    (U[3] => U_DATA[3]) = (0:0:0, 0:0:0);
    (U[40] => U_DATA[40]) = (0:0:0, 0:0:0);
    (U[41] => U_DATA[41]) = (0:0:0, 0:0:0);
    (U[42] => U_DATA[42]) = (0:0:0, 0:0:0);
    (U[43] => U_DATA[43]) = (0:0:0, 0:0:0);
    (U[4] => U_DATA[4]) = (0:0:0, 0:0:0);
    (U[5] => U_DATA[5]) = (0:0:0, 0:0:0);
    (U[6] => U_DATA[6]) = (0:0:0, 0:0:0);
    (U[7] => U_DATA[7]) = (0:0:0, 0:0:0);
    (U[8] => U_DATA[8]) = (0:0:0, 0:0:0);
    (U[9] => U_DATA[9]) = (0:0:0, 0:0:0);
    (V[0] => V_DATA[0]) = (0:0:0, 0:0:0);
    (V[10] => V_DATA[10]) = (0:0:0, 0:0:0);
    (V[11] => V_DATA[11]) = (0:0:0, 0:0:0);
    (V[12] => V_DATA[12]) = (0:0:0, 0:0:0);
    (V[13] => V_DATA[13]) = (0:0:0, 0:0:0);
    (V[14] => V_DATA[14]) = (0:0:0, 0:0:0);
    (V[15] => V_DATA[15]) = (0:0:0, 0:0:0);
    (V[16] => V_DATA[16]) = (0:0:0, 0:0:0);
    (V[17] => V_DATA[17]) = (0:0:0, 0:0:0);
    (V[18] => V_DATA[18]) = (0:0:0, 0:0:0);
    (V[19] => V_DATA[19]) = (0:0:0, 0:0:0);
    (V[20] => V_DATA[20]) = (0:0:0, 0:0:0);
    (V[21] => V_DATA[21]) = (0:0:0, 0:0:0);
    (V[22] => V_DATA[22]) = (0:0:0, 0:0:0);
    (V[23] => V_DATA[23]) = (0:0:0, 0:0:0);
    (V[24] => V_DATA[24]) = (0:0:0, 0:0:0);
    (V[25] => V_DATA[25]) = (0:0:0, 0:0:0);
    (V[26] => V_DATA[26]) = (0:0:0, 0:0:0);
    (V[27] => V_DATA[27]) = (0:0:0, 0:0:0);
    (V[28] => V_DATA[28]) = (0:0:0, 0:0:0);
    (V[29] => V_DATA[29]) = (0:0:0, 0:0:0);
    (V[30] => V_DATA[30]) = (0:0:0, 0:0:0);
    (V[31] => V_DATA[31]) = (0:0:0, 0:0:0);
    (V[32] => V_DATA[32]) = (0:0:0, 0:0:0);
    (V[33] => V_DATA[33]) = (0:0:0, 0:0:0);
    (V[34] => V_DATA[34]) = (0:0:0, 0:0:0);
    (V[35] => V_DATA[35]) = (0:0:0, 0:0:0);
    (V[36] => V_DATA[36]) = (0:0:0, 0:0:0);
    (V[37] => V_DATA[37]) = (0:0:0, 0:0:0);
    (V[38] => V_DATA[38]) = (0:0:0, 0:0:0);
    (V[39] => V_DATA[39]) = (0:0:0, 0:0:0);
    (V[40] => V_DATA[40]) = (0:0:0, 0:0:0);
    (V[41] => V_DATA[41]) = (0:0:0, 0:0:0);
    (V[42] => V_DATA[42]) = (0:0:0, 0:0:0);
    (V[43] => V_DATA[43]) = (0:0:0, 0:0:0);
    (V[4] => V_DATA[4]) = (0:0:0, 0:0:0);
    (V[5] => V_DATA[5]) = (0:0:0, 0:0:0);
    (V[6] => V_DATA[6]) = (0:0:0, 0:0:0);
    (V[7] => V_DATA[7]) = (0:0:0, 0:0:0);
    (V[8] => V_DATA[8]) = (0:0:0, 0:0:0);
    (V[9] => V_DATA[9]) = (0:0:0, 0:0:0);
`ifdef XIL_TIMING
    $setuphold (negedge CLK, negedge CEM, 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, CEM_delay);
    $setuphold (negedge CLK, negedge RSTM, 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, RSTM_delay);
    $setuphold (negedge CLK, negedge U[0], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, U_delay[0]);
    $setuphold (negedge CLK, negedge U[10], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, U_delay[10]);
    $setuphold (negedge CLK, negedge U[11], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, U_delay[11]);
    $setuphold (negedge CLK, negedge U[12], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, U_delay[12]);
    $setuphold (negedge CLK, negedge U[13], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, U_delay[13]);
    $setuphold (negedge CLK, negedge U[14], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, U_delay[14]);
    $setuphold (negedge CLK, negedge U[15], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, U_delay[15]);
    $setuphold (negedge CLK, negedge U[16], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, U_delay[16]);
    $setuphold (negedge CLK, negedge U[17], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, U_delay[17]);
    $setuphold (negedge CLK, negedge U[18], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, U_delay[18]);
    $setuphold (negedge CLK, negedge U[19], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, U_delay[19]);
    $setuphold (negedge CLK, negedge U[1], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, U_delay[1]);
    $setuphold (negedge CLK, negedge U[20], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, U_delay[20]);
    $setuphold (negedge CLK, negedge U[21], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, U_delay[21]);
    $setuphold (negedge CLK, negedge U[22], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, U_delay[22]);
    $setuphold (negedge CLK, negedge U[23], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, U_delay[23]);
    $setuphold (negedge CLK, negedge U[24], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, U_delay[24]);
    $setuphold (negedge CLK, negedge U[25], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, U_delay[25]);
    $setuphold (negedge CLK, negedge U[26], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, U_delay[26]);
    $setuphold (negedge CLK, negedge U[27], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, U_delay[27]);
    $setuphold (negedge CLK, negedge U[28], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, U_delay[28]);
    $setuphold (negedge CLK, negedge U[29], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, U_delay[29]);
    $setuphold (negedge CLK, negedge U[2], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, U_delay[2]);
    $setuphold (negedge CLK, negedge U[30], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, U_delay[30]);
    $setuphold (negedge CLK, negedge U[31], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, U_delay[31]);
    $setuphold (negedge CLK, negedge U[32], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, U_delay[32]);
    $setuphold (negedge CLK, negedge U[33], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, U_delay[33]);
    $setuphold (negedge CLK, negedge U[34], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, U_delay[34]);
    $setuphold (negedge CLK, negedge U[35], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, U_delay[35]);
    $setuphold (negedge CLK, negedge U[36], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, U_delay[36]);
    $setuphold (negedge CLK, negedge U[37], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, U_delay[37]);
    $setuphold (negedge CLK, negedge U[38], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, U_delay[38]);
    $setuphold (negedge CLK, negedge U[39], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, U_delay[39]);
    $setuphold (negedge CLK, negedge U[3], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, U_delay[3]);
    $setuphold (negedge CLK, negedge U[40], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, U_delay[40]);
    $setuphold (negedge CLK, negedge U[41], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, U_delay[41]);
    $setuphold (negedge CLK, negedge U[42], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, U_delay[42]);
    $setuphold (negedge CLK, negedge U[43], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, U_delay[43]);
    $setuphold (negedge CLK, negedge U[4], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, U_delay[4]);
    $setuphold (negedge CLK, negedge U[5], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, U_delay[5]);
    $setuphold (negedge CLK, negedge U[6], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, U_delay[6]);
    $setuphold (negedge CLK, negedge U[7], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, U_delay[7]);
    $setuphold (negedge CLK, negedge U[8], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, U_delay[8]);
    $setuphold (negedge CLK, negedge U[9], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, U_delay[9]);
    $setuphold (negedge CLK, negedge V[0], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, V_delay[0]);
    $setuphold (negedge CLK, negedge V[10], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, V_delay[10]);
    $setuphold (negedge CLK, negedge V[11], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, V_delay[11]);
    $setuphold (negedge CLK, negedge V[12], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, V_delay[12]);
    $setuphold (negedge CLK, negedge V[13], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, V_delay[13]);
    $setuphold (negedge CLK, negedge V[14], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, V_delay[14]);
    $setuphold (negedge CLK, negedge V[15], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, V_delay[15]);
    $setuphold (negedge CLK, negedge V[16], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, V_delay[16]);
    $setuphold (negedge CLK, negedge V[17], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, V_delay[17]);
    $setuphold (negedge CLK, negedge V[18], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, V_delay[18]);
    $setuphold (negedge CLK, negedge V[19], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, V_delay[19]);
    $setuphold (negedge CLK, negedge V[20], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, V_delay[20]);
    $setuphold (negedge CLK, negedge V[21], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, V_delay[21]);
    $setuphold (negedge CLK, negedge V[22], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, V_delay[22]);
    $setuphold (negedge CLK, negedge V[23], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, V_delay[23]);
    $setuphold (negedge CLK, negedge V[24], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, V_delay[24]);
    $setuphold (negedge CLK, negedge V[25], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, V_delay[25]);
    $setuphold (negedge CLK, negedge V[26], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, V_delay[26]);
    $setuphold (negedge CLK, negedge V[27], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, V_delay[27]);
    $setuphold (negedge CLK, negedge V[28], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, V_delay[28]);
    $setuphold (negedge CLK, negedge V[29], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, V_delay[29]);
    $setuphold (negedge CLK, negedge V[30], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, V_delay[30]);
    $setuphold (negedge CLK, negedge V[31], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, V_delay[31]);
    $setuphold (negedge CLK, negedge V[32], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, V_delay[32]);
    $setuphold (negedge CLK, negedge V[33], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, V_delay[33]);
    $setuphold (negedge CLK, negedge V[34], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, V_delay[34]);
    $setuphold (negedge CLK, negedge V[35], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, V_delay[35]);
    $setuphold (negedge CLK, negedge V[36], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, V_delay[36]);
    $setuphold (negedge CLK, negedge V[37], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, V_delay[37]);
    $setuphold (negedge CLK, negedge V[38], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, V_delay[38]);
    $setuphold (negedge CLK, negedge V[39], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, V_delay[39]);
    $setuphold (negedge CLK, negedge V[40], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, V_delay[40]);
    $setuphold (negedge CLK, negedge V[41], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, V_delay[41]);
    $setuphold (negedge CLK, negedge V[42], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, V_delay[42]);
    $setuphold (negedge CLK, negedge V[43], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, V_delay[43]);
    $setuphold (negedge CLK, negedge V[4], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, V_delay[4]);
    $setuphold (negedge CLK, negedge V[5], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, V_delay[5]);
    $setuphold (negedge CLK, negedge V[6], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, V_delay[6]);
    $setuphold (negedge CLK, negedge V[7], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, V_delay[7]);
    $setuphold (negedge CLK, negedge V[8], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, V_delay[8]);
    $setuphold (negedge CLK, negedge V[9], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, V_delay[9]);
    $setuphold (negedge CLK, posedge CEM, 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, CEM_delay);
    $setuphold (negedge CLK, posedge RSTM, 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, RSTM_delay);
    $setuphold (negedge CLK, posedge U[0], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, U_delay[0]);
    $setuphold (negedge CLK, posedge U[10], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, U_delay[10]);
    $setuphold (negedge CLK, posedge U[11], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, U_delay[11]);
    $setuphold (negedge CLK, posedge U[12], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, U_delay[12]);
    $setuphold (negedge CLK, posedge U[13], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, U_delay[13]);
    $setuphold (negedge CLK, posedge U[14], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, U_delay[14]);
    $setuphold (negedge CLK, posedge U[15], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, U_delay[15]);
    $setuphold (negedge CLK, posedge U[16], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, U_delay[16]);
    $setuphold (negedge CLK, posedge U[17], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, U_delay[17]);
    $setuphold (negedge CLK, posedge U[18], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, U_delay[18]);
    $setuphold (negedge CLK, posedge U[19], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, U_delay[19]);
    $setuphold (negedge CLK, posedge U[1], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, U_delay[1]);
    $setuphold (negedge CLK, posedge U[20], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, U_delay[20]);
    $setuphold (negedge CLK, posedge U[21], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, U_delay[21]);
    $setuphold (negedge CLK, posedge U[22], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, U_delay[22]);
    $setuphold (negedge CLK, posedge U[23], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, U_delay[23]);
    $setuphold (negedge CLK, posedge U[24], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, U_delay[24]);
    $setuphold (negedge CLK, posedge U[25], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, U_delay[25]);
    $setuphold (negedge CLK, posedge U[26], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, U_delay[26]);
    $setuphold (negedge CLK, posedge U[27], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, U_delay[27]);
    $setuphold (negedge CLK, posedge U[28], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, U_delay[28]);
    $setuphold (negedge CLK, posedge U[29], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, U_delay[29]);
    $setuphold (negedge CLK, posedge U[2], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, U_delay[2]);
    $setuphold (negedge CLK, posedge U[30], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, U_delay[30]);
    $setuphold (negedge CLK, posedge U[31], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, U_delay[31]);
    $setuphold (negedge CLK, posedge U[32], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, U_delay[32]);
    $setuphold (negedge CLK, posedge U[33], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, U_delay[33]);
    $setuphold (negedge CLK, posedge U[34], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, U_delay[34]);
    $setuphold (negedge CLK, posedge U[35], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, U_delay[35]);
    $setuphold (negedge CLK, posedge U[36], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, U_delay[36]);
    $setuphold (negedge CLK, posedge U[37], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, U_delay[37]);
    $setuphold (negedge CLK, posedge U[38], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, U_delay[38]);
    $setuphold (negedge CLK, posedge U[39], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, U_delay[39]);
    $setuphold (negedge CLK, posedge U[3], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, U_delay[3]);
    $setuphold (negedge CLK, posedge U[40], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, U_delay[40]);
    $setuphold (negedge CLK, posedge U[41], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, U_delay[41]);
    $setuphold (negedge CLK, posedge U[42], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, U_delay[42]);
    $setuphold (negedge CLK, posedge U[43], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, U_delay[43]);
    $setuphold (negedge CLK, posedge U[4], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, U_delay[4]);
    $setuphold (negedge CLK, posedge U[5], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, U_delay[5]);
    $setuphold (negedge CLK, posedge U[6], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, U_delay[6]);
    $setuphold (negedge CLK, posedge U[7], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, U_delay[7]);
    $setuphold (negedge CLK, posedge U[8], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, U_delay[8]);
    $setuphold (negedge CLK, posedge U[9], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, U_delay[9]);
    $setuphold (negedge CLK, posedge V[0], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, V_delay[0]);
    $setuphold (negedge CLK, posedge V[10], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, V_delay[10]);
    $setuphold (negedge CLK, posedge V[11], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, V_delay[11]);
    $setuphold (negedge CLK, posedge V[12], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, V_delay[12]);
    $setuphold (negedge CLK, posedge V[13], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, V_delay[13]);
    $setuphold (negedge CLK, posedge V[14], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, V_delay[14]);
    $setuphold (negedge CLK, posedge V[15], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, V_delay[15]);
    $setuphold (negedge CLK, posedge V[16], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, V_delay[16]);
    $setuphold (negedge CLK, posedge V[17], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, V_delay[17]);
    $setuphold (negedge CLK, posedge V[18], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, V_delay[18]);
    $setuphold (negedge CLK, posedge V[19], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, V_delay[19]);
    $setuphold (negedge CLK, posedge V[20], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, V_delay[20]);
    $setuphold (negedge CLK, posedge V[21], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, V_delay[21]);
    $setuphold (negedge CLK, posedge V[22], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, V_delay[22]);
    $setuphold (negedge CLK, posedge V[23], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, V_delay[23]);
    $setuphold (negedge CLK, posedge V[24], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, V_delay[24]);
    $setuphold (negedge CLK, posedge V[25], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, V_delay[25]);
    $setuphold (negedge CLK, posedge V[26], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, V_delay[26]);
    $setuphold (negedge CLK, posedge V[27], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, V_delay[27]);
    $setuphold (negedge CLK, posedge V[28], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, V_delay[28]);
    $setuphold (negedge CLK, posedge V[29], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, V_delay[29]);
    $setuphold (negedge CLK, posedge V[30], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, V_delay[30]);
    $setuphold (negedge CLK, posedge V[31], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, V_delay[31]);
    $setuphold (negedge CLK, posedge V[32], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, V_delay[32]);
    $setuphold (negedge CLK, posedge V[33], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, V_delay[33]);
    $setuphold (negedge CLK, posedge V[34], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, V_delay[34]);
    $setuphold (negedge CLK, posedge V[35], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, V_delay[35]);
    $setuphold (negedge CLK, posedge V[36], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, V_delay[36]);
    $setuphold (negedge CLK, posedge V[37], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, V_delay[37]);
    $setuphold (negedge CLK, posedge V[38], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, V_delay[38]);
    $setuphold (negedge CLK, posedge V[39], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, V_delay[39]);
    $setuphold (negedge CLK, posedge V[40], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, V_delay[40]);
    $setuphold (negedge CLK, posedge V[41], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, V_delay[41]);
    $setuphold (negedge CLK, posedge V[42], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, V_delay[42]);
    $setuphold (negedge CLK, posedge V[43], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, V_delay[43]);
    $setuphold (negedge CLK, posedge V[4], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, V_delay[4]);
    $setuphold (negedge CLK, posedge V[5], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, V_delay[5]);
    $setuphold (negedge CLK, posedge V[6], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, V_delay[6]);
    $setuphold (negedge CLK, posedge V[7], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, V_delay[7]);
    $setuphold (negedge CLK, posedge V[8], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, V_delay[8]);
    $setuphold (negedge CLK, posedge V[9], 0:0:0, 0:0:0, notifier, clk_en_n, clk_en_n, CLK_delay, V_delay[9]);
    $setuphold (posedge CLK, negedge CEM, 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, CEM_delay);
    $setuphold (posedge CLK, negedge RSTM, 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, RSTM_delay);
    $setuphold (posedge CLK, negedge U[0], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, U_delay[0]);
    $setuphold (posedge CLK, negedge U[10], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, U_delay[10]);
    $setuphold (posedge CLK, negedge U[11], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, U_delay[11]);
    $setuphold (posedge CLK, negedge U[12], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, U_delay[12]);
    $setuphold (posedge CLK, negedge U[13], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, U_delay[13]);
    $setuphold (posedge CLK, negedge U[14], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, U_delay[14]);
    $setuphold (posedge CLK, negedge U[15], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, U_delay[15]);
    $setuphold (posedge CLK, negedge U[16], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, U_delay[16]);
    $setuphold (posedge CLK, negedge U[17], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, U_delay[17]);
    $setuphold (posedge CLK, negedge U[18], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, U_delay[18]);
    $setuphold (posedge CLK, negedge U[19], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, U_delay[19]);
    $setuphold (posedge CLK, negedge U[1], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, U_delay[1]);
    $setuphold (posedge CLK, negedge U[20], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, U_delay[20]);
    $setuphold (posedge CLK, negedge U[21], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, U_delay[21]);
    $setuphold (posedge CLK, negedge U[22], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, U_delay[22]);
    $setuphold (posedge CLK, negedge U[23], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, U_delay[23]);
    $setuphold (posedge CLK, negedge U[24], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, U_delay[24]);
    $setuphold (posedge CLK, negedge U[25], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, U_delay[25]);
    $setuphold (posedge CLK, negedge U[26], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, U_delay[26]);
    $setuphold (posedge CLK, negedge U[27], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, U_delay[27]);
    $setuphold (posedge CLK, negedge U[28], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, U_delay[28]);
    $setuphold (posedge CLK, negedge U[29], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, U_delay[29]);
    $setuphold (posedge CLK, negedge U[2], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, U_delay[2]);
    $setuphold (posedge CLK, negedge U[30], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, U_delay[30]);
    $setuphold (posedge CLK, negedge U[31], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, U_delay[31]);
    $setuphold (posedge CLK, negedge U[32], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, U_delay[32]);
    $setuphold (posedge CLK, negedge U[33], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, U_delay[33]);
    $setuphold (posedge CLK, negedge U[34], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, U_delay[34]);
    $setuphold (posedge CLK, negedge U[35], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, U_delay[35]);
    $setuphold (posedge CLK, negedge U[36], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, U_delay[36]);
    $setuphold (posedge CLK, negedge U[37], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, U_delay[37]);
    $setuphold (posedge CLK, negedge U[38], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, U_delay[38]);
    $setuphold (posedge CLK, negedge U[39], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, U_delay[39]);
    $setuphold (posedge CLK, negedge U[3], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, U_delay[3]);
    $setuphold (posedge CLK, negedge U[40], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, U_delay[40]);
    $setuphold (posedge CLK, negedge U[41], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, U_delay[41]);
    $setuphold (posedge CLK, negedge U[42], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, U_delay[42]);
    $setuphold (posedge CLK, negedge U[43], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, U_delay[43]);
    $setuphold (posedge CLK, negedge U[4], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, U_delay[4]);
    $setuphold (posedge CLK, negedge U[5], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, U_delay[5]);
    $setuphold (posedge CLK, negedge U[6], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, U_delay[6]);
    $setuphold (posedge CLK, negedge U[7], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, U_delay[7]);
    $setuphold (posedge CLK, negedge U[8], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, U_delay[8]);
    $setuphold (posedge CLK, negedge U[9], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, U_delay[9]);
    $setuphold (posedge CLK, negedge V[0], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, V_delay[0]);
    $setuphold (posedge CLK, negedge V[10], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, V_delay[10]);
    $setuphold (posedge CLK, negedge V[11], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, V_delay[11]);
    $setuphold (posedge CLK, negedge V[12], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, V_delay[12]);
    $setuphold (posedge CLK, negedge V[13], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, V_delay[13]);
    $setuphold (posedge CLK, negedge V[14], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, V_delay[14]);
    $setuphold (posedge CLK, negedge V[15], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, V_delay[15]);
    $setuphold (posedge CLK, negedge V[16], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, V_delay[16]);
    $setuphold (posedge CLK, negedge V[17], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, V_delay[17]);
    $setuphold (posedge CLK, negedge V[18], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, V_delay[18]);
    $setuphold (posedge CLK, negedge V[19], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, V_delay[19]);
    $setuphold (posedge CLK, negedge V[20], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, V_delay[20]);
    $setuphold (posedge CLK, negedge V[21], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, V_delay[21]);
    $setuphold (posedge CLK, negedge V[22], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, V_delay[22]);
    $setuphold (posedge CLK, negedge V[23], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, V_delay[23]);
    $setuphold (posedge CLK, negedge V[24], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, V_delay[24]);
    $setuphold (posedge CLK, negedge V[25], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, V_delay[25]);
    $setuphold (posedge CLK, negedge V[26], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, V_delay[26]);
    $setuphold (posedge CLK, negedge V[27], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, V_delay[27]);
    $setuphold (posedge CLK, negedge V[28], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, V_delay[28]);
    $setuphold (posedge CLK, negedge V[29], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, V_delay[29]);
    $setuphold (posedge CLK, negedge V[30], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, V_delay[30]);
    $setuphold (posedge CLK, negedge V[31], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, V_delay[31]);
    $setuphold (posedge CLK, negedge V[32], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, V_delay[32]);
    $setuphold (posedge CLK, negedge V[33], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, V_delay[33]);
    $setuphold (posedge CLK, negedge V[34], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, V_delay[34]);
    $setuphold (posedge CLK, negedge V[35], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, V_delay[35]);
    $setuphold (posedge CLK, negedge V[36], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, V_delay[36]);
    $setuphold (posedge CLK, negedge V[37], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, V_delay[37]);
    $setuphold (posedge CLK, negedge V[38], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, V_delay[38]);
    $setuphold (posedge CLK, negedge V[39], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, V_delay[39]);
    $setuphold (posedge CLK, negedge V[40], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, V_delay[40]);
    $setuphold (posedge CLK, negedge V[41], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, V_delay[41]);
    $setuphold (posedge CLK, negedge V[42], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, V_delay[42]);
    $setuphold (posedge CLK, negedge V[43], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, V_delay[43]);
    $setuphold (posedge CLK, negedge V[4], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, V_delay[4]);
    $setuphold (posedge CLK, negedge V[5], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, V_delay[5]);
    $setuphold (posedge CLK, negedge V[6], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, V_delay[6]);
    $setuphold (posedge CLK, negedge V[7], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, V_delay[7]);
    $setuphold (posedge CLK, negedge V[8], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, V_delay[8]);
    $setuphold (posedge CLK, negedge V[9], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, V_delay[9]);
    $setuphold (posedge CLK, posedge CEM, 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, CEM_delay);
    $setuphold (posedge CLK, posedge RSTM, 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, RSTM_delay);
    $setuphold (posedge CLK, posedge U[0], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, U_delay[0]);
    $setuphold (posedge CLK, posedge U[10], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, U_delay[10]);
    $setuphold (posedge CLK, posedge U[11], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, U_delay[11]);
    $setuphold (posedge CLK, posedge U[12], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, U_delay[12]);
    $setuphold (posedge CLK, posedge U[13], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, U_delay[13]);
    $setuphold (posedge CLK, posedge U[14], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, U_delay[14]);
    $setuphold (posedge CLK, posedge U[15], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, U_delay[15]);
    $setuphold (posedge CLK, posedge U[16], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, U_delay[16]);
    $setuphold (posedge CLK, posedge U[17], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, U_delay[17]);
    $setuphold (posedge CLK, posedge U[18], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, U_delay[18]);
    $setuphold (posedge CLK, posedge U[19], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, U_delay[19]);
    $setuphold (posedge CLK, posedge U[1], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, U_delay[1]);
    $setuphold (posedge CLK, posedge U[20], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, U_delay[20]);
    $setuphold (posedge CLK, posedge U[21], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, U_delay[21]);
    $setuphold (posedge CLK, posedge U[22], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, U_delay[22]);
    $setuphold (posedge CLK, posedge U[23], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, U_delay[23]);
    $setuphold (posedge CLK, posedge U[24], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, U_delay[24]);
    $setuphold (posedge CLK, posedge U[25], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, U_delay[25]);
    $setuphold (posedge CLK, posedge U[26], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, U_delay[26]);
    $setuphold (posedge CLK, posedge U[27], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, U_delay[27]);
    $setuphold (posedge CLK, posedge U[28], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, U_delay[28]);
    $setuphold (posedge CLK, posedge U[29], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, U_delay[29]);
    $setuphold (posedge CLK, posedge U[2], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, U_delay[2]);
    $setuphold (posedge CLK, posedge U[30], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, U_delay[30]);
    $setuphold (posedge CLK, posedge U[31], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, U_delay[31]);
    $setuphold (posedge CLK, posedge U[32], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, U_delay[32]);
    $setuphold (posedge CLK, posedge U[33], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, U_delay[33]);
    $setuphold (posedge CLK, posedge U[34], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, U_delay[34]);
    $setuphold (posedge CLK, posedge U[35], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, U_delay[35]);
    $setuphold (posedge CLK, posedge U[36], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, U_delay[36]);
    $setuphold (posedge CLK, posedge U[37], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, U_delay[37]);
    $setuphold (posedge CLK, posedge U[38], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, U_delay[38]);
    $setuphold (posedge CLK, posedge U[39], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, U_delay[39]);
    $setuphold (posedge CLK, posedge U[3], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, U_delay[3]);
    $setuphold (posedge CLK, posedge U[40], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, U_delay[40]);
    $setuphold (posedge CLK, posedge U[41], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, U_delay[41]);
    $setuphold (posedge CLK, posedge U[42], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, U_delay[42]);
    $setuphold (posedge CLK, posedge U[43], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, U_delay[43]);
    $setuphold (posedge CLK, posedge U[4], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, U_delay[4]);
    $setuphold (posedge CLK, posedge U[5], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, U_delay[5]);
    $setuphold (posedge CLK, posedge U[6], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, U_delay[6]);
    $setuphold (posedge CLK, posedge U[7], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, U_delay[7]);
    $setuphold (posedge CLK, posedge U[8], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, U_delay[8]);
    $setuphold (posedge CLK, posedge U[9], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, U_delay[9]);
    $setuphold (posedge CLK, posedge V[0], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, V_delay[0]);
    $setuphold (posedge CLK, posedge V[10], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, V_delay[10]);
    $setuphold (posedge CLK, posedge V[11], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, V_delay[11]);
    $setuphold (posedge CLK, posedge V[12], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, V_delay[12]);
    $setuphold (posedge CLK, posedge V[13], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, V_delay[13]);
    $setuphold (posedge CLK, posedge V[14], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, V_delay[14]);
    $setuphold (posedge CLK, posedge V[15], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, V_delay[15]);
    $setuphold (posedge CLK, posedge V[16], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, V_delay[16]);
    $setuphold (posedge CLK, posedge V[17], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, V_delay[17]);
    $setuphold (posedge CLK, posedge V[18], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, V_delay[18]);
    $setuphold (posedge CLK, posedge V[19], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, V_delay[19]);
    $setuphold (posedge CLK, posedge V[20], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, V_delay[20]);
    $setuphold (posedge CLK, posedge V[21], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, V_delay[21]);
    $setuphold (posedge CLK, posedge V[22], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, V_delay[22]);
    $setuphold (posedge CLK, posedge V[23], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, V_delay[23]);
    $setuphold (posedge CLK, posedge V[24], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, V_delay[24]);
    $setuphold (posedge CLK, posedge V[25], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, V_delay[25]);
    $setuphold (posedge CLK, posedge V[26], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, V_delay[26]);
    $setuphold (posedge CLK, posedge V[27], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, V_delay[27]);
    $setuphold (posedge CLK, posedge V[28], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, V_delay[28]);
    $setuphold (posedge CLK, posedge V[29], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, V_delay[29]);
    $setuphold (posedge CLK, posedge V[30], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, V_delay[30]);
    $setuphold (posedge CLK, posedge V[31], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, V_delay[31]);
    $setuphold (posedge CLK, posedge V[32], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, V_delay[32]);
    $setuphold (posedge CLK, posedge V[33], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, V_delay[33]);
    $setuphold (posedge CLK, posedge V[34], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, V_delay[34]);
    $setuphold (posedge CLK, posedge V[35], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, V_delay[35]);
    $setuphold (posedge CLK, posedge V[36], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, V_delay[36]);
    $setuphold (posedge CLK, posedge V[37], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, V_delay[37]);
    $setuphold (posedge CLK, posedge V[38], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, V_delay[38]);
    $setuphold (posedge CLK, posedge V[39], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, V_delay[39]);
    $setuphold (posedge CLK, posedge V[40], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, V_delay[40]);
    $setuphold (posedge CLK, posedge V[41], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, V_delay[41]);
    $setuphold (posedge CLK, posedge V[42], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, V_delay[42]);
    $setuphold (posedge CLK, posedge V[43], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, V_delay[43]);
    $setuphold (posedge CLK, posedge V[4], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, V_delay[4]);
    $setuphold (posedge CLK, posedge V[5], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, V_delay[5]);
    $setuphold (posedge CLK, posedge V[6], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, V_delay[6]);
    $setuphold (posedge CLK, posedge V[7], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, V_delay[7]);
    $setuphold (posedge CLK, posedge V[8], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, V_delay[8]);
    $setuphold (posedge CLK, posedge V[9], 0:0:0, 0:0:0, notifier, clk_en_p, clk_en_p, CLK_delay, V_delay[9]);
`endif
    specparam PATHPULSE$ = 0;
  endspecify
`endif
endmodule