module s12;
 final begin
    $write("*-* All Finished *-*\n");
 end
endmodule