module bug810 #(
		/*parameter*/ int unsigned DW = 32);
endmodule