module bug815 (
	       test_if bad[2]);
endmodule