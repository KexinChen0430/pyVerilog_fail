module header
	// Internal signals
	// Generated Signal List
	// End of Generated Signal List
	// %COMPILER_OPTS%
	// Generated Signal Assignments
	// Generated Instances and Port Mappings
		// Generated Instance Port Map for inst_eba
		inst_eba_e inst_eba (
		);
		// End of Generated Instance Port Map for inst_eba
		// Generated Instance Port Map for inst_ebb
		inst_ebb_e inst_ebb (
		);
		// End of Generated Instance Port Map for inst_ebb
		// Generated Instance Port Map for inst_ebc
		inst_ebc_e inst_ebc (
		);
		// End of Generated Instance Port Map for inst_ebc
endmodule