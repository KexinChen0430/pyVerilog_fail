module  ng8cf0c(
   sys_clk,
   rst_n,
   pse18cc,
   jrc662,
   zk63316,
   lf198b2,
   yxcc596,
   os62cb4,
   fp165a1,
   xyb2d0e,
   ba96872,
   wlb4393,
   uxa1c9c,
   vke4e4,
   ay5cd66,
   `ifdef EN_VC0
      hq93919,
      ri9c8cb,
      tue465a,
   `endif
   `ifdef EN_VC1
      sj232d3,
      hd1969c,
      uicb4e7,
   `endif
   `ifdef EN_VC2
      pf5a739,
      end39ce,
      tw9ce75,
   `endif
   `ifdef EN_VC3
      kde73aa,
      ux39d54,
      kqceaa5,
   `endif
   `ifdef EN_VC4
      ip75528,
      ntaa944,
      al54a27,
   `endif
   `ifdef EN_VC5
      lfa513c,
      hd289e7,
      al44f3e,
   `endif
   `ifdef EN_VC6
      hd279f5,
      an3cfaf,
      ipe7d7d,
   `endif
   `ifdef EN_VC7
      gq3ebed,
      ykf5f68,
      phafb41,
   `endif
   os7da0f,
   qted079,
   ww683cd,
   tx_vsd_data,
   yx4e2a2,
   al7fcee,
   xw69c54,
   jce1a71,
   zx74783,
   qia3c1e,
   tw1e0f1,
   icf078a,
   ls83c50,
   ls1e282,
   wlb4ebf,
   xya75fd,
   lqe4a1a,
   ba250d2,
   an3c4c4,
   ene2624,
   mec4930,
   jpd27c8,
   do93e46,
   mt9f233,
   xjc264f,
   jr1327f,
   cm46737,
   sj23425,
   ec1a12c,
   tud0960,
   hd84b02,
   gqb98bf
   );
`ifdef LW1
parameter LANE_WIDTH = 1 ;
`else
`ifdef LW2
parameter LANE_WIDTH = 2 ;
`else
`ifdef LW4
parameter LANE_WIDTH = 4 ;
`else
parameter LANE_WIDTH = 1 ;
`endif
`endif
`endif
parameter D_WIDTH = 16 ;
parameter K27_7 = 8'hFB ;
parameter K28_0 = 8'h1C ;
parameter K28_2 = 8'h5C ;
parameter K28_3 = 8'h7C ;
parameter K28_5 = 8'hBC ;
parameter K29_7 = 8'hFD ;
parameter K30_7 = 8'hFE ;
parameter K23_7 = 8'hF7 ;
parameter K28_1 = 8'h3C ;
parameter D5_2  = 8'h45 ;
parameter D10_2 = 8'h4A ;
parameter D21_5 = 8'hB5 ;
parameter D26_5 = 8'hBA ;
parameter COM = K28_5 ;
parameter STP = K27_7 ;
parameter SDP = K28_2 ;
parameter END = K29_7 ;
parameter EDB = K30_7 ;
parameter SKP = K28_0 ;
parameter IDL = K28_3 ;
parameter PAD = K23_7 ;
parameter FTS = K28_1 ;
parameter OS_WIDTH      = 4 ;
parameter OS_T1_LIP_LAP = 4'd0 ;
parameter OS_T2_LIP_LAP = 4'd1 ;
parameter OS_COMPLI     = 4'd2 ;
parameter OS_T1         = 4'd3 ;
parameter OS_T2         = 4'd4 ;
parameter OS_IDLE       = 4'd5 ;
parameter OS_EIDLE      = 4'd6 ;
parameter OS_NFTS       = 4'd7 ;
parameter OS_BEACON     = 4'd8 ;
parameter DSM_WIDTH    = 2 ;
parameter PSM_WIDTH    = 2 ;
parameter RSM_WIDTH    = 2 ;
parameter L0SM_WIDTH   = 2 ;
parameter L0sTSM_WIDTH = 2 ;
parameter L0sRSM_WIDTH = 2 ;
parameter L1SM_WIDTH   = 1 ;
parameter L2SM_WIDTH   = 1 ;
parameter DISM_WIDTH   = 2 ;
parameter LBSM_WIDTH   = 2 ;
parameter HRSM_WIDTH   = 1 ;
parameter CFGSM_WIDTH  = 2 ;
parameter MSM_WIDTH    = 3 ;
parameter DETECT    = 4'd0 ;
parameter POLLING   = 4'd1 ;
parameter CONFIG    = 4'd2 ;
parameter L0        = 4'd3 ;
parameter L0s       = 4'd4 ;
parameter L1        = 4'd5 ;
parameter L2        = 4'd6 ;
parameter RECOVERY  = 4'd7 ;
parameter LOOPBACK  = 4'd8 ;
parameter HOTRST    = 4'd9 ;
parameter DISABLED  = 4'd10 ;
`ifdef VC1
parameter FADDR = 3 ;
`else
`ifdef VC2
parameter FADDR = 3 ;
`else
`ifdef VC3
parameter FADDR = 5 ;
`else
`ifdef VC4
parameter FADDR = 5 ;
`else
parameter FADDR = 6 ;
`endif
`endif
`endif
`endif
`ifdef VC1
parameter  wjcc96b=2;
parameter  fn64b5d=7;
parameter  fc25aee       =  3'b011;
parameter  hd2d772  =  3'b111;
parameter  fn6bb97     =  3'b000;
parameter  ne5dcbf    =  3'b001;
parameter  neee5fa   =  3'b010;
`else
`ifdef VC2
parameter  wjcc96b=2;
parameter  fn64b5d=7;
parameter  fc25aee       =  3'b011;
parameter  hd2d772  =  3'b111;
parameter  fn6bb97     =  3'b000;
parameter  ne5dcbf    =  3'b001;
parameter  neee5fa   =  3'b010;
parameter  ksf3af     =  3'b100;
parameter  lq79d79    =  3'b101;
parameter  qgcebcb   =  3'b110;
`else
`ifdef VC3
parameter  wjcc96b=3;
parameter  fn64b5d=15;
parameter  fc25aee       =  4'b0011;
parameter  hd2d772  =  4'b1111;
parameter  fn6bb97     =  4'b0000;
parameter  ne5dcbf    =  4'b0001;
parameter  neee5fa   =  4'b0010;
parameter  ksf3af     =  4'b0100;
parameter  lq79d79    =  4'b0101;
parameter  qgcebcb   =  4'b0110;
parameter  ea5307d     =  4'b1000;
parameter  ou983e8    =  4'b1001;
parameter  ykc1f41   =  4'b1010;
`else
`ifdef VC4
parameter  wjcc96b=3;
parameter  fn64b5d=15;
parameter  fc25aee       =  4'b0011;
parameter  hd2d772  =  4'b1111;
parameter  fn6bb97     =  4'b0000;
parameter  ne5dcbf    =  4'b0001;
parameter  neee5fa   =  4'b0010;
parameter  ksf3af     =  4'b0100;
parameter  lq79d79    =  4'b0101;
parameter  qgcebcb   =  4'b0110;
parameter  ea5307d     =  4'b1000;
parameter  ou983e8    =  4'b1001;
parameter  ykc1f41   =  4'b1010;
parameter  shcc581     =  4'b1100;
parameter  su62c0c    =  4'b1101;
parameter  lf16061   =  4'b1110;
`else
parameter  wjcc96b=4;
parameter  fn64b5d=31;
parameter  fc25aee       =  5'b00011;
parameter  hd2d772  =  5'b11111;
parameter  fn6bb97     =  5'b00000;
parameter  ne5dcbf    =  5'b00001;
parameter  neee5fa   =  5'b00010;
parameter  ksf3af     =  5'b00100;
parameter  lq79d79    =  5'b00101;
parameter  qgcebcb   =  5'b00110;
parameter  ea5307d     =  5'b01000;
parameter  ou983e8    =  5'b01001;
parameter  ykc1f41   =  5'b01010;
parameter  shcc581     =  5'b01100;
parameter  su62c0c    =  5'b01101;
parameter  lf16061   =  5'b01110;
parameter  uic1c8f     =  5'b10000;
parameter  jee479    =  5'b10001;
parameter  cm723cb   =  5'b10010;
parameter  vx91e59     =  5'b10100;
parameter  wl8f2ce    =  5'b10101;
parameter  dm79675   =  5'b10110;
parameter  aycb3aa     =  5'b11000;
parameter  ic59d51    =  5'b11001;
parameter  ykcea88   =  5'b11010;
parameter  qt75440     =  5'b11100;
parameter  zzaa204    =  5'b11101;
parameter  of51026   =  5'b11110;
`endif
`endif
`endif
`endif
parameter uvc3724   = 2'b00;
parameter je1b925  = 2'b01;
parameter mrdc92b = 2'b10;
input                     sys_clk;
input                     rst_n;
input  [13:0]             pse18cc;
input                     jrc662;
input                     zk63316;
input                     lf198b2;
input  [2:0]              yxcc596;
input  [1:0]              os62cb4;
input                     fp165a1;
input  [2:0]              xyb2d0e;
input  [1:0]              ba96872;
input  [`NUM_VC -1:0]     wlb4393;
input  [`NUM_VC -1:0]     uxa1c9c;
input  [`NUM_VC -1:0]     vke4e4;
input [(`NUM_VC*3)-1:0]   ay5cd66;
`ifdef EN_VC0
input  [23:0]             hq93919;
input  [23:0]             ri9c8cb;
input  [23:0]             tue465a;
`endif
`ifdef EN_VC1
input  [23:0]             sj232d3;
input  [23:0]             hd1969c;
input  [23:0]             uicb4e7;
`endif
`ifdef EN_VC2
input  [23:0]             pf5a739;
input  [23:0]             end39ce;
input  [23:0]             tw9ce75;
`endif
`ifdef EN_VC3
input  [23:0]             kde73aa;
input  [23:0]             ux39d54;
input  [23:0]             kqceaa5;
`endif
`ifdef EN_VC4
input  [23:0]             ip75528;
input  [23:0]             ntaa944;
input  [23:0]             al54a27;
`endif
`ifdef EN_VC5
input  [23:0]             lfa513c;
input  [23:0]             hd289e7;
input  [23:0]             al44f3e;
`endif
`ifdef EN_VC6
input  [23:0]             hd279f5;
input  [23:0]             an3cfaf;
input  [23:0]             ipe7d7d;
`endif
`ifdef EN_VC7
input  [23:0]             gq3ebed;
input  [23:0]             ykf5f68;
input  [23:0]             phafb41;
`endif
input                     os7da0f;
input                     ww683cd;
input  [2:0]              qted079;
input  [23:0]             tx_vsd_data;
input                     yx4e2a2;
input                     al7fcee;
input                     xw69c54;
input  [11:0]             jce1a71;
input                     zx74783;
input                     qia3c1e;
input  [2:0]              tw1e0f1;
input                     icf078a;
input  [1:0]              ls83c50;
input  [`NUM_VC -1:0]     ls1e282;
input                     wlb4ebf;
input                     xya75fd;
input                     lqe4a1a;
output [FADDR:0]          ba250d2;
output                    an3c4c4;
output                    ene2624;
output [3:0]              mec4930;
output [`NUM_VC -1:0]     jpd27c8;
output [`NUM_VC -1:0]     do93e46;
output [`NUM_VC -1:0]     mt9f233;
output                    xjc264f;
output                    jr1327f;
output                    cm46737;
output                    sj23425;
output                    ec1a12c;
output [31:0]             tud0960;
output [31:0]             hd84b02;
output                    gqb98bf;
reg    [FADDR:0]          ba250d2;
reg                       an3c4c4;
reg                       ene2624;
reg    [3:0]              mec4930;
reg    [`NUM_VC -1:0]     jpd27c8;
reg    [`NUM_VC -1:0]     do93e46;
reg    [`NUM_VC -1:0]     mt9f233;
reg                       xjc264f;
reg                       jr1327f;
wire                      cm46737;
reg                       ec1a12c;
reg                       vi42b97;
reg                       gqb98bf;
reg                       sj23425;
reg    [`NUM_VC -1:0]     kq72e84;
reg  [31:0]               aa97420[0:`NUM_VC -1];
reg  [31:0]               lfba100[0:`NUM_VC -1];
reg  [31:0]               rgd0807[0:`NUM_VC -1];
reg  [`NUM_VC -1:0]       rv8403a;
reg  [`NUM_VC -1:0]       hq201d6;
reg  [`NUM_VC -1:0]       ymeb3;
reg  [`NUM_VC -1:0]       qv7599;
reg  [`NUM_VC -1:0]       do3accd;
reg  [`NUM_VC -1:0]       czd666a;
reg  [`NUM_VC -1:0]       ymb3354;
reg  [`NUM_VC -1:0]       ng99aa1;
reg  [`NUM_VC -1:0]       pfcd50a;
reg  [`NUM_VC -1:0]       wj6a856;
reg  [`NUM_VC -1:0]       uv542b5;
reg                       sja15ad;
reg                       iead6d;
reg  [31:0]               tud0960;
reg  [wjcc96b:0]            doada0f;
reg                       su6d07a;
reg                       me683d1;
reg  [wjcc96b:0]            swf44d;
reg  [wjcc96b:0]            qgd134d;
reg  [1:0]                ls89a69 [0:`NUM_VC -1];
reg  [1:0]                tu4d34b [0:`NUM_VC -1];
reg  [1:0]                by69a5a [0:`NUM_VC -1];
reg                       dm4d2d2;
reg                       dm69692;
reg  [wjcc96b:0]            vv5a49d;
reg  [wjcc96b:0]            qi92776;
reg                       hq93bb0;
reg                       qi9dd83;
reg  [31:0]               hd84b02;
reg  [31:0]               jc760c3;
reg  [31:0]               zzb061b;
reg                       ri830de;
reg                       mt186f3;
reg                       kdc379d;
reg                       hq1bced;
reg                       uide76b;
reg  [31:0]               thf3b58;
reg                       uk9dac6;
reg                       shed630;
reg                       pf6b185;
reg                       lq58c2e;
reg                       yxc6172;
reg  [wjcc96b:0]            ux85cab;
reg  [wjcc96b:0]            go72ae8 [fn64b5d:0];
reg  [wjcc96b:0]            lq5d02d;
reg  [wjcc96b:0]            rt40b5d;
reg  [wjcc96b:0]            jr2d779;
reg  [wjcc96b:0]            lq5de7f;
reg                       wwef3fa;
reg  [wjcc96b:0]            xwcfe83;
reg                       ip7f41a;
reg  [wjcc96b:0]            vid06a9;
reg  [wjcc96b:0]            wy1aa5b [fn64b5d:0];
reg  [wjcc96b:0]            uv4b659;
reg  [wjcc96b:0]            wjd966c;
reg  [wjcc96b:0]            kq59b29;
reg  [wjcc96b:0]            ps6ca47;
reg                       mr6523a;
reg  [wjcc96b:0]            ho48ead;
reg  [13:0]               ne4756b;
reg                       fc3ab5b;
reg                       rgd5ada;
reg                       puad6d2;
reg                       rt6b693;
reg  [3:0]                cz5b49e;
reg  [3:0]                dmda4f4;
reg  [3:0]                nrd27a2;
reg  [3:0]                je93d16;
reg  [FADDR:0]            lqf459f;
reg                       jea2cfa;
reg    [FADDR:0]          oub3e9e;
reg    [FADDR:0]          ykfa784;
reg    [FADDR:0]          db9e10d;
integer                   kqf086e, hd84371, ec21b8e, yzdc70, vv6e385, jp71c2e;
reg  [wjcc96b:0]            cz70bbf [`NUM_VC -1:0];
reg  [wjcc96b:0]            ie2efed [`NUM_VC -1:0];
reg  [wjcc96b:0]            dbbfb48 [`NUM_VC -1:0];
wire [wjcc96b:0]            yxed235;
wire [wjcc96b:0]            tu48d6b;
wire [wjcc96b:0]            hq35ad8;
`ifdef VC1
`else
`ifdef VC2
`else
`ifdef VC3
`else
`ifdef VC4
`else
`endif
`endif
`endif
`endif
`ifdef EN_VC0
wire [2:0] hof43fe = 3'b000;
`endif
`ifdef EN_VC1
wire [2:0] epa1ff2 = ay5cd66[5:3];
`endif
`ifdef EN_VC2
wire [2:0] wyff94 = ay5cd66[8:6];
`endif
`ifdef EN_VC3
wire [2:0] al7fca0 = ay5cd66[11:9];
`endif
`ifdef EN_VC4
wire [2:0] dmfe504 = ay5cd66[14:12];
`endif
`ifdef EN_VC5
wire [2:0] gbf2823 = ay5cd66[17:15];
`endif
`ifdef EN_VC6
wire [2:0] xl9411c = ay5cd66[20:18];
`endif
`ifdef EN_VC7
wire [2:0] rva08e7 = ay5cd66[23:21];
`endif
`ifdef EN_VC0
`endif
`ifdef EN_VC1
`endif
`ifdef EN_VC2
`endif
`ifdef EN_VC3
`endif
`ifdef EN_VC4
`endif
`ifdef EN_VC5
`endif
`ifdef EN_VC6
`endif
`ifdef EN_VC7
`endif
`ifdef EN_VC0
`endif
`ifdef EN_VC1
`endif
`ifdef EN_VC2
`endif
`ifdef EN_VC3
`endif
`ifdef EN_VC4
`endif
`ifdef EN_VC5
`endif
`ifdef EN_VC6
`endif
`ifdef EN_VC7
`endif
wire [1:0]  off2268  = ls89a69[0];
wire [1:0]  ng89a2f  = tu4d34b[0];
wire [1:0]  yk68bda  = by69a5a[0];
wire [31:0]  je2f687     = aa97420[0];
wire [31:0]  neda1d7    = lfba100[0];
wire [31:0]  ie875d2   = rgd0807[0];
reg [13 : 0] ldd748a;
reg vxba456;
reg vvd22b7;
reg xl915be;
reg [2 : 0] qv8adf7;
reg [1 : 0] cm56fbc;
reg dob7de1;
reg [2 : 0] yzbef0a;
reg [1 : 0] off7854;
reg [`NUM_VC - 1 : 0] gqbc2a4;
reg [`NUM_VC - 1 : 0] zke1520;
reg [`NUM_VC - 1 : 0] mga903;
reg [(`NUM_VC * 3) - 1 : 0] cz75325;
reg uxa40c4;
reg [2 : 0] zm20625;
reg ph312b;
reg [23 : 0] wl1895f;
reg ldd88f4;
reg wwc47a6;
reg co2bf0b;
reg [11 : 0] rt5f859;
reg zxfc2cf;
reg vie167e;
reg [2 : 0] hqb3f3;
reg me59f9b;
reg [1 : 0] facfcd8;
reg [`NUM_VC - 1 : 0] vv7e6c2;
reg vvf3617;
reg rv9b0bf;
reg vvd85fe;
reg fnc2ff7;
reg [`NUM_VC - 1 : 0] qv17fbe;
reg [`NUM_VC - 1 : 0] ntbfdf5;
reg [`NUM_VC - 1 : 0] dmfefae;
reg [`NUM_VC - 1 : 0] czf7d72;
reg [`NUM_VC - 1 : 0] qvbeb94;
reg [`NUM_VC - 1 : 0] ayf5ca4;
reg [`NUM_VC - 1 : 0] epae521;
reg [`NUM_VC - 1 : 0] ay7290c;
reg [`NUM_VC - 1 : 0] bn94860;
reg [`NUM_VC - 1 : 0] sja4306;
reg [`NUM_VC - 1 : 0] ie21835;
reg [`NUM_VC - 1 : 0] fpc1a8;
reg uv60d46;
reg xl6a34;
reg [wjcc96b : 0] xya8d32;
reg ww46992;
reg uk34c90;
reg [wjcc96b : 0] ph32408;
reg [wjcc96b : 0] yz90238;
reg zz811c5;
reg ux8e2e;
reg [wjcc96b : 0] hd38bab;
reg [wjcc96b : 0] ou2eafb;
reg ip757d9;
reg mtabecc;
reg [31 : 0] th5f665;
reg [31 : 0] jcfb32e;
reg czd9973;
reg enccb9c;
reg qt65ce5;
reg ou2e72c;
reg dm73960;
reg [31 : 0] xy9cb02;
reg ose5812;
reg an2c090;
reg al60485;
reg wl242d;
reg an1216d;
reg [wjcc96b : 0] mt85b64;
reg [wjcc96b : 0] me6d92e;
reg [wjcc96b : 0] xj64b82;
reg [wjcc96b : 0] mg2e0b2;
reg [wjcc96b : 0] gq82c84;
reg zz16420;
reg [wjcc96b : 0] mt90833;
reg db8419c;
reg [wjcc96b : 0] lf6732;
reg [wjcc96b : 0] xy9ccbc;
reg [wjcc96b : 0] zz32f16;
reg [wjcc96b : 0] ksbc5b1;
reg [wjcc96b : 0] tj16c45;
reg ieb622f;
reg [wjcc96b : 0] wy88bcc;
reg [13 : 0] fn45e61;
reg tw2f30f;
reg rg7987a;
reg ofcc3d3;
reg pf61e9c;
reg [3 : 0] gqf4e6;
reg [3 : 0] gb7a731;
reg [3 : 0] end398d;
reg [3 : 0] tw9cc6d;
reg [FADDR : 0] aa31b56;
reg co8dab1;
reg [FADDR : 0] kd6ac49;
reg [FADDR : 0] kfb1268;
reg [FADDR : 0] me49a22;
reg [wjcc96b : 0] me6888a;
reg [wjcc96b : 0] lf22284;
reg [wjcc96b : 0] wl8a133;
reg [1 : 0] fn5099d;
reg [1 : 0] zz84cee;
reg [1 : 0] yz26777;
reg [31 : 0] cb33bbc;
reg [31 : 0] ou9dde4;
reg [31 : 0] vieef20;
reg [2047:0] necf6c2;
wire [106:0] ld7b613;
`ifdef LW1
`else
`ifdef LW2
`else
`ifdef LW4
`else
`endif
`endif
`endif
`ifdef VC1
`else
`ifdef VC2
`else
`ifdef VC3
`else
`ifdef VC4
`else
`endif
`endif
`endif
`endif
`ifdef VC1
`else
`ifdef VC2
`else
`ifdef VC3
`else
`ifdef VC4
`else
`endif
`endif
`endif
`endif
`ifdef EN_VC0
`endif
`ifdef EN_VC1
`endif
`ifdef EN_VC2
`endif
`ifdef EN_VC3
`endif
`ifdef EN_VC4
`endif
`ifdef EN_VC5
`endif
`ifdef EN_VC6
`endif
`ifdef EN_VC7
`endif
`ifdef VC1
`else
`ifdef VC2
`else
`ifdef VC3
`else
`ifdef VC4
`else
`endif
`endif
`endif
`endif
`ifdef EN_VC0
`endif
`ifdef EN_VC1
`endif
`ifdef EN_VC2
`endif
`ifdef EN_VC3
`endif
`ifdef EN_VC4
`endif
`ifdef EN_VC5
`endif
`ifdef EN_VC6
`endif
`ifdef EN_VC7
`endif
`ifdef EN_VC0
`endif
`ifdef EN_VC1
`endif
`ifdef EN_VC2
`endif
`ifdef EN_VC3
`endif
`ifdef EN_VC4
`endif
`ifdef EN_VC5
`endif
`ifdef EN_VC6
`endif
`ifdef EN_VC7
`endif
`ifdef EN_VC0
`endif
`ifdef EN_VC1
`endif
`ifdef EN_VC2
`endif
`ifdef EN_VC3
`endif
`ifdef EN_VC4
`endif
`ifdef EN_VC5
`endif
`ifdef EN_VC6
`endif
`ifdef EN_VC7
`endif
localparam qgdb09f = 107,nrd84f8 = 32'hfdffd42b;
localparam [31:0] thc27c7 = nrd84f8;
localparam mt9f1ff = nrd84f8 & 4'hf;
localparam [11:0] fnc7fe5 = 'h7ff;
wire  [(1 << mt9f1ff)  -1:0] suff972;
reg    [qgdb09f-1:0] cme5c87;
reg [mt9f1ff-1:0] qg721c0 [0:1];
reg [mt9f1ff-1:0] ym8700c;
reg rv38061;
integer jcc030e;
integer vk1872;
`ifdef LW1
`else
`ifdef LW2
`else
`ifdef LW4
`else
`endif
`endif
`endif
`ifdef VC1
`else
`ifdef VC2
`else
`ifdef VC3
`else
`ifdef VC4
`else
`endif
`endif
`endif
`endif
`ifdef VC1
`else
`ifdef VC2
`else
`ifdef VC3
`else
`ifdef VC4
`else
`endif
`endif
`endif
`endif
`ifdef EN_VC0
`endif
`ifdef EN_VC1
`endif
`ifdef EN_VC2
`endif
`ifdef EN_VC3
`endif
`ifdef EN_VC4
`endif
`ifdef EN_VC5
`endif
`ifdef EN_VC6
`endif
`ifdef EN_VC7
`endif
`ifdef VC1
`else
`ifdef VC2
`else
`ifdef VC3
`else
`ifdef VC4
`else
`endif
`endif
`endif
`endif
`ifdef EN_VC0
`endif
`ifdef EN_VC1
`endif
`ifdef EN_VC2
`endif
`ifdef EN_VC3
`endif
`ifdef EN_VC4
`endif
`ifdef EN_VC5
`endif
`ifdef EN_VC6
`endif
`ifdef EN_VC7
`endif
`ifdef EN_VC0
`endif
`ifdef EN_VC1
`endif
`ifdef EN_VC2
`endif
`ifdef EN_VC3
`endif
`ifdef EN_VC4
`endif
`ifdef EN_VC5
`endif
`ifdef EN_VC6
`endif
`ifdef EN_VC7
`endif
`ifdef EN_VC0
`endif
`ifdef EN_VC1
`endif
`ifdef EN_VC2
`endif
`ifdef EN_VC3
`endif
`ifdef EN_VC4
`endif
`ifdef EN_VC5
`endif
`ifdef EN_VC6
`endif
`ifdef EN_VC7
`endif
`ifdef LW1
`else
`ifdef LW2
`else
`ifdef LW4
`else
`endif
`endif
`endif
`ifdef VC1
`else
`ifdef VC2
`else
`ifdef VC3
`else
`ifdef VC4
`else
`endif
`endif
`endif
`endif
`ifdef VC1
`else
`ifdef VC2
`else
`ifdef VC3
`else
`ifdef VC4
`else
`endif
`endif
`endif
`endif
`ifdef EN_VC0
`endif
`ifdef EN_VC1
`endif
`ifdef EN_VC2
`endif
`ifdef EN_VC3
`endif
`ifdef EN_VC4
`endif
`ifdef EN_VC5
`endif
`ifdef EN_VC6
`endif
`ifdef EN_VC7
`endif
always @(posedge sys_clk or negedge rst_n) begin   if (rst_n == 1'b0) begin      zzb061b      <= 32'd0;      ri830de   <= 1'b0;      mt186f3 <= 1'b0;      kdc379d     <= 1'b0;      hq1bced      <= 1'b0;      uide76b        <= 1'b0;   end   else begin            if(ldd88f4 || wwc47a6 || co2bf0b)         zzb061b[11:0]  <= rt5f859;      zzb061b[23:12] <= 12'h000;              if(ldd88f4)         zzb061b[31:24]  <= 8'b0001_0000;          else if(((wwc47a6 || vvd85fe) && !dm73960) || co2bf0b)         zzb061b[31:24]  <= 8'b0000_0000;
            hq1bced  <= (ldd88f4 || wwc47a6 || vvd85fe) ? 1'b1 : 1'b0;            if(zz16420 && (mt90833 == hd2d772))         uide76b <= 1'b0;      else if(ldd88f4)         uide76b <= 1'b1;
            if(zz16420 && (mt90833 == hd2d772))         kdc379d <= 1'b0;      else if(ou2e72c)         kdc379d <= 1'b1;            ri830de  <= ou2e72c & !qt65ce5;            mt186f3  <= czd9973 | uk34c90;   end
end
`ifdef VC1
   assign yxed235  = {1'b0, cm56fbc};           assign tu48d6b  = {1'b0, off7854};   assign hq35ad8 = {1'b0, facfcd8};
`else
`ifdef VC2
      assign yxed235  = {qv8adf7[0], cm56fbc};      assign tu48d6b  = {yzbef0a[0], off7854};      assign hq35ad8 = {hqb3f3[0], facfcd8};
`else
`ifdef VC3
         assign yxed235  = {qv8adf7[1:0], cm56fbc};         assign tu48d6b  = {yzbef0a[1:0], off7854};         assign hq35ad8 = {hqb3f3[1:0], facfcd8};
`else
`ifdef VC4
            assign yxed235  = {qv8adf7[1:0], cm56fbc};              assign tu48d6b  = {yzbef0a[1:0], off7854};              assign hq35ad8 = {hqb3f3[1:0], facfcd8};
`else
            assign yxed235  = {qv8adf7, cm56fbc};                  assign tu48d6b  = {yzbef0a, off7854};                  assign hq35ad8 = {hqb3f3, facfcd8};
`endif
`endif
`endif
`endif
always @(posedge sys_clk or negedge rst_n) begin   if (rst_n == 1'b0) begin      yxc6172   <= 1'b0;      ux85cab       <= 0;      for(kqf086e=0; kqf086e<=fn64b5d; kqf086e=kqf086e+1)         go72ae8[kqf086e]     <= 0;      lq5d02d       <= 0;      rt40b5d     <= 0;      jr2d779    <= 0;   end   else begin                        lq5d02d <= me6888a;            rt40b5d  <= me6d92e;            if(czd9973)         jr2d779 <= hd2d772;      else         jr2d779 <= (uk34c90) ? yz90238 : xj64b82;            yxc6172  <= |ntbfdf5;                  if(an1216d || enccb9c)         ux85cab  <= mt85b64 + 1;      if(an1216d || enccb9c)         go72ae8[mt85b64]  <= mg2e0b2;   end
end
always @(posedge sys_clk or negedge rst_n) begin   if (rst_n == 1'b0) begin      for(hd84371=0; hd84371<`NUM_VC; hd84371=hd84371+1) begin                  ls89a69[hd84371]       <= 2'b01;         tu4d34b[hd84371]      <= 2'b01;         by69a5a[hd84371]     <= 2'b01;      end      su6d07a         <= 1'b0;      me683d1       <= 1'b0;      swf44d         <= 0;      qgd134d       <= 0;      xjc264f           <= 1'b1;      fc3ab5b         <= 1'b1;   end   else begin
                        for(hd84371=0; hd84371<`NUM_VC; hd84371=hd84371+1) begin         if((hqb3f3 == hd84371) && (zxfc2cf || vie167e)) begin            if(me59f9b) begin                  ls89a69[hd84371]   <= 2'b11;               tu4d34b[hd84371]  <= 2'b11;               by69a5a[hd84371] <= 2'b11;            end            else begin                 ls89a69[hd84371]   <= 2'b01;               tu4d34b[hd84371]  <= 2'b01;               by69a5a[hd84371] <= 2'b01;            end         end                  else if(!qv17fbe[hd84371]) begin                          if(!gqbc2a4[hd84371])               ls89a69[hd84371]   <= 2'b10;                if(!zke1520[hd84371])               tu4d34b[hd84371]  <= 2'b10;                if(!mga903[hd84371])               by69a5a[hd84371] <= 2'b10;             end      end            su6d07a   <= zxfc2cf;      if(zxfc2cf)            swf44d   <= wl8a133;            me683d1  <= ww46992;      qgd134d  <= ph32408;
                  if(zxfc2cf)         xjc264f  <= 1'b0;      else if(zz16420 && (mt90833 == ph32408))         xjc264f  <= 1'b1;
      fc3ab5b  <= xjc264f;   end
end
always @(posedge sys_clk or negedge rst_n) begin   if (rst_n == 1'b0) begin      dm4d2d2        <= 1'b0;      dm69692      <= 1'b0;      vv5a49d        <= 0;      qi92776      <= 0;      jr1327f          <= 1'b1;         end   else begin            dm4d2d2   <= vie167e;      if(vie167e)            vv5a49d   <= wl8a133;            dm69692  <= zz811c5;      qi92776  <= hd38bab;
                  if(vie167e)         jr1327f  <= 1'b0;      else if(ieb622f && (wy88bcc == hd38bab))         jr1327f  <= 1'b1;
         end
end
always @(posedge sys_clk or negedge rst_n) begin   if (rst_n == 1'b0) begin      puad6d2          <= 1'b0;      rt6b693          <= 1'b0;      cz5b49e          <= 0;      dmda4f4     <= 0;      nrd27a2     <= 0;      je93d16     <= 0;   end   else begin      puad6d2 <= 1'b0;      rt6b693 <= 1'b0;      if(vxba456 || ofcc3d3) begin         if(an1216d || enccb9c || vvd22b7)             puad6d2     <= 1'b1;         else begin            rt6b693     <= 1'b1;            cz5b49e     <= gqf4e6 + 3'b001;            end      end      dmda4f4 <= gqf4e6;      nrd27a2 <= gb7a731;      je93d16 <= end398d;   end
end
always @(posedge sys_clk or negedge rst_n) begin   if (rst_n == 1'b0) begin      rgd5ada            <= 1'b0;      ba250d2       <= 0;      oub3e9e  <= 0;      ykfa784       <= 0;      mec4930       <= 0;      lqf459f             <= 0;      jea2cfa       <= 1'b0;   end   else begin      rgd5ada       <= an1216d | enccb9c;      ba250d2  <= aa31b56;      jea2cfa  <= vvd22b7;      if(vvd22b7)          mec4930 <= tw9cc6d;        oub3e9e <= ~ba250d2 + 1;              if((an1216d || enccb9c) && vvd22b7)          ykfa784  <= kd6ac49 + 1;              else         ykfa784  <= kd6ac49;        lqf459f <= aa31b56 + me49a22;   end
end
always @(kfb1268 or rg7987a or pf61e9c or co8dab1) begin      case({rg7987a, pf61e9c, co8dab1})         3'b100,         3'b010   : db9e10d = 1;            3'b001,         3'b101   : db9e10d = kfb1268;         default  : db9e10d = 0;      endcase
end
always @(posedge sys_clk or negedge rst_n) begin   if (rst_n == 1'b0) begin      sj23425     <= 1'b0;      doada0f       <= 0;      an3c4c4     <= 1'b0;      wwef3fa     <= 1'b0;      lq5de7f     <= 0;      xwcfe83   <= 0;      ene2624     <= 1'b0;      mr6523a     <= 1'b0;      ps6ca47     <= 0;      ho48ead   <= 0;   end   else begin            sj23425   <= zz16420 || ieb622f;         if(rv9b0bf)         doada0f    <= wy1aa5b[tj16c45];      else         doada0f    <= go72ae8[gq82c84];            an3c4c4   <= (mt85b64 != gq82c84) ? 1'b1 : 1'b0;      xwcfe83 <= go72ae8[gq82c84];      wwef3fa     <= 1'b0;      if(vvf3617) begin         wwef3fa     <= 1'b1;         lq5de7f     <= gq82c84 + 1;      end            ene2624   <= (lf6732 != tj16c45) ? 1'b1 : 1'b0;      ho48ead <= wy1aa5b[tj16c45];      mr6523a     <= 1'b0;      if(rv9b0bf) begin         mr6523a     <= 1'b1;         ps6ca47     <= tj16c45 + 1;      end   end
end
always @(posedge sys_clk or negedge rst_n) begin   if (rst_n == 1'b0) begin      lq58c2e          <= 1'b0;      pf6b185         <= 1'b0;      uk9dac6       <= 1'b0;      shed630       <= 1'b0;      gqb98bf      <= 1'b0;      ne4756b <= 14'd0;   end   else begin            lq58c2e  <= (co2bf0b && !qt65ce5) ? 1'b1 : 1'b0;            if((ieb622f && (wy88bcc == hd2d772)) || (zz16420 && (mt90833 == hd2d772)))         pf6b185 <= 1'b0;      else if(wl242d)         pf6b185 <= 1'b1;            uk9dac6  <= wl242d & !al60485;            shed630    <= ose5812 | mtabecc | ux8e2e;                  if(al60485)         ne4756b <= fn45e61 + 1;      else         ne4756b <= 14'd0;
      if(fn45e61 == ldd748a)         gqb98bf  <= 1'b1;      else         gqb98bf  <= 1'b0;   end
end
always @(posedge sys_clk or negedge rst_n) begin   if (rst_n == 1'b0) begin      ip7f41a    <= 1'b0;      vid06a9     <= 0;      for(ec21b8e=0; ec21b8e<=fn64b5d; ec21b8e=ec21b8e+1)         wy1aa5b[ec21b8e]     <= 0;      uv4b659       <= 0;      wjd966c     <= 0;      kq59b29    <= 0;   end   else begin                        uv4b659 <= lf22284;            wjd966c  <= xy9ccbc;            if(mtabecc)         kq59b29  <= fc25aee;      else if(ux8e2e)         kq59b29  <= ou2eafb;      else         kq59b29 <= (ose5812) ? hd2d772 : zz32f16;                ip7f41a  <= |dmfefae;                  if(db8419c || an2c090)         vid06a9  <= lf6732 + 1;      if(db8419c || an2c090)         wy1aa5b[lf6732]  <= ksbc5b1;   end
end
always @(posedge sys_clk or negedge rst_n) begin   if (rst_n == 1'b0) begin      hq93bb0      <= 1'b0;      qi9dd83    <= 1'b0;      jc760c3     <= 32'd0;      hd84b02 <= 32'd0;      ec1a12c  <= 1'b0;      vi42b97  <= 1'b0;   end   else begin            hq93bb0 <= uxa40c4 || ph312b;      if(uxa40c4)          jc760c3   <= {5'b00100, zm20625, 24'd0};      else if(ph312b)           jc760c3   <= {8'b00110000, wl1895f};            qi9dd83  <= ip757d9;      if((wy88bcc == fc25aee) && rv9b0bf)         hd84b02 <= th5f665;            vi42b97  <= ((wy88bcc == fc25aee) && rv9b0bf)  ? 1'b1 : 1'b0;      ec1a12c       <= fnc2ff7;   end
end
assign cm46737 = ec1a12c;
`ifdef EN_VC0
   always @(ls89a69[0] or tu4d34b[0] or by69a5a[0] or      hof43fe or hq93919 or ri9c8cb or tue465a) begin      aa97420[0]   = {ls89a69[0], 2'b00, 1'b0, hof43fe, hq93919};      lfba100[0]  = {tu4d34b[0], 2'b01, 1'b0, hof43fe, ri9c8cb};      rgd0807[0] = {by69a5a[0], 2'b10, 1'b0, hof43fe, tue465a};   end
`endif
`ifdef EN_VC1
   always @(ls89a69[1] or tu4d34b[1] or by69a5a[1] or      epa1ff2 or sj232d3 or hd1969c or uicb4e7) begin      aa97420[1]   = {ls89a69[1], 2'b00, 1'b0, epa1ff2, sj232d3};      lfba100[1]  = {tu4d34b[1], 2'b01, 1'b0, epa1ff2, hd1969c};      rgd0807[1] = {by69a5a[1], 2'b10, 1'b0, epa1ff2, uicb4e7};   end
`endif
`ifdef EN_VC2
   always @(ls89a69[2] or tu4d34b[2] or by69a5a[2] or      wyff94 or pf5a739 or end39ce or tw9ce75) begin      aa97420[2]   = {ls89a69[2], 2'b00, 1'b0, wyff94, pf5a739};      lfba100[2]  = {tu4d34b[2], 2'b01, 1'b0, wyff94, end39ce};      rgd0807[2] = {by69a5a[2], 2'b10, 1'b0, wyff94, tw9ce75};   end
`endif
`ifdef EN_VC3
   always @(ls89a69[3] or tu4d34b[3] or by69a5a[3] or      al7fca0 or kde73aa or ux39d54 or kqceaa5) begin      aa97420[3]   = {ls89a69[3], 2'b00, 1'b0, al7fca0, kde73aa};      lfba100[3]  = {tu4d34b[3], 2'b01, 1'b0, al7fca0, ux39d54};      rgd0807[3] = {by69a5a[3], 2'b10, 1'b0, al7fca0, kqceaa5};   end
`endif
`ifdef EN_VC4
   always @(ls89a69[4] or tu4d34b[4] or by69a5a[4] or      dmfe504 or ip75528 or ntaa944 or al54a27) begin      aa97420[4]   = {ls89a69[4], 2'b00, 1'b0, dmfe504, ip75528};      lfba100[4]  = {tu4d34b[4], 2'b01, 1'b0, dmfe504, ntaa944};      rgd0807[4] = {by69a5a[4], 2'b10, 1'b0, dmfe504, al54a27};   end
`endif
`ifdef EN_VC5
   always @(ls89a69[5] or tu4d34b[5] or by69a5a[5] or      gbf2823 or lfa513c or hd289e7 or al44f3e) begin      aa97420[5]   = {ls89a69[5], 2'b00, 1'b0, gbf2823, lfa513c};      lfba100[5]  = {tu4d34b[5], 2'b01, 1'b0, gbf2823, hd289e7};      rgd0807[5] = {by69a5a[5], 2'b10, 1'b0, gbf2823, al44f3e};   end
`endif
`ifdef EN_VC6
   always @(ls89a69[6] or tu4d34b[6] or by69a5a[6] or      xl9411c or hd279f5 or an3cfaf or ipe7d7d) begin      aa97420[6]   = {ls89a69[6], 2'b00, 1'b0, xl9411c, hd279f5};      lfba100[6]  = {tu4d34b[6], 2'b01, 1'b0, xl9411c, an3cfaf};      rgd0807[6] = {by69a5a[6], 2'b10, 1'b0, xl9411c, ipe7d7d};   end
`endif
`ifdef EN_VC7
   always @(ls89a69[7] or tu4d34b[7] or by69a5a[7] or      rva08e7 or gq3ebed or ykf5f68 or phafb41) begin      aa97420[7]   = {ls89a69[7], 2'b00, 1'b0, rva08e7, gq3ebed};      lfba100[7]  = {tu4d34b[7], 2'b01, 1'b0, rva08e7, ykf5f68};      rgd0807[7] = {by69a5a[7], 2'b10, 1'b0, rva08e7, phafb41};   end
`endif
always @(posedge sys_clk or negedge rst_n) begin   if (rst_n == 1'b0) begin      tud0960   <= 32'd0;   end   else begin      case(xya8d32[wjcc96b:0])
`ifdef EN_VC0
            fn6bb97     : tud0960  <= aa97420[0];            ne5dcbf    : tud0960  <= lfba100[0];            neee5fa   : tud0960  <= rgd0807[0];
`endif
`ifdef EN_VC1
            ksf3af     : tud0960  <= aa97420[1];            lq79d79    : tud0960  <= lfba100[1];            qgcebcb   : tud0960  <= rgd0807[1];
`endif
`ifdef EN_VC2
            ea5307d     : tud0960  <= aa97420[2];            ou983e8    : tud0960  <= lfba100[2];            ykc1f41   : tud0960  <= rgd0807[2];
`endif
`ifdef EN_VC3
            shcc581     : tud0960  <= aa97420[3];            su62c0c    : tud0960  <= lfba100[3];            lf16061   : tud0960  <= rgd0807[3];
`endif
`ifdef EN_VC4
            uic1c8f     : tud0960  <= aa97420[4];            jee479    : tud0960  <= lfba100[4];            cm723cb   : tud0960  <= rgd0807[4];
`endif
`ifdef EN_VC5
            vx91e59     : tud0960  <= aa97420[5];            wl8f2ce    : tud0960  <= lfba100[5];            dm79675   : tud0960  <= rgd0807[5];
`endif
`ifdef EN_VC6
            aycb3aa     : tud0960  <= aa97420[6];            ic59d51    : tud0960  <= lfba100[6];            ykcea88   : tud0960  <= rgd0807[6];
`endif
`ifdef EN_VC7
            qt75440     : tud0960  <= aa97420[7];            zzaa204    : tud0960  <= lfba100[7];            of51026   : tud0960  <= rgd0807[7];
`endif
         default  : tud0960  <= jcfb32e;       endcase   end
end
`ifdef EN_VC0
always @(posedge sys_clk or negedge rst_n) begin   if (rst_n == 1'b0) begin      cz70bbf[0]   <= fn6bb97;      ie2efed[0]  <= ne5dcbf;      dbbfb48[0] <= neee5fa;   end   else begin      cz70bbf[0]   <= fn6bb97;      ie2efed[0]  <= ne5dcbf;      dbbfb48[0] <= neee5fa;   end
end
`endif
`ifdef EN_VC1
always @(posedge sys_clk or negedge rst_n) begin   if (rst_n == 1'b0) begin      cz70bbf[1]   <= ksf3af;      ie2efed[1]  <= lq79d79;      dbbfb48[1] <= qgcebcb;   end   else begin      cz70bbf[1]   <= ksf3af;      ie2efed[1]  <= lq79d79;      dbbfb48[1] <= qgcebcb;   end
end
`endif
`ifdef EN_VC2
always @(posedge sys_clk or negedge rst_n) begin   if (rst_n == 1'b0) begin      cz70bbf[2]   <= ea5307d;      ie2efed[2]  <= ou983e8;      dbbfb48[2] <= ykc1f41;   end   else begin      cz70bbf[2]   <= ea5307d;      ie2efed[2]  <= ou983e8;      dbbfb48[2] <= ykc1f41;   end
end
`endif
`ifdef EN_VC3
always @(posedge sys_clk or negedge rst_n) begin   if (rst_n == 1'b0) begin      cz70bbf[3]   <= shcc581;      ie2efed[3]  <= su62c0c;      dbbfb48[3] <= lf16061;   end   else begin      cz70bbf[3]   <= shcc581;      ie2efed[3]  <= su62c0c;      dbbfb48[3] <= lf16061;   end
end
`endif
`ifdef EN_VC4
always @(posedge sys_clk or negedge rst_n) begin   if (rst_n == 1'b0) begin      cz70bbf[4]   <= uic1c8f;      ie2efed[4]  <= jee479;      dbbfb48[4] <= cm723cb;   end   else begin      cz70bbf[4]   <= uic1c8f;      ie2efed[4]  <= jee479;      dbbfb48[4] <= cm723cb;   end
end
`endif
`ifdef EN_VC5
always @(posedge sys_clk or negedge rst_n) begin   if (rst_n == 1'b0) begin      cz70bbf[5]   <= vx91e59;      ie2efed[5]  <= wl8f2ce;      dbbfb48[5] <= dm79675;   end   else begin      cz70bbf[5]   <= vx91e59;      ie2efed[5]  <= wl8f2ce;      dbbfb48[5] <= dm79675;   end
end
`endif
`ifdef EN_VC6
always @(posedge sys_clk or negedge rst_n) begin   if (rst_n == 1'b0) begin      cz70bbf[6]   <= aycb3aa;      ie2efed[6]  <= ic59d51;      dbbfb48[6] <= ykcea88;   end   else begin      cz70bbf[6]   <= aycb3aa;      ie2efed[6]  <= ic59d51;      dbbfb48[6] <= ykcea88;   end
end
`endif
`ifdef EN_VC7
always @(posedge sys_clk or negedge rst_n) begin   if (rst_n == 1'b0) begin      cz70bbf[7]   <= qt75440;      ie2efed[7]  <= zzaa204;      dbbfb48[7] <= of51026;   end   else begin      cz70bbf[7]   <= qt75440;      ie2efed[7]  <= zzaa204;      dbbfb48[7] <= of51026;   end
end
`endif
always @(posedge sys_clk or negedge rst_n) begin   if (rst_n == 1'b0) begin      for(yzdc70=0; yzdc70<`NUM_VC; yzdc70=yzdc70+1) begin         ymeb3[yzdc70]   <= 1'b0;         qv7599[yzdc70]  <= 1'b0;         do3accd[yzdc70] <= 1'b0;         czd666a[yzdc70]  <= 1'b0;         ymb3354[yzdc70] <= 1'b0;         ng99aa1[yzdc70]<= 1'b0;         pfcd50a[yzdc70]  <= 1'b0;         wj6a856[yzdc70] <= 1'b0;         uv542b5[yzdc70]<= 1'b0;      end      sja15ad     <= 1'b0;      iead6d     <= 1'b0;      rv8403a   <= 0;      hq201d6   <= 0;   end   else begin      sja15ad  <= xl915be;      iead6d  <= dob7de1;      for(yzdc70=0; yzdc70<`NUM_VC; yzdc70=yzdc70+1) begin                  ymeb3[yzdc70]   <= 1'b0;         qv7599[yzdc70]  <= 1'b0;         do3accd[yzdc70] <= 1'b0;         if((xl915be && qv8adf7 == yzdc70) || (dob7de1 && yzbef0a == yzdc70)) begin            case(cm56fbc)               uvc3724   : ymeb3[yzdc70]   <= 1'b1;               je1b925  : qv7599[yzdc70]  <= 1'b1;               mrdc92b : do3accd[yzdc70] <= 1'b1;            endcase         end                                    if(zz16420 && (mt90833 == cz70bbf[yzdc70]))            czd666a[yzdc70] <= 1'b0;         else if(czf7d72[yzdc70] && uv60d46)            czd666a[yzdc70] <= 1'b1;         if(zz16420 && (mt90833 == ie2efed[yzdc70]))            ymb3354[yzdc70] <= 1'b0;         else if(qvbeb94[yzdc70] && uv60d46)            ymb3354[yzdc70] <= 1'b1;         if(zz16420 && (mt90833 == dbbfb48[yzdc70]))            ng99aa1[yzdc70] <= 1'b0;         else if(ayf5ca4[yzdc70] && uv60d46)            ng99aa1[yzdc70] <= 1'b1;                  rv8403a[yzdc70]    <= uv60d46 & ((czf7d72[yzdc70] & !epae521[yzdc70]) |                          (qvbeb94[yzdc70] & !ay7290c[yzdc70]) | (ayf5ca4[yzdc70] & !bn94860[yzdc70]));                           if(ieb622f && (wy88bcc == cz70bbf[yzdc70]))            pfcd50a[yzdc70] <= 1'b0;                  else if(czf7d72[yzdc70] && xl6a34 && !epae521[yzdc70])            pfcd50a[yzdc70] <= 1'b1;         if(ieb622f && (wy88bcc == ie2efed[yzdc70]))            wj6a856[yzdc70] <= 1'b0;         else if(qvbeb94[yzdc70] && xl6a34 && !ay7290c[yzdc70])            wj6a856[yzdc70] <= 1'b1;         if(ieb622f && (wy88bcc == dbbfb48[yzdc70]))            uv542b5[yzdc70] <= 1'b0;         else if(ayf5ca4[yzdc70] && xl6a34 && !bn94860[yzdc70])            uv542b5[yzdc70] <= 1'b1;                  hq201d6[yzdc70]    <= xl6a34 & ((czf7d72[yzdc70] & !epae521[yzdc70] & !sja4306[yzdc70]) |                          (qvbeb94[yzdc70] & !ay7290c[yzdc70] & !ie21835[yzdc70]) |                          (ayf5ca4[yzdc70] & !bn94860[yzdc70] & !fpc1a8[yzdc70]));      end    end
end
always @(posedge sys_clk or negedge rst_n) begin   if (rst_n == 1'b0) begin      jpd27c8   <= 0;      do93e46  <= 0;      mt9f233 <= 0;   end   else begin      for(vv6e385=0; vv6e385<`NUM_VC; vv6e385=vv6e385+1) begin         jpd27c8[vv6e385]   <= 1'b0;         do93e46[vv6e385]  <= 1'b0;         mt9f233[vv6e385] <= 1'b0;         if((zz16420 && (mt90833 == cz70bbf[vv6e385])) ||            (ieb622f && (wy88bcc == cz70bbf[vv6e385])))            jpd27c8[vv6e385] <= 1'b1;         if((zz16420 && (mt90833 == ie2efed[vv6e385])) ||            (ieb622f && (wy88bcc == ie2efed[vv6e385])))            do93e46[vv6e385] <= 1'b1;         if((zz16420 && (mt90833 == dbbfb48[vv6e385])) ||            (ieb622f && (wy88bcc == dbbfb48[vv6e385])))            mt9f233[vv6e385] <= 1'b1;      end   end
end
always @(posedge sys_clk or negedge rst_n) begin   if (rst_n == 1'b0) begin      kq72e84 <= 1;   end   else begin      for(jp71c2e=0; jp71c2e<`NUM_VC; jp71c2e=jp71c2e+1) begin         if(vv7e6c2[jp71c2e])            kq72e84[jp71c2e] <= 1'b1;         else if(!vv7e6c2[jp71c2e] && (mt9f233[jp71c2e] || co2bf0b || ldd88f4))            kq72e84[jp71c2e] <= 1'b0;      end   end
end
always@* begin ldd748a<={pse18cc>>1,ld7b613[0]};vxba456<=ld7b613[1];vvd22b7<=ld7b613[2];xl915be<=ld7b613[3];qv8adf7<={yxcc596>>1,ld7b613[4]};cm56fbc<={os62cb4>>1,ld7b613[5]};dob7de1<=ld7b613[6];yzbef0a<={xyb2d0e>>1,ld7b613[7]};off7854<={ba96872>>1,ld7b613[8]};gqbc2a4<={wlb4393>>1,ld7b613[9]};zke1520<={uxa1c9c>>1,ld7b613[10]};mga903<={vke4e4>>1,ld7b613[11]};cz75325<={ay5cd66>>1,ld7b613[12]};uxa40c4<=ld7b613[13];zm20625<={qted079>>1,ld7b613[14]};ph312b<=ld7b613[15];wl1895f<={tx_vsd_data>>1,ld7b613[16]};ldd88f4<=ld7b613[17];wwc47a6<=ld7b613[18];co2bf0b<=ld7b613[19];rt5f859<={jce1a71>>1,ld7b613[20]};zxfc2cf<=ld7b613[21];vie167e<=ld7b613[22];hqb3f3<={tw1e0f1>>1,ld7b613[23]};me59f9b<=ld7b613[24];facfcd8<={ls83c50>>1,ld7b613[25]};vv7e6c2<={ls1e282>>1,ld7b613[26]};vvf3617<=ld7b613[27];rv9b0bf<=ld7b613[28];vvd85fe<=ld7b613[29];fnc2ff7<=ld7b613[30];qv17fbe<={kq72e84>>1,ld7b613[31]};ntbfdf5<={rv8403a>>1,ld7b613[32]};dmfefae<={hq201d6>>1,ld7b613[33]};czf7d72<={ymeb3>>1,ld7b613[34]};qvbeb94<={qv7599>>1,ld7b613[35]};ayf5ca4<={do3accd>>1,ld7b613[36]};epae521<={czd666a>>1,ld7b613[37]};ay7290c<={ymb3354>>1,ld7b613[38]};bn94860<={ng99aa1>>1,ld7b613[39]};sja4306<={pfcd50a>>1,ld7b613[40]};ie21835<={wj6a856>>1,ld7b613[41]};fpc1a8<={uv542b5>>1,ld7b613[42]};uv60d46<=ld7b613[43];xl6a34<=ld7b613[44];xya8d32<={doada0f>>1,ld7b613[45]};ww46992<=ld7b613[46];uk34c90<=ld7b613[47];ph32408<={swf44d>>1,ld7b613[48]};yz90238<={qgd134d>>1,ld7b613[49]};zz811c5<=ld7b613[50];ux8e2e<=ld7b613[51];hd38bab<={vv5a49d>>1,ld7b613[52]};ou2eafb<={qi92776>>1,ld7b613[53]};ip757d9<=ld7b613[54];mtabecc<=ld7b613[55];th5f665<={jc760c3>>1,ld7b613[56]};jcfb32e<={zzb061b>>1,ld7b613[57]};czd9973<=ld7b613[58];enccb9c<=ld7b613[59];qt65ce5<=ld7b613[60];ou2e72c<=ld7b613[61];dm73960<=ld7b613[62];xy9cb02<={thf3b58>>1,ld7b613[63]};ose5812<=ld7b613[64];an2c090<=ld7b613[65];al60485<=ld7b613[66];wl242d<=ld7b613[67];an1216d<=ld7b613[68];mt85b64<={ux85cab>>1,ld7b613[69]};me6d92e<={lq5d02d>>1,ld7b613[70]};xj64b82<={rt40b5d>>1,ld7b613[71]};mg2e0b2<={jr2d779>>1,ld7b613[72]};gq82c84<={lq5de7f>>1,ld7b613[73]};zz16420<=ld7b613[74];mt90833<={xwcfe83>>1,ld7b613[75]};db8419c<=ld7b613[76];lf6732<={vid06a9>>1,ld7b613[77]};xy9ccbc<={uv4b659>>1,ld7b613[78]};zz32f16<={wjd966c>>1,ld7b613[79]};ksbc5b1<={kq59b29>>1,ld7b613[80]};tj16c45<={ps6ca47>>1,ld7b613[81]};ieb622f<=ld7b613[82];wy88bcc<={ho48ead>>1,ld7b613[83]};fn45e61<={ne4756b>>1,ld7b613[84]};tw2f30f<=ld7b613[85];rg7987a<=ld7b613[86];ofcc3d3<=ld7b613[87];pf61e9c<=ld7b613[88];gqf4e6<={cz5b49e>>1,ld7b613[89]};gb7a731<={dmda4f4>>1,ld7b613[90]};end398d<={nrd27a2>>1,ld7b613[91]};tw9cc6d<={je93d16>>1,ld7b613[92]};aa31b56<={lqf459f>>1,ld7b613[93]};co8dab1<=ld7b613[94];kd6ac49<={oub3e9e>>1,ld7b613[95]};kfb1268<={ykfa784>>1,ld7b613[96]};me49a22<={db9e10d>>1,ld7b613[97]};me6888a<={yxed235>>1,ld7b613[98]};lf22284<={tu48d6b>>1,ld7b613[99]};wl8a133<={hq35ad8>>1,ld7b613[100]};fn5099d<={off2268>>1,ld7b613[101]};zz84cee<={ng89a2f>>1,ld7b613[102]};yz26777<={yk68bda>>1,ld7b613[103]};cb33bbc<={je2f687>>1,ld7b613[104]};ou9dde4<={neda1d7>>1,ld7b613[105]};vieef20<={ie875d2>>1,ld7b613[106]};end
always@* begin necf6c2[2047]<=jrc662;necf6c2[2046]<=zk63316;necf6c2[2045]<=lq5d02d[0];necf6c2[2044]<=lf198b2;necf6c2[2043]<=rt40b5d[0];necf6c2[2041]<=yxcc596[0];necf6c2[2038]<=jr2d779[0];necf6c2[2035]<=os62cb4[0];necf6c2[2029]<=zzb061b[0];necf6c2[2028]<=lq5de7f[0];necf6c2[2022]<=fp165a1;necf6c2[2011]<=ri830de;necf6c2[2009]<=wwef3fa;necf6c2[1996]<=xyb2d0e[0];necf6c2[1986]<=je2f687[0];necf6c2[1974]<=mt186f3;necf6c2[1971]<=xwcfe83[0];necf6c2[1945]<=ba96872[0];necf6c2[1943]<=qgd134d[0];necf6c2[1924]<=neda1d7[0];necf6c2[1922]<=ls83c50[0];necf6c2[1901]<=kdc379d;necf6c2[1895]<=ip7f41a;necf6c2[1857]<=ne4756b[0];necf6c2[1842]<=wlb4393[0];necf6c2[1839]<=dm4d2d2;necf6c2[1800]<=ie875d2[0];necf6c2[1797]<=ls1e282[0];necf6c2[1791]<=lq58c2e;necf6c2[1784]<=off2268[0];necf6c2[1778]<=su6d07a;necf6c2[1776]<=qia3c1e;necf6c2[1759]<=uk9dac6;necf6c2[1755]<=hq1bced;necf6c2[1742]<=vid06a9[0];necf6c2[1677]<=jea2cfa;necf6c2[1667]<=fc3ab5b;necf6c2[1652]<=kq59b29[0];necf6c2[1637]<=uxa1c9c[0];necf6c2[1631]<=dm69692;necf6c2[1622]<=qted079[0];necf6c2[1546]<=wlb4ebf;necf6c2[1535]<=yxc6172;necf6c2[1531]<=qi9dd83;necf6c2[1520]<=ng89a2f[0];necf6c2[1509]<=me683d1;necf6c2[1504]<=tw1e0f1[0];necf6c2[1471]<=shed630;necf6c2[1468]<=jce1a71[0];necf6c2[1463]<=uide76b;necf6c2[1437]<=uv4b659[0];necf6c2[1391]<=al7fcee;necf6c2[1312]<=ymeb3[0];necf6c2[1307]<=oub3e9e[0];necf6c2[1286]<=rgd5ada;necf6c2[1256]<=ps6ca47[0];necf6c2[1226]<=vke4e4[0];necf6c2[1215]<=vv5a49d[0];necf6c2[1197]<=ww683cd;necf6c2[1153]<=do3accd[0];necf6c2[1135]<=db9e10d[0];necf6c2[1050]<=rt6b693;necf6c2[1044]<=xya75fd;necf6c2[1037]<=ng99aa1[0];necf6c2[1023]<=pse18cc[0];necf6c2[1022]<=ux85cab[0];necf6c2[1014]<=jc760c3[0];necf6c2[993]<=yk68bda[0];necf6c2[971]<=swf44d[0];necf6c2[961]<=icf078a;necf6c2[928]<=ho48ead[0];necf6c2[895]<=pf6b185;necf6c2[892]<=hq35ad8[0];necf6c2[889]<=doada0f[0];necf6c2[888]<=zx74783;necf6c2[879]<=thf3b58[0];necf6c2[838]<=lqf459f[0];necf6c2[826]<=wjd966c[0];necf6c2[811]<=os7da0f;necf6c2[765]<=hq93bb0;necf6c2[734]<=xw69c54;necf6c2[695]<=yx4e2a2;necf6c2[656]<=hq201d6[0];necf6c2[576]<=qv7599[0];necf6c2[567]<=ykfa784[0];necf6c2[525]<=puad6d2;necf6c2[518]<=ymb3354[0];necf6c2[464]<=mr6523a;necf6c2[446]<=tu48d6b[0];necf6c2[444]<=iead6d;necf6c2[419]<=je93d16[0];necf6c2[405]<=ay5cd66[0];necf6c2[382]<=qi92776[0];necf6c2[347]<=tx_vsd_data[0];necf6c2[328]<=rv8403a[0];necf6c2[259]<=czd666a[0];necf6c2[223]<=yxed235[0];necf6c2[222]<=sja15ad;necf6c2[209]<=nrd27a2[0];necf6c2[164]<=kq72e84[0];necf6c2[111]<=uv542b5[0];necf6c2[104]<=dmda4f4[0];necf6c2[82]<=vi42b97;necf6c2[55]<=wj6a856[0];necf6c2[52]<=cz5b49e[0];necf6c2[41]<=lqe4a1a;necf6c2[27]<=pfcd50a[0];end         assign suff972 = necf6c2,ld7b613 = cme5c87;   initial begin   jcc030e = $fopen(".fred");   $fdisplay( jcc030e, "%3h\n%3h", (thc27c7 >> 4) & fnc7fe5, (thc27c7 >> (mt9f1ff+4)) & fnc7fe5 );   $fclose(jcc030e);   $readmemh(".fred", qg721c0);   end   always @ (suff972) begin   ym8700c = qg721c0[1];       for (vk1872=0; vk1872<qgdb09f; vk1872=vk1872+1) begin           cme5c87[vk1872] = suff972[ym8700c];       rv38061  = ^(ym8700c & qg721c0[0]);       ym8700c =  {ym8700c, rv38061};       end   end
endmodule