module header
	// Internal signals
		// Generated Signal List
		// End of Generated Signal List
	// %COMPILER_OPTS%
	// Generated Signal Assignments
	// Generated Instances
	// wiring ...
	// Generated Instances and Port Mappings
		// Generated Instance Port Map for i_avfb_top_rs
		avfb_top_rs i_avfb_top_rs (
		);
		// End of Generated Instance Port Map for i_avfb_top_rs
endmodule