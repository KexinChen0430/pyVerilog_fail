module ram (WrAddress, RdAddress, Data, WE, RdClock, RdClockEn, Reset,
    WrClock, WrClockEn, Q)/* synthesis NGD_DRC_MASK=1 */;
    input wire [13:0] WrAddress;
    input wire [13:0] RdAddress;
    input wire [7:0] Data;
    input wire WE;
    input wire RdClock;
    input wire RdClockEn;
    input wire Reset;
    input wire WrClock;
    input wire WrClockEn;
    output wire [7:0] Q;
    wire scuba_vhi;
    wire scuba_vlo;
    wire raddr13_ff;
    wire mdout1_1_0;
    wire mdout1_0_0;
    wire mdout1_1_1;
    wire mdout1_0_1;
    wire mdout1_1_2;
    wire mdout1_0_2;
    wire mdout1_1_3;
    wire mdout1_0_3;
    wire mdout1_1_4;
    wire mdout1_0_4;
    wire mdout1_1_5;
    wire mdout1_0_5;
    wire mdout1_1_6;
    wire mdout1_0_6;
    wire raddr13_ff2;
    wire mdout1_1_7;
    wire mdout1_0_7;
    VHI scuba_vhi_inst (.Z(scuba_vhi));
    defparam ram_0_0_15.INIT_DATA = "STATIC" ;
    defparam ram_0_0_15.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam ram_0_0_15.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_0_15.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_0_15.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_0_15.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_0_15.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_0_15.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_0_15.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_0_15.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_0_15.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_0_15.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_0_15.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_0_15.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_0_15.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_0_15.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_0_15.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_0_15.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_0_15.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_0_15.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_0_15.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_0_15.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_0_15.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_0_15.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_0_15.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_0_15.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_0_15.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_0_15.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_0_15.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_0_15.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_0_15.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_0_15.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_0_15.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_0_15.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_0_15.CSDECODE_B = "0b000" ;
    defparam ram_0_0_15.CSDECODE_A = "0b000" ;
    defparam ram_0_0_15.WRITEMODE_B = "NORMAL" ;
    defparam ram_0_0_15.WRITEMODE_A = "NORMAL" ;
    defparam ram_0_0_15.GSR = "ENABLED" ;
    defparam ram_0_0_15.RESETMODE = "SYNC" ;
    defparam ram_0_0_15.REGMODE_B = "OUTREG" ;
    defparam ram_0_0_15.REGMODE_A = "OUTREG" ;
    defparam ram_0_0_15.DATA_WIDTH_B = 1 ;
    defparam ram_0_0_15.DATA_WIDTH_A = 1 ;
    DP8KC ram_0_0_15 (.DIA8(scuba_vlo), .DIA7(scuba_vlo), .DIA6(scuba_vlo),
        .DIA5(scuba_vlo), .DIA4(scuba_vlo), .DIA3(scuba_vlo), .DIA2(scuba_vlo),
        .DIA1(Data[0]), .DIA0(scuba_vlo), .ADA12(WrAddress[12]), .ADA11(WrAddress[11]),
        .ADA10(WrAddress[10]), .ADA9(WrAddress[9]), .ADA8(WrAddress[8]),
        .ADA7(WrAddress[7]), .ADA6(WrAddress[6]), .ADA5(WrAddress[5]), .ADA4(WrAddress[4]),
        .ADA3(WrAddress[3]), .ADA2(WrAddress[2]), .ADA1(WrAddress[1]), .ADA0(WrAddress[0]),
        .CEA(WrClockEn), .OCEA(WrClockEn), .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo),
        .CSA1(scuba_vlo), .CSA0(WrAddress[13]), .RSTA(Reset), .DIB8(scuba_vlo),
        .DIB7(scuba_vlo), .DIB6(scuba_vlo), .DIB5(scuba_vlo), .DIB4(scuba_vlo),
        .DIB3(scuba_vlo), .DIB2(scuba_vlo), .DIB1(scuba_vlo), .DIB0(scuba_vlo),
        .ADB12(RdAddress[12]), .ADB11(RdAddress[11]), .ADB10(RdAddress[10]),
        .ADB9(RdAddress[9]), .ADB8(RdAddress[8]), .ADB7(RdAddress[7]), .ADB6(RdAddress[6]),
        .ADB5(RdAddress[5]), .ADB4(RdAddress[4]), .ADB3(RdAddress[3]), .ADB2(RdAddress[2]),
        .ADB1(RdAddress[1]), .ADB0(RdAddress[0]), .CEB(RdClockEn), .OCEB(RdClockEn),
        .CLKB(RdClock), .WEB(scuba_vlo), .CSB2(scuba_vlo), .CSB1(scuba_vlo),
        .CSB0(RdAddress[13]), .RSTB(Reset), .DOA8(), .DOA7(), .DOA6(), .DOA5(),
        .DOA4(), .DOA3(), .DOA2(), .DOA1(), .DOA0(), .DOB8(), .DOB7(), .DOB6(),
        .DOB5(), .DOB4(), .DOB3(), .DOB2(), .DOB1(), .DOB0(mdout1_0_0))
             /* synthesis MEM_LPC_FILE="ram.lpc" */
             /* synthesis MEM_INIT_FILE="INIT_ALL_0s" */;
    defparam ram_0_1_14.INIT_DATA = "STATIC" ;
    defparam ram_0_1_14.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam ram_0_1_14.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_1_14.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_1_14.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_1_14.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_1_14.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_1_14.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_1_14.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_1_14.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_1_14.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_1_14.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_1_14.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_1_14.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_1_14.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_1_14.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_1_14.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_1_14.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_1_14.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_1_14.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_1_14.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_1_14.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_1_14.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_1_14.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_1_14.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_1_14.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_1_14.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_1_14.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_1_14.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_1_14.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_1_14.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_1_14.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_1_14.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_1_14.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_1_14.CSDECODE_B = "0b000" ;
    defparam ram_0_1_14.CSDECODE_A = "0b000" ;
    defparam ram_0_1_14.WRITEMODE_B = "NORMAL" ;
    defparam ram_0_1_14.WRITEMODE_A = "NORMAL" ;
    defparam ram_0_1_14.GSR = "ENABLED" ;
    defparam ram_0_1_14.RESETMODE = "SYNC" ;
    defparam ram_0_1_14.REGMODE_B = "OUTREG" ;
    defparam ram_0_1_14.REGMODE_A = "OUTREG" ;
    defparam ram_0_1_14.DATA_WIDTH_B = 1 ;
    defparam ram_0_1_14.DATA_WIDTH_A = 1 ;
    DP8KC ram_0_1_14 (.DIA8(scuba_vlo), .DIA7(scuba_vlo), .DIA6(scuba_vlo),
        .DIA5(scuba_vlo), .DIA4(scuba_vlo), .DIA3(scuba_vlo), .DIA2(scuba_vlo),
        .DIA1(Data[1]), .DIA0(scuba_vlo), .ADA12(WrAddress[12]), .ADA11(WrAddress[11]),
        .ADA10(WrAddress[10]), .ADA9(WrAddress[9]), .ADA8(WrAddress[8]),
        .ADA7(WrAddress[7]), .ADA6(WrAddress[6]), .ADA5(WrAddress[5]), .ADA4(WrAddress[4]),
        .ADA3(WrAddress[3]), .ADA2(WrAddress[2]), .ADA1(WrAddress[1]), .ADA0(WrAddress[0]),
        .CEA(WrClockEn), .OCEA(WrClockEn), .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo),
        .CSA1(scuba_vlo), .CSA0(WrAddress[13]), .RSTA(Reset), .DIB8(scuba_vlo),
        .DIB7(scuba_vlo), .DIB6(scuba_vlo), .DIB5(scuba_vlo), .DIB4(scuba_vlo),
        .DIB3(scuba_vlo), .DIB2(scuba_vlo), .DIB1(scuba_vlo), .DIB0(scuba_vlo),
        .ADB12(RdAddress[12]), .ADB11(RdAddress[11]), .ADB10(RdAddress[10]),
        .ADB9(RdAddress[9]), .ADB8(RdAddress[8]), .ADB7(RdAddress[7]), .ADB6(RdAddress[6]),
        .ADB5(RdAddress[5]), .ADB4(RdAddress[4]), .ADB3(RdAddress[3]), .ADB2(RdAddress[2]),
        .ADB1(RdAddress[1]), .ADB0(RdAddress[0]), .CEB(RdClockEn), .OCEB(RdClockEn),
        .CLKB(RdClock), .WEB(scuba_vlo), .CSB2(scuba_vlo), .CSB1(scuba_vlo),
        .CSB0(RdAddress[13]), .RSTB(Reset), .DOA8(), .DOA7(), .DOA6(), .DOA5(),
        .DOA4(), .DOA3(), .DOA2(), .DOA1(), .DOA0(), .DOB8(), .DOB7(), .DOB6(),
        .DOB5(), .DOB4(), .DOB3(), .DOB2(), .DOB1(), .DOB0(mdout1_0_1))
             /* synthesis MEM_LPC_FILE="ram.lpc" */
             /* synthesis MEM_INIT_FILE="INIT_ALL_0s" */;
    defparam ram_0_2_13.INIT_DATA = "STATIC" ;
    defparam ram_0_2_13.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam ram_0_2_13.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_2_13.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_2_13.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_2_13.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_2_13.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_2_13.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_2_13.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_2_13.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_2_13.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_2_13.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_2_13.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_2_13.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_2_13.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_2_13.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_2_13.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_2_13.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_2_13.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_2_13.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_2_13.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_2_13.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_2_13.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_2_13.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_2_13.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_2_13.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_2_13.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_2_13.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_2_13.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_2_13.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_2_13.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_2_13.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_2_13.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_2_13.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_2_13.CSDECODE_B = "0b000" ;
    defparam ram_0_2_13.CSDECODE_A = "0b000" ;
    defparam ram_0_2_13.WRITEMODE_B = "NORMAL" ;
    defparam ram_0_2_13.WRITEMODE_A = "NORMAL" ;
    defparam ram_0_2_13.GSR = "ENABLED" ;
    defparam ram_0_2_13.RESETMODE = "SYNC" ;
    defparam ram_0_2_13.REGMODE_B = "OUTREG" ;
    defparam ram_0_2_13.REGMODE_A = "OUTREG" ;
    defparam ram_0_2_13.DATA_WIDTH_B = 1 ;
    defparam ram_0_2_13.DATA_WIDTH_A = 1 ;
    DP8KC ram_0_2_13 (.DIA8(scuba_vlo), .DIA7(scuba_vlo), .DIA6(scuba_vlo),
        .DIA5(scuba_vlo), .DIA4(scuba_vlo), .DIA3(scuba_vlo), .DIA2(scuba_vlo),
        .DIA1(Data[2]), .DIA0(scuba_vlo), .ADA12(WrAddress[12]), .ADA11(WrAddress[11]),
        .ADA10(WrAddress[10]), .ADA9(WrAddress[9]), .ADA8(WrAddress[8]),
        .ADA7(WrAddress[7]), .ADA6(WrAddress[6]), .ADA5(WrAddress[5]), .ADA4(WrAddress[4]),
        .ADA3(WrAddress[3]), .ADA2(WrAddress[2]), .ADA1(WrAddress[1]), .ADA0(WrAddress[0]),
        .CEA(WrClockEn), .OCEA(WrClockEn), .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo),
        .CSA1(scuba_vlo), .CSA0(WrAddress[13]), .RSTA(Reset), .DIB8(scuba_vlo),
        .DIB7(scuba_vlo), .DIB6(scuba_vlo), .DIB5(scuba_vlo), .DIB4(scuba_vlo),
        .DIB3(scuba_vlo), .DIB2(scuba_vlo), .DIB1(scuba_vlo), .DIB0(scuba_vlo),
        .ADB12(RdAddress[12]), .ADB11(RdAddress[11]), .ADB10(RdAddress[10]),
        .ADB9(RdAddress[9]), .ADB8(RdAddress[8]), .ADB7(RdAddress[7]), .ADB6(RdAddress[6]),
        .ADB5(RdAddress[5]), .ADB4(RdAddress[4]), .ADB3(RdAddress[3]), .ADB2(RdAddress[2]),
        .ADB1(RdAddress[1]), .ADB0(RdAddress[0]), .CEB(RdClockEn), .OCEB(RdClockEn),
        .CLKB(RdClock), .WEB(scuba_vlo), .CSB2(scuba_vlo), .CSB1(scuba_vlo),
        .CSB0(RdAddress[13]), .RSTB(Reset), .DOA8(), .DOA7(), .DOA6(), .DOA5(),
        .DOA4(), .DOA3(), .DOA2(), .DOA1(), .DOA0(), .DOB8(), .DOB7(), .DOB6(),
        .DOB5(), .DOB4(), .DOB3(), .DOB2(), .DOB1(), .DOB0(mdout1_0_2))
             /* synthesis MEM_LPC_FILE="ram.lpc" */
             /* synthesis MEM_INIT_FILE="INIT_ALL_0s" */;
    defparam ram_0_3_12.INIT_DATA = "STATIC" ;
    defparam ram_0_3_12.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam ram_0_3_12.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_3_12.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_3_12.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_3_12.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_3_12.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_3_12.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_3_12.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_3_12.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_3_12.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_3_12.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_3_12.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_3_12.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_3_12.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_3_12.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_3_12.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_3_12.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_3_12.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_3_12.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_3_12.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_3_12.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_3_12.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_3_12.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_3_12.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_3_12.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_3_12.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_3_12.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_3_12.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_3_12.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_3_12.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_3_12.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_3_12.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_3_12.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_3_12.CSDECODE_B = "0b000" ;
    defparam ram_0_3_12.CSDECODE_A = "0b000" ;
    defparam ram_0_3_12.WRITEMODE_B = "NORMAL" ;
    defparam ram_0_3_12.WRITEMODE_A = "NORMAL" ;
    defparam ram_0_3_12.GSR = "ENABLED" ;
    defparam ram_0_3_12.RESETMODE = "SYNC" ;
    defparam ram_0_3_12.REGMODE_B = "OUTREG" ;
    defparam ram_0_3_12.REGMODE_A = "OUTREG" ;
    defparam ram_0_3_12.DATA_WIDTH_B = 1 ;
    defparam ram_0_3_12.DATA_WIDTH_A = 1 ;
    DP8KC ram_0_3_12 (.DIA8(scuba_vlo), .DIA7(scuba_vlo), .DIA6(scuba_vlo),
        .DIA5(scuba_vlo), .DIA4(scuba_vlo), .DIA3(scuba_vlo), .DIA2(scuba_vlo),
        .DIA1(Data[3]), .DIA0(scuba_vlo), .ADA12(WrAddress[12]), .ADA11(WrAddress[11]),
        .ADA10(WrAddress[10]), .ADA9(WrAddress[9]), .ADA8(WrAddress[8]),
        .ADA7(WrAddress[7]), .ADA6(WrAddress[6]), .ADA5(WrAddress[5]), .ADA4(WrAddress[4]),
        .ADA3(WrAddress[3]), .ADA2(WrAddress[2]), .ADA1(WrAddress[1]), .ADA0(WrAddress[0]),
        .CEA(WrClockEn), .OCEA(WrClockEn), .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo),
        .CSA1(scuba_vlo), .CSA0(WrAddress[13]), .RSTA(Reset), .DIB8(scuba_vlo),
        .DIB7(scuba_vlo), .DIB6(scuba_vlo), .DIB5(scuba_vlo), .DIB4(scuba_vlo),
        .DIB3(scuba_vlo), .DIB2(scuba_vlo), .DIB1(scuba_vlo), .DIB0(scuba_vlo),
        .ADB12(RdAddress[12]), .ADB11(RdAddress[11]), .ADB10(RdAddress[10]),
        .ADB9(RdAddress[9]), .ADB8(RdAddress[8]), .ADB7(RdAddress[7]), .ADB6(RdAddress[6]),
        .ADB5(RdAddress[5]), .ADB4(RdAddress[4]), .ADB3(RdAddress[3]), .ADB2(RdAddress[2]),
        .ADB1(RdAddress[1]), .ADB0(RdAddress[0]), .CEB(RdClockEn), .OCEB(RdClockEn),
        .CLKB(RdClock), .WEB(scuba_vlo), .CSB2(scuba_vlo), .CSB1(scuba_vlo),
        .CSB0(RdAddress[13]), .RSTB(Reset), .DOA8(), .DOA7(), .DOA6(), .DOA5(),
        .DOA4(), .DOA3(), .DOA2(), .DOA1(), .DOA0(), .DOB8(), .DOB7(), .DOB6(),
        .DOB5(), .DOB4(), .DOB3(), .DOB2(), .DOB1(), .DOB0(mdout1_0_3))
             /* synthesis MEM_LPC_FILE="ram.lpc" */
             /* synthesis MEM_INIT_FILE="INIT_ALL_0s" */;
    defparam ram_0_4_11.INIT_DATA = "STATIC" ;
    defparam ram_0_4_11.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam ram_0_4_11.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_4_11.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_4_11.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_4_11.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_4_11.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_4_11.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_4_11.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_4_11.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_4_11.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_4_11.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_4_11.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_4_11.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_4_11.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_4_11.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_4_11.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_4_11.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_4_11.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_4_11.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_4_11.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_4_11.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_4_11.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_4_11.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_4_11.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_4_11.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_4_11.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_4_11.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_4_11.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_4_11.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_4_11.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_4_11.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_4_11.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_4_11.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_4_11.CSDECODE_B = "0b000" ;
    defparam ram_0_4_11.CSDECODE_A = "0b000" ;
    defparam ram_0_4_11.WRITEMODE_B = "NORMAL" ;
    defparam ram_0_4_11.WRITEMODE_A = "NORMAL" ;
    defparam ram_0_4_11.GSR = "ENABLED" ;
    defparam ram_0_4_11.RESETMODE = "SYNC" ;
    defparam ram_0_4_11.REGMODE_B = "OUTREG" ;
    defparam ram_0_4_11.REGMODE_A = "OUTREG" ;
    defparam ram_0_4_11.DATA_WIDTH_B = 1 ;
    defparam ram_0_4_11.DATA_WIDTH_A = 1 ;
    DP8KC ram_0_4_11 (.DIA8(scuba_vlo), .DIA7(scuba_vlo), .DIA6(scuba_vlo),
        .DIA5(scuba_vlo), .DIA4(scuba_vlo), .DIA3(scuba_vlo), .DIA2(scuba_vlo),
        .DIA1(Data[4]), .DIA0(scuba_vlo), .ADA12(WrAddress[12]), .ADA11(WrAddress[11]),
        .ADA10(WrAddress[10]), .ADA9(WrAddress[9]), .ADA8(WrAddress[8]),
        .ADA7(WrAddress[7]), .ADA6(WrAddress[6]), .ADA5(WrAddress[5]), .ADA4(WrAddress[4]),
        .ADA3(WrAddress[3]), .ADA2(WrAddress[2]), .ADA1(WrAddress[1]), .ADA0(WrAddress[0]),
        .CEA(WrClockEn), .OCEA(WrClockEn), .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo),
        .CSA1(scuba_vlo), .CSA0(WrAddress[13]), .RSTA(Reset), .DIB8(scuba_vlo),
        .DIB7(scuba_vlo), .DIB6(scuba_vlo), .DIB5(scuba_vlo), .DIB4(scuba_vlo),
        .DIB3(scuba_vlo), .DIB2(scuba_vlo), .DIB1(scuba_vlo), .DIB0(scuba_vlo),
        .ADB12(RdAddress[12]), .ADB11(RdAddress[11]), .ADB10(RdAddress[10]),
        .ADB9(RdAddress[9]), .ADB8(RdAddress[8]), .ADB7(RdAddress[7]), .ADB6(RdAddress[6]),
        .ADB5(RdAddress[5]), .ADB4(RdAddress[4]), .ADB3(RdAddress[3]), .ADB2(RdAddress[2]),
        .ADB1(RdAddress[1]), .ADB0(RdAddress[0]), .CEB(RdClockEn), .OCEB(RdClockEn),
        .CLKB(RdClock), .WEB(scuba_vlo), .CSB2(scuba_vlo), .CSB1(scuba_vlo),
        .CSB0(RdAddress[13]), .RSTB(Reset), .DOA8(), .DOA7(), .DOA6(), .DOA5(),
        .DOA4(), .DOA3(), .DOA2(), .DOA1(), .DOA0(), .DOB8(), .DOB7(), .DOB6(),
        .DOB5(), .DOB4(), .DOB3(), .DOB2(), .DOB1(), .DOB0(mdout1_0_4))
             /* synthesis MEM_LPC_FILE="ram.lpc" */
             /* synthesis MEM_INIT_FILE="INIT_ALL_0s" */;
    defparam ram_0_5_10.INIT_DATA = "STATIC" ;
    defparam ram_0_5_10.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam ram_0_5_10.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_5_10.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_5_10.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_5_10.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_5_10.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_5_10.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_5_10.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_5_10.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_5_10.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_5_10.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_5_10.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_5_10.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_5_10.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_5_10.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_5_10.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_5_10.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_5_10.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_5_10.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_5_10.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_5_10.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_5_10.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_5_10.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_5_10.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_5_10.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_5_10.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_5_10.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_5_10.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_5_10.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_5_10.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_5_10.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_5_10.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_5_10.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_5_10.CSDECODE_B = "0b000" ;
    defparam ram_0_5_10.CSDECODE_A = "0b000" ;
    defparam ram_0_5_10.WRITEMODE_B = "NORMAL" ;
    defparam ram_0_5_10.WRITEMODE_A = "NORMAL" ;
    defparam ram_0_5_10.GSR = "ENABLED" ;
    defparam ram_0_5_10.RESETMODE = "SYNC" ;
    defparam ram_0_5_10.REGMODE_B = "OUTREG" ;
    defparam ram_0_5_10.REGMODE_A = "OUTREG" ;
    defparam ram_0_5_10.DATA_WIDTH_B = 1 ;
    defparam ram_0_5_10.DATA_WIDTH_A = 1 ;
    DP8KC ram_0_5_10 (.DIA8(scuba_vlo), .DIA7(scuba_vlo), .DIA6(scuba_vlo),
        .DIA5(scuba_vlo), .DIA4(scuba_vlo), .DIA3(scuba_vlo), .DIA2(scuba_vlo),
        .DIA1(Data[5]), .DIA0(scuba_vlo), .ADA12(WrAddress[12]), .ADA11(WrAddress[11]),
        .ADA10(WrAddress[10]), .ADA9(WrAddress[9]), .ADA8(WrAddress[8]),
        .ADA7(WrAddress[7]), .ADA6(WrAddress[6]), .ADA5(WrAddress[5]), .ADA4(WrAddress[4]),
        .ADA3(WrAddress[3]), .ADA2(WrAddress[2]), .ADA1(WrAddress[1]), .ADA0(WrAddress[0]),
        .CEA(WrClockEn), .OCEA(WrClockEn), .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo),
        .CSA1(scuba_vlo), .CSA0(WrAddress[13]), .RSTA(Reset), .DIB8(scuba_vlo),
        .DIB7(scuba_vlo), .DIB6(scuba_vlo), .DIB5(scuba_vlo), .DIB4(scuba_vlo),
        .DIB3(scuba_vlo), .DIB2(scuba_vlo), .DIB1(scuba_vlo), .DIB0(scuba_vlo),
        .ADB12(RdAddress[12]), .ADB11(RdAddress[11]), .ADB10(RdAddress[10]),
        .ADB9(RdAddress[9]), .ADB8(RdAddress[8]), .ADB7(RdAddress[7]), .ADB6(RdAddress[6]),
        .ADB5(RdAddress[5]), .ADB4(RdAddress[4]), .ADB3(RdAddress[3]), .ADB2(RdAddress[2]),
        .ADB1(RdAddress[1]), .ADB0(RdAddress[0]), .CEB(RdClockEn), .OCEB(RdClockEn),
        .CLKB(RdClock), .WEB(scuba_vlo), .CSB2(scuba_vlo), .CSB1(scuba_vlo),
        .CSB0(RdAddress[13]), .RSTB(Reset), .DOA8(), .DOA7(), .DOA6(), .DOA5(),
        .DOA4(), .DOA3(), .DOA2(), .DOA1(), .DOA0(), .DOB8(), .DOB7(), .DOB6(),
        .DOB5(), .DOB4(), .DOB3(), .DOB2(), .DOB1(), .DOB0(mdout1_0_5))
             /* synthesis MEM_LPC_FILE="ram.lpc" */
             /* synthesis MEM_INIT_FILE="INIT_ALL_0s" */;
    defparam ram_0_6_9.INIT_DATA = "STATIC" ;
    defparam ram_0_6_9.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam ram_0_6_9.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_6_9.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_6_9.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_6_9.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_6_9.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_6_9.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_6_9.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_6_9.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_6_9.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_6_9.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_6_9.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_6_9.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_6_9.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_6_9.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_6_9.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_6_9.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_6_9.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_6_9.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_6_9.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_6_9.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_6_9.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_6_9.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_6_9.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_6_9.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_6_9.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_6_9.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_6_9.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_6_9.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_6_9.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_6_9.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_6_9.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_6_9.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_6_9.CSDECODE_B = "0b000" ;
    defparam ram_0_6_9.CSDECODE_A = "0b000" ;
    defparam ram_0_6_9.WRITEMODE_B = "NORMAL" ;
    defparam ram_0_6_9.WRITEMODE_A = "NORMAL" ;
    defparam ram_0_6_9.GSR = "ENABLED" ;
    defparam ram_0_6_9.RESETMODE = "SYNC" ;
    defparam ram_0_6_9.REGMODE_B = "OUTREG" ;
    defparam ram_0_6_9.REGMODE_A = "OUTREG" ;
    defparam ram_0_6_9.DATA_WIDTH_B = 1 ;
    defparam ram_0_6_9.DATA_WIDTH_A = 1 ;
    DP8KC ram_0_6_9 (.DIA8(scuba_vlo), .DIA7(scuba_vlo), .DIA6(scuba_vlo),
        .DIA5(scuba_vlo), .DIA4(scuba_vlo), .DIA3(scuba_vlo), .DIA2(scuba_vlo),
        .DIA1(Data[6]), .DIA0(scuba_vlo), .ADA12(WrAddress[12]), .ADA11(WrAddress[11]),
        .ADA10(WrAddress[10]), .ADA9(WrAddress[9]), .ADA8(WrAddress[8]),
        .ADA7(WrAddress[7]), .ADA6(WrAddress[6]), .ADA5(WrAddress[5]), .ADA4(WrAddress[4]),
        .ADA3(WrAddress[3]), .ADA2(WrAddress[2]), .ADA1(WrAddress[1]), .ADA0(WrAddress[0]),
        .CEA(WrClockEn), .OCEA(WrClockEn), .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo),
        .CSA1(scuba_vlo), .CSA0(WrAddress[13]), .RSTA(Reset), .DIB8(scuba_vlo),
        .DIB7(scuba_vlo), .DIB6(scuba_vlo), .DIB5(scuba_vlo), .DIB4(scuba_vlo),
        .DIB3(scuba_vlo), .DIB2(scuba_vlo), .DIB1(scuba_vlo), .DIB0(scuba_vlo),
        .ADB12(RdAddress[12]), .ADB11(RdAddress[11]), .ADB10(RdAddress[10]),
        .ADB9(RdAddress[9]), .ADB8(RdAddress[8]), .ADB7(RdAddress[7]), .ADB6(RdAddress[6]),
        .ADB5(RdAddress[5]), .ADB4(RdAddress[4]), .ADB3(RdAddress[3]), .ADB2(RdAddress[2]),
        .ADB1(RdAddress[1]), .ADB0(RdAddress[0]), .CEB(RdClockEn), .OCEB(RdClockEn),
        .CLKB(RdClock), .WEB(scuba_vlo), .CSB2(scuba_vlo), .CSB1(scuba_vlo),
        .CSB0(RdAddress[13]), .RSTB(Reset), .DOA8(), .DOA7(), .DOA6(), .DOA5(),
        .DOA4(), .DOA3(), .DOA2(), .DOA1(), .DOA0(), .DOB8(), .DOB7(), .DOB6(),
        .DOB5(), .DOB4(), .DOB3(), .DOB2(), .DOB1(), .DOB0(mdout1_0_6))
             /* synthesis MEM_LPC_FILE="ram.lpc" */
             /* synthesis MEM_INIT_FILE="INIT_ALL_0s" */;
    defparam ram_0_7_8.INIT_DATA = "STATIC" ;
    defparam ram_0_7_8.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam ram_0_7_8.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_7_8.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_7_8.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_7_8.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_7_8.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_7_8.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_7_8.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_7_8.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_7_8.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_7_8.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_7_8.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_7_8.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_7_8.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_7_8.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_7_8.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_7_8.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_7_8.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_7_8.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_7_8.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_7_8.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_7_8.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_7_8.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_7_8.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_7_8.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_7_8.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_7_8.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_7_8.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_7_8.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_7_8.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_7_8.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_7_8.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_7_8.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_0_7_8.CSDECODE_B = "0b000" ;
    defparam ram_0_7_8.CSDECODE_A = "0b000" ;
    defparam ram_0_7_8.WRITEMODE_B = "NORMAL" ;
    defparam ram_0_7_8.WRITEMODE_A = "NORMAL" ;
    defparam ram_0_7_8.GSR = "ENABLED" ;
    defparam ram_0_7_8.RESETMODE = "SYNC" ;
    defparam ram_0_7_8.REGMODE_B = "OUTREG" ;
    defparam ram_0_7_8.REGMODE_A = "OUTREG" ;
    defparam ram_0_7_8.DATA_WIDTH_B = 1 ;
    defparam ram_0_7_8.DATA_WIDTH_A = 1 ;
    DP8KC ram_0_7_8 (.DIA8(scuba_vlo), .DIA7(scuba_vlo), .DIA6(scuba_vlo),
        .DIA5(scuba_vlo), .DIA4(scuba_vlo), .DIA3(scuba_vlo), .DIA2(scuba_vlo),
        .DIA1(Data[7]), .DIA0(scuba_vlo), .ADA12(WrAddress[12]), .ADA11(WrAddress[11]),
        .ADA10(WrAddress[10]), .ADA9(WrAddress[9]), .ADA8(WrAddress[8]),
        .ADA7(WrAddress[7]), .ADA6(WrAddress[6]), .ADA5(WrAddress[5]), .ADA4(WrAddress[4]),
        .ADA3(WrAddress[3]), .ADA2(WrAddress[2]), .ADA1(WrAddress[1]), .ADA0(WrAddress[0]),
        .CEA(WrClockEn), .OCEA(WrClockEn), .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo),
        .CSA1(scuba_vlo), .CSA0(WrAddress[13]), .RSTA(Reset), .DIB8(scuba_vlo),
        .DIB7(scuba_vlo), .DIB6(scuba_vlo), .DIB5(scuba_vlo), .DIB4(scuba_vlo),
        .DIB3(scuba_vlo), .DIB2(scuba_vlo), .DIB1(scuba_vlo), .DIB0(scuba_vlo),
        .ADB12(RdAddress[12]), .ADB11(RdAddress[11]), .ADB10(RdAddress[10]),
        .ADB9(RdAddress[9]), .ADB8(RdAddress[8]), .ADB7(RdAddress[7]), .ADB6(RdAddress[6]),
        .ADB5(RdAddress[5]), .ADB4(RdAddress[4]), .ADB3(RdAddress[3]), .ADB2(RdAddress[2]),
        .ADB1(RdAddress[1]), .ADB0(RdAddress[0]), .CEB(RdClockEn), .OCEB(RdClockEn),
        .CLKB(RdClock), .WEB(scuba_vlo), .CSB2(scuba_vlo), .CSB1(scuba_vlo),
        .CSB0(RdAddress[13]), .RSTB(Reset), .DOA8(), .DOA7(), .DOA6(), .DOA5(),
        .DOA4(), .DOA3(), .DOA2(), .DOA1(), .DOA0(), .DOB8(), .DOB7(), .DOB6(),
        .DOB5(), .DOB4(), .DOB3(), .DOB2(), .DOB1(), .DOB0(mdout1_0_7))
             /* synthesis MEM_LPC_FILE="ram.lpc" */
             /* synthesis MEM_INIT_FILE="INIT_ALL_0s" */;
    defparam ram_1_0_7.INIT_DATA = "STATIC" ;
    defparam ram_1_0_7.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam ram_1_0_7.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_0_7.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_0_7.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_0_7.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_0_7.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_0_7.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_0_7.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_0_7.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_0_7.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_0_7.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_0_7.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_0_7.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_0_7.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_0_7.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_0_7.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_0_7.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_0_7.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_0_7.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_0_7.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_0_7.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_0_7.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_0_7.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_0_7.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_0_7.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_0_7.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_0_7.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_0_7.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_0_7.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_0_7.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_0_7.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_0_7.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_0_7.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_0_7.CSDECODE_B = "0b001" ;
    defparam ram_1_0_7.CSDECODE_A = "0b001" ;
    defparam ram_1_0_7.WRITEMODE_B = "NORMAL" ;
    defparam ram_1_0_7.WRITEMODE_A = "NORMAL" ;
    defparam ram_1_0_7.GSR = "ENABLED" ;
    defparam ram_1_0_7.RESETMODE = "SYNC" ;
    defparam ram_1_0_7.REGMODE_B = "OUTREG" ;
    defparam ram_1_0_7.REGMODE_A = "OUTREG" ;
    defparam ram_1_0_7.DATA_WIDTH_B = 1 ;
    defparam ram_1_0_7.DATA_WIDTH_A = 1 ;
    DP8KC ram_1_0_7 (.DIA8(scuba_vlo), .DIA7(scuba_vlo), .DIA6(scuba_vlo),
        .DIA5(scuba_vlo), .DIA4(scuba_vlo), .DIA3(scuba_vlo), .DIA2(scuba_vlo),
        .DIA1(Data[0]), .DIA0(scuba_vlo), .ADA12(WrAddress[12]), .ADA11(WrAddress[11]),
        .ADA10(WrAddress[10]), .ADA9(WrAddress[9]), .ADA8(WrAddress[8]),
        .ADA7(WrAddress[7]), .ADA6(WrAddress[6]), .ADA5(WrAddress[5]), .ADA4(WrAddress[4]),
        .ADA3(WrAddress[3]), .ADA2(WrAddress[2]), .ADA1(WrAddress[1]), .ADA0(WrAddress[0]),
        .CEA(WrClockEn), .OCEA(WrClockEn), .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo),
        .CSA1(scuba_vlo), .CSA0(WrAddress[13]), .RSTA(Reset), .DIB8(scuba_vlo),
        .DIB7(scuba_vlo), .DIB6(scuba_vlo), .DIB5(scuba_vlo), .DIB4(scuba_vlo),
        .DIB3(scuba_vlo), .DIB2(scuba_vlo), .DIB1(scuba_vlo), .DIB0(scuba_vlo),
        .ADB12(RdAddress[12]), .ADB11(RdAddress[11]), .ADB10(RdAddress[10]),
        .ADB9(RdAddress[9]), .ADB8(RdAddress[8]), .ADB7(RdAddress[7]), .ADB6(RdAddress[6]),
        .ADB5(RdAddress[5]), .ADB4(RdAddress[4]), .ADB3(RdAddress[3]), .ADB2(RdAddress[2]),
        .ADB1(RdAddress[1]), .ADB0(RdAddress[0]), .CEB(RdClockEn), .OCEB(RdClockEn),
        .CLKB(RdClock), .WEB(scuba_vlo), .CSB2(scuba_vlo), .CSB1(scuba_vlo),
        .CSB0(RdAddress[13]), .RSTB(Reset), .DOA8(), .DOA7(), .DOA6(), .DOA5(),
        .DOA4(), .DOA3(), .DOA2(), .DOA1(), .DOA0(), .DOB8(), .DOB7(), .DOB6(),
        .DOB5(), .DOB4(), .DOB3(), .DOB2(), .DOB1(), .DOB0(mdout1_1_0))
             /* synthesis MEM_LPC_FILE="ram.lpc" */
             /* synthesis MEM_INIT_FILE="INIT_ALL_0s" */;
    defparam ram_1_1_6.INIT_DATA = "STATIC" ;
    defparam ram_1_1_6.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam ram_1_1_6.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_1_6.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_1_6.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_1_6.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_1_6.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_1_6.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_1_6.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_1_6.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_1_6.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_1_6.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_1_6.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_1_6.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_1_6.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_1_6.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_1_6.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_1_6.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_1_6.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_1_6.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_1_6.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_1_6.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_1_6.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_1_6.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_1_6.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_1_6.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_1_6.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_1_6.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_1_6.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_1_6.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_1_6.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_1_6.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_1_6.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_1_6.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_1_6.CSDECODE_B = "0b001" ;
    defparam ram_1_1_6.CSDECODE_A = "0b001" ;
    defparam ram_1_1_6.WRITEMODE_B = "NORMAL" ;
    defparam ram_1_1_6.WRITEMODE_A = "NORMAL" ;
    defparam ram_1_1_6.GSR = "ENABLED" ;
    defparam ram_1_1_6.RESETMODE = "SYNC" ;
    defparam ram_1_1_6.REGMODE_B = "OUTREG" ;
    defparam ram_1_1_6.REGMODE_A = "OUTREG" ;
    defparam ram_1_1_6.DATA_WIDTH_B = 1 ;
    defparam ram_1_1_6.DATA_WIDTH_A = 1 ;
    DP8KC ram_1_1_6 (.DIA8(scuba_vlo), .DIA7(scuba_vlo), .DIA6(scuba_vlo),
        .DIA5(scuba_vlo), .DIA4(scuba_vlo), .DIA3(scuba_vlo), .DIA2(scuba_vlo),
        .DIA1(Data[1]), .DIA0(scuba_vlo), .ADA12(WrAddress[12]), .ADA11(WrAddress[11]),
        .ADA10(WrAddress[10]), .ADA9(WrAddress[9]), .ADA8(WrAddress[8]),
        .ADA7(WrAddress[7]), .ADA6(WrAddress[6]), .ADA5(WrAddress[5]), .ADA4(WrAddress[4]),
        .ADA3(WrAddress[3]), .ADA2(WrAddress[2]), .ADA1(WrAddress[1]), .ADA0(WrAddress[0]),
        .CEA(WrClockEn), .OCEA(WrClockEn), .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo),
        .CSA1(scuba_vlo), .CSA0(WrAddress[13]), .RSTA(Reset), .DIB8(scuba_vlo),
        .DIB7(scuba_vlo), .DIB6(scuba_vlo), .DIB5(scuba_vlo), .DIB4(scuba_vlo),
        .DIB3(scuba_vlo), .DIB2(scuba_vlo), .DIB1(scuba_vlo), .DIB0(scuba_vlo),
        .ADB12(RdAddress[12]), .ADB11(RdAddress[11]), .ADB10(RdAddress[10]),
        .ADB9(RdAddress[9]), .ADB8(RdAddress[8]), .ADB7(RdAddress[7]), .ADB6(RdAddress[6]),
        .ADB5(RdAddress[5]), .ADB4(RdAddress[4]), .ADB3(RdAddress[3]), .ADB2(RdAddress[2]),
        .ADB1(RdAddress[1]), .ADB0(RdAddress[0]), .CEB(RdClockEn), .OCEB(RdClockEn),
        .CLKB(RdClock), .WEB(scuba_vlo), .CSB2(scuba_vlo), .CSB1(scuba_vlo),
        .CSB0(RdAddress[13]), .RSTB(Reset), .DOA8(), .DOA7(), .DOA6(), .DOA5(),
        .DOA4(), .DOA3(), .DOA2(), .DOA1(), .DOA0(), .DOB8(), .DOB7(), .DOB6(),
        .DOB5(), .DOB4(), .DOB3(), .DOB2(), .DOB1(), .DOB0(mdout1_1_1))
             /* synthesis MEM_LPC_FILE="ram.lpc" */
             /* synthesis MEM_INIT_FILE="INIT_ALL_0s" */;
    defparam ram_1_2_5.INIT_DATA = "STATIC" ;
    defparam ram_1_2_5.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam ram_1_2_5.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_2_5.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_2_5.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_2_5.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_2_5.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_2_5.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_2_5.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_2_5.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_2_5.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_2_5.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_2_5.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_2_5.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_2_5.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_2_5.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_2_5.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_2_5.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_2_5.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_2_5.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_2_5.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_2_5.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_2_5.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_2_5.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_2_5.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_2_5.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_2_5.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_2_5.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_2_5.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_2_5.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_2_5.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_2_5.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_2_5.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_2_5.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_2_5.CSDECODE_B = "0b001" ;
    defparam ram_1_2_5.CSDECODE_A = "0b001" ;
    defparam ram_1_2_5.WRITEMODE_B = "NORMAL" ;
    defparam ram_1_2_5.WRITEMODE_A = "NORMAL" ;
    defparam ram_1_2_5.GSR = "ENABLED" ;
    defparam ram_1_2_5.RESETMODE = "SYNC" ;
    defparam ram_1_2_5.REGMODE_B = "OUTREG" ;
    defparam ram_1_2_5.REGMODE_A = "OUTREG" ;
    defparam ram_1_2_5.DATA_WIDTH_B = 1 ;
    defparam ram_1_2_5.DATA_WIDTH_A = 1 ;
    DP8KC ram_1_2_5 (.DIA8(scuba_vlo), .DIA7(scuba_vlo), .DIA6(scuba_vlo),
        .DIA5(scuba_vlo), .DIA4(scuba_vlo), .DIA3(scuba_vlo), .DIA2(scuba_vlo),
        .DIA1(Data[2]), .DIA0(scuba_vlo), .ADA12(WrAddress[12]), .ADA11(WrAddress[11]),
        .ADA10(WrAddress[10]), .ADA9(WrAddress[9]), .ADA8(WrAddress[8]),
        .ADA7(WrAddress[7]), .ADA6(WrAddress[6]), .ADA5(WrAddress[5]), .ADA4(WrAddress[4]),
        .ADA3(WrAddress[3]), .ADA2(WrAddress[2]), .ADA1(WrAddress[1]), .ADA0(WrAddress[0]),
        .CEA(WrClockEn), .OCEA(WrClockEn), .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo),
        .CSA1(scuba_vlo), .CSA0(WrAddress[13]), .RSTA(Reset), .DIB8(scuba_vlo),
        .DIB7(scuba_vlo), .DIB6(scuba_vlo), .DIB5(scuba_vlo), .DIB4(scuba_vlo),
        .DIB3(scuba_vlo), .DIB2(scuba_vlo), .DIB1(scuba_vlo), .DIB0(scuba_vlo),
        .ADB12(RdAddress[12]), .ADB11(RdAddress[11]), .ADB10(RdAddress[10]),
        .ADB9(RdAddress[9]), .ADB8(RdAddress[8]), .ADB7(RdAddress[7]), .ADB6(RdAddress[6]),
        .ADB5(RdAddress[5]), .ADB4(RdAddress[4]), .ADB3(RdAddress[3]), .ADB2(RdAddress[2]),
        .ADB1(RdAddress[1]), .ADB0(RdAddress[0]), .CEB(RdClockEn), .OCEB(RdClockEn),
        .CLKB(RdClock), .WEB(scuba_vlo), .CSB2(scuba_vlo), .CSB1(scuba_vlo),
        .CSB0(RdAddress[13]), .RSTB(Reset), .DOA8(), .DOA7(), .DOA6(), .DOA5(),
        .DOA4(), .DOA3(), .DOA2(), .DOA1(), .DOA0(), .DOB8(), .DOB7(), .DOB6(),
        .DOB5(), .DOB4(), .DOB3(), .DOB2(), .DOB1(), .DOB0(mdout1_1_2))
             /* synthesis MEM_LPC_FILE="ram.lpc" */
             /* synthesis MEM_INIT_FILE="INIT_ALL_0s" */;
    defparam ram_1_3_4.INIT_DATA = "STATIC" ;
    defparam ram_1_3_4.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam ram_1_3_4.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_3_4.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_3_4.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_3_4.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_3_4.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_3_4.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_3_4.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_3_4.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_3_4.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_3_4.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_3_4.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_3_4.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_3_4.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_3_4.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_3_4.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_3_4.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_3_4.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_3_4.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_3_4.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_3_4.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_3_4.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_3_4.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_3_4.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_3_4.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_3_4.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_3_4.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_3_4.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_3_4.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_3_4.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_3_4.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_3_4.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_3_4.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_3_4.CSDECODE_B = "0b001" ;
    defparam ram_1_3_4.CSDECODE_A = "0b001" ;
    defparam ram_1_3_4.WRITEMODE_B = "NORMAL" ;
    defparam ram_1_3_4.WRITEMODE_A = "NORMAL" ;
    defparam ram_1_3_4.GSR = "ENABLED" ;
    defparam ram_1_3_4.RESETMODE = "SYNC" ;
    defparam ram_1_3_4.REGMODE_B = "OUTREG" ;
    defparam ram_1_3_4.REGMODE_A = "OUTREG" ;
    defparam ram_1_3_4.DATA_WIDTH_B = 1 ;
    defparam ram_1_3_4.DATA_WIDTH_A = 1 ;
    DP8KC ram_1_3_4 (.DIA8(scuba_vlo), .DIA7(scuba_vlo), .DIA6(scuba_vlo),
        .DIA5(scuba_vlo), .DIA4(scuba_vlo), .DIA3(scuba_vlo), .DIA2(scuba_vlo),
        .DIA1(Data[3]), .DIA0(scuba_vlo), .ADA12(WrAddress[12]), .ADA11(WrAddress[11]),
        .ADA10(WrAddress[10]), .ADA9(WrAddress[9]), .ADA8(WrAddress[8]),
        .ADA7(WrAddress[7]), .ADA6(WrAddress[6]), .ADA5(WrAddress[5]), .ADA4(WrAddress[4]),
        .ADA3(WrAddress[3]), .ADA2(WrAddress[2]), .ADA1(WrAddress[1]), .ADA0(WrAddress[0]),
        .CEA(WrClockEn), .OCEA(WrClockEn), .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo),
        .CSA1(scuba_vlo), .CSA0(WrAddress[13]), .RSTA(Reset), .DIB8(scuba_vlo),
        .DIB7(scuba_vlo), .DIB6(scuba_vlo), .DIB5(scuba_vlo), .DIB4(scuba_vlo),
        .DIB3(scuba_vlo), .DIB2(scuba_vlo), .DIB1(scuba_vlo), .DIB0(scuba_vlo),
        .ADB12(RdAddress[12]), .ADB11(RdAddress[11]), .ADB10(RdAddress[10]),
        .ADB9(RdAddress[9]), .ADB8(RdAddress[8]), .ADB7(RdAddress[7]), .ADB6(RdAddress[6]),
        .ADB5(RdAddress[5]), .ADB4(RdAddress[4]), .ADB3(RdAddress[3]), .ADB2(RdAddress[2]),
        .ADB1(RdAddress[1]), .ADB0(RdAddress[0]), .CEB(RdClockEn), .OCEB(RdClockEn),
        .CLKB(RdClock), .WEB(scuba_vlo), .CSB2(scuba_vlo), .CSB1(scuba_vlo),
        .CSB0(RdAddress[13]), .RSTB(Reset), .DOA8(), .DOA7(), .DOA6(), .DOA5(),
        .DOA4(), .DOA3(), .DOA2(), .DOA1(), .DOA0(), .DOB8(), .DOB7(), .DOB6(),
        .DOB5(), .DOB4(), .DOB3(), .DOB2(), .DOB1(), .DOB0(mdout1_1_3))
             /* synthesis MEM_LPC_FILE="ram.lpc" */
             /* synthesis MEM_INIT_FILE="INIT_ALL_0s" */;
    defparam ram_1_4_3.INIT_DATA = "STATIC" ;
    defparam ram_1_4_3.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam ram_1_4_3.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_4_3.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_4_3.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_4_3.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_4_3.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_4_3.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_4_3.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_4_3.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_4_3.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_4_3.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_4_3.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_4_3.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_4_3.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_4_3.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_4_3.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_4_3.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_4_3.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_4_3.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_4_3.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_4_3.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_4_3.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_4_3.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_4_3.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_4_3.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_4_3.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_4_3.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_4_3.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_4_3.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_4_3.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_4_3.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_4_3.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_4_3.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_4_3.CSDECODE_B = "0b001" ;
    defparam ram_1_4_3.CSDECODE_A = "0b001" ;
    defparam ram_1_4_3.WRITEMODE_B = "NORMAL" ;
    defparam ram_1_4_3.WRITEMODE_A = "NORMAL" ;
    defparam ram_1_4_3.GSR = "ENABLED" ;
    defparam ram_1_4_3.RESETMODE = "SYNC" ;
    defparam ram_1_4_3.REGMODE_B = "OUTREG" ;
    defparam ram_1_4_3.REGMODE_A = "OUTREG" ;
    defparam ram_1_4_3.DATA_WIDTH_B = 1 ;
    defparam ram_1_4_3.DATA_WIDTH_A = 1 ;
    DP8KC ram_1_4_3 (.DIA8(scuba_vlo), .DIA7(scuba_vlo), .DIA6(scuba_vlo),
        .DIA5(scuba_vlo), .DIA4(scuba_vlo), .DIA3(scuba_vlo), .DIA2(scuba_vlo),
        .DIA1(Data[4]), .DIA0(scuba_vlo), .ADA12(WrAddress[12]), .ADA11(WrAddress[11]),
        .ADA10(WrAddress[10]), .ADA9(WrAddress[9]), .ADA8(WrAddress[8]),
        .ADA7(WrAddress[7]), .ADA6(WrAddress[6]), .ADA5(WrAddress[5]), .ADA4(WrAddress[4]),
        .ADA3(WrAddress[3]), .ADA2(WrAddress[2]), .ADA1(WrAddress[1]), .ADA0(WrAddress[0]),
        .CEA(WrClockEn), .OCEA(WrClockEn), .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo),
        .CSA1(scuba_vlo), .CSA0(WrAddress[13]), .RSTA(Reset), .DIB8(scuba_vlo),
        .DIB7(scuba_vlo), .DIB6(scuba_vlo), .DIB5(scuba_vlo), .DIB4(scuba_vlo),
        .DIB3(scuba_vlo), .DIB2(scuba_vlo), .DIB1(scuba_vlo), .DIB0(scuba_vlo),
        .ADB12(RdAddress[12]), .ADB11(RdAddress[11]), .ADB10(RdAddress[10]),
        .ADB9(RdAddress[9]), .ADB8(RdAddress[8]), .ADB7(RdAddress[7]), .ADB6(RdAddress[6]),
        .ADB5(RdAddress[5]), .ADB4(RdAddress[4]), .ADB3(RdAddress[3]), .ADB2(RdAddress[2]),
        .ADB1(RdAddress[1]), .ADB0(RdAddress[0]), .CEB(RdClockEn), .OCEB(RdClockEn),
        .CLKB(RdClock), .WEB(scuba_vlo), .CSB2(scuba_vlo), .CSB1(scuba_vlo),
        .CSB0(RdAddress[13]), .RSTB(Reset), .DOA8(), .DOA7(), .DOA6(), .DOA5(),
        .DOA4(), .DOA3(), .DOA2(), .DOA1(), .DOA0(), .DOB8(), .DOB7(), .DOB6(),
        .DOB5(), .DOB4(), .DOB3(), .DOB2(), .DOB1(), .DOB0(mdout1_1_4))
             /* synthesis MEM_LPC_FILE="ram.lpc" */
             /* synthesis MEM_INIT_FILE="INIT_ALL_0s" */;
    defparam ram_1_5_2.INIT_DATA = "STATIC" ;
    defparam ram_1_5_2.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam ram_1_5_2.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_5_2.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_5_2.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_5_2.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_5_2.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_5_2.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_5_2.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_5_2.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_5_2.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_5_2.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_5_2.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_5_2.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_5_2.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_5_2.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_5_2.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_5_2.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_5_2.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_5_2.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_5_2.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_5_2.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_5_2.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_5_2.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_5_2.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_5_2.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_5_2.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_5_2.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_5_2.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_5_2.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_5_2.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_5_2.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_5_2.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_5_2.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_5_2.CSDECODE_B = "0b001" ;
    defparam ram_1_5_2.CSDECODE_A = "0b001" ;
    defparam ram_1_5_2.WRITEMODE_B = "NORMAL" ;
    defparam ram_1_5_2.WRITEMODE_A = "NORMAL" ;
    defparam ram_1_5_2.GSR = "ENABLED" ;
    defparam ram_1_5_2.RESETMODE = "SYNC" ;
    defparam ram_1_5_2.REGMODE_B = "OUTREG" ;
    defparam ram_1_5_2.REGMODE_A = "OUTREG" ;
    defparam ram_1_5_2.DATA_WIDTH_B = 1 ;
    defparam ram_1_5_2.DATA_WIDTH_A = 1 ;
    DP8KC ram_1_5_2 (.DIA8(scuba_vlo), .DIA7(scuba_vlo), .DIA6(scuba_vlo),
        .DIA5(scuba_vlo), .DIA4(scuba_vlo), .DIA3(scuba_vlo), .DIA2(scuba_vlo),
        .DIA1(Data[5]), .DIA0(scuba_vlo), .ADA12(WrAddress[12]), .ADA11(WrAddress[11]),
        .ADA10(WrAddress[10]), .ADA9(WrAddress[9]), .ADA8(WrAddress[8]),
        .ADA7(WrAddress[7]), .ADA6(WrAddress[6]), .ADA5(WrAddress[5]), .ADA4(WrAddress[4]),
        .ADA3(WrAddress[3]), .ADA2(WrAddress[2]), .ADA1(WrAddress[1]), .ADA0(WrAddress[0]),
        .CEA(WrClockEn), .OCEA(WrClockEn), .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo),
        .CSA1(scuba_vlo), .CSA0(WrAddress[13]), .RSTA(Reset), .DIB8(scuba_vlo),
        .DIB7(scuba_vlo), .DIB6(scuba_vlo), .DIB5(scuba_vlo), .DIB4(scuba_vlo),
        .DIB3(scuba_vlo), .DIB2(scuba_vlo), .DIB1(scuba_vlo), .DIB0(scuba_vlo),
        .ADB12(RdAddress[12]), .ADB11(RdAddress[11]), .ADB10(RdAddress[10]),
        .ADB9(RdAddress[9]), .ADB8(RdAddress[8]), .ADB7(RdAddress[7]), .ADB6(RdAddress[6]),
        .ADB5(RdAddress[5]), .ADB4(RdAddress[4]), .ADB3(RdAddress[3]), .ADB2(RdAddress[2]),
        .ADB1(RdAddress[1]), .ADB0(RdAddress[0]), .CEB(RdClockEn), .OCEB(RdClockEn),
        .CLKB(RdClock), .WEB(scuba_vlo), .CSB2(scuba_vlo), .CSB1(scuba_vlo),
        .CSB0(RdAddress[13]), .RSTB(Reset), .DOA8(), .DOA7(), .DOA6(), .DOA5(),
        .DOA4(), .DOA3(), .DOA2(), .DOA1(), .DOA0(), .DOB8(), .DOB7(), .DOB6(),
        .DOB5(), .DOB4(), .DOB3(), .DOB2(), .DOB1(), .DOB0(mdout1_1_5))
             /* synthesis MEM_LPC_FILE="ram.lpc" */
             /* synthesis MEM_INIT_FILE="INIT_ALL_0s" */;
    defparam ram_1_6_1.INIT_DATA = "STATIC" ;
    defparam ram_1_6_1.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam ram_1_6_1.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_6_1.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_6_1.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_6_1.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_6_1.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_6_1.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_6_1.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_6_1.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_6_1.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_6_1.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_6_1.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_6_1.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_6_1.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_6_1.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_6_1.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_6_1.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_6_1.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_6_1.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_6_1.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_6_1.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_6_1.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_6_1.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_6_1.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_6_1.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_6_1.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_6_1.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_6_1.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_6_1.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_6_1.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_6_1.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_6_1.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_6_1.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_6_1.CSDECODE_B = "0b001" ;
    defparam ram_1_6_1.CSDECODE_A = "0b001" ;
    defparam ram_1_6_1.WRITEMODE_B = "NORMAL" ;
    defparam ram_1_6_1.WRITEMODE_A = "NORMAL" ;
    defparam ram_1_6_1.GSR = "ENABLED" ;
    defparam ram_1_6_1.RESETMODE = "SYNC" ;
    defparam ram_1_6_1.REGMODE_B = "OUTREG" ;
    defparam ram_1_6_1.REGMODE_A = "OUTREG" ;
    defparam ram_1_6_1.DATA_WIDTH_B = 1 ;
    defparam ram_1_6_1.DATA_WIDTH_A = 1 ;
    DP8KC ram_1_6_1 (.DIA8(scuba_vlo), .DIA7(scuba_vlo), .DIA6(scuba_vlo),
        .DIA5(scuba_vlo), .DIA4(scuba_vlo), .DIA3(scuba_vlo), .DIA2(scuba_vlo),
        .DIA1(Data[6]), .DIA0(scuba_vlo), .ADA12(WrAddress[12]), .ADA11(WrAddress[11]),
        .ADA10(WrAddress[10]), .ADA9(WrAddress[9]), .ADA8(WrAddress[8]),
        .ADA7(WrAddress[7]), .ADA6(WrAddress[6]), .ADA5(WrAddress[5]), .ADA4(WrAddress[4]),
        .ADA3(WrAddress[3]), .ADA2(WrAddress[2]), .ADA1(WrAddress[1]), .ADA0(WrAddress[0]),
        .CEA(WrClockEn), .OCEA(WrClockEn), .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo),
        .CSA1(scuba_vlo), .CSA0(WrAddress[13]), .RSTA(Reset), .DIB8(scuba_vlo),
        .DIB7(scuba_vlo), .DIB6(scuba_vlo), .DIB5(scuba_vlo), .DIB4(scuba_vlo),
        .DIB3(scuba_vlo), .DIB2(scuba_vlo), .DIB1(scuba_vlo), .DIB0(scuba_vlo),
        .ADB12(RdAddress[12]), .ADB11(RdAddress[11]), .ADB10(RdAddress[10]),
        .ADB9(RdAddress[9]), .ADB8(RdAddress[8]), .ADB7(RdAddress[7]), .ADB6(RdAddress[6]),
        .ADB5(RdAddress[5]), .ADB4(RdAddress[4]), .ADB3(RdAddress[3]), .ADB2(RdAddress[2]),
        .ADB1(RdAddress[1]), .ADB0(RdAddress[0]), .CEB(RdClockEn), .OCEB(RdClockEn),
        .CLKB(RdClock), .WEB(scuba_vlo), .CSB2(scuba_vlo), .CSB1(scuba_vlo),
        .CSB0(RdAddress[13]), .RSTB(Reset), .DOA8(), .DOA7(), .DOA6(), .DOA5(),
        .DOA4(), .DOA3(), .DOA2(), .DOA1(), .DOA0(), .DOB8(), .DOB7(), .DOB6(),
        .DOB5(), .DOB4(), .DOB3(), .DOB2(), .DOB1(), .DOB0(mdout1_1_6))
             /* synthesis MEM_LPC_FILE="ram.lpc" */
             /* synthesis MEM_INIT_FILE="INIT_ALL_0s" */;
    defparam ram_1_7_0.INIT_DATA = "STATIC" ;
    defparam ram_1_7_0.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam ram_1_7_0.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_7_0.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_7_0.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_7_0.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_7_0.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_7_0.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_7_0.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_7_0.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_7_0.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_7_0.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_7_0.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_7_0.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_7_0.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_7_0.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_7_0.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_7_0.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_7_0.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_7_0.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_7_0.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_7_0.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_7_0.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_7_0.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_7_0.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_7_0.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_7_0.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_7_0.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_7_0.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_7_0.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_7_0.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_7_0.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_7_0.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_7_0.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram_1_7_0.CSDECODE_B = "0b001" ;
    defparam ram_1_7_0.CSDECODE_A = "0b001" ;
    defparam ram_1_7_0.WRITEMODE_B = "NORMAL" ;
    defparam ram_1_7_0.WRITEMODE_A = "NORMAL" ;
    defparam ram_1_7_0.GSR = "ENABLED" ;
    defparam ram_1_7_0.RESETMODE = "SYNC" ;
    defparam ram_1_7_0.REGMODE_B = "OUTREG" ;
    defparam ram_1_7_0.REGMODE_A = "OUTREG" ;
    defparam ram_1_7_0.DATA_WIDTH_B = 1 ;
    defparam ram_1_7_0.DATA_WIDTH_A = 1 ;
    DP8KC ram_1_7_0 (.DIA8(scuba_vlo), .DIA7(scuba_vlo), .DIA6(scuba_vlo),
        .DIA5(scuba_vlo), .DIA4(scuba_vlo), .DIA3(scuba_vlo), .DIA2(scuba_vlo),
        .DIA1(Data[7]), .DIA0(scuba_vlo), .ADA12(WrAddress[12]), .ADA11(WrAddress[11]),
        .ADA10(WrAddress[10]), .ADA9(WrAddress[9]), .ADA8(WrAddress[8]),
        .ADA7(WrAddress[7]), .ADA6(WrAddress[6]), .ADA5(WrAddress[5]), .ADA4(WrAddress[4]),
        .ADA3(WrAddress[3]), .ADA2(WrAddress[2]), .ADA1(WrAddress[1]), .ADA0(WrAddress[0]),
        .CEA(WrClockEn), .OCEA(WrClockEn), .CLKA(WrClock), .WEA(WE), .CSA2(scuba_vlo),
        .CSA1(scuba_vlo), .CSA0(WrAddress[13]), .RSTA(Reset), .DIB8(scuba_vlo),
        .DIB7(scuba_vlo), .DIB6(scuba_vlo), .DIB5(scuba_vlo), .DIB4(scuba_vlo),
        .DIB3(scuba_vlo), .DIB2(scuba_vlo), .DIB1(scuba_vlo), .DIB0(scuba_vlo),
        .ADB12(RdAddress[12]), .ADB11(RdAddress[11]), .ADB10(RdAddress[10]),
        .ADB9(RdAddress[9]), .ADB8(RdAddress[8]), .ADB7(RdAddress[7]), .ADB6(RdAddress[6]),
        .ADB5(RdAddress[5]), .ADB4(RdAddress[4]), .ADB3(RdAddress[3]), .ADB2(RdAddress[2]),
        .ADB1(RdAddress[1]), .ADB0(RdAddress[0]), .CEB(RdClockEn), .OCEB(RdClockEn),
        .CLKB(RdClock), .WEB(scuba_vlo), .CSB2(scuba_vlo), .CSB1(scuba_vlo),
        .CSB0(RdAddress[13]), .RSTB(Reset), .DOA8(), .DOA7(), .DOA6(), .DOA5(),
        .DOA4(), .DOA3(), .DOA2(), .DOA1(), .DOA0(), .DOB8(), .DOB7(), .DOB6(),
        .DOB5(), .DOB4(), .DOB3(), .DOB2(), .DOB1(), .DOB0(mdout1_1_7))
             /* synthesis MEM_LPC_FILE="ram.lpc" */
             /* synthesis MEM_INIT_FILE="INIT_ALL_0s" */;
    FD1P3DX FF_1 (.D(RdAddress[13]), .SP(RdClockEn), .CK(RdClock), .CD(scuba_vlo),
        .Q(raddr13_ff))
             /* synthesis GSR="ENABLED" */;
    VLO scuba_vlo_inst (.Z(scuba_vlo));
    FD1P3DX FF_0 (.D(raddr13_ff), .SP(RdClockEn), .CK(RdClock), .CD(scuba_vlo),
        .Q(raddr13_ff2))
             /* synthesis GSR="ENABLED" */;
    MUX21 mux_7 (.D0(mdout1_0_0), .D1(mdout1_1_0), .SD(raddr13_ff2), .Z(Q[0]));
    MUX21 mux_6 (.D0(mdout1_0_1), .D1(mdout1_1_1), .SD(raddr13_ff2), .Z(Q[1]));
    MUX21 mux_5 (.D0(mdout1_0_2), .D1(mdout1_1_2), .SD(raddr13_ff2), .Z(Q[2]));
    MUX21 mux_4 (.D0(mdout1_0_3), .D1(mdout1_1_3), .SD(raddr13_ff2), .Z(Q[3]));
    MUX21 mux_3 (.D0(mdout1_0_4), .D1(mdout1_1_4), .SD(raddr13_ff2), .Z(Q[4]));
    MUX21 mux_2 (.D0(mdout1_0_5), .D1(mdout1_1_5), .SD(raddr13_ff2), .Z(Q[5]));
    MUX21 mux_1 (.D0(mdout1_0_6), .D1(mdout1_1_6), .SD(raddr13_ff2), .Z(Q[6]));
    MUX21 mux_0 (.D0(mdout1_0_7), .D1(mdout1_1_7), .SD(raddr13_ff2), .Z(Q[7]));
    // exemplar begin
    // exemplar attribute ram_0_0_15 MEM_LPC_FILE ram.lpc
    // exemplar attribute ram_0_0_15 MEM_INIT_FILE INIT_ALL_0s
    // exemplar attribute ram_0_1_14 MEM_LPC_FILE ram.lpc
    // exemplar attribute ram_0_1_14 MEM_INIT_FILE INIT_ALL_0s
    // exemplar attribute ram_0_2_13 MEM_LPC_FILE ram.lpc
    // exemplar attribute ram_0_2_13 MEM_INIT_FILE INIT_ALL_0s
    // exemplar attribute ram_0_3_12 MEM_LPC_FILE ram.lpc
    // exemplar attribute ram_0_3_12 MEM_INIT_FILE INIT_ALL_0s
    // exemplar attribute ram_0_4_11 MEM_LPC_FILE ram.lpc
    // exemplar attribute ram_0_4_11 MEM_INIT_FILE INIT_ALL_0s
    // exemplar attribute ram_0_5_10 MEM_LPC_FILE ram.lpc
    // exemplar attribute ram_0_5_10 MEM_INIT_FILE INIT_ALL_0s
    // exemplar attribute ram_0_6_9 MEM_LPC_FILE ram.lpc
    // exemplar attribute ram_0_6_9 MEM_INIT_FILE INIT_ALL_0s
    // exemplar attribute ram_0_7_8 MEM_LPC_FILE ram.lpc
    // exemplar attribute ram_0_7_8 MEM_INIT_FILE INIT_ALL_0s
    // exemplar attribute ram_1_0_7 MEM_LPC_FILE ram.lpc
    // exemplar attribute ram_1_0_7 MEM_INIT_FILE INIT_ALL_0s
    // exemplar attribute ram_1_1_6 MEM_LPC_FILE ram.lpc
    // exemplar attribute ram_1_1_6 MEM_INIT_FILE INIT_ALL_0s
    // exemplar attribute ram_1_2_5 MEM_LPC_FILE ram.lpc
    // exemplar attribute ram_1_2_5 MEM_INIT_FILE INIT_ALL_0s
    // exemplar attribute ram_1_3_4 MEM_LPC_FILE ram.lpc
    // exemplar attribute ram_1_3_4 MEM_INIT_FILE INIT_ALL_0s
    // exemplar attribute ram_1_4_3 MEM_LPC_FILE ram.lpc
    // exemplar attribute ram_1_4_3 MEM_INIT_FILE INIT_ALL_0s
    // exemplar attribute ram_1_5_2 MEM_LPC_FILE ram.lpc
    // exemplar attribute ram_1_5_2 MEM_INIT_FILE INIT_ALL_0s
    // exemplar attribute ram_1_6_1 MEM_LPC_FILE ram.lpc
    // exemplar attribute ram_1_6_1 MEM_INIT_FILE INIT_ALL_0s
    // exemplar attribute ram_1_7_0 MEM_LPC_FILE ram.lpc
    // exemplar attribute ram_1_7_0 MEM_INIT_FILE INIT_ALL_0s
    // exemplar attribute FF_1 GSR ENABLED
    // exemplar attribute FF_0 GSR ENABLED
    // exemplar end
endmodule