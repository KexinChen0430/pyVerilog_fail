module
cabac_binarization cabac_binarization_u0(
				//input
				.clk							(clk						),
				.rst_n							(rst_n						),
				.cabac_start_i					(start_d1_r					),
				.slice_type_i					(mb_type_i					),
				.mb_x_total_i					(mb_x_total_i				),
				.mb_y_total_i					(mb_y_total_i				),
				.mb_x_i							(mb_x_i						),
				.mb_y_i							(mb_y_i						),
			    .param_qp_i                     (param_qp_i                 ),
			    .sao_i                          (sao_i                      ),
				.luma_mode_i  			        (luma_mode_i  		        ),
				.chroma_mode_i                  (chroma_mode_i              ),
				.inter_cu_part_size_i			(mb_p_pu_mode_i				),
                .merge_flag_i                   (merge_flag_i               ),
                .merge_idx_i                    (merge_idx_i                ),
                .cu_skip_flag_i                 (cu_skip_flag_i             ),
            	.cu_split_flag_i				(mb_partition_i				),
				.luma_cbf_i						(cbf_y_w   				    ),
				.cr_cbf_i						(cbf_v_w				    ),
				.cb_cbf_i						(cbf_u_w				    ),
				.lcu_qp_i						(qp_i						),
				.coeff_data_i					(tq_rdata_i					),
				.cu_mvd_i						(mb_mvd_rdata_i				),
//                .mvd_idx_i                      (mvd_idx_i                  ),
				.table_build_end_i				(table_build_end_w			),
				.no_bit_flag_i					(no_bit_flag_w				),
				//output
				.slice_init_flag_o				(slice_init_flag_w			),
  				.cu_luma_mode_ren_o             (cu_luma_mode_ren_w         ),
                .cu_luma_mode_raddr_o           (cu_luma_mode_raddr_w       ),
                .cu_chroma_mode_ren_o           (cu_chroma_mode_ren_w       ),
                .cu_chroma_mode_raddr_o         (cu_chroma_mode_raddr_w     ),
				.cu_mvd_ren_o                   (cu_mvd_ren_w               ),
				.cu_mvd_raddr_o					(cu_mvd_raddr_w				),
				.cu_coeff_raddr_o				(cu_coeff_raddr_w			),
				.cu_coeff_ren_o					(cu_coeff_ren_w				),
				.cabac_mb_done_o				(cabac_mb_done_w			),
                .cabac_slice_done_o				(cabac_slice_done_w			),
				.coeff_type_o                   (coeff_type_w               ),
                .binary_pair_0_o				(ctx_pair_0_w				),
                .binary_pair_1_o				(ctx_pair_1_w				),
                .binary_pair_2_o				(ctx_pair_2_w				),
                .binary_pair_3_o				(ctx_pair_3_w				),
				.binary_pair_valid_num_o        (valid_num_bin_pair_w       ),
                .cabac_curr_state_o				(cabac_curr_state_w			)
);
//      slice initial
cabac_slice_init cabac_slice_init_u0(
				.clk							(clk					),
				.rst_n							(rst_n					),
				.start_slice_init_i				(slice_init_flag_w		),
				.slice_type_i					(mb_type_i				),
				.slice_qp_i						(slice_qp_r				),
				.table_build_end_o				(table_build_end_w		),
				.w_en_ctx_state_0_o				(w_en_ctx_state_0_w		),
    			.w_addr_ctx_state_0_o			(w_addr_ctx_state_0_w	),
    			.w_data_ctx_state_0_o			(w_data_ctx_state_0_w	),
    			.w_en_ctx_state_1_o				(w_en_ctx_state_1_w		),
    			.w_addr_ctx_state_1_o			(w_addr_ctx_state_1_w	),
    			.w_data_ctx_state_1_o			(w_data_ctx_state_1_w	),
    			.w_en_ctx_state_2_o				(w_en_ctx_state_2_w		),
    			.w_addr_ctx_state_2_o			(w_addr_ctx_state_2_w	),
    			.w_data_ctx_state_2_o			(w_data_ctx_state_2_w	),
    			.w_en_ctx_state_3_o				(w_en_ctx_state_3_w		),
    			.w_addr_ctx_state_3_o			(w_addr_ctx_state_3_w	),
    			.w_data_ctx_state_3_o			(w_data_ctx_state_3_w	),
    			.w_en_ctx_state_4_o				(w_en_ctx_state_4_w		),
    			.w_addr_ctx_state_4_o			(w_addr_ctx_state_4_w	),
    			.w_data_ctx_state_4_o			(w_data_ctx_state_4_w	)
);
//        modeling
cabac_modeling cabac_modeling_u0(
				//input
				.clk 							(clk						),
				.rst_n							(rst_n						),
                .modeling_pair_0_i				(ctx_pair_0_w				),
                .modeling_pair_1_i				(ctx_pair_1_w				),
                .modeling_pair_2_i				(ctx_pair_2_w				),
                .modeling_pair_3_i				(ctx_pair_3_w				),
                .valid_num_modeling_i			(valid_num_bin_pair_w       ),
                .cabac_start_i					(start_d1_r					),
                .slice_qp_i						(slice_qp_r					),
                .slice_type_i					(mb_type_i					),
                .first_mb_flag_i				(first_mb_flag_r			),
                .w_en_ctx_state_0_i				(w_en_ctx_state_0_w			),
    			.w_addr_ctx_state_0_i			(w_addr_ctx_state_0_w		),
    			.w_data_ctx_state_0_i			(w_data_ctx_state_0_w		),
    			.w_en_ctx_state_1_i				(w_en_ctx_state_1_w			),
    			.w_addr_ctx_state_1_i			(w_addr_ctx_state_1_w		),
    			.w_data_ctx_state_1_i			(w_data_ctx_state_1_w		),
    			.w_en_ctx_state_2_i				(w_en_ctx_state_2_w			),
    			.w_addr_ctx_state_2_i			(w_addr_ctx_state_2_w		),
    			.w_data_ctx_state_2_i			(w_data_ctx_state_2_w		),
    			.w_en_ctx_state_3_i				(w_en_ctx_state_3_w			),
    			.w_addr_ctx_state_3_i			(w_addr_ctx_state_3_w		),
    			.w_data_ctx_state_3_i			(w_data_ctx_state_3_w		),
    			.w_en_ctx_state_4_i				(w_en_ctx_state_4_w			),
    			.w_addr_ctx_state_4_i			(w_addr_ctx_state_4_w		),
    			.w_data_ctx_state_4_i			(w_data_ctx_state_4_w		),
                //output
                .modeling_ctx_pair_0_o			(modeling_ctx_pair_0_w		),
                .modeling_ctx_pair_1_o			(modeling_ctx_pair_1_w		),
                .modeling_ctx_pair_2_o			(modeling_ctx_pair_2_w		),
                .modeling_ctx_pair_3_o			(modeling_ctx_pair_3_w		),
                .valid_num_modeling_o			(valid_num_bae_w			)
);
//        bae
cabac_bae     cabac_bae_u0(
                .clk                            ( clk                       ),
                .rst_n                          ( rst_n                     ),
                .table_build_end_i 		        ( table_build_end_w         ),
                .bae_ctx_pair_0_i               ( modeling_ctx_pair_0_w     ),
                .bae_ctx_pair_1_i               ( modeling_ctx_pair_1_w     ),
                .bae_ctx_pair_2_i               ( modeling_ctx_pair_2_w     ),
                .bae_ctx_pair_3_i               ( modeling_ctx_pair_3_w     ),
                .bae_output_byte_o              ( output_byte_w			    ),
                .output_byte_en_o               ( output_byte_en_w		    ),
                .no_bit_flag_o			        ( no_bit_flag_w             )
);
endmodule