module ram2048x16 (Clock, ClockEn, Reset, WE, Address, Data, Q)/* synthesis NGD_DRC_MASK=1 */;
    input wire Clock;
    input wire ClockEn;
    input wire Reset;
    input wire WE;
    input wire [10:0] Address;
    input wire [15:0] Data;
    output wire [15:0] Q;
    wire scuba_vhi;
    wire scuba_vlo;
    defparam ram2048x16_0_0_3.INIT_DATA = "STATIC" ;
    defparam ram2048x16_0_0_3.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam ram2048x16_0_0_3.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_0_3.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_0_3.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_0_3.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_0_3.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_0_3.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_0_3.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_0_3.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_0_3.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_0_3.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_0_3.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_0_3.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_0_3.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_0_3.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_0_3.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_0_3.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_0_3.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_0_3.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_0_3.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_0_3.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_0_3.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_0_3.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_0_3.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_0_3.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_0_3.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_0_3.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_0_3.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_0_3.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_0_3.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_0_3.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_0_3.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_0_3.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_0_3.CSDECODE_B = "0b111" ;
    defparam ram2048x16_0_0_3.CSDECODE_A = "0b000" ;
    defparam ram2048x16_0_0_3.WRITEMODE_B = "NORMAL" ;
    defparam ram2048x16_0_0_3.WRITEMODE_A = "NORMAL" ;
    defparam ram2048x16_0_0_3.GSR = "ENABLED" ;
    defparam ram2048x16_0_0_3.RESETMODE = "ASYNC" ;
    defparam ram2048x16_0_0_3.REGMODE_B = "NOREG" ;
    defparam ram2048x16_0_0_3.REGMODE_A = "OUTREG" ;
    defparam ram2048x16_0_0_3.DATA_WIDTH_B = 4 ;
    defparam ram2048x16_0_0_3.DATA_WIDTH_A = 4 ;
    DP8KC ram2048x16_0_0_3 (.DIA8(scuba_vlo), .DIA7(scuba_vlo), .DIA6(scuba_vlo),
        .DIA5(scuba_vlo), .DIA4(scuba_vlo), .DIA3(Data[3]), .DIA2(Data[2]),
        .DIA1(Data[1]), .DIA0(Data[0]), .ADA12(Address[10]), .ADA11(Address[9]),
        .ADA10(Address[8]), .ADA9(Address[7]), .ADA8(Address[6]), .ADA7(Address[5]),
        .ADA6(Address[4]), .ADA5(Address[3]), .ADA4(Address[2]), .ADA3(Address[1]),
        .ADA2(Address[0]), .ADA1(scuba_vlo), .ADA0(scuba_vlo), .CEA(ClockEn),
        .OCEA(ClockEn), .CLKA(Clock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo),
        .CSA0(scuba_vlo), .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo),
        .DIB6(scuba_vlo), .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo),
        .DIB2(scuba_vlo), .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(scuba_vlo),
        .ADB11(scuba_vlo), .ADB10(scuba_vlo), .ADB9(scuba_vlo), .ADB8(scuba_vlo),
        .ADB7(scuba_vlo), .ADB6(scuba_vlo), .ADB5(scuba_vlo), .ADB4(scuba_vlo),
        .ADB3(scuba_vlo), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo),
        .CEB(scuba_vhi), .OCEB(scuba_vhi), .CLKB(scuba_vlo), .WEB(scuba_vlo),
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(scuba_vlo),
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(Q[3]), .DOA2(Q[2]),
        .DOA1(Q[1]), .DOA0(Q[0]), .DOB8(), .DOB7(), .DOB6(), .DOB5(), .DOB4(),
        .DOB3(), .DOB2(), .DOB1(), .DOB0())
             /* synthesis MEM_LPC_FILE="ram2048x16.lpc" */
             /* synthesis MEM_INIT_FILE="INIT_ALL_0s" */;
    defparam ram2048x16_0_1_2.INIT_DATA = "STATIC" ;
    defparam ram2048x16_0_1_2.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam ram2048x16_0_1_2.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_1_2.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_1_2.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_1_2.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_1_2.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_1_2.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_1_2.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_1_2.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_1_2.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_1_2.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_1_2.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_1_2.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_1_2.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_1_2.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_1_2.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_1_2.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_1_2.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_1_2.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_1_2.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_1_2.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_1_2.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_1_2.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_1_2.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_1_2.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_1_2.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_1_2.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_1_2.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_1_2.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_1_2.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_1_2.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_1_2.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_1_2.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_1_2.CSDECODE_B = "0b111" ;
    defparam ram2048x16_0_1_2.CSDECODE_A = "0b000" ;
    defparam ram2048x16_0_1_2.WRITEMODE_B = "NORMAL" ;
    defparam ram2048x16_0_1_2.WRITEMODE_A = "NORMAL" ;
    defparam ram2048x16_0_1_2.GSR = "ENABLED" ;
    defparam ram2048x16_0_1_2.RESETMODE = "ASYNC" ;
    defparam ram2048x16_0_1_2.REGMODE_B = "NOREG" ;
    defparam ram2048x16_0_1_2.REGMODE_A = "OUTREG" ;
    defparam ram2048x16_0_1_2.DATA_WIDTH_B = 4 ;
    defparam ram2048x16_0_1_2.DATA_WIDTH_A = 4 ;
    DP8KC ram2048x16_0_1_2 (.DIA8(scuba_vlo), .DIA7(scuba_vlo), .DIA6(scuba_vlo),
        .DIA5(scuba_vlo), .DIA4(scuba_vlo), .DIA3(Data[7]), .DIA2(Data[6]),
        .DIA1(Data[5]), .DIA0(Data[4]), .ADA12(Address[10]), .ADA11(Address[9]),
        .ADA10(Address[8]), .ADA9(Address[7]), .ADA8(Address[6]), .ADA7(Address[5]),
        .ADA6(Address[4]), .ADA5(Address[3]), .ADA4(Address[2]), .ADA3(Address[1]),
        .ADA2(Address[0]), .ADA1(scuba_vlo), .ADA0(scuba_vlo), .CEA(ClockEn),
        .OCEA(ClockEn), .CLKA(Clock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo),
        .CSA0(scuba_vlo), .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo),
        .DIB6(scuba_vlo), .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo),
        .DIB2(scuba_vlo), .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(scuba_vlo),
        .ADB11(scuba_vlo), .ADB10(scuba_vlo), .ADB9(scuba_vlo), .ADB8(scuba_vlo),
        .ADB7(scuba_vlo), .ADB6(scuba_vlo), .ADB5(scuba_vlo), .ADB4(scuba_vlo),
        .ADB3(scuba_vlo), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo),
        .CEB(scuba_vhi), .OCEB(scuba_vhi), .CLKB(scuba_vlo), .WEB(scuba_vlo),
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(scuba_vlo),
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(Q[7]), .DOA2(Q[6]),
        .DOA1(Q[5]), .DOA0(Q[4]), .DOB8(), .DOB7(), .DOB6(), .DOB5(), .DOB4(),
        .DOB3(), .DOB2(), .DOB1(), .DOB0())
             /* synthesis MEM_LPC_FILE="ram2048x16.lpc" */
             /* synthesis MEM_INIT_FILE="INIT_ALL_0s" */;
    defparam ram2048x16_0_2_1.INIT_DATA = "STATIC" ;
    defparam ram2048x16_0_2_1.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam ram2048x16_0_2_1.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_2_1.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_2_1.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_2_1.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_2_1.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_2_1.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_2_1.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_2_1.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_2_1.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_2_1.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_2_1.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_2_1.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_2_1.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_2_1.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_2_1.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_2_1.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_2_1.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_2_1.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_2_1.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_2_1.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_2_1.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_2_1.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_2_1.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_2_1.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_2_1.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_2_1.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_2_1.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_2_1.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_2_1.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_2_1.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_2_1.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_2_1.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_2_1.CSDECODE_B = "0b111" ;
    defparam ram2048x16_0_2_1.CSDECODE_A = "0b000" ;
    defparam ram2048x16_0_2_1.WRITEMODE_B = "NORMAL" ;
    defparam ram2048x16_0_2_1.WRITEMODE_A = "NORMAL" ;
    defparam ram2048x16_0_2_1.GSR = "ENABLED" ;
    defparam ram2048x16_0_2_1.RESETMODE = "ASYNC" ;
    defparam ram2048x16_0_2_1.REGMODE_B = "NOREG" ;
    defparam ram2048x16_0_2_1.REGMODE_A = "OUTREG" ;
    defparam ram2048x16_0_2_1.DATA_WIDTH_B = 4 ;
    defparam ram2048x16_0_2_1.DATA_WIDTH_A = 4 ;
    DP8KC ram2048x16_0_2_1 (.DIA8(scuba_vlo), .DIA7(scuba_vlo), .DIA6(scuba_vlo),
        .DIA5(scuba_vlo), .DIA4(scuba_vlo), .DIA3(Data[11]), .DIA2(Data[10]),
        .DIA1(Data[9]), .DIA0(Data[8]), .ADA12(Address[10]), .ADA11(Address[9]),
        .ADA10(Address[8]), .ADA9(Address[7]), .ADA8(Address[6]), .ADA7(Address[5]),
        .ADA6(Address[4]), .ADA5(Address[3]), .ADA4(Address[2]), .ADA3(Address[1]),
        .ADA2(Address[0]), .ADA1(scuba_vlo), .ADA0(scuba_vlo), .CEA(ClockEn),
        .OCEA(ClockEn), .CLKA(Clock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo),
        .CSA0(scuba_vlo), .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo),
        .DIB6(scuba_vlo), .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo),
        .DIB2(scuba_vlo), .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(scuba_vlo),
        .ADB11(scuba_vlo), .ADB10(scuba_vlo), .ADB9(scuba_vlo), .ADB8(scuba_vlo),
        .ADB7(scuba_vlo), .ADB6(scuba_vlo), .ADB5(scuba_vlo), .ADB4(scuba_vlo),
        .ADB3(scuba_vlo), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo),
        .CEB(scuba_vhi), .OCEB(scuba_vhi), .CLKB(scuba_vlo), .WEB(scuba_vlo),
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(scuba_vlo),
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(Q[11]), .DOA2(Q[10]),
        .DOA1(Q[9]), .DOA0(Q[8]), .DOB8(), .DOB7(), .DOB6(), .DOB5(), .DOB4(),
        .DOB3(), .DOB2(), .DOB1(), .DOB0())
             /* synthesis MEM_LPC_FILE="ram2048x16.lpc" */
             /* synthesis MEM_INIT_FILE="INIT_ALL_0s" */;
    VHI scuba_vhi_inst (.Z(scuba_vhi));
    VLO scuba_vlo_inst (.Z(scuba_vlo));
    defparam ram2048x16_0_3_0.INIT_DATA = "STATIC" ;
    defparam ram2048x16_0_3_0.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam ram2048x16_0_3_0.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_3_0.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_3_0.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_3_0.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_3_0.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_3_0.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_3_0.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_3_0.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_3_0.INITVAL_17 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_3_0.INITVAL_16 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_3_0.INITVAL_15 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_3_0.INITVAL_14 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_3_0.INITVAL_13 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_3_0.INITVAL_12 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_3_0.INITVAL_11 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_3_0.INITVAL_10 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_3_0.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_3_0.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_3_0.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_3_0.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_3_0.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_3_0.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_3_0.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_3_0.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_3_0.INITVAL_07 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_3_0.INITVAL_06 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_3_0.INITVAL_05 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_3_0.INITVAL_04 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_3_0.INITVAL_03 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_3_0.INITVAL_02 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_3_0.INITVAL_01 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_3_0.INITVAL_00 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam ram2048x16_0_3_0.CSDECODE_B = "0b111" ;
    defparam ram2048x16_0_3_0.CSDECODE_A = "0b000" ;
    defparam ram2048x16_0_3_0.WRITEMODE_B = "NORMAL" ;
    defparam ram2048x16_0_3_0.WRITEMODE_A = "NORMAL" ;
    defparam ram2048x16_0_3_0.GSR = "ENABLED" ;
    defparam ram2048x16_0_3_0.RESETMODE = "ASYNC" ;
    defparam ram2048x16_0_3_0.REGMODE_B = "NOREG" ;
    defparam ram2048x16_0_3_0.REGMODE_A = "OUTREG" ;
    defparam ram2048x16_0_3_0.DATA_WIDTH_B = 4 ;
    defparam ram2048x16_0_3_0.DATA_WIDTH_A = 4 ;
    DP8KC ram2048x16_0_3_0 (.DIA8(scuba_vlo), .DIA7(scuba_vlo), .DIA6(scuba_vlo),
        .DIA5(scuba_vlo), .DIA4(scuba_vlo), .DIA3(Data[15]), .DIA2(Data[14]),
        .DIA1(Data[13]), .DIA0(Data[12]), .ADA12(Address[10]), .ADA11(Address[9]),
        .ADA10(Address[8]), .ADA9(Address[7]), .ADA8(Address[6]), .ADA7(Address[5]),
        .ADA6(Address[4]), .ADA5(Address[3]), .ADA4(Address[2]), .ADA3(Address[1]),
        .ADA2(Address[0]), .ADA1(scuba_vlo), .ADA0(scuba_vlo), .CEA(ClockEn),
        .OCEA(ClockEn), .CLKA(Clock), .WEA(WE), .CSA2(scuba_vlo), .CSA1(scuba_vlo),
        .CSA0(scuba_vlo), .RSTA(Reset), .DIB8(scuba_vlo), .DIB7(scuba_vlo),
        .DIB6(scuba_vlo), .DIB5(scuba_vlo), .DIB4(scuba_vlo), .DIB3(scuba_vlo),
        .DIB2(scuba_vlo), .DIB1(scuba_vlo), .DIB0(scuba_vlo), .ADB12(scuba_vlo),
        .ADB11(scuba_vlo), .ADB10(scuba_vlo), .ADB9(scuba_vlo), .ADB8(scuba_vlo),
        .ADB7(scuba_vlo), .ADB6(scuba_vlo), .ADB5(scuba_vlo), .ADB4(scuba_vlo),
        .ADB3(scuba_vlo), .ADB2(scuba_vlo), .ADB1(scuba_vlo), .ADB0(scuba_vlo),
        .CEB(scuba_vhi), .OCEB(scuba_vhi), .CLKB(scuba_vlo), .WEB(scuba_vlo),
        .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo), .RSTB(scuba_vlo),
        .DOA8(), .DOA7(), .DOA6(), .DOA5(), .DOA4(), .DOA3(Q[15]), .DOA2(Q[14]),
        .DOA1(Q[13]), .DOA0(Q[12]), .DOB8(), .DOB7(), .DOB6(), .DOB5(),
        .DOB4(), .DOB3(), .DOB2(), .DOB1(), .DOB0())
             /* synthesis MEM_LPC_FILE="ram2048x16.lpc" */
             /* synthesis MEM_INIT_FILE="INIT_ALL_0s" */;
    // exemplar begin
    // exemplar attribute ram2048x16_0_0_3 MEM_LPC_FILE ram2048x16.lpc
    // exemplar attribute ram2048x16_0_0_3 MEM_INIT_FILE INIT_ALL_0s
    // exemplar attribute ram2048x16_0_1_2 MEM_LPC_FILE ram2048x16.lpc
    // exemplar attribute ram2048x16_0_1_2 MEM_INIT_FILE INIT_ALL_0s
    // exemplar attribute ram2048x16_0_2_1 MEM_LPC_FILE ram2048x16.lpc
    // exemplar attribute ram2048x16_0_2_1 MEM_INIT_FILE INIT_ALL_0s
    // exemplar attribute ram2048x16_0_3_0 MEM_LPC_FILE ram2048x16.lpc
    // exemplar attribute ram2048x16_0_3_0 MEM_INIT_FILE INIT_ALL_0s
    // exemplar end
endmodule