module multiplier64fp (
  clk, ce, rdy, a, b, result
)/* synthesis syn_black_box syn_noprune=1 */;
  input clk;
  input ce;
  output rdy;
  input [63 : 0] a;
  input [63 : 0] b;
  output [63 : 0] result;
  // synthesis translate_off
  wire \U0/op_inst/FLT_PT_OP/MULT.OP/OP/sign_op ;
  wire \NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/HND_SHK/RDY ;
  wire sig00000001;
  wire sig00000002;
  wire sig00000003;
  wire sig00000004;
  wire sig00000005;
  wire sig00000006;
  wire sig00000007;
  wire sig00000008;
  wire sig00000009;
  wire sig0000000a;
  wire sig0000000b;
  wire sig0000000c;
  wire sig0000000d;
  wire sig0000000e;
  wire sig0000000f;
  wire sig00000010;
  wire sig00000011;
  wire sig00000012;
  wire sig00000013;
  wire sig00000014;
  wire sig00000015;
  wire sig00000016;
  wire sig00000017;
  wire sig00000018;
  wire sig00000019;
  wire sig0000001a;
  wire sig0000001b;
  wire sig0000001c;
  wire sig0000001d;
  wire sig0000001e;
  wire sig0000001f;
  wire sig00000020;
  wire sig00000021;
  wire sig00000022;
  wire sig00000023;
  wire sig00000024;
  wire sig00000025;
  wire sig00000026;
  wire sig00000027;
  wire sig00000028;
  wire sig00000029;
  wire sig0000002a;
  wire sig0000002b;
  wire sig0000002c;
  wire sig0000002d;
  wire sig0000002e;
  wire sig0000002f;
  wire sig00000030;
  wire sig00000031;
  wire sig00000032;
  wire sig00000033;
  wire sig00000034;
  wire sig00000035;
  wire sig00000036;
  wire sig00000037;
  wire sig00000038;
  wire sig00000039;
  wire sig0000003a;
  wire sig0000003b;
  wire sig0000003c;
  wire sig0000003d;
  wire sig0000003e;
  wire sig0000003f;
  wire sig00000040;
  wire sig00000041;
  wire sig00000042;
  wire sig00000043;
  wire sig00000044;
  wire sig00000045;
  wire sig00000046;
  wire sig00000047;
  wire sig00000048;
  wire sig00000049;
  wire sig0000004a;
  wire sig0000004b;
  wire sig0000004c;
  wire sig0000004d;
  wire sig0000004e;
  wire sig0000004f;
  wire sig00000050;
  wire sig00000051;
  wire sig00000052;
  wire sig00000053;
  wire sig00000054;
  wire sig00000055;
  wire sig00000056;
  wire sig00000057;
  wire sig00000058;
  wire sig00000059;
  wire sig0000005a;
  wire sig0000005b;
  wire sig0000005c;
  wire sig0000005d;
  wire sig0000005e;
  wire sig0000005f;
  wire sig00000060;
  wire sig00000061;
  wire sig00000062;
  wire sig00000063;
  wire sig00000064;
  wire sig00000065;
  wire sig00000066;
  wire sig00000067;
  wire sig00000068;
  wire sig00000069;
  wire sig0000006a;
  wire sig0000006b;
  wire sig0000006c;
  wire sig0000006d;
  wire sig0000006e;
  wire sig0000006f;
  wire sig00000070;
  wire sig00000071;
  wire sig00000072;
  wire sig00000073;
  wire sig00000074;
  wire sig00000075;
  wire sig00000076;
  wire sig00000077;
  wire sig00000078;
  wire sig00000079;
  wire sig0000007a;
  wire sig0000007b;
  wire sig0000007c;
  wire sig0000007d;
  wire sig0000007e;
  wire sig0000007f;
  wire sig00000080;
  wire sig00000081;
  wire sig00000082;
  wire sig00000083;
  wire sig00000084;
  wire sig00000085;
  wire sig00000086;
  wire sig00000087;
  wire sig00000088;
  wire sig00000089;
  wire sig0000008a;
  wire sig0000008b;
  wire sig0000008c;
  wire sig0000008d;
  wire sig0000008e;
  wire sig0000008f;
  wire sig00000090;
  wire sig00000091;
  wire sig00000092;
  wire sig00000093;
  wire sig00000094;
  wire sig00000095;
  wire sig00000096;
  wire sig00000097;
  wire sig00000098;
  wire sig00000099;
  wire sig0000009a;
  wire sig0000009b;
  wire sig0000009c;
  wire sig0000009d;
  wire sig0000009e;
  wire sig0000009f;
  wire sig000000a0;
  wire sig000000a1;
  wire sig000000a2;
  wire sig000000a3;
  wire sig000000a4;
  wire sig000000a5;
  wire sig000000a6;
  wire sig000000a7;
  wire sig000000a8;
  wire sig000000a9;
  wire sig000000aa;
  wire sig000000ab;
  wire sig000000ac;
  wire sig000000ad;
  wire sig000000ae;
  wire sig000000af;
  wire sig000000b0;
  wire sig000000b1;
  wire sig000000b2;
  wire sig000000b3;
  wire sig000000b4;
  wire sig000000b5;
  wire sig000000b6;
  wire sig000000b7;
  wire sig000000b8;
  wire sig000000b9;
  wire sig000000ba;
  wire sig000000bb;
  wire sig000000bc;
  wire sig000000bd;
  wire sig000000be;
  wire sig000000bf;
  wire sig000000c0;
  wire sig000000c1;
  wire sig000000c2;
  wire sig000000c3;
  wire sig000000c4;
  wire sig000000c5;
  wire sig000000c6;
  wire sig000000c7;
  wire sig000000c8;
  wire sig000000c9;
  wire sig000000ca;
  wire sig000000cb;
  wire sig000000cc;
  wire sig000000cd;
  wire sig000000ce;
  wire sig000000cf;
  wire sig000000d0;
  wire sig000000d1;
  wire sig000000d2;
  wire sig000000d3;
  wire sig000000d4;
  wire sig000000d5;
  wire sig000000d6;
  wire sig000000d7;
  wire sig000000d8;
  wire sig000000d9;
  wire sig000000da;
  wire sig000000db;
  wire sig000000dc;
  wire sig000000dd;
  wire sig000000de;
  wire sig000000df;
  wire sig000000e0;
  wire sig000000e1;
  wire sig000000e2;
  wire sig000000e3;
  wire sig000000e4;
  wire sig000000e5;
  wire sig000000e6;
  wire sig000000e7;
  wire sig000000e8;
  wire sig000000e9;
  wire sig000000ea;
  wire sig000000eb;
  wire sig000000ec;
  wire sig000000ed;
  wire sig000000ee;
  wire sig000000ef;
  wire sig000000f0;
  wire sig000000f1;
  wire sig000000f2;
  wire sig000000f3;
  wire sig000000f4;
  wire sig000000f5;
  wire sig000000f6;
  wire sig000000f7;
  wire sig000000f8;
  wire sig000000f9;
  wire sig000000fa;
  wire sig000000fb;
  wire sig000000fc;
  wire sig000000fd;
  wire sig000000fe;
  wire sig000000ff;
  wire sig00000100;
  wire sig00000101;
  wire sig00000102;
  wire sig00000103;
  wire sig00000104;
  wire sig00000105;
  wire sig00000106;
  wire sig00000107;
  wire sig00000108;
  wire sig00000109;
  wire sig0000010a;
  wire sig0000010b;
  wire sig0000010c;
  wire sig0000010d;
  wire sig0000010e;
  wire sig0000010f;
  wire sig00000110;
  wire sig00000111;
  wire sig00000112;
  wire sig00000113;
  wire sig00000114;
  wire sig00000115;
  wire sig00000116;
  wire sig00000117;
  wire sig00000118;
  wire sig00000119;
  wire sig0000011a;
  wire sig0000011b;
  wire sig0000011c;
  wire sig0000011d;
  wire sig0000011e;
  wire sig0000011f;
  wire sig00000120;
  wire sig00000121;
  wire sig00000122;
  wire sig00000123;
  wire sig00000124;
  wire sig00000125;
  wire sig00000126;
  wire sig00000127;
  wire sig00000128;
  wire sig00000129;
  wire sig0000012a;
  wire sig0000012b;
  wire sig0000012c;
  wire sig0000012d;
  wire sig0000012e;
  wire sig0000012f;
  wire sig00000130;
  wire sig00000131;
  wire sig00000132;
  wire sig00000133;
  wire sig00000134;
  wire sig00000135;
  wire sig00000136;
  wire sig00000137;
  wire sig00000138;
  wire sig00000139;
  wire sig0000013a;
  wire sig0000013b;
  wire sig0000013c;
  wire sig0000013d;
  wire sig0000013e;
  wire sig0000013f;
  wire sig00000140;
  wire sig00000141;
  wire sig00000142;
  wire sig00000143;
  wire sig00000144;
  wire sig00000145;
  wire sig00000146;
  wire sig00000147;
  wire sig00000148;
  wire sig00000149;
  wire sig0000014a;
  wire sig0000014b;
  wire sig0000014c;
  wire sig0000014d;
  wire sig0000014e;
  wire sig0000014f;
  wire sig00000150;
  wire sig00000151;
  wire sig00000152;
  wire sig00000153;
  wire sig00000154;
  wire sig00000155;
  wire sig00000156;
  wire sig00000157;
  wire sig00000158;
  wire sig00000159;
  wire sig0000015a;
  wire sig0000015b;
  wire sig0000015c;
  wire sig0000015d;
  wire sig0000015e;
  wire sig0000015f;
  wire sig00000160;
  wire sig00000161;
  wire sig00000162;
  wire sig00000163;
  wire sig00000164;
  wire sig00000165;
  wire sig00000166;
  wire sig00000167;
  wire sig00000168;
  wire sig00000169;
  wire sig0000016a;
  wire sig0000016b;
  wire sig0000016c;
  wire sig0000016d;
  wire sig0000016e;
  wire sig0000016f;
  wire sig00000170;
  wire sig00000171;
  wire sig00000172;
  wire sig00000173;
  wire sig00000174;
  wire sig00000175;
  wire sig00000176;
  wire sig00000177;
  wire sig00000178;
  wire sig00000179;
  wire sig0000017a;
  wire sig0000017b;
  wire sig0000017c;
  wire sig0000017d;
  wire sig0000017e;
  wire sig0000017f;
  wire sig00000180;
  wire sig00000181;
  wire sig00000182;
  wire sig00000183;
  wire sig00000184;
  wire sig00000185;
  wire sig00000186;
  wire sig00000187;
  wire sig00000188;
  wire sig00000189;
  wire sig0000018a;
  wire sig0000018b;
  wire sig0000018c;
  wire sig0000018d;
  wire sig0000018e;
  wire sig0000018f;
  wire sig00000190;
  wire sig00000191;
  wire sig00000192;
  wire sig00000193;
  wire sig00000194;
  wire sig00000195;
  wire sig00000196;
  wire sig00000197;
  wire sig00000198;
  wire sig00000199;
  wire sig0000019a;
  wire sig0000019b;
  wire sig0000019c;
  wire sig0000019d;
  wire sig0000019e;
  wire sig0000019f;
  wire sig000001a0;
  wire sig000001a1;
  wire sig000001a2;
  wire sig000001a3;
  wire sig000001a4;
  wire sig000001a5;
  wire sig000001a6;
  wire sig000001a7;
  wire sig000001a8;
  wire sig000001a9;
  wire sig000001aa;
  wire sig000001ab;
  wire sig000001ac;
  wire sig000001ad;
  wire sig000001ae;
  wire sig000001af;
  wire sig000001b0;
  wire sig000001b1;
  wire sig000001b2;
  wire sig000001b3;
  wire sig000001b4;
  wire sig000001b5;
  wire sig000001b6;
  wire sig000001b7;
  wire sig000001b8;
  wire sig000001b9;
  wire sig000001ba;
  wire sig000001bb;
  wire sig000001bc;
  wire sig000001bd;
  wire sig000001be;
  wire sig000001bf;
  wire sig000001c0;
  wire sig000001c1;
  wire sig000001c2;
  wire sig000001c3;
  wire sig000001c4;
  wire sig000001c5;
  wire sig000001c6;
  wire sig000001c7;
  wire sig000001c8;
  wire sig000001c9;
  wire sig000001ca;
  wire sig000001cb;
  wire sig000001cc;
  wire sig000001cd;
  wire sig000001ce;
  wire sig000001cf;
  wire sig000001d0;
  wire sig000001d1;
  wire sig000001d2;
  wire sig000001d3;
  wire sig000001d4;
  wire sig000001d5;
  wire sig000001d6;
  wire sig000001d7;
  wire sig000001d8;
  wire sig000001d9;
  wire sig000001da;
  wire sig000001db;
  wire sig000001dc;
  wire sig000001dd;
  wire sig000001de;
  wire sig000001df;
  wire sig000001e0;
  wire sig000001e1;
  wire sig000001e2;
  wire sig000001e3;
  wire sig000001e4;
  wire sig000001e5;
  wire sig000001e6;
  wire sig000001e7;
  wire sig000001e8;
  wire sig000001e9;
  wire sig000001ea;
  wire sig000001eb;
  wire sig000001ec;
  wire sig000001ed;
  wire sig000001ee;
  wire sig000001ef;
  wire sig000001f0;
  wire sig000001f1;
  wire sig000001f2;
  wire sig000001f3;
  wire sig000001f4;
  wire sig000001f5;
  wire sig000001f6;
  wire sig000001f7;
  wire sig000001f8;
  wire sig000001f9;
  wire sig000001fa;
  wire sig000001fb;
  wire sig000001fc;
  wire sig000001fd;
  wire sig000001fe;
  wire sig000001ff;
  wire sig00000200;
  wire sig00000201;
  wire sig00000202;
  wire sig00000203;
  wire sig00000204;
  wire sig00000205;
  wire sig00000206;
  wire sig00000207;
  wire sig00000208;
  wire sig00000209;
  wire sig0000020a;
  wire sig0000020b;
  wire sig0000020c;
  wire sig0000020d;
  wire sig0000020e;
  wire sig0000020f;
  wire sig00000210;
  wire sig00000211;
  wire sig00000212;
  wire sig00000213;
  wire sig00000214;
  wire sig00000215;
  wire sig00000216;
  wire sig00000217;
  wire sig00000218;
  wire sig00000219;
  wire sig0000021a;
  wire sig0000021b;
  wire sig0000021c;
  wire sig0000021d;
  wire sig0000021e;
  wire sig0000021f;
  wire sig00000220;
  wire sig00000221;
  wire sig00000222;
  wire sig00000223;
  wire sig00000224;
  wire sig00000225;
  wire sig00000226;
  wire sig00000227;
  wire sig00000228;
  wire sig00000229;
  wire sig0000022a;
  wire sig0000022b;
  wire sig0000022c;
  wire sig0000022d;
  wire sig0000022e;
  wire sig0000022f;
  wire sig00000230;
  wire sig00000231;
  wire sig00000232;
  wire sig00000233;
  wire sig00000234;
  wire sig00000235;
  wire sig00000236;
  wire sig00000237;
  wire sig00000238;
  wire sig00000239;
  wire sig0000023a;
  wire sig0000023b;
  wire sig0000023c;
  wire sig0000023d;
  wire sig0000023e;
  wire sig0000023f;
  wire sig00000240;
  wire sig00000241;
  wire sig00000242;
  wire sig00000243;
  wire sig00000244;
  wire sig00000245;
  wire sig00000246;
  wire sig00000247;
  wire sig00000248;
  wire sig00000249;
  wire sig0000024a;
  wire sig0000024b;
  wire sig0000024c;
  wire sig0000024d;
  wire sig0000024e;
  wire sig0000024f;
  wire sig00000250;
  wire sig00000251;
  wire sig00000252;
  wire sig00000253;
  wire sig00000254;
  wire sig00000255;
  wire sig00000256;
  wire sig00000257;
  wire sig00000258;
  wire sig00000259;
  wire sig0000025a;
  wire sig0000025b;
  wire sig0000025c;
  wire sig0000025d;
  wire sig0000025e;
  wire sig0000025f;
  wire sig00000260;
  wire sig00000261;
  wire sig00000262;
  wire sig00000263;
  wire sig00000264;
  wire sig00000265;
  wire sig00000266;
  wire sig00000267;
  wire sig00000268;
  wire sig00000269;
  wire sig0000026a;
  wire sig0000026b;
  wire sig0000026c;
  wire sig0000026d;
  wire sig0000026e;
  wire sig0000026f;
  wire sig00000270;
  wire sig00000271;
  wire sig00000272;
  wire sig00000273;
  wire sig00000274;
  wire sig00000275;
  wire sig00000276;
  wire sig00000277;
  wire sig00000278;
  wire sig00000279;
  wire sig0000027a;
  wire sig0000027b;
  wire sig0000027c;
  wire sig0000027d;
  wire sig0000027e;
  wire sig0000027f;
  wire sig00000280;
  wire sig00000281;
  wire sig00000282;
  wire sig00000283;
  wire sig00000284;
  wire sig00000285;
  wire sig00000286;
  wire sig00000287;
  wire sig00000288;
  wire sig00000289;
  wire sig0000028a;
  wire sig0000028b;
  wire sig0000028c;
  wire sig0000028d;
  wire sig0000028e;
  wire sig0000028f;
  wire sig00000290;
  wire sig00000291;
  wire sig00000292;
  wire sig00000293;
  wire sig00000294;
  wire sig00000295;
  wire sig00000296;
  wire sig00000297;
  wire sig00000298;
  wire sig00000299;
  wire sig0000029a;
  wire sig0000029b;
  wire sig0000029c;
  wire sig0000029d;
  wire sig0000029e;
  wire sig0000029f;
  wire sig000002a0;
  wire sig000002a1;
  wire sig000002a2;
  wire sig000002a3;
  wire sig000002a4;
  wire sig000002a5;
  wire sig000002a6;
  wire sig000002a7;
  wire sig000002a8;
  wire sig000002a9;
  wire sig000002aa;
  wire sig000002ab;
  wire sig000002ac;
  wire sig000002ad;
  wire sig000002ae;
  wire sig000002af;
  wire sig000002b0;
  wire sig000002b1;
  wire sig000002b2;
  wire sig000002b3;
  wire sig000002b4;
  wire sig000002b5;
  wire sig000002b6;
  wire sig000002b7;
  wire sig000002b8;
  wire sig000002b9;
  wire sig000002ba;
  wire sig000002bb;
  wire sig000002bc;
  wire sig000002bd;
  wire sig000002be;
  wire sig000002bf;
  wire sig000002c0;
  wire sig000002c1;
  wire sig000002c2;
  wire sig000002c3;
  wire sig000002c4;
  wire sig000002c5;
  wire sig000002c6;
  wire sig000002c7;
  wire sig000002c8;
  wire sig000002c9;
  wire sig000002ca;
  wire sig000002cb;
  wire sig000002cc;
  wire sig000002cd;
  wire sig000002ce;
  wire sig000002cf;
  wire sig000002d0;
  wire sig000002d1;
  wire sig000002d2;
  wire sig000002d3;
  wire sig000002d4;
  wire sig000002d5;
  wire sig000002d6;
  wire sig000002d7;
  wire sig000002d8;
  wire sig000002d9;
  wire sig000002da;
  wire sig000002db;
  wire sig000002dc;
  wire sig000002dd;
  wire sig000002de;
  wire sig000002df;
  wire sig000002e0;
  wire sig000002e1;
  wire sig000002e2;
  wire sig000002e3;
  wire sig000002e4;
  wire sig000002e5;
  wire sig000002e6;
  wire sig000002e7;
  wire sig000002e8;
  wire sig000002e9;
  wire sig000002ea;
  wire sig000002eb;
  wire sig000002ec;
  wire sig000002ed;
  wire sig000002ee;
  wire sig000002ef;
  wire sig000002f0;
  wire sig000002f1;
  wire sig000002f2;
  wire sig000002f3;
  wire sig000002f4;
  wire sig000002f5;
  wire sig000002f6;
  wire sig000002f7;
  wire sig000002f8;
  wire sig000002f9;
  wire sig000002fa;
  wire sig000002fb;
  wire sig000002fc;
  wire sig000002fd;
  wire sig000002fe;
  wire sig000002ff;
  wire sig00000300;
  wire sig00000301;
  wire sig00000302;
  wire sig00000303;
  wire sig00000304;
  wire sig00000305;
  wire sig00000306;
  wire sig00000307;
  wire sig00000308;
  wire sig00000309;
  wire sig0000030a;
  wire sig0000030b;
  wire sig0000030c;
  wire sig0000030d;
  wire sig0000030e;
  wire sig0000030f;
  wire sig00000310;
  wire sig00000311;
  wire sig00000312;
  wire sig00000313;
  wire sig00000314;
  wire sig00000315;
  wire sig00000316;
  wire sig00000317;
  wire sig00000318;
  wire sig00000319;
  wire sig0000031a;
  wire sig0000031b;
  wire sig0000031c;
  wire sig0000031d;
  wire sig0000031e;
  wire sig0000031f;
  wire sig00000320;
  wire sig00000321;
  wire sig00000322;
  wire sig00000323;
  wire sig00000324;
  wire sig00000325;
  wire sig00000326;
  wire sig00000327;
  wire sig00000328;
  wire sig00000329;
  wire sig0000032a;
  wire sig0000032b;
  wire sig0000032c;
  wire sig0000032d;
  wire sig0000032e;
  wire sig0000032f;
  wire sig00000330;
  wire sig00000331;
  wire sig00000332;
  wire sig00000333;
  wire sig00000334;
  wire sig00000335;
  wire sig00000336;
  wire sig00000337;
  wire sig00000338;
  wire sig00000339;
  wire sig0000033a;
  wire sig0000033b;
  wire sig0000033c;
  wire sig0000033d;
  wire sig0000033e;
  wire sig0000033f;
  wire sig00000340;
  wire sig00000341;
  wire sig00000342;
  wire sig00000343;
  wire sig00000344;
  wire sig00000345;
  wire sig00000346;
  wire sig00000347;
  wire sig00000348;
  wire sig00000349;
  wire sig0000034a;
  wire sig0000034b;
  wire sig0000034c;
  wire sig0000034d;
  wire sig0000034e;
  wire sig0000034f;
  wire sig00000350;
  wire sig00000351;
  wire sig00000352;
  wire sig00000353;
  wire sig00000354;
  wire sig00000355;
  wire sig00000356;
  wire sig00000357;
  wire sig00000358;
  wire sig00000359;
  wire sig0000035a;
  wire sig0000035b;
  wire sig0000035c;
  wire sig0000035d;
  wire sig0000035e;
  wire sig0000035f;
  wire sig00000360;
  wire sig00000361;
  wire sig00000362;
  wire sig00000363;
  wire sig00000364;
  wire sig00000365;
  wire sig00000366;
  wire sig00000367;
  wire sig00000368;
  wire sig00000369;
  wire sig0000036a;
  wire sig0000036b;
  wire sig0000036c;
  wire sig0000036d;
  wire sig0000036e;
  wire sig0000036f;
  wire sig00000370;
  wire sig00000371;
  wire sig00000372;
  wire sig00000373;
  wire sig00000374;
  wire sig00000375;
  wire sig00000376;
  wire sig00000377;
  wire sig00000378;
  wire sig00000379;
  wire sig0000037a;
  wire sig0000037b;
  wire sig0000037c;
  wire sig0000037d;
  wire sig0000037e;
  wire sig0000037f;
  wire sig00000380;
  wire sig00000381;
  wire sig00000382;
  wire sig00000383;
  wire sig00000384;
  wire sig00000385;
  wire sig00000386;
  wire sig00000387;
  wire sig00000388;
  wire sig00000389;
  wire sig0000038a;
  wire sig0000038b;
  wire sig0000038c;
  wire sig0000038d;
  wire sig0000038e;
  wire sig0000038f;
  wire sig00000390;
  wire sig00000391;
  wire sig00000392;
  wire sig00000393;
  wire sig00000394;
  wire sig00000395;
  wire sig00000396;
  wire sig00000397;
  wire sig00000398;
  wire sig00000399;
  wire sig0000039a;
  wire sig0000039b;
  wire sig0000039c;
  wire sig0000039d;
  wire sig0000039e;
  wire sig0000039f;
  wire sig000003a0;
  wire sig000003a1;
  wire sig000003a2;
  wire sig000003a3;
  wire sig000003a4;
  wire sig000003a5;
  wire sig000003a6;
  wire sig000003a7;
  wire sig000003a8;
  wire sig000003a9;
  wire sig000003aa;
  wire sig000003ab;
  wire sig000003ac;
  wire sig000003ad;
  wire sig000003ae;
  wire sig000003af;
  wire sig000003b0;
  wire sig000003b1;
  wire sig000003b2;
  wire sig000003b3;
  wire sig000003b4;
  wire sig000003b5;
  wire sig000003b6;
  wire sig000003b7;
  wire sig000003b8;
  wire sig000003b9;
  wire sig000003ba;
  wire sig000003bb;
  wire sig000003bc;
  wire sig000003bd;
  wire sig000003be;
  wire sig000003bf;
  wire sig000003c0;
  wire sig000003c1;
  wire sig000003c2;
  wire sig000003c3;
  wire sig000003c4;
  wire sig000003c5;
  wire sig000003c6;
  wire sig000003c7;
  wire sig000003c8;
  wire sig000003c9;
  wire sig000003ca;
  wire sig000003cb;
  wire sig000003cc;
  wire sig000003cd;
  wire sig000003ce;
  wire sig000003cf;
  wire sig000003d0;
  wire sig000003d1;
  wire sig000003d2;
  wire sig000003d3;
  wire sig000003d4;
  wire sig000003d5;
  wire sig000003d6;
  wire sig000003d7;
  wire sig000003d8;
  wire sig000003d9;
  wire sig000003da;
  wire sig000003db;
  wire sig000003dc;
  wire sig000003dd;
  wire sig000003de;
  wire sig000003df;
  wire sig000003e0;
  wire sig000003e1;
  wire sig000003e2;
  wire sig000003e3;
  wire sig000003e4;
  wire sig000003e5;
  wire sig000003e6;
  wire sig000003e7;
  wire sig000003e8;
  wire sig000003e9;
  wire sig000003ea;
  wire sig000003eb;
  wire sig000003ec;
  wire sig000003ed;
  wire sig000003ee;
  wire sig000003ef;
  wire sig000003f0;
  wire sig000003f1;
  wire sig000003f2;
  wire sig000003f3;
  wire sig000003f4;
  wire sig000003f5;
  wire sig000003f6;
  wire sig000003f7;
  wire sig000003f8;
  wire sig000003f9;
  wire sig000003fa;
  wire sig000003fb;
  wire sig000003fc;
  wire sig000003fd;
  wire sig000003fe;
  wire sig000003ff;
  wire sig00000400;
  wire sig00000401;
  wire sig00000402;
  wire sig00000403;
  wire sig00000404;
  wire sig00000405;
  wire sig00000406;
  wire sig00000407;
  wire sig00000408;
  wire sig00000409;
  wire sig0000040a;
  wire sig0000040b;
  wire sig0000040c;
  wire sig0000040d;
  wire sig0000040e;
  wire sig0000040f;
  wire sig00000410;
  wire sig00000411;
  wire sig00000412;
  wire sig00000413;
  wire sig00000414;
  wire sig00000415;
  wire sig00000416;
  wire sig00000417;
  wire sig00000418;
  wire sig00000419;
  wire sig0000041a;
  wire sig0000041b;
  wire sig0000041c;
  wire sig0000041d;
  wire sig0000041e;
  wire sig0000041f;
  wire sig00000420;
  wire sig00000421;
  wire sig00000422;
  wire sig00000423;
  wire sig00000424;
  wire sig00000425;
  wire sig00000426;
  wire sig00000427;
  wire sig00000428;
  wire sig00000429;
  wire sig0000042a;
  wire sig0000042b;
  wire sig0000042c;
  wire sig0000042d;
  wire sig0000042e;
  wire sig0000042f;
  wire sig00000430;
  wire sig00000431;
  wire sig00000432;
  wire sig00000433;
  wire sig00000434;
  wire sig00000435;
  wire sig00000436;
  wire sig00000437;
  wire sig00000438;
  wire sig00000439;
  wire sig0000043a;
  wire sig0000043b;
  wire sig0000043c;
  wire sig0000043d;
  wire sig0000043e;
  wire sig0000043f;
  wire sig00000440;
  wire sig00000441;
  wire sig00000442;
  wire sig00000443;
  wire sig00000444;
  wire sig00000445;
  wire sig00000446;
  wire sig00000447;
  wire sig00000448;
  wire sig00000449;
  wire sig0000044a;
  wire sig0000044b;
  wire sig0000044c;
  wire sig0000044d;
  wire sig0000044e;
  wire sig0000044f;
  wire sig00000450;
  wire sig00000451;
  wire sig00000452;
  wire sig00000453;
  wire sig00000454;
  wire sig00000455;
  wire sig00000456;
  wire sig00000457;
  wire sig00000458;
  wire sig00000459;
  wire sig0000045a;
  wire sig0000045b;
  wire sig0000045c;
  wire sig0000045d;
  wire sig0000045e;
  wire sig0000045f;
  wire sig00000460;
  wire sig00000461;
  wire sig00000462;
  wire sig00000463;
  wire sig00000464;
  wire sig00000465;
  wire sig00000466;
  wire sig00000467;
  wire sig00000468;
  wire sig00000469;
  wire sig0000046a;
  wire sig0000046b;
  wire sig0000046c;
  wire sig0000046d;
  wire sig0000046e;
  wire sig0000046f;
  wire sig00000470;
  wire sig00000471;
  wire sig00000472;
  wire sig00000473;
  wire sig00000474;
  wire sig00000475;
  wire sig00000476;
  wire sig00000477;
  wire sig00000478;
  wire sig00000479;
  wire sig0000047a;
  wire sig0000047b;
  wire sig0000047c;
  wire sig0000047d;
  wire sig0000047e;
  wire sig0000047f;
  wire sig00000480;
  wire sig00000481;
  wire sig00000482;
  wire sig00000483;
  wire sig00000484;
  wire sig00000485;
  wire sig00000486;
  wire sig00000487;
  wire sig00000488;
  wire sig00000489;
  wire sig0000048a;
  wire sig0000048b;
  wire sig0000048c;
  wire sig0000048d;
  wire sig0000048e;
  wire sig0000048f;
  wire sig00000490;
  wire sig00000491;
  wire sig00000492;
  wire sig00000493;
  wire sig00000494;
  wire sig00000495;
  wire sig00000496;
  wire sig00000497;
  wire sig00000498;
  wire sig00000499;
  wire sig0000049a;
  wire sig0000049b;
  wire sig0000049c;
  wire sig0000049d;
  wire sig0000049e;
  wire sig0000049f;
  wire sig000004a0;
  wire sig000004a1;
  wire sig000004a2;
  wire sig000004a3;
  wire sig000004a4;
  wire sig000004a5;
  wire sig000004a6;
  wire sig000004a7;
  wire sig000004a8;
  wire sig000004a9;
  wire sig000004aa;
  wire sig000004ab;
  wire sig000004ac;
  wire sig000004ad;
  wire sig000004ae;
  wire sig000004af;
  wire sig000004b0;
  wire sig000004b1;
  wire sig000004b2;
  wire sig000004b3;
  wire sig000004b4;
  wire sig000004b5;
  wire sig000004b6;
  wire sig000004b7;
  wire sig000004b8;
  wire sig000004b9;
  wire sig000004ba;
  wire sig000004bb;
  wire sig000004bc;
  wire sig000004bd;
  wire sig000004be;
  wire sig000004bf;
  wire sig000004c0;
  wire sig000004c1;
  wire sig000004c2;
  wire sig000004c3;
  wire sig000004c4;
  wire sig000004c5;
  wire sig000004c6;
  wire sig000004c7;
  wire sig000004c8;
  wire sig000004c9;
  wire sig000004ca;
  wire sig000004cb;
  wire sig000004cc;
  wire sig000004cd;
  wire sig000004ce;
  wire sig000004cf;
  wire sig000004d0;
  wire sig000004d1;
  wire sig000004d2;
  wire sig000004d3;
  wire sig000004d4;
  wire sig000004d5;
  wire sig000004d6;
  wire sig000004d7;
  wire sig000004d8;
  wire sig000004d9;
  wire sig000004da;
  wire sig000004db;
  wire sig000004dc;
  wire sig000004dd;
  wire sig000004de;
  wire sig000004df;
  wire sig000004e0;
  wire sig000004e1;
  wire sig000004e2;
  wire sig000004e3;
  wire sig000004e4;
  wire sig000004e5;
  wire sig000004e6;
  wire sig000004e7;
  wire sig000004e8;
  wire sig000004e9;
  wire sig000004ea;
  wire sig000004eb;
  wire sig000004ec;
  wire sig000004ed;
  wire sig000004ee;
  wire sig000004ef;
  wire sig000004f0;
  wire sig000004f1;
  wire sig000004f2;
  wire sig000004f3;
  wire sig000004f4;
  wire sig000004f5;
  wire sig000004f6;
  wire sig000004f7;
  wire sig000004f8;
  wire sig000004f9;
  wire sig000004fa;
  wire sig000004fb;
  wire sig000004fc;
  wire sig000004fd;
  wire sig000004fe;
  wire sig000004ff;
  wire sig00000500;
  wire sig00000501;
  wire sig00000502;
  wire sig00000503;
  wire sig00000504;
  wire sig00000505;
  wire sig00000506;
  wire sig00000507;
  wire sig00000508;
  wire sig00000509;
  wire sig0000050a;
  wire sig0000050b;
  wire sig0000050c;
  wire sig0000050d;
  wire sig0000050e;
  wire sig0000050f;
  wire sig00000510;
  wire sig00000511;
  wire sig00000512;
  wire sig00000513;
  wire sig00000514;
  wire sig00000515;
  wire sig00000516;
  wire sig00000517;
  wire sig00000518;
  wire sig00000519;
  wire sig0000051a;
  wire sig0000051b;
  wire sig0000051c;
  wire sig0000051d;
  wire sig0000051e;
  wire sig0000051f;
  wire sig00000520;
  wire sig00000521;
  wire sig00000522;
  wire sig00000523;
  wire sig00000524;
  wire sig00000525;
  wire sig00000526;
  wire sig00000527;
  wire sig00000528;
  wire sig00000529;
  wire sig0000052a;
  wire sig0000052b;
  wire sig0000052c;
  wire sig0000052d;
  wire sig0000052e;
  wire sig0000052f;
  wire sig00000530;
  wire sig00000531;
  wire sig00000532;
  wire sig00000533;
  wire sig00000534;
  wire sig00000535;
  wire sig00000536;
  wire sig00000537;
  wire sig00000538;
  wire sig00000539;
  wire sig0000053a;
  wire sig0000053b;
  wire sig0000053c;
  wire sig0000053d;
  wire sig0000053e;
  wire sig0000053f;
  wire sig00000540;
  wire sig00000541;
  wire sig00000542;
  wire sig00000543;
  wire sig00000544;
  wire sig00000545;
  wire sig00000546;
  wire sig00000547;
  wire sig00000548;
  wire sig00000549;
  wire sig0000054a;
  wire sig0000054b;
  wire sig0000054c;
  wire sig0000054d;
  wire sig0000054e;
  wire sig0000054f;
  wire sig00000550;
  wire sig00000551;
  wire sig00000552;
  wire sig00000553;
  wire sig00000554;
  wire sig00000555;
  wire sig00000556;
  wire sig00000557;
  wire sig00000558;
  wire sig00000559;
  wire sig0000055a;
  wire sig0000055b;
  wire sig0000055c;
  wire sig0000055d;
  wire sig0000055e;
  wire sig0000055f;
  wire sig00000560;
  wire sig00000561;
  wire sig00000562;
  wire sig00000563;
  wire sig00000564;
  wire sig00000565;
  wire sig00000566;
  wire sig00000567;
  wire sig00000568;
  wire sig00000569;
  wire sig0000056a;
  wire sig0000056b;
  wire sig0000056c;
  wire sig0000056d;
  wire sig0000056e;
  wire sig0000056f;
  wire sig00000570;
  wire sig00000571;
  wire sig00000572;
  wire sig00000573;
  wire sig00000574;
  wire sig00000575;
  wire sig00000576;
  wire sig00000577;
  wire sig00000578;
  wire sig00000579;
  wire sig0000057a;
  wire sig0000057b;
  wire sig0000057c;
  wire sig0000057d;
  wire sig0000057e;
  wire sig0000057f;
  wire sig00000580;
  wire sig00000581;
  wire sig00000582;
  wire sig00000583;
  wire sig00000584;
  wire sig00000585;
  wire sig00000586;
  wire sig00000587;
  wire sig00000588;
  wire sig00000589;
  wire sig0000058a;
  wire sig0000058b;
  wire sig0000058c;
  wire sig0000058d;
  wire sig0000058e;
  wire sig0000058f;
  wire sig00000590;
  wire sig00000591;
  wire sig00000592;
  wire sig00000593;
  wire sig00000594;
  wire sig00000595;
  wire sig00000596;
  wire sig00000597;
  wire sig00000598;
  wire sig00000599;
  wire sig0000059a;
  wire sig0000059b;
  wire sig0000059c;
  wire sig0000059d;
  wire sig0000059e;
  wire sig0000059f;
  wire sig000005a0;
  wire sig000005a1;
  wire sig000005a2;
  wire sig000005a3;
  wire sig000005a4;
  wire sig000005a5;
  wire sig000005a6;
  wire sig000005a7;
  wire sig000005a8;
  wire sig000005a9;
  wire sig000005aa;
  wire sig000005ab;
  wire sig000005ac;
  wire sig000005ad;
  wire sig000005ae;
  wire sig000005af;
  wire sig000005b0;
  wire sig000005b1;
  wire sig000005b2;
  wire sig000005b3;
  wire sig000005b4;
  wire sig000005b5;
  wire sig000005b6;
  wire sig000005b7;
  wire sig000005b8;
  wire sig000005b9;
  wire sig000005ba;
  wire sig000005bb;
  wire sig000005bc;
  wire sig000005bd;
  wire sig000005be;
  wire sig000005bf;
  wire sig000005c0;
  wire sig000005c1;
  wire sig000005c2;
  wire sig000005c3;
  wire sig000005c4;
  wire sig000005c5;
  wire sig000005c6;
  wire sig000005c7;
  wire sig000005c8;
  wire sig000005c9;
  wire sig000005ca;
  wire sig000005cb;
  wire sig000005cc;
  wire sig000005cd;
  wire sig000005ce;
  wire sig000005cf;
  wire sig000005d0;
  wire sig000005d1;
  wire sig000005d2;
  wire sig000005d3;
  wire sig000005d4;
  wire sig000005d5;
  wire sig000005d6;
  wire sig000005d7;
  wire sig000005d8;
  wire sig000005d9;
  wire sig000005da;
  wire sig000005db;
  wire sig000005dc;
  wire sig000005dd;
  wire sig000005de;
  wire sig000005df;
  wire sig000005e0;
  wire sig000005e1;
  wire sig000005e2;
  wire sig000005e3;
  wire sig000005e4;
  wire sig000005e5;
  wire sig000005e6;
  wire sig000005e7;
  wire sig000005e8;
  wire sig000005e9;
  wire sig000005ea;
  wire sig000005eb;
  wire sig000005ec;
  wire sig000005ed;
  wire sig000005ee;
  wire sig000005ef;
  wire sig000005f0;
  wire sig000005f1;
  wire sig000005f2;
  wire sig000005f3;
  wire sig000005f4;
  wire sig000005f5;
  wire sig000005f6;
  wire sig000005f7;
  wire sig000005f8;
  wire sig000005f9;
  wire sig000005fa;
  wire sig000005fb;
  wire sig000005fc;
  wire sig000005fd;
  wire sig000005fe;
  wire sig000005ff;
  wire sig00000600;
  wire sig00000601;
  wire sig00000602;
  wire sig00000603;
  wire sig00000604;
  wire sig00000605;
  wire sig00000606;
  wire sig00000607;
  wire sig00000608;
  wire sig00000609;
  wire sig0000060a;
  wire sig0000060b;
  wire sig0000060c;
  wire sig0000060d;
  wire sig0000060e;
  wire sig0000060f;
  wire sig00000610;
  wire sig00000611;
  wire sig00000612;
  wire sig00000613;
  wire sig00000614;
  wire sig00000615;
  wire sig00000616;
  wire sig00000617;
  wire sig00000618;
  wire sig00000619;
  wire sig0000061a;
  wire sig0000061b;
  wire sig0000061c;
  wire sig0000061d;
  wire sig0000061e;
  wire sig0000061f;
  wire sig00000620;
  wire sig00000621;
  wire sig00000622;
  wire sig00000623;
  wire sig00000624;
  wire sig00000625;
  wire sig00000626;
  wire sig00000627;
  wire sig00000628;
  wire sig00000629;
  wire sig0000062a;
  wire sig0000062b;
  wire sig0000062c;
  wire sig0000062d;
  wire sig0000062e;
  wire sig0000062f;
  wire sig00000630;
  wire sig00000631;
  wire sig00000632;
  wire NLW_blk0000010f_O_UNCONNECTED;
  wire NLW_blk00000273_Q15_UNCONNECTED;
  wire NLW_blk00000275_Q15_UNCONNECTED;
  wire NLW_blk00000277_Q15_UNCONNECTED;
  wire NLW_blk00000279_Q15_UNCONNECTED;
  wire NLW_blk0000027b_Q15_UNCONNECTED;
  wire NLW_blk0000027d_Q15_UNCONNECTED;
  wire NLW_blk0000027f_Q15_UNCONNECTED;
  wire NLW_blk00000281_Q15_UNCONNECTED;
  wire NLW_blk00000283_Q15_UNCONNECTED;
  wire NLW_blk00000285_Q15_UNCONNECTED;
  wire NLW_blk00000287_Q15_UNCONNECTED;
  wire NLW_blk00000289_Q15_UNCONNECTED;
  wire NLW_blk0000028b_Q15_UNCONNECTED;
  wire NLW_blk0000028d_Q15_UNCONNECTED;
  wire NLW_blk0000028f_Q15_UNCONNECTED;
  wire NLW_blk00000291_Q15_UNCONNECTED;
  wire NLW_blk00000293_Q15_UNCONNECTED;
  wire NLW_blk00000295_Q15_UNCONNECTED;
  wire NLW_blk00000297_Q15_UNCONNECTED;
  wire NLW_blk00000299_Q15_UNCONNECTED;
  wire NLW_blk0000029b_Q15_UNCONNECTED;
  wire NLW_blk0000029d_Q15_UNCONNECTED;
  wire NLW_blk0000029f_Q15_UNCONNECTED;
  wire NLW_blk000002a1_Q15_UNCONNECTED;
  wire NLW_blk000002a3_Q15_UNCONNECTED;
  wire NLW_blk000002a5_Q15_UNCONNECTED;
  wire NLW_blk000002a7_Q15_UNCONNECTED;
  wire NLW_blk000002a9_Q15_UNCONNECTED;
  wire NLW_blk000002ab_Q15_UNCONNECTED;
  wire NLW_blk000002ad_Q15_UNCONNECTED;
  wire NLW_blk000002af_Q15_UNCONNECTED;
  wire NLW_blk000002b1_Q15_UNCONNECTED;
  wire NLW_blk000002b3_Q15_UNCONNECTED;
  wire NLW_blk000002b5_Q15_UNCONNECTED;
  wire NLW_blk000002b7_Q15_UNCONNECTED;
  wire NLW_blk000002b9_Q15_UNCONNECTED;
  wire NLW_blk000002bb_Q15_UNCONNECTED;
  wire NLW_blk000002bd_Q15_UNCONNECTED;
  wire NLW_blk000002bf_Q15_UNCONNECTED;
  wire NLW_blk000002c1_Q15_UNCONNECTED;
  wire NLW_blk000002c3_Q15_UNCONNECTED;
  wire NLW_blk000002c5_Q15_UNCONNECTED;
  wire NLW_blk000002c7_Q15_UNCONNECTED;
  wire NLW_blk000002c9_Q15_UNCONNECTED;
  wire NLW_blk000002cb_Q15_UNCONNECTED;
  wire NLW_blk000002cd_Q15_UNCONNECTED;
  wire NLW_blk000002cf_Q15_UNCONNECTED;
  wire NLW_blk000002d1_Q15_UNCONNECTED;
  wire NLW_blk000002d3_Q15_UNCONNECTED;
  wire NLW_blk000002d5_Q15_UNCONNECTED;
  wire NLW_blk000002d7_Q15_UNCONNECTED;
  wire NLW_blk000002d9_Q15_UNCONNECTED;
  wire NLW_blk000002db_Q15_UNCONNECTED;
  wire NLW_blk000002dd_Q15_UNCONNECTED;
  wire NLW_blk000002df_Q15_UNCONNECTED;
  wire NLW_blk000002e1_Q15_UNCONNECTED;
  wire NLW_blk000002e3_Q15_UNCONNECTED;
  wire NLW_blk000002e5_Q15_UNCONNECTED;
  wire NLW_blk000002e7_Q15_UNCONNECTED;
  wire NLW_blk000002e9_Q15_UNCONNECTED;
  wire NLW_blk000002eb_Q15_UNCONNECTED;
  wire NLW_blk000002ed_Q15_UNCONNECTED;
  wire NLW_blk000002ef_Q15_UNCONNECTED;
  wire NLW_blk000002f1_Q15_UNCONNECTED;
  wire NLW_blk000002f3_Q15_UNCONNECTED;
  wire NLW_blk000002f5_Q15_UNCONNECTED;
  wire NLW_blk000002f7_Q15_UNCONNECTED;
  wire NLW_blk000002f9_Q15_UNCONNECTED;
  wire NLW_blk000002fb_Q15_UNCONNECTED;
  wire NLW_blk000002fd_Q15_UNCONNECTED;
  wire NLW_blk000002ff_Q15_UNCONNECTED;
  wire NLW_blk00000301_Q15_UNCONNECTED;
  wire NLW_blk00000303_Q15_UNCONNECTED;
  wire NLW_blk00000305_Q15_UNCONNECTED;
  wire NLW_blk00000307_Q15_UNCONNECTED;
  wire NLW_blk00000309_Q15_UNCONNECTED;
  wire NLW_blk0000030b_Q15_UNCONNECTED;
  wire NLW_blk0000030d_Q15_UNCONNECTED;
  wire NLW_blk0000030f_Q15_UNCONNECTED;
  wire NLW_blk00000311_Q15_UNCONNECTED;
  wire NLW_blk00000313_Q15_UNCONNECTED;
  wire NLW_blk00000315_Q15_UNCONNECTED;
  wire NLW_blk00000317_Q15_UNCONNECTED;
  wire NLW_blk00000319_Q15_UNCONNECTED;
  wire NLW_blk0000031b_Q15_UNCONNECTED;
  wire NLW_blk0000031d_Q15_UNCONNECTED;
  wire NLW_blk0000031f_Q15_UNCONNECTED;
  wire NLW_blk00000321_Q15_UNCONNECTED;
  wire NLW_blk00000323_Q15_UNCONNECTED;
  wire NLW_blk00000325_Q15_UNCONNECTED;
  wire NLW_blk00000327_Q15_UNCONNECTED;
  wire NLW_blk00000329_Q15_UNCONNECTED;
  wire NLW_blk0000032b_Q15_UNCONNECTED;
  wire NLW_blk0000032d_Q15_UNCONNECTED;
  wire NLW_blk0000032f_Q15_UNCONNECTED;
  wire NLW_blk00000331_Q15_UNCONNECTED;
  wire NLW_blk00000333_Q15_UNCONNECTED;
  wire NLW_blk00000335_Q15_UNCONNECTED;
  wire NLW_blk00000337_Q15_UNCONNECTED;
  wire NLW_blk00000339_Q15_UNCONNECTED;
  wire NLW_blk0000033b_Q15_UNCONNECTED;
  wire NLW_blk0000033d_Q15_UNCONNECTED;
  wire NLW_blk0000033f_Q15_UNCONNECTED;
  wire NLW_blk00000341_Q15_UNCONNECTED;
  wire NLW_blk00000343_Q15_UNCONNECTED;
  wire NLW_blk00000345_Q15_UNCONNECTED;
  wire NLW_blk00000347_Q15_UNCONNECTED;
  wire NLW_blk00000349_Q15_UNCONNECTED;
  wire NLW_blk0000034b_Q15_UNCONNECTED;
  wire NLW_blk0000034d_Q15_UNCONNECTED;
  wire NLW_blk0000034f_Q15_UNCONNECTED;
  wire NLW_blk00000351_Q15_UNCONNECTED;
  wire NLW_blk00000353_Q15_UNCONNECTED;
  wire NLW_blk00000355_Q15_UNCONNECTED;
  wire NLW_blk00000357_Q15_UNCONNECTED;
  wire NLW_blk00000359_Q15_UNCONNECTED;
  wire NLW_blk0000035b_Q15_UNCONNECTED;
  wire NLW_blk0000035d_Q15_UNCONNECTED;
  wire NLW_blk0000035f_Q15_UNCONNECTED;
  wire NLW_blk00000361_Q15_UNCONNECTED;
  wire NLW_blk00000363_Q15_UNCONNECTED;
  wire NLW_blk00000365_Q15_UNCONNECTED;
  wire NLW_blk00000367_Q15_UNCONNECTED;
  wire NLW_blk00000369_Q15_UNCONNECTED;
  wire NLW_blk0000036b_Q15_UNCONNECTED;
  wire NLW_blk0000036d_Q15_UNCONNECTED;
  wire NLW_blk0000036f_Q15_UNCONNECTED;
  wire NLW_blk00000371_Q15_UNCONNECTED;
  wire NLW_blk00000373_Q15_UNCONNECTED;
  wire NLW_blk00000375_Q15_UNCONNECTED;
  wire NLW_blk00000377_Q15_UNCONNECTED;
  wire NLW_blk00000379_Q15_UNCONNECTED;
  wire NLW_blk0000037b_Q15_UNCONNECTED;
  wire NLW_blk0000037d_Q15_UNCONNECTED;
  wire NLW_blk0000037f_Q15_UNCONNECTED;
  wire NLW_blk00000381_Q15_UNCONNECTED;
  wire NLW_blk00000383_Q15_UNCONNECTED;
  wire NLW_blk00000385_Q15_UNCONNECTED;
  wire NLW_blk00000387_Q15_UNCONNECTED;
  wire NLW_blk00000389_Q15_UNCONNECTED;
  wire NLW_blk0000038b_Q15_UNCONNECTED;
  wire NLW_blk0000038d_Q15_UNCONNECTED;
  wire NLW_blk0000038f_Q15_UNCONNECTED;
  wire NLW_blk00000391_Q15_UNCONNECTED;
  wire NLW_blk00000393_Q15_UNCONNECTED;
  wire NLW_blk00000395_Q15_UNCONNECTED;
  wire NLW_blk00000397_Q15_UNCONNECTED;
  wire NLW_blk00000399_Q15_UNCONNECTED;
  wire NLW_blk0000039b_Q15_UNCONNECTED;
  wire NLW_blk0000039d_Q15_UNCONNECTED;
  wire NLW_blk0000039f_Q15_UNCONNECTED;
  wire NLW_blk000003a1_Q15_UNCONNECTED;
  wire NLW_blk000003a3_Q15_UNCONNECTED;
  wire NLW_blk000003a5_Q15_UNCONNECTED;
  wire NLW_blk000003a7_Q15_UNCONNECTED;
  wire NLW_blk000003a9_Q15_UNCONNECTED;
  wire NLW_blk000003ab_Q15_UNCONNECTED;
  wire NLW_blk000003ad_Q15_UNCONNECTED;
  wire NLW_blk000003af_Q15_UNCONNECTED;
  wire NLW_blk000003b1_Q15_UNCONNECTED;
  wire NLW_blk000003b3_Q15_UNCONNECTED;
  wire NLW_blk000003b5_Q15_UNCONNECTED;
  wire NLW_blk000003b7_Q15_UNCONNECTED;
  wire NLW_blk000003b9_Q15_UNCONNECTED;
  wire NLW_blk000003bb_Q15_UNCONNECTED;
  wire NLW_blk000003bd_Q15_UNCONNECTED;
  wire NLW_blk000003bf_Q15_UNCONNECTED;
  wire NLW_blk000003c1_Q15_UNCONNECTED;
  wire NLW_blk000003c3_Q15_UNCONNECTED;
  wire NLW_blk000003c5_Q15_UNCONNECTED;
  wire NLW_blk000003c7_Q15_UNCONNECTED;
  wire NLW_blk000003c9_Q15_UNCONNECTED;
  wire NLW_blk000003cb_Q15_UNCONNECTED;
  wire NLW_blk000003cd_Q15_UNCONNECTED;
  wire NLW_blk000003cf_Q15_UNCONNECTED;
  wire NLW_blk000003d1_Q15_UNCONNECTED;
  wire NLW_blk000003d3_Q15_UNCONNECTED;
  wire NLW_blk000003d5_Q15_UNCONNECTED;
  wire NLW_blk000003d7_Q15_UNCONNECTED;
  wire NLW_blk000003d9_Q15_UNCONNECTED;
  wire NLW_blk000003db_Q15_UNCONNECTED;
  wire NLW_blk000003dd_Q15_UNCONNECTED;
  wire NLW_blk000003df_Q15_UNCONNECTED;
  wire NLW_blk000003e1_Q15_UNCONNECTED;
  wire NLW_blk000003e3_Q15_UNCONNECTED;
  wire NLW_blk000003e5_Q15_UNCONNECTED;
  wire NLW_blk000003e7_Q15_UNCONNECTED;
  wire NLW_blk000003e9_Q15_UNCONNECTED;
  wire NLW_blk000003eb_Q15_UNCONNECTED;
  wire NLW_blk000003ed_Q15_UNCONNECTED;
  wire NLW_blk000003ef_Q15_UNCONNECTED;
  wire NLW_blk000003f1_Q15_UNCONNECTED;
  wire NLW_blk000003f3_Q15_UNCONNECTED;
  wire NLW_blk000003f5_Q15_UNCONNECTED;
  wire NLW_blk000003f7_Q15_UNCONNECTED;
  wire NLW_blk000003f9_Q15_UNCONNECTED;
  wire NLW_blk000003fb_Q15_UNCONNECTED;
  wire NLW_blk000003fd_Q15_UNCONNECTED;
  wire NLW_blk000003ff_Q15_UNCONNECTED;
  wire NLW_blk00000401_Q15_UNCONNECTED;
  wire NLW_blk00000403_Q15_UNCONNECTED;
  wire NLW_blk00000405_Q15_UNCONNECTED;
  wire NLW_blk00000407_Q15_UNCONNECTED;
  wire NLW_blk00000409_Q15_UNCONNECTED;
  wire NLW_blk0000040b_Q15_UNCONNECTED;
  wire \NLW_blk0000040d_PCOUT<47>_UNCONNECTED ;
  wire \NLW_blk0000040d_PCOUT<46>_UNCONNECTED ;
  wire \NLW_blk0000040d_PCOUT<45>_UNCONNECTED ;
  wire \NLW_blk0000040d_PCOUT<44>_UNCONNECTED ;
  wire \NLW_blk0000040d_PCOUT<43>_UNCONNECTED ;
  wire \NLW_blk0000040d_PCOUT<42>_UNCONNECTED ;
  wire \NLW_blk0000040d_PCOUT<41>_UNCONNECTED ;
  wire \NLW_blk0000040d_PCOUT<40>_UNCONNECTED ;
  wire \NLW_blk0000040d_PCOUT<39>_UNCONNECTED ;
  wire \NLW_blk0000040d_PCOUT<38>_UNCONNECTED ;
  wire \NLW_blk0000040d_PCOUT<37>_UNCONNECTED ;
  wire \NLW_blk0000040d_PCOUT<36>_UNCONNECTED ;
  wire \NLW_blk0000040d_PCOUT<35>_UNCONNECTED ;
  wire \NLW_blk0000040d_PCOUT<34>_UNCONNECTED ;
  wire \NLW_blk0000040d_PCOUT<33>_UNCONNECTED ;
  wire \NLW_blk0000040d_PCOUT<32>_UNCONNECTED ;
  wire \NLW_blk0000040d_PCOUT<31>_UNCONNECTED ;
  wire \NLW_blk0000040d_PCOUT<30>_UNCONNECTED ;
  wire \NLW_blk0000040d_PCOUT<29>_UNCONNECTED ;
  wire \NLW_blk0000040d_PCOUT<28>_UNCONNECTED ;
  wire \NLW_blk0000040d_PCOUT<27>_UNCONNECTED ;
  wire \NLW_blk0000040d_PCOUT<26>_UNCONNECTED ;
  wire \NLW_blk0000040d_PCOUT<25>_UNCONNECTED ;
  wire \NLW_blk0000040d_PCOUT<24>_UNCONNECTED ;
  wire \NLW_blk0000040d_PCOUT<23>_UNCONNECTED ;
  wire \NLW_blk0000040d_PCOUT<22>_UNCONNECTED ;
  wire \NLW_blk0000040d_PCOUT<21>_UNCONNECTED ;
  wire \NLW_blk0000040d_PCOUT<20>_UNCONNECTED ;
  wire \NLW_blk0000040d_PCOUT<19>_UNCONNECTED ;
  wire \NLW_blk0000040d_PCOUT<18>_UNCONNECTED ;
  wire \NLW_blk0000040d_PCOUT<17>_UNCONNECTED ;
  wire \NLW_blk0000040d_PCOUT<16>_UNCONNECTED ;
  wire \NLW_blk0000040d_PCOUT<15>_UNCONNECTED ;
  wire \NLW_blk0000040d_PCOUT<14>_UNCONNECTED ;
  wire \NLW_blk0000040d_PCOUT<13>_UNCONNECTED ;
  wire \NLW_blk0000040d_PCOUT<12>_UNCONNECTED ;
  wire \NLW_blk0000040d_PCOUT<11>_UNCONNECTED ;
  wire \NLW_blk0000040d_PCOUT<10>_UNCONNECTED ;
  wire \NLW_blk0000040d_PCOUT<9>_UNCONNECTED ;
  wire \NLW_blk0000040d_PCOUT<8>_UNCONNECTED ;
  wire \NLW_blk0000040d_PCOUT<7>_UNCONNECTED ;
  wire \NLW_blk0000040d_PCOUT<6>_UNCONNECTED ;
  wire \NLW_blk0000040d_PCOUT<5>_UNCONNECTED ;
  wire \NLW_blk0000040d_PCOUT<4>_UNCONNECTED ;
  wire \NLW_blk0000040d_PCOUT<3>_UNCONNECTED ;
  wire \NLW_blk0000040d_PCOUT<2>_UNCONNECTED ;
  wire \NLW_blk0000040d_PCOUT<1>_UNCONNECTED ;
  wire \NLW_blk0000040d_PCOUT<0>_UNCONNECTED ;
  wire NLW_blk0000040d_PATTERNBDETECT_UNCONNECTED;
  wire NLW_blk0000040d_MULTSIGNOUT_UNCONNECTED;
  wire NLW_blk0000040d_CARRYCASCOUT_UNCONNECTED;
  wire NLW_blk0000040d_UNDERFLOW_UNCONNECTED;
  wire NLW_blk0000040d_PATTERNDETECT_UNCONNECTED;
  wire NLW_blk0000040d_OVERFLOW_UNCONNECTED;
  wire \NLW_blk0000040d_ACOUT<29>_UNCONNECTED ;
  wire \NLW_blk0000040d_ACOUT<28>_UNCONNECTED ;
  wire \NLW_blk0000040d_ACOUT<27>_UNCONNECTED ;
  wire \NLW_blk0000040d_ACOUT<26>_UNCONNECTED ;
  wire \NLW_blk0000040d_ACOUT<25>_UNCONNECTED ;
  wire \NLW_blk0000040d_ACOUT<24>_UNCONNECTED ;
  wire \NLW_blk0000040d_ACOUT<23>_UNCONNECTED ;
  wire \NLW_blk0000040d_ACOUT<22>_UNCONNECTED ;
  wire \NLW_blk0000040d_ACOUT<21>_UNCONNECTED ;
  wire \NLW_blk0000040d_ACOUT<20>_UNCONNECTED ;
  wire \NLW_blk0000040d_ACOUT<19>_UNCONNECTED ;
  wire \NLW_blk0000040d_ACOUT<18>_UNCONNECTED ;
  wire \NLW_blk0000040d_ACOUT<17>_UNCONNECTED ;
  wire \NLW_blk0000040d_ACOUT<16>_UNCONNECTED ;
  wire \NLW_blk0000040d_ACOUT<15>_UNCONNECTED ;
  wire \NLW_blk0000040d_ACOUT<14>_UNCONNECTED ;
  wire \NLW_blk0000040d_ACOUT<13>_UNCONNECTED ;
  wire \NLW_blk0000040d_ACOUT<12>_UNCONNECTED ;
  wire \NLW_blk0000040d_ACOUT<11>_UNCONNECTED ;
  wire \NLW_blk0000040d_ACOUT<10>_UNCONNECTED ;
  wire \NLW_blk0000040d_ACOUT<9>_UNCONNECTED ;
  wire \NLW_blk0000040d_ACOUT<8>_UNCONNECTED ;
  wire \NLW_blk0000040d_ACOUT<7>_UNCONNECTED ;
  wire \NLW_blk0000040d_ACOUT<6>_UNCONNECTED ;
  wire \NLW_blk0000040d_ACOUT<5>_UNCONNECTED ;
  wire \NLW_blk0000040d_ACOUT<4>_UNCONNECTED ;
  wire \NLW_blk0000040d_ACOUT<3>_UNCONNECTED ;
  wire \NLW_blk0000040d_ACOUT<2>_UNCONNECTED ;
  wire \NLW_blk0000040d_ACOUT<1>_UNCONNECTED ;
  wire \NLW_blk0000040d_ACOUT<0>_UNCONNECTED ;
  wire \NLW_blk0000040d_CARRYOUT<3>_UNCONNECTED ;
  wire \NLW_blk0000040d_CARRYOUT<2>_UNCONNECTED ;
  wire \NLW_blk0000040d_CARRYOUT<1>_UNCONNECTED ;
  wire \NLW_blk0000040d_CARRYOUT<0>_UNCONNECTED ;
  wire \NLW_blk0000040d_BCOUT<17>_UNCONNECTED ;
  wire \NLW_blk0000040d_BCOUT<16>_UNCONNECTED ;
  wire \NLW_blk0000040d_BCOUT<15>_UNCONNECTED ;
  wire \NLW_blk0000040d_BCOUT<14>_UNCONNECTED ;
  wire \NLW_blk0000040d_BCOUT<13>_UNCONNECTED ;
  wire \NLW_blk0000040d_BCOUT<12>_UNCONNECTED ;
  wire \NLW_blk0000040d_BCOUT<11>_UNCONNECTED ;
  wire \NLW_blk0000040d_BCOUT<10>_UNCONNECTED ;
  wire \NLW_blk0000040d_BCOUT<9>_UNCONNECTED ;
  wire \NLW_blk0000040d_BCOUT<8>_UNCONNECTED ;
  wire \NLW_blk0000040d_BCOUT<7>_UNCONNECTED ;
  wire \NLW_blk0000040d_BCOUT<6>_UNCONNECTED ;
  wire \NLW_blk0000040d_BCOUT<5>_UNCONNECTED ;
  wire \NLW_blk0000040d_BCOUT<4>_UNCONNECTED ;
  wire \NLW_blk0000040d_BCOUT<3>_UNCONNECTED ;
  wire \NLW_blk0000040d_BCOUT<2>_UNCONNECTED ;
  wire \NLW_blk0000040d_BCOUT<1>_UNCONNECTED ;
  wire \NLW_blk0000040d_BCOUT<0>_UNCONNECTED ;
  wire \NLW_blk0000040d_P<47>_UNCONNECTED ;
  wire \NLW_blk0000040d_P<46>_UNCONNECTED ;
  wire \NLW_blk0000040d_P<45>_UNCONNECTED ;
  wire \NLW_blk0000040d_P<44>_UNCONNECTED ;
  wire \NLW_blk0000040d_P<43>_UNCONNECTED ;
  wire \NLW_blk0000040d_P<42>_UNCONNECTED ;
  wire \NLW_blk0000040d_P<41>_UNCONNECTED ;
  wire \NLW_blk0000040d_P<40>_UNCONNECTED ;
  wire \NLW_blk0000040d_P<39>_UNCONNECTED ;
  wire \NLW_blk0000040d_P<38>_UNCONNECTED ;
  wire \NLW_blk0000040d_P<37>_UNCONNECTED ;
  wire \NLW_blk0000040d_P<36>_UNCONNECTED ;
  wire \NLW_blk0000040d_P<35>_UNCONNECTED ;
  wire \NLW_blk0000040d_P<34>_UNCONNECTED ;
  wire \NLW_blk0000040d_P<33>_UNCONNECTED ;
  wire \NLW_blk0000040d_P<32>_UNCONNECTED ;
  wire \NLW_blk0000040d_P<31>_UNCONNECTED ;
  wire \NLW_blk0000040d_P<30>_UNCONNECTED ;
  wire \NLW_blk0000040d_P<29>_UNCONNECTED ;
  wire \NLW_blk0000040d_P<28>_UNCONNECTED ;
  wire \NLW_blk0000040d_P<27>_UNCONNECTED ;
  wire \NLW_blk0000040d_P<26>_UNCONNECTED ;
  wire \NLW_blk0000040d_P<25>_UNCONNECTED ;
  wire \NLW_blk0000040d_P<24>_UNCONNECTED ;
  wire \NLW_blk0000040d_P<23>_UNCONNECTED ;
  wire \NLW_blk0000040d_P<22>_UNCONNECTED ;
  wire \NLW_blk0000040d_P<21>_UNCONNECTED ;
  wire NLW_blk0000040e_PATTERNBDETECT_UNCONNECTED;
  wire NLW_blk0000040e_MULTSIGNOUT_UNCONNECTED;
  wire NLW_blk0000040e_CARRYCASCOUT_UNCONNECTED;
  wire NLW_blk0000040e_UNDERFLOW_UNCONNECTED;
  wire NLW_blk0000040e_PATTERNDETECT_UNCONNECTED;
  wire NLW_blk0000040e_OVERFLOW_UNCONNECTED;
  wire \NLW_blk0000040e_CARRYOUT<3>_UNCONNECTED ;
  wire \NLW_blk0000040e_CARRYOUT<2>_UNCONNECTED ;
  wire \NLW_blk0000040e_CARRYOUT<1>_UNCONNECTED ;
  wire \NLW_blk0000040e_CARRYOUT<0>_UNCONNECTED ;
  wire \NLW_blk0000040e_BCOUT<17>_UNCONNECTED ;
  wire \NLW_blk0000040e_BCOUT<16>_UNCONNECTED ;
  wire \NLW_blk0000040e_BCOUT<15>_UNCONNECTED ;
  wire \NLW_blk0000040e_BCOUT<14>_UNCONNECTED ;
  wire \NLW_blk0000040e_BCOUT<13>_UNCONNECTED ;
  wire \NLW_blk0000040e_BCOUT<12>_UNCONNECTED ;
  wire \NLW_blk0000040e_BCOUT<11>_UNCONNECTED ;
  wire \NLW_blk0000040e_BCOUT<10>_UNCONNECTED ;
  wire \NLW_blk0000040e_BCOUT<9>_UNCONNECTED ;
  wire \NLW_blk0000040e_BCOUT<8>_UNCONNECTED ;
  wire \NLW_blk0000040e_BCOUT<7>_UNCONNECTED ;
  wire \NLW_blk0000040e_BCOUT<6>_UNCONNECTED ;
  wire \NLW_blk0000040e_BCOUT<5>_UNCONNECTED ;
  wire \NLW_blk0000040e_BCOUT<4>_UNCONNECTED ;
  wire \NLW_blk0000040e_BCOUT<3>_UNCONNECTED ;
  wire \NLW_blk0000040e_BCOUT<2>_UNCONNECTED ;
  wire \NLW_blk0000040e_BCOUT<1>_UNCONNECTED ;
  wire \NLW_blk0000040e_BCOUT<0>_UNCONNECTED ;
  wire \NLW_blk0000040e_P<47>_UNCONNECTED ;
  wire \NLW_blk0000040e_P<46>_UNCONNECTED ;
  wire \NLW_blk0000040e_P<45>_UNCONNECTED ;
  wire \NLW_blk0000040e_P<44>_UNCONNECTED ;
  wire \NLW_blk0000040e_P<43>_UNCONNECTED ;
  wire \NLW_blk0000040e_P<42>_UNCONNECTED ;
  wire \NLW_blk0000040e_P<41>_UNCONNECTED ;
  wire \NLW_blk0000040e_P<40>_UNCONNECTED ;
  wire \NLW_blk0000040e_P<39>_UNCONNECTED ;
  wire \NLW_blk0000040e_P<38>_UNCONNECTED ;
  wire \NLW_blk0000040e_P<37>_UNCONNECTED ;
  wire \NLW_blk0000040e_P<36>_UNCONNECTED ;
  wire \NLW_blk0000040e_P<35>_UNCONNECTED ;
  wire \NLW_blk0000040e_P<34>_UNCONNECTED ;
  wire \NLW_blk0000040e_P<33>_UNCONNECTED ;
  wire \NLW_blk0000040e_P<32>_UNCONNECTED ;
  wire \NLW_blk0000040e_P<31>_UNCONNECTED ;
  wire \NLW_blk0000040e_P<30>_UNCONNECTED ;
  wire \NLW_blk0000040e_P<29>_UNCONNECTED ;
  wire \NLW_blk0000040e_P<28>_UNCONNECTED ;
  wire \NLW_blk0000040e_P<27>_UNCONNECTED ;
  wire \NLW_blk0000040e_P<26>_UNCONNECTED ;
  wire \NLW_blk0000040e_P<25>_UNCONNECTED ;
  wire \NLW_blk0000040e_P<24>_UNCONNECTED ;
  wire \NLW_blk0000040e_P<23>_UNCONNECTED ;
  wire \NLW_blk0000040e_P<22>_UNCONNECTED ;
  wire \NLW_blk0000040e_P<21>_UNCONNECTED ;
  wire \NLW_blk0000040e_P<20>_UNCONNECTED ;
  wire \NLW_blk0000040e_P<19>_UNCONNECTED ;
  wire \NLW_blk0000040e_P<18>_UNCONNECTED ;
  wire \NLW_blk0000040e_P<17>_UNCONNECTED ;
  wire NLW_blk0000040f_PATTERNBDETECT_UNCONNECTED;
  wire NLW_blk0000040f_MULTSIGNOUT_UNCONNECTED;
  wire NLW_blk0000040f_CARRYCASCOUT_UNCONNECTED;
  wire NLW_blk0000040f_UNDERFLOW_UNCONNECTED;
  wire NLW_blk0000040f_PATTERNDETECT_UNCONNECTED;
  wire NLW_blk0000040f_OVERFLOW_UNCONNECTED;
  wire \NLW_blk0000040f_CARRYOUT<3>_UNCONNECTED ;
  wire \NLW_blk0000040f_CARRYOUT<2>_UNCONNECTED ;
  wire \NLW_blk0000040f_CARRYOUT<1>_UNCONNECTED ;
  wire \NLW_blk0000040f_CARRYOUT<0>_UNCONNECTED ;
  wire \NLW_blk0000040f_BCOUT<17>_UNCONNECTED ;
  wire \NLW_blk0000040f_BCOUT<16>_UNCONNECTED ;
  wire \NLW_blk0000040f_BCOUT<15>_UNCONNECTED ;
  wire \NLW_blk0000040f_BCOUT<14>_UNCONNECTED ;
  wire \NLW_blk0000040f_BCOUT<13>_UNCONNECTED ;
  wire \NLW_blk0000040f_BCOUT<12>_UNCONNECTED ;
  wire \NLW_blk0000040f_BCOUT<11>_UNCONNECTED ;
  wire \NLW_blk0000040f_BCOUT<10>_UNCONNECTED ;
  wire \NLW_blk0000040f_BCOUT<9>_UNCONNECTED ;
  wire \NLW_blk0000040f_BCOUT<8>_UNCONNECTED ;
  wire \NLW_blk0000040f_BCOUT<7>_UNCONNECTED ;
  wire \NLW_blk0000040f_BCOUT<6>_UNCONNECTED ;
  wire \NLW_blk0000040f_BCOUT<5>_UNCONNECTED ;
  wire \NLW_blk0000040f_BCOUT<4>_UNCONNECTED ;
  wire \NLW_blk0000040f_BCOUT<3>_UNCONNECTED ;
  wire \NLW_blk0000040f_BCOUT<2>_UNCONNECTED ;
  wire \NLW_blk0000040f_BCOUT<1>_UNCONNECTED ;
  wire \NLW_blk0000040f_BCOUT<0>_UNCONNECTED ;
  wire \NLW_blk0000040f_P<47>_UNCONNECTED ;
  wire \NLW_blk0000040f_P<46>_UNCONNECTED ;
  wire \NLW_blk0000040f_P<45>_UNCONNECTED ;
  wire \NLW_blk0000040f_P<44>_UNCONNECTED ;
  wire \NLW_blk0000040f_P<43>_UNCONNECTED ;
  wire \NLW_blk0000040f_P<42>_UNCONNECTED ;
  wire \NLW_blk0000040f_P<41>_UNCONNECTED ;
  wire \NLW_blk0000040f_P<40>_UNCONNECTED ;
  wire \NLW_blk0000040f_P<39>_UNCONNECTED ;
  wire \NLW_blk0000040f_P<38>_UNCONNECTED ;
  wire \NLW_blk0000040f_P<37>_UNCONNECTED ;
  wire \NLW_blk0000040f_P<36>_UNCONNECTED ;
  wire \NLW_blk0000040f_P<35>_UNCONNECTED ;
  wire \NLW_blk0000040f_P<34>_UNCONNECTED ;
  wire \NLW_blk0000040f_P<33>_UNCONNECTED ;
  wire \NLW_blk0000040f_P<32>_UNCONNECTED ;
  wire \NLW_blk0000040f_P<31>_UNCONNECTED ;
  wire \NLW_blk0000040f_P<30>_UNCONNECTED ;
  wire \NLW_blk0000040f_P<29>_UNCONNECTED ;
  wire \NLW_blk0000040f_P<28>_UNCONNECTED ;
  wire \NLW_blk0000040f_P<27>_UNCONNECTED ;
  wire \NLW_blk0000040f_P<26>_UNCONNECTED ;
  wire \NLW_blk0000040f_P<25>_UNCONNECTED ;
  wire \NLW_blk0000040f_P<24>_UNCONNECTED ;
  wire \NLW_blk0000040f_P<23>_UNCONNECTED ;
  wire \NLW_blk0000040f_P<22>_UNCONNECTED ;
  wire \NLW_blk0000040f_P<21>_UNCONNECTED ;
  wire \NLW_blk0000040f_P<20>_UNCONNECTED ;
  wire \NLW_blk0000040f_P<19>_UNCONNECTED ;
  wire \NLW_blk0000040f_P<18>_UNCONNECTED ;
  wire \NLW_blk0000040f_P<17>_UNCONNECTED ;
  wire NLW_blk00000410_PATTERNBDETECT_UNCONNECTED;
  wire NLW_blk00000410_MULTSIGNOUT_UNCONNECTED;
  wire NLW_blk00000410_CARRYCASCOUT_UNCONNECTED;
  wire NLW_blk00000410_UNDERFLOW_UNCONNECTED;
  wire NLW_blk00000410_PATTERNDETECT_UNCONNECTED;
  wire NLW_blk00000410_OVERFLOW_UNCONNECTED;
  wire \NLW_blk00000410_ACOUT<29>_UNCONNECTED ;
  wire \NLW_blk00000410_ACOUT<28>_UNCONNECTED ;
  wire \NLW_blk00000410_ACOUT<27>_UNCONNECTED ;
  wire \NLW_blk00000410_ACOUT<26>_UNCONNECTED ;
  wire \NLW_blk00000410_ACOUT<25>_UNCONNECTED ;
  wire \NLW_blk00000410_ACOUT<24>_UNCONNECTED ;
  wire \NLW_blk00000410_ACOUT<23>_UNCONNECTED ;
  wire \NLW_blk00000410_ACOUT<22>_UNCONNECTED ;
  wire \NLW_blk00000410_ACOUT<21>_UNCONNECTED ;
  wire \NLW_blk00000410_ACOUT<20>_UNCONNECTED ;
  wire \NLW_blk00000410_ACOUT<19>_UNCONNECTED ;
  wire \NLW_blk00000410_ACOUT<18>_UNCONNECTED ;
  wire \NLW_blk00000410_ACOUT<17>_UNCONNECTED ;
  wire \NLW_blk00000410_ACOUT<16>_UNCONNECTED ;
  wire \NLW_blk00000410_ACOUT<15>_UNCONNECTED ;
  wire \NLW_blk00000410_ACOUT<14>_UNCONNECTED ;
  wire \NLW_blk00000410_ACOUT<13>_UNCONNECTED ;
  wire \NLW_blk00000410_ACOUT<12>_UNCONNECTED ;
  wire \NLW_blk00000410_ACOUT<11>_UNCONNECTED ;
  wire \NLW_blk00000410_ACOUT<10>_UNCONNECTED ;
  wire \NLW_blk00000410_ACOUT<9>_UNCONNECTED ;
  wire \NLW_blk00000410_ACOUT<8>_UNCONNECTED ;
  wire \NLW_blk00000410_ACOUT<7>_UNCONNECTED ;
  wire \NLW_blk00000410_ACOUT<6>_UNCONNECTED ;
  wire \NLW_blk00000410_ACOUT<5>_UNCONNECTED ;
  wire \NLW_blk00000410_ACOUT<4>_UNCONNECTED ;
  wire \NLW_blk00000410_ACOUT<3>_UNCONNECTED ;
  wire \NLW_blk00000410_ACOUT<2>_UNCONNECTED ;
  wire \NLW_blk00000410_ACOUT<1>_UNCONNECTED ;
  wire \NLW_blk00000410_ACOUT<0>_UNCONNECTED ;
  wire \NLW_blk00000410_CARRYOUT<3>_UNCONNECTED ;
  wire \NLW_blk00000410_CARRYOUT<2>_UNCONNECTED ;
  wire \NLW_blk00000410_CARRYOUT<1>_UNCONNECTED ;
  wire \NLW_blk00000410_CARRYOUT<0>_UNCONNECTED ;
  wire \NLW_blk00000410_BCOUT<17>_UNCONNECTED ;
  wire \NLW_blk00000410_BCOUT<16>_UNCONNECTED ;
  wire \NLW_blk00000410_BCOUT<15>_UNCONNECTED ;
  wire \NLW_blk00000410_BCOUT<14>_UNCONNECTED ;
  wire \NLW_blk00000410_BCOUT<13>_UNCONNECTED ;
  wire \NLW_blk00000410_BCOUT<12>_UNCONNECTED ;
  wire \NLW_blk00000410_BCOUT<11>_UNCONNECTED ;
  wire \NLW_blk00000410_BCOUT<10>_UNCONNECTED ;
  wire \NLW_blk00000410_BCOUT<9>_UNCONNECTED ;
  wire \NLW_blk00000410_BCOUT<8>_UNCONNECTED ;
  wire \NLW_blk00000410_BCOUT<7>_UNCONNECTED ;
  wire \NLW_blk00000410_BCOUT<6>_UNCONNECTED ;
  wire \NLW_blk00000410_BCOUT<5>_UNCONNECTED ;
  wire \NLW_blk00000410_BCOUT<4>_UNCONNECTED ;
  wire \NLW_blk00000410_BCOUT<3>_UNCONNECTED ;
  wire \NLW_blk00000410_BCOUT<2>_UNCONNECTED ;
  wire \NLW_blk00000410_BCOUT<1>_UNCONNECTED ;
  wire \NLW_blk00000410_BCOUT<0>_UNCONNECTED ;
  wire \NLW_blk00000410_P<47>_UNCONNECTED ;
  wire \NLW_blk00000410_P<46>_UNCONNECTED ;
  wire \NLW_blk00000410_P<45>_UNCONNECTED ;
  wire \NLW_blk00000410_P<44>_UNCONNECTED ;
  wire \NLW_blk00000410_P<43>_UNCONNECTED ;
  wire \NLW_blk00000410_P<42>_UNCONNECTED ;
  wire \NLW_blk00000410_P<41>_UNCONNECTED ;
  wire \NLW_blk00000410_P<40>_UNCONNECTED ;
  wire \NLW_blk00000410_P<39>_UNCONNECTED ;
  wire \NLW_blk00000410_P<38>_UNCONNECTED ;
  wire \NLW_blk00000410_P<37>_UNCONNECTED ;
  wire \NLW_blk00000410_P<36>_UNCONNECTED ;
  wire \NLW_blk00000410_P<35>_UNCONNECTED ;
  wire \NLW_blk00000410_P<34>_UNCONNECTED ;
  wire \NLW_blk00000410_P<33>_UNCONNECTED ;
  wire \NLW_blk00000410_P<32>_UNCONNECTED ;
  wire \NLW_blk00000410_P<31>_UNCONNECTED ;
  wire \NLW_blk00000410_P<30>_UNCONNECTED ;
  wire \NLW_blk00000410_P<29>_UNCONNECTED ;
  wire \NLW_blk00000410_P<28>_UNCONNECTED ;
  wire \NLW_blk00000410_P<27>_UNCONNECTED ;
  wire \NLW_blk00000410_P<26>_UNCONNECTED ;
  wire \NLW_blk00000410_P<25>_UNCONNECTED ;
  wire \NLW_blk00000410_P<24>_UNCONNECTED ;
  wire \NLW_blk00000410_P<23>_UNCONNECTED ;
  wire \NLW_blk00000410_P<22>_UNCONNECTED ;
  wire \NLW_blk00000410_P<21>_UNCONNECTED ;
  wire \NLW_blk00000410_P<20>_UNCONNECTED ;
  wire \NLW_blk00000410_P<19>_UNCONNECTED ;
  wire \NLW_blk00000410_P<18>_UNCONNECTED ;
  wire \NLW_blk00000410_P<17>_UNCONNECTED ;
  wire \NLW_blk00000410_P<16>_UNCONNECTED ;
  wire \NLW_blk00000410_P<15>_UNCONNECTED ;
  wire \NLW_blk00000410_P<14>_UNCONNECTED ;
  wire \NLW_blk00000410_P<13>_UNCONNECTED ;
  wire \NLW_blk00000410_P<12>_UNCONNECTED ;
  wire \NLW_blk00000410_P<11>_UNCONNECTED ;
  wire \NLW_blk00000410_P<10>_UNCONNECTED ;
  wire \NLW_blk00000410_P<9>_UNCONNECTED ;
  wire \NLW_blk00000410_P<8>_UNCONNECTED ;
  wire \NLW_blk00000410_P<7>_UNCONNECTED ;
  wire \NLW_blk00000410_P<6>_UNCONNECTED ;
  wire \NLW_blk00000410_P<5>_UNCONNECTED ;
  wire \NLW_blk00000410_P<4>_UNCONNECTED ;
  wire \NLW_blk00000410_P<3>_UNCONNECTED ;
  wire \NLW_blk00000410_P<2>_UNCONNECTED ;
  wire \NLW_blk00000410_P<1>_UNCONNECTED ;
  wire \NLW_blk00000410_P<0>_UNCONNECTED ;
  wire NLW_blk00000411_PATTERNBDETECT_UNCONNECTED;
  wire NLW_blk00000411_MULTSIGNOUT_UNCONNECTED;
  wire NLW_blk00000411_CARRYCASCOUT_UNCONNECTED;
  wire NLW_blk00000411_UNDERFLOW_UNCONNECTED;
  wire NLW_blk00000411_OVERFLOW_UNCONNECTED;
  wire \NLW_blk00000411_CARRYOUT<3>_UNCONNECTED ;
  wire \NLW_blk00000411_CARRYOUT<2>_UNCONNECTED ;
  wire \NLW_blk00000411_CARRYOUT<1>_UNCONNECTED ;
  wire \NLW_blk00000411_CARRYOUT<0>_UNCONNECTED ;
  wire \NLW_blk00000411_BCOUT<17>_UNCONNECTED ;
  wire \NLW_blk00000411_BCOUT<16>_UNCONNECTED ;
  wire \NLW_blk00000411_BCOUT<15>_UNCONNECTED ;
  wire \NLW_blk00000411_BCOUT<14>_UNCONNECTED ;
  wire \NLW_blk00000411_BCOUT<13>_UNCONNECTED ;
  wire \NLW_blk00000411_BCOUT<12>_UNCONNECTED ;
  wire \NLW_blk00000411_BCOUT<11>_UNCONNECTED ;
  wire \NLW_blk00000411_BCOUT<10>_UNCONNECTED ;
  wire \NLW_blk00000411_BCOUT<9>_UNCONNECTED ;
  wire \NLW_blk00000411_BCOUT<8>_UNCONNECTED ;
  wire \NLW_blk00000411_BCOUT<7>_UNCONNECTED ;
  wire \NLW_blk00000411_BCOUT<6>_UNCONNECTED ;
  wire \NLW_blk00000411_BCOUT<5>_UNCONNECTED ;
  wire \NLW_blk00000411_BCOUT<4>_UNCONNECTED ;
  wire \NLW_blk00000411_BCOUT<3>_UNCONNECTED ;
  wire \NLW_blk00000411_BCOUT<2>_UNCONNECTED ;
  wire \NLW_blk00000411_BCOUT<1>_UNCONNECTED ;
  wire \NLW_blk00000411_BCOUT<0>_UNCONNECTED ;
  wire \NLW_blk00000411_P<47>_UNCONNECTED ;
  wire \NLW_blk00000411_P<46>_UNCONNECTED ;
  wire \NLW_blk00000411_P<45>_UNCONNECTED ;
  wire \NLW_blk00000411_P<44>_UNCONNECTED ;
  wire \NLW_blk00000411_P<43>_UNCONNECTED ;
  wire \NLW_blk00000411_P<42>_UNCONNECTED ;
  wire \NLW_blk00000411_P<41>_UNCONNECTED ;
  wire \NLW_blk00000411_P<40>_UNCONNECTED ;
  wire \NLW_blk00000411_P<39>_UNCONNECTED ;
  wire \NLW_blk00000411_P<38>_UNCONNECTED ;
  wire \NLW_blk00000411_P<37>_UNCONNECTED ;
  wire \NLW_blk00000411_P<36>_UNCONNECTED ;
  wire \NLW_blk00000411_P<35>_UNCONNECTED ;
  wire \NLW_blk00000411_P<34>_UNCONNECTED ;
  wire \NLW_blk00000411_P<33>_UNCONNECTED ;
  wire \NLW_blk00000411_P<32>_UNCONNECTED ;
  wire \NLW_blk00000411_P<31>_UNCONNECTED ;
  wire \NLW_blk00000411_P<30>_UNCONNECTED ;
  wire \NLW_blk00000411_P<29>_UNCONNECTED ;
  wire \NLW_blk00000411_P<28>_UNCONNECTED ;
  wire \NLW_blk00000411_P<27>_UNCONNECTED ;
  wire \NLW_blk00000411_P<26>_UNCONNECTED ;
  wire \NLW_blk00000411_P<25>_UNCONNECTED ;
  wire \NLW_blk00000411_P<24>_UNCONNECTED ;
  wire \NLW_blk00000411_P<23>_UNCONNECTED ;
  wire \NLW_blk00000411_P<22>_UNCONNECTED ;
  wire \NLW_blk00000411_P<21>_UNCONNECTED ;
  wire \NLW_blk00000411_P<20>_UNCONNECTED ;
  wire \NLW_blk00000411_P<19>_UNCONNECTED ;
  wire \NLW_blk00000411_P<18>_UNCONNECTED ;
  wire \NLW_blk00000411_P<17>_UNCONNECTED ;
  wire \NLW_blk00000411_P<16>_UNCONNECTED ;
  wire \NLW_blk00000411_P<15>_UNCONNECTED ;
  wire \NLW_blk00000411_P<14>_UNCONNECTED ;
  wire \NLW_blk00000411_P<13>_UNCONNECTED ;
  wire \NLW_blk00000411_P<12>_UNCONNECTED ;
  wire \NLW_blk00000411_P<11>_UNCONNECTED ;
  wire \NLW_blk00000411_P<10>_UNCONNECTED ;
  wire \NLW_blk00000411_P<9>_UNCONNECTED ;
  wire \NLW_blk00000411_P<8>_UNCONNECTED ;
  wire \NLW_blk00000411_P<7>_UNCONNECTED ;
  wire \NLW_blk00000411_P<6>_UNCONNECTED ;
  wire \NLW_blk00000411_P<5>_UNCONNECTED ;
  wire \NLW_blk00000411_P<4>_UNCONNECTED ;
  wire \NLW_blk00000411_P<3>_UNCONNECTED ;
  wire \NLW_blk00000411_P<2>_UNCONNECTED ;
  wire \NLW_blk00000411_P<1>_UNCONNECTED ;
  wire \NLW_blk00000411_P<0>_UNCONNECTED ;
  wire NLW_blk00000412_PATTERNBDETECT_UNCONNECTED;
  wire NLW_blk00000412_MULTSIGNOUT_UNCONNECTED;
  wire NLW_blk00000412_CARRYCASCOUT_UNCONNECTED;
  wire NLW_blk00000412_UNDERFLOW_UNCONNECTED;
  wire NLW_blk00000412_PATTERNDETECT_UNCONNECTED;
  wire NLW_blk00000412_OVERFLOW_UNCONNECTED;
  wire \NLW_blk00000412_ACOUT<29>_UNCONNECTED ;
  wire \NLW_blk00000412_ACOUT<28>_UNCONNECTED ;
  wire \NLW_blk00000412_ACOUT<27>_UNCONNECTED ;
  wire \NLW_blk00000412_ACOUT<26>_UNCONNECTED ;
  wire \NLW_blk00000412_ACOUT<25>_UNCONNECTED ;
  wire \NLW_blk00000412_ACOUT<24>_UNCONNECTED ;
  wire \NLW_blk00000412_ACOUT<23>_UNCONNECTED ;
  wire \NLW_blk00000412_ACOUT<22>_UNCONNECTED ;
  wire \NLW_blk00000412_ACOUT<21>_UNCONNECTED ;
  wire \NLW_blk00000412_ACOUT<20>_UNCONNECTED ;
  wire \NLW_blk00000412_ACOUT<19>_UNCONNECTED ;
  wire \NLW_blk00000412_ACOUT<18>_UNCONNECTED ;
  wire \NLW_blk00000412_ACOUT<17>_UNCONNECTED ;
  wire \NLW_blk00000412_ACOUT<16>_UNCONNECTED ;
  wire \NLW_blk00000412_ACOUT<15>_UNCONNECTED ;
  wire \NLW_blk00000412_ACOUT<14>_UNCONNECTED ;
  wire \NLW_blk00000412_ACOUT<13>_UNCONNECTED ;
  wire \NLW_blk00000412_ACOUT<12>_UNCONNECTED ;
  wire \NLW_blk00000412_ACOUT<11>_UNCONNECTED ;
  wire \NLW_blk00000412_ACOUT<10>_UNCONNECTED ;
  wire \NLW_blk00000412_ACOUT<9>_UNCONNECTED ;
  wire \NLW_blk00000412_ACOUT<8>_UNCONNECTED ;
  wire \NLW_blk00000412_ACOUT<7>_UNCONNECTED ;
  wire \NLW_blk00000412_ACOUT<6>_UNCONNECTED ;
  wire \NLW_blk00000412_ACOUT<5>_UNCONNECTED ;
  wire \NLW_blk00000412_ACOUT<4>_UNCONNECTED ;
  wire \NLW_blk00000412_ACOUT<3>_UNCONNECTED ;
  wire \NLW_blk00000412_ACOUT<2>_UNCONNECTED ;
  wire \NLW_blk00000412_ACOUT<1>_UNCONNECTED ;
  wire \NLW_blk00000412_ACOUT<0>_UNCONNECTED ;
  wire \NLW_blk00000412_CARRYOUT<3>_UNCONNECTED ;
  wire \NLW_blk00000412_CARRYOUT<2>_UNCONNECTED ;
  wire \NLW_blk00000412_CARRYOUT<1>_UNCONNECTED ;
  wire \NLW_blk00000412_CARRYOUT<0>_UNCONNECTED ;
  wire \NLW_blk00000412_BCOUT<17>_UNCONNECTED ;
  wire \NLW_blk00000412_BCOUT<16>_UNCONNECTED ;
  wire \NLW_blk00000412_BCOUT<15>_UNCONNECTED ;
  wire \NLW_blk00000412_BCOUT<14>_UNCONNECTED ;
  wire \NLW_blk00000412_BCOUT<13>_UNCONNECTED ;
  wire \NLW_blk00000412_BCOUT<12>_UNCONNECTED ;
  wire \NLW_blk00000412_BCOUT<11>_UNCONNECTED ;
  wire \NLW_blk00000412_BCOUT<10>_UNCONNECTED ;
  wire \NLW_blk00000412_BCOUT<9>_UNCONNECTED ;
  wire \NLW_blk00000412_BCOUT<8>_UNCONNECTED ;
  wire \NLW_blk00000412_BCOUT<7>_UNCONNECTED ;
  wire \NLW_blk00000412_BCOUT<6>_UNCONNECTED ;
  wire \NLW_blk00000412_BCOUT<5>_UNCONNECTED ;
  wire \NLW_blk00000412_BCOUT<4>_UNCONNECTED ;
  wire \NLW_blk00000412_BCOUT<3>_UNCONNECTED ;
  wire \NLW_blk00000412_BCOUT<2>_UNCONNECTED ;
  wire \NLW_blk00000412_BCOUT<1>_UNCONNECTED ;
  wire \NLW_blk00000412_BCOUT<0>_UNCONNECTED ;
  wire \NLW_blk00000412_P<47>_UNCONNECTED ;
  wire \NLW_blk00000412_P<46>_UNCONNECTED ;
  wire \NLW_blk00000412_P<45>_UNCONNECTED ;
  wire \NLW_blk00000412_P<44>_UNCONNECTED ;
  wire \NLW_blk00000412_P<43>_UNCONNECTED ;
  wire \NLW_blk00000412_P<42>_UNCONNECTED ;
  wire \NLW_blk00000412_P<41>_UNCONNECTED ;
  wire \NLW_blk00000412_P<40>_UNCONNECTED ;
  wire \NLW_blk00000412_P<39>_UNCONNECTED ;
  wire \NLW_blk00000412_P<38>_UNCONNECTED ;
  wire \NLW_blk00000412_P<37>_UNCONNECTED ;
  wire \NLW_blk00000412_P<36>_UNCONNECTED ;
  wire \NLW_blk00000412_P<35>_UNCONNECTED ;
  wire \NLW_blk00000412_P<34>_UNCONNECTED ;
  wire \NLW_blk00000412_P<33>_UNCONNECTED ;
  wire \NLW_blk00000412_P<32>_UNCONNECTED ;
  wire \NLW_blk00000412_P<31>_UNCONNECTED ;
  wire \NLW_blk00000412_P<30>_UNCONNECTED ;
  wire \NLW_blk00000412_P<29>_UNCONNECTED ;
  wire \NLW_blk00000412_P<28>_UNCONNECTED ;
  wire \NLW_blk00000412_P<27>_UNCONNECTED ;
  wire \NLW_blk00000412_P<26>_UNCONNECTED ;
  wire \NLW_blk00000412_P<25>_UNCONNECTED ;
  wire \NLW_blk00000412_P<24>_UNCONNECTED ;
  wire \NLW_blk00000412_P<23>_UNCONNECTED ;
  wire \NLW_blk00000412_P<22>_UNCONNECTED ;
  wire \NLW_blk00000412_P<21>_UNCONNECTED ;
  wire \NLW_blk00000412_P<20>_UNCONNECTED ;
  wire \NLW_blk00000412_P<19>_UNCONNECTED ;
  wire \NLW_blk00000412_P<18>_UNCONNECTED ;
  wire \NLW_blk00000412_P<17>_UNCONNECTED ;
  wire \NLW_blk00000412_P<16>_UNCONNECTED ;
  wire \NLW_blk00000412_P<15>_UNCONNECTED ;
  wire \NLW_blk00000412_P<14>_UNCONNECTED ;
  wire \NLW_blk00000412_P<13>_UNCONNECTED ;
  wire \NLW_blk00000412_P<12>_UNCONNECTED ;
  wire \NLW_blk00000412_P<11>_UNCONNECTED ;
  wire \NLW_blk00000412_P<10>_UNCONNECTED ;
  wire \NLW_blk00000412_P<9>_UNCONNECTED ;
  wire \NLW_blk00000412_P<8>_UNCONNECTED ;
  wire \NLW_blk00000412_P<7>_UNCONNECTED ;
  wire \NLW_blk00000412_P<6>_UNCONNECTED ;
  wire \NLW_blk00000412_P<5>_UNCONNECTED ;
  wire \NLW_blk00000412_P<4>_UNCONNECTED ;
  wire \NLW_blk00000412_P<3>_UNCONNECTED ;
  wire \NLW_blk00000412_P<2>_UNCONNECTED ;
  wire \NLW_blk00000412_P<1>_UNCONNECTED ;
  wire \NLW_blk00000412_P<0>_UNCONNECTED ;
  wire NLW_blk00000413_PATTERNBDETECT_UNCONNECTED;
  wire NLW_blk00000413_MULTSIGNOUT_UNCONNECTED;
  wire NLW_blk00000413_CARRYCASCOUT_UNCONNECTED;
  wire NLW_blk00000413_UNDERFLOW_UNCONNECTED;
  wire NLW_blk00000413_PATTERNDETECT_UNCONNECTED;
  wire NLW_blk00000413_OVERFLOW_UNCONNECTED;
  wire \NLW_blk00000413_ACOUT<29>_UNCONNECTED ;
  wire \NLW_blk00000413_ACOUT<28>_UNCONNECTED ;
  wire \NLW_blk00000413_ACOUT<27>_UNCONNECTED ;
  wire \NLW_blk00000413_ACOUT<26>_UNCONNECTED ;
  wire \NLW_blk00000413_ACOUT<25>_UNCONNECTED ;
  wire \NLW_blk00000413_ACOUT<24>_UNCONNECTED ;
  wire \NLW_blk00000413_ACOUT<23>_UNCONNECTED ;
  wire \NLW_blk00000413_ACOUT<22>_UNCONNECTED ;
  wire \NLW_blk00000413_ACOUT<21>_UNCONNECTED ;
  wire \NLW_blk00000413_ACOUT<20>_UNCONNECTED ;
  wire \NLW_blk00000413_ACOUT<19>_UNCONNECTED ;
  wire \NLW_blk00000413_ACOUT<18>_UNCONNECTED ;
  wire \NLW_blk00000413_ACOUT<17>_UNCONNECTED ;
  wire \NLW_blk00000413_ACOUT<16>_UNCONNECTED ;
  wire \NLW_blk00000413_ACOUT<15>_UNCONNECTED ;
  wire \NLW_blk00000413_ACOUT<14>_UNCONNECTED ;
  wire \NLW_blk00000413_ACOUT<13>_UNCONNECTED ;
  wire \NLW_blk00000413_ACOUT<12>_UNCONNECTED ;
  wire \NLW_blk00000413_ACOUT<11>_UNCONNECTED ;
  wire \NLW_blk00000413_ACOUT<10>_UNCONNECTED ;
  wire \NLW_blk00000413_ACOUT<9>_UNCONNECTED ;
  wire \NLW_blk00000413_ACOUT<8>_UNCONNECTED ;
  wire \NLW_blk00000413_ACOUT<7>_UNCONNECTED ;
  wire \NLW_blk00000413_ACOUT<6>_UNCONNECTED ;
  wire \NLW_blk00000413_ACOUT<5>_UNCONNECTED ;
  wire \NLW_blk00000413_ACOUT<4>_UNCONNECTED ;
  wire \NLW_blk00000413_ACOUT<3>_UNCONNECTED ;
  wire \NLW_blk00000413_ACOUT<2>_UNCONNECTED ;
  wire \NLW_blk00000413_ACOUT<1>_UNCONNECTED ;
  wire \NLW_blk00000413_ACOUT<0>_UNCONNECTED ;
  wire \NLW_blk00000413_CARRYOUT<3>_UNCONNECTED ;
  wire \NLW_blk00000413_CARRYOUT<2>_UNCONNECTED ;
  wire \NLW_blk00000413_CARRYOUT<1>_UNCONNECTED ;
  wire \NLW_blk00000413_CARRYOUT<0>_UNCONNECTED ;
  wire \NLW_blk00000413_BCOUT<17>_UNCONNECTED ;
  wire \NLW_blk00000413_BCOUT<16>_UNCONNECTED ;
  wire \NLW_blk00000413_BCOUT<15>_UNCONNECTED ;
  wire \NLW_blk00000413_BCOUT<14>_UNCONNECTED ;
  wire \NLW_blk00000413_BCOUT<13>_UNCONNECTED ;
  wire \NLW_blk00000413_BCOUT<12>_UNCONNECTED ;
  wire \NLW_blk00000413_BCOUT<11>_UNCONNECTED ;
  wire \NLW_blk00000413_BCOUT<10>_UNCONNECTED ;
  wire \NLW_blk00000413_BCOUT<9>_UNCONNECTED ;
  wire \NLW_blk00000413_BCOUT<8>_UNCONNECTED ;
  wire \NLW_blk00000413_BCOUT<7>_UNCONNECTED ;
  wire \NLW_blk00000413_BCOUT<6>_UNCONNECTED ;
  wire \NLW_blk00000413_BCOUT<5>_UNCONNECTED ;
  wire \NLW_blk00000413_BCOUT<4>_UNCONNECTED ;
  wire \NLW_blk00000413_BCOUT<3>_UNCONNECTED ;
  wire \NLW_blk00000413_BCOUT<2>_UNCONNECTED ;
  wire \NLW_blk00000413_BCOUT<1>_UNCONNECTED ;
  wire \NLW_blk00000413_BCOUT<0>_UNCONNECTED ;
  wire \NLW_blk00000413_P<47>_UNCONNECTED ;
  wire \NLW_blk00000413_P<46>_UNCONNECTED ;
  wire \NLW_blk00000413_P<45>_UNCONNECTED ;
  wire \NLW_blk00000413_P<44>_UNCONNECTED ;
  wire \NLW_blk00000413_P<43>_UNCONNECTED ;
  wire \NLW_blk00000413_P<42>_UNCONNECTED ;
  wire \NLW_blk00000413_P<41>_UNCONNECTED ;
  wire \NLW_blk00000413_P<40>_UNCONNECTED ;
  wire \NLW_blk00000413_P<39>_UNCONNECTED ;
  wire \NLW_blk00000413_P<38>_UNCONNECTED ;
  wire \NLW_blk00000413_P<37>_UNCONNECTED ;
  wire \NLW_blk00000413_P<36>_UNCONNECTED ;
  wire \NLW_blk00000413_P<35>_UNCONNECTED ;
  wire \NLW_blk00000413_P<34>_UNCONNECTED ;
  wire \NLW_blk00000413_P<33>_UNCONNECTED ;
  wire \NLW_blk00000413_P<32>_UNCONNECTED ;
  wire \NLW_blk00000413_P<31>_UNCONNECTED ;
  wire \NLW_blk00000413_P<30>_UNCONNECTED ;
  wire \NLW_blk00000413_P<29>_UNCONNECTED ;
  wire \NLW_blk00000413_P<28>_UNCONNECTED ;
  wire \NLW_blk00000413_P<27>_UNCONNECTED ;
  wire \NLW_blk00000413_P<26>_UNCONNECTED ;
  wire \NLW_blk00000413_P<25>_UNCONNECTED ;
  wire \NLW_blk00000413_P<24>_UNCONNECTED ;
  wire \NLW_blk00000413_P<23>_UNCONNECTED ;
  wire \NLW_blk00000413_P<22>_UNCONNECTED ;
  wire \NLW_blk00000413_P<21>_UNCONNECTED ;
  wire \NLW_blk00000413_P<20>_UNCONNECTED ;
  wire \NLW_blk00000413_P<19>_UNCONNECTED ;
  wire \NLW_blk00000413_P<18>_UNCONNECTED ;
  wire \NLW_blk00000413_P<17>_UNCONNECTED ;
  wire \NLW_blk00000413_P<16>_UNCONNECTED ;
  wire \NLW_blk00000413_P<15>_UNCONNECTED ;
  wire \NLW_blk00000413_P<14>_UNCONNECTED ;
  wire \NLW_blk00000413_P<13>_UNCONNECTED ;
  wire \NLW_blk00000413_P<12>_UNCONNECTED ;
  wire \NLW_blk00000413_P<11>_UNCONNECTED ;
  wire \NLW_blk00000413_P<10>_UNCONNECTED ;
  wire \NLW_blk00000413_P<9>_UNCONNECTED ;
  wire \NLW_blk00000413_P<8>_UNCONNECTED ;
  wire \NLW_blk00000413_P<7>_UNCONNECTED ;
  wire \NLW_blk00000413_P<6>_UNCONNECTED ;
  wire \NLW_blk00000413_P<5>_UNCONNECTED ;
  wire \NLW_blk00000413_P<4>_UNCONNECTED ;
  wire \NLW_blk00000413_P<3>_UNCONNECTED ;
  wire \NLW_blk00000413_P<2>_UNCONNECTED ;
  wire \NLW_blk00000413_P<1>_UNCONNECTED ;
  wire \NLW_blk00000413_P<0>_UNCONNECTED ;
  wire NLW_blk00000414_PATTERNBDETECT_UNCONNECTED;
  wire NLW_blk00000414_MULTSIGNOUT_UNCONNECTED;
  wire NLW_blk00000414_CARRYCASCOUT_UNCONNECTED;
  wire NLW_blk00000414_UNDERFLOW_UNCONNECTED;
  wire NLW_blk00000414_OVERFLOW_UNCONNECTED;
  wire \NLW_blk00000414_ACOUT<29>_UNCONNECTED ;
  wire \NLW_blk00000414_ACOUT<28>_UNCONNECTED ;
  wire \NLW_blk00000414_ACOUT<27>_UNCONNECTED ;
  wire \NLW_blk00000414_ACOUT<26>_UNCONNECTED ;
  wire \NLW_blk00000414_ACOUT<25>_UNCONNECTED ;
  wire \NLW_blk00000414_ACOUT<24>_UNCONNECTED ;
  wire \NLW_blk00000414_ACOUT<23>_UNCONNECTED ;
  wire \NLW_blk00000414_ACOUT<22>_UNCONNECTED ;
  wire \NLW_blk00000414_ACOUT<21>_UNCONNECTED ;
  wire \NLW_blk00000414_ACOUT<20>_UNCONNECTED ;
  wire \NLW_blk00000414_ACOUT<19>_UNCONNECTED ;
  wire \NLW_blk00000414_ACOUT<18>_UNCONNECTED ;
  wire \NLW_blk00000414_ACOUT<17>_UNCONNECTED ;
  wire \NLW_blk00000414_ACOUT<16>_UNCONNECTED ;
  wire \NLW_blk00000414_ACOUT<15>_UNCONNECTED ;
  wire \NLW_blk00000414_ACOUT<14>_UNCONNECTED ;
  wire \NLW_blk00000414_ACOUT<13>_UNCONNECTED ;
  wire \NLW_blk00000414_ACOUT<12>_UNCONNECTED ;
  wire \NLW_blk00000414_ACOUT<11>_UNCONNECTED ;
  wire \NLW_blk00000414_ACOUT<10>_UNCONNECTED ;
  wire \NLW_blk00000414_ACOUT<9>_UNCONNECTED ;
  wire \NLW_blk00000414_ACOUT<8>_UNCONNECTED ;
  wire \NLW_blk00000414_ACOUT<7>_UNCONNECTED ;
  wire \NLW_blk00000414_ACOUT<6>_UNCONNECTED ;
  wire \NLW_blk00000414_ACOUT<5>_UNCONNECTED ;
  wire \NLW_blk00000414_ACOUT<4>_UNCONNECTED ;
  wire \NLW_blk00000414_ACOUT<3>_UNCONNECTED ;
  wire \NLW_blk00000414_ACOUT<2>_UNCONNECTED ;
  wire \NLW_blk00000414_ACOUT<1>_UNCONNECTED ;
  wire \NLW_blk00000414_ACOUT<0>_UNCONNECTED ;
  wire \NLW_blk00000414_CARRYOUT<3>_UNCONNECTED ;
  wire \NLW_blk00000414_CARRYOUT<2>_UNCONNECTED ;
  wire \NLW_blk00000414_CARRYOUT<1>_UNCONNECTED ;
  wire \NLW_blk00000414_CARRYOUT<0>_UNCONNECTED ;
  wire \NLW_blk00000414_P<47>_UNCONNECTED ;
  wire \NLW_blk00000414_P<46>_UNCONNECTED ;
  wire \NLW_blk00000414_P<45>_UNCONNECTED ;
  wire \NLW_blk00000414_P<44>_UNCONNECTED ;
  wire \NLW_blk00000414_P<43>_UNCONNECTED ;
  wire \NLW_blk00000414_P<42>_UNCONNECTED ;
  wire \NLW_blk00000414_P<41>_UNCONNECTED ;
  wire \NLW_blk00000414_P<40>_UNCONNECTED ;
  wire \NLW_blk00000414_P<39>_UNCONNECTED ;
  wire \NLW_blk00000414_P<38>_UNCONNECTED ;
  wire \NLW_blk00000414_P<37>_UNCONNECTED ;
  wire \NLW_blk00000414_P<36>_UNCONNECTED ;
  wire \NLW_blk00000414_P<35>_UNCONNECTED ;
  wire \NLW_blk00000414_P<34>_UNCONNECTED ;
  wire \NLW_blk00000414_P<33>_UNCONNECTED ;
  wire \NLW_blk00000414_P<32>_UNCONNECTED ;
  wire \NLW_blk00000414_P<31>_UNCONNECTED ;
  wire \NLW_blk00000414_P<30>_UNCONNECTED ;
  wire \NLW_blk00000414_P<29>_UNCONNECTED ;
  wire \NLW_blk00000414_P<28>_UNCONNECTED ;
  wire \NLW_blk00000414_P<27>_UNCONNECTED ;
  wire \NLW_blk00000414_P<26>_UNCONNECTED ;
  wire \NLW_blk00000414_P<25>_UNCONNECTED ;
  wire \NLW_blk00000414_P<24>_UNCONNECTED ;
  wire \NLW_blk00000414_P<23>_UNCONNECTED ;
  wire \NLW_blk00000414_P<22>_UNCONNECTED ;
  wire \NLW_blk00000414_P<21>_UNCONNECTED ;
  wire \NLW_blk00000414_P<20>_UNCONNECTED ;
  wire \NLW_blk00000414_P<19>_UNCONNECTED ;
  wire \NLW_blk00000414_P<18>_UNCONNECTED ;
  wire \NLW_blk00000414_P<17>_UNCONNECTED ;
  wire \NLW_blk00000414_P<16>_UNCONNECTED ;
  wire \NLW_blk00000414_P<15>_UNCONNECTED ;
  wire \NLW_blk00000414_P<14>_UNCONNECTED ;
  wire \NLW_blk00000414_P<13>_UNCONNECTED ;
  wire \NLW_blk00000414_P<12>_UNCONNECTED ;
  wire \NLW_blk00000414_P<11>_UNCONNECTED ;
  wire \NLW_blk00000414_P<10>_UNCONNECTED ;
  wire \NLW_blk00000414_P<9>_UNCONNECTED ;
  wire \NLW_blk00000414_P<8>_UNCONNECTED ;
  wire \NLW_blk00000414_P<7>_UNCONNECTED ;
  wire \NLW_blk00000414_P<6>_UNCONNECTED ;
  wire \NLW_blk00000414_P<5>_UNCONNECTED ;
  wire \NLW_blk00000414_P<4>_UNCONNECTED ;
  wire \NLW_blk00000414_P<3>_UNCONNECTED ;
  wire \NLW_blk00000414_P<2>_UNCONNECTED ;
  wire \NLW_blk00000414_P<1>_UNCONNECTED ;
  wire \NLW_blk00000414_P<0>_UNCONNECTED ;
  wire NLW_blk00000415_PATTERNBDETECT_UNCONNECTED;
  wire NLW_blk00000415_MULTSIGNOUT_UNCONNECTED;
  wire NLW_blk00000415_CARRYCASCOUT_UNCONNECTED;
  wire NLW_blk00000415_UNDERFLOW_UNCONNECTED;
  wire NLW_blk00000415_PATTERNDETECT_UNCONNECTED;
  wire NLW_blk00000415_OVERFLOW_UNCONNECTED;
  wire \NLW_blk00000415_ACOUT<29>_UNCONNECTED ;
  wire \NLW_blk00000415_ACOUT<28>_UNCONNECTED ;
  wire \NLW_blk00000415_ACOUT<27>_UNCONNECTED ;
  wire \NLW_blk00000415_ACOUT<26>_UNCONNECTED ;
  wire \NLW_blk00000415_ACOUT<25>_UNCONNECTED ;
  wire \NLW_blk00000415_ACOUT<24>_UNCONNECTED ;
  wire \NLW_blk00000415_ACOUT<23>_UNCONNECTED ;
  wire \NLW_blk00000415_ACOUT<22>_UNCONNECTED ;
  wire \NLW_blk00000415_ACOUT<21>_UNCONNECTED ;
  wire \NLW_blk00000415_ACOUT<20>_UNCONNECTED ;
  wire \NLW_blk00000415_ACOUT<19>_UNCONNECTED ;
  wire \NLW_blk00000415_ACOUT<18>_UNCONNECTED ;
  wire \NLW_blk00000415_ACOUT<17>_UNCONNECTED ;
  wire \NLW_blk00000415_ACOUT<16>_UNCONNECTED ;
  wire \NLW_blk00000415_ACOUT<15>_UNCONNECTED ;
  wire \NLW_blk00000415_ACOUT<14>_UNCONNECTED ;
  wire \NLW_blk00000415_ACOUT<13>_UNCONNECTED ;
  wire \NLW_blk00000415_ACOUT<12>_UNCONNECTED ;
  wire \NLW_blk00000415_ACOUT<11>_UNCONNECTED ;
  wire \NLW_blk00000415_ACOUT<10>_UNCONNECTED ;
  wire \NLW_blk00000415_ACOUT<9>_UNCONNECTED ;
  wire \NLW_blk00000415_ACOUT<8>_UNCONNECTED ;
  wire \NLW_blk00000415_ACOUT<7>_UNCONNECTED ;
  wire \NLW_blk00000415_ACOUT<6>_UNCONNECTED ;
  wire \NLW_blk00000415_ACOUT<5>_UNCONNECTED ;
  wire \NLW_blk00000415_ACOUT<4>_UNCONNECTED ;
  wire \NLW_blk00000415_ACOUT<3>_UNCONNECTED ;
  wire \NLW_blk00000415_ACOUT<2>_UNCONNECTED ;
  wire \NLW_blk00000415_ACOUT<1>_UNCONNECTED ;
  wire \NLW_blk00000415_ACOUT<0>_UNCONNECTED ;
  wire \NLW_blk00000415_CARRYOUT<3>_UNCONNECTED ;
  wire \NLW_blk00000415_CARRYOUT<2>_UNCONNECTED ;
  wire \NLW_blk00000415_CARRYOUT<1>_UNCONNECTED ;
  wire \NLW_blk00000415_CARRYOUT<0>_UNCONNECTED ;
  wire \NLW_blk00000415_BCOUT<17>_UNCONNECTED ;
  wire \NLW_blk00000415_BCOUT<16>_UNCONNECTED ;
  wire \NLW_blk00000415_BCOUT<15>_UNCONNECTED ;
  wire \NLW_blk00000415_BCOUT<14>_UNCONNECTED ;
  wire \NLW_blk00000415_BCOUT<13>_UNCONNECTED ;
  wire \NLW_blk00000415_BCOUT<12>_UNCONNECTED ;
  wire \NLW_blk00000415_BCOUT<11>_UNCONNECTED ;
  wire \NLW_blk00000415_BCOUT<10>_UNCONNECTED ;
  wire \NLW_blk00000415_BCOUT<9>_UNCONNECTED ;
  wire \NLW_blk00000415_BCOUT<8>_UNCONNECTED ;
  wire \NLW_blk00000415_BCOUT<7>_UNCONNECTED ;
  wire \NLW_blk00000415_BCOUT<6>_UNCONNECTED ;
  wire \NLW_blk00000415_BCOUT<5>_UNCONNECTED ;
  wire \NLW_blk00000415_BCOUT<4>_UNCONNECTED ;
  wire \NLW_blk00000415_BCOUT<3>_UNCONNECTED ;
  wire \NLW_blk00000415_BCOUT<2>_UNCONNECTED ;
  wire \NLW_blk00000415_BCOUT<1>_UNCONNECTED ;
  wire \NLW_blk00000415_BCOUT<0>_UNCONNECTED ;
  wire \NLW_blk00000415_P<47>_UNCONNECTED ;
  wire \NLW_blk00000415_P<46>_UNCONNECTED ;
  wire \NLW_blk00000415_P<45>_UNCONNECTED ;
  wire \NLW_blk00000415_P<44>_UNCONNECTED ;
  wire \NLW_blk00000415_P<43>_UNCONNECTED ;
  wire \NLW_blk00000415_P<42>_UNCONNECTED ;
  wire \NLW_blk00000415_P<41>_UNCONNECTED ;
  wire \NLW_blk00000415_P<40>_UNCONNECTED ;
  wire \NLW_blk00000415_P<39>_UNCONNECTED ;
  wire \NLW_blk00000415_P<38>_UNCONNECTED ;
  wire \NLW_blk00000415_P<37>_UNCONNECTED ;
  wire \NLW_blk00000415_P<36>_UNCONNECTED ;
  wire \NLW_blk00000415_P<35>_UNCONNECTED ;
  wire \NLW_blk00000415_P<34>_UNCONNECTED ;
  wire \NLW_blk00000415_P<33>_UNCONNECTED ;
  wire \NLW_blk00000415_P<32>_UNCONNECTED ;
  wire \NLW_blk00000415_P<31>_UNCONNECTED ;
  wire \NLW_blk00000415_P<30>_UNCONNECTED ;
  wire \NLW_blk00000415_P<29>_UNCONNECTED ;
  wire \NLW_blk00000415_P<28>_UNCONNECTED ;
  wire \NLW_blk00000415_P<27>_UNCONNECTED ;
  wire \NLW_blk00000415_P<26>_UNCONNECTED ;
  wire \NLW_blk00000415_P<25>_UNCONNECTED ;
  wire \NLW_blk00000415_P<24>_UNCONNECTED ;
  wire \NLW_blk00000415_P<23>_UNCONNECTED ;
  wire \NLW_blk00000415_P<22>_UNCONNECTED ;
  wire \NLW_blk00000415_P<21>_UNCONNECTED ;
  wire \NLW_blk00000415_P<20>_UNCONNECTED ;
  wire \NLW_blk00000415_P<19>_UNCONNECTED ;
  wire \NLW_blk00000415_P<18>_UNCONNECTED ;
  wire \NLW_blk00000415_P<17>_UNCONNECTED ;
  wire \NLW_blk00000415_P<16>_UNCONNECTED ;
  wire \NLW_blk00000415_P<15>_UNCONNECTED ;
  wire \NLW_blk00000415_P<14>_UNCONNECTED ;
  wire \NLW_blk00000415_P<13>_UNCONNECTED ;
  wire \NLW_blk00000415_P<12>_UNCONNECTED ;
  wire \NLW_blk00000415_P<11>_UNCONNECTED ;
  wire \NLW_blk00000415_P<10>_UNCONNECTED ;
  wire \NLW_blk00000415_P<9>_UNCONNECTED ;
  wire \NLW_blk00000415_P<8>_UNCONNECTED ;
  wire \NLW_blk00000415_P<7>_UNCONNECTED ;
  wire \NLW_blk00000415_P<6>_UNCONNECTED ;
  wire \NLW_blk00000415_P<5>_UNCONNECTED ;
  wire \NLW_blk00000415_P<4>_UNCONNECTED ;
  wire \NLW_blk00000415_P<3>_UNCONNECTED ;
  wire \NLW_blk00000415_P<2>_UNCONNECTED ;
  wire \NLW_blk00000415_P<1>_UNCONNECTED ;
  wire \NLW_blk00000415_P<0>_UNCONNECTED ;
  wire NLW_blk00000416_PATTERNBDETECT_UNCONNECTED;
  wire NLW_blk00000416_MULTSIGNOUT_UNCONNECTED;
  wire NLW_blk00000416_CARRYCASCOUT_UNCONNECTED;
  wire NLW_blk00000416_UNDERFLOW_UNCONNECTED;
  wire NLW_blk00000416_OVERFLOW_UNCONNECTED;
  wire \NLW_blk00000416_ACOUT<29>_UNCONNECTED ;
  wire \NLW_blk00000416_ACOUT<28>_UNCONNECTED ;
  wire \NLW_blk00000416_ACOUT<27>_UNCONNECTED ;
  wire \NLW_blk00000416_ACOUT<26>_UNCONNECTED ;
  wire \NLW_blk00000416_ACOUT<25>_UNCONNECTED ;
  wire \NLW_blk00000416_ACOUT<24>_UNCONNECTED ;
  wire \NLW_blk00000416_ACOUT<23>_UNCONNECTED ;
  wire \NLW_blk00000416_ACOUT<22>_UNCONNECTED ;
  wire \NLW_blk00000416_ACOUT<21>_UNCONNECTED ;
  wire \NLW_blk00000416_ACOUT<20>_UNCONNECTED ;
  wire \NLW_blk00000416_ACOUT<19>_UNCONNECTED ;
  wire \NLW_blk00000416_ACOUT<18>_UNCONNECTED ;
  wire \NLW_blk00000416_ACOUT<17>_UNCONNECTED ;
  wire \NLW_blk00000416_ACOUT<16>_UNCONNECTED ;
  wire \NLW_blk00000416_ACOUT<15>_UNCONNECTED ;
  wire \NLW_blk00000416_ACOUT<14>_UNCONNECTED ;
  wire \NLW_blk00000416_ACOUT<13>_UNCONNECTED ;
  wire \NLW_blk00000416_ACOUT<12>_UNCONNECTED ;
  wire \NLW_blk00000416_ACOUT<11>_UNCONNECTED ;
  wire \NLW_blk00000416_ACOUT<10>_UNCONNECTED ;
  wire \NLW_blk00000416_ACOUT<9>_UNCONNECTED ;
  wire \NLW_blk00000416_ACOUT<8>_UNCONNECTED ;
  wire \NLW_blk00000416_ACOUT<7>_UNCONNECTED ;
  wire \NLW_blk00000416_ACOUT<6>_UNCONNECTED ;
  wire \NLW_blk00000416_ACOUT<5>_UNCONNECTED ;
  wire \NLW_blk00000416_ACOUT<4>_UNCONNECTED ;
  wire \NLW_blk00000416_ACOUT<3>_UNCONNECTED ;
  wire \NLW_blk00000416_ACOUT<2>_UNCONNECTED ;
  wire \NLW_blk00000416_ACOUT<1>_UNCONNECTED ;
  wire \NLW_blk00000416_ACOUT<0>_UNCONNECTED ;
  wire \NLW_blk00000416_CARRYOUT<3>_UNCONNECTED ;
  wire \NLW_blk00000416_CARRYOUT<2>_UNCONNECTED ;
  wire \NLW_blk00000416_CARRYOUT<1>_UNCONNECTED ;
  wire \NLW_blk00000416_CARRYOUT<0>_UNCONNECTED ;
  wire \NLW_blk00000416_P<47>_UNCONNECTED ;
  wire \NLW_blk00000416_P<46>_UNCONNECTED ;
  wire \NLW_blk00000416_P<45>_UNCONNECTED ;
  wire \NLW_blk00000416_P<44>_UNCONNECTED ;
  wire \NLW_blk00000416_P<43>_UNCONNECTED ;
  wire \NLW_blk00000416_P<42>_UNCONNECTED ;
  wire \NLW_blk00000416_P<41>_UNCONNECTED ;
  wire \NLW_blk00000416_P<40>_UNCONNECTED ;
  wire \NLW_blk00000416_P<39>_UNCONNECTED ;
  wire \NLW_blk00000416_P<38>_UNCONNECTED ;
  wire \NLW_blk00000416_P<37>_UNCONNECTED ;
  wire \NLW_blk00000416_P<36>_UNCONNECTED ;
  wire \NLW_blk00000416_P<35>_UNCONNECTED ;
  wire \NLW_blk00000416_P<34>_UNCONNECTED ;
  wire \NLW_blk00000416_P<33>_UNCONNECTED ;
  wire \NLW_blk00000416_P<32>_UNCONNECTED ;
  wire \NLW_blk00000416_P<31>_UNCONNECTED ;
  wire \NLW_blk00000416_P<30>_UNCONNECTED ;
  wire \NLW_blk00000416_P<29>_UNCONNECTED ;
  wire \NLW_blk00000416_P<28>_UNCONNECTED ;
  wire \NLW_blk00000416_P<27>_UNCONNECTED ;
  wire \NLW_blk00000416_P<26>_UNCONNECTED ;
  wire \NLW_blk00000416_P<25>_UNCONNECTED ;
  wire \NLW_blk00000416_P<24>_UNCONNECTED ;
  wire \NLW_blk00000416_P<23>_UNCONNECTED ;
  wire \NLW_blk00000416_P<22>_UNCONNECTED ;
  wire \NLW_blk00000416_P<21>_UNCONNECTED ;
  wire \NLW_blk00000416_P<20>_UNCONNECTED ;
  wire \NLW_blk00000416_P<19>_UNCONNECTED ;
  wire \NLW_blk00000416_P<18>_UNCONNECTED ;
  wire \NLW_blk00000416_P<17>_UNCONNECTED ;
  wire \NLW_blk00000416_P<16>_UNCONNECTED ;
  wire \NLW_blk00000416_P<15>_UNCONNECTED ;
  wire \NLW_blk00000416_P<14>_UNCONNECTED ;
  wire \NLW_blk00000416_P<13>_UNCONNECTED ;
  wire \NLW_blk00000416_P<12>_UNCONNECTED ;
  wire \NLW_blk00000416_P<11>_UNCONNECTED ;
  wire \NLW_blk00000416_P<10>_UNCONNECTED ;
  wire \NLW_blk00000416_P<9>_UNCONNECTED ;
  wire \NLW_blk00000416_P<8>_UNCONNECTED ;
  wire \NLW_blk00000416_P<7>_UNCONNECTED ;
  wire \NLW_blk00000416_P<6>_UNCONNECTED ;
  wire \NLW_blk00000416_P<5>_UNCONNECTED ;
  wire \NLW_blk00000416_P<4>_UNCONNECTED ;
  wire \NLW_blk00000416_P<3>_UNCONNECTED ;
  wire \NLW_blk00000416_P<2>_UNCONNECTED ;
  wire \NLW_blk00000416_P<1>_UNCONNECTED ;
  wire \NLW_blk00000416_P<0>_UNCONNECTED ;
  wire [10 : 0] \NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/exp_op ;
  wire [51 : 0] \NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op ;
  assign
    result[63] = \U0/op_inst/FLT_PT_OP/MULT.OP/OP/sign_op ,
    result[62] = \NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/exp_op [10],
    result[61] = \NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/exp_op [9],
    result[60] = \NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/exp_op [8],
    result[59] = \NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/exp_op [7],
    result[58] = \NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/exp_op [6],
    result[57] = \NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/exp_op [5],
    result[56] = \NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/exp_op [4],
    result[55] = \NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/exp_op [3],
    result[54] = \NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/exp_op [2],
    result[53] = \NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/exp_op [1],
    result[52] = \NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/exp_op [0],
    result[51] = \NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [51],
    result[50] = \NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [50],
    result[49] = \NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [49],
    result[48] = \NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [48],
    result[47] = \NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [47],
    result[46] = \NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [46],
    result[45] = \NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [45],
    result[44] = \NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [44],
    result[43] = \NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [43],
    result[42] = \NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [42],
    result[41] = \NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [41],
    result[40] = \NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [40],
    result[39] = \NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [39],
    result[38] = \NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [38],
    result[37] = \NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [37],
    result[36] = \NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [36],
    result[35] = \NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [35],
    result[34] = \NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [34],
    result[33] = \NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [33],
    result[32] = \NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [32],
    result[31] = \NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [31],
    result[30] = \NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [30],
    result[29] = \NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [29],
    result[28] = \NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [28],
    result[27] = \NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [27],
    result[26] = \NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [26],
    result[25] = \NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [25],
    result[24] = \NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [24],
    result[23] = \NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [23],
    result[22] = \NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [22],
    result[21] = \NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [21],
    result[20] = \NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [20],
    result[19] = \NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [19],
    result[18] = \NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [18],
    result[17] = \NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [17],
    result[16] = \NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [16],
    result[15] = \NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [15],
    result[14] = \NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [14],
    result[13] = \NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [13],
    result[12] = \NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [12],
    result[11] = \NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [11],
    result[10] = \NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [10],
    result[9] = \NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [9],
    result[8] = \NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [8],
    result[7] = \NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [7],
    result[6] = \NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [6],
    result[5] = \NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [5],
    result[4] = \NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [4],
    result[3] = \NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [3],
    result[2] = \NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [2],
    result[1] = \NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [1],
    result[0] = \NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [0],
    rdy = \NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/HND_SHK/RDY ;
  VCC   blk00000001 (
    .P(sig00000001)
  );
  GND   blk00000002 (
    .G(sig00000461)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000003 (
    .C(clk),
    .CE(ce),
    .D(sig00000091),
    .Q(sig0000007e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000004 (
    .C(clk),
    .CE(ce),
    .D(sig00000092),
    .Q(sig0000007b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000005 (
    .C(clk),
    .CE(ce),
    .D(sig0000009f),
    .Q(sig0000007f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000006 (
    .C(clk),
    .CE(ce),
    .D(sig0000008f),
    .Q(sig000000a2)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000007 (
    .C(clk),
    .CE(ce),
    .D(sig00000090),
    .Q(sig0000009a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000008 (
    .C(clk),
    .CE(ce),
    .D(sig00000083),
    .Q(sig000000a3)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000009 (
    .C(clk),
    .CE(ce),
    .D(sig00000082),
    .Q(sig000000a4)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000000a (
    .C(clk),
    .CE(ce),
    .D(sig00000081),
    .Q(sig000000a6)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000000b (
    .C(clk),
    .CE(ce),
    .D(sig00000080),
    .Q(sig000000a7)
  );
  XORCY   blk0000000c (
    .CI(sig000000b7),
    .LI(sig00000461),
    .O(sig000000b5)
  );
  XORCY   blk0000000d (
    .CI(sig000000b9),
    .LI(sig0000008e),
    .O(sig000000b6)
  );
  MUXCY   blk0000000e (
    .CI(sig000000b9),
    .DI(b[62]),
    .S(sig0000008e),
    .O(sig000000b7)
  );
  XORCY   blk0000000f (
    .CI(sig000000bb),
    .LI(sig0000008d),
    .O(sig000000b8)
  );
  MUXCY   blk00000010 (
    .CI(sig000000bb),
    .DI(b[61]),
    .S(sig0000008d),
    .O(sig000000b9)
  );
  XORCY   blk00000011 (
    .CI(sig000000bd),
    .LI(sig0000008c),
    .O(sig000000ba)
  );
  MUXCY   blk00000012 (
    .CI(sig000000bd),
    .DI(b[60]),
    .S(sig0000008c),
    .O(sig000000bb)
  );
  XORCY   blk00000013 (
    .CI(sig000000bf),
    .LI(sig0000008b),
    .O(sig000000bc)
  );
  MUXCY   blk00000014 (
    .CI(sig000000bf),
    .DI(b[59]),
    .S(sig0000008b),
    .O(sig000000bd)
  );
  XORCY   blk00000015 (
    .CI(sig000000c1),
    .LI(sig0000008a),
    .O(sig000000be)
  );
  MUXCY   blk00000016 (
    .CI(sig000000c1),
    .DI(b[58]),
    .S(sig0000008a),
    .O(sig000000bf)
  );
  XORCY   blk00000017 (
    .CI(sig000000c3),
    .LI(sig00000089),
    .O(sig000000c0)
  );
  MUXCY   blk00000018 (
    .CI(sig000000c3),
    .DI(b[57]),
    .S(sig00000089),
    .O(sig000000c1)
  );
  XORCY   blk00000019 (
    .CI(sig000000c5),
    .LI(sig00000088),
    .O(sig000000c2)
  );
  MUXCY   blk0000001a (
    .CI(sig000000c5),
    .DI(b[56]),
    .S(sig00000088),
    .O(sig000000c3)
  );
  XORCY   blk0000001b (
    .CI(sig000000c7),
    .LI(sig00000087),
    .O(sig000000c4)
  );
  MUXCY   blk0000001c (
    .CI(sig000000c7),
    .DI(b[55]),
    .S(sig00000087),
    .O(sig000000c5)
  );
  XORCY   blk0000001d (
    .CI(sig000000c9),
    .LI(sig00000086),
    .O(sig000000c6)
  );
  MUXCY   blk0000001e (
    .CI(sig000000c9),
    .DI(b[54]),
    .S(sig00000086),
    .O(sig000000c7)
  );
  XORCY   blk0000001f (
    .CI(sig000000cb),
    .LI(sig00000085),
    .O(sig000000c8)
  );
  MUXCY   blk00000020 (
    .CI(sig000000cb),
    .DI(b[53]),
    .S(sig00000085),
    .O(sig000000c9)
  );
  XORCY   blk00000021 (
    .CI(sig00000001),
    .LI(sig00000084),
    .O(sig000000ca)
  );
  MUXCY   blk00000022 (
    .CI(sig00000001),
    .DI(b[52]),
    .S(sig00000084),
    .O(sig000000cb)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000023 (
    .C(clk),
    .CE(ce),
    .D(sig000000b5),
    .Q(sig000000a9)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000024 (
    .C(clk),
    .CE(ce),
    .D(sig000000b6),
    .Q(sig000000b4)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000025 (
    .C(clk),
    .CE(ce),
    .D(sig000000b8),
    .Q(sig000000b3)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000026 (
    .C(clk),
    .CE(ce),
    .D(sig000000ba),
    .Q(sig000000b2)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000027 (
    .C(clk),
    .CE(ce),
    .D(sig000000bc),
    .Q(sig000000b1)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000028 (
    .C(clk),
    .CE(ce),
    .D(sig000000be),
    .Q(sig000000b0)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000029 (
    .C(clk),
    .CE(ce),
    .D(sig000000c0),
    .Q(sig000000af)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000002a (
    .C(clk),
    .CE(ce),
    .D(sig000000c2),
    .Q(sig000000ae)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000002b (
    .C(clk),
    .CE(ce),
    .D(sig000000c4),
    .Q(sig000000ad)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000002c (
    .C(clk),
    .CE(ce),
    .D(sig000000c6),
    .Q(sig000000ac)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000002d (
    .C(clk),
    .CE(ce),
    .D(sig000000c8),
    .Q(sig000000ab)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000002e (
    .C(clk),
    .CE(ce),
    .D(sig000000ca),
    .Q(sig000000aa)
  );
  MUXCY   blk0000002f (
    .CI(sig000000df),
    .DI(sig00000461),
    .S(sig000000dd),
    .O(sig000000de)
  );
  MUXCY   blk00000030 (
    .CI(sig000000e0),
    .DI(sig00000461),
    .S(sig000000d5),
    .O(sig000000df)
  );
  MUXCY   blk00000031 (
    .CI(sig000000e1),
    .DI(sig00000461),
    .S(sig000000d6),
    .O(sig000000e0)
  );
  MUXCY   blk00000032 (
    .CI(sig000000e2),
    .DI(sig00000461),
    .S(sig000000d7),
    .O(sig000000e1)
  );
  MUXCY   blk00000033 (
    .CI(sig000000e3),
    .DI(sig00000461),
    .S(sig000000d8),
    .O(sig000000e2)
  );
  MUXCY   blk00000034 (
    .CI(sig000000e4),
    .DI(sig00000461),
    .S(sig000000d9),
    .O(sig000000e3)
  );
  MUXCY   blk00000035 (
    .CI(sig000000e5),
    .DI(sig00000461),
    .S(sig000000da),
    .O(sig000000e4)
  );
  MUXCY   blk00000036 (
    .CI(sig000000e6),
    .DI(sig00000461),
    .S(sig000000db),
    .O(sig000000e5)
  );
  MUXCY   blk00000037 (
    .CI(sig00000001),
    .DI(sig00000461),
    .S(sig000000dc),
    .O(sig000000e6)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000038 (
    .C(clk),
    .CE(ce),
    .D(sig000000de),
    .Q(sig000000a5)
  );
  MUXCY   blk00000039 (
    .CI(sig000000e8),
    .DI(sig00000461),
    .S(sig000000d4),
    .O(sig000000e7)
  );
  MUXCY   blk0000003a (
    .CI(sig000000e9),
    .DI(sig00000461),
    .S(sig000000cc),
    .O(sig000000e8)
  );
  MUXCY   blk0000003b (
    .CI(sig000000ea),
    .DI(sig00000461),
    .S(sig000000cd),
    .O(sig000000e9)
  );
  MUXCY   blk0000003c (
    .CI(sig000000eb),
    .DI(sig00000461),
    .S(sig000000ce),
    .O(sig000000ea)
  );
  MUXCY   blk0000003d (
    .CI(sig000000ec),
    .DI(sig00000461),
    .S(sig000000cf),
    .O(sig000000eb)
  );
  MUXCY   blk0000003e (
    .CI(sig000000ed),
    .DI(sig00000461),
    .S(sig000000d0),
    .O(sig000000ec)
  );
  MUXCY   blk0000003f (
    .CI(sig000000ee),
    .DI(sig00000461),
    .S(sig000000d1),
    .O(sig000000ed)
  );
  MUXCY   blk00000040 (
    .CI(sig000000ef),
    .DI(sig00000461),
    .S(sig000000d2),
    .O(sig000000ee)
  );
  MUXCY   blk00000041 (
    .CI(sig00000001),
    .DI(sig00000461),
    .S(sig000000d3),
    .O(sig000000ef)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000042 (
    .C(clk),
    .CE(ce),
    .D(sig000000e7),
    .Q(sig000000a8)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000043 (
    .C(clk),
    .CE(ce),
    .D(sig00000097),
    .Q(sig000000f1)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000044 (
    .C(clk),
    .CE(ce),
    .D(sig00000096),
    .Q(sig000000f0)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000045 (
    .C(clk),
    .CE(ce),
    .D(sig000000f2),
    .Q(sig0000009f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000046 (
    .C(clk),
    .CE(ce),
    .D(sig000000f3),
    .Q(sig000000f2)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000047 (
    .C(clk),
    .CE(ce),
    .D(sig000000f4),
    .Q(sig000000f3)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000048 (
    .C(clk),
    .CE(ce),
    .D(sig000000f5),
    .Q(sig000000f4)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000049 (
    .C(clk),
    .CE(ce),
    .D(sig000000f6),
    .Q(sig000000f5)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000004a (
    .C(clk),
    .CE(ce),
    .D(sig000000f7),
    .Q(sig000000f6)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000004b (
    .C(clk),
    .CE(ce),
    .D(sig000000f8),
    .Q(sig000000f7)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000004c (
    .C(clk),
    .CE(ce),
    .D(sig000000f9),
    .Q(sig000000f8)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000004d (
    .C(clk),
    .CE(ce),
    .D(sig000000fa),
    .Q(sig000000f9)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000004e (
    .C(clk),
    .CE(ce),
    .D(sig000000fb),
    .Q(sig000000fa)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000004f (
    .C(clk),
    .CE(ce),
    .D(sig00000098),
    .Q(sig000000fb)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000050 (
    .C(clk),
    .CE(ce),
    .D(sig00000095),
    .Q(sig000000ff)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000051 (
    .C(clk),
    .CE(ce),
    .D(sig00000099),
    .Q(sig000000fe)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000052 (
    .C(clk),
    .CE(ce),
    .D(sig00000093),
    .Q(sig000000fd)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000053 (
    .C(clk),
    .CE(ce),
    .D(sig00000094),
    .Q(sig000000fc)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000054 (
    .C(clk),
    .CE(ce),
    .D(sig0000007e),
    .Q(sig00000007)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000055 (
    .C(clk),
    .CE(ce),
    .D(sig0000007b),
    .Q(sig00000005)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000056 (
    .C(clk),
    .CE(ce),
    .D(sig00000079),
    .Q(sig00000003)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000057 (
    .C(clk),
    .CE(ce),
    .D(sig0000007c),
    .Q(sig00000004)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000058 (
    .C(clk),
    .CE(ce),
    .D(sig0000007d),
    .Q(sig00000006)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000059 (
    .C(clk),
    .CE(ce),
    .D(sig000001c5),
    .Q(sig00000148)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000005a (
    .C(clk),
    .CE(ce),
    .D(sig000001c6),
    .Q(sig000001a2)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000005b (
    .C(clk),
    .CE(ce),
    .D(a[16]),
    .Q(sig000001a3)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000005c (
    .C(clk),
    .CE(ce),
    .D(a[15]),
    .Q(sig000001a4)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000005d (
    .C(clk),
    .CE(ce),
    .D(a[14]),
    .Q(sig000001a5)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000005e (
    .C(clk),
    .CE(ce),
    .D(a[13]),
    .Q(sig000001a6)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000005f (
    .C(clk),
    .CE(ce),
    .D(a[12]),
    .Q(sig000001a7)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000060 (
    .C(clk),
    .CE(ce),
    .D(a[11]),
    .Q(sig000001a8)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000061 (
    .C(clk),
    .CE(ce),
    .D(a[10]),
    .Q(sig000001a9)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000062 (
    .C(clk),
    .CE(ce),
    .D(a[9]),
    .Q(sig000001aa)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000063 (
    .C(clk),
    .CE(ce),
    .D(a[8]),
    .Q(sig000001ab)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000064 (
    .C(clk),
    .CE(ce),
    .D(a[7]),
    .Q(sig000001ac)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000065 (
    .C(clk),
    .CE(ce),
    .D(a[6]),
    .Q(sig000001ad)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000066 (
    .C(clk),
    .CE(ce),
    .D(a[5]),
    .Q(sig000001ae)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000067 (
    .C(clk),
    .CE(ce),
    .D(a[4]),
    .Q(sig000001af)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000068 (
    .C(clk),
    .CE(ce),
    .D(a[3]),
    .Q(sig000001b0)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000069 (
    .C(clk),
    .CE(ce),
    .D(a[2]),
    .Q(sig000001b1)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000006a (
    .C(clk),
    .CE(ce),
    .D(a[1]),
    .Q(sig000001b2)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000006b (
    .C(clk),
    .CE(ce),
    .D(a[0]),
    .Q(sig000001b3)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000006c (
    .C(clk),
    .CE(ce),
    .D(b[33]),
    .Q(sig000001b4)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000006d (
    .C(clk),
    .CE(ce),
    .D(b[32]),
    .Q(sig000001b5)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000006e (
    .C(clk),
    .CE(ce),
    .D(b[31]),
    .Q(sig000001b6)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000006f (
    .C(clk),
    .CE(ce),
    .D(b[30]),
    .Q(sig000001b7)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000070 (
    .C(clk),
    .CE(ce),
    .D(b[29]),
    .Q(sig000001b8)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000071 (
    .C(clk),
    .CE(ce),
    .D(b[28]),
    .Q(sig000001b9)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000072 (
    .C(clk),
    .CE(ce),
    .D(b[27]),
    .Q(sig000001ba)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000073 (
    .C(clk),
    .CE(ce),
    .D(b[26]),
    .Q(sig000001bb)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000074 (
    .C(clk),
    .CE(ce),
    .D(b[25]),
    .Q(sig000001bc)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000075 (
    .C(clk),
    .CE(ce),
    .D(b[24]),
    .Q(sig000001bd)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000076 (
    .C(clk),
    .CE(ce),
    .D(b[23]),
    .Q(sig000001be)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000077 (
    .C(clk),
    .CE(ce),
    .D(b[22]),
    .Q(sig000001bf)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000078 (
    .C(clk),
    .CE(ce),
    .D(b[21]),
    .Q(sig000001c0)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000079 (
    .C(clk),
    .CE(ce),
    .D(b[20]),
    .Q(sig000001c1)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000007a (
    .C(clk),
    .CE(ce),
    .D(b[19]),
    .Q(sig000001c2)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000007b (
    .C(clk),
    .CE(ce),
    .D(b[18]),
    .Q(sig000001c3)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000007c (
    .C(clk),
    .CE(ce),
    .D(b[17]),
    .Q(sig000001c4)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000007d (
    .C(clk),
    .CE(ce),
    .D(sig000001d1),
    .Q(sig0000001d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000007e (
    .C(clk),
    .CE(ce),
    .D(sig000001d0),
    .Q(sig0000001e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000007f (
    .C(clk),
    .CE(ce),
    .D(sig000001cf),
    .Q(sig0000001f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000080 (
    .C(clk),
    .CE(ce),
    .D(sig000001ce),
    .Q(sig00000020)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000081 (
    .C(clk),
    .CE(ce),
    .D(sig000001cd),
    .Q(sig00000021)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000082 (
    .C(clk),
    .CE(ce),
    .D(sig000001cc),
    .Q(sig00000022)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000083 (
    .C(clk),
    .CE(ce),
    .D(sig000001cb),
    .Q(sig00000023)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000084 (
    .C(clk),
    .CE(ce),
    .D(sig000001ca),
    .Q(sig00000024)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000085 (
    .C(clk),
    .CE(ce),
    .D(sig000001c9),
    .Q(sig00000025)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000086 (
    .C(clk),
    .CE(ce),
    .D(sig000001c8),
    .Q(sig00000026)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000087 (
    .C(clk),
    .CE(ce),
    .D(sig000001c7),
    .Q(sig00000027)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000088 (
    .C(clk),
    .CE(ce),
    .D(sig00000550),
    .Q(sig0000016d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000089 (
    .C(clk),
    .CE(ce),
    .D(sig0000016d),
    .Q(sig00000149)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000008a (
    .C(clk),
    .CE(ce),
    .D(sig00000002),
    .Q(sig00000460)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000008b (
    .C(clk),
    .CE(ce),
    .D(sig00000008),
    .Q(sig00000437)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000008c (
    .C(clk),
    .CE(ce),
    .D(sig00000009),
    .Q(sig0000047c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000008d (
    .C(clk),
    .CE(ce),
    .D(sig0000000a),
    .Q(sig0000047b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000008e (
    .C(clk),
    .CE(ce),
    .D(sig0000000b),
    .Q(sig0000047a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000008f (
    .C(clk),
    .CE(ce),
    .D(sig0000000c),
    .Q(sig00000479)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000090 (
    .C(clk),
    .CE(ce),
    .D(sig0000000d),
    .Q(sig00000478)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000091 (
    .C(clk),
    .CE(ce),
    .D(sig0000000e),
    .Q(sig00000477)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000092 (
    .C(clk),
    .CE(ce),
    .D(sig0000000f),
    .Q(sig00000476)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000093 (
    .C(clk),
    .CE(ce),
    .D(sig00000010),
    .Q(sig00000475)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000094 (
    .C(clk),
    .CE(ce),
    .D(sig00000011),
    .Q(sig00000474)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000095 (
    .C(clk),
    .CE(ce),
    .D(sig00000012),
    .Q(sig00000473)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000096 (
    .C(clk),
    .CE(ce),
    .D(sig00000013),
    .Q(sig00000472)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000097 (
    .C(clk),
    .CE(ce),
    .D(sig00000014),
    .Q(sig00000471)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000098 (
    .C(clk),
    .CE(ce),
    .D(sig00000015),
    .Q(sig00000470)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000099 (
    .C(clk),
    .CE(ce),
    .D(sig00000016),
    .Q(sig0000046f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000009a (
    .C(clk),
    .CE(ce),
    .D(sig00000017),
    .Q(sig0000046e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000009b (
    .C(clk),
    .CE(ce),
    .D(sig00000018),
    .Q(sig0000046d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000009c (
    .C(clk),
    .CE(ce),
    .D(sig00000019),
    .Q(sig0000046c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000009d (
    .C(clk),
    .CE(ce),
    .D(sig0000001a),
    .Q(sig0000046b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000009e (
    .C(clk),
    .CE(ce),
    .D(sig0000001b),
    .Q(sig0000046a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000009f (
    .C(clk),
    .CE(ce),
    .D(sig0000001c),
    .Q(sig00000469)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000a0 (
    .C(clk),
    .CE(ce),
    .D(sig0000001d),
    .Q(sig00000462)
  );
  MUXCY   blk000000a1 (
    .CI(sig00000001),
    .DI(sig00000461),
    .S(sig00000481),
    .O(sig0000047e)
  );
  MUXCY   blk000000a2 (
    .CI(sig0000047e),
    .DI(sig00000461),
    .S(sig00000461),
    .O(sig0000047f)
  );
  MUXCY   blk000000a3 (
    .CI(sig0000047f),
    .DI(sig00000001),
    .S(sig00000480),
    .O(sig0000045f)
  );
  XORCY   blk000000a4 (
    .CI(sig00000484),
    .LI(sig00000461),
    .O(sig00000482)
  );
  XORCY   blk000000a5 (
    .CI(sig00000486),
    .LI(sig00000451),
    .O(sig00000483)
  );
  MUXCY   blk000000a6 (
    .CI(sig00000486),
    .DI(sig00000461),
    .S(sig00000451),
    .O(sig00000484)
  );
  XORCY   blk000000a7 (
    .CI(sig00000488),
    .LI(sig00000450),
    .O(sig00000485)
  );
  MUXCY   blk000000a8 (
    .CI(sig00000488),
    .DI(sig00000461),
    .S(sig00000450),
    .O(sig00000486)
  );
  XORCY   blk000000a9 (
    .CI(sig0000048a),
    .LI(sig0000044f),
    .O(sig00000487)
  );
  MUXCY   blk000000aa (
    .CI(sig0000048a),
    .DI(sig00000461),
    .S(sig0000044f),
    .O(sig00000488)
  );
  XORCY   blk000000ab (
    .CI(sig0000048c),
    .LI(sig0000044e),
    .O(sig00000489)
  );
  MUXCY   blk000000ac (
    .CI(sig0000048c),
    .DI(sig00000461),
    .S(sig0000044e),
    .O(sig0000048a)
  );
  XORCY   blk000000ad (
    .CI(sig0000048e),
    .LI(sig0000044d),
    .O(sig0000048b)
  );
  MUXCY   blk000000ae (
    .CI(sig0000048e),
    .DI(sig00000461),
    .S(sig0000044d),
    .O(sig0000048c)
  );
  XORCY   blk000000af (
    .CI(sig00000490),
    .LI(sig0000044c),
    .O(sig0000048d)
  );
  MUXCY   blk000000b0 (
    .CI(sig00000490),
    .DI(sig00000461),
    .S(sig0000044c),
    .O(sig0000048e)
  );
  XORCY   blk000000b1 (
    .CI(sig00000492),
    .LI(sig0000044b),
    .O(sig0000048f)
  );
  MUXCY   blk000000b2 (
    .CI(sig00000492),
    .DI(sig00000461),
    .S(sig0000044b),
    .O(sig00000490)
  );
  XORCY   blk000000b3 (
    .CI(sig00000494),
    .LI(sig0000044a),
    .O(sig00000491)
  );
  MUXCY   blk000000b4 (
    .CI(sig00000494),
    .DI(sig00000461),
    .S(sig0000044a),
    .O(sig00000492)
  );
  XORCY   blk000000b5 (
    .CI(sig00000496),
    .LI(sig00000449),
    .O(sig00000493)
  );
  MUXCY   blk000000b6 (
    .CI(sig00000496),
    .DI(sig00000461),
    .S(sig00000449),
    .O(sig00000494)
  );
  XORCY   blk000000b7 (
    .CI(sig00000498),
    .LI(sig00000448),
    .O(sig00000495)
  );
  MUXCY   blk000000b8 (
    .CI(sig00000498),
    .DI(sig00000461),
    .S(sig00000448),
    .O(sig00000496)
  );
  XORCY   blk000000b9 (
    .CI(sig0000049a),
    .LI(sig00000447),
    .O(sig00000497)
  );
  MUXCY   blk000000ba (
    .CI(sig0000049a),
    .DI(sig00000461),
    .S(sig00000447),
    .O(sig00000498)
  );
  XORCY   blk000000bb (
    .CI(sig0000049c),
    .LI(sig00000446),
    .O(sig00000499)
  );
  MUXCY   blk000000bc (
    .CI(sig0000049c),
    .DI(sig00000461),
    .S(sig00000446),
    .O(sig0000049a)
  );
  XORCY   blk000000bd (
    .CI(sig0000049e),
    .LI(sig00000445),
    .O(sig0000049b)
  );
  MUXCY   blk000000be (
    .CI(sig0000049e),
    .DI(sig00000461),
    .S(sig00000445),
    .O(sig0000049c)
  );
  XORCY   blk000000bf (
    .CI(sig000004a0),
    .LI(sig00000444),
    .O(sig0000049d)
  );
  MUXCY   blk000000c0 (
    .CI(sig000004a0),
    .DI(sig00000461),
    .S(sig00000444),
    .O(sig0000049e)
  );
  XORCY   blk000000c1 (
    .CI(sig000004a2),
    .LI(sig00000443),
    .O(sig0000049f)
  );
  MUXCY   blk000000c2 (
    .CI(sig000004a2),
    .DI(sig00000461),
    .S(sig00000443),
    .O(sig000004a0)
  );
  XORCY   blk000000c3 (
    .CI(sig000004a4),
    .LI(sig00000442),
    .O(sig000004a1)
  );
  MUXCY   blk000000c4 (
    .CI(sig000004a4),
    .DI(sig00000461),
    .S(sig00000442),
    .O(sig000004a2)
  );
  XORCY   blk000000c5 (
    .CI(sig000004a6),
    .LI(sig00000441),
    .O(sig000004a3)
  );
  MUXCY   blk000000c6 (
    .CI(sig000004a6),
    .DI(sig00000461),
    .S(sig00000441),
    .O(sig000004a4)
  );
  XORCY   blk000000c7 (
    .CI(sig000004a8),
    .LI(sig00000440),
    .O(sig000004a5)
  );
  MUXCY   blk000000c8 (
    .CI(sig000004a8),
    .DI(sig00000461),
    .S(sig00000440),
    .O(sig000004a6)
  );
  XORCY   blk000000c9 (
    .CI(sig000004aa),
    .LI(sig0000043f),
    .O(sig000004a7)
  );
  MUXCY   blk000000ca (
    .CI(sig000004aa),
    .DI(sig00000461),
    .S(sig0000043f),
    .O(sig000004a8)
  );
  XORCY   blk000000cb (
    .CI(sig000004ac),
    .LI(sig0000043e),
    .O(sig000004a9)
  );
  MUXCY   blk000000cc (
    .CI(sig000004ac),
    .DI(sig00000461),
    .S(sig0000043e),
    .O(sig000004aa)
  );
  XORCY   blk000000cd (
    .CI(sig000004ae),
    .LI(sig0000043d),
    .O(sig000004ab)
  );
  MUXCY   blk000000ce (
    .CI(sig000004ae),
    .DI(sig00000461),
    .S(sig0000043d),
    .O(sig000004ac)
  );
  XORCY   blk000000cf (
    .CI(sig000004b0),
    .LI(sig0000043c),
    .O(sig000004ad)
  );
  MUXCY   blk000000d0 (
    .CI(sig000004b0),
    .DI(sig00000461),
    .S(sig0000043c),
    .O(sig000004ae)
  );
  XORCY   blk000000d1 (
    .CI(sig000004b2),
    .LI(sig0000043b),
    .O(sig000004af)
  );
  MUXCY   blk000000d2 (
    .CI(sig000004b2),
    .DI(sig00000461),
    .S(sig0000043b),
    .O(sig000004b0)
  );
  XORCY   blk000000d3 (
    .CI(sig000004b4),
    .LI(sig0000043a),
    .O(sig000004b1)
  );
  MUXCY   blk000000d4 (
    .CI(sig000004b4),
    .DI(sig00000461),
    .S(sig0000043a),
    .O(sig000004b2)
  );
  XORCY   blk000000d5 (
    .CI(sig000004b6),
    .LI(sig00000439),
    .O(sig000004b3)
  );
  MUXCY   blk000000d6 (
    .CI(sig000004b6),
    .DI(sig00000461),
    .S(sig00000439),
    .O(sig000004b4)
  );
  XORCY   blk000000d7 (
    .CI(sig0000045f),
    .LI(sig00000438),
    .O(sig000004b5)
  );
  MUXCY   blk000000d8 (
    .CI(sig0000045f),
    .DI(sig00000461),
    .S(sig00000438),
    .O(sig000004b6)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000d9 (
    .C(clk),
    .CE(ce),
    .D(sig00000482),
    .Q(sig0000045e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000da (
    .C(clk),
    .CE(ce),
    .D(sig000004d0),
    .Q(sig00000054)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000db (
    .C(clk),
    .CE(ce),
    .D(sig000004cf),
    .Q(sig00000055)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000dc (
    .C(clk),
    .CE(ce),
    .D(sig000004ce),
    .Q(sig00000056)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000dd (
    .C(clk),
    .CE(ce),
    .D(sig000004cd),
    .Q(sig00000057)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000de (
    .C(clk),
    .CE(ce),
    .D(sig000004cc),
    .Q(sig00000058)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000df (
    .C(clk),
    .CE(ce),
    .D(sig000004cb),
    .Q(sig00000059)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000e0 (
    .C(clk),
    .CE(ce),
    .D(sig000004ca),
    .Q(sig0000005a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000e1 (
    .C(clk),
    .CE(ce),
    .D(sig000004c9),
    .Q(sig0000005b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000e2 (
    .C(clk),
    .CE(ce),
    .D(sig000004c8),
    .Q(sig0000005c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000e3 (
    .C(clk),
    .CE(ce),
    .D(sig000004c7),
    .Q(sig0000005d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000e4 (
    .C(clk),
    .CE(ce),
    .D(sig000004c6),
    .Q(sig0000005e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000e5 (
    .C(clk),
    .CE(ce),
    .D(sig000004c5),
    .Q(sig0000005f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000e6 (
    .C(clk),
    .CE(ce),
    .D(sig000004c4),
    .Q(sig00000060)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000e7 (
    .C(clk),
    .CE(ce),
    .D(sig000004c3),
    .Q(sig00000061)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000e8 (
    .C(clk),
    .CE(ce),
    .D(sig000004c2),
    .Q(sig00000062)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000e9 (
    .C(clk),
    .CE(ce),
    .D(sig000004c1),
    .Q(sig00000063)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000ea (
    .C(clk),
    .CE(ce),
    .D(sig000004c0),
    .Q(sig00000064)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000eb (
    .C(clk),
    .CE(ce),
    .D(sig000004bf),
    .Q(sig00000065)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000ec (
    .C(clk),
    .CE(ce),
    .D(sig000004be),
    .Q(sig00000066)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000ed (
    .C(clk),
    .CE(ce),
    .D(sig000004bd),
    .Q(sig00000067)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000ee (
    .C(clk),
    .CE(ce),
    .D(sig000004bc),
    .Q(sig00000068)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000ef (
    .C(clk),
    .CE(ce),
    .D(sig000004bb),
    .Q(sig00000069)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000f0 (
    .C(clk),
    .CE(ce),
    .D(sig000004ba),
    .Q(sig0000006a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000f1 (
    .C(clk),
    .CE(ce),
    .D(sig000004b9),
    .Q(sig0000006b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000f2 (
    .C(clk),
    .CE(ce),
    .D(sig000004b8),
    .Q(sig0000006c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000f3 (
    .C(clk),
    .CE(ce),
    .D(sig000004b7),
    .Q(sig0000006d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000f4 (
    .C(clk),
    .CE(ce),
    .D(sig00000483),
    .Q(sig000004d0)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000f5 (
    .C(clk),
    .CE(ce),
    .D(sig00000485),
    .Q(sig000004cf)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000f6 (
    .C(clk),
    .CE(ce),
    .D(sig00000487),
    .Q(sig000004ce)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000f7 (
    .C(clk),
    .CE(ce),
    .D(sig00000489),
    .Q(sig000004cd)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000f8 (
    .C(clk),
    .CE(ce),
    .D(sig0000048b),
    .Q(sig000004cc)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000f9 (
    .C(clk),
    .CE(ce),
    .D(sig0000048d),
    .Q(sig000004cb)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000fa (
    .C(clk),
    .CE(ce),
    .D(sig0000048f),
    .Q(sig000004ca)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000fb (
    .C(clk),
    .CE(ce),
    .D(sig00000491),
    .Q(sig000004c9)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000fc (
    .C(clk),
    .CE(ce),
    .D(sig00000493),
    .Q(sig000004c8)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000fd (
    .C(clk),
    .CE(ce),
    .D(sig00000495),
    .Q(sig000004c7)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000fe (
    .C(clk),
    .CE(ce),
    .D(sig00000497),
    .Q(sig000004c6)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000ff (
    .C(clk),
    .CE(ce),
    .D(sig00000499),
    .Q(sig000004c5)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000100 (
    .C(clk),
    .CE(ce),
    .D(sig0000049b),
    .Q(sig000004c4)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000101 (
    .C(clk),
    .CE(ce),
    .D(sig0000049d),
    .Q(sig000004c3)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000102 (
    .C(clk),
    .CE(ce),
    .D(sig0000049f),
    .Q(sig000004c2)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000103 (
    .C(clk),
    .CE(ce),
    .D(sig000004a1),
    .Q(sig000004c1)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000104 (
    .C(clk),
    .CE(ce),
    .D(sig000004a3),
    .Q(sig000004c0)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000105 (
    .C(clk),
    .CE(ce),
    .D(sig000004a5),
    .Q(sig000004bf)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000106 (
    .C(clk),
    .CE(ce),
    .D(sig000004a7),
    .Q(sig000004be)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000107 (
    .C(clk),
    .CE(ce),
    .D(sig000004a9),
    .Q(sig000004bd)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000108 (
    .C(clk),
    .CE(ce),
    .D(sig000004ab),
    .Q(sig000004bc)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000109 (
    .C(clk),
    .CE(ce),
    .D(sig000004ad),
    .Q(sig000004bb)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000010a (
    .C(clk),
    .CE(ce),
    .D(sig000004af),
    .Q(sig000004ba)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000010b (
    .C(clk),
    .CE(ce),
    .D(sig000004b1),
    .Q(sig000004b9)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000010c (
    .C(clk),
    .CE(ce),
    .D(sig000004b3),
    .Q(sig000004b8)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000010d (
    .C(clk),
    .CE(ce),
    .D(sig000004b5),
    .Q(sig000004b7)
  );
  XORCY   blk0000010e (
    .CI(sig000004d2),
    .LI(sig00000461),
    .O(sig000004d1)
  );
  XORCY   blk0000010f (
    .CI(sig000004d4),
    .LI(sig0000041c),
    .O(NLW_blk0000010f_O_UNCONNECTED)
  );
  MUXCY   blk00000110 (
    .CI(sig000004d4),
    .DI(sig00000001),
    .S(sig0000041c),
    .O(sig000004d2)
  );
  XORCY   blk00000111 (
    .CI(sig000004d6),
    .LI(sig00000436),
    .O(sig000004d3)
  );
  MUXCY   blk00000112 (
    .CI(sig000004d6),
    .DI(sig00000461),
    .S(sig00000436),
    .O(sig000004d4)
  );
  XORCY   blk00000113 (
    .CI(sig000004d8),
    .LI(sig00000435),
    .O(sig000004d5)
  );
  MUXCY   blk00000114 (
    .CI(sig000004d8),
    .DI(sig00000461),
    .S(sig00000435),
    .O(sig000004d6)
  );
  XORCY   blk00000115 (
    .CI(sig000004da),
    .LI(sig00000434),
    .O(sig000004d7)
  );
  MUXCY   blk00000116 (
    .CI(sig000004da),
    .DI(sig00000461),
    .S(sig00000434),
    .O(sig000004d8)
  );
  XORCY   blk00000117 (
    .CI(sig000004dc),
    .LI(sig00000433),
    .O(sig000004d9)
  );
  MUXCY   blk00000118 (
    .CI(sig000004dc),
    .DI(sig00000461),
    .S(sig00000433),
    .O(sig000004da)
  );
  XORCY   blk00000119 (
    .CI(sig000004de),
    .LI(sig00000432),
    .O(sig000004db)
  );
  MUXCY   blk0000011a (
    .CI(sig000004de),
    .DI(sig00000461),
    .S(sig00000432),
    .O(sig000004dc)
  );
  XORCY   blk0000011b (
    .CI(sig000004e0),
    .LI(sig00000431),
    .O(sig000004dd)
  );
  MUXCY   blk0000011c (
    .CI(sig000004e0),
    .DI(sig00000461),
    .S(sig00000431),
    .O(sig000004de)
  );
  XORCY   blk0000011d (
    .CI(sig000004e2),
    .LI(sig00000430),
    .O(sig000004df)
  );
  MUXCY   blk0000011e (
    .CI(sig000004e2),
    .DI(sig00000461),
    .S(sig00000430),
    .O(sig000004e0)
  );
  XORCY   blk0000011f (
    .CI(sig000004e4),
    .LI(sig0000042f),
    .O(sig000004e1)
  );
  MUXCY   blk00000120 (
    .CI(sig000004e4),
    .DI(sig00000461),
    .S(sig0000042f),
    .O(sig000004e2)
  );
  XORCY   blk00000121 (
    .CI(sig000004e6),
    .LI(sig0000042e),
    .O(sig000004e3)
  );
  MUXCY   blk00000122 (
    .CI(sig000004e6),
    .DI(sig00000461),
    .S(sig0000042e),
    .O(sig000004e4)
  );
  XORCY   blk00000123 (
    .CI(sig000004e8),
    .LI(sig0000042d),
    .O(sig000004e5)
  );
  MUXCY   blk00000124 (
    .CI(sig000004e8),
    .DI(sig00000461),
    .S(sig0000042d),
    .O(sig000004e6)
  );
  XORCY   blk00000125 (
    .CI(sig000004ea),
    .LI(sig0000042c),
    .O(sig000004e7)
  );
  MUXCY   blk00000126 (
    .CI(sig000004ea),
    .DI(sig00000461),
    .S(sig0000042c),
    .O(sig000004e8)
  );
  XORCY   blk00000127 (
    .CI(sig000004ec),
    .LI(sig0000042b),
    .O(sig000004e9)
  );
  MUXCY   blk00000128 (
    .CI(sig000004ec),
    .DI(sig00000461),
    .S(sig0000042b),
    .O(sig000004ea)
  );
  XORCY   blk00000129 (
    .CI(sig000004ee),
    .LI(sig0000042a),
    .O(sig000004eb)
  );
  MUXCY   blk0000012a (
    .CI(sig000004ee),
    .DI(sig00000461),
    .S(sig0000042a),
    .O(sig000004ec)
  );
  XORCY   blk0000012b (
    .CI(sig000004f0),
    .LI(sig00000429),
    .O(sig000004ed)
  );
  MUXCY   blk0000012c (
    .CI(sig000004f0),
    .DI(sig00000461),
    .S(sig00000429),
    .O(sig000004ee)
  );
  XORCY   blk0000012d (
    .CI(sig000004f2),
    .LI(sig00000428),
    .O(sig000004ef)
  );
  MUXCY   blk0000012e (
    .CI(sig000004f2),
    .DI(sig00000461),
    .S(sig00000428),
    .O(sig000004f0)
  );
  XORCY   blk0000012f (
    .CI(sig000004f4),
    .LI(sig00000427),
    .O(sig000004f1)
  );
  MUXCY   blk00000130 (
    .CI(sig000004f4),
    .DI(sig00000461),
    .S(sig00000427),
    .O(sig000004f2)
  );
  XORCY   blk00000131 (
    .CI(sig000004f6),
    .LI(sig00000426),
    .O(sig000004f3)
  );
  MUXCY   blk00000132 (
    .CI(sig000004f6),
    .DI(sig00000461),
    .S(sig00000426),
    .O(sig000004f4)
  );
  XORCY   blk00000133 (
    .CI(sig000004f8),
    .LI(sig00000425),
    .O(sig000004f5)
  );
  MUXCY   blk00000134 (
    .CI(sig000004f8),
    .DI(sig00000461),
    .S(sig00000425),
    .O(sig000004f6)
  );
  XORCY   blk00000135 (
    .CI(sig000004fa),
    .LI(sig00000424),
    .O(sig000004f7)
  );
  MUXCY   blk00000136 (
    .CI(sig000004fa),
    .DI(sig00000461),
    .S(sig00000424),
    .O(sig000004f8)
  );
  XORCY   blk00000137 (
    .CI(sig000004fc),
    .LI(sig00000423),
    .O(sig000004f9)
  );
  MUXCY   blk00000138 (
    .CI(sig000004fc),
    .DI(sig00000461),
    .S(sig00000423),
    .O(sig000004fa)
  );
  XORCY   blk00000139 (
    .CI(sig000004fe),
    .LI(sig00000422),
    .O(sig000004fb)
  );
  MUXCY   blk0000013a (
    .CI(sig000004fe),
    .DI(sig00000461),
    .S(sig00000422),
    .O(sig000004fc)
  );
  XORCY   blk0000013b (
    .CI(sig00000500),
    .LI(sig00000421),
    .O(sig000004fd)
  );
  MUXCY   blk0000013c (
    .CI(sig00000500),
    .DI(sig00000461),
    .S(sig00000421),
    .O(sig000004fe)
  );
  XORCY   blk0000013d (
    .CI(sig00000502),
    .LI(sig00000420),
    .O(sig000004ff)
  );
  MUXCY   blk0000013e (
    .CI(sig00000502),
    .DI(sig00000461),
    .S(sig00000420),
    .O(sig00000500)
  );
  XORCY   blk0000013f (
    .CI(sig00000504),
    .LI(sig0000041f),
    .O(sig00000501)
  );
  MUXCY   blk00000140 (
    .CI(sig00000504),
    .DI(sig00000461),
    .S(sig0000041f),
    .O(sig00000502)
  );
  XORCY   blk00000141 (
    .CI(sig00000506),
    .LI(sig0000041e),
    .O(sig00000503)
  );
  MUXCY   blk00000142 (
    .CI(sig00000506),
    .DI(sig00000461),
    .S(sig0000041e),
    .O(sig00000504)
  );
  XORCY   blk00000143 (
    .CI(sig0000045e),
    .LI(sig0000041d),
    .O(sig00000505)
  );
  MUXCY   blk00000144 (
    .CI(sig0000045e),
    .DI(sig00000461),
    .S(sig0000041d),
    .O(sig00000506)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000145 (
    .C(clk),
    .CE(ce),
    .D(sig000004d1),
    .Q(sig0000045d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000146 (
    .C(clk),
    .CE(ce),
    .D(sig000004d3),
    .Q(sig0000003a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000147 (
    .C(clk),
    .CE(ce),
    .D(sig000004d5),
    .Q(sig0000003b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000148 (
    .C(clk),
    .CE(ce),
    .D(sig000004d7),
    .Q(sig0000003c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000149 (
    .C(clk),
    .CE(ce),
    .D(sig000004d9),
    .Q(sig0000003d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000014a (
    .C(clk),
    .CE(ce),
    .D(sig000004db),
    .Q(sig0000003e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000014b (
    .C(clk),
    .CE(ce),
    .D(sig000004dd),
    .Q(sig0000003f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000014c (
    .C(clk),
    .CE(ce),
    .D(sig000004df),
    .Q(sig00000040)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000014d (
    .C(clk),
    .CE(ce),
    .D(sig000004e1),
    .Q(sig00000041)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000014e (
    .C(clk),
    .CE(ce),
    .D(sig000004e3),
    .Q(sig00000042)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000014f (
    .C(clk),
    .CE(ce),
    .D(sig000004e5),
    .Q(sig00000043)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000150 (
    .C(clk),
    .CE(ce),
    .D(sig000004e7),
    .Q(sig00000044)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000151 (
    .C(clk),
    .CE(ce),
    .D(sig000004e9),
    .Q(sig00000045)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000152 (
    .C(clk),
    .CE(ce),
    .D(sig000004eb),
    .Q(sig00000046)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000153 (
    .C(clk),
    .CE(ce),
    .D(sig000004ed),
    .Q(sig00000047)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000154 (
    .C(clk),
    .CE(ce),
    .D(sig000004ef),
    .Q(sig00000048)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000155 (
    .C(clk),
    .CE(ce),
    .D(sig000004f1),
    .Q(sig00000049)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000156 (
    .C(clk),
    .CE(ce),
    .D(sig000004f3),
    .Q(sig0000004a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000157 (
    .C(clk),
    .CE(ce),
    .D(sig000004f5),
    .Q(sig0000004b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000158 (
    .C(clk),
    .CE(ce),
    .D(sig000004f7),
    .Q(sig0000004c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000159 (
    .C(clk),
    .CE(ce),
    .D(sig000004f9),
    .Q(sig0000004d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000015a (
    .C(clk),
    .CE(ce),
    .D(sig000004fb),
    .Q(sig0000004e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000015b (
    .C(clk),
    .CE(ce),
    .D(sig000004fd),
    .Q(sig0000004f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000015c (
    .C(clk),
    .CE(ce),
    .D(sig000004ff),
    .Q(sig00000050)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000015d (
    .C(clk),
    .CE(ce),
    .D(sig00000501),
    .Q(sig00000051)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000015e (
    .C(clk),
    .CE(ce),
    .D(sig00000503),
    .Q(sig00000052)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000015f (
    .C(clk),
    .CE(ce),
    .D(sig00000505),
    .Q(sig00000053)
  );
  XORCY   blk00000160 (
    .CI(sig00000507),
    .LI(sig0000045c),
    .O(sig0000006e)
  );
  XORCY   blk00000161 (
    .CI(sig00000508),
    .LI(sig0000055b),
    .O(sig0000006f)
  );
  MUXCY   blk00000162 (
    .CI(sig00000508),
    .DI(sig00000461),
    .S(sig0000055b),
    .O(sig00000507)
  );
  XORCY   blk00000163 (
    .CI(sig00000509),
    .LI(sig0000055c),
    .O(sig00000070)
  );
  MUXCY   blk00000164 (
    .CI(sig00000509),
    .DI(sig00000461),
    .S(sig0000055c),
    .O(sig00000508)
  );
  XORCY   blk00000165 (
    .CI(sig0000050a),
    .LI(sig0000055d),
    .O(sig00000071)
  );
  MUXCY   blk00000166 (
    .CI(sig0000050a),
    .DI(sig00000461),
    .S(sig0000055d),
    .O(sig00000509)
  );
  XORCY   blk00000167 (
    .CI(sig0000050b),
    .LI(sig0000055e),
    .O(sig00000072)
  );
  MUXCY   blk00000168 (
    .CI(sig0000050b),
    .DI(sig00000461),
    .S(sig0000055e),
    .O(sig0000050a)
  );
  XORCY   blk00000169 (
    .CI(sig0000050c),
    .LI(sig0000055f),
    .O(sig00000073)
  );
  MUXCY   blk0000016a (
    .CI(sig0000050c),
    .DI(sig00000461),
    .S(sig0000055f),
    .O(sig0000050b)
  );
  XORCY   blk0000016b (
    .CI(sig0000050d),
    .LI(sig00000560),
    .O(sig00000074)
  );
  MUXCY   blk0000016c (
    .CI(sig0000050d),
    .DI(sig00000461),
    .S(sig00000560),
    .O(sig0000050c)
  );
  XORCY   blk0000016d (
    .CI(sig0000050e),
    .LI(sig00000561),
    .O(sig00000075)
  );
  MUXCY   blk0000016e (
    .CI(sig0000050e),
    .DI(sig00000461),
    .S(sig00000561),
    .O(sig0000050d)
  );
  XORCY   blk0000016f (
    .CI(sig0000050f),
    .LI(sig00000562),
    .O(sig00000076)
  );
  MUXCY   blk00000170 (
    .CI(sig0000050f),
    .DI(sig00000461),
    .S(sig00000562),
    .O(sig0000050e)
  );
  XORCY   blk00000171 (
    .CI(sig00000510),
    .LI(sig00000563),
    .O(sig00000077)
  );
  MUXCY   blk00000172 (
    .CI(sig00000510),
    .DI(sig00000461),
    .S(sig00000563),
    .O(sig0000050f)
  );
  XORCY   blk00000173 (
    .CI(sig0000045d),
    .LI(sig00000564),
    .O(sig00000078)
  );
  MUXCY   blk00000174 (
    .CI(sig0000045d),
    .DI(sig00000461),
    .S(sig00000564),
    .O(sig00000510)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000175 (
    .C(clk),
    .D(sig00000544),
    .Q(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [51])
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000176 (
    .C(clk),
    .D(sig00000543),
    .Q(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [50])
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000177 (
    .C(clk),
    .D(sig00000542),
    .Q(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [49])
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000178 (
    .C(clk),
    .D(sig00000541),
    .Q(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [48])
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000179 (
    .C(clk),
    .D(sig00000540),
    .Q(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [47])
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000017a (
    .C(clk),
    .D(sig0000053f),
    .Q(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [46])
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000017b (
    .C(clk),
    .D(sig0000053e),
    .Q(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [45])
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000017c (
    .C(clk),
    .D(sig0000053d),
    .Q(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [44])
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000017d (
    .C(clk),
    .D(sig0000053c),
    .Q(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [43])
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000017e (
    .C(clk),
    .D(sig0000053b),
    .Q(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [42])
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000017f (
    .C(clk),
    .D(sig0000053a),
    .Q(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [41])
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000180 (
    .C(clk),
    .D(sig00000539),
    .Q(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [40])
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000181 (
    .C(clk),
    .D(sig00000538),
    .Q(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [39])
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000182 (
    .C(clk),
    .D(sig00000537),
    .Q(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [38])
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000183 (
    .C(clk),
    .D(sig00000536),
    .Q(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [37])
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000184 (
    .C(clk),
    .D(sig00000535),
    .Q(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [36])
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000185 (
    .C(clk),
    .D(sig00000534),
    .Q(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [35])
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000186 (
    .C(clk),
    .D(sig00000533),
    .Q(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [34])
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000187 (
    .C(clk),
    .D(sig00000532),
    .Q(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [33])
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000188 (
    .C(clk),
    .D(sig00000531),
    .Q(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [32])
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000189 (
    .C(clk),
    .D(sig00000530),
    .Q(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [31])
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000018a (
    .C(clk),
    .D(sig0000052f),
    .Q(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [30])
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000018b (
    .C(clk),
    .D(sig0000052e),
    .Q(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [29])
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000018c (
    .C(clk),
    .D(sig0000052d),
    .Q(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [28])
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000018d (
    .C(clk),
    .D(sig0000052c),
    .Q(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [27])
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000018e (
    .C(clk),
    .D(sig0000052b),
    .Q(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [26])
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000018f (
    .C(clk),
    .D(sig0000052a),
    .Q(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [25])
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000190 (
    .C(clk),
    .D(sig00000529),
    .Q(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [24])
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000191 (
    .C(clk),
    .D(sig00000528),
    .Q(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [23])
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000192 (
    .C(clk),
    .D(sig00000527),
    .Q(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [22])
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000193 (
    .C(clk),
    .D(sig00000526),
    .Q(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [21])
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000194 (
    .C(clk),
    .D(sig00000525),
    .Q(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [20])
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000195 (
    .C(clk),
    .D(sig00000524),
    .Q(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [19])
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000196 (
    .C(clk),
    .D(sig00000523),
    .Q(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [18])
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000197 (
    .C(clk),
    .D(sig00000522),
    .Q(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [17])
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000198 (
    .C(clk),
    .D(sig00000521),
    .Q(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [16])
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000199 (
    .C(clk),
    .D(sig00000520),
    .Q(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [15])
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000019a (
    .C(clk),
    .D(sig0000051f),
    .Q(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [14])
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000019b (
    .C(clk),
    .D(sig0000051e),
    .Q(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [13])
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000019c (
    .C(clk),
    .D(sig0000051d),
    .Q(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [12])
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000019d (
    .C(clk),
    .D(sig0000051c),
    .Q(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [11])
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000019e (
    .C(clk),
    .D(sig0000051b),
    .Q(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [10])
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000019f (
    .C(clk),
    .D(sig0000051a),
    .Q(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [9])
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001a0 (
    .C(clk),
    .D(sig00000519),
    .Q(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [8])
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001a1 (
    .C(clk),
    .D(sig00000518),
    .Q(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [7])
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001a2 (
    .C(clk),
    .D(sig00000517),
    .Q(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [6])
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001a3 (
    .C(clk),
    .D(sig00000516),
    .Q(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [5])
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001a4 (
    .C(clk),
    .D(sig00000515),
    .Q(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [4])
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001a5 (
    .C(clk),
    .D(sig00000514),
    .Q(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [3])
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001a6 (
    .C(clk),
    .D(sig00000513),
    .Q(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [2])
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001a7 (
    .C(clk),
    .D(sig00000512),
    .Q(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [1])
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001a8 (
    .C(clk),
    .D(sig00000511),
    .Q(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [0])
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001a9 (
    .C(clk),
    .D(sig0000054f),
    .Q(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/exp_op [10])
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001aa (
    .C(clk),
    .D(sig0000054e),
    .Q(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/exp_op [9])
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001ab (
    .C(clk),
    .D(sig0000054d),
    .Q(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/exp_op [8])
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001ac (
    .C(clk),
    .D(sig0000054c),
    .Q(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/exp_op [7])
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001ad (
    .C(clk),
    .D(sig0000054b),
    .Q(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/exp_op [6])
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001ae (
    .C(clk),
    .D(sig0000054a),
    .Q(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/exp_op [5])
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001af (
    .C(clk),
    .D(sig00000549),
    .Q(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/exp_op [4])
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001b0 (
    .C(clk),
    .D(sig00000548),
    .Q(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/exp_op [3])
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001b1 (
    .C(clk),
    .D(sig00000547),
    .Q(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/exp_op [2])
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001b2 (
    .C(clk),
    .D(sig00000546),
    .Q(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/exp_op [1])
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001b3 (
    .C(clk),
    .D(sig00000545),
    .Q(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/exp_op [0])
  );
  LUT6 #(
    .INIT ( 64'hFFFFFFFF11101010 ))
  blk000001b4 (
    .I0(sig0000009b),
    .I1(sig000000a1),
    .I2(sig0000009c),
    .I3(sig0000009e),
    .I4(sig00000008),
    .I5(sig000000a0),
    .O(sig00000091)
  );
  LUT6 #(
    .INIT ( 64'h0202020202000202 ))
  blk000001b5 (
    .I0(sig0000009d),
    .I1(sig000000a0),
    .I2(sig000000a1),
    .I3(sig0000009b),
    .I4(sig00000008),
    .I5(sig0000009c),
    .O(sig00000090)
  );
  LUT6 #(
    .INIT ( 64'h153E113215141110 ))
  blk000001b6 (
    .I0(sig000000a4),
    .I1(sig000000a7),
    .I2(sig000000a3),
    .I3(sig000000a6),
    .I4(sig000000a8),
    .I5(sig000000a5),
    .O(sig00000097)
  );
  LUT3 #(
    .INIT ( 8'h04 ))
  blk000001b7 (
    .I0(sig0000007e),
    .I1(sig0000007b),
    .I2(sig0000009a),
    .O(sig00000079)
  );
  LUT4 #(
    .INIT ( 16'hF888 ))
  blk000001b8 (
    .I0(sig000000b4),
    .I1(sig000000a9),
    .I2(sig000000aa),
    .I3(sig0000007a),
    .O(sig00000094)
  );
  LUT3 #(
    .INIT ( 8'h10 ))
  blk000001b9 (
    .I0(sig000000aa),
    .I1(sig000000b4),
    .I2(sig0000007a),
    .O(sig00000099)
  );
  LUT2 #(
    .INIT ( 4'hE ))
  blk000001ba (
    .I0(sig000000a4),
    .I1(sig000000a7),
    .O(sig00000096)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk000001bb (
    .I0(a[63]),
    .I1(b[63]),
    .O(sig0000008f)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk000001bc (
    .I0(a[52]),
    .I1(b[52]),
    .O(sig00000084)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk000001bd (
    .I0(a[53]),
    .I1(b[53]),
    .O(sig00000085)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk000001be (
    .I0(a[54]),
    .I1(b[54]),
    .O(sig00000086)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk000001bf (
    .I0(a[55]),
    .I1(b[55]),
    .O(sig00000087)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk000001c0 (
    .I0(a[56]),
    .I1(b[56]),
    .O(sig00000088)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk000001c1 (
    .I0(a[57]),
    .I1(b[57]),
    .O(sig00000089)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk000001c2 (
    .I0(a[58]),
    .I1(b[58]),
    .O(sig0000008a)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk000001c3 (
    .I0(a[59]),
    .I1(b[59]),
    .O(sig0000008b)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk000001c4 (
    .I0(a[60]),
    .I1(b[60]),
    .O(sig0000008c)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk000001c5 (
    .I0(a[61]),
    .I1(b[61]),
    .O(sig0000008d)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk000001c6 (
    .I0(a[62]),
    .I1(b[62]),
    .O(sig0000008e)
  );
  LUT2 #(
    .INIT ( 4'hE ))
  blk000001c7 (
    .I0(sig0000007b),
    .I1(sig0000007e),
    .O(sig0000007c)
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  blk000001c8 (
    .I0(sig0000007e),
    .I1(sig0000007b),
    .O(sig0000007d)
  );
  LUT2 #(
    .INIT ( 4'h1 ))
  blk000001c9 (
    .I0(sig000000a9),
    .I1(sig000000b4),
    .O(sig00000093)
  );
  LUT6 #(
    .INIT ( 64'h0000000000000001 ))
  blk000001ca (
    .I0(a[42]),
    .I1(a[43]),
    .I2(a[44]),
    .I3(a[45]),
    .I4(a[46]),
    .I5(a[47]),
    .O(sig000000cc)
  );
  LUT6 #(
    .INIT ( 64'h0000000000000001 ))
  blk000001cb (
    .I0(a[36]),
    .I1(a[37]),
    .I2(a[38]),
    .I3(a[39]),
    .I4(a[40]),
    .I5(a[41]),
    .O(sig000000cd)
  );
  LUT6 #(
    .INIT ( 64'h0000000000000001 ))
  blk000001cc (
    .I0(a[30]),
    .I1(a[31]),
    .I2(a[32]),
    .I3(a[33]),
    .I4(a[34]),
    .I5(a[35]),
    .O(sig000000ce)
  );
  LUT6 #(
    .INIT ( 64'h0000000000000001 ))
  blk000001cd (
    .I0(a[24]),
    .I1(a[25]),
    .I2(a[26]),
    .I3(a[27]),
    .I4(a[28]),
    .I5(a[29]),
    .O(sig000000cf)
  );
  LUT6 #(
    .INIT ( 64'h0000000000000001 ))
  blk000001ce (
    .I0(a[18]),
    .I1(a[19]),
    .I2(a[20]),
    .I3(a[21]),
    .I4(a[22]),
    .I5(a[23]),
    .O(sig000000d0)
  );
  LUT6 #(
    .INIT ( 64'h0000000000000001 ))
  blk000001cf (
    .I0(a[12]),
    .I1(a[13]),
    .I2(a[14]),
    .I3(a[15]),
    .I4(a[16]),
    .I5(a[17]),
    .O(sig000000d1)
  );
  LUT6 #(
    .INIT ( 64'h0000000000000001 ))
  blk000001d0 (
    .I0(a[6]),
    .I1(a[7]),
    .I2(a[8]),
    .I3(a[9]),
    .I4(a[10]),
    .I5(a[11]),
    .O(sig000000d2)
  );
  LUT6 #(
    .INIT ( 64'h0000000000000001 ))
  blk000001d1 (
    .I0(a[0]),
    .I1(a[1]),
    .I2(a[2]),
    .I3(a[3]),
    .I4(a[4]),
    .I5(a[5]),
    .O(sig000000d3)
  );
  LUT4 #(
    .INIT ( 16'h0001 ))
  blk000001d2 (
    .I0(a[48]),
    .I1(a[49]),
    .I2(a[50]),
    .I3(a[51]),
    .O(sig000000d4)
  );
  LUT6 #(
    .INIT ( 64'h0000000000000001 ))
  blk000001d3 (
    .I0(b[42]),
    .I1(b[43]),
    .I2(b[44]),
    .I3(b[45]),
    .I4(b[46]),
    .I5(b[47]),
    .O(sig000000d5)
  );
  LUT6 #(
    .INIT ( 64'h0000000000000001 ))
  blk000001d4 (
    .I0(b[36]),
    .I1(b[37]),
    .I2(b[38]),
    .I3(b[39]),
    .I4(b[40]),
    .I5(b[41]),
    .O(sig000000d6)
  );
  LUT6 #(
    .INIT ( 64'h0000000000000001 ))
  blk000001d5 (
    .I0(b[30]),
    .I1(b[31]),
    .I2(b[32]),
    .I3(b[33]),
    .I4(b[34]),
    .I5(b[35]),
    .O(sig000000d7)
  );
  LUT6 #(
    .INIT ( 64'h0000000000000001 ))
  blk000001d6 (
    .I0(b[24]),
    .I1(b[25]),
    .I2(b[26]),
    .I3(b[27]),
    .I4(b[28]),
    .I5(b[29]),
    .O(sig000000d8)
  );
  LUT6 #(
    .INIT ( 64'h0000000000000001 ))
  blk000001d7 (
    .I0(b[18]),
    .I1(b[19]),
    .I2(b[20]),
    .I3(b[21]),
    .I4(b[22]),
    .I5(b[23]),
    .O(sig000000d9)
  );
  LUT6 #(
    .INIT ( 64'h0000000000000001 ))
  blk000001d8 (
    .I0(b[12]),
    .I1(b[13]),
    .I2(b[14]),
    .I3(b[15]),
    .I4(b[16]),
    .I5(b[17]),
    .O(sig000000da)
  );
  LUT6 #(
    .INIT ( 64'h0000000000000001 ))
  blk000001d9 (
    .I0(b[6]),
    .I1(b[7]),
    .I2(b[8]),
    .I3(b[9]),
    .I4(b[10]),
    .I5(b[11]),
    .O(sig000000db)
  );
  LUT6 #(
    .INIT ( 64'h0000000000000001 ))
  blk000001da (
    .I0(b[0]),
    .I1(b[1]),
    .I2(b[2]),
    .I3(b[3]),
    .I4(b[4]),
    .I5(b[5]),
    .O(sig000000dc)
  );
  LUT4 #(
    .INIT ( 16'h0001 ))
  blk000001db (
    .I0(b[48]),
    .I1(b[49]),
    .I2(b[50]),
    .I3(b[51]),
    .O(sig000000dd)
  );
  LUT2 #(
    .INIT ( 4'h8 ))
  blk000001dc (
    .I0(sig00000364),
    .I1(sig000002b5),
    .O(sig000001c5)
  );
  LUT2 #(
    .INIT ( 4'h8 ))
  blk000001dd (
    .I0(sig00000365),
    .I1(sig000003d8),
    .O(sig000001c6)
  );
  LUT3 #(
    .INIT ( 8'hAC ))
  blk000001de (
    .I0(sig00000462),
    .I1(sig00000463),
    .I2(sig00000460),
    .O(sig0000041d)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000001df (
    .I0(sig0000046d),
    .I1(sig0000046c),
    .I2(sig00000460),
    .O(sig00000427)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000001e0 (
    .I0(sig0000046e),
    .I1(sig0000046d),
    .I2(sig00000460),
    .O(sig00000428)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000001e1 (
    .I0(sig0000046f),
    .I1(sig0000046e),
    .I2(sig00000460),
    .O(sig00000429)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000001e2 (
    .I0(sig00000470),
    .I1(sig0000046f),
    .I2(sig00000460),
    .O(sig0000042a)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000001e3 (
    .I0(sig00000471),
    .I1(sig00000470),
    .I2(sig00000460),
    .O(sig0000042b)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000001e4 (
    .I0(sig00000472),
    .I1(sig00000471),
    .I2(sig00000460),
    .O(sig0000042c)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000001e5 (
    .I0(sig00000473),
    .I1(sig00000472),
    .I2(sig00000460),
    .O(sig0000042d)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000001e6 (
    .I0(sig00000474),
    .I1(sig00000473),
    .I2(sig00000460),
    .O(sig0000042e)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000001e7 (
    .I0(sig00000475),
    .I1(sig00000474),
    .I2(sig00000460),
    .O(sig0000042f)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000001e8 (
    .I0(sig00000476),
    .I1(sig00000475),
    .I2(sig00000460),
    .O(sig00000430)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000001e9 (
    .I0(sig00000464),
    .I1(sig00000463),
    .I2(sig00000460),
    .O(sig0000041e)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk000001ea (
    .I0(sig00000460),
    .I1(sig00000476),
    .I2(sig00000477),
    .O(sig00000431)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk000001eb (
    .I0(sig00000460),
    .I1(sig00000477),
    .I2(sig00000478),
    .O(sig00000432)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk000001ec (
    .I0(sig00000460),
    .I1(sig00000478),
    .I2(sig00000479),
    .O(sig00000433)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk000001ed (
    .I0(sig00000460),
    .I1(sig00000479),
    .I2(sig0000047a),
    .O(sig00000434)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk000001ee (
    .I0(sig00000460),
    .I1(sig0000047a),
    .I2(sig0000047b),
    .O(sig00000435)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk000001ef (
    .I0(sig00000460),
    .I1(sig0000047b),
    .I2(sig0000047c),
    .O(sig00000436)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000001f0 (
    .I0(sig00000465),
    .I1(sig00000464),
    .I2(sig00000460),
    .O(sig0000041f)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000001f1 (
    .I0(sig00000466),
    .I1(sig00000465),
    .I2(sig00000460),
    .O(sig00000420)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000001f2 (
    .I0(sig00000467),
    .I1(sig00000466),
    .I2(sig00000460),
    .O(sig00000421)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000001f3 (
    .I0(sig00000468),
    .I1(sig00000467),
    .I2(sig00000460),
    .O(sig00000422)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000001f4 (
    .I0(sig00000469),
    .I1(sig00000468),
    .I2(sig00000460),
    .O(sig00000423)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000001f5 (
    .I0(sig0000046a),
    .I1(sig00000469),
    .I2(sig00000460),
    .O(sig00000424)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000001f6 (
    .I0(sig0000046b),
    .I1(sig0000046a),
    .I2(sig00000460),
    .O(sig00000425)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000001f7 (
    .I0(sig0000046c),
    .I1(sig0000046b),
    .I2(sig00000460),
    .O(sig00000426)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk000001f8 (
    .I0(sig00000550),
    .I1(sig0000047d),
    .O(sig0000045c)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000001f9 (
    .I0(sig00000037),
    .I1(sig00000036),
    .I2(sig00000008),
    .O(sig00000438)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000001fa (
    .I0(sig0000002d),
    .I1(sig0000002c),
    .I2(sig00000008),
    .O(sig00000442)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000001fb (
    .I0(sig0000002c),
    .I1(sig0000002b),
    .I2(sig00000008),
    .O(sig00000443)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000001fc (
    .I0(sig0000002b),
    .I1(sig0000002a),
    .I2(sig00000008),
    .O(sig00000444)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000001fd (
    .I0(sig0000002a),
    .I1(sig00000029),
    .I2(sig00000008),
    .O(sig00000445)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000001fe (
    .I0(sig00000029),
    .I1(sig00000028),
    .I2(sig00000008),
    .O(sig00000446)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000001ff (
    .I0(sig00000028),
    .I1(sig00000027),
    .I2(sig00000008),
    .O(sig00000447)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000200 (
    .I0(sig00000027),
    .I1(sig00000026),
    .I2(sig00000008),
    .O(sig00000448)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000201 (
    .I0(sig00000026),
    .I1(sig00000025),
    .I2(sig00000008),
    .O(sig00000449)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000202 (
    .I0(sig00000025),
    .I1(sig00000024),
    .I2(sig00000008),
    .O(sig0000044a)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000203 (
    .I0(sig00000024),
    .I1(sig00000023),
    .I2(sig00000008),
    .O(sig0000044b)
  );
  LUT3 #(
    .INIT ( 8'hAC ))
  blk00000204 (
    .I0(sig00000035),
    .I1(sig00000036),
    .I2(sig00000008),
    .O(sig00000439)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000205 (
    .I0(sig00000023),
    .I1(sig00000022),
    .I2(sig00000008),
    .O(sig0000044c)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000206 (
    .I0(sig00000022),
    .I1(sig00000021),
    .I2(sig00000008),
    .O(sig0000044d)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000207 (
    .I0(sig00000021),
    .I1(sig00000020),
    .I2(sig00000008),
    .O(sig0000044e)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000208 (
    .I0(sig00000020),
    .I1(sig0000001f),
    .I2(sig00000008),
    .O(sig0000044f)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000209 (
    .I0(sig0000001f),
    .I1(sig0000001e),
    .I2(sig00000008),
    .O(sig00000450)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk0000020a (
    .I0(sig00000008),
    .I1(sig0000001d),
    .I2(sig0000001e),
    .O(sig00000451)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk0000020b (
    .I0(sig00000035),
    .I1(sig00000034),
    .I2(sig00000008),
    .O(sig0000043a)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk0000020c (
    .I0(sig00000034),
    .I1(sig00000033),
    .I2(sig00000008),
    .O(sig0000043b)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk0000020d (
    .I0(sig00000033),
    .I1(sig00000032),
    .I2(sig00000008),
    .O(sig0000043c)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk0000020e (
    .I0(sig00000032),
    .I1(sig00000031),
    .I2(sig00000008),
    .O(sig0000043d)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk0000020f (
    .I0(sig00000031),
    .I1(sig00000030),
    .I2(sig00000008),
    .O(sig0000043e)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000210 (
    .I0(sig00000030),
    .I1(sig0000002f),
    .I2(sig00000008),
    .O(sig0000043f)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000211 (
    .I0(sig0000002f),
    .I1(sig0000002e),
    .I2(sig00000008),
    .O(sig00000440)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000212 (
    .I0(sig0000002e),
    .I1(sig0000002d),
    .I2(sig00000008),
    .O(sig00000441)
  );
  LUT5 #(
    .INIT ( 32'h0455FFDD ))
  blk00000213 (
    .I0(sig00000038),
    .I1(sig00000039),
    .I2(sig00000036),
    .I3(sig00000008),
    .I4(sig00000037),
    .O(sig00000480)
  );
  LUT3 #(
    .INIT ( 8'hEF ))
  blk00000214 (
    .I0(sig00000037),
    .I1(sig00000038),
    .I2(sig00000039),
    .O(sig00000481)
  );
  LUT5 #(
    .INIT ( 32'h44EE44E4 ))
  blk00000215 (
    .I0(ce),
    .I1(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/exp_op [1]),
    .I2(sig00000007),
    .I3(sig00000003),
    .I4(sig00000077),
    .O(sig00000546)
  );
  LUT5 #(
    .INIT ( 32'h44EE44E4 ))
  blk00000216 (
    .I0(ce),
    .I1(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/exp_op [3]),
    .I2(sig00000007),
    .I3(sig00000003),
    .I4(sig00000075),
    .O(sig00000548)
  );
  LUT5 #(
    .INIT ( 32'h44EE44E4 ))
  blk00000217 (
    .I0(ce),
    .I1(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/exp_op [4]),
    .I2(sig00000007),
    .I3(sig00000003),
    .I4(sig00000074),
    .O(sig00000549)
  );
  LUT5 #(
    .INIT ( 32'h44EE44E4 ))
  blk00000218 (
    .I0(ce),
    .I1(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/exp_op [2]),
    .I2(sig00000007),
    .I3(sig00000003),
    .I4(sig00000076),
    .O(sig00000547)
  );
  LUT5 #(
    .INIT ( 32'h44EE44E4 ))
  blk00000219 (
    .I0(ce),
    .I1(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/exp_op [6]),
    .I2(sig00000007),
    .I3(sig00000003),
    .I4(sig00000072),
    .O(sig0000054b)
  );
  LUT5 #(
    .INIT ( 32'h44EE44E4 ))
  blk0000021a (
    .I0(ce),
    .I1(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/exp_op [7]),
    .I2(sig00000007),
    .I3(sig00000003),
    .I4(sig00000071),
    .O(sig0000054c)
  );
  LUT5 #(
    .INIT ( 32'h44EE44E4 ))
  blk0000021b (
    .I0(ce),
    .I1(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/exp_op [9]),
    .I2(sig00000007),
    .I3(sig00000003),
    .I4(sig0000006f),
    .O(sig0000054e)
  );
  LUT5 #(
    .INIT ( 32'h44EE44E4 ))
  blk0000021c (
    .I0(ce),
    .I1(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/exp_op [10]),
    .I2(sig00000007),
    .I3(sig00000003),
    .I4(sig0000006e),
    .O(sig0000054f)
  );
  LUT5 #(
    .INIT ( 32'h44EE44E4 ))
  blk0000021d (
    .I0(ce),
    .I1(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/exp_op [5]),
    .I2(sig00000007),
    .I3(sig00000003),
    .I4(sig00000073),
    .O(sig0000054a)
  );
  LUT5 #(
    .INIT ( 32'h44EE44E4 ))
  blk0000021e (
    .I0(ce),
    .I1(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/exp_op [8]),
    .I2(sig00000007),
    .I3(sig00000003),
    .I4(sig00000070),
    .O(sig0000054d)
  );
  LUT4 #(
    .INIT ( 16'h7520 ))
  blk0000021f (
    .I0(ce),
    .I1(sig00000004),
    .I2(sig0000006c),
    .I3(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [1]),
    .O(sig00000512)
  );
  LUT4 #(
    .INIT ( 16'h7520 ))
  blk00000220 (
    .I0(ce),
    .I1(sig00000004),
    .I2(sig0000006b),
    .I3(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [2]),
    .O(sig00000513)
  );
  LUT4 #(
    .INIT ( 16'h7520 ))
  blk00000221 (
    .I0(ce),
    .I1(sig00000004),
    .I2(sig0000006d),
    .I3(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [0]),
    .O(sig00000511)
  );
  LUT4 #(
    .INIT ( 16'h7520 ))
  blk00000222 (
    .I0(ce),
    .I1(sig00000004),
    .I2(sig00000069),
    .I3(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [4]),
    .O(sig00000515)
  );
  LUT4 #(
    .INIT ( 16'h7520 ))
  blk00000223 (
    .I0(ce),
    .I1(sig00000004),
    .I2(sig00000068),
    .I3(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [5]),
    .O(sig00000516)
  );
  LUT4 #(
    .INIT ( 16'h7520 ))
  blk00000224 (
    .I0(ce),
    .I1(sig00000004),
    .I2(sig0000006a),
    .I3(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [3]),
    .O(sig00000514)
  );
  LUT4 #(
    .INIT ( 16'h7520 ))
  blk00000225 (
    .I0(ce),
    .I1(sig00000004),
    .I2(sig00000066),
    .I3(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [7]),
    .O(sig00000518)
  );
  LUT4 #(
    .INIT ( 16'h7520 ))
  blk00000226 (
    .I0(ce),
    .I1(sig00000004),
    .I2(sig00000065),
    .I3(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [8]),
    .O(sig00000519)
  );
  LUT4 #(
    .INIT ( 16'h7520 ))
  blk00000227 (
    .I0(ce),
    .I1(sig00000004),
    .I2(sig00000067),
    .I3(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [6]),
    .O(sig00000517)
  );
  LUT4 #(
    .INIT ( 16'h7520 ))
  blk00000228 (
    .I0(ce),
    .I1(sig00000004),
    .I2(sig00000063),
    .I3(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [10]),
    .O(sig0000051b)
  );
  LUT4 #(
    .INIT ( 16'h7520 ))
  blk00000229 (
    .I0(ce),
    .I1(sig00000004),
    .I2(sig00000062),
    .I3(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [11]),
    .O(sig0000051c)
  );
  LUT4 #(
    .INIT ( 16'h7520 ))
  blk0000022a (
    .I0(ce),
    .I1(sig00000004),
    .I2(sig00000064),
    .I3(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [9]),
    .O(sig0000051a)
  );
  LUT4 #(
    .INIT ( 16'h7520 ))
  blk0000022b (
    .I0(ce),
    .I1(sig00000004),
    .I2(sig0000005f),
    .I3(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [14]),
    .O(sig0000051f)
  );
  LUT4 #(
    .INIT ( 16'h7520 ))
  blk0000022c (
    .I0(ce),
    .I1(sig00000004),
    .I2(sig00000061),
    .I3(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [12]),
    .O(sig0000051d)
  );
  LUT4 #(
    .INIT ( 16'h7520 ))
  blk0000022d (
    .I0(ce),
    .I1(sig00000004),
    .I2(sig00000060),
    .I3(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [13]),
    .O(sig0000051e)
  );
  LUT4 #(
    .INIT ( 16'h7520 ))
  blk0000022e (
    .I0(ce),
    .I1(sig00000004),
    .I2(sig0000005d),
    .I3(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [16]),
    .O(sig00000521)
  );
  LUT4 #(
    .INIT ( 16'h7520 ))
  blk0000022f (
    .I0(ce),
    .I1(sig00000004),
    .I2(sig0000005c),
    .I3(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [17]),
    .O(sig00000522)
  );
  LUT4 #(
    .INIT ( 16'h7520 ))
  blk00000230 (
    .I0(ce),
    .I1(sig00000004),
    .I2(sig0000005e),
    .I3(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [15]),
    .O(sig00000520)
  );
  LUT4 #(
    .INIT ( 16'h7520 ))
  blk00000231 (
    .I0(ce),
    .I1(sig00000004),
    .I2(sig0000005a),
    .I3(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [19]),
    .O(sig00000524)
  );
  LUT4 #(
    .INIT ( 16'h7520 ))
  blk00000232 (
    .I0(ce),
    .I1(sig00000004),
    .I2(sig00000059),
    .I3(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [20]),
    .O(sig00000525)
  );
  LUT4 #(
    .INIT ( 16'h7520 ))
  blk00000233 (
    .I0(ce),
    .I1(sig00000004),
    .I2(sig0000005b),
    .I3(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [18]),
    .O(sig00000523)
  );
  LUT4 #(
    .INIT ( 16'h7520 ))
  blk00000234 (
    .I0(ce),
    .I1(sig00000004),
    .I2(sig00000056),
    .I3(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [23]),
    .O(sig00000528)
  );
  LUT4 #(
    .INIT ( 16'h7520 ))
  blk00000235 (
    .I0(ce),
    .I1(sig00000004),
    .I2(sig00000058),
    .I3(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [21]),
    .O(sig00000526)
  );
  LUT4 #(
    .INIT ( 16'h7520 ))
  blk00000236 (
    .I0(ce),
    .I1(sig00000004),
    .I2(sig00000057),
    .I3(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [22]),
    .O(sig00000527)
  );
  LUT4 #(
    .INIT ( 16'h7520 ))
  blk00000237 (
    .I0(ce),
    .I1(sig00000004),
    .I2(sig00000054),
    .I3(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [25]),
    .O(sig0000052a)
  );
  LUT4 #(
    .INIT ( 16'h7520 ))
  blk00000238 (
    .I0(ce),
    .I1(sig00000004),
    .I2(sig00000053),
    .I3(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [26]),
    .O(sig0000052b)
  );
  LUT4 #(
    .INIT ( 16'h7520 ))
  blk00000239 (
    .I0(ce),
    .I1(sig00000004),
    .I2(sig00000055),
    .I3(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [24]),
    .O(sig00000529)
  );
  LUT4 #(
    .INIT ( 16'h7520 ))
  blk0000023a (
    .I0(ce),
    .I1(sig00000004),
    .I2(sig00000051),
    .I3(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [28]),
    .O(sig0000052d)
  );
  LUT4 #(
    .INIT ( 16'h7520 ))
  blk0000023b (
    .I0(ce),
    .I1(sig00000004),
    .I2(sig00000050),
    .I3(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [29]),
    .O(sig0000052e)
  );
  LUT4 #(
    .INIT ( 16'h7520 ))
  blk0000023c (
    .I0(ce),
    .I1(sig00000004),
    .I2(sig00000052),
    .I3(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [27]),
    .O(sig0000052c)
  );
  LUT4 #(
    .INIT ( 16'h7520 ))
  blk0000023d (
    .I0(ce),
    .I1(sig00000004),
    .I2(sig0000004d),
    .I3(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [32]),
    .O(sig00000531)
  );
  LUT4 #(
    .INIT ( 16'h7520 ))
  blk0000023e (
    .I0(ce),
    .I1(sig00000004),
    .I2(sig0000004f),
    .I3(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [30]),
    .O(sig0000052f)
  );
  LUT4 #(
    .INIT ( 16'h7520 ))
  blk0000023f (
    .I0(ce),
    .I1(sig00000004),
    .I2(sig0000004e),
    .I3(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [31]),
    .O(sig00000530)
  );
  LUT4 #(
    .INIT ( 16'h7520 ))
  blk00000240 (
    .I0(ce),
    .I1(sig00000004),
    .I2(sig0000004b),
    .I3(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [34]),
    .O(sig00000533)
  );
  LUT4 #(
    .INIT ( 16'h7520 ))
  blk00000241 (
    .I0(ce),
    .I1(sig00000004),
    .I2(sig0000004a),
    .I3(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [35]),
    .O(sig00000534)
  );
  LUT4 #(
    .INIT ( 16'h7520 ))
  blk00000242 (
    .I0(ce),
    .I1(sig00000004),
    .I2(sig0000004c),
    .I3(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [33]),
    .O(sig00000532)
  );
  LUT4 #(
    .INIT ( 16'h7520 ))
  blk00000243 (
    .I0(ce),
    .I1(sig00000004),
    .I2(sig00000048),
    .I3(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [37]),
    .O(sig00000536)
  );
  LUT4 #(
    .INIT ( 16'h7520 ))
  blk00000244 (
    .I0(ce),
    .I1(sig00000004),
    .I2(sig00000047),
    .I3(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [38]),
    .O(sig00000537)
  );
  LUT4 #(
    .INIT ( 16'h7520 ))
  blk00000245 (
    .I0(ce),
    .I1(sig00000004),
    .I2(sig00000049),
    .I3(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [36]),
    .O(sig00000535)
  );
  LUT4 #(
    .INIT ( 16'h7520 ))
  blk00000246 (
    .I0(ce),
    .I1(sig00000004),
    .I2(sig00000044),
    .I3(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [41]),
    .O(sig0000053a)
  );
  LUT4 #(
    .INIT ( 16'h7520 ))
  blk00000247 (
    .I0(ce),
    .I1(sig00000004),
    .I2(sig00000046),
    .I3(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [39]),
    .O(sig00000538)
  );
  LUT4 #(
    .INIT ( 16'h7520 ))
  blk00000248 (
    .I0(ce),
    .I1(sig00000004),
    .I2(sig00000045),
    .I3(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [40]),
    .O(sig00000539)
  );
  LUT4 #(
    .INIT ( 16'h7520 ))
  blk00000249 (
    .I0(ce),
    .I1(sig00000004),
    .I2(sig00000042),
    .I3(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [43]),
    .O(sig0000053c)
  );
  LUT4 #(
    .INIT ( 16'h7520 ))
  blk0000024a (
    .I0(ce),
    .I1(sig00000004),
    .I2(sig00000041),
    .I3(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [44]),
    .O(sig0000053d)
  );
  LUT4 #(
    .INIT ( 16'h7520 ))
  blk0000024b (
    .I0(ce),
    .I1(sig00000004),
    .I2(sig00000043),
    .I3(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [42]),
    .O(sig0000053b)
  );
  LUT4 #(
    .INIT ( 16'h7520 ))
  blk0000024c (
    .I0(ce),
    .I1(sig00000004),
    .I2(sig0000003f),
    .I3(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [46]),
    .O(sig0000053f)
  );
  LUT4 #(
    .INIT ( 16'h7520 ))
  blk0000024d (
    .I0(ce),
    .I1(sig00000004),
    .I2(sig0000003e),
    .I3(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [47]),
    .O(sig00000540)
  );
  LUT4 #(
    .INIT ( 16'h7520 ))
  blk0000024e (
    .I0(ce),
    .I1(sig00000004),
    .I2(sig00000040),
    .I3(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [45]),
    .O(sig0000053e)
  );
  LUT4 #(
    .INIT ( 16'h7520 ))
  blk0000024f (
    .I0(ce),
    .I1(sig00000004),
    .I2(sig0000003b),
    .I3(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [50]),
    .O(sig00000543)
  );
  LUT4 #(
    .INIT ( 16'h7520 ))
  blk00000250 (
    .I0(ce),
    .I1(sig00000004),
    .I2(sig0000003d),
    .I3(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [48]),
    .O(sig00000541)
  );
  LUT4 #(
    .INIT ( 16'h7520 ))
  blk00000251 (
    .I0(ce),
    .I1(sig00000004),
    .I2(sig0000003c),
    .I3(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [49]),
    .O(sig00000542)
  );
  LUT5 #(
    .INIT ( 32'h77752220 ))
  blk00000252 (
    .I0(ce),
    .I1(sig00000003),
    .I2(sig00000007),
    .I3(sig00000078),
    .I4(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/exp_op [0]),
    .O(sig00000545)
  );
  LUT5 #(
    .INIT ( 32'h77752220 ))
  blk00000253 (
    .I0(ce),
    .I1(sig00000005),
    .I2(sig00000006),
    .I3(sig0000003a),
    .I4(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/MULT.OP/OP/mant_op [51]),
    .O(sig00000544)
  );
  LUT2 #(
    .INIT ( 4'h1 ))
  blk00000254 (
    .I0(sig0000009b),
    .I1(sig0000009c),
    .O(sig00000552)
  );
  LUT6 #(
    .INIT ( 64'hFFFFFFFF51554055 ))
  blk00000255 (
    .I0(sig000000a0),
    .I1(sig00000008),
    .I2(sig0000009e),
    .I3(sig00000552),
    .I4(sig0000009d),
    .I5(sig000000a1),
    .O(sig00000092)
  );
  LUT2 #(
    .INIT ( 4'hB ))
  blk00000256 (
    .I0(sig000000a6),
    .I1(sig000000a5),
    .O(sig00000553)
  );
  LUT6 #(
    .INIT ( 64'h0020202000AAAAAA ))
  blk00000257 (
    .I0(sig000000a2),
    .I1(sig000000a3),
    .I2(sig000000a8),
    .I3(sig00000553),
    .I4(sig000000a4),
    .I5(sig000000a7),
    .O(sig00000098)
  );
  LUT5 #(
    .INIT ( 32'h80000000 ))
  blk00000258 (
    .I0(sig000000ab),
    .I1(sig000000ae),
    .I2(sig000000ad),
    .I3(sig000000ac),
    .I4(sig000000a9),
    .O(sig00000554)
  );
  LUT6 #(
    .INIT ( 64'h8000000000000000 ))
  blk00000259 (
    .I0(sig000000b0),
    .I1(sig000000af),
    .I2(sig000000b3),
    .I3(sig000000b2),
    .I4(sig000000b1),
    .I5(sig00000554),
    .O(sig0000007a)
  );
  LUT6 #(
    .INIT ( 64'h8000000000000000 ))
  blk0000025a (
    .I0(a[57]),
    .I1(a[56]),
    .I2(a[55]),
    .I3(a[54]),
    .I4(a[53]),
    .I5(a[52]),
    .O(sig00000555)
  );
  LUT6 #(
    .INIT ( 64'h8000000000000000 ))
  blk0000025b (
    .I0(a[62]),
    .I1(a[61]),
    .I2(a[60]),
    .I3(a[59]),
    .I4(a[58]),
    .I5(sig00000555),
    .O(sig00000080)
  );
  LUT6 #(
    .INIT ( 64'hFFFFFFFFFFFFFFFE ))
  blk0000025c (
    .I0(a[57]),
    .I1(a[56]),
    .I2(a[55]),
    .I3(a[54]),
    .I4(a[53]),
    .I5(a[52]),
    .O(sig00000556)
  );
  LUT6 #(
    .INIT ( 64'h0000000000000001 ))
  blk0000025d (
    .I0(a[62]),
    .I1(a[61]),
    .I2(a[60]),
    .I3(a[59]),
    .I4(a[58]),
    .I5(sig00000556),
    .O(sig00000081)
  );
  LUT6 #(
    .INIT ( 64'h8000000000000000 ))
  blk0000025e (
    .I0(b[57]),
    .I1(b[56]),
    .I2(b[55]),
    .I3(b[54]),
    .I4(b[53]),
    .I5(b[52]),
    .O(sig00000557)
  );
  LUT6 #(
    .INIT ( 64'h8000000000000000 ))
  blk0000025f (
    .I0(b[62]),
    .I1(b[61]),
    .I2(b[60]),
    .I3(b[59]),
    .I4(b[58]),
    .I5(sig00000557),
    .O(sig00000082)
  );
  LUT6 #(
    .INIT ( 64'hFFFFFFFFFFFFFFFE ))
  blk00000260 (
    .I0(b[57]),
    .I1(b[56]),
    .I2(b[55]),
    .I3(b[54]),
    .I4(b[53]),
    .I5(b[52]),
    .O(sig00000558)
  );
  LUT6 #(
    .INIT ( 64'h0000000000000001 ))
  blk00000261 (
    .I0(b[62]),
    .I1(b[61]),
    .I2(b[60]),
    .I3(b[59]),
    .I4(b[58]),
    .I5(sig00000558),
    .O(sig00000083)
  );
  LUT6 #(
    .INIT ( 64'h0000000000010000 ))
  blk00000262 (
    .I0(sig000000aa),
    .I1(sig000000ab),
    .I2(sig000000ac),
    .I3(sig000000ad),
    .I4(sig000000b4),
    .I5(sig000000ae),
    .O(sig00000559)
  );
  LUT6 #(
    .INIT ( 64'h0000000000000001 ))
  blk00000263 (
    .I0(sig000000b0),
    .I1(sig000000af),
    .I2(sig000000b1),
    .I3(sig000000b2),
    .I4(sig000000b3),
    .I5(sig000000a9),
    .O(sig0000055a)
  );
  LUT2 #(
    .INIT ( 4'h8 ))
  blk00000264 (
    .I0(sig00000559),
    .I1(sig0000055a),
    .O(sig00000095)
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  blk00000265 (
    .I0(sig0000045b),
    .O(sig0000055b)
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  blk00000266 (
    .I0(sig0000045a),
    .O(sig0000055c)
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  blk00000267 (
    .I0(sig00000459),
    .O(sig0000055d)
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  blk00000268 (
    .I0(sig00000458),
    .O(sig0000055e)
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  blk00000269 (
    .I0(sig00000457),
    .O(sig0000055f)
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  blk0000026a (
    .I0(sig00000456),
    .O(sig00000560)
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  blk0000026b (
    .I0(sig00000455),
    .O(sig00000561)
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  blk0000026c (
    .I0(sig00000454),
    .O(sig00000562)
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  blk0000026d (
    .I0(sig00000453),
    .O(sig00000563)
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  blk0000026e (
    .I0(sig00000452),
    .O(sig00000564)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk0000026f (
    .I0(ce),
    .I1(sig00000551),
    .I2(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/HND_SHK/RDY ),
    .O(sig00000565)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000270 (
    .C(clk),
    .D(sig00000565),
    .Q(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/HND_SHK/RDY )
  );
  INV   blk00000271 (
    .I(sig00000008),
    .O(sig00000002)
  );
  INV   blk00000272 (
    .I(sig00000437),
    .O(sig0000041c)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000273 (
    .A0(sig00000461),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000001),
    .CE(ce),
    .CLK(clk),
    .D(sig000000f1),
    .Q(sig00000566),
    .Q15(NLW_blk00000273_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000274 (
    .C(clk),
    .CE(ce),
    .D(sig00000566),
    .Q(sig000000a1)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000275 (
    .A0(sig00000461),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000001),
    .CE(ce),
    .CLK(clk),
    .D(sig000000f0),
    .Q(sig00000567),
    .Q15(NLW_blk00000275_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000276 (
    .C(clk),
    .CE(ce),
    .D(sig00000567),
    .Q(sig000000a0)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000277 (
    .A0(sig00000461),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000001),
    .CE(ce),
    .CLK(clk),
    .D(sig000000ff),
    .Q(sig00000568),
    .Q15(NLW_blk00000277_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000278 (
    .C(clk),
    .CE(ce),
    .D(sig00000568),
    .Q(sig0000009d)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000279 (
    .A0(sig00000461),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000001),
    .CE(ce),
    .CLK(clk),
    .D(sig000000fe),
    .Q(sig00000569),
    .Q15(NLW_blk00000279_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000027a (
    .C(clk),
    .CE(ce),
    .D(sig00000569),
    .Q(sig0000009e)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk0000027b (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig00000148),
    .Q(sig0000056a),
    .Q15(NLW_blk0000027b_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000027c (
    .C(clk),
    .CE(ce),
    .D(sig0000056a),
    .Q(sig00000039)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk0000027d (
    .A0(sig00000461),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000001),
    .CE(ce),
    .CLK(clk),
    .D(sig000000fd),
    .Q(sig0000056b),
    .Q15(NLW_blk0000027d_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000027e (
    .C(clk),
    .CE(ce),
    .D(sig0000056b),
    .Q(sig0000009b)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk0000027f (
    .A0(sig00000461),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000001),
    .CE(ce),
    .CLK(clk),
    .D(sig000000fc),
    .Q(sig0000056c),
    .Q15(NLW_blk0000027f_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000280 (
    .C(clk),
    .CE(ce),
    .D(sig0000056c),
    .Q(sig0000009c)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000281 (
    .A0(sig00000461),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(a[33]),
    .Q(sig0000056d),
    .Q15(NLW_blk00000281_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000282 (
    .C(clk),
    .CE(ce),
    .D(sig0000056d),
    .Q(sig00000191)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000283 (
    .A0(sig00000461),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig000001a2),
    .Q(sig0000056e),
    .Q15(NLW_blk00000283_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000284 (
    .C(clk),
    .CE(ce),
    .D(sig0000056e),
    .Q(sig00000364)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000285 (
    .A0(sig00000461),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig000003d9),
    .Q(sig0000056f),
    .Q15(NLW_blk00000285_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000286 (
    .C(clk),
    .CE(ce),
    .D(sig0000056f),
    .Q(sig000003d8)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000287 (
    .A0(sig00000461),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(a[30]),
    .Q(sig00000570),
    .Q15(NLW_blk00000287_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000288 (
    .C(clk),
    .CE(ce),
    .D(sig00000570),
    .Q(sig00000194)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000289 (
    .A0(sig00000461),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(a[32]),
    .Q(sig00000571),
    .Q15(NLW_blk00000289_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000028a (
    .C(clk),
    .CE(ce),
    .D(sig00000571),
    .Q(sig00000192)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk0000028b (
    .A0(sig00000461),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(a[31]),
    .Q(sig00000572),
    .Q15(NLW_blk0000028b_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000028c (
    .C(clk),
    .CE(ce),
    .D(sig00000572),
    .Q(sig00000193)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk0000028d (
    .A0(sig00000461),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(a[29]),
    .Q(sig00000573),
    .Q15(NLW_blk0000028d_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000028e (
    .C(clk),
    .CE(ce),
    .D(sig00000573),
    .Q(sig00000195)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk0000028f (
    .A0(sig00000461),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(a[28]),
    .Q(sig00000574),
    .Q15(NLW_blk0000028f_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000290 (
    .C(clk),
    .CE(ce),
    .D(sig00000574),
    .Q(sig00000196)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000291 (
    .A0(sig00000461),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(a[27]),
    .Q(sig00000575),
    .Q15(NLW_blk00000291_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000292 (
    .C(clk),
    .CE(ce),
    .D(sig00000575),
    .Q(sig00000197)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000293 (
    .A0(sig00000461),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(a[26]),
    .Q(sig00000576),
    .Q15(NLW_blk00000293_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000294 (
    .C(clk),
    .CE(ce),
    .D(sig00000576),
    .Q(sig00000198)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000295 (
    .A0(sig00000461),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(a[23]),
    .Q(sig00000577),
    .Q15(NLW_blk00000295_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000296 (
    .C(clk),
    .CE(ce),
    .D(sig00000577),
    .Q(sig0000019b)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000297 (
    .A0(sig00000461),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(a[25]),
    .Q(sig00000578),
    .Q15(NLW_blk00000297_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000298 (
    .C(clk),
    .CE(ce),
    .D(sig00000578),
    .Q(sig00000199)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000299 (
    .A0(sig00000461),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(a[24]),
    .Q(sig00000579),
    .Q15(NLW_blk00000299_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000029a (
    .C(clk),
    .CE(ce),
    .D(sig00000579),
    .Q(sig0000019a)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk0000029b (
    .A0(sig00000461),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(a[20]),
    .Q(sig0000057a),
    .Q15(NLW_blk0000029b_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000029c (
    .C(clk),
    .CE(ce),
    .D(sig0000057a),
    .Q(sig0000019e)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk0000029d (
    .A0(sig00000461),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(a[22]),
    .Q(sig0000057b),
    .Q15(NLW_blk0000029d_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000029e (
    .C(clk),
    .CE(ce),
    .D(sig0000057b),
    .Q(sig0000019c)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk0000029f (
    .A0(sig00000461),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(a[21]),
    .Q(sig0000057c),
    .Q15(NLW_blk0000029f_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002a0 (
    .C(clk),
    .CE(ce),
    .D(sig0000057c),
    .Q(sig0000019d)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000002a1 (
    .A0(sig00000461),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(a[17]),
    .Q(sig0000057d),
    .Q15(NLW_blk000002a1_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002a2 (
    .C(clk),
    .CE(ce),
    .D(sig0000057d),
    .Q(sig000001a1)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000002a3 (
    .A0(sig00000461),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(a[19]),
    .Q(sig0000057e),
    .Q15(NLW_blk000002a3_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002a4 (
    .C(clk),
    .CE(ce),
    .D(sig0000057e),
    .Q(sig0000019f)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000002a5 (
    .A0(sig00000461),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(a[18]),
    .Q(sig0000057f),
    .Q15(NLW_blk000002a5_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002a6 (
    .C(clk),
    .CE(ce),
    .D(sig0000057f),
    .Q(sig000001a0)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000002a7 (
    .A0(sig00000461),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig00000236),
    .Q(sig00000580),
    .Q15(NLW_blk000002a7_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002a8 (
    .C(clk),
    .CE(ce),
    .D(sig00000580),
    .Q(sig00000028)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000002a9 (
    .A0(sig00000461),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig00000235),
    .Q(sig00000581),
    .Q15(NLW_blk000002a9_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002aa (
    .C(clk),
    .CE(ce),
    .D(sig00000581),
    .Q(sig00000029)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000002ab (
    .A0(sig00000461),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig00000234),
    .Q(sig00000582),
    .Q15(NLW_blk000002ab_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002ac (
    .C(clk),
    .CE(ce),
    .D(sig00000582),
    .Q(sig0000002a)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000002ad (
    .A0(sig00000461),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig00000233),
    .Q(sig00000583),
    .Q15(NLW_blk000002ad_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002ae (
    .C(clk),
    .CE(ce),
    .D(sig00000583),
    .Q(sig0000002b)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000002af (
    .A0(sig00000461),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig00000230),
    .Q(sig00000584),
    .Q15(NLW_blk000002af_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002b0 (
    .C(clk),
    .CE(ce),
    .D(sig00000584),
    .Q(sig0000002e)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000002b1 (
    .A0(sig00000461),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig00000232),
    .Q(sig00000585),
    .Q15(NLW_blk000002b1_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002b2 (
    .C(clk),
    .CE(ce),
    .D(sig00000585),
    .Q(sig0000002c)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000002b3 (
    .A0(sig00000461),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig00000231),
    .Q(sig00000586),
    .Q15(NLW_blk000002b3_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002b4 (
    .C(clk),
    .CE(ce),
    .D(sig00000586),
    .Q(sig0000002d)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000002b5 (
    .A0(sig00000461),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig0000022d),
    .Q(sig00000587),
    .Q15(NLW_blk000002b5_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002b6 (
    .C(clk),
    .CE(ce),
    .D(sig00000587),
    .Q(sig00000031)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000002b7 (
    .A0(sig00000461),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig0000022f),
    .Q(sig00000588),
    .Q15(NLW_blk000002b7_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002b8 (
    .C(clk),
    .CE(ce),
    .D(sig00000588),
    .Q(sig0000002f)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000002b9 (
    .A0(sig00000461),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig0000022e),
    .Q(sig00000589),
    .Q15(NLW_blk000002b9_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002ba (
    .C(clk),
    .CE(ce),
    .D(sig00000589),
    .Q(sig00000030)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000002bb (
    .A0(sig00000461),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig0000022a),
    .Q(sig0000058a),
    .Q15(NLW_blk000002bb_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002bc (
    .C(clk),
    .CE(ce),
    .D(sig0000058a),
    .Q(sig00000034)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000002bd (
    .A0(sig00000461),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig0000022c),
    .Q(sig0000058b),
    .Q15(NLW_blk000002bd_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002be (
    .C(clk),
    .CE(ce),
    .D(sig0000058b),
    .Q(sig00000032)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000002bf (
    .A0(sig00000461),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig0000022b),
    .Q(sig0000058c),
    .Q15(NLW_blk000002bf_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002c0 (
    .C(clk),
    .CE(ce),
    .D(sig0000058c),
    .Q(sig00000033)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000002c1 (
    .A0(sig00000461),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig00000229),
    .Q(sig0000058d),
    .Q15(NLW_blk000002c1_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002c2 (
    .C(clk),
    .CE(ce),
    .D(sig0000058d),
    .Q(sig00000035)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000002c3 (
    .A0(sig00000461),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig00000228),
    .Q(sig0000058e),
    .Q15(NLW_blk000002c3_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002c4 (
    .C(clk),
    .CE(ce),
    .D(sig0000058e),
    .Q(sig00000036)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000002c5 (
    .A0(sig00000461),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig00000227),
    .Q(sig0000058f),
    .Q15(NLW_blk000002c5_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002c6 (
    .C(clk),
    .CE(ce),
    .D(sig0000058f),
    .Q(sig00000037)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000002c7 (
    .A0(sig00000461),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig00000226),
    .Q(sig00000590),
    .Q15(NLW_blk000002c7_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002c8 (
    .C(clk),
    .CE(ce),
    .D(sig00000590),
    .Q(sig00000038)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000002c9 (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(a[49]),
    .Q(sig00000591),
    .Q15(NLW_blk000002c9_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002ca (
    .C(clk),
    .CE(ce),
    .D(sig00000591),
    .Q(sig00000170)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000002cb (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(a[51]),
    .Q(sig00000592),
    .Q15(NLW_blk000002cb_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002cc (
    .C(clk),
    .CE(ce),
    .D(sig00000592),
    .Q(sig0000016e)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000002cd (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(a[50]),
    .Q(sig00000593),
    .Q15(NLW_blk000002cd_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002ce (
    .C(clk),
    .CE(ce),
    .D(sig00000593),
    .Q(sig0000016f)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000002cf (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(a[46]),
    .Q(sig00000594),
    .Q15(NLW_blk000002cf_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002d0 (
    .C(clk),
    .CE(ce),
    .D(sig00000594),
    .Q(sig00000173)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000002d1 (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(a[48]),
    .Q(sig00000595),
    .Q15(NLW_blk000002d1_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002d2 (
    .C(clk),
    .CE(ce),
    .D(sig00000595),
    .Q(sig00000171)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000002d3 (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(a[47]),
    .Q(sig00000596),
    .Q15(NLW_blk000002d3_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002d4 (
    .C(clk),
    .CE(ce),
    .D(sig00000596),
    .Q(sig00000172)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000002d5 (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(a[43]),
    .Q(sig00000597),
    .Q15(NLW_blk000002d5_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002d6 (
    .C(clk),
    .CE(ce),
    .D(sig00000597),
    .Q(sig00000176)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000002d7 (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(a[45]),
    .Q(sig00000598),
    .Q15(NLW_blk000002d7_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002d8 (
    .C(clk),
    .CE(ce),
    .D(sig00000598),
    .Q(sig00000174)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000002d9 (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(a[44]),
    .Q(sig00000599),
    .Q15(NLW_blk000002d9_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002da (
    .C(clk),
    .CE(ce),
    .D(sig00000599),
    .Q(sig00000175)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000002db (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(a[42]),
    .Q(sig0000059a),
    .Q15(NLW_blk000002db_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002dc (
    .C(clk),
    .CE(ce),
    .D(sig0000059a),
    .Q(sig00000177)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000002dd (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(a[41]),
    .Q(sig0000059b),
    .Q15(NLW_blk000002dd_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002de (
    .C(clk),
    .CE(ce),
    .D(sig0000059b),
    .Q(sig00000178)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000002df (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(a[40]),
    .Q(sig0000059c),
    .Q15(NLW_blk000002df_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002e0 (
    .C(clk),
    .CE(ce),
    .D(sig0000059c),
    .Q(sig00000179)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000002e1 (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(a[39]),
    .Q(sig0000059d),
    .Q15(NLW_blk000002e1_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002e2 (
    .C(clk),
    .CE(ce),
    .D(sig0000059d),
    .Q(sig0000017a)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000002e3 (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(a[36]),
    .Q(sig0000059e),
    .Q15(NLW_blk000002e3_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002e4 (
    .C(clk),
    .CE(ce),
    .D(sig0000059e),
    .Q(sig0000017d)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000002e5 (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(a[38]),
    .Q(sig0000059f),
    .Q15(NLW_blk000002e5_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002e6 (
    .C(clk),
    .CE(ce),
    .D(sig0000059f),
    .Q(sig0000017b)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000002e7 (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(a[37]),
    .Q(sig000005a0),
    .Q15(NLW_blk000002e7_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002e8 (
    .C(clk),
    .CE(ce),
    .D(sig000005a0),
    .Q(sig0000017c)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000002e9 (
    .A0(sig00000461),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig00000001),
    .Q(sig000005a1),
    .Q15(NLW_blk000002e9_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002ea (
    .C(clk),
    .CE(ce),
    .D(sig000005a1),
    .Q(sig00000550)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000002eb (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(a[35]),
    .Q(sig000005a2),
    .Q15(NLW_blk000002eb_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002ec (
    .C(clk),
    .CE(ce),
    .D(sig000005a2),
    .Q(sig0000017e)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000002ed (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(a[34]),
    .Q(sig000005a3),
    .Q15(NLW_blk000002ed_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002ee (
    .C(clk),
    .CE(ce),
    .D(sig000005a3),
    .Q(sig0000017f)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000002ef (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(b[14]),
    .Q(sig000005a4),
    .Q15(NLW_blk000002ef_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002f0 (
    .C(clk),
    .CE(ce),
    .D(sig000005a4),
    .Q(sig00000182)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000002f1 (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(b[16]),
    .Q(sig000005a5),
    .Q15(NLW_blk000002f1_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002f2 (
    .C(clk),
    .CE(ce),
    .D(sig000005a5),
    .Q(sig00000180)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000002f3 (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(b[15]),
    .Q(sig000005a6),
    .Q15(NLW_blk000002f3_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002f4 (
    .C(clk),
    .CE(ce),
    .D(sig000005a6),
    .Q(sig00000181)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000002f5 (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(b[13]),
    .Q(sig000005a7),
    .Q15(NLW_blk000002f5_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002f6 (
    .C(clk),
    .CE(ce),
    .D(sig000005a7),
    .Q(sig00000183)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000002f7 (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(b[12]),
    .Q(sig000005a8),
    .Q15(NLW_blk000002f7_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002f8 (
    .C(clk),
    .CE(ce),
    .D(sig000005a8),
    .Q(sig00000184)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000002f9 (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(b[11]),
    .Q(sig000005a9),
    .Q15(NLW_blk000002f9_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002fa (
    .C(clk),
    .CE(ce),
    .D(sig000005a9),
    .Q(sig00000185)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000002fb (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(b[10]),
    .Q(sig000005aa),
    .Q15(NLW_blk000002fb_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002fc (
    .C(clk),
    .CE(ce),
    .D(sig000005aa),
    .Q(sig00000186)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000002fd (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(b[7]),
    .Q(sig000005ab),
    .Q15(NLW_blk000002fd_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002fe (
    .C(clk),
    .CE(ce),
    .D(sig000005ab),
    .Q(sig00000189)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000002ff (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(b[9]),
    .Q(sig000005ac),
    .Q15(NLW_blk000002ff_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000300 (
    .C(clk),
    .CE(ce),
    .D(sig000005ac),
    .Q(sig00000187)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000301 (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(b[8]),
    .Q(sig000005ad),
    .Q15(NLW_blk00000301_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000302 (
    .C(clk),
    .CE(ce),
    .D(sig000005ad),
    .Q(sig00000188)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000303 (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(b[4]),
    .Q(sig000005ae),
    .Q15(NLW_blk00000303_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000304 (
    .C(clk),
    .CE(ce),
    .D(sig000005ae),
    .Q(sig0000018c)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000305 (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(b[6]),
    .Q(sig000005af),
    .Q15(NLW_blk00000305_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000306 (
    .C(clk),
    .CE(ce),
    .D(sig000005af),
    .Q(sig0000018a)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000307 (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(b[5]),
    .Q(sig000005b0),
    .Q15(NLW_blk00000307_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000308 (
    .C(clk),
    .CE(ce),
    .D(sig000005b0),
    .Q(sig0000018b)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000309 (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(b[1]),
    .Q(sig000005b1),
    .Q15(NLW_blk00000309_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000030a (
    .C(clk),
    .CE(ce),
    .D(sig000005b1),
    .Q(sig0000018f)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk0000030b (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(b[3]),
    .Q(sig000005b2),
    .Q15(NLW_blk0000030b_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000030c (
    .C(clk),
    .CE(ce),
    .D(sig000005b2),
    .Q(sig0000018d)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk0000030d (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(b[2]),
    .Q(sig000005b3),
    .Q15(NLW_blk0000030d_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000030e (
    .C(clk),
    .CE(ce),
    .D(sig000005b3),
    .Q(sig0000018e)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk0000030f (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(b[0]),
    .Q(sig000005b4),
    .Q15(NLW_blk0000030f_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000310 (
    .C(clk),
    .CE(ce),
    .D(sig000005b4),
    .Q(sig00000190)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000311 (
    .A0(sig00000461),
    .A1(sig00000001),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(b[51]),
    .Q(sig000005b5),
    .Q15(NLW_blk00000311_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000312 (
    .C(clk),
    .CE(ce),
    .D(sig000005b5),
    .Q(sig0000014a)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000313 (
    .A0(sig00000461),
    .A1(sig00000001),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(b[50]),
    .Q(sig000005b6),
    .Q15(NLW_blk00000313_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000314 (
    .C(clk),
    .CE(ce),
    .D(sig000005b6),
    .Q(sig0000014b)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000315 (
    .A0(sig00000461),
    .A1(sig00000001),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(b[49]),
    .Q(sig000005b7),
    .Q15(NLW_blk00000315_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000316 (
    .C(clk),
    .CE(ce),
    .D(sig000005b7),
    .Q(sig0000014c)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000317 (
    .A0(sig00000461),
    .A1(sig00000001),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(b[46]),
    .Q(sig000005b8),
    .Q15(NLW_blk00000317_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000318 (
    .C(clk),
    .CE(ce),
    .D(sig000005b8),
    .Q(sig0000014f)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000319 (
    .A0(sig00000461),
    .A1(sig00000001),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(b[48]),
    .Q(sig000005b9),
    .Q15(NLW_blk00000319_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000031a (
    .C(clk),
    .CE(ce),
    .D(sig000005b9),
    .Q(sig0000014d)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk0000031b (
    .A0(sig00000461),
    .A1(sig00000001),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(b[47]),
    .Q(sig000005ba),
    .Q15(NLW_blk0000031b_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000031c (
    .C(clk),
    .CE(ce),
    .D(sig000005ba),
    .Q(sig0000014e)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk0000031d (
    .A0(sig00000461),
    .A1(sig00000001),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(b[43]),
    .Q(sig000005bb),
    .Q15(NLW_blk0000031d_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000031e (
    .C(clk),
    .CE(ce),
    .D(sig000005bb),
    .Q(sig00000152)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk0000031f (
    .A0(sig00000461),
    .A1(sig00000001),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(b[45]),
    .Q(sig000005bc),
    .Q15(NLW_blk0000031f_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000320 (
    .C(clk),
    .CE(ce),
    .D(sig000005bc),
    .Q(sig00000150)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000321 (
    .A0(sig00000461),
    .A1(sig00000001),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(b[44]),
    .Q(sig000005bd),
    .Q15(NLW_blk00000321_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000322 (
    .C(clk),
    .CE(ce),
    .D(sig000005bd),
    .Q(sig00000151)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000323 (
    .A0(sig00000461),
    .A1(sig00000001),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(b[40]),
    .Q(sig000005be),
    .Q15(NLW_blk00000323_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000324 (
    .C(clk),
    .CE(ce),
    .D(sig000005be),
    .Q(sig00000155)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000325 (
    .A0(sig00000461),
    .A1(sig00000001),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(b[42]),
    .Q(sig000005bf),
    .Q15(NLW_blk00000325_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000326 (
    .C(clk),
    .CE(ce),
    .D(sig000005bf),
    .Q(sig00000153)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000327 (
    .A0(sig00000461),
    .A1(sig00000001),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(b[41]),
    .Q(sig000005c0),
    .Q15(NLW_blk00000327_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000328 (
    .C(clk),
    .CE(ce),
    .D(sig000005c0),
    .Q(sig00000154)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000329 (
    .A0(sig00000461),
    .A1(sig00000001),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(b[37]),
    .Q(sig000005c1),
    .Q15(NLW_blk00000329_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000032a (
    .C(clk),
    .CE(ce),
    .D(sig000005c1),
    .Q(sig00000158)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk0000032b (
    .A0(sig00000461),
    .A1(sig00000001),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(b[39]),
    .Q(sig000005c2),
    .Q15(NLW_blk0000032b_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000032c (
    .C(clk),
    .CE(ce),
    .D(sig000005c2),
    .Q(sig00000156)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk0000032d (
    .A0(sig00000461),
    .A1(sig00000001),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(b[38]),
    .Q(sig000005c3),
    .Q15(NLW_blk0000032d_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000032e (
    .C(clk),
    .CE(ce),
    .D(sig000005c3),
    .Q(sig00000157)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk0000032f (
    .A0(sig00000461),
    .A1(sig00000001),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(b[34]),
    .Q(sig000005c4),
    .Q15(NLW_blk0000032f_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000330 (
    .C(clk),
    .CE(ce),
    .D(sig000005c4),
    .Q(sig0000015b)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000331 (
    .A0(sig00000461),
    .A1(sig00000001),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(b[36]),
    .Q(sig000005c5),
    .Q15(NLW_blk00000331_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000332 (
    .C(clk),
    .CE(ce),
    .D(sig000005c5),
    .Q(sig00000159)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000333 (
    .A0(sig00000461),
    .A1(sig00000001),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(b[35]),
    .Q(sig000005c6),
    .Q15(NLW_blk00000333_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000334 (
    .C(clk),
    .CE(ce),
    .D(sig000005c6),
    .Q(sig0000015a)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000335 (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig000001a5),
    .Q(sig000005c7),
    .Q15(NLW_blk00000335_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000336 (
    .C(clk),
    .CE(ce),
    .D(sig000005c7),
    .Q(sig0000015e)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000337 (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig000001a3),
    .Q(sig000005c8),
    .Q15(NLW_blk00000337_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000338 (
    .C(clk),
    .CE(ce),
    .D(sig000005c8),
    .Q(sig0000015c)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000339 (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig000001a4),
    .Q(sig000005c9),
    .Q15(NLW_blk00000339_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000033a (
    .C(clk),
    .CE(ce),
    .D(sig000005c9),
    .Q(sig0000015d)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk0000033b (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig000001a8),
    .Q(sig000005ca),
    .Q15(NLW_blk0000033b_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000033c (
    .C(clk),
    .CE(ce),
    .D(sig000005ca),
    .Q(sig00000161)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk0000033d (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig000001a6),
    .Q(sig000005cb),
    .Q15(NLW_blk0000033d_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000033e (
    .C(clk),
    .CE(ce),
    .D(sig000005cb),
    .Q(sig0000015f)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk0000033f (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig000001a7),
    .Q(sig000005cc),
    .Q15(NLW_blk0000033f_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000340 (
    .C(clk),
    .CE(ce),
    .D(sig000005cc),
    .Q(sig00000160)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000341 (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig000001a9),
    .Q(sig000005cd),
    .Q15(NLW_blk00000341_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000342 (
    .C(clk),
    .CE(ce),
    .D(sig000005cd),
    .Q(sig00000162)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000343 (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig000001aa),
    .Q(sig000005ce),
    .Q15(NLW_blk00000343_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000344 (
    .C(clk),
    .CE(ce),
    .D(sig000005ce),
    .Q(sig00000163)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000345 (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig000001ab),
    .Q(sig000005cf),
    .Q15(NLW_blk00000345_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000346 (
    .C(clk),
    .CE(ce),
    .D(sig000005cf),
    .Q(sig00000164)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000347 (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig000001ac),
    .Q(sig000005d0),
    .Q15(NLW_blk00000347_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000348 (
    .C(clk),
    .CE(ce),
    .D(sig000005d0),
    .Q(sig00000165)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000349 (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig000001af),
    .Q(sig000005d1),
    .Q15(NLW_blk00000349_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000034a (
    .C(clk),
    .CE(ce),
    .D(sig000005d1),
    .Q(sig00000168)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk0000034b (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig000001ad),
    .Q(sig000005d2),
    .Q15(NLW_blk0000034b_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000034c (
    .C(clk),
    .CE(ce),
    .D(sig000005d2),
    .Q(sig00000166)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk0000034d (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig000001ae),
    .Q(sig000005d3),
    .Q15(NLW_blk0000034d_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000034e (
    .C(clk),
    .CE(ce),
    .D(sig000005d3),
    .Q(sig00000167)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk0000034f (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig000001b2),
    .Q(sig000005d4),
    .Q15(NLW_blk0000034f_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000350 (
    .C(clk),
    .CE(ce),
    .D(sig000005d4),
    .Q(sig0000016b)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000351 (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig000001b0),
    .Q(sig000005d5),
    .Q15(NLW_blk00000351_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000352 (
    .C(clk),
    .CE(ce),
    .D(sig000005d5),
    .Q(sig00000169)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000353 (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig000001b1),
    .Q(sig000005d6),
    .Q15(NLW_blk00000353_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000354 (
    .C(clk),
    .CE(ce),
    .D(sig000005d6),
    .Q(sig0000016a)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000355 (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig000001b3),
    .Q(sig000005d7),
    .Q15(NLW_blk00000355_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000356 (
    .C(clk),
    .CE(ce),
    .D(sig000005d7),
    .Q(sig0000016c)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000357 (
    .A0(sig00000461),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig00000149),
    .Q(sig000005d8),
    .Q15(NLW_blk00000357_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000358 (
    .C(clk),
    .CE(ce),
    .D(sig000005d8),
    .Q(sig00000113)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000359 (
    .A0(sig00000001),
    .A1(sig00000001),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig000001b4),
    .Q(sig000005d9),
    .Q15(NLW_blk00000359_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000035a (
    .C(clk),
    .CE(ce),
    .D(sig000005d9),
    .Q(sig00000126)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk0000035b (
    .A0(sig00000001),
    .A1(sig00000001),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig000001b7),
    .Q(sig000005da),
    .Q15(NLW_blk0000035b_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000035c (
    .C(clk),
    .CE(ce),
    .D(sig000005da),
    .Q(sig00000129)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk0000035d (
    .A0(sig00000001),
    .A1(sig00000001),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig000001b5),
    .Q(sig000005db),
    .Q15(NLW_blk0000035d_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000035e (
    .C(clk),
    .CE(ce),
    .D(sig000005db),
    .Q(sig00000127)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk0000035f (
    .A0(sig00000001),
    .A1(sig00000001),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig000001b6),
    .Q(sig000005dc),
    .Q15(NLW_blk0000035f_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000360 (
    .C(clk),
    .CE(ce),
    .D(sig000005dc),
    .Q(sig00000128)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000361 (
    .A0(sig00000001),
    .A1(sig00000001),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig000001b8),
    .Q(sig000005dd),
    .Q15(NLW_blk00000361_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000362 (
    .C(clk),
    .CE(ce),
    .D(sig000005dd),
    .Q(sig0000012a)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000363 (
    .A0(sig00000001),
    .A1(sig00000001),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig000001b9),
    .Q(sig000005de),
    .Q15(NLW_blk00000363_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000364 (
    .C(clk),
    .CE(ce),
    .D(sig000005de),
    .Q(sig0000012b)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000365 (
    .A0(sig00000001),
    .A1(sig00000001),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig000001ba),
    .Q(sig000005df),
    .Q15(NLW_blk00000365_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000366 (
    .C(clk),
    .CE(ce),
    .D(sig000005df),
    .Q(sig0000012c)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000367 (
    .A0(sig00000001),
    .A1(sig00000001),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig000001bb),
    .Q(sig000005e0),
    .Q15(NLW_blk00000367_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000368 (
    .C(clk),
    .CE(ce),
    .D(sig000005e0),
    .Q(sig0000012d)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000369 (
    .A0(sig00000001),
    .A1(sig00000001),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig000001be),
    .Q(sig000005e1),
    .Q15(NLW_blk00000369_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000036a (
    .C(clk),
    .CE(ce),
    .D(sig000005e1),
    .Q(sig00000130)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk0000036b (
    .A0(sig00000001),
    .A1(sig00000001),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig000001bc),
    .Q(sig000005e2),
    .Q15(NLW_blk0000036b_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000036c (
    .C(clk),
    .CE(ce),
    .D(sig000005e2),
    .Q(sig0000012e)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk0000036d (
    .A0(sig00000001),
    .A1(sig00000001),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig000001bd),
    .Q(sig000005e3),
    .Q15(NLW_blk0000036d_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000036e (
    .C(clk),
    .CE(ce),
    .D(sig000005e3),
    .Q(sig0000012f)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk0000036f (
    .A0(sig00000001),
    .A1(sig00000001),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig000001c1),
    .Q(sig000005e4),
    .Q15(NLW_blk0000036f_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000370 (
    .C(clk),
    .CE(ce),
    .D(sig000005e4),
    .Q(sig00000133)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000371 (
    .A0(sig00000001),
    .A1(sig00000001),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig000001bf),
    .Q(sig000005e5),
    .Q15(NLW_blk00000371_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000372 (
    .C(clk),
    .CE(ce),
    .D(sig000005e5),
    .Q(sig00000131)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000373 (
    .A0(sig00000001),
    .A1(sig00000001),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig000001c0),
    .Q(sig000005e6),
    .Q15(NLW_blk00000373_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000374 (
    .C(clk),
    .CE(ce),
    .D(sig000005e6),
    .Q(sig00000132)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000375 (
    .A0(sig00000001),
    .A1(sig00000001),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig000001c4),
    .Q(sig000005e7),
    .Q15(NLW_blk00000375_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000376 (
    .C(clk),
    .CE(ce),
    .D(sig000005e7),
    .Q(sig00000136)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000377 (
    .A0(sig00000001),
    .A1(sig00000001),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig000001c2),
    .Q(sig000005e8),
    .Q15(NLW_blk00000377_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000378 (
    .C(clk),
    .CE(ce),
    .D(sig000005e8),
    .Q(sig00000134)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000379 (
    .A0(sig00000001),
    .A1(sig00000001),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig000001c3),
    .Q(sig000005e9),
    .Q15(NLW_blk00000379_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000037a (
    .C(clk),
    .CE(ce),
    .D(sig000005e9),
    .Q(sig00000135)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk0000037b (
    .A0(sig00000001),
    .A1(sig00000001),
    .A2(sig00000461),
    .A3(sig00000001),
    .CE(ce),
    .CLK(clk),
    .D(sig000000b4),
    .Q(sig000005ea),
    .Q15(NLW_blk0000037b_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000037c (
    .C(clk),
    .CE(ce),
    .D(sig000005ea),
    .Q(sig0000047d)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk0000037d (
    .A0(sig00000001),
    .A1(sig00000001),
    .A2(sig00000461),
    .A3(sig00000001),
    .CE(ce),
    .CLK(clk),
    .D(sig000000b1),
    .Q(sig000005eb),
    .Q15(NLW_blk0000037d_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000037e (
    .C(clk),
    .CE(ce),
    .D(sig000005eb),
    .Q(sig00000459)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk0000037f (
    .A0(sig00000001),
    .A1(sig00000001),
    .A2(sig00000461),
    .A3(sig00000001),
    .CE(ce),
    .CLK(clk),
    .D(sig000000b3),
    .Q(sig000005ec),
    .Q15(NLW_blk0000037f_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000380 (
    .C(clk),
    .CE(ce),
    .D(sig000005ec),
    .Q(sig0000045b)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000381 (
    .A0(sig00000001),
    .A1(sig00000001),
    .A2(sig00000461),
    .A3(sig00000001),
    .CE(ce),
    .CLK(clk),
    .D(sig000000b2),
    .Q(sig000005ed),
    .Q15(NLW_blk00000381_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000382 (
    .C(clk),
    .CE(ce),
    .D(sig000005ed),
    .Q(sig0000045a)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000383 (
    .A0(sig00000001),
    .A1(sig00000001),
    .A2(sig00000461),
    .A3(sig00000001),
    .CE(ce),
    .CLK(clk),
    .D(sig000000ae),
    .Q(sig000005ee),
    .Q15(NLW_blk00000383_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000384 (
    .C(clk),
    .CE(ce),
    .D(sig000005ee),
    .Q(sig00000456)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000385 (
    .A0(sig00000001),
    .A1(sig00000001),
    .A2(sig00000461),
    .A3(sig00000001),
    .CE(ce),
    .CLK(clk),
    .D(sig000000b0),
    .Q(sig000005ef),
    .Q15(NLW_blk00000385_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000386 (
    .C(clk),
    .CE(ce),
    .D(sig000005ef),
    .Q(sig00000458)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000387 (
    .A0(sig00000001),
    .A1(sig00000001),
    .A2(sig00000461),
    .A3(sig00000001),
    .CE(ce),
    .CLK(clk),
    .D(sig000000af),
    .Q(sig000005f0),
    .Q15(NLW_blk00000387_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000388 (
    .C(clk),
    .CE(ce),
    .D(sig000005f0),
    .Q(sig00000457)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000389 (
    .A0(sig00000001),
    .A1(sig00000001),
    .A2(sig00000461),
    .A3(sig00000001),
    .CE(ce),
    .CLK(clk),
    .D(sig000000ab),
    .Q(sig000005f1),
    .Q15(NLW_blk00000389_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000038a (
    .C(clk),
    .CE(ce),
    .D(sig000005f1),
    .Q(sig00000453)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk0000038b (
    .A0(sig00000001),
    .A1(sig00000001),
    .A2(sig00000461),
    .A3(sig00000001),
    .CE(ce),
    .CLK(clk),
    .D(sig000000ad),
    .Q(sig000005f2),
    .Q15(NLW_blk0000038b_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000038c (
    .C(clk),
    .CE(ce),
    .D(sig000005f2),
    .Q(sig00000455)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk0000038d (
    .A0(sig00000001),
    .A1(sig00000001),
    .A2(sig00000461),
    .A3(sig00000001),
    .CE(ce),
    .CLK(clk),
    .D(sig000000ac),
    .Q(sig000005f3),
    .Q15(NLW_blk0000038d_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000038e (
    .C(clk),
    .CE(ce),
    .D(sig000005f3),
    .Q(sig00000454)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk0000038f (
    .A0(sig00000461),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig000001d6),
    .Q(sig000005f4),
    .Q15(NLW_blk0000038f_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000390 (
    .C(clk),
    .CE(ce),
    .D(sig000005f4),
    .Q(sig00000467)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000391 (
    .A0(sig00000001),
    .A1(sig00000001),
    .A2(sig00000461),
    .A3(sig00000001),
    .CE(ce),
    .CLK(clk),
    .D(sig000000aa),
    .Q(sig000005f5),
    .Q15(NLW_blk00000391_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000392 (
    .C(clk),
    .CE(ce),
    .D(sig000005f5),
    .Q(sig00000452)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000393 (
    .A0(sig00000461),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig000001d7),
    .Q(sig000005f6),
    .Q15(NLW_blk00000393_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000394 (
    .C(clk),
    .CE(ce),
    .D(sig000005f6),
    .Q(sig00000468)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000395 (
    .A0(sig00000461),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig000001d3),
    .Q(sig000005f7),
    .Q15(NLW_blk00000395_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000396 (
    .C(clk),
    .CE(ce),
    .D(sig000005f7),
    .Q(sig00000464)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000397 (
    .A0(sig00000461),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig000001d5),
    .Q(sig000005f8),
    .Q15(NLW_blk00000397_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000398 (
    .C(clk),
    .CE(ce),
    .D(sig000005f8),
    .Q(sig00000466)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000399 (
    .A0(sig00000461),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig000001d4),
    .Q(sig000005f9),
    .Q15(NLW_blk00000399_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000039a (
    .C(clk),
    .CE(ce),
    .D(sig000005f9),
    .Q(sig00000465)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk0000039b (
    .A0(sig00000461),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig0000007f),
    .Q(sig000005fa),
    .Q15(NLW_blk0000039b_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000039c (
    .C(clk),
    .CE(ce),
    .D(sig000005fa),
    .Q(\U0/op_inst/FLT_PT_OP/MULT.OP/OP/sign_op )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk0000039d (
    .A0(sig00000461),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig000001d2),
    .Q(sig000005fb),
    .Q15(NLW_blk0000039d_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000039e (
    .C(clk),
    .CE(ce),
    .D(sig000005fb),
    .Q(sig00000463)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk0000039f (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig00000192),
    .Q(sig000005fc),
    .Q15(NLW_blk0000039f_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003a0 (
    .C(clk),
    .CE(ce),
    .D(sig000005fc),
    .Q(sig00000138)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000003a1 (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig00000191),
    .Q(sig000005fd),
    .Q15(NLW_blk000003a1_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003a2 (
    .C(clk),
    .CE(ce),
    .D(sig000005fd),
    .Q(sig00000137)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000003a3 (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig00000193),
    .Q(sig000005fe),
    .Q15(NLW_blk000003a3_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003a4 (
    .C(clk),
    .CE(ce),
    .D(sig000005fe),
    .Q(sig00000139)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000003a5 (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig00000194),
    .Q(sig000005ff),
    .Q15(NLW_blk000003a5_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003a6 (
    .C(clk),
    .CE(ce),
    .D(sig000005ff),
    .Q(sig0000013a)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000003a7 (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig00000195),
    .Q(sig00000600),
    .Q15(NLW_blk000003a7_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003a8 (
    .C(clk),
    .CE(ce),
    .D(sig00000600),
    .Q(sig0000013b)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000003a9 (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig00000196),
    .Q(sig00000601),
    .Q15(NLW_blk000003a9_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003aa (
    .C(clk),
    .CE(ce),
    .D(sig00000601),
    .Q(sig0000013c)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000003ab (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig00000199),
    .Q(sig00000602),
    .Q15(NLW_blk000003ab_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003ac (
    .C(clk),
    .CE(ce),
    .D(sig00000602),
    .Q(sig0000013f)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000003ad (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig00000197),
    .Q(sig00000603),
    .Q15(NLW_blk000003ad_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003ae (
    .C(clk),
    .CE(ce),
    .D(sig00000603),
    .Q(sig0000013d)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000003af (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig00000198),
    .Q(sig00000604),
    .Q15(NLW_blk000003af_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003b0 (
    .C(clk),
    .CE(ce),
    .D(sig00000604),
    .Q(sig0000013e)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000003b1 (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig0000019c),
    .Q(sig00000605),
    .Q15(NLW_blk000003b1_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003b2 (
    .C(clk),
    .CE(ce),
    .D(sig00000605),
    .Q(sig00000142)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000003b3 (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig0000019a),
    .Q(sig00000606),
    .Q15(NLW_blk000003b3_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003b4 (
    .C(clk),
    .CE(ce),
    .D(sig00000606),
    .Q(sig00000140)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000003b5 (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig0000019b),
    .Q(sig00000607),
    .Q15(NLW_blk000003b5_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003b6 (
    .C(clk),
    .CE(ce),
    .D(sig00000607),
    .Q(sig00000141)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000003b7 (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig0000019f),
    .Q(sig00000608),
    .Q15(NLW_blk000003b7_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003b8 (
    .C(clk),
    .CE(ce),
    .D(sig00000608),
    .Q(sig00000145)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000003b9 (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig0000019d),
    .Q(sig00000609),
    .Q15(NLW_blk000003b9_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003ba (
    .C(clk),
    .CE(ce),
    .D(sig00000609),
    .Q(sig00000143)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000003bb (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig0000019e),
    .Q(sig0000060a),
    .Q15(NLW_blk000003bb_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003bc (
    .C(clk),
    .CE(ce),
    .D(sig0000060a),
    .Q(sig00000144)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000003bd (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig000001a0),
    .Q(sig0000060b),
    .Q15(NLW_blk000003bd_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003be (
    .C(clk),
    .CE(ce),
    .D(sig0000060b),
    .Q(sig00000146)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000003bf (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig000001a1),
    .Q(sig0000060c),
    .Q15(NLW_blk000003bf_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003c0 (
    .C(clk),
    .CE(ce),
    .D(sig0000060c),
    .Q(sig00000147)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000003c1 (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig0000016e),
    .Q(sig0000060d),
    .Q15(NLW_blk000003c1_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003c2 (
    .C(clk),
    .CE(ce),
    .D(sig0000060d),
    .Q(sig00000114)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000003c3 (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig00000171),
    .Q(sig0000060e),
    .Q15(NLW_blk000003c3_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003c4 (
    .C(clk),
    .CE(ce),
    .D(sig0000060e),
    .Q(sig00000117)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000003c5 (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig0000016f),
    .Q(sig0000060f),
    .Q15(NLW_blk000003c5_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003c6 (
    .C(clk),
    .CE(ce),
    .D(sig0000060f),
    .Q(sig00000115)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000003c7 (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig00000170),
    .Q(sig00000610),
    .Q15(NLW_blk000003c7_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003c8 (
    .C(clk),
    .CE(ce),
    .D(sig00000610),
    .Q(sig00000116)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000003c9 (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig00000174),
    .Q(sig00000611),
    .Q15(NLW_blk000003c9_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003ca (
    .C(clk),
    .CE(ce),
    .D(sig00000611),
    .Q(sig0000011a)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000003cb (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig00000172),
    .Q(sig00000612),
    .Q15(NLW_blk000003cb_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003cc (
    .C(clk),
    .CE(ce),
    .D(sig00000612),
    .Q(sig00000118)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000003cd (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig00000173),
    .Q(sig00000613),
    .Q15(NLW_blk000003cd_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003ce (
    .C(clk),
    .CE(ce),
    .D(sig00000613),
    .Q(sig00000119)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000003cf (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig00000177),
    .Q(sig00000614),
    .Q15(NLW_blk000003cf_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003d0 (
    .C(clk),
    .CE(ce),
    .D(sig00000614),
    .Q(sig0000011d)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000003d1 (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig00000175),
    .Q(sig00000615),
    .Q15(NLW_blk000003d1_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003d2 (
    .C(clk),
    .CE(ce),
    .D(sig00000615),
    .Q(sig0000011b)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000003d3 (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig00000176),
    .Q(sig00000616),
    .Q15(NLW_blk000003d3_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003d4 (
    .C(clk),
    .CE(ce),
    .D(sig00000616),
    .Q(sig0000011c)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000003d5 (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig0000017a),
    .Q(sig00000617),
    .Q15(NLW_blk000003d5_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003d6 (
    .C(clk),
    .CE(ce),
    .D(sig00000617),
    .Q(sig00000120)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000003d7 (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig00000178),
    .Q(sig00000618),
    .Q15(NLW_blk000003d7_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003d8 (
    .C(clk),
    .CE(ce),
    .D(sig00000618),
    .Q(sig0000011e)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000003d9 (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig00000179),
    .Q(sig00000619),
    .Q15(NLW_blk000003d9_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003da (
    .C(clk),
    .CE(ce),
    .D(sig00000619),
    .Q(sig0000011f)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000003db (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig0000017d),
    .Q(sig0000061a),
    .Q15(NLW_blk000003db_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003dc (
    .C(clk),
    .CE(ce),
    .D(sig0000061a),
    .Q(sig00000123)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000003dd (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig0000017b),
    .Q(sig0000061b),
    .Q15(NLW_blk000003dd_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003de (
    .C(clk),
    .CE(ce),
    .D(sig0000061b),
    .Q(sig00000121)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000003df (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig0000017c),
    .Q(sig0000061c),
    .Q15(NLW_blk000003df_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003e0 (
    .C(clk),
    .CE(ce),
    .D(sig0000061c),
    .Q(sig00000122)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000003e1 (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig0000017e),
    .Q(sig0000061d),
    .Q15(NLW_blk000003e1_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003e2 (
    .C(clk),
    .CE(ce),
    .D(sig0000061d),
    .Q(sig00000124)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000003e3 (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig0000017f),
    .Q(sig0000061e),
    .Q15(NLW_blk000003e3_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003e4 (
    .C(clk),
    .CE(ce),
    .D(sig0000061e),
    .Q(sig00000125)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000003e5 (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig0000014b),
    .Q(sig0000061f),
    .Q15(NLW_blk000003e5_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003e6 (
    .C(clk),
    .CE(ce),
    .D(sig0000061f),
    .Q(sig00000102)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000003e7 (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig0000014c),
    .Q(sig00000620),
    .Q15(NLW_blk000003e7_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003e8 (
    .C(clk),
    .CE(ce),
    .D(sig00000620),
    .Q(sig00000103)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000003e9 (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig0000014d),
    .Q(sig00000621),
    .Q15(NLW_blk000003e9_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003ea (
    .C(clk),
    .CE(ce),
    .D(sig00000621),
    .Q(sig00000104)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000003eb (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig0000014e),
    .Q(sig00000622),
    .Q15(NLW_blk000003eb_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003ec (
    .C(clk),
    .CE(ce),
    .D(sig00000622),
    .Q(sig00000105)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000003ed (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig00000151),
    .Q(sig00000623),
    .Q15(NLW_blk000003ed_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003ee (
    .C(clk),
    .CE(ce),
    .D(sig00000623),
    .Q(sig00000108)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000003ef (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig0000014f),
    .Q(sig00000624),
    .Q15(NLW_blk000003ef_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003f0 (
    .C(clk),
    .CE(ce),
    .D(sig00000624),
    .Q(sig00000106)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000003f1 (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig00000150),
    .Q(sig00000625),
    .Q15(NLW_blk000003f1_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003f2 (
    .C(clk),
    .CE(ce),
    .D(sig00000625),
    .Q(sig00000107)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000003f3 (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig00000154),
    .Q(sig00000626),
    .Q15(NLW_blk000003f3_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003f4 (
    .C(clk),
    .CE(ce),
    .D(sig00000626),
    .Q(sig0000010b)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000003f5 (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig00000152),
    .Q(sig00000627),
    .Q15(NLW_blk000003f5_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003f6 (
    .C(clk),
    .CE(ce),
    .D(sig00000627),
    .Q(sig00000109)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000003f7 (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig00000153),
    .Q(sig00000628),
    .Q15(NLW_blk000003f7_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003f8 (
    .C(clk),
    .CE(ce),
    .D(sig00000628),
    .Q(sig0000010a)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000003f9 (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig00000157),
    .Q(sig00000629),
    .Q15(NLW_blk000003f9_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003fa (
    .C(clk),
    .CE(ce),
    .D(sig00000629),
    .Q(sig0000010e)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000003fb (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig00000155),
    .Q(sig0000062a),
    .Q15(NLW_blk000003fb_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003fc (
    .C(clk),
    .CE(ce),
    .D(sig0000062a),
    .Q(sig0000010c)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000003fd (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig00000156),
    .Q(sig0000062b),
    .Q15(NLW_blk000003fd_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003fe (
    .C(clk),
    .CE(ce),
    .D(sig0000062b),
    .Q(sig0000010d)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000003ff (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig00000158),
    .Q(sig0000062c),
    .Q15(NLW_blk000003ff_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000400 (
    .C(clk),
    .CE(ce),
    .D(sig0000062c),
    .Q(sig0000010f)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000401 (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig00000159),
    .Q(sig0000062d),
    .Q15(NLW_blk00000401_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000402 (
    .C(clk),
    .CE(ce),
    .D(sig0000062d),
    .Q(sig00000110)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000403 (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig0000015a),
    .Q(sig0000062e),
    .Q15(NLW_blk00000403_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000404 (
    .C(clk),
    .CE(ce),
    .D(sig0000062e),
    .Q(sig00000111)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000405 (
    .A0(sig00000001),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig0000015b),
    .Q(sig0000062f),
    .Q15(NLW_blk00000405_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000406 (
    .C(clk),
    .CE(ce),
    .D(sig0000062f),
    .Q(sig00000112)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000407 (
    .A0(sig00000461),
    .A1(sig00000461),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig00000113),
    .Q(sig00000630),
    .Q15(NLW_blk00000407_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000408 (
    .C(clk),
    .CE(ce),
    .D(sig00000630),
    .Q(sig00000100)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000409 (
    .A0(sig00000461),
    .A1(sig00000001),
    .A2(sig00000461),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig0000014a),
    .Q(sig00000631),
    .Q15(NLW_blk00000409_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000040a (
    .C(clk),
    .CE(ce),
    .D(sig00000631),
    .Q(sig00000101)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk0000040b (
    .A0(sig00000461),
    .A1(sig00000461),
    .A2(sig00000001),
    .A3(sig00000461),
    .CE(ce),
    .CLK(clk),
    .D(sig00000100),
    .Q(sig00000632),
    .Q15(NLW_blk0000040b_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000040c (
    .C(clk),
    .CE(ce),
    .D(sig00000632),
    .Q(sig00000551)
  );
  DSP48E #(
    .ACASCREG ( 1 ),
    .ALUMODEREG ( 0 ),
    .AREG ( 1 ),
    .AUTORESET_PATTERN_DETECT ( "FALSE" ),
    .AUTORESET_PATTERN_DETECT_OPTINV ( "MATCH" ),
    .A_INPUT ( "CASCADE" ),
    .BCASCREG ( 2 ),
    .BREG ( 2 ),
    .B_INPUT ( "DIRECT" ),
    .CARRYINREG ( 0 ),
    .CARRYINSELREG ( 0 ),
    .CREG ( 0 ),
    .MASK ( 48'h3FFFFFFFFFFF ),
    .MREG ( 1 ),
    .MULTCARRYINREG ( 0 ),
    .OPMODEREG ( 0 ),
    .PATTERN ( 48'h000000000000 ),
    .PREG ( 1 ),
    .SEL_MASK ( "MASK" ),
    .SEL_PATTERN ( "PATTERN" ),
    .SEL_ROUNDING_MASK ( "SEL_MASK" ),
    .SIM_MODE ( "SAFE" ),
    .USE_MULT ( "MULT_S" ),
    .USE_PATTERN_DETECT ( "NO_PATDET" ),
    .USE_SIMD ( "ONE48" ))
  blk0000040d (
    .CEM(ce),
    .CLK(clk),
    .PATTERNBDETECT(NLW_blk0000040d_PATTERNBDETECT_UNCONNECTED),
    .RSTC(sig00000461),
    .CEB1(ce),
    .MULTSIGNOUT(NLW_blk0000040d_MULTSIGNOUT_UNCONNECTED),
    .CEC(sig00000461),
    .RSTM(sig00000461),
    .MULTSIGNIN(sig00000461),
    .CEB2(ce),
    .RSTCTRL(sig00000461),
    .CEP(ce),
    .CARRYCASCOUT(NLW_blk0000040d_CARRYCASCOUT_UNCONNECTED),
    .RSTA(sig00000461),
    .CECARRYIN(sig00000461),
    .UNDERFLOW(NLW_blk0000040d_UNDERFLOW_UNCONNECTED),
    .PATTERNDETECT(NLW_blk0000040d_PATTERNDETECT_UNCONNECTED),
    .RSTALUMODE(sig00000461),
    .RSTALLCARRYIN(sig00000461),
    .CEALUMODE(sig00000461),
    .CEA2(ce),
    .CEA1(sig00000461),
    .RSTB(sig00000461),
    .CEMULTCARRYIN(sig00000461),
    .OVERFLOW(NLW_blk0000040d_OVERFLOW_UNCONNECTED),
    .CECTRL(sig00000461),
    .CARRYIN(sig00000461),
    .CARRYCASCIN(sig00000461),
    .RSTP(sig00000461),
    .CARRYINSEL({sig00000461, sig00000461, sig00000461}),
    .OPMODE({sig00000001, sig00000461, sig00000001, sig00000461, sig00000001, sig00000461, sig00000001}),
    .PCIN({sig00000207, sig00000206, sig00000205, sig00000204, sig00000203, sig00000202, sig00000201, sig00000200, sig000001ff, sig000001fe,
sig000001fd, sig000001fc, sig000001fb, sig000001fa, sig000001f9, sig000001f8, sig000001f7, sig000001f6, sig000001f5, sig000001f4, sig000001f3,
sig000001f2, sig000001f1, sig000001f0, sig000001ef, sig000001ee, sig000001ed, sig000001ec, sig000001eb, sig000001ea, sig000001e9, sig000001e8,
sig000001e7, sig000001e6, sig000001e5, sig000001e4, sig000001e3, sig000001e2, sig000001e1, sig000001e0, sig000001df, sig000001de, sig000001dd,
sig000001dc, sig000001db, sig000001da, sig000001d9, sig000001d8}),
    .B({sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461
, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000100, sig00000101}),
    .P({\NLW_blk0000040d_P<47>_UNCONNECTED , \NLW_blk0000040d_P<46>_UNCONNECTED , \NLW_blk0000040d_P<45>_UNCONNECTED ,
\NLW_blk0000040d_P<44>_UNCONNECTED , \NLW_blk0000040d_P<43>_UNCONNECTED , \NLW_blk0000040d_P<42>_UNCONNECTED , \NLW_blk0000040d_P<41>_UNCONNECTED ,
\NLW_blk0000040d_P<40>_UNCONNECTED , \NLW_blk0000040d_P<39>_UNCONNECTED , \NLW_blk0000040d_P<38>_UNCONNECTED , \NLW_blk0000040d_P<37>_UNCONNECTED ,
\NLW_blk0000040d_P<36>_UNCONNECTED , \NLW_blk0000040d_P<35>_UNCONNECTED , \NLW_blk0000040d_P<34>_UNCONNECTED , \NLW_blk0000040d_P<33>_UNCONNECTED ,
\NLW_blk0000040d_P<32>_UNCONNECTED , \NLW_blk0000040d_P<31>_UNCONNECTED , \NLW_blk0000040d_P<30>_UNCONNECTED , \NLW_blk0000040d_P<29>_UNCONNECTED ,
\NLW_blk0000040d_P<28>_UNCONNECTED , \NLW_blk0000040d_P<27>_UNCONNECTED , \NLW_blk0000040d_P<26>_UNCONNECTED , \NLW_blk0000040d_P<25>_UNCONNECTED ,
\NLW_blk0000040d_P<24>_UNCONNECTED , \NLW_blk0000040d_P<23>_UNCONNECTED , \NLW_blk0000040d_P<22>_UNCONNECTED , \NLW_blk0000040d_P<21>_UNCONNECTED ,
sig00000008, sig00000009, sig0000000a, sig0000000b, sig0000000c, sig0000000d, sig0000000e, sig0000000f, sig00000010, sig00000011, sig00000012,
sig00000013, sig00000014, sig00000015, sig00000016, sig00000017, sig00000018, sig00000019, sig0000001a, sig0000001b, sig0000001c}),
    .PCOUT({\NLW_blk0000040d_PCOUT<47>_UNCONNECTED , \NLW_blk0000040d_PCOUT<46>_UNCONNECTED , \NLW_blk0000040d_PCOUT<45>_UNCONNECTED ,
\NLW_blk0000040d_PCOUT<44>_UNCONNECTED , \NLW_blk0000040d_PCOUT<43>_UNCONNECTED , \NLW_blk0000040d_PCOUT<42>_UNCONNECTED ,
\NLW_blk0000040d_PCOUT<41>_UNCONNECTED , \NLW_blk0000040d_PCOUT<40>_UNCONNECTED , \NLW_blk0000040d_PCOUT<39>_UNCONNECTED ,
\NLW_blk0000040d_PCOUT<38>_UNCONNECTED , \NLW_blk0000040d_PCOUT<37>_UNCONNECTED , \NLW_blk0000040d_PCOUT<36>_UNCONNECTED ,
\NLW_blk0000040d_PCOUT<35>_UNCONNECTED , \NLW_blk0000040d_PCOUT<34>_UNCONNECTED , \NLW_blk0000040d_PCOUT<33>_UNCONNECTED ,
\NLW_blk0000040d_PCOUT<32>_UNCONNECTED , \NLW_blk0000040d_PCOUT<31>_UNCONNECTED , \NLW_blk0000040d_PCOUT<30>_UNCONNECTED ,
\NLW_blk0000040d_PCOUT<29>_UNCONNECTED , \NLW_blk0000040d_PCOUT<28>_UNCONNECTED , \NLW_blk0000040d_PCOUT<27>_UNCONNECTED ,
\NLW_blk0000040d_PCOUT<26>_UNCONNECTED , \NLW_blk0000040d_PCOUT<25>_UNCONNECTED , \NLW_blk0000040d_PCOUT<24>_UNCONNECTED ,
\NLW_blk0000040d_PCOUT<23>_UNCONNECTED , \NLW_blk0000040d_PCOUT<22>_UNCONNECTED , \NLW_blk0000040d_PCOUT<21>_UNCONNECTED ,
\NLW_blk0000040d_PCOUT<20>_UNCONNECTED , \NLW_blk0000040d_PCOUT<19>_UNCONNECTED , \NLW_blk0000040d_PCOUT<18>_UNCONNECTED ,
\NLW_blk0000040d_PCOUT<17>_UNCONNECTED , \NLW_blk0000040d_PCOUT<16>_UNCONNECTED , \NLW_blk0000040d_PCOUT<15>_UNCONNECTED ,
\NLW_blk0000040d_PCOUT<14>_UNCONNECTED , \NLW_blk0000040d_PCOUT<13>_UNCONNECTED , \NLW_blk0000040d_PCOUT<12>_UNCONNECTED ,
\NLW_blk0000040d_PCOUT<11>_UNCONNECTED , \NLW_blk0000040d_PCOUT<10>_UNCONNECTED , \NLW_blk0000040d_PCOUT<9>_UNCONNECTED ,
\NLW_blk0000040d_PCOUT<8>_UNCONNECTED , \NLW_blk0000040d_PCOUT<7>_UNCONNECTED , \NLW_blk0000040d_PCOUT<6>_UNCONNECTED ,
\NLW_blk0000040d_PCOUT<5>_UNCONNECTED , \NLW_blk0000040d_PCOUT<4>_UNCONNECTED , \NLW_blk0000040d_PCOUT<3>_UNCONNECTED ,
\NLW_blk0000040d_PCOUT<2>_UNCONNECTED , \NLW_blk0000040d_PCOUT<1>_UNCONNECTED , \NLW_blk0000040d_PCOUT<0>_UNCONNECTED }),
    .ACIN({sig00000225, sig00000224, sig00000223, sig00000222, sig00000221, sig00000220, sig0000021f, sig0000021e, sig0000021d, sig0000021c,
sig0000021b, sig0000021a, sig00000219, sig00000218, sig00000217, sig00000216, sig00000215, sig00000214, sig00000213, sig00000212, sig00000211,
sig00000210, sig0000020f, sig0000020e, sig0000020d, sig0000020c, sig0000020b, sig0000020a, sig00000209, sig00000208}),
    .ACOUT({\NLW_blk0000040d_ACOUT<29>_UNCONNECTED , \NLW_blk0000040d_ACOUT<28>_UNCONNECTED , \NLW_blk0000040d_ACOUT<27>_UNCONNECTED ,
\NLW_blk0000040d_ACOUT<26>_UNCONNECTED , \NLW_blk0000040d_ACOUT<25>_UNCONNECTED , \NLW_blk0000040d_ACOUT<24>_UNCONNECTED ,
\NLW_blk0000040d_ACOUT<23>_UNCONNECTED , \NLW_blk0000040d_ACOUT<22>_UNCONNECTED , \NLW_blk0000040d_ACOUT<21>_UNCONNECTED ,
\NLW_blk0000040d_ACOUT<20>_UNCONNECTED , \NLW_blk0000040d_ACOUT<19>_UNCONNECTED , \NLW_blk0000040d_ACOUT<18>_UNCONNECTED ,
\NLW_blk0000040d_ACOUT<17>_UNCONNECTED , \NLW_blk0000040d_ACOUT<16>_UNCONNECTED , \NLW_blk0000040d_ACOUT<15>_UNCONNECTED ,
\NLW_blk0000040d_ACOUT<14>_UNCONNECTED , \NLW_blk0000040d_ACOUT<13>_UNCONNECTED , \NLW_blk0000040d_ACOUT<12>_UNCONNECTED ,
\NLW_blk0000040d_ACOUT<11>_UNCONNECTED , \NLW_blk0000040d_ACOUT<10>_UNCONNECTED , \NLW_blk0000040d_ACOUT<9>_UNCONNECTED ,
\NLW_blk0000040d_ACOUT<8>_UNCONNECTED , \NLW_blk0000040d_ACOUT<7>_UNCONNECTED , \NLW_blk0000040d_ACOUT<6>_UNCONNECTED ,
\NLW_blk0000040d_ACOUT<5>_UNCONNECTED , \NLW_blk0000040d_ACOUT<4>_UNCONNECTED , \NLW_blk0000040d_ACOUT<3>_UNCONNECTED ,
\NLW_blk0000040d_ACOUT<2>_UNCONNECTED , \NLW_blk0000040d_ACOUT<1>_UNCONNECTED , \NLW_blk0000040d_ACOUT<0>_UNCONNECTED }),
    .ALUMODE({sig00000461, sig00000461, sig00000461, sig00000461}),
    .C({sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461
, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461,
sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461,
sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461,
sig00000461, sig00000461, sig00000461, sig00000461}),
    .CARRYOUT({\NLW_blk0000040d_CARRYOUT<3>_UNCONNECTED , \NLW_blk0000040d_CARRYOUT<2>_UNCONNECTED , \NLW_blk0000040d_CARRYOUT<1>_UNCONNECTED ,
\NLW_blk0000040d_CARRYOUT<0>_UNCONNECTED }),
    .BCIN({sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461,
sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461}),
    .BCOUT({\NLW_blk0000040d_BCOUT<17>_UNCONNECTED , \NLW_blk0000040d_BCOUT<16>_UNCONNECTED , \NLW_blk0000040d_BCOUT<15>_UNCONNECTED ,
\NLW_blk0000040d_BCOUT<14>_UNCONNECTED , \NLW_blk0000040d_BCOUT<13>_UNCONNECTED , \NLW_blk0000040d_BCOUT<12>_UNCONNECTED ,
\NLW_blk0000040d_BCOUT<11>_UNCONNECTED , \NLW_blk0000040d_BCOUT<10>_UNCONNECTED , \NLW_blk0000040d_BCOUT<9>_UNCONNECTED ,
\NLW_blk0000040d_BCOUT<8>_UNCONNECTED , \NLW_blk0000040d_BCOUT<7>_UNCONNECTED , \NLW_blk0000040d_BCOUT<6>_UNCONNECTED ,
\NLW_blk0000040d_BCOUT<5>_UNCONNECTED , \NLW_blk0000040d_BCOUT<4>_UNCONNECTED , \NLW_blk0000040d_BCOUT<3>_UNCONNECTED ,
\NLW_blk0000040d_BCOUT<2>_UNCONNECTED , \NLW_blk0000040d_BCOUT<1>_UNCONNECTED , \NLW_blk0000040d_BCOUT<0>_UNCONNECTED }),
    .A({sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461
, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461,
sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461})
  );
  DSP48E #(
    .ACASCREG ( 1 ),
    .ALUMODEREG ( 0 ),
    .AREG ( 1 ),
    .AUTORESET_PATTERN_DETECT ( "FALSE" ),
    .AUTORESET_PATTERN_DETECT_OPTINV ( "MATCH" ),
    .A_INPUT ( "CASCADE" ),
    .BCASCREG ( 2 ),
    .BREG ( 2 ),
    .B_INPUT ( "DIRECT" ),
    .CARRYINREG ( 0 ),
    .CARRYINSELREG ( 0 ),
    .CREG ( 0 ),
    .MASK ( 48'h3FFFFFFFFFFF ),
    .MREG ( 1 ),
    .MULTCARRYINREG ( 0 ),
    .OPMODEREG ( 0 ),
    .PATTERN ( 48'h000000000000 ),
    .PREG ( 1 ),
    .SEL_MASK ( "MASK" ),
    .SEL_PATTERN ( "PATTERN" ),
    .SEL_ROUNDING_MASK ( "SEL_MASK" ),
    .SIM_MODE ( "SAFE" ),
    .USE_MULT ( "MULT_S" ),
    .USE_PATTERN_DETECT ( "NO_PATDET" ),
    .USE_SIMD ( "ONE48" ))
  blk0000040e (
    .CEM(ce),
    .CLK(clk),
    .PATTERNBDETECT(NLW_blk0000040e_PATTERNBDETECT_UNCONNECTED),
    .RSTC(sig00000461),
    .CEB1(ce),
    .MULTSIGNOUT(NLW_blk0000040e_MULTSIGNOUT_UNCONNECTED),
    .CEC(sig00000461),
    .RSTM(sig00000461),
    .MULTSIGNIN(sig00000461),
    .CEB2(ce),
    .RSTCTRL(sig00000461),
    .CEP(ce),
    .CARRYCASCOUT(NLW_blk0000040e_CARRYCASCOUT_UNCONNECTED),
    .RSTA(sig00000461),
    .CECARRYIN(sig00000461),
    .UNDERFLOW(NLW_blk0000040e_UNDERFLOW_UNCONNECTED),
    .PATTERNDETECT(NLW_blk0000040e_PATTERNDETECT_UNCONNECTED),
    .RSTALUMODE(sig00000461),
    .RSTALLCARRYIN(sig00000461),
    .CEALUMODE(sig00000461),
    .CEA2(ce),
    .CEA1(sig00000461),
    .RSTB(sig00000461),
    .CEMULTCARRYIN(sig00000461),
    .OVERFLOW(NLW_blk0000040e_OVERFLOW_UNCONNECTED),
    .CECTRL(sig00000461),
    .CARRYIN(sig00000461),
    .CARRYCASCIN(sig00000461),
    .RSTP(sig00000461),
    .CARRYINSEL({sig00000461, sig00000461, sig00000461}),
    .ACOUT({sig00000225, sig00000224, sig00000223, sig00000222, sig00000221, sig00000220, sig0000021f, sig0000021e, sig0000021d, sig0000021c,
sig0000021b, sig0000021a, sig00000219, sig00000218, sig00000217, sig00000216, sig00000215, sig00000214, sig00000213, sig00000212, sig00000211,
sig00000210, sig0000020f, sig0000020e, sig0000020d, sig0000020c, sig0000020b, sig0000020a, sig00000209, sig00000208}),
    .OPMODE({sig00000001, sig00000461, sig00000001, sig00000461, sig00000001, sig00000461, sig00000001}),
    .PCIN({sig00000266, sig00000265, sig00000264, sig00000263, sig00000262, sig00000261, sig00000260, sig0000025f, sig0000025e, sig0000025d,
sig0000025c, sig0000025b, sig0000025a, sig00000259, sig00000258, sig00000257, sig00000256, sig00000255, sig00000254, sig00000253, sig00000252,
sig00000251, sig00000250, sig0000024f, sig0000024e, sig0000024d, sig0000024c, sig0000024b, sig0000024a, sig00000249, sig00000248, sig00000247,
sig00000246, sig00000245, sig00000244, sig00000243, sig00000242, sig00000241, sig00000240, sig0000023f, sig0000023e, sig0000023d, sig0000023c,
sig0000023b, sig0000023a, sig00000239, sig00000238, sig00000237}),
    .B({sig00000461, sig00000102, sig00000103, sig00000104, sig00000105, sig00000106, sig00000107, sig00000108, sig00000109, sig0000010a, sig0000010b
, sig0000010c, sig0000010d, sig0000010e, sig0000010f, sig00000110, sig00000111, sig00000112}),
    .P({\NLW_blk0000040e_P<47>_UNCONNECTED , \NLW_blk0000040e_P<46>_UNCONNECTED , \NLW_blk0000040e_P<45>_UNCONNECTED ,
\NLW_blk0000040e_P<44>_UNCONNECTED , \NLW_blk0000040e_P<43>_UNCONNECTED , \NLW_blk0000040e_P<42>_UNCONNECTED , \NLW_blk0000040e_P<41>_UNCONNECTED ,
\NLW_blk0000040e_P<40>_UNCONNECTED , \NLW_blk0000040e_P<39>_UNCONNECTED , \NLW_blk0000040e_P<38>_UNCONNECTED , \NLW_blk0000040e_P<37>_UNCONNECTED ,
\NLW_blk0000040e_P<36>_UNCONNECTED , \NLW_blk0000040e_P<35>_UNCONNECTED , \NLW_blk0000040e_P<34>_UNCONNECTED , \NLW_blk0000040e_P<33>_UNCONNECTED ,
\NLW_blk0000040e_P<32>_UNCONNECTED , \NLW_blk0000040e_P<31>_UNCONNECTED , \NLW_blk0000040e_P<30>_UNCONNECTED , \NLW_blk0000040e_P<29>_UNCONNECTED ,
\NLW_blk0000040e_P<28>_UNCONNECTED , \NLW_blk0000040e_P<27>_UNCONNECTED , \NLW_blk0000040e_P<26>_UNCONNECTED , \NLW_blk0000040e_P<25>_UNCONNECTED ,
\NLW_blk0000040e_P<24>_UNCONNECTED , \NLW_blk0000040e_P<23>_UNCONNECTED , \NLW_blk0000040e_P<22>_UNCONNECTED , \NLW_blk0000040e_P<21>_UNCONNECTED ,
\NLW_blk0000040e_P<20>_UNCONNECTED , \NLW_blk0000040e_P<19>_UNCONNECTED , \NLW_blk0000040e_P<18>_UNCONNECTED , \NLW_blk0000040e_P<17>_UNCONNECTED ,
sig000001d7, sig000001d6, sig000001d5, sig000001d4, sig000001d3, sig000001d2, sig000001d1, sig000001d0, sig000001cf, sig000001ce, sig000001cd,
sig000001cc, sig000001cb, sig000001ca, sig000001c9, sig000001c8, sig000001c7}),
    .PCOUT({sig00000207, sig00000206, sig00000205, sig00000204, sig00000203, sig00000202, sig00000201, sig00000200, sig000001ff, sig000001fe,
sig000001fd, sig000001fc, sig000001fb, sig000001fa, sig000001f9, sig000001f8, sig000001f7, sig000001f6, sig000001f5, sig000001f4, sig000001f3,
sig000001f2, sig000001f1, sig000001f0, sig000001ef, sig000001ee, sig000001ed, sig000001ec, sig000001eb, sig000001ea, sig000001e9, sig000001e8,
sig000001e7, sig000001e6, sig000001e5, sig000001e4, sig000001e3, sig000001e2, sig000001e1, sig000001e0, sig000001df, sig000001de, sig000001dd,
sig000001dc, sig000001db, sig000001da, sig000001d9, sig000001d8}),
    .ACIN({sig00000284, sig00000283, sig00000282, sig00000281, sig00000280, sig0000027f, sig0000027e, sig0000027d, sig0000027c, sig0000027b,
sig0000027a, sig00000279, sig00000278, sig00000277, sig00000276, sig00000275, sig00000274, sig00000273, sig00000272, sig00000271, sig00000270,
sig0000026f, sig0000026e, sig0000026d, sig0000026c, sig0000026b, sig0000026a, sig00000269, sig00000268, sig00000267}),
    .ALUMODE({sig00000461, sig00000461, sig00000461, sig00000461}),
    .C({sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461
, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461,
sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461,
sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461,
sig00000461, sig00000461, sig00000461, sig00000461}),
    .CARRYOUT({\NLW_blk0000040e_CARRYOUT<3>_UNCONNECTED , \NLW_blk0000040e_CARRYOUT<2>_UNCONNECTED , \NLW_blk0000040e_CARRYOUT<1>_UNCONNECTED ,
\NLW_blk0000040e_CARRYOUT<0>_UNCONNECTED }),
    .BCIN({sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461,
sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461}),
    .BCOUT({\NLW_blk0000040e_BCOUT<17>_UNCONNECTED , \NLW_blk0000040e_BCOUT<16>_UNCONNECTED , \NLW_blk0000040e_BCOUT<15>_UNCONNECTED ,
\NLW_blk0000040e_BCOUT<14>_UNCONNECTED , \NLW_blk0000040e_BCOUT<13>_UNCONNECTED , \NLW_blk0000040e_BCOUT<12>_UNCONNECTED ,
\NLW_blk0000040e_BCOUT<11>_UNCONNECTED , \NLW_blk0000040e_BCOUT<10>_UNCONNECTED , \NLW_blk0000040e_BCOUT<9>_UNCONNECTED ,
\NLW_blk0000040e_BCOUT<8>_UNCONNECTED , \NLW_blk0000040e_BCOUT<7>_UNCONNECTED , \NLW_blk0000040e_BCOUT<6>_UNCONNECTED ,
\NLW_blk0000040e_BCOUT<5>_UNCONNECTED , \NLW_blk0000040e_BCOUT<4>_UNCONNECTED , \NLW_blk0000040e_BCOUT<3>_UNCONNECTED ,
\NLW_blk0000040e_BCOUT<2>_UNCONNECTED , \NLW_blk0000040e_BCOUT<1>_UNCONNECTED , \NLW_blk0000040e_BCOUT<0>_UNCONNECTED }),
    .A({sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461
, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461,
sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461})
  );
  DSP48E #(
    .ACASCREG ( 2 ),
    .ALUMODEREG ( 0 ),
    .AREG ( 2 ),
    .AUTORESET_PATTERN_DETECT ( "FALSE" ),
    .AUTORESET_PATTERN_DETECT_OPTINV ( "MATCH" ),
    .A_INPUT ( "DIRECT" ),
    .BCASCREG ( 2 ),
    .BREG ( 2 ),
    .B_INPUT ( "DIRECT" ),
    .CARRYINREG ( 0 ),
    .CARRYINSELREG ( 0 ),
    .CREG ( 0 ),
    .MASK ( 48'h3FFFFFFFFFFF ),
    .MREG ( 1 ),
    .MULTCARRYINREG ( 0 ),
    .OPMODEREG ( 0 ),
    .PATTERN ( 48'h000000000000 ),
    .PREG ( 1 ),
    .SEL_MASK ( "MASK" ),
    .SEL_PATTERN ( "PATTERN" ),
    .SEL_ROUNDING_MASK ( "SEL_MASK" ),
    .SIM_MODE ( "SAFE" ),
    .USE_MULT ( "MULT_S" ),
    .USE_PATTERN_DETECT ( "NO_PATDET" ),
    .USE_SIMD ( "ONE48" ))
  blk0000040f (
    .CEM(ce),
    .CLK(clk),
    .PATTERNBDETECT(NLW_blk0000040f_PATTERNBDETECT_UNCONNECTED),
    .RSTC(sig00000461),
    .CEB1(ce),
    .MULTSIGNOUT(NLW_blk0000040f_MULTSIGNOUT_UNCONNECTED),
    .CEC(sig00000461),
    .RSTM(sig00000461),
    .MULTSIGNIN(sig00000461),
    .CEB2(ce),
    .RSTCTRL(sig00000461),
    .CEP(ce),
    .CARRYCASCOUT(NLW_blk0000040f_CARRYCASCOUT_UNCONNECTED),
    .RSTA(sig00000461),
    .CECARRYIN(sig00000461),
    .UNDERFLOW(NLW_blk0000040f_UNDERFLOW_UNCONNECTED),
    .PATTERNDETECT(NLW_blk0000040f_PATTERNDETECT_UNCONNECTED),
    .RSTALUMODE(sig00000461),
    .RSTALLCARRYIN(sig00000461),
    .CEALUMODE(sig00000461),
    .CEA2(ce),
    .CEA1(ce),
    .RSTB(sig00000461),
    .CEMULTCARRYIN(sig00000461),
    .OVERFLOW(NLW_blk0000040f_OVERFLOW_UNCONNECTED),
    .CECTRL(sig00000461),
    .CARRYIN(sig00000461),
    .CARRYCASCIN(sig00000461),
    .RSTP(sig00000461),
    .CARRYINSEL({sig00000461, sig00000461, sig00000461}),
    .ACOUT({sig00000284, sig00000283, sig00000282, sig00000281, sig00000280, sig0000027f, sig0000027e, sig0000027d, sig0000027c, sig0000027b,
sig0000027a, sig00000279, sig00000278, sig00000277, sig00000276, sig00000275, sig00000274, sig00000273, sig00000272, sig00000271, sig00000270,
sig0000026f, sig0000026e, sig0000026d, sig0000026c, sig0000026b, sig0000026a, sig00000269, sig00000268, sig00000267}),
    .OPMODE({sig00000461, sig00000461, sig00000001, sig00000461, sig00000001, sig00000461, sig00000001}),
    .PCIN({sig000002b4, sig000002b3, sig000002b2, sig000002b1, sig000002b0, sig000002af, sig000002ae, sig000002ad, sig000002ac, sig000002ab,
sig000002aa, sig000002a9, sig000002a8, sig000002a7, sig000002a6, sig000002a5, sig000002a4, sig000002a3, sig000002a2, sig000002a1, sig000002a0,
sig0000029f, sig0000029e, sig0000029d, sig0000029c, sig0000029b, sig0000029a, sig00000299, sig00000298, sig00000297, sig00000296, sig00000295,
sig00000294, sig00000293, sig00000292, sig00000291, sig00000290, sig0000028f, sig0000028e, sig0000028d, sig0000028c, sig0000028b, sig0000028a,
sig00000289, sig00000288, sig00000287, sig00000286, sig00000285}),
    .B({sig00000461, sig00000126, sig00000127, sig00000128, sig00000129, sig0000012a, sig0000012b, sig0000012c, sig0000012d, sig0000012e, sig0000012f
, sig00000130, sig00000131, sig00000132, sig00000133, sig00000134, sig00000135, sig00000136}),
    .P({\NLW_blk0000040f_P<47>_UNCONNECTED , \NLW_blk0000040f_P<46>_UNCONNECTED , \NLW_blk0000040f_P<45>_UNCONNECTED ,
\NLW_blk0000040f_P<44>_UNCONNECTED , \NLW_blk0000040f_P<43>_UNCONNECTED , \NLW_blk0000040f_P<42>_UNCONNECTED , \NLW_blk0000040f_P<41>_UNCONNECTED ,
\NLW_blk0000040f_P<40>_UNCONNECTED , \NLW_blk0000040f_P<39>_UNCONNECTED , \NLW_blk0000040f_P<38>_UNCONNECTED , \NLW_blk0000040f_P<37>_UNCONNECTED ,
\NLW_blk0000040f_P<36>_UNCONNECTED , \NLW_blk0000040f_P<35>_UNCONNECTED , \NLW_blk0000040f_P<34>_UNCONNECTED , \NLW_blk0000040f_P<33>_UNCONNECTED ,
\NLW_blk0000040f_P<32>_UNCONNECTED , \NLW_blk0000040f_P<31>_UNCONNECTED , \NLW_blk0000040f_P<30>_UNCONNECTED , \NLW_blk0000040f_P<29>_UNCONNECTED ,
\NLW_blk0000040f_P<28>_UNCONNECTED , \NLW_blk0000040f_P<27>_UNCONNECTED , \NLW_blk0000040f_P<26>_UNCONNECTED , \NLW_blk0000040f_P<25>_UNCONNECTED ,
\NLW_blk0000040f_P<24>_UNCONNECTED , \NLW_blk0000040f_P<23>_UNCONNECTED , \NLW_blk0000040f_P<22>_UNCONNECTED , \NLW_blk0000040f_P<21>_UNCONNECTED ,
\NLW_blk0000040f_P<20>_UNCONNECTED , \NLW_blk0000040f_P<19>_UNCONNECTED , \NLW_blk0000040f_P<18>_UNCONNECTED , \NLW_blk0000040f_P<17>_UNCONNECTED ,
sig00000236, sig00000235, sig00000234, sig00000233, sig00000232, sig00000231, sig00000230, sig0000022f, sig0000022e, sig0000022d, sig0000022c,
sig0000022b, sig0000022a, sig00000229, sig00000228, sig00000227, sig00000226}),
    .A({sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461
, sig00000113, sig00000114, sig00000115, sig00000116, sig00000117, sig00000118, sig00000119, sig0000011a, sig0000011b, sig0000011c, sig0000011d,
sig0000011e, sig0000011f, sig00000120, sig00000121, sig00000122, sig00000123, sig00000124, sig00000125}),
    .PCOUT({sig00000266, sig00000265, sig00000264, sig00000263, sig00000262, sig00000261, sig00000260, sig0000025f, sig0000025e, sig0000025d,
sig0000025c, sig0000025b, sig0000025a, sig00000259, sig00000258, sig00000257, sig00000256, sig00000255, sig00000254, sig00000253, sig00000252,
sig00000251, sig00000250, sig0000024f, sig0000024e, sig0000024d, sig0000024c, sig0000024b, sig0000024a, sig00000249, sig00000248, sig00000247,
sig00000246, sig00000245, sig00000244, sig00000243, sig00000242, sig00000241, sig00000240, sig0000023f, sig0000023e, sig0000023d, sig0000023c,
sig0000023b, sig0000023a, sig00000239, sig00000238, sig00000237}),
    .ALUMODE({sig00000461, sig00000461, sig00000461, sig00000461}),
    .C({sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461
, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461,
sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461,
sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461,
sig00000461, sig00000461, sig00000461, sig00000461}),
    .CARRYOUT({\NLW_blk0000040f_CARRYOUT<3>_UNCONNECTED , \NLW_blk0000040f_CARRYOUT<2>_UNCONNECTED , \NLW_blk0000040f_CARRYOUT<1>_UNCONNECTED ,
\NLW_blk0000040f_CARRYOUT<0>_UNCONNECTED }),
    .BCIN({sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461,
sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461}),
    .BCOUT({\NLW_blk0000040f_BCOUT<17>_UNCONNECTED , \NLW_blk0000040f_BCOUT<16>_UNCONNECTED , \NLW_blk0000040f_BCOUT<15>_UNCONNECTED ,
\NLW_blk0000040f_BCOUT<14>_UNCONNECTED , \NLW_blk0000040f_BCOUT<13>_UNCONNECTED , \NLW_blk0000040f_BCOUT<12>_UNCONNECTED ,
\NLW_blk0000040f_BCOUT<11>_UNCONNECTED , \NLW_blk0000040f_BCOUT<10>_UNCONNECTED , \NLW_blk0000040f_BCOUT<9>_UNCONNECTED ,
\NLW_blk0000040f_BCOUT<8>_UNCONNECTED , \NLW_blk0000040f_BCOUT<7>_UNCONNECTED , \NLW_blk0000040f_BCOUT<6>_UNCONNECTED ,
\NLW_blk0000040f_BCOUT<5>_UNCONNECTED , \NLW_blk0000040f_BCOUT<4>_UNCONNECTED , \NLW_blk0000040f_BCOUT<3>_UNCONNECTED ,
\NLW_blk0000040f_BCOUT<2>_UNCONNECTED , \NLW_blk0000040f_BCOUT<1>_UNCONNECTED , \NLW_blk0000040f_BCOUT<0>_UNCONNECTED }),
    .ACIN({sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461,
sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461,
sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461})
  );
  DSP48E #(
    .ACASCREG ( 1 ),
    .ALUMODEREG ( 0 ),
    .AREG ( 1 ),
    .AUTORESET_PATTERN_DETECT ( "FALSE" ),
    .AUTORESET_PATTERN_DETECT_OPTINV ( "MATCH" ),
    .A_INPUT ( "CASCADE" ),
    .BCASCREG ( 2 ),
    .BREG ( 2 ),
    .B_INPUT ( "DIRECT" ),
    .CARRYINREG ( 0 ),
    .CARRYINSELREG ( 0 ),
    .CREG ( 0 ),
    .MASK ( 48'h3FFFFFFFFFFF ),
    .MREG ( 1 ),
    .MULTCARRYINREG ( 0 ),
    .OPMODEREG ( 0 ),
    .PATTERN ( 48'h000000000000 ),
    .PREG ( 1 ),
    .SEL_MASK ( "MASK" ),
    .SEL_PATTERN ( "PATTERN" ),
    .SEL_ROUNDING_MASK ( "SEL_MASK" ),
    .SIM_MODE ( "SAFE" ),
    .USE_MULT ( "MULT_S" ),
    .USE_PATTERN_DETECT ( "NO_PATDET" ),
    .USE_SIMD ( "ONE48" ))
  blk00000410 (
    .CEM(ce),
    .CLK(clk),
    .PATTERNBDETECT(NLW_blk00000410_PATTERNBDETECT_UNCONNECTED),
    .RSTC(sig00000461),
    .CEB1(ce),
    .MULTSIGNOUT(NLW_blk00000410_MULTSIGNOUT_UNCONNECTED),
    .CEC(sig00000461),
    .RSTM(sig00000461),
    .MULTSIGNIN(sig00000461),
    .CEB2(ce),
    .RSTCTRL(sig00000461),
    .CEP(ce),
    .CARRYCASCOUT(NLW_blk00000410_CARRYCASCOUT_UNCONNECTED),
    .RSTA(sig00000461),
    .CECARRYIN(sig00000461),
    .UNDERFLOW(NLW_blk00000410_UNDERFLOW_UNCONNECTED),
    .PATTERNDETECT(NLW_blk00000410_PATTERNDETECT_UNCONNECTED),
    .RSTALUMODE(sig00000461),
    .RSTALLCARRYIN(sig00000461),
    .CEALUMODE(sig00000461),
    .CEA2(ce),
    .CEA1(sig00000461),
    .RSTB(sig00000461),
    .CEMULTCARRYIN(sig00000461),
    .OVERFLOW(NLW_blk00000410_OVERFLOW_UNCONNECTED),
    .CECTRL(sig00000461),
    .CARRYIN(sig00000461),
    .CARRYCASCIN(sig00000461),
    .RSTP(sig00000461),
    .CARRYINSEL({sig00000461, sig00000461, sig00000461}),
    .OPMODE({sig00000001, sig00000461, sig00000001, sig00000461, sig00000001, sig00000461, sig00000001}),
    .PCIN({sig000002e5, sig000002e4, sig000002e3, sig000002e2, sig000002e1, sig000002e0, sig000002df, sig000002de, sig000002dd, sig000002dc,
sig000002db, sig000002da, sig000002d9, sig000002d8, sig000002d7, sig000002d6, sig000002d5, sig000002d4, sig000002d3, sig000002d2, sig000002d1,
sig000002d0, sig000002cf, sig000002ce, sig000002cd, sig000002cc, sig000002cb, sig000002ca, sig000002c9, sig000002c8, sig000002c7, sig000002c6,
sig000002c5, sig000002c4, sig000002c3, sig000002c2, sig000002c1, sig000002c0, sig000002bf, sig000002be, sig000002bd, sig000002bc, sig000002bb,
sig000002ba, sig000002b9, sig000002b8, sig000002b7, sig000002b6}),
    .B({sig00000461, sig00000137, sig00000138, sig00000139, sig0000013a, sig0000013b, sig0000013c, sig0000013d, sig0000013e, sig0000013f, sig00000140
, sig00000141, sig00000142, sig00000143, sig00000144, sig00000145, sig00000146, sig00000147}),
    .PCOUT({sig000002b4, sig000002b3, sig000002b2, sig000002b1, sig000002b0, sig000002af, sig000002ae, sig000002ad, sig000002ac, sig000002ab,
sig000002aa, sig000002a9, sig000002a8, sig000002a7, sig000002a6, sig000002a5, sig000002a4, sig000002a3, sig000002a2, sig000002a1, sig000002a0,
sig0000029f, sig0000029e, sig0000029d, sig0000029c, sig0000029b, sig0000029a, sig00000299, sig00000298, sig00000297, sig00000296, sig00000295,
sig00000294, sig00000293, sig00000292, sig00000291, sig00000290, sig0000028f, sig0000028e, sig0000028d, sig0000028c, sig0000028b, sig0000028a,
sig00000289, sig00000288, sig00000287, sig00000286, sig00000285}),
    .ACIN({sig00000303, sig00000302, sig00000301, sig00000300, sig000002ff, sig000002fe, sig000002fd, sig000002fc, sig000002fb, sig000002fa,
sig000002f9, sig000002f8, sig000002f7, sig000002f6, sig000002f5, sig000002f4, sig000002f3, sig000002f2, sig000002f1, sig000002f0, sig000002ef,
sig000002ee, sig000002ed, sig000002ec, sig000002eb, sig000002ea, sig000002e9, sig000002e8, sig000002e7, sig000002e6}),
    .ACOUT({\NLW_blk00000410_ACOUT<29>_UNCONNECTED , \NLW_blk00000410_ACOUT<28>_UNCONNECTED , \NLW_blk00000410_ACOUT<27>_UNCONNECTED ,
\NLW_blk00000410_ACOUT<26>_UNCONNECTED , \NLW_blk00000410_ACOUT<25>_UNCONNECTED , \NLW_blk00000410_ACOUT<24>_UNCONNECTED ,
\NLW_blk00000410_ACOUT<23>_UNCONNECTED , \NLW_blk00000410_ACOUT<22>_UNCONNECTED , \NLW_blk00000410_ACOUT<21>_UNCONNECTED ,
\NLW_blk00000410_ACOUT<20>_UNCONNECTED , \NLW_blk00000410_ACOUT<19>_UNCONNECTED , \NLW_blk00000410_ACOUT<18>_UNCONNECTED ,
\NLW_blk00000410_ACOUT<17>_UNCONNECTED , \NLW_blk00000410_ACOUT<16>_UNCONNECTED , \NLW_blk00000410_ACOUT<15>_UNCONNECTED ,
\NLW_blk00000410_ACOUT<14>_UNCONNECTED , \NLW_blk00000410_ACOUT<13>_UNCONNECTED , \NLW_blk00000410_ACOUT<12>_UNCONNECTED ,
\NLW_blk00000410_ACOUT<11>_UNCONNECTED , \NLW_blk00000410_ACOUT<10>_UNCONNECTED , \NLW_blk00000410_ACOUT<9>_UNCONNECTED ,
\NLW_blk00000410_ACOUT<8>_UNCONNECTED , \NLW_blk00000410_ACOUT<7>_UNCONNECTED , \NLW_blk00000410_ACOUT<6>_UNCONNECTED ,
\NLW_blk00000410_ACOUT<5>_UNCONNECTED , \NLW_blk00000410_ACOUT<4>_UNCONNECTED , \NLW_blk00000410_ACOUT<3>_UNCONNECTED ,
\NLW_blk00000410_ACOUT<2>_UNCONNECTED , \NLW_blk00000410_ACOUT<1>_UNCONNECTED , \NLW_blk00000410_ACOUT<0>_UNCONNECTED }),
    .ALUMODE({sig00000461, sig00000461, sig00000461, sig00000461}),
    .C({sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461
, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461,
sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461,
sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461,
sig00000461, sig00000461, sig00000461, sig00000461}),
    .CARRYOUT({\NLW_blk00000410_CARRYOUT<3>_UNCONNECTED , \NLW_blk00000410_CARRYOUT<2>_UNCONNECTED , \NLW_blk00000410_CARRYOUT<1>_UNCONNECTED ,
\NLW_blk00000410_CARRYOUT<0>_UNCONNECTED }),
    .BCIN({sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461,
sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461}),
    .BCOUT({\NLW_blk00000410_BCOUT<17>_UNCONNECTED , \NLW_blk00000410_BCOUT<16>_UNCONNECTED , \NLW_blk00000410_BCOUT<15>_UNCONNECTED ,
\NLW_blk00000410_BCOUT<14>_UNCONNECTED , \NLW_blk00000410_BCOUT<13>_UNCONNECTED , \NLW_blk00000410_BCOUT<12>_UNCONNECTED ,
\NLW_blk00000410_BCOUT<11>_UNCONNECTED , \NLW_blk00000410_BCOUT<10>_UNCONNECTED , \NLW_blk00000410_BCOUT<9>_UNCONNECTED ,
\NLW_blk00000410_BCOUT<8>_UNCONNECTED , \NLW_blk00000410_BCOUT<7>_UNCONNECTED , \NLW_blk00000410_BCOUT<6>_UNCONNECTED ,
\NLW_blk00000410_BCOUT<5>_UNCONNECTED , \NLW_blk00000410_BCOUT<4>_UNCONNECTED , \NLW_blk00000410_BCOUT<3>_UNCONNECTED ,
\NLW_blk00000410_BCOUT<2>_UNCONNECTED , \NLW_blk00000410_BCOUT<1>_UNCONNECTED , \NLW_blk00000410_BCOUT<0>_UNCONNECTED }),
    .P({\NLW_blk00000410_P<47>_UNCONNECTED , \NLW_blk00000410_P<46>_UNCONNECTED , \NLW_blk00000410_P<45>_UNCONNECTED ,
\NLW_blk00000410_P<44>_UNCONNECTED , \NLW_blk00000410_P<43>_UNCONNECTED , \NLW_blk00000410_P<42>_UNCONNECTED , \NLW_blk00000410_P<41>_UNCONNECTED ,
\NLW_blk00000410_P<40>_UNCONNECTED , \NLW_blk00000410_P<39>_UNCONNECTED , \NLW_blk00000410_P<38>_UNCONNECTED , \NLW_blk00000410_P<37>_UNCONNECTED ,
\NLW_blk00000410_P<36>_UNCONNECTED , \NLW_blk00000410_P<35>_UNCONNECTED , \NLW_blk00000410_P<34>_UNCONNECTED , \NLW_blk00000410_P<33>_UNCONNECTED ,
\NLW_blk00000410_P<32>_UNCONNECTED , \NLW_blk00000410_P<31>_UNCONNECTED , \NLW_blk00000410_P<30>_UNCONNECTED , \NLW_blk00000410_P<29>_UNCONNECTED ,
\NLW_blk00000410_P<28>_UNCONNECTED , \NLW_blk00000410_P<27>_UNCONNECTED , \NLW_blk00000410_P<26>_UNCONNECTED , \NLW_blk00000410_P<25>_UNCONNECTED ,
\NLW_blk00000410_P<24>_UNCONNECTED , \NLW_blk00000410_P<23>_UNCONNECTED , \NLW_blk00000410_P<22>_UNCONNECTED , \NLW_blk00000410_P<21>_UNCONNECTED ,
\NLW_blk00000410_P<20>_UNCONNECTED , \NLW_blk00000410_P<19>_UNCONNECTED , \NLW_blk00000410_P<18>_UNCONNECTED , \NLW_blk00000410_P<17>_UNCONNECTED ,
\NLW_blk00000410_P<16>_UNCONNECTED , \NLW_blk00000410_P<15>_UNCONNECTED , \NLW_blk00000410_P<14>_UNCONNECTED , \NLW_blk00000410_P<13>_UNCONNECTED ,
\NLW_blk00000410_P<12>_UNCONNECTED , \NLW_blk00000410_P<11>_UNCONNECTED , \NLW_blk00000410_P<10>_UNCONNECTED , \NLW_blk00000410_P<9>_UNCONNECTED ,
\NLW_blk00000410_P<8>_UNCONNECTED , \NLW_blk00000410_P<7>_UNCONNECTED , \NLW_blk00000410_P<6>_UNCONNECTED , \NLW_blk00000410_P<5>_UNCONNECTED ,
\NLW_blk00000410_P<4>_UNCONNECTED , \NLW_blk00000410_P<3>_UNCONNECTED , \NLW_blk00000410_P<2>_UNCONNECTED , \NLW_blk00000410_P<1>_UNCONNECTED ,
\NLW_blk00000410_P<0>_UNCONNECTED }),
    .A({sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461
, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461,
sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461})
  );
  DSP48E #(
    .ACASCREG ( 2 ),
    .ALUMODEREG ( 0 ),
    .AREG ( 2 ),
    .AUTORESET_PATTERN_DETECT ( "FALSE" ),
    .AUTORESET_PATTERN_DETECT_OPTINV ( "MATCH" ),
    .A_INPUT ( "DIRECT" ),
    .BCASCREG ( 2 ),
    .BREG ( 2 ),
    .B_INPUT ( "DIRECT" ),
    .CARRYINREG ( 0 ),
    .CARRYINSELREG ( 0 ),
    .CREG ( 0 ),
    .MASK ( 48'hFFFFFFFE0000 ),
    .MREG ( 1 ),
    .MULTCARRYINREG ( 0 ),
    .OPMODEREG ( 0 ),
    .PATTERN ( 48'h000000000000 ),
    .PREG ( 1 ),
    .SEL_MASK ( "MASK" ),
    .SEL_PATTERN ( "PATTERN" ),
    .SEL_ROUNDING_MASK ( "SEL_MASK" ),
    .SIM_MODE ( "SAFE" ),
    .USE_MULT ( "MULT_S" ),
    .USE_PATTERN_DETECT ( "PATDET" ),
    .USE_SIMD ( "ONE48" ))
  blk00000411 (
    .CEM(ce),
    .PATTERNDETECT(sig000002b5),
    .CLK(clk),
    .PATTERNBDETECT(NLW_blk00000411_PATTERNBDETECT_UNCONNECTED),
    .RSTC(sig00000461),
    .CEB1(ce),
    .MULTSIGNOUT(NLW_blk00000411_MULTSIGNOUT_UNCONNECTED),
    .CEC(sig00000461),
    .RSTM(sig00000461),
    .MULTSIGNIN(sig00000461),
    .CEB2(ce),
    .RSTCTRL(sig00000461),
    .CEP(ce),
    .CARRYCASCOUT(NLW_blk00000411_CARRYCASCOUT_UNCONNECTED),
    .RSTA(sig00000461),
    .CECARRYIN(sig00000461),
    .UNDERFLOW(NLW_blk00000411_UNDERFLOW_UNCONNECTED),
    .RSTALUMODE(sig00000461),
    .RSTALLCARRYIN(sig00000461),
    .CEALUMODE(sig00000461),
    .CEA2(ce),
    .CEA1(ce),
    .RSTB(sig00000461),
    .CEMULTCARRYIN(sig00000461),
    .OVERFLOW(NLW_blk00000411_OVERFLOW_UNCONNECTED),
    .CECTRL(sig00000461),
    .CARRYIN(sig00000461),
    .CARRYCASCIN(sig00000461),
    .RSTP(sig00000461),
    .CARRYINSEL({sig00000461, sig00000461, sig00000461}),
    .ACOUT({sig00000303, sig00000302, sig00000301, sig00000300, sig000002ff, sig000002fe, sig000002fd, sig000002fc, sig000002fb, sig000002fa,
sig000002f9, sig000002f8, sig000002f7, sig000002f6, sig000002f5, sig000002f4, sig000002f3, sig000002f2, sig000002f1, sig000002f0, sig000002ef,
sig000002ee, sig000002ed, sig000002ec, sig000002eb, sig000002ea, sig000002e9, sig000002e8, sig000002e7, sig000002e6}),
    .OPMODE({sig00000461, sig00000461, sig00000001, sig00000461, sig00000001, sig00000461, sig00000001}),
    .PCIN({sig00000333, sig00000332, sig00000331, sig00000330, sig0000032f, sig0000032e, sig0000032d, sig0000032c, sig0000032b, sig0000032a,
sig00000329, sig00000328, sig00000327, sig00000326, sig00000325, sig00000324, sig00000323, sig00000322, sig00000321, sig00000320, sig0000031f,
sig0000031e, sig0000031d, sig0000031c, sig0000031b, sig0000031a, sig00000319, sig00000318, sig00000317, sig00000316, sig00000315, sig00000314,
sig00000313, sig00000312, sig00000311, sig00000310, sig0000030f, sig0000030e, sig0000030d, sig0000030c, sig0000030b, sig0000030a, sig00000309,
sig00000308, sig00000307, sig00000306, sig00000305, sig00000304}),
    .B({sig00000461, sig0000015c, sig0000015d, sig0000015e, sig0000015f, sig00000160, sig00000161, sig00000162, sig00000163, sig00000164, sig00000165
, sig00000166, sig00000167, sig00000168, sig00000169, sig0000016a, sig0000016b, sig0000016c}),
    .A({sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461
, sig00000149, sig0000014a, sig0000014b, sig0000014c, sig0000014d, sig0000014e, sig0000014f, sig00000150, sig00000151, sig00000152, sig00000153,
sig00000154, sig00000155, sig00000156, sig00000157, sig00000158, sig00000159, sig0000015a, sig0000015b}),
    .PCOUT({sig000002e5, sig000002e4, sig000002e3, sig000002e2, sig000002e1, sig000002e0, sig000002df, sig000002de, sig000002dd, sig000002dc,
sig000002db, sig000002da, sig000002d9, sig000002d8, sig000002d7, sig000002d6, sig000002d5, sig000002d4, sig000002d3, sig000002d2, sig000002d1,
sig000002d0, sig000002cf, sig000002ce, sig000002cd, sig000002cc, sig000002cb, sig000002ca, sig000002c9, sig000002c8, sig000002c7, sig000002c6,
sig000002c5, sig000002c4, sig000002c3, sig000002c2, sig000002c1, sig000002c0, sig000002bf, sig000002be, sig000002bd, sig000002bc, sig000002bb,
sig000002ba, sig000002b9, sig000002b8, sig000002b7, sig000002b6}),
    .ALUMODE({sig00000461, sig00000461, sig00000461, sig00000461}),
    .C({sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461
, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461,
sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461,
sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461,
sig00000461, sig00000461, sig00000461, sig00000461}),
    .CARRYOUT({\NLW_blk00000411_CARRYOUT<3>_UNCONNECTED , \NLW_blk00000411_CARRYOUT<2>_UNCONNECTED , \NLW_blk00000411_CARRYOUT<1>_UNCONNECTED ,
\NLW_blk00000411_CARRYOUT<0>_UNCONNECTED }),
    .BCIN({sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461,
sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461}),
    .BCOUT({\NLW_blk00000411_BCOUT<17>_UNCONNECTED , \NLW_blk00000411_BCOUT<16>_UNCONNECTED , \NLW_blk00000411_BCOUT<15>_UNCONNECTED ,
\NLW_blk00000411_BCOUT<14>_UNCONNECTED , \NLW_blk00000411_BCOUT<13>_UNCONNECTED , \NLW_blk00000411_BCOUT<12>_UNCONNECTED ,
\NLW_blk00000411_BCOUT<11>_UNCONNECTED , \NLW_blk00000411_BCOUT<10>_UNCONNECTED , \NLW_blk00000411_BCOUT<9>_UNCONNECTED ,
\NLW_blk00000411_BCOUT<8>_UNCONNECTED , \NLW_blk00000411_BCOUT<7>_UNCONNECTED , \NLW_blk00000411_BCOUT<6>_UNCONNECTED ,
\NLW_blk00000411_BCOUT<5>_UNCONNECTED , \NLW_blk00000411_BCOUT<4>_UNCONNECTED , \NLW_blk00000411_BCOUT<3>_UNCONNECTED ,
\NLW_blk00000411_BCOUT<2>_UNCONNECTED , \NLW_blk00000411_BCOUT<1>_UNCONNECTED , \NLW_blk00000411_BCOUT<0>_UNCONNECTED }),
    .P({\NLW_blk00000411_P<47>_UNCONNECTED , \NLW_blk00000411_P<46>_UNCONNECTED , \NLW_blk00000411_P<45>_UNCONNECTED ,
\NLW_blk00000411_P<44>_UNCONNECTED , \NLW_blk00000411_P<43>_UNCONNECTED , \NLW_blk00000411_P<42>_UNCONNECTED , \NLW_blk00000411_P<41>_UNCONNECTED ,
\NLW_blk00000411_P<40>_UNCONNECTED , \NLW_blk00000411_P<39>_UNCONNECTED , \NLW_blk00000411_P<38>_UNCONNECTED , \NLW_blk00000411_P<37>_UNCONNECTED ,
\NLW_blk00000411_P<36>_UNCONNECTED , \NLW_blk00000411_P<35>_UNCONNECTED , \NLW_blk00000411_P<34>_UNCONNECTED , \NLW_blk00000411_P<33>_UNCONNECTED ,
\NLW_blk00000411_P<32>_UNCONNECTED , \NLW_blk00000411_P<31>_UNCONNECTED , \NLW_blk00000411_P<30>_UNCONNECTED , \NLW_blk00000411_P<29>_UNCONNECTED ,
\NLW_blk00000411_P<28>_UNCONNECTED , \NLW_blk00000411_P<27>_UNCONNECTED , \NLW_blk00000411_P<26>_UNCONNECTED , \NLW_blk00000411_P<25>_UNCONNECTED ,
\NLW_blk00000411_P<24>_UNCONNECTED , \NLW_blk00000411_P<23>_UNCONNECTED , \NLW_blk00000411_P<22>_UNCONNECTED , \NLW_blk00000411_P<21>_UNCONNECTED ,
\NLW_blk00000411_P<20>_UNCONNECTED , \NLW_blk00000411_P<19>_UNCONNECTED , \NLW_blk00000411_P<18>_UNCONNECTED , \NLW_blk00000411_P<17>_UNCONNECTED ,
\NLW_blk00000411_P<16>_UNCONNECTED , \NLW_blk00000411_P<15>_UNCONNECTED , \NLW_blk00000411_P<14>_UNCONNECTED , \NLW_blk00000411_P<13>_UNCONNECTED ,
\NLW_blk00000411_P<12>_UNCONNECTED , \NLW_blk00000411_P<11>_UNCONNECTED , \NLW_blk00000411_P<10>_UNCONNECTED , \NLW_blk00000411_P<9>_UNCONNECTED ,
\NLW_blk00000411_P<8>_UNCONNECTED , \NLW_blk00000411_P<7>_UNCONNECTED , \NLW_blk00000411_P<6>_UNCONNECTED , \NLW_blk00000411_P<5>_UNCONNECTED ,
\NLW_blk00000411_P<4>_UNCONNECTED , \NLW_blk00000411_P<3>_UNCONNECTED , \NLW_blk00000411_P<2>_UNCONNECTED , \NLW_blk00000411_P<1>_UNCONNECTED ,
\NLW_blk00000411_P<0>_UNCONNECTED }),
    .ACIN({sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461,
sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461,
sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461})
  );
  DSP48E #(
    .ACASCREG ( 2 ),
    .ALUMODEREG ( 0 ),
    .AREG ( 2 ),
    .AUTORESET_PATTERN_DETECT ( "FALSE" ),
    .AUTORESET_PATTERN_DETECT_OPTINV ( "MATCH" ),
    .A_INPUT ( "DIRECT" ),
    .BCASCREG ( 2 ),
    .BREG ( 2 ),
    .B_INPUT ( "DIRECT" ),
    .CARRYINREG ( 0 ),
    .CARRYINSELREG ( 0 ),
    .CREG ( 0 ),
    .MASK ( 48'h3FFFFFFFFFFF ),
    .MREG ( 1 ),
    .MULTCARRYINREG ( 0 ),
    .OPMODEREG ( 0 ),
    .PATTERN ( 48'h000000000000 ),
    .PREG ( 1 ),
    .SEL_MASK ( "MASK" ),
    .SEL_PATTERN ( "PATTERN" ),
    .SEL_ROUNDING_MASK ( "SEL_MASK" ),
    .SIM_MODE ( "SAFE" ),
    .USE_MULT ( "MULT_S" ),
    .USE_PATTERN_DETECT ( "NO_PATDET" ),
    .USE_SIMD ( "ONE48" ))
  blk00000412 (
    .CEM(ce),
    .CLK(clk),
    .PATTERNBDETECT(NLW_blk00000412_PATTERNBDETECT_UNCONNECTED),
    .RSTC(sig00000461),
    .CEB1(ce),
    .MULTSIGNOUT(NLW_blk00000412_MULTSIGNOUT_UNCONNECTED),
    .CEC(sig00000461),
    .RSTM(sig00000461),
    .MULTSIGNIN(sig00000461),
    .CEB2(ce),
    .RSTCTRL(sig00000461),
    .CEP(ce),
    .CARRYCASCOUT(NLW_blk00000412_CARRYCASCOUT_UNCONNECTED),
    .RSTA(sig00000461),
    .CECARRYIN(sig00000461),
    .UNDERFLOW(NLW_blk00000412_UNDERFLOW_UNCONNECTED),
    .PATTERNDETECT(NLW_blk00000412_PATTERNDETECT_UNCONNECTED),
    .RSTALUMODE(sig00000461),
    .RSTALLCARRYIN(sig00000461),
    .CEALUMODE(sig00000461),
    .CEA2(ce),
    .CEA1(ce),
    .RSTB(sig00000461),
    .CEMULTCARRYIN(sig00000461),
    .OVERFLOW(NLW_blk00000412_OVERFLOW_UNCONNECTED),
    .CECTRL(sig00000461),
    .CARRYIN(sig00000461),
    .CARRYCASCIN(sig00000461),
    .RSTP(sig00000461),
    .CARRYINSEL({sig00000461, sig00000461, sig00000461}),
    .OPMODE({sig00000461, sig00000461, sig00000001, sig00000461, sig00000001, sig00000461, sig00000001}),
    .PCIN({sig00000363, sig00000362, sig00000361, sig00000360, sig0000035f, sig0000035e, sig0000035d, sig0000035c, sig0000035b, sig0000035a,
sig00000359, sig00000358, sig00000357, sig00000356, sig00000355, sig00000354, sig00000353, sig00000352, sig00000351, sig00000350, sig0000034f,
sig0000034e, sig0000034d, sig0000034c, sig0000034b, sig0000034a, sig00000349, sig00000348, sig00000347, sig00000346, sig00000345, sig00000344,
sig00000343, sig00000342, sig00000341, sig00000340, sig0000033f, sig0000033e, sig0000033d, sig0000033c, sig0000033b, sig0000033a, sig00000339,
sig00000338, sig00000337, sig00000336, sig00000335, sig00000334}),
    .B({sig00000461, sig00000180, sig00000181, sig00000182, sig00000183, sig00000184, sig00000185, sig00000186, sig00000187, sig00000188, sig00000189
, sig0000018a, sig0000018b, sig0000018c, sig0000018d, sig0000018e, sig0000018f, sig00000190}),
    .A({sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461
, sig0000016d, sig0000016e, sig0000016f, sig00000170, sig00000171, sig00000172, sig00000173, sig00000174, sig00000175, sig00000176, sig00000177,
sig00000178, sig00000179, sig0000017a, sig0000017b, sig0000017c, sig0000017d, sig0000017e, sig0000017f}),
    .PCOUT({sig00000333, sig00000332, sig00000331, sig00000330, sig0000032f, sig0000032e, sig0000032d, sig0000032c, sig0000032b, sig0000032a,
sig00000329, sig00000328, sig00000327, sig00000326, sig00000325, sig00000324, sig00000323, sig00000322, sig00000321, sig00000320, sig0000031f,
sig0000031e, sig0000031d, sig0000031c, sig0000031b, sig0000031a, sig00000319, sig00000318, sig00000317, sig00000316, sig00000315, sig00000314,
sig00000313, sig00000312, sig00000311, sig00000310, sig0000030f, sig0000030e, sig0000030d, sig0000030c, sig0000030b, sig0000030a, sig00000309,
sig00000308, sig00000307, sig00000306, sig00000305, sig00000304}),
    .ACOUT({\NLW_blk00000412_ACOUT<29>_UNCONNECTED , \NLW_blk00000412_ACOUT<28>_UNCONNECTED , \NLW_blk00000412_ACOUT<27>_UNCONNECTED ,
\NLW_blk00000412_ACOUT<26>_UNCONNECTED , \NLW_blk00000412_ACOUT<25>_UNCONNECTED , \NLW_blk00000412_ACOUT<24>_UNCONNECTED ,
\NLW_blk00000412_ACOUT<23>_UNCONNECTED , \NLW_blk00000412_ACOUT<22>_UNCONNECTED , \NLW_blk00000412_ACOUT<21>_UNCONNECTED ,
\NLW_blk00000412_ACOUT<20>_UNCONNECTED , \NLW_blk00000412_ACOUT<19>_UNCONNECTED , \NLW_blk00000412_ACOUT<18>_UNCONNECTED ,
\NLW_blk00000412_ACOUT<17>_UNCONNECTED , \NLW_blk00000412_ACOUT<16>_UNCONNECTED , \NLW_blk00000412_ACOUT<15>_UNCONNECTED ,
\NLW_blk00000412_ACOUT<14>_UNCONNECTED , \NLW_blk00000412_ACOUT<13>_UNCONNECTED , \NLW_blk00000412_ACOUT<12>_UNCONNECTED ,
\NLW_blk00000412_ACOUT<11>_UNCONNECTED , \NLW_blk00000412_ACOUT<10>_UNCONNECTED , \NLW_blk00000412_ACOUT<9>_UNCONNECTED ,
\NLW_blk00000412_ACOUT<8>_UNCONNECTED , \NLW_blk00000412_ACOUT<7>_UNCONNECTED , \NLW_blk00000412_ACOUT<6>_UNCONNECTED ,
\NLW_blk00000412_ACOUT<5>_UNCONNECTED , \NLW_blk00000412_ACOUT<4>_UNCONNECTED , \NLW_blk00000412_ACOUT<3>_UNCONNECTED ,
\NLW_blk00000412_ACOUT<2>_UNCONNECTED , \NLW_blk00000412_ACOUT<1>_UNCONNECTED , \NLW_blk00000412_ACOUT<0>_UNCONNECTED }),
    .ALUMODE({sig00000461, sig00000461, sig00000461, sig00000461}),
    .C({sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461
, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461,
sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461,
sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461,
sig00000461, sig00000461, sig00000461, sig00000461}),
    .CARRYOUT({\NLW_blk00000412_CARRYOUT<3>_UNCONNECTED , \NLW_blk00000412_CARRYOUT<2>_UNCONNECTED , \NLW_blk00000412_CARRYOUT<1>_UNCONNECTED ,
\NLW_blk00000412_CARRYOUT<0>_UNCONNECTED }),
    .BCIN({sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461,
sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461}),
    .BCOUT({\NLW_blk00000412_BCOUT<17>_UNCONNECTED , \NLW_blk00000412_BCOUT<16>_UNCONNECTED , \NLW_blk00000412_BCOUT<15>_UNCONNECTED ,
\NLW_blk00000412_BCOUT<14>_UNCONNECTED , \NLW_blk00000412_BCOUT<13>_UNCONNECTED , \NLW_blk00000412_BCOUT<12>_UNCONNECTED ,
\NLW_blk00000412_BCOUT<11>_UNCONNECTED , \NLW_blk00000412_BCOUT<10>_UNCONNECTED , \NLW_blk00000412_BCOUT<9>_UNCONNECTED ,
\NLW_blk00000412_BCOUT<8>_UNCONNECTED , \NLW_blk00000412_BCOUT<7>_UNCONNECTED , \NLW_blk00000412_BCOUT<6>_UNCONNECTED ,
\NLW_blk00000412_BCOUT<5>_UNCONNECTED , \NLW_blk00000412_BCOUT<4>_UNCONNECTED , \NLW_blk00000412_BCOUT<3>_UNCONNECTED ,
\NLW_blk00000412_BCOUT<2>_UNCONNECTED , \NLW_blk00000412_BCOUT<1>_UNCONNECTED , \NLW_blk00000412_BCOUT<0>_UNCONNECTED }),
    .P({\NLW_blk00000412_P<47>_UNCONNECTED , \NLW_blk00000412_P<46>_UNCONNECTED , \NLW_blk00000412_P<45>_UNCONNECTED ,
\NLW_blk00000412_P<44>_UNCONNECTED , \NLW_blk00000412_P<43>_UNCONNECTED , \NLW_blk00000412_P<42>_UNCONNECTED , \NLW_blk00000412_P<41>_UNCONNECTED ,
\NLW_blk00000412_P<40>_UNCONNECTED , \NLW_blk00000412_P<39>_UNCONNECTED , \NLW_blk00000412_P<38>_UNCONNECTED , \NLW_blk00000412_P<37>_UNCONNECTED ,
\NLW_blk00000412_P<36>_UNCONNECTED , \NLW_blk00000412_P<35>_UNCONNECTED , \NLW_blk00000412_P<34>_UNCONNECTED , \NLW_blk00000412_P<33>_UNCONNECTED ,
\NLW_blk00000412_P<32>_UNCONNECTED , \NLW_blk00000412_P<31>_UNCONNECTED , \NLW_blk00000412_P<30>_UNCONNECTED , \NLW_blk00000412_P<29>_UNCONNECTED ,
\NLW_blk00000412_P<28>_UNCONNECTED , \NLW_blk00000412_P<27>_UNCONNECTED , \NLW_blk00000412_P<26>_UNCONNECTED , \NLW_blk00000412_P<25>_UNCONNECTED ,
\NLW_blk00000412_P<24>_UNCONNECTED , \NLW_blk00000412_P<23>_UNCONNECTED , \NLW_blk00000412_P<22>_UNCONNECTED , \NLW_blk00000412_P<21>_UNCONNECTED ,
\NLW_blk00000412_P<20>_UNCONNECTED , \NLW_blk00000412_P<19>_UNCONNECTED , \NLW_blk00000412_P<18>_UNCONNECTED , \NLW_blk00000412_P<17>_UNCONNECTED ,
\NLW_blk00000412_P<16>_UNCONNECTED , \NLW_blk00000412_P<15>_UNCONNECTED , \NLW_blk00000412_P<14>_UNCONNECTED , \NLW_blk00000412_P<13>_UNCONNECTED ,
\NLW_blk00000412_P<12>_UNCONNECTED , \NLW_blk00000412_P<11>_UNCONNECTED , \NLW_blk00000412_P<10>_UNCONNECTED , \NLW_blk00000412_P<9>_UNCONNECTED ,
\NLW_blk00000412_P<8>_UNCONNECTED , \NLW_blk00000412_P<7>_UNCONNECTED , \NLW_blk00000412_P<6>_UNCONNECTED , \NLW_blk00000412_P<5>_UNCONNECTED ,
\NLW_blk00000412_P<4>_UNCONNECTED , \NLW_blk00000412_P<3>_UNCONNECTED , \NLW_blk00000412_P<2>_UNCONNECTED , \NLW_blk00000412_P<1>_UNCONNECTED ,
\NLW_blk00000412_P<0>_UNCONNECTED }),
    .ACIN({sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461,
sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461,
sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461})
  );
  DSP48E #(
    .ACASCREG ( 2 ),
    .ALUMODEREG ( 0 ),
    .AREG ( 2 ),
    .AUTORESET_PATTERN_DETECT ( "FALSE" ),
    .AUTORESET_PATTERN_DETECT_OPTINV ( "MATCH" ),
    .A_INPUT ( "DIRECT" ),
    .BCASCREG ( 1 ),
    .BREG ( 1 ),
    .B_INPUT ( "CASCADE" ),
    .CARRYINREG ( 0 ),
    .CARRYINSELREG ( 0 ),
    .CREG ( 0 ),
    .MASK ( 48'h3FFFFFFFFFFF ),
    .MREG ( 1 ),
    .MULTCARRYINREG ( 0 ),
    .OPMODEREG ( 0 ),
    .PATTERN ( 48'h000000000000 ),
    .PREG ( 1 ),
    .SEL_MASK ( "MASK" ),
    .SEL_PATTERN ( "PATTERN" ),
    .SEL_ROUNDING_MASK ( "SEL_MASK" ),
    .SIM_MODE ( "SAFE" ),
    .USE_MULT ( "MULT_S" ),
    .USE_PATTERN_DETECT ( "NO_PATDET" ),
    .USE_SIMD ( "ONE48" ))
  blk00000413 (
    .CEM(ce),
    .CLK(clk),
    .PATTERNBDETECT(NLW_blk00000413_PATTERNBDETECT_UNCONNECTED),
    .RSTC(sig00000461),
    .CEB1(sig00000461),
    .MULTSIGNOUT(NLW_blk00000413_MULTSIGNOUT_UNCONNECTED),
    .CEC(sig00000461),
    .RSTM(sig00000461),
    .MULTSIGNIN(sig00000461),
    .CEB2(ce),
    .RSTCTRL(sig00000461),
    .CEP(ce),
    .CARRYCASCOUT(NLW_blk00000413_CARRYCASCOUT_UNCONNECTED),
    .RSTA(sig00000461),
    .CECARRYIN(sig00000461),
    .UNDERFLOW(NLW_blk00000413_UNDERFLOW_UNCONNECTED),
    .PATTERNDETECT(NLW_blk00000413_PATTERNDETECT_UNCONNECTED),
    .RSTALUMODE(sig00000461),
    .RSTALLCARRYIN(sig00000461),
    .CEALUMODE(sig00000461),
    .CEA2(ce),
    .CEA1(ce),
    .RSTB(sig00000461),
    .CEMULTCARRYIN(sig00000461),
    .OVERFLOW(NLW_blk00000413_OVERFLOW_UNCONNECTED),
    .CECTRL(sig00000461),
    .CARRYIN(sig00000461),
    .CARRYCASCIN(sig00000461),
    .RSTP(sig00000461),
    .CARRYINSEL({sig00000461, sig00000461, sig00000461}),
    .OPMODE({sig00000001, sig00000461, sig00000001, sig00000461, sig00000001, sig00000461, sig00000001}),
    .PCIN({sig00000395, sig00000394, sig00000393, sig00000392, sig00000391, sig00000390, sig0000038f, sig0000038e, sig0000038d, sig0000038c,
sig0000038b, sig0000038a, sig00000389, sig00000388, sig00000387, sig00000386, sig00000385, sig00000384, sig00000383, sig00000382, sig00000381,
sig00000380, sig0000037f, sig0000037e, sig0000037d, sig0000037c, sig0000037b, sig0000037a, sig00000379, sig00000378, sig00000377, sig00000376,
sig00000375, sig00000374, sig00000373, sig00000372, sig00000371, sig00000370, sig0000036f, sig0000036e, sig0000036d, sig0000036c, sig0000036b,
sig0000036a, sig00000369, sig00000368, sig00000367, sig00000366}),
    .BCIN({sig000003a7, sig000003a6, sig000003a5, sig000003a4, sig000003a3, sig000003a2, sig000003a1, sig000003a0, sig0000039f, sig0000039e,
sig0000039d, sig0000039c, sig0000039b, sig0000039a, sig00000399, sig00000398, sig00000397, sig00000396}),
    .A({sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461
, sig00000461, sig00000461, sig00000191, sig00000192, sig00000193, sig00000194, sig00000195, sig00000196, sig00000197, sig00000198, sig00000199,
sig0000019a, sig0000019b, sig0000019c, sig0000019d, sig0000019e, sig0000019f, sig000001a0, sig000001a1}),
    .PCOUT({sig00000363, sig00000362, sig00000361, sig00000360, sig0000035f, sig0000035e, sig0000035d, sig0000035c, sig0000035b, sig0000035a,
sig00000359, sig00000358, sig00000357, sig00000356, sig00000355, sig00000354, sig00000353, sig00000352, sig00000351, sig00000350, sig0000034f,
sig0000034e, sig0000034d, sig0000034c, sig0000034b, sig0000034a, sig00000349, sig00000348, sig00000347, sig00000346, sig00000345, sig00000344,
sig00000343, sig00000342, sig00000341, sig00000340, sig0000033f, sig0000033e, sig0000033d, sig0000033c, sig0000033b, sig0000033a, sig00000339,
sig00000338, sig00000337, sig00000336, sig00000335, sig00000334}),
    .ACOUT({\NLW_blk00000413_ACOUT<29>_UNCONNECTED , \NLW_blk00000413_ACOUT<28>_UNCONNECTED , \NLW_blk00000413_ACOUT<27>_UNCONNECTED ,
\NLW_blk00000413_ACOUT<26>_UNCONNECTED , \NLW_blk00000413_ACOUT<25>_UNCONNECTED , \NLW_blk00000413_ACOUT<24>_UNCONNECTED ,
\NLW_blk00000413_ACOUT<23>_UNCONNECTED , \NLW_blk00000413_ACOUT<22>_UNCONNECTED , \NLW_blk00000413_ACOUT<21>_UNCONNECTED ,
\NLW_blk00000413_ACOUT<20>_UNCONNECTED , \NLW_blk00000413_ACOUT<19>_UNCONNECTED , \NLW_blk00000413_ACOUT<18>_UNCONNECTED ,
\NLW_blk00000413_ACOUT<17>_UNCONNECTED , \NLW_blk00000413_ACOUT<16>_UNCONNECTED , \NLW_blk00000413_ACOUT<15>_UNCONNECTED ,
\NLW_blk00000413_ACOUT<14>_UNCONNECTED , \NLW_blk00000413_ACOUT<13>_UNCONNECTED , \NLW_blk00000413_ACOUT<12>_UNCONNECTED ,
\NLW_blk00000413_ACOUT<11>_UNCONNECTED , \NLW_blk00000413_ACOUT<10>_UNCONNECTED , \NLW_blk00000413_ACOUT<9>_UNCONNECTED ,
\NLW_blk00000413_ACOUT<8>_UNCONNECTED , \NLW_blk00000413_ACOUT<7>_UNCONNECTED , \NLW_blk00000413_ACOUT<6>_UNCONNECTED ,
\NLW_blk00000413_ACOUT<5>_UNCONNECTED , \NLW_blk00000413_ACOUT<4>_UNCONNECTED , \NLW_blk00000413_ACOUT<3>_UNCONNECTED ,
\NLW_blk00000413_ACOUT<2>_UNCONNECTED , \NLW_blk00000413_ACOUT<1>_UNCONNECTED , \NLW_blk00000413_ACOUT<0>_UNCONNECTED }),
    .ALUMODE({sig00000461, sig00000461, sig00000461, sig00000461}),
    .C({sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461
, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461,
sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461,
sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461,
sig00000461, sig00000461, sig00000461, sig00000461}),
    .CARRYOUT({\NLW_blk00000413_CARRYOUT<3>_UNCONNECTED , \NLW_blk00000413_CARRYOUT<2>_UNCONNECTED , \NLW_blk00000413_CARRYOUT<1>_UNCONNECTED ,
\NLW_blk00000413_CARRYOUT<0>_UNCONNECTED }),
    .B({sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461
, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461}),
    .BCOUT({\NLW_blk00000413_BCOUT<17>_UNCONNECTED , \NLW_blk00000413_BCOUT<16>_UNCONNECTED , \NLW_blk00000413_BCOUT<15>_UNCONNECTED ,
\NLW_blk00000413_BCOUT<14>_UNCONNECTED , \NLW_blk00000413_BCOUT<13>_UNCONNECTED , \NLW_blk00000413_BCOUT<12>_UNCONNECTED ,
\NLW_blk00000413_BCOUT<11>_UNCONNECTED , \NLW_blk00000413_BCOUT<10>_UNCONNECTED , \NLW_blk00000413_BCOUT<9>_UNCONNECTED ,
\NLW_blk00000413_BCOUT<8>_UNCONNECTED , \NLW_blk00000413_BCOUT<7>_UNCONNECTED , \NLW_blk00000413_BCOUT<6>_UNCONNECTED ,
\NLW_blk00000413_BCOUT<5>_UNCONNECTED , \NLW_blk00000413_BCOUT<4>_UNCONNECTED , \NLW_blk00000413_BCOUT<3>_UNCONNECTED ,
\NLW_blk00000413_BCOUT<2>_UNCONNECTED , \NLW_blk00000413_BCOUT<1>_UNCONNECTED , \NLW_blk00000413_BCOUT<0>_UNCONNECTED }),
    .P({\NLW_blk00000413_P<47>_UNCONNECTED , \NLW_blk00000413_P<46>_UNCONNECTED , \NLW_blk00000413_P<45>_UNCONNECTED ,
\NLW_blk00000413_P<44>_UNCONNECTED , \NLW_blk00000413_P<43>_UNCONNECTED , \NLW_blk00000413_P<42>_UNCONNECTED , \NLW_blk00000413_P<41>_UNCONNECTED ,
\NLW_blk00000413_P<40>_UNCONNECTED , \NLW_blk00000413_P<39>_UNCONNECTED , \NLW_blk00000413_P<38>_UNCONNECTED , \NLW_blk00000413_P<37>_UNCONNECTED ,
\NLW_blk00000413_P<36>_UNCONNECTED , \NLW_blk00000413_P<35>_UNCONNECTED , \NLW_blk00000413_P<34>_UNCONNECTED , \NLW_blk00000413_P<33>_UNCONNECTED ,
\NLW_blk00000413_P<32>_UNCONNECTED , \NLW_blk00000413_P<31>_UNCONNECTED , \NLW_blk00000413_P<30>_UNCONNECTED , \NLW_blk00000413_P<29>_UNCONNECTED ,
\NLW_blk00000413_P<28>_UNCONNECTED , \NLW_blk00000413_P<27>_UNCONNECTED , \NLW_blk00000413_P<26>_UNCONNECTED , \NLW_blk00000413_P<25>_UNCONNECTED ,
\NLW_blk00000413_P<24>_UNCONNECTED , \NLW_blk00000413_P<23>_UNCONNECTED , \NLW_blk00000413_P<22>_UNCONNECTED , \NLW_blk00000413_P<21>_UNCONNECTED ,
\NLW_blk00000413_P<20>_UNCONNECTED , \NLW_blk00000413_P<19>_UNCONNECTED , \NLW_blk00000413_P<18>_UNCONNECTED , \NLW_blk00000413_P<17>_UNCONNECTED ,
\NLW_blk00000413_P<16>_UNCONNECTED , \NLW_blk00000413_P<15>_UNCONNECTED , \NLW_blk00000413_P<14>_UNCONNECTED , \NLW_blk00000413_P<13>_UNCONNECTED ,
\NLW_blk00000413_P<12>_UNCONNECTED , \NLW_blk00000413_P<11>_UNCONNECTED , \NLW_blk00000413_P<10>_UNCONNECTED , \NLW_blk00000413_P<9>_UNCONNECTED ,
\NLW_blk00000413_P<8>_UNCONNECTED , \NLW_blk00000413_P<7>_UNCONNECTED , \NLW_blk00000413_P<6>_UNCONNECTED , \NLW_blk00000413_P<5>_UNCONNECTED ,
\NLW_blk00000413_P<4>_UNCONNECTED , \NLW_blk00000413_P<3>_UNCONNECTED , \NLW_blk00000413_P<2>_UNCONNECTED , \NLW_blk00000413_P<1>_UNCONNECTED ,
\NLW_blk00000413_P<0>_UNCONNECTED }),
    .ACIN({sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461,
sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461,
sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461})
  );
  DSP48E #(
    .ACASCREG ( 2 ),
    .ALUMODEREG ( 0 ),
    .AREG ( 2 ),
    .AUTORESET_PATTERN_DETECT ( "FALSE" ),
    .AUTORESET_PATTERN_DETECT_OPTINV ( "MATCH" ),
    .A_INPUT ( "DIRECT" ),
    .BCASCREG ( 2 ),
    .BREG ( 2 ),
    .B_INPUT ( "DIRECT" ),
    .CARRYINREG ( 0 ),
    .CARRYINSELREG ( 0 ),
    .CREG ( 0 ),
    .MASK ( 48'hFFFFFFFE0000 ),
    .MREG ( 1 ),
    .MULTCARRYINREG ( 0 ),
    .OPMODEREG ( 0 ),
    .PATTERN ( 48'h000000000000 ),
    .PREG ( 1 ),
    .SEL_MASK ( "MASK" ),
    .SEL_PATTERN ( "PATTERN" ),
    .SEL_ROUNDING_MASK ( "SEL_MASK" ),
    .SIM_MODE ( "SAFE" ),
    .USE_MULT ( "MULT_S" ),
    .USE_PATTERN_DETECT ( "PATDET" ),
    .USE_SIMD ( "ONE48" ))
  blk00000414 (
    .CEM(ce),
    .PATTERNDETECT(sig00000365),
    .CLK(clk),
    .PATTERNBDETECT(NLW_blk00000414_PATTERNBDETECT_UNCONNECTED),
    .RSTC(sig00000461),
    .CEB1(ce),
    .MULTSIGNOUT(NLW_blk00000414_MULTSIGNOUT_UNCONNECTED),
    .CEC(sig00000461),
    .RSTM(sig00000461),
    .MULTSIGNIN(sig00000461),
    .CEB2(ce),
    .RSTCTRL(sig00000461),
    .CEP(ce),
    .CARRYCASCOUT(NLW_blk00000414_CARRYCASCOUT_UNCONNECTED),
    .RSTA(sig00000461),
    .CECARRYIN(sig00000461),
    .UNDERFLOW(NLW_blk00000414_UNDERFLOW_UNCONNECTED),
    .RSTALUMODE(sig00000461),
    .RSTALLCARRYIN(sig00000461),
    .CEALUMODE(sig00000461),
    .CEA2(ce),
    .CEA1(ce),
    .RSTB(sig00000461),
    .CEMULTCARRYIN(sig00000461),
    .OVERFLOW(NLW_blk00000414_OVERFLOW_UNCONNECTED),
    .CECTRL(sig00000461),
    .CARRYIN(sig00000461),
    .CARRYCASCIN(sig00000461),
    .RSTP(sig00000461),
    .CARRYINSEL({sig00000461, sig00000461, sig00000461}),
    .OPMODE({sig00000461, sig00000461, sig00000001, sig00000461, sig00000001, sig00000461, sig00000001}),
    .PCIN({sig000003d7, sig000003d6, sig000003d5, sig000003d4, sig000003d3, sig000003d2, sig000003d1, sig000003d0, sig000003cf, sig000003ce,
sig000003cd, sig000003cc, sig000003cb, sig000003ca, sig000003c9, sig000003c8, sig000003c7, sig000003c6, sig000003c5, sig000003c4, sig000003c3,
sig000003c2, sig000003c1, sig000003c0, sig000003bf, sig000003be, sig000003bd, sig000003bc, sig000003bb, sig000003ba, sig000003b9, sig000003b8,
sig000003b7, sig000003b6, sig000003b5, sig000003b4, sig000003b3, sig000003b2, sig000003b1, sig000003b0, sig000003af, sig000003ae, sig000003ad,
sig000003ac, sig000003ab, sig000003aa, sig000003a9, sig000003a8}),
    .B({sig00000461, sig000001b4, sig000001b5, sig000001b6, sig000001b7, sig000001b8, sig000001b9, sig000001ba, sig000001bb, sig000001bc, sig000001bd
, sig000001be, sig000001bf, sig000001c0, sig000001c1, sig000001c2, sig000001c3, sig000001c4}),
    .BCOUT({sig000003a7, sig000003a6, sig000003a5, sig000003a4, sig000003a3, sig000003a2, sig000003a1, sig000003a0, sig0000039f, sig0000039e,
sig0000039d, sig0000039c, sig0000039b, sig0000039a, sig00000399, sig00000398, sig00000397, sig00000396}),
    .A({sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461
, sig00000461, sig00000461, sig000001a3, sig000001a4, sig000001a5, sig000001a6, sig000001a7, sig000001a8, sig000001a9, sig000001aa, sig000001ab,
sig000001ac, sig000001ad, sig000001ae, sig000001af, sig000001b0, sig000001b1, sig000001b2, sig000001b3}),
    .PCOUT({sig00000395, sig00000394, sig00000393, sig00000392, sig00000391, sig00000390, sig0000038f, sig0000038e, sig0000038d, sig0000038c,
sig0000038b, sig0000038a, sig00000389, sig00000388, sig00000387, sig00000386, sig00000385, sig00000384, sig00000383, sig00000382, sig00000381,
sig00000380, sig0000037f, sig0000037e, sig0000037d, sig0000037c, sig0000037b, sig0000037a, sig00000379, sig00000378, sig00000377, sig00000376,
sig00000375, sig00000374, sig00000373, sig00000372, sig00000371, sig00000370, sig0000036f, sig0000036e, sig0000036d, sig0000036c, sig0000036b,
sig0000036a, sig00000369, sig00000368, sig00000367, sig00000366}),
    .ACOUT({\NLW_blk00000414_ACOUT<29>_UNCONNECTED , \NLW_blk00000414_ACOUT<28>_UNCONNECTED , \NLW_blk00000414_ACOUT<27>_UNCONNECTED ,
\NLW_blk00000414_ACOUT<26>_UNCONNECTED , \NLW_blk00000414_ACOUT<25>_UNCONNECTED , \NLW_blk00000414_ACOUT<24>_UNCONNECTED ,
\NLW_blk00000414_ACOUT<23>_UNCONNECTED , \NLW_blk00000414_ACOUT<22>_UNCONNECTED , \NLW_blk00000414_ACOUT<21>_UNCONNECTED ,
\NLW_blk00000414_ACOUT<20>_UNCONNECTED , \NLW_blk00000414_ACOUT<19>_UNCONNECTED , \NLW_blk00000414_ACOUT<18>_UNCONNECTED ,
\NLW_blk00000414_ACOUT<17>_UNCONNECTED , \NLW_blk00000414_ACOUT<16>_UNCONNECTED , \NLW_blk00000414_ACOUT<15>_UNCONNECTED ,
\NLW_blk00000414_ACOUT<14>_UNCONNECTED , \NLW_blk00000414_ACOUT<13>_UNCONNECTED , \NLW_blk00000414_ACOUT<12>_UNCONNECTED ,
\NLW_blk00000414_ACOUT<11>_UNCONNECTED , \NLW_blk00000414_ACOUT<10>_UNCONNECTED , \NLW_blk00000414_ACOUT<9>_UNCONNECTED ,
\NLW_blk00000414_ACOUT<8>_UNCONNECTED , \NLW_blk00000414_ACOUT<7>_UNCONNECTED , \NLW_blk00000414_ACOUT<6>_UNCONNECTED ,
\NLW_blk00000414_ACOUT<5>_UNCONNECTED , \NLW_blk00000414_ACOUT<4>_UNCONNECTED , \NLW_blk00000414_ACOUT<3>_UNCONNECTED ,
\NLW_blk00000414_ACOUT<2>_UNCONNECTED , \NLW_blk00000414_ACOUT<1>_UNCONNECTED , \NLW_blk00000414_ACOUT<0>_UNCONNECTED }),
    .ALUMODE({sig00000461, sig00000461, sig00000461, sig00000461}),
    .C({sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461
, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461,
sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461,
sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461,
sig00000461, sig00000461, sig00000461, sig00000461}),
    .CARRYOUT({\NLW_blk00000414_CARRYOUT<3>_UNCONNECTED , \NLW_blk00000414_CARRYOUT<2>_UNCONNECTED , \NLW_blk00000414_CARRYOUT<1>_UNCONNECTED ,
\NLW_blk00000414_CARRYOUT<0>_UNCONNECTED }),
    .BCIN({sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461,
sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461}),
    .P({\NLW_blk00000414_P<47>_UNCONNECTED , \NLW_blk00000414_P<46>_UNCONNECTED , \NLW_blk00000414_P<45>_UNCONNECTED ,
\NLW_blk00000414_P<44>_UNCONNECTED , \NLW_blk00000414_P<43>_UNCONNECTED , \NLW_blk00000414_P<42>_UNCONNECTED , \NLW_blk00000414_P<41>_UNCONNECTED ,
\NLW_blk00000414_P<40>_UNCONNECTED , \NLW_blk00000414_P<39>_UNCONNECTED , \NLW_blk00000414_P<38>_UNCONNECTED , \NLW_blk00000414_P<37>_UNCONNECTED ,
\NLW_blk00000414_P<36>_UNCONNECTED , \NLW_blk00000414_P<35>_UNCONNECTED , \NLW_blk00000414_P<34>_UNCONNECTED , \NLW_blk00000414_P<33>_UNCONNECTED ,
\NLW_blk00000414_P<32>_UNCONNECTED , \NLW_blk00000414_P<31>_UNCONNECTED , \NLW_blk00000414_P<30>_UNCONNECTED , \NLW_blk00000414_P<29>_UNCONNECTED ,
\NLW_blk00000414_P<28>_UNCONNECTED , \NLW_blk00000414_P<27>_UNCONNECTED , \NLW_blk00000414_P<26>_UNCONNECTED , \NLW_blk00000414_P<25>_UNCONNECTED ,
\NLW_blk00000414_P<24>_UNCONNECTED , \NLW_blk00000414_P<23>_UNCONNECTED , \NLW_blk00000414_P<22>_UNCONNECTED , \NLW_blk00000414_P<21>_UNCONNECTED ,
\NLW_blk00000414_P<20>_UNCONNECTED , \NLW_blk00000414_P<19>_UNCONNECTED , \NLW_blk00000414_P<18>_UNCONNECTED , \NLW_blk00000414_P<17>_UNCONNECTED ,
\NLW_blk00000414_P<16>_UNCONNECTED , \NLW_blk00000414_P<15>_UNCONNECTED , \NLW_blk00000414_P<14>_UNCONNECTED , \NLW_blk00000414_P<13>_UNCONNECTED ,
\NLW_blk00000414_P<12>_UNCONNECTED , \NLW_blk00000414_P<11>_UNCONNECTED , \NLW_blk00000414_P<10>_UNCONNECTED , \NLW_blk00000414_P<9>_UNCONNECTED ,
\NLW_blk00000414_P<8>_UNCONNECTED , \NLW_blk00000414_P<7>_UNCONNECTED , \NLW_blk00000414_P<6>_UNCONNECTED , \NLW_blk00000414_P<5>_UNCONNECTED ,
\NLW_blk00000414_P<4>_UNCONNECTED , \NLW_blk00000414_P<3>_UNCONNECTED , \NLW_blk00000414_P<2>_UNCONNECTED , \NLW_blk00000414_P<1>_UNCONNECTED ,
\NLW_blk00000414_P<0>_UNCONNECTED }),
    .ACIN({sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461,
sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461,
sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461})
  );
  DSP48E #(
    .ACASCREG ( 2 ),
    .ALUMODEREG ( 0 ),
    .AREG ( 2 ),
    .AUTORESET_PATTERN_DETECT ( "FALSE" ),
    .AUTORESET_PATTERN_DETECT_OPTINV ( "MATCH" ),
    .A_INPUT ( "DIRECT" ),
    .BCASCREG ( 1 ),
    .BREG ( 1 ),
    .B_INPUT ( "CASCADE" ),
    .CARRYINREG ( 0 ),
    .CARRYINSELREG ( 0 ),
    .CREG ( 0 ),
    .MASK ( 48'h3FFFFFFFFFFF ),
    .MREG ( 1 ),
    .MULTCARRYINREG ( 0 ),
    .OPMODEREG ( 0 ),
    .PATTERN ( 48'h000000000000 ),
    .PREG ( 1 ),
    .SEL_MASK ( "MASK" ),
    .SEL_PATTERN ( "PATTERN" ),
    .SEL_ROUNDING_MASK ( "SEL_MASK" ),
    .SIM_MODE ( "SAFE" ),
    .USE_MULT ( "MULT_S" ),
    .USE_PATTERN_DETECT ( "NO_PATDET" ),
    .USE_SIMD ( "ONE48" ))
  blk00000415 (
    .CEM(ce),
    .CLK(clk),
    .PATTERNBDETECT(NLW_blk00000415_PATTERNBDETECT_UNCONNECTED),
    .RSTC(sig00000461),
    .CEB1(sig00000461),
    .MULTSIGNOUT(NLW_blk00000415_MULTSIGNOUT_UNCONNECTED),
    .CEC(sig00000461),
    .RSTM(sig00000461),
    .MULTSIGNIN(sig00000461),
    .CEB2(ce),
    .RSTCTRL(sig00000461),
    .CEP(ce),
    .CARRYCASCOUT(NLW_blk00000415_CARRYCASCOUT_UNCONNECTED),
    .RSTA(sig00000461),
    .CECARRYIN(sig00000461),
    .UNDERFLOW(NLW_blk00000415_UNDERFLOW_UNCONNECTED),
    .PATTERNDETECT(NLW_blk00000415_PATTERNDETECT_UNCONNECTED),
    .RSTALUMODE(sig00000461),
    .RSTALLCARRYIN(sig00000461),
    .CEALUMODE(sig00000461),
    .CEA2(ce),
    .CEA1(ce),
    .RSTB(sig00000461),
    .CEMULTCARRYIN(sig00000461),
    .OVERFLOW(NLW_blk00000415_OVERFLOW_UNCONNECTED),
    .CECTRL(sig00000461),
    .CARRYIN(sig00000461),
    .CARRYCASCIN(sig00000461),
    .RSTP(sig00000461),
    .CARRYINSEL({sig00000461, sig00000461, sig00000461}),
    .OPMODE({sig00000001, sig00000461, sig00000001, sig00000461, sig00000001, sig00000461, sig00000001}),
    .PCIN({sig00000409, sig00000408, sig00000407, sig00000406, sig00000405, sig00000404, sig00000403, sig00000402, sig00000401, sig00000400,
sig000003ff, sig000003fe, sig000003fd, sig000003fc, sig000003fb, sig000003fa, sig000003f9, sig000003f8, sig000003f7, sig000003f6, sig000003f5,
sig000003f4, sig000003f3, sig000003f2, sig000003f1, sig000003f0, sig000003ef, sig000003ee, sig000003ed, sig000003ec, sig000003eb, sig000003ea,
sig000003e9, sig000003e8, sig000003e7, sig000003e6, sig000003e5, sig000003e4, sig000003e3, sig000003e2, sig000003e1, sig000003e0, sig000003df,
sig000003de, sig000003dd, sig000003dc, sig000003db, sig000003da}),
    .BCIN({sig0000041b, sig0000041a, sig00000419, sig00000418, sig00000417, sig00000416, sig00000415, sig00000414, sig00000413, sig00000412,
sig00000411, sig00000410, sig0000040f, sig0000040e, sig0000040d, sig0000040c, sig0000040b, sig0000040a}),
    .A({sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461
, sig00000461, sig00000461, a[33], a[32], a[31], a[30], a[29], a[28], a[27], a[26], a[25], a[24], a[23], a[22], a[21], a[20], a[19], a[18], a[17]}),
    .PCOUT({sig000003d7, sig000003d6, sig000003d5, sig000003d4, sig000003d3, sig000003d2, sig000003d1, sig000003d0, sig000003cf, sig000003ce,
sig000003cd, sig000003cc, sig000003cb, sig000003ca, sig000003c9, sig000003c8, sig000003c7, sig000003c6, sig000003c5, sig000003c4, sig000003c3,
sig000003c2, sig000003c1, sig000003c0, sig000003bf, sig000003be, sig000003bd, sig000003bc, sig000003bb, sig000003ba, sig000003b9, sig000003b8,
sig000003b7, sig000003b6, sig000003b5, sig000003b4, sig000003b3, sig000003b2, sig000003b1, sig000003b0, sig000003af, sig000003ae, sig000003ad,
sig000003ac, sig000003ab, sig000003aa, sig000003a9, sig000003a8}),
    .ACOUT({\NLW_blk00000415_ACOUT<29>_UNCONNECTED , \NLW_blk00000415_ACOUT<28>_UNCONNECTED , \NLW_blk00000415_ACOUT<27>_UNCONNECTED ,
\NLW_blk00000415_ACOUT<26>_UNCONNECTED , \NLW_blk00000415_ACOUT<25>_UNCONNECTED , \NLW_blk00000415_ACOUT<24>_UNCONNECTED ,
\NLW_blk00000415_ACOUT<23>_UNCONNECTED , \NLW_blk00000415_ACOUT<22>_UNCONNECTED , \NLW_blk00000415_ACOUT<21>_UNCONNECTED ,
\NLW_blk00000415_ACOUT<20>_UNCONNECTED , \NLW_blk00000415_ACOUT<19>_UNCONNECTED , \NLW_blk00000415_ACOUT<18>_UNCONNECTED ,
\NLW_blk00000415_ACOUT<17>_UNCONNECTED , \NLW_blk00000415_ACOUT<16>_UNCONNECTED , \NLW_blk00000415_ACOUT<15>_UNCONNECTED ,
\NLW_blk00000415_ACOUT<14>_UNCONNECTED , \NLW_blk00000415_ACOUT<13>_UNCONNECTED , \NLW_blk00000415_ACOUT<12>_UNCONNECTED ,
\NLW_blk00000415_ACOUT<11>_UNCONNECTED , \NLW_blk00000415_ACOUT<10>_UNCONNECTED , \NLW_blk00000415_ACOUT<9>_UNCONNECTED ,
\NLW_blk00000415_ACOUT<8>_UNCONNECTED , \NLW_blk00000415_ACOUT<7>_UNCONNECTED , \NLW_blk00000415_ACOUT<6>_UNCONNECTED ,
\NLW_blk00000415_ACOUT<5>_UNCONNECTED , \NLW_blk00000415_ACOUT<4>_UNCONNECTED , \NLW_blk00000415_ACOUT<3>_UNCONNECTED ,
\NLW_blk00000415_ACOUT<2>_UNCONNECTED , \NLW_blk00000415_ACOUT<1>_UNCONNECTED , \NLW_blk00000415_ACOUT<0>_UNCONNECTED }),
    .ALUMODE({sig00000461, sig00000461, sig00000461, sig00000461}),
    .C({sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461
, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461,
sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461,
sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461,
sig00000461, sig00000461, sig00000461, sig00000461}),
    .CARRYOUT({\NLW_blk00000415_CARRYOUT<3>_UNCONNECTED , \NLW_blk00000415_CARRYOUT<2>_UNCONNECTED , \NLW_blk00000415_CARRYOUT<1>_UNCONNECTED ,
\NLW_blk00000415_CARRYOUT<0>_UNCONNECTED }),
    .B({sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461
, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461}),
    .BCOUT({\NLW_blk00000415_BCOUT<17>_UNCONNECTED , \NLW_blk00000415_BCOUT<16>_UNCONNECTED , \NLW_blk00000415_BCOUT<15>_UNCONNECTED ,
\NLW_blk00000415_BCOUT<14>_UNCONNECTED , \NLW_blk00000415_BCOUT<13>_UNCONNECTED , \NLW_blk00000415_BCOUT<12>_UNCONNECTED ,
\NLW_blk00000415_BCOUT<11>_UNCONNECTED , \NLW_blk00000415_BCOUT<10>_UNCONNECTED , \NLW_blk00000415_BCOUT<9>_UNCONNECTED ,
\NLW_blk00000415_BCOUT<8>_UNCONNECTED , \NLW_blk00000415_BCOUT<7>_UNCONNECTED , \NLW_blk00000415_BCOUT<6>_UNCONNECTED ,
\NLW_blk00000415_BCOUT<5>_UNCONNECTED , \NLW_blk00000415_BCOUT<4>_UNCONNECTED , \NLW_blk00000415_BCOUT<3>_UNCONNECTED ,
\NLW_blk00000415_BCOUT<2>_UNCONNECTED , \NLW_blk00000415_BCOUT<1>_UNCONNECTED , \NLW_blk00000415_BCOUT<0>_UNCONNECTED }),
    .P({\NLW_blk00000415_P<47>_UNCONNECTED , \NLW_blk00000415_P<46>_UNCONNECTED , \NLW_blk00000415_P<45>_UNCONNECTED ,
\NLW_blk00000415_P<44>_UNCONNECTED , \NLW_blk00000415_P<43>_UNCONNECTED , \NLW_blk00000415_P<42>_UNCONNECTED , \NLW_blk00000415_P<41>_UNCONNECTED ,
\NLW_blk00000415_P<40>_UNCONNECTED , \NLW_blk00000415_P<39>_UNCONNECTED , \NLW_blk00000415_P<38>_UNCONNECTED , \NLW_blk00000415_P<37>_UNCONNECTED ,
\NLW_blk00000415_P<36>_UNCONNECTED , \NLW_blk00000415_P<35>_UNCONNECTED , \NLW_blk00000415_P<34>_UNCONNECTED , \NLW_blk00000415_P<33>_UNCONNECTED ,
\NLW_blk00000415_P<32>_UNCONNECTED , \NLW_blk00000415_P<31>_UNCONNECTED , \NLW_blk00000415_P<30>_UNCONNECTED , \NLW_blk00000415_P<29>_UNCONNECTED ,
\NLW_blk00000415_P<28>_UNCONNECTED , \NLW_blk00000415_P<27>_UNCONNECTED , \NLW_blk00000415_P<26>_UNCONNECTED , \NLW_blk00000415_P<25>_UNCONNECTED ,
\NLW_blk00000415_P<24>_UNCONNECTED , \NLW_blk00000415_P<23>_UNCONNECTED , \NLW_blk00000415_P<22>_UNCONNECTED , \NLW_blk00000415_P<21>_UNCONNECTED ,
\NLW_blk00000415_P<20>_UNCONNECTED , \NLW_blk00000415_P<19>_UNCONNECTED , \NLW_blk00000415_P<18>_UNCONNECTED , \NLW_blk00000415_P<17>_UNCONNECTED ,
\NLW_blk00000415_P<16>_UNCONNECTED , \NLW_blk00000415_P<15>_UNCONNECTED , \NLW_blk00000415_P<14>_UNCONNECTED , \NLW_blk00000415_P<13>_UNCONNECTED ,
\NLW_blk00000415_P<12>_UNCONNECTED , \NLW_blk00000415_P<11>_UNCONNECTED , \NLW_blk00000415_P<10>_UNCONNECTED , \NLW_blk00000415_P<9>_UNCONNECTED ,
\NLW_blk00000415_P<8>_UNCONNECTED , \NLW_blk00000415_P<7>_UNCONNECTED , \NLW_blk00000415_P<6>_UNCONNECTED , \NLW_blk00000415_P<5>_UNCONNECTED ,
\NLW_blk00000415_P<4>_UNCONNECTED , \NLW_blk00000415_P<3>_UNCONNECTED , \NLW_blk00000415_P<2>_UNCONNECTED , \NLW_blk00000415_P<1>_UNCONNECTED ,
\NLW_blk00000415_P<0>_UNCONNECTED }),
    .ACIN({sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461,
sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461,
sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461})
  );
  DSP48E #(
    .ACASCREG ( 1 ),
    .ALUMODEREG ( 0 ),
    .AREG ( 1 ),
    .AUTORESET_PATTERN_DETECT ( "FALSE" ),
    .AUTORESET_PATTERN_DETECT_OPTINV ( "MATCH" ),
    .A_INPUT ( "DIRECT" ),
    .BCASCREG ( 1 ),
    .BREG ( 1 ),
    .B_INPUT ( "DIRECT" ),
    .CARRYINREG ( 0 ),
    .CARRYINSELREG ( 0 ),
    .CREG ( 0 ),
    .MASK ( 48'hFFFFFFFE0000 ),
    .MREG ( 1 ),
    .MULTCARRYINREG ( 0 ),
    .OPMODEREG ( 0 ),
    .PATTERN ( 48'h000000000000 ),
    .PREG ( 1 ),
    .SEL_MASK ( "MASK" ),
    .SEL_PATTERN ( "PATTERN" ),
    .SEL_ROUNDING_MASK ( "SEL_MASK" ),
    .SIM_MODE ( "SAFE" ),
    .USE_MULT ( "MULT_S" ),
    .USE_PATTERN_DETECT ( "PATDET" ),
    .USE_SIMD ( "ONE48" ))
  blk00000416 (
    .CEM(ce),
    .PATTERNDETECT(sig000003d9),
    .CLK(clk),
    .PATTERNBDETECT(NLW_blk00000416_PATTERNBDETECT_UNCONNECTED),
    .RSTC(sig00000461),
    .CEB1(sig00000461),
    .MULTSIGNOUT(NLW_blk00000416_MULTSIGNOUT_UNCONNECTED),
    .CEC(sig00000461),
    .RSTM(sig00000461),
    .MULTSIGNIN(sig00000461),
    .CEB2(ce),
    .RSTCTRL(sig00000461),
    .CEP(ce),
    .CARRYCASCOUT(NLW_blk00000416_CARRYCASCOUT_UNCONNECTED),
    .RSTA(sig00000461),
    .CECARRYIN(sig00000461),
    .UNDERFLOW(NLW_blk00000416_UNDERFLOW_UNCONNECTED),
    .RSTALUMODE(sig00000461),
    .RSTALLCARRYIN(sig00000461),
    .CEALUMODE(sig00000461),
    .CEA2(ce),
    .CEA1(sig00000461),
    .RSTB(sig00000461),
    .CEMULTCARRYIN(sig00000461),
    .OVERFLOW(NLW_blk00000416_OVERFLOW_UNCONNECTED),
    .CECTRL(sig00000461),
    .CARRYIN(sig00000461),
    .CARRYCASCIN(sig00000461),
    .RSTP(sig00000461),
    .CARRYINSEL({sig00000461, sig00000461, sig00000461}),
    .OPMODE({sig00000461, sig00000461, sig00000461, sig00000461, sig00000001, sig00000461, sig00000001}),
    .B({sig00000461, b[16], b[15], b[14], b[13], b[12], b[11], b[10], b[9], b[8], b[7], b[6], b[5], b[4], b[3], b[2], b[1], b[0]}),
    .BCOUT({sig0000041b, sig0000041a, sig00000419, sig00000418, sig00000417, sig00000416, sig00000415, sig00000414, sig00000413, sig00000412,
sig00000411, sig00000410, sig0000040f, sig0000040e, sig0000040d, sig0000040c, sig0000040b, sig0000040a}),
    .A({sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461
, sig00000461, sig00000461, a[16], a[15], a[14], a[13], a[12], a[11], a[10], a[9], a[8], a[7], a[6], a[5], a[4], a[3], a[2], a[1], a[0]}),
    .PCOUT({sig00000409, sig00000408, sig00000407, sig00000406, sig00000405, sig00000404, sig00000403, sig00000402, sig00000401, sig00000400,
sig000003ff, sig000003fe, sig000003fd, sig000003fc, sig000003fb, sig000003fa, sig000003f9, sig000003f8, sig000003f7, sig000003f6, sig000003f5,
sig000003f4, sig000003f3, sig000003f2, sig000003f1, sig000003f0, sig000003ef, sig000003ee, sig000003ed, sig000003ec, sig000003eb, sig000003ea,
sig000003e9, sig000003e8, sig000003e7, sig000003e6, sig000003e5, sig000003e4, sig000003e3, sig000003e2, sig000003e1, sig000003e0, sig000003df,
sig000003de, sig000003dd, sig000003dc, sig000003db, sig000003da}),
    .ACOUT({\NLW_blk00000416_ACOUT<29>_UNCONNECTED , \NLW_blk00000416_ACOUT<28>_UNCONNECTED , \NLW_blk00000416_ACOUT<27>_UNCONNECTED ,
\NLW_blk00000416_ACOUT<26>_UNCONNECTED , \NLW_blk00000416_ACOUT<25>_UNCONNECTED , \NLW_blk00000416_ACOUT<24>_UNCONNECTED ,
\NLW_blk00000416_ACOUT<23>_UNCONNECTED , \NLW_blk00000416_ACOUT<22>_UNCONNECTED , \NLW_blk00000416_ACOUT<21>_UNCONNECTED ,
\NLW_blk00000416_ACOUT<20>_UNCONNECTED , \NLW_blk00000416_ACOUT<19>_UNCONNECTED , \NLW_blk00000416_ACOUT<18>_UNCONNECTED ,
\NLW_blk00000416_ACOUT<17>_UNCONNECTED , \NLW_blk00000416_ACOUT<16>_UNCONNECTED , \NLW_blk00000416_ACOUT<15>_UNCONNECTED ,
\NLW_blk00000416_ACOUT<14>_UNCONNECTED , \NLW_blk00000416_ACOUT<13>_UNCONNECTED , \NLW_blk00000416_ACOUT<12>_UNCONNECTED ,
\NLW_blk00000416_ACOUT<11>_UNCONNECTED , \NLW_blk00000416_ACOUT<10>_UNCONNECTED , \NLW_blk00000416_ACOUT<9>_UNCONNECTED ,
\NLW_blk00000416_ACOUT<8>_UNCONNECTED , \NLW_blk00000416_ACOUT<7>_UNCONNECTED , \NLW_blk00000416_ACOUT<6>_UNCONNECTED ,
\NLW_blk00000416_ACOUT<5>_UNCONNECTED , \NLW_blk00000416_ACOUT<4>_UNCONNECTED , \NLW_blk00000416_ACOUT<3>_UNCONNECTED ,
\NLW_blk00000416_ACOUT<2>_UNCONNECTED , \NLW_blk00000416_ACOUT<1>_UNCONNECTED , \NLW_blk00000416_ACOUT<0>_UNCONNECTED }),
    .PCIN({sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461,
sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461,
sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461,
sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461,
sig00000461, sig00000461, sig00000461, sig00000461, sig00000461}),
    .ALUMODE({sig00000461, sig00000461, sig00000461, sig00000461}),
    .C({sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461
, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461,
sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461,
sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461,
sig00000461, sig00000461, sig00000461, sig00000461}),
    .CARRYOUT({\NLW_blk00000416_CARRYOUT<3>_UNCONNECTED , \NLW_blk00000416_CARRYOUT<2>_UNCONNECTED , \NLW_blk00000416_CARRYOUT<1>_UNCONNECTED ,
\NLW_blk00000416_CARRYOUT<0>_UNCONNECTED }),
    .BCIN({sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461,
sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461}),
    .P({\NLW_blk00000416_P<47>_UNCONNECTED , \NLW_blk00000416_P<46>_UNCONNECTED , \NLW_blk00000416_P<45>_UNCONNECTED ,
\NLW_blk00000416_P<44>_UNCONNECTED , \NLW_blk00000416_P<43>_UNCONNECTED , \NLW_blk00000416_P<42>_UNCONNECTED , \NLW_blk00000416_P<41>_UNCONNECTED ,
\NLW_blk00000416_P<40>_UNCONNECTED , \NLW_blk00000416_P<39>_UNCONNECTED , \NLW_blk00000416_P<38>_UNCONNECTED , \NLW_blk00000416_P<37>_UNCONNECTED ,
\NLW_blk00000416_P<36>_UNCONNECTED , \NLW_blk00000416_P<35>_UNCONNECTED , \NLW_blk00000416_P<34>_UNCONNECTED , \NLW_blk00000416_P<33>_UNCONNECTED ,
\NLW_blk00000416_P<32>_UNCONNECTED , \NLW_blk00000416_P<31>_UNCONNECTED , \NLW_blk00000416_P<30>_UNCONNECTED , \NLW_blk00000416_P<29>_UNCONNECTED ,
\NLW_blk00000416_P<28>_UNCONNECTED , \NLW_blk00000416_P<27>_UNCONNECTED , \NLW_blk00000416_P<26>_UNCONNECTED , \NLW_blk00000416_P<25>_UNCONNECTED ,
\NLW_blk00000416_P<24>_UNCONNECTED , \NLW_blk00000416_P<23>_UNCONNECTED , \NLW_blk00000416_P<22>_UNCONNECTED , \NLW_blk00000416_P<21>_UNCONNECTED ,
\NLW_blk00000416_P<20>_UNCONNECTED , \NLW_blk00000416_P<19>_UNCONNECTED , \NLW_blk00000416_P<18>_UNCONNECTED , \NLW_blk00000416_P<17>_UNCONNECTED ,
\NLW_blk00000416_P<16>_UNCONNECTED , \NLW_blk00000416_P<15>_UNCONNECTED , \NLW_blk00000416_P<14>_UNCONNECTED , \NLW_blk00000416_P<13>_UNCONNECTED ,
\NLW_blk00000416_P<12>_UNCONNECTED , \NLW_blk00000416_P<11>_UNCONNECTED , \NLW_blk00000416_P<10>_UNCONNECTED , \NLW_blk00000416_P<9>_UNCONNECTED ,
\NLW_blk00000416_P<8>_UNCONNECTED , \NLW_blk00000416_P<7>_UNCONNECTED , \NLW_blk00000416_P<6>_UNCONNECTED , \NLW_blk00000416_P<5>_UNCONNECTED ,
\NLW_blk00000416_P<4>_UNCONNECTED , \NLW_blk00000416_P<3>_UNCONNECTED , \NLW_blk00000416_P<2>_UNCONNECTED , \NLW_blk00000416_P<1>_UNCONNECTED ,
\NLW_blk00000416_P<0>_UNCONNECTED }),
    .ACIN({sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461,
sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461,
sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461, sig00000461})
  );
// synthesis translate_on
endmodule