module works only with 16/32/64 gtx input data width");
            $finish;
        end
endgenerate
// set data outputs to gtx
assign  txdata_out    = txdata;
assign  txcharisk_out = txcharisk;
*/
endmodule