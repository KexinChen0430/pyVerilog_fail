module outputs
  wire [63 : 0] slave_rdata;
  wire [3 : 0] slave_bid, slave_rid;
  wire [1 : 0] slave_bresp, slave_rresp;
  wire RDY_set_addr_map,
       slave_arready,
       slave_awready,
       slave_bvalid,
       slave_rlast,
       slave_rvalid,
       slave_wready;
  // register rg_addr_base
  reg [63 : 0] rg_addr_base;
  wire [63 : 0] rg_addr_base$D_IN;
  wire rg_addr_base$EN;
  // register rg_addr_lim
  reg [63 : 0] rg_addr_lim;
  wire [63 : 0] rg_addr_lim$D_IN;
  wire rg_addr_lim$EN;
  // register rg_module_ready
  reg rg_module_ready;
  wire rg_module_ready$D_IN, rg_module_ready$EN;
  // ports of submodule slave_xactor_f_rd_addr
  wire [96 : 0] slave_xactor_f_rd_addr$D_IN, slave_xactor_f_rd_addr$D_OUT;
  wire slave_xactor_f_rd_addr$CLR,
       slave_xactor_f_rd_addr$DEQ,
       slave_xactor_f_rd_addr$EMPTY_N,
       slave_xactor_f_rd_addr$ENQ,
       slave_xactor_f_rd_addr$FULL_N;
  // ports of submodule slave_xactor_f_rd_data
  wire [70 : 0] slave_xactor_f_rd_data$D_IN, slave_xactor_f_rd_data$D_OUT;
  wire slave_xactor_f_rd_data$CLR,
       slave_xactor_f_rd_data$DEQ,
       slave_xactor_f_rd_data$EMPTY_N,
       slave_xactor_f_rd_data$ENQ,
       slave_xactor_f_rd_data$FULL_N;
  // ports of submodule slave_xactor_f_wr_addr
  wire [96 : 0] slave_xactor_f_wr_addr$D_IN, slave_xactor_f_wr_addr$D_OUT;
  wire slave_xactor_f_wr_addr$CLR,
       slave_xactor_f_wr_addr$DEQ,
       slave_xactor_f_wr_addr$EMPTY_N,
       slave_xactor_f_wr_addr$ENQ,
       slave_xactor_f_wr_addr$FULL_N;
  // ports of submodule slave_xactor_f_wr_data
  wire [72 : 0] slave_xactor_f_wr_data$D_IN;
  wire slave_xactor_f_wr_data$CLR,
       slave_xactor_f_wr_data$DEQ,
       slave_xactor_f_wr_data$EMPTY_N,
       slave_xactor_f_wr_data$ENQ,
       slave_xactor_f_wr_data$FULL_N;
  // ports of submodule slave_xactor_f_wr_resp
  wire [5 : 0] slave_xactor_f_wr_resp$D_IN, slave_xactor_f_wr_resp$D_OUT;
  wire slave_xactor_f_wr_resp$CLR,
       slave_xactor_f_wr_resp$DEQ,
       slave_xactor_f_wr_resp$EMPTY_N,
       slave_xactor_f_wr_resp$ENQ,
       slave_xactor_f_wr_resp$FULL_N;
  // rule scheduling signals
  wire CAN_FIRE_RL_rl_process_rd_req,
       CAN_FIRE_RL_rl_process_wr_req,
       CAN_FIRE_set_addr_map,
       CAN_FIRE_slave_m_arvalid,
       CAN_FIRE_slave_m_awvalid,
       CAN_FIRE_slave_m_bready,
       CAN_FIRE_slave_m_rready,
       CAN_FIRE_slave_m_wvalid,
       WILL_FIRE_RL_rl_process_rd_req,
       WILL_FIRE_RL_rl_process_wr_req,
       WILL_FIRE_set_addr_map,
       WILL_FIRE_slave_m_arvalid,
       WILL_FIRE_slave_m_awvalid,
       WILL_FIRE_slave_m_bready,
       WILL_FIRE_slave_m_rready,
       WILL_FIRE_slave_m_wvalid;
  // declarations used by system tasks
  // synopsys translate_off
  reg [31 : 0] v__h808;
  reg [31 : 0] v__h8925;
  reg [31 : 0] v__h9218;
  reg [31 : 0] v__h9328;
  reg [31 : 0] v__h802;
  reg [31 : 0] v__h8919;
  reg [31 : 0] v__h9212;
  reg [31 : 0] v__h9322;
  // synopsys translate_on
  // remaining internal signals
  reg [63 : 0] data64__h987;
  reg [31 : 0] CASE_byte_addr05_16_0x0_24_0x0_32_0x54040000_4_ETC__q1,
	       CASE_byte_addr05_16_0x28067_24_0x80000000_32_0_ETC__q2;
  wire [63 : 0] byte_addr__h705, rdata__h924;
  wire [1 : 0] rdr_rresp__h957;
  wire NOT_slave_xactor_f_rd_addr_first_BITS_31_TO_29_ETC___d18,
       NOT_slave_xactor_f_wr_addr_first__208_BITS_31__ETC___d1218;
  // action method set_addr_map
  assign RDY_set_addr_map = 1'd1 ;
  assign CAN_FIRE_set_addr_map = 1'd1 ;
  assign WILL_FIRE_set_addr_map = EN_set_addr_map ;
  // action method slave_m_awvalid
  assign CAN_FIRE_slave_m_awvalid = 1'd1 ;
  assign WILL_FIRE_slave_m_awvalid = 1'd1 ;
  // value method slave_m_awready
  assign slave_awready = slave_xactor_f_wr_addr$FULL_N ;
  // action method slave_m_wvalid
  assign CAN_FIRE_slave_m_wvalid = 1'd1 ;
  assign WILL_FIRE_slave_m_wvalid = 1'd1 ;
  // value method slave_m_wready
  assign slave_wready = slave_xactor_f_wr_data$FULL_N ;
  // value method slave_m_bvalid
  assign slave_bvalid = slave_xactor_f_wr_resp$EMPTY_N ;
  // value method slave_m_bid
  assign slave_bid = slave_xactor_f_wr_resp$D_OUT[5:2] ;
  // value method slave_m_bresp
  assign slave_bresp = slave_xactor_f_wr_resp$D_OUT[1:0] ;
  // action method slave_m_bready
  assign CAN_FIRE_slave_m_bready = 1'd1 ;
  assign WILL_FIRE_slave_m_bready = 1'd1 ;
  // action method slave_m_arvalid
  assign CAN_FIRE_slave_m_arvalid = 1'd1 ;
  assign WILL_FIRE_slave_m_arvalid = 1'd1 ;
  // value method slave_m_arready
  assign slave_arready = slave_xactor_f_rd_addr$FULL_N ;
  // value method slave_m_rvalid
  assign slave_rvalid = slave_xactor_f_rd_data$EMPTY_N ;
  // value method slave_m_rid
  assign slave_rid = slave_xactor_f_rd_data$D_OUT[70:67] ;
  // value method slave_m_rdata
  assign slave_rdata = slave_xactor_f_rd_data$D_OUT[66:3] ;
  // value method slave_m_rresp
  assign slave_rresp = slave_xactor_f_rd_data$D_OUT[2:1] ;
  // value method slave_m_rlast
  assign slave_rlast = slave_xactor_f_rd_data$D_OUT[0] ;
  // action method slave_m_rready
  assign CAN_FIRE_slave_m_rready = 1'd1 ;
  assign WILL_FIRE_slave_m_rready = 1'd1 ;
  // submodule slave_xactor_f_rd_addr
  FIFO2 #(.width(32'd97), .guarded(32'd1)) slave_xactor_f_rd_addr(.RST(RST_N),
								  .CLK(CLK),
								  .D_IN(slave_xactor_f_rd_addr$D_IN),
								  .ENQ(slave_xactor_f_rd_addr$ENQ),
								  .DEQ(slave_xactor_f_rd_addr$DEQ),
								  .CLR(slave_xactor_f_rd_addr$CLR),
								  .D_OUT(slave_xactor_f_rd_addr$D_OUT),
								  .FULL_N(slave_xactor_f_rd_addr$FULL_N),
								  .EMPTY_N(slave_xactor_f_rd_addr$EMPTY_N));
  // submodule slave_xactor_f_rd_data
  FIFO2 #(.width(32'd71), .guarded(32'd1)) slave_xactor_f_rd_data(.RST(RST_N),
								  .CLK(CLK),
								  .D_IN(slave_xactor_f_rd_data$D_IN),
								  .ENQ(slave_xactor_f_rd_data$ENQ),
								  .DEQ(slave_xactor_f_rd_data$DEQ),
								  .CLR(slave_xactor_f_rd_data$CLR),
								  .D_OUT(slave_xactor_f_rd_data$D_OUT),
								  .FULL_N(slave_xactor_f_rd_data$FULL_N),
								  .EMPTY_N(slave_xactor_f_rd_data$EMPTY_N));
  // submodule slave_xactor_f_wr_addr
  FIFO2 #(.width(32'd97), .guarded(32'd1)) slave_xactor_f_wr_addr(.RST(RST_N),
								  .CLK(CLK),
								  .D_IN(slave_xactor_f_wr_addr$D_IN),
								  .ENQ(slave_xactor_f_wr_addr$ENQ),
								  .DEQ(slave_xactor_f_wr_addr$DEQ),
								  .CLR(slave_xactor_f_wr_addr$CLR),
								  .D_OUT(slave_xactor_f_wr_addr$D_OUT),
								  .FULL_N(slave_xactor_f_wr_addr$FULL_N),
								  .EMPTY_N(slave_xactor_f_wr_addr$EMPTY_N));
  // submodule slave_xactor_f_wr_data
  FIFO2 #(.width(32'd73), .guarded(32'd1)) slave_xactor_f_wr_data(.RST(RST_N),
								  .CLK(CLK),
								  .D_IN(slave_xactor_f_wr_data$D_IN),
								  .ENQ(slave_xactor_f_wr_data$ENQ),
								  .DEQ(slave_xactor_f_wr_data$DEQ),
								  .CLR(slave_xactor_f_wr_data$CLR),
								  .D_OUT(),
								  .FULL_N(slave_xactor_f_wr_data$FULL_N),
								  .EMPTY_N(slave_xactor_f_wr_data$EMPTY_N));
  // submodule slave_xactor_f_wr_resp
  FIFO2 #(.width(32'd6), .guarded(32'd1)) slave_xactor_f_wr_resp(.RST(RST_N),
								 .CLK(CLK),
								 .D_IN(slave_xactor_f_wr_resp$D_IN),
								 .ENQ(slave_xactor_f_wr_resp$ENQ),
								 .DEQ(slave_xactor_f_wr_resp$DEQ),
								 .CLR(slave_xactor_f_wr_resp$CLR),
								 .D_OUT(slave_xactor_f_wr_resp$D_OUT),
								 .FULL_N(slave_xactor_f_wr_resp$FULL_N),
								 .EMPTY_N(slave_xactor_f_wr_resp$EMPTY_N));
  // rule RL_rl_process_rd_req
  assign CAN_FIRE_RL_rl_process_rd_req =
	     slave_xactor_f_rd_addr$EMPTY_N &&
	     slave_xactor_f_rd_data$FULL_N &&
	     rg_module_ready ;
  assign WILL_FIRE_RL_rl_process_rd_req = CAN_FIRE_RL_rl_process_rd_req ;
  // rule RL_rl_process_wr_req
  assign CAN_FIRE_RL_rl_process_wr_req =
	     slave_xactor_f_wr_addr$EMPTY_N &&
	     slave_xactor_f_wr_data$EMPTY_N &&
	     slave_xactor_f_wr_resp$FULL_N &&
	     rg_module_ready ;
  assign WILL_FIRE_RL_rl_process_wr_req = CAN_FIRE_RL_rl_process_wr_req ;
  // register rg_addr_base
  assign rg_addr_base$D_IN = set_addr_map_addr_base ;
  assign rg_addr_base$EN = EN_set_addr_map ;
  // register rg_addr_lim
  assign rg_addr_lim$D_IN = set_addr_map_addr_lim ;
  assign rg_addr_lim$EN = EN_set_addr_map ;
  // register rg_module_ready
  assign rg_module_ready$D_IN = 1'd1 ;
  assign rg_module_ready$EN = EN_set_addr_map ;
  // submodule slave_xactor_f_rd_addr
  assign slave_xactor_f_rd_addr$D_IN =
	     { slave_arid,
	       slave_araddr,
	       slave_arlen,
	       slave_arsize,
	       slave_arburst,
	       slave_arlock,
	       slave_arcache,
	       slave_arprot,
	       slave_arqos,
	       slave_arregion } ;
  assign slave_xactor_f_rd_addr$ENQ =
	     slave_arvalid && slave_xactor_f_rd_addr$FULL_N ;
  assign slave_xactor_f_rd_addr$DEQ = CAN_FIRE_RL_rl_process_rd_req ;
  assign slave_xactor_f_rd_addr$CLR = 1'b0 ;
  // submodule slave_xactor_f_rd_data
  assign slave_xactor_f_rd_data$D_IN =
	     { slave_xactor_f_rd_addr$D_OUT[96:93],
	       rdata__h924,
	       rdr_rresp__h957,
	       1'd1 } ;
  assign slave_xactor_f_rd_data$ENQ = CAN_FIRE_RL_rl_process_rd_req ;
  assign slave_xactor_f_rd_data$DEQ =
	     slave_rready && slave_xactor_f_rd_data$EMPTY_N ;
  assign slave_xactor_f_rd_data$CLR = 1'b0 ;
  // submodule slave_xactor_f_wr_addr
  assign slave_xactor_f_wr_addr$D_IN =
	     { slave_awid,
	       slave_awaddr,
	       slave_awlen,
	       slave_awsize,
	       slave_awburst,
	       slave_awlock,
	       slave_awcache,
	       slave_awprot,
	       slave_awqos,
	       slave_awregion } ;
  assign slave_xactor_f_wr_addr$ENQ =
	     slave_awvalid && slave_xactor_f_wr_addr$FULL_N ;
  assign slave_xactor_f_wr_addr$DEQ = CAN_FIRE_RL_rl_process_wr_req ;
  assign slave_xactor_f_wr_addr$CLR = 1'b0 ;
  // submodule slave_xactor_f_wr_data
  assign slave_xactor_f_wr_data$D_IN =
	     { slave_wdata, slave_wstrb, slave_wlast } ;
  assign slave_xactor_f_wr_data$ENQ =
	     slave_wvalid && slave_xactor_f_wr_data$FULL_N ;
  assign slave_xactor_f_wr_data$DEQ = CAN_FIRE_RL_rl_process_wr_req ;
  assign slave_xactor_f_wr_data$CLR = 1'b0 ;
  // submodule slave_xactor_f_wr_resp
  assign slave_xactor_f_wr_resp$D_IN =
	     { slave_xactor_f_wr_addr$D_OUT[96:93],
	       NOT_slave_xactor_f_wr_addr_first__208_BITS_31__ETC___d1218 ?
		 2'b10 :
		 2'b0 } ;
  assign slave_xactor_f_wr_resp$ENQ = CAN_FIRE_RL_rl_process_wr_req ;
  assign slave_xactor_f_wr_resp$DEQ =
	     slave_bready && slave_xactor_f_wr_resp$EMPTY_N ;
  assign slave_xactor_f_wr_resp$CLR = 1'b0 ;
  // remaining internal signals
  assign NOT_slave_xactor_f_rd_addr_first_BITS_31_TO_29_ETC___d18 =
	     slave_xactor_f_rd_addr$D_OUT[31:29] != 3'b0 ||
	     rg_addr_base > slave_xactor_f_rd_addr$D_OUT[92:29] ||
	     slave_xactor_f_rd_addr$D_OUT[92:29] >= rg_addr_lim ;
  assign NOT_slave_xactor_f_wr_addr_first__208_BITS_31__ETC___d1218 =
	     slave_xactor_f_wr_addr$D_OUT[31:29] != 3'b0 ||
	     rg_addr_base > slave_xactor_f_wr_addr$D_OUT[92:29] ||
	     slave_xactor_f_wr_addr$D_OUT[92:29] >= rg_addr_lim ;
  assign byte_addr__h705 =
	     slave_xactor_f_rd_addr$D_OUT[92:29] - rg_addr_base ;
  assign rdata__h924 =
	     NOT_slave_xactor_f_rd_addr_first_BITS_31_TO_29_ETC___d18 ?
	       64'd0 :
	       data64__h987 ;
  assign rdr_rresp__h957 =
	     NOT_slave_xactor_f_rd_addr_first_BITS_31_TO_29_ETC___d18 ?
	       2'b10 :
	       2'b0 ;
  always@(byte_addr__h705)
  begin
    case (byte_addr__h705)
      64'd16,
      64'd24,
      64'd56,
      64'd72,
      64'd80,
      64'd88,
      64'd200,
      64'd232,
      64'd312,
      64'd424,
      64'd448,
      64'd600,
      64'd728,
      64'd1136,
      64'd1144,
      64'd1152,
      64'd1160,
      64'd1168,
      64'd1176,
      64'd1184,
      64'd1192,
      64'd1200,
      64'd1208,
      64'd1216,
      64'd1224,
      64'd1232,
      64'd1240,
      64'd1248,
      64'd1256,
      64'd1264,
      64'd1272,
      64'd1280,
      64'd1288,
      64'd1296,
      64'd1304,
      64'd1312,
      64'd1320,
      64'd1328,
      64'd1336,
      64'd1344,
      64'd1352,
      64'd1360,
      64'd1368,
      64'd1376,
      64'd1384,
      64'd1392,
      64'd1400,
      64'd1408,
      64'd1416,
      64'd1424,
      64'd1432,
      64'd1440,
      64'd1448,
      64'd1456,
      64'd1464,
      64'd1472,
      64'd1480,
      64'd1488,
      64'd1496,
      64'd1504,
      64'd1512,
      64'd1520,
      64'd1528,
      64'd1536,
      64'd1544,
      64'd1552,
      64'd1560,
      64'd1568,
      64'd1576,
      64'd1584,
      64'd1592,
      64'd1600,
      64'd1608,
      64'd1616,
      64'd1624,
      64'd1632,
      64'd1640,
      64'd1648,
      64'd1656,
      64'd1664,
      64'd1672,
      64'd1680,
      64'd1688,
      64'd1696,
      64'd1704,
      64'd1712,
      64'd1720,
      64'd1728,
      64'd1736,
      64'd1744,
      64'd1752,
      64'd1760,
      64'd1768,
      64'd1776,
      64'd1784,
      64'd1792,
      64'd1800,
      64'd1808,
      64'd1816,
      64'd1824,
      64'd1832,
      64'd1840,
      64'd1848,
      64'd1856,
      64'd1864,
      64'd1872,
      64'd1880,
      64'd1888,
      64'd1896,
      64'd1904,
      64'd1912,
      64'd1920,
      64'd1928,
      64'd1936,
      64'd1944,
      64'd1952,
      64'd1960,
      64'd1968,
      64'd1976,
      64'd1984,
      64'd1992,
      64'd2000,
      64'd2008,
      64'd2016,
      64'd2024,
      64'd2032,
      64'd2040,
      64'd2048,
      64'd2056,
      64'd2064,
      64'd2072,
      64'd2080,
      64'd2088,
      64'd2096,
      64'd2104,
      64'd2112,
      64'd2120,
      64'd2128,
      64'd2136,
      64'd2144,
      64'd2152,
      64'd2160,
      64'd2168,
      64'd2176,
      64'd2184,
      64'd2192,
      64'd2200,
      64'd2208,
      64'd2216,
      64'd2224,
      64'd2232,
      64'd2240,
      64'd2248,
      64'd2256,
      64'd2264,
      64'd2272,
      64'd2280,
      64'd2288,
      64'd2296,
      64'd2304,
      64'd2312,
      64'd2320,
      64'd2328,
      64'd2336,
      64'd2344,
      64'd2352,
      64'd2360,
      64'd2368,
      64'd2376,
      64'd2384,
      64'd2392,
      64'd2400,
      64'd2408,
      64'd2416,
      64'd2424,
      64'd2432,
      64'd2440,
      64'd2448,
      64'd2456,
      64'd2464,
      64'd2472,
      64'd2480,
      64'd2488,
      64'd2496,
      64'd2504,
      64'd2512,
      64'd2520,
      64'd2528,
      64'd2536,
      64'd2544,
      64'd2552,
      64'd2560,
      64'd2568,
      64'd2576,
      64'd2584,
      64'd2592,
      64'd2600,
      64'd2608,
      64'd2616,
      64'd2624,
      64'd2632,
      64'd2640,
      64'd2648,
      64'd2656,
      64'd2664,
      64'd2672,
      64'd2680,
      64'd2688,
      64'd2696,
      64'd2704,
      64'd2712,
      64'd2720,
      64'd2728,
      64'd2736,
      64'd2744,
      64'd2752,
      64'd2760,
      64'd2768,
      64'd2776,
      64'd2784,
      64'd2792,
      64'd2800,
      64'd2808,
      64'd2816,
      64'd2824,
      64'd2832,
      64'd2840,
      64'd2848,
      64'd2856,
      64'd2864,
      64'd2872,
      64'd2880,
      64'd2888,
      64'd2896,
      64'd2904,
      64'd2912,
      64'd2920,
      64'd2928,
      64'd2936,
      64'd2944,
      64'd2952,
      64'd2960,
      64'd2968,
      64'd2976,
      64'd2984,
      64'd2992,
      64'd3000,
      64'd3008,
      64'd3016,
      64'd3024,
      64'd3032,
      64'd3040,
      64'd3048,
      64'd3056,
      64'd3064,
      64'd3072,
      64'd3080,
      64'd3088,
      64'd3096,
      64'd3104,
      64'd3112,
      64'd3120,
      64'd3128,
      64'd3136,
      64'd3144,
      64'd3152,
      64'd3160,
      64'd3168,
      64'd3176,
      64'd3184,
      64'd3192,
      64'd3200,
      64'd3208,
      64'd3216,
      64'd3224,
      64'd3232,
      64'd3240,
      64'd3248,
      64'd3256,
      64'd3264,
      64'd3272,
      64'd3280,
      64'd3288,
      64'd3296,
      64'd3304,
      64'd3312,
      64'd3320,
      64'd3328,
      64'd3336,
      64'd3344,
      64'd3352,
      64'd3360,
      64'd3368,
      64'd3376,
      64'd3384,
      64'd3392,
      64'd3400,
      64'd3408,
      64'd3416,
      64'd3424,
      64'd3432,
      64'd3440,
      64'd3448,
      64'd3456,
      64'd3464,
      64'd3472,
      64'd3480,
      64'd3488,
      64'd3496,
      64'd3504,
      64'd3512,
      64'd3520,
      64'd3528,
      64'd3536,
      64'd3544,
      64'd3552,
      64'd3560,
      64'd3568,
      64'd3576,
      64'd3584,
      64'd3592,
      64'd3600,
      64'd3608,
      64'd3616,
      64'd3624,
      64'd3632,
      64'd3640,
      64'd3648,
      64'd3656,
      64'd3664,
      64'd3672,
      64'd3680,
      64'd3688,
      64'd3696,
      64'd3704,
      64'd3712,
      64'd3720,
      64'd3728,
      64'd3736,
      64'd3744,
      64'd3752,
      64'd3760,
      64'd3768,
      64'd3776,
      64'd3784,
      64'd3792,
      64'd3800,
      64'd3808,
      64'd3816,
      64'd3824,
      64'd3832,
      64'd3840,
      64'd3848,
      64'd3856,
      64'd3864,
      64'd3872,
      64'd3880,
      64'd3888,
      64'd3896,
      64'd3904,
      64'd3912,
      64'd3920,
      64'd3928,
      64'd3936,
      64'd3944,
      64'd3952,
      64'd3960,
      64'd3968,
      64'd3976,
      64'd3984,
      64'd3992,
      64'd4000,
      64'd4008,
      64'd4016,
      64'd4024,
      64'd4032,
      64'd4040,
      64'd4048,
      64'd4056,
      64'd4064,
      64'd4072,
      64'd4080,
      64'd4088:
	  CASE_byte_addr05_16_0x0_24_0x0_32_0x54040000_4_ETC__q1 = 32'h0;
      64'd32:
	  CASE_byte_addr05_16_0x0_24_0x0_32_0x54040000_4_ETC__q1 =
	      32'h54040000;
      64'd40:
	  CASE_byte_addr05_16_0x0_24_0x0_32_0x54040000_4_ETC__q1 =
	      32'h88030000;
      64'd48:
	  CASE_byte_addr05_16_0x0_24_0x0_32_0x54040000_4_ETC__q1 =
	      32'h11000000;
      64'd64:
	  CASE_byte_addr05_16_0x0_24_0x0_32_0x54040000_4_ETC__q1 =
	      32'h50030000;
      64'd96,
      64'd112,
      64'd208,
      64'd224,
      64'd240,
      64'd432,
      64'd488,
      64'd872,
      64'd888:
	  CASE_byte_addr05_16_0x0_24_0x0_32_0x54040000_4_ETC__q1 =
	      32'h04000000;
      64'd104, 64'd120, 64'd504, 64'd792, 64'd920:
	  CASE_byte_addr05_16_0x0_24_0x0_32_0x54040000_4_ETC__q1 =
	      32'h02000000;
      64'd128:
	  CASE_byte_addr05_16_0x0_24_0x0_32_0x54040000_4_ETC__q1 =
	      32'h16000000;
      64'd136:
	  CASE_byte_addr05_16_0x0_24_0x0_32_0x54040000_4_ETC__q1 =
	      32'h62626375;
      64'd144:
	  CASE_byte_addr05_16_0x0_24_0x0_32_0x54040000_4_ETC__q1 =
	      32'h656B6970;
      64'd152:
	  CASE_byte_addr05_16_0x0_24_0x0_32_0x54040000_4_ETC__q1 =
	      32'h65642D65;
      64'd160,
      64'd264,
      64'd280,
      64'd296,
      64'd336,
      64'd360,
      64'd384,
      64'd456,
      64'd552,
      64'd592,
      64'd608,
      64'd624,
      64'd672,
      64'd704,
      64'd760,
      64'd816,
      64'd840,
      64'd880:
	  CASE_byte_addr05_16_0x0_24_0x0_32_0x54040000_4_ETC__q1 =
	      32'h03000000;
      64'd168:
	  CASE_byte_addr05_16_0x0_24_0x0_32_0x54040000_4_ETC__q1 =
	      32'h26000000;
      64'd176, 64'd640:
	  CASE_byte_addr05_16_0x0_24_0x0_32_0x54040000_4_ETC__q1 =
	      32'h732C7261;
      64'd184, 64'd648:
	  CASE_byte_addr05_16_0x0_24_0x0_32_0x54040000_4_ETC__q1 =
	      32'h7261622D;
      64'd192,
      64'd216,
      64'd400,
      64'd440,
      64'd496,
      64'd512,
      64'd584,
      64'd744,
      64'd752,
      64'd912:
	  CASE_byte_addr05_16_0x0_24_0x0_32_0x54040000_4_ETC__q1 =
	      32'h01000000;
      64'd248, 64'd896:
	  CASE_byte_addr05_16_0x0_24_0x0_32_0x54040000_4_ETC__q1 =
	      32'h80969800;
      64'd256:
	  CASE_byte_addr05_16_0x0_24_0x0_32_0x54040000_4_ETC__q1 =
	      32'h40757063;
      64'd272:
	  CASE_byte_addr05_16_0x0_24_0x0_32_0x54040000_4_ETC__q1 =
	      32'h3F000000;
      64'd288, 64'd560, 64'd768, 64'd848:
	  CASE_byte_addr05_16_0x0_24_0x0_32_0x54040000_4_ETC__q1 =
	      32'h4B000000;
      64'd304:
	  CASE_byte_addr05_16_0x0_24_0x0_32_0x54040000_4_ETC__q1 =
	      32'h4F000000;
      64'd320:
	  CASE_byte_addr05_16_0x0_24_0x0_32_0x54040000_4_ETC__q1 =
	      32'h06000000;
      64'd328:
	  CASE_byte_addr05_16_0x0_24_0x0_32_0x54040000_4_ETC__q1 =
	      32'h63736972;
      64'd344:
	  CASE_byte_addr05_16_0x0_24_0x0_32_0x54040000_4_ETC__q1 =
	      32'h56000000;
      64'd352:
	  CASE_byte_addr05_16_0x0_24_0x0_32_0x54040000_4_ETC__q1 =
	      32'h75616D69;
      64'd368:
	  CASE_byte_addr05_16_0x0_24_0x0_32_0x54040000_4_ETC__q1 =
	      32'h60000000;
      64'd376:
	  CASE_byte_addr05_16_0x0_24_0x0_32_0x54040000_4_ETC__q1 =
	      32'h76732C76;
      64'd392:
	  CASE_byte_addr05_16_0x0_24_0x0_32_0x54040000_4_ETC__q1 =
	      32'h69000000;
      64'd408:
	  CASE_byte_addr05_16_0x0_24_0x0_32_0x54040000_4_ETC__q1 =
	      32'h70757272;
      64'd416:
	  CASE_byte_addr05_16_0x0_24_0x0_32_0x54040000_4_ETC__q1 =
	      32'h6F72746E;
      64'd464, 64'd632, 64'd712, 64'd824:
	  CASE_byte_addr05_16_0x0_24_0x0_32_0x54040000_4_ETC__q1 =
	      32'h1B000000;
      64'd472:
	  CASE_byte_addr05_16_0x0_24_0x0_32_0x54040000_4_ETC__q1 =
	      32'h70632C76;
      64'd480:
	  CASE_byte_addr05_16_0x0_24_0x0_32_0x54040000_4_ETC__q1 =
	      32'h00006374;
      64'd520:
	  CASE_byte_addr05_16_0x0_24_0x0_32_0x54040000_4_ETC__q1 =
	      32'h38407972;
      64'd528:
	  CASE_byte_addr05_16_0x0_24_0x0_32_0x54040000_4_ETC__q1 =
	      32'h00303030;
      64'd536:
	  CASE_byte_addr05_16_0x0_24_0x0_32_0x54040000_4_ETC__q1 =
	      32'h07000000;
      64'd544:
	  CASE_byte_addr05_16_0x0_24_0x0_32_0x54040000_4_ETC__q1 =
	      32'h6F6D656D;
      64'd568:
	  CASE_byte_addr05_16_0x0_24_0x0_32_0x54040000_4_ETC__q1 =
	      32'h00000080;
      64'd576:
	  CASE_byte_addr05_16_0x0_24_0x0_32_0x54040000_4_ETC__q1 =
	      32'h00000010;
      64'd616:
	  CASE_byte_addr05_16_0x0_24_0x0_32_0x54040000_4_ETC__q1 =
	      32'h0F000000;
      64'd656:
	  CASE_byte_addr05_16_0x0_24_0x0_32_0x54040000_4_ETC__q1 =
	      32'h69730063;
      64'd664:
	  CASE_byte_addr05_16_0x0_24_0x0_32_0x54040000_4_ETC__q1 =
	      32'h7375622D;
      64'd680:
	  CASE_byte_addr05_16_0x0_24_0x0_32_0x54040000_4_ETC__q1 =
	      32'hA7000000;
      64'd688:
	  CASE_byte_addr05_16_0x0_24_0x0_32_0x54040000_4_ETC__q1 =
	      32'h6E696C63;
      64'd696, 64'd808:
	  CASE_byte_addr05_16_0x0_24_0x0_32_0x54040000_4_ETC__q1 =
	      32'h30303030;
      64'd720:
	  CASE_byte_addr05_16_0x0_24_0x0_32_0x54040000_4_ETC__q1 =
	      32'h6C632C76;
      64'd736:
	  CASE_byte_addr05_16_0x0_24_0x0_32_0x54040000_4_ETC__q1 =
	      32'h10000000;
      64'd776:
	  CASE_byte_addr05_16_0x0_24_0x0_32_0x54040000_4_ETC__q1 =
	      32'h00000002;
      64'd784:
	  CASE_byte_addr05_16_0x0_24_0x0_32_0x54040000_4_ETC__q1 =
	      32'h00000C00;
      64'd800:
	  CASE_byte_addr05_16_0x0_24_0x0_32_0x54040000_4_ETC__q1 =
	      32'h74726175;
      64'd832:
	  CASE_byte_addr05_16_0x0_24_0x0_32_0x54040000_4_ETC__q1 =
	      32'h61303535;
      64'd856:
	  CASE_byte_addr05_16_0x0_24_0x0_32_0x54040000_4_ETC__q1 =
	      32'h000000C0;
      64'd864:
	  CASE_byte_addr05_16_0x0_24_0x0_32_0x54040000_4_ETC__q1 =
	      32'h40000000;
      64'd904:
	  CASE_byte_addr05_16_0x0_24_0x0_32_0x54040000_4_ETC__q1 =
	      32'h08000000;
      64'd928:
	  CASE_byte_addr05_16_0x0_24_0x0_32_0x54040000_4_ETC__q1 =
	      32'h09000000;
      64'd936:
	  CASE_byte_addr05_16_0x0_24_0x0_32_0x54040000_4_ETC__q1 =
	      32'h73736572;
      64'd944:
	  CASE_byte_addr05_16_0x0_24_0x0_32_0x54040000_4_ETC__q1 =
	      32'h2300736C;
      64'd952:
	  CASE_byte_addr05_16_0x0_24_0x0_32_0x54040000_4_ETC__q1 =
	      32'h6C65632D;
      64'd960:
	  CASE_byte_addr05_16_0x0_24_0x0_32_0x54040000_4_ETC__q1 =
	      32'h61706D6F;
      64'd968:
	  CASE_byte_addr05_16_0x0_24_0x0_32_0x54040000_4_ETC__q1 =
	      32'h6F6D0065;
      64'd976:
	  CASE_byte_addr05_16_0x0_24_0x0_32_0x54040000_4_ETC__q1 =
	      32'h656D6974;
      64'd984:
	  CASE_byte_addr05_16_0x0_24_0x0_32_0x54040000_4_ETC__q1 =
	      32'h6572662D;
      64'd992:
	  CASE_byte_addr05_16_0x0_24_0x0_32_0x54040000_4_ETC__q1 =
	      32'h64007963;
      64'd1000:
	  CASE_byte_addr05_16_0x0_24_0x0_32_0x54040000_4_ETC__q1 =
	      32'h79745F65;
      64'd1008:
	  CASE_byte_addr05_16_0x0_24_0x0_32_0x54040000_4_ETC__q1 =
	      32'h73006765;
      64'd1016:
	  CASE_byte_addr05_16_0x0_24_0x0_32_0x54040000_4_ETC__q1 =
	      32'h69720073;
      64'd1024:
	  CASE_byte_addr05_16_0x0_24_0x0_32_0x54040000_4_ETC__q1 =
	      32'h00617369;
      64'd1032:
	  CASE_byte_addr05_16_0x0_24_0x0_32_0x54040000_4_ETC__q1 =
	      32'h65707974;
      64'd1040:
	  CASE_byte_addr05_16_0x0_24_0x0_32_0x54040000_4_ETC__q1 =
	      32'h662D6B63;
      64'd1048:
	  CASE_byte_addr05_16_0x0_24_0x0_32_0x54040000_4_ETC__q1 =
	      32'h79636E65;
      64'd1056, 64'd1072:
	  CASE_byte_addr05_16_0x0_24_0x0_32_0x54040000_4_ETC__q1 =
	      32'h72726574;
      64'd1064:
	  CASE_byte_addr05_16_0x0_24_0x0_32_0x54040000_4_ETC__q1 =
	      32'h6C6C6563;
      64'd1080:
	  CASE_byte_addr05_16_0x0_24_0x0_32_0x54040000_4_ETC__q1 =
	      32'h746E6F63;
      64'd1088:
	  CASE_byte_addr05_16_0x0_24_0x0_32_0x54040000_4_ETC__q1 =
	      32'h70007265;
      64'd1096:
	  CASE_byte_addr05_16_0x0_24_0x0_32_0x54040000_4_ETC__q1 =
	      32'h7200656C;
      64'd1104:
	  CASE_byte_addr05_16_0x0_24_0x0_32_0x54040000_4_ETC__q1 =
	      32'h6E690073;
      64'd1112:
	  CASE_byte_addr05_16_0x0_24_0x0_32_0x54040000_4_ETC__q1 =
	      32'h73747075;
      64'd1120:
	  CASE_byte_addr05_16_0x0_24_0x0_32_0x54040000_4_ETC__q1 =
	      32'h65646E65;
      64'd1128:
	  CASE_byte_addr05_16_0x0_24_0x0_32_0x54040000_4_ETC__q1 =
	      32'h68732D67;
      default: CASE_byte_addr05_16_0x0_24_0x0_32_0x54040000_4_ETC__q1 =
		   32'hAAAAAAAA;
    endcase
  end
  always@(byte_addr__h705)
  begin
    case (byte_addr__h705)
      64'd16:
	  CASE_byte_addr05_16_0x28067_24_0x80000000_32_0_ETC__q2 =
	      32'h00028067;
      64'd24:
	  CASE_byte_addr05_16_0x28067_24_0x80000000_32_0_ETC__q2 =
	      32'h80000000;
      64'd32:
	  CASE_byte_addr05_16_0x28067_24_0x80000000_32_0_ETC__q2 =
	      32'hEDFE0DD0;
      64'd40:
	  CASE_byte_addr05_16_0x28067_24_0x80000000_32_0_ETC__q2 =
	      32'h38000000;
      64'd48:
	  CASE_byte_addr05_16_0x28067_24_0x80000000_32_0_ETC__q2 =
	      32'h28000000;
      64'd56, 64'd560, 64'd768, 64'd848:
	  CASE_byte_addr05_16_0x28067_24_0x80000000_32_0_ETC__q2 =
	      32'h10000000;
      64'd64:
	  CASE_byte_addr05_16_0x28067_24_0x80000000_32_0_ETC__q2 =
	      32'hCC000000;
      64'd72,
      64'd80,
      64'd104,
      64'd216,
      64'd296,
      64'd568,
      64'd576,
      64'd672,
      64'd680,
      64'd776,
      64'd784,
      64'd840,
      64'd856,
      64'd864,
      64'd1144,
      64'd1152,
      64'd1160,
      64'd1168,
      64'd1176,
      64'd1184,
      64'd1192,
      64'd1200,
      64'd1208,
      64'd1216,
      64'd1224,
      64'd1232,
      64'd1240,
      64'd1248,
      64'd1256,
      64'd1264,
      64'd1272,
      64'd1280,
      64'd1288,
      64'd1296,
      64'd1304,
      64'd1312,
      64'd1320,
      64'd1328,
      64'd1336,
      64'd1344,
      64'd1352,
      64'd1360,
      64'd1368,
      64'd1376,
      64'd1384,
      64'd1392,
      64'd1400,
      64'd1408,
      64'd1416,
      64'd1424,
      64'd1432,
      64'd1440,
      64'd1448,
      64'd1456,
      64'd1464,
      64'd1472,
      64'd1480,
      64'd1488,
      64'd1496,
      64'd1504,
      64'd1512,
      64'd1520,
      64'd1528,
      64'd1536,
      64'd1544,
      64'd1552,
      64'd1560,
      64'd1568,
      64'd1576,
      64'd1584,
      64'd1592,
      64'd1600,
      64'd1608,
      64'd1616,
      64'd1624,
      64'd1632,
      64'd1640,
      64'd1648,
      64'd1656,
      64'd1664,
      64'd1672,
      64'd1680,
      64'd1688,
      64'd1696,
      64'd1704,
      64'd1712,
      64'd1720,
      64'd1728,
      64'd1736,
      64'd1744,
      64'd1752,
      64'd1760,
      64'd1768,
      64'd1776,
      64'd1784,
      64'd1792,
      64'd1800,
      64'd1808,
      64'd1816,
      64'd1824,
      64'd1832,
      64'd1840,
      64'd1848,
      64'd1856,
      64'd1864,
      64'd1872,
      64'd1880,
      64'd1888,
      64'd1896,
      64'd1904,
      64'd1912,
      64'd1920,
      64'd1928,
      64'd1936,
      64'd1944,
      64'd1952,
      64'd1960,
      64'd1968,
      64'd1976,
      64'd1984,
      64'd1992,
      64'd2000,
      64'd2008,
      64'd2016,
      64'd2024,
      64'd2032,
      64'd2040,
      64'd2048,
      64'd2056,
      64'd2064,
      64'd2072,
      64'd2080,
      64'd2088,
      64'd2096,
      64'd2104,
      64'd2112,
      64'd2120,
      64'd2128,
      64'd2136,
      64'd2144,
      64'd2152,
      64'd2160,
      64'd2168,
      64'd2176,
      64'd2184,
      64'd2192,
      64'd2200,
      64'd2208,
      64'd2216,
      64'd2224,
      64'd2232,
      64'd2240,
      64'd2248,
      64'd2256,
      64'd2264,
      64'd2272,
      64'd2280,
      64'd2288,
      64'd2296,
      64'd2304,
      64'd2312,
      64'd2320,
      64'd2328,
      64'd2336,
      64'd2344,
      64'd2352,
      64'd2360,
      64'd2368,
      64'd2376,
      64'd2384,
      64'd2392,
      64'd2400,
      64'd2408,
      64'd2416,
      64'd2424,
      64'd2432,
      64'd2440,
      64'd2448,
      64'd2456,
      64'd2464,
      64'd2472,
      64'd2480,
      64'd2488,
      64'd2496,
      64'd2504,
      64'd2512,
      64'd2520,
      64'd2528,
      64'd2536,
      64'd2544,
      64'd2552,
      64'd2560,
      64'd2568,
      64'd2576,
      64'd2584,
      64'd2592,
      64'd2600,
      64'd2608,
      64'd2616,
      64'd2624,
      64'd2632,
      64'd2640,
      64'd2648,
      64'd2656,
      64'd2664,
      64'd2672,
      64'd2680,
      64'd2688,
      64'd2696,
      64'd2704,
      64'd2712,
      64'd2720,
      64'd2728,
      64'd2736,
      64'd2744,
      64'd2752,
      64'd2760,
      64'd2768,
      64'd2776,
      64'd2784,
      64'd2792,
      64'd2800,
      64'd2808,
      64'd2816,
      64'd2824,
      64'd2832,
      64'd2840,
      64'd2848,
      64'd2856,
      64'd2864,
      64'd2872,
      64'd2880,
      64'd2888,
      64'd2896,
      64'd2904,
      64'd2912,
      64'd2920,
      64'd2928,
      64'd2936,
      64'd2944,
      64'd2952,
      64'd2960,
      64'd2968,
      64'd2976,
      64'd2984,
      64'd2992,
      64'd3000,
      64'd3008,
      64'd3016,
      64'd3024,
      64'd3032,
      64'd3040,
      64'd3048,
      64'd3056,
      64'd3064,
      64'd3072,
      64'd3080,
      64'd3088,
      64'd3096,
      64'd3104,
      64'd3112,
      64'd3120,
      64'd3128,
      64'd3136,
      64'd3144,
      64'd3152,
      64'd3160,
      64'd3168,
      64'd3176,
      64'd3184,
      64'd3192,
      64'd3200,
      64'd3208,
      64'd3216,
      64'd3224,
      64'd3232,
      64'd3240,
      64'd3248,
      64'd3256,
      64'd3264,
      64'd3272,
      64'd3280,
      64'd3288,
      64'd3296,
      64'd3304,
      64'd3312,
      64'd3320,
      64'd3328,
      64'd3336,
      64'd3344,
      64'd3352,
      64'd3360,
      64'd3368,
      64'd3376,
      64'd3384,
      64'd3392,
      64'd3400,
      64'd3408,
      64'd3416,
      64'd3424,
      64'd3432,
      64'd3440,
      64'd3448,
      64'd3456,
      64'd3464,
      64'd3472,
      64'd3480,
      64'd3488,
      64'd3496,
      64'd3504,
      64'd3512,
      64'd3520,
      64'd3528,
      64'd3536,
      64'd3544,
      64'd3552,
      64'd3560,
      64'd3568,
      64'd3576,
      64'd3584,
      64'd3592,
      64'd3600,
      64'd3608,
      64'd3616,
      64'd3624,
      64'd3632,
      64'd3640,
      64'd3648,
      64'd3656,
      64'd3664,
      64'd3672,
      64'd3680,
      64'd3688,
      64'd3696,
      64'd3704,
      64'd3712,
      64'd3720,
      64'd3728,
      64'd3736,
      64'd3744,
      64'd3752,
      64'd3760,
      64'd3768,
      64'd3776,
      64'd3784,
      64'd3792,
      64'd3800,
      64'd3808,
      64'd3816,
      64'd3824,
      64'd3832,
      64'd3840,
      64'd3848,
      64'd3856,
      64'd3864,
      64'd3872,
      64'd3880,
      64'd3888,
      64'd3896,
      64'd3904,
      64'd3912,
      64'd3920,
      64'd3928,
      64'd3936,
      64'd3944,
      64'd3952,
      64'd3960,
      64'd3968,
      64'd3976,
      64'd3984,
      64'd3992,
      64'd4000,
      64'd4008,
      64'd4016,
      64'd4024,
      64'd4032,
      64'd4040,
      64'd4048,
      64'd4056,
      64'd4064,
      64'd4072,
      64'd4080,
      64'd4088:
	  CASE_byte_addr05_16_0x28067_24_0x80000000_32_0_ETC__q2 = 32'h0;
      64'd88, 64'd256, 64'd688, 64'd800:
	  CASE_byte_addr05_16_0x28067_24_0x80000000_32_0_ETC__q2 =
	      32'h01000000;
      64'd96,
      64'd112,
      64'd128,
      64'd208,
      64'd224,
      64'd240,
      64'd320,
      64'd432,
      64'd448,
      64'd488,
      64'd536,
      64'd736,
      64'd752,
      64'd872,
      64'd888,
      64'd904:
	  CASE_byte_addr05_16_0x28067_24_0x80000000_32_0_ETC__q2 =
	      32'h03000000;
      64'd120, 64'd232, 64'd464:
	  CASE_byte_addr05_16_0x28067_24_0x80000000_32_0_ETC__q2 =
	      32'h0F000000;
      64'd136, 64'd328:
	  CASE_byte_addr05_16_0x28067_24_0x80000000_32_0_ETC__q2 =
	      32'h1B000000;
      64'd144:
	  CASE_byte_addr05_16_0x28067_24_0x80000000_32_0_ETC__q2 =
	      32'h732C7261;
      64'd152:
	  CASE_byte_addr05_16_0x28067_24_0x80000000_32_0_ETC__q2 =
	      32'h7261622D;
      64'd160, 64'd336:
	  CASE_byte_addr05_16_0x28067_24_0x80000000_32_0_ETC__q2 =
	      32'h00000076;
      64'd168:
	  CASE_byte_addr05_16_0x28067_24_0x80000000_32_0_ETC__q2 =
	      32'h12000000;
      64'd176, 64'd640:
	  CASE_byte_addr05_16_0x28067_24_0x80000000_32_0_ETC__q2 =
	      32'h62626375;
      64'd184, 64'd648:
	  CASE_byte_addr05_16_0x28067_24_0x80000000_32_0_ETC__q2 =
	      32'h656B6970;
      64'd192:
	  CASE_byte_addr05_16_0x28067_24_0x80000000_32_0_ETC__q2 =
	      32'h00000065;
      64'd200:
	  CASE_byte_addr05_16_0x28067_24_0x80000000_32_0_ETC__q2 =
	      32'h73757063;
      64'd248:
	  CASE_byte_addr05_16_0x28067_24_0x80000000_32_0_ETC__q2 =
	      32'h2C000000;
      64'd264, 64'd704, 64'd816:
	  CASE_byte_addr05_16_0x28067_24_0x80000000_32_0_ETC__q2 =
	      32'h00000030;
      64'd272, 64'd288, 64'd392, 64'd600, 64'd616:
	  CASE_byte_addr05_16_0x28067_24_0x80000000_32_0_ETC__q2 =
	      32'h04000000;
      64'd280:
	  CASE_byte_addr05_16_0x28067_24_0x80000000_32_0_ETC__q2 =
	      32'h00757063;
      64'd304:
	  CASE_byte_addr05_16_0x28067_24_0x80000000_32_0_ETC__q2 =
	      32'h05000000;
      64'd312:
	  CASE_byte_addr05_16_0x28067_24_0x80000000_32_0_ETC__q2 =
	      32'h79616B6F;
      64'd344:
	  CASE_byte_addr05_16_0x28067_24_0x80000000_32_0_ETC__q2 =
	      32'h0A000000;
      64'd352:
	  CASE_byte_addr05_16_0x28067_24_0x80000000_32_0_ETC__q2 =
	      32'h32337672;
      64'd360:
	  CASE_byte_addr05_16_0x28067_24_0x80000000_32_0_ETC__q2 =
	      32'h00000073;
      64'd368, 64'd920:
	  CASE_byte_addr05_16_0x28067_24_0x80000000_32_0_ETC__q2 =
	      32'h0B000000;
      64'd376, 64'd472, 64'd720:
	  CASE_byte_addr05_16_0x28067_24_0x80000000_32_0_ETC__q2 =
	      32'h63736972;
      64'd384:
	  CASE_byte_addr05_16_0x28067_24_0x80000000_32_0_ETC__q2 =
	      32'h00003233;
      64'd400:
	  CASE_byte_addr05_16_0x28067_24_0x80000000_32_0_ETC__q2 =
	      32'h80969800;
      64'd408:
	  CASE_byte_addr05_16_0x28067_24_0x80000000_32_0_ETC__q2 =
	      32'h65746E69;
      64'd416:
	  CASE_byte_addr05_16_0x28067_24_0x80000000_32_0_ETC__q2 =
	      32'h6F632D74;
      64'd424:
	  CASE_byte_addr05_16_0x28067_24_0x80000000_32_0_ETC__q2 =
	      32'h72656C6C;
      64'd440:
	  CASE_byte_addr05_16_0x28067_24_0x80000000_32_0_ETC__q2 =
	      32'h79000000;
      64'd456:
	  CASE_byte_addr05_16_0x28067_24_0x80000000_32_0_ETC__q2 =
	      32'h8A000000;
      64'd480:
	  CASE_byte_addr05_16_0x28067_24_0x80000000_32_0_ETC__q2 =
	      32'h6E692D75;
      64'd496:
	  CASE_byte_addr05_16_0x28067_24_0x80000000_32_0_ETC__q2 =
	      32'h9F000000;
      64'd504, 64'd512, 64'd584, 64'd608, 64'd624, 64'd792, 64'd928:
	  CASE_byte_addr05_16_0x28067_24_0x80000000_32_0_ETC__q2 =
	      32'h02000000;
      64'd520:
	  CASE_byte_addr05_16_0x28067_24_0x80000000_32_0_ETC__q2 =
	      32'h6F6D656D;
      64'd528:
	  CASE_byte_addr05_16_0x28067_24_0x80000000_32_0_ETC__q2 =
	      32'h30303030;
      64'd544:
	  CASE_byte_addr05_16_0x28067_24_0x80000000_32_0_ETC__q2 =
	      32'h3F000000;
      64'd552:
	  CASE_byte_addr05_16_0x28067_24_0x80000000_32_0_ETC__q2 =
	      32'h00007972;
      64'd592:
	  CASE_byte_addr05_16_0x28067_24_0x80000000_32_0_ETC__q2 =
	      32'h00636F73;
      64'd632:
	  CASE_byte_addr05_16_0x28067_24_0x80000000_32_0_ETC__q2 =
	      32'h21000000;
      64'd656:
	  CASE_byte_addr05_16_0x28067_24_0x80000000_32_0_ETC__q2 =
	      32'h6F732D65;
      64'd664:
	  CASE_byte_addr05_16_0x28067_24_0x80000000_32_0_ETC__q2 =
	      32'h656C706D;
      64'd696:
	  CASE_byte_addr05_16_0x28067_24_0x80000000_32_0_ETC__q2 =
	      32'h30324074;
      64'd712:
	  CASE_byte_addr05_16_0x28067_24_0x80000000_32_0_ETC__q2 =
	      32'h0D000000;
      64'd728:
	  CASE_byte_addr05_16_0x28067_24_0x80000000_32_0_ETC__q2 =
	      32'h30746E69;
      64'd744, 64'd912:
	  CASE_byte_addr05_16_0x28067_24_0x80000000_32_0_ETC__q2 =
	      32'hAE000000;
      64'd760:
	  CASE_byte_addr05_16_0x28067_24_0x80000000_32_0_ETC__q2 =
	      32'h07000000;
      64'd808:
	  CASE_byte_addr05_16_0x28067_24_0x80000000_32_0_ETC__q2 =
	      32'h30306340;
      64'd824:
	  CASE_byte_addr05_16_0x28067_24_0x80000000_32_0_ETC__q2 =
	      32'h09000000;
      64'd832:
	  CASE_byte_addr05_16_0x28067_24_0x80000000_32_0_ETC__q2 =
	      32'h3631736E;
      64'd880:
	  CASE_byte_addr05_16_0x28067_24_0x80000000_32_0_ETC__q2 =
	      32'hC2000000;
      64'd896:
	  CASE_byte_addr05_16_0x28067_24_0x80000000_32_0_ETC__q2 =
	      32'h69000000;
      64'd936:
	  CASE_byte_addr05_16_0x28067_24_0x80000000_32_0_ETC__q2 =
	      32'h64646123;
      64'd944:
	  CASE_byte_addr05_16_0x28067_24_0x80000000_32_0_ETC__q2 =
	      32'h6C65632D;
      64'd952:
	  CASE_byte_addr05_16_0x28067_24_0x80000000_32_0_ETC__q2 =
	      32'h657A6973;
      64'd960:
	  CASE_byte_addr05_16_0x28067_24_0x80000000_32_0_ETC__q2 =
	      32'h6300736C;
      64'd968:
	  CASE_byte_addr05_16_0x28067_24_0x80000000_32_0_ETC__q2 =
	      32'h6C626974;
      64'd976:
	  CASE_byte_addr05_16_0x28067_24_0x80000000_32_0_ETC__q2 =
	      32'h006C6564;
      64'd984:
	  CASE_byte_addr05_16_0x28067_24_0x80000000_32_0_ETC__q2 =
	      32'h65736162;
      64'd992:
	  CASE_byte_addr05_16_0x28067_24_0x80000000_32_0_ETC__q2 =
	      32'h6E657571;
      64'd1000:
	  CASE_byte_addr05_16_0x28067_24_0x80000000_32_0_ETC__q2 =
	      32'h63697665;
      64'd1008:
	  CASE_byte_addr05_16_0x28067_24_0x80000000_32_0_ETC__q2 =
	      32'h72006570;
      64'd1016:
	  CASE_byte_addr05_16_0x28067_24_0x80000000_32_0_ETC__q2 =
	      32'h75746174;
      64'd1024:
	  CASE_byte_addr05_16_0x28067_24_0x80000000_32_0_ETC__q2 =
	      32'h2C766373;
      64'd1032:
	  CASE_byte_addr05_16_0x28067_24_0x80000000_32_0_ETC__q2 =
	      32'h2D756D6D;
      64'd1040:
	  CASE_byte_addr05_16_0x28067_24_0x80000000_32_0_ETC__q2 =
	      32'h6F6C6300;
      64'd1048:
	  CASE_byte_addr05_16_0x28067_24_0x80000000_32_0_ETC__q2 =
	      32'h75716572;
      64'd1056:
	  CASE_byte_addr05_16_0x28067_24_0x80000000_32_0_ETC__q2 =
	      32'h6E692300;
      64'd1064, 64'd1080:
	  CASE_byte_addr05_16_0x28067_24_0x80000000_32_0_ETC__q2 =
	      32'h2D747075;
      64'd1072:
	  CASE_byte_addr05_16_0x28067_24_0x80000000_32_0_ETC__q2 =
	      32'h6E690073;
      64'd1088:
	  CASE_byte_addr05_16_0x28067_24_0x80000000_32_0_ETC__q2 =
	      32'h6C6C6F72;
      64'd1096:
	  CASE_byte_addr05_16_0x28067_24_0x80000000_32_0_ETC__q2 =
	      32'h646E6168;
      64'd1104:
	  CASE_byte_addr05_16_0x28067_24_0x80000000_32_0_ETC__q2 =
	      32'h65676E61;
      64'd1112:
	  CASE_byte_addr05_16_0x28067_24_0x80000000_32_0_ETC__q2 =
	      32'h72726574;
      64'd1120:
	  CASE_byte_addr05_16_0x28067_24_0x80000000_32_0_ETC__q2 =
	      32'h7478652D;
      64'd1128:
	  CASE_byte_addr05_16_0x28067_24_0x80000000_32_0_ETC__q2 =
	      32'h65720064;
      64'd1136:
	  CASE_byte_addr05_16_0x28067_24_0x80000000_32_0_ETC__q2 =
	      32'h00746669;
      default: CASE_byte_addr05_16_0x28067_24_0x80000000_32_0_ETC__q2 =
		   32'hAAAAAAAA;
    endcase
  end
  always@(byte_addr__h705 or
	  CASE_byte_addr05_16_0x0_24_0x0_32_0x54040000_4_ETC__q1 or
	  CASE_byte_addr05_16_0x28067_24_0x80000000_32_0_ETC__q2)
  begin
    case (byte_addr__h705)
      64'd0: data64__h987 = 64'h0202859300000297;
      64'd8: data64__h987 = 64'h0182A283F1402573;
      default: data64__h987 =
		   { CASE_byte_addr05_16_0x0_24_0x0_32_0x54040000_4_ETC__q1,
		     CASE_byte_addr05_16_0x28067_24_0x80000000_32_0_ETC__q2 };
    endcase
  end
  // handling of inlined registers
  always@(posedge CLK)
  begin
    if (RST_N == `BSV_RESET_VALUE)
      begin
        rg_module_ready <= `BSV_ASSIGNMENT_DELAY 1'd0;
      end
    else
      begin
        if (rg_module_ready$EN)
	  rg_module_ready <= `BSV_ASSIGNMENT_DELAY rg_module_ready$D_IN;
      end
    if (rg_addr_base$EN)
      rg_addr_base <= `BSV_ASSIGNMENT_DELAY rg_addr_base$D_IN;
    if (rg_addr_lim$EN) rg_addr_lim <= `BSV_ASSIGNMENT_DELAY rg_addr_lim$D_IN;
  end
  // synopsys translate_off
  `ifdef BSV_NO_INITIAL_BLOCKS
  `else // not BSV_NO_INITIAL_BLOCKS
  initial
  begin
    rg_addr_base = 64'hAAAAAAAAAAAAAAAA;
    rg_addr_lim = 64'hAAAAAAAAAAAAAAAA;
    rg_module_ready = 1'h0;
  end
  `endif // BSV_NO_INITIAL_BLOCKS
  // synopsys translate_on
  // handling of system tasks
  // synopsys translate_off
  always@(negedge CLK)
  begin
    #0;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_rd_req &&
	  NOT_slave_xactor_f_rd_addr_first_BITS_31_TO_29_ETC___d18)
	begin
	  v__h808 = $stime;
	  #0;
	end
    v__h802 = v__h808 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_rd_req &&
	  NOT_slave_xactor_f_rd_addr_first_BITS_31_TO_29_ETC___d18)
	$display("%0d: ERROR: Boot_ROM.rl_process_rd_req: unrecognized addr",
		 v__h802);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_rd_req &&
	  NOT_slave_xactor_f_rd_addr_first_BITS_31_TO_29_ETC___d18)
	$write("    ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_rd_req &&
	  NOT_slave_xactor_f_rd_addr_first_BITS_31_TO_29_ETC___d18)
	$write("AXI4_Rd_Addr { ", "arid: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_rd_req &&
	  NOT_slave_xactor_f_rd_addr_first_BITS_31_TO_29_ETC___d18)
	$write("'h%h", slave_xactor_f_rd_addr$D_OUT[96:93]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_rd_req &&
	  NOT_slave_xactor_f_rd_addr_first_BITS_31_TO_29_ETC___d18)
	$write(", ", "araddr: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_rd_req &&
	  NOT_slave_xactor_f_rd_addr_first_BITS_31_TO_29_ETC___d18)
	$write("'h%h", slave_xactor_f_rd_addr$D_OUT[92:29]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_rd_req &&
	  NOT_slave_xactor_f_rd_addr_first_BITS_31_TO_29_ETC___d18)
	$write(", ", "arlen: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_rd_req &&
	  NOT_slave_xactor_f_rd_addr_first_BITS_31_TO_29_ETC___d18)
	$write("'h%h", slave_xactor_f_rd_addr$D_OUT[28:21]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_rd_req &&
	  NOT_slave_xactor_f_rd_addr_first_BITS_31_TO_29_ETC___d18)
	$write(", ", "arsize: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_rd_req &&
	  NOT_slave_xactor_f_rd_addr_first_BITS_31_TO_29_ETC___d18)
	$write("'h%h", slave_xactor_f_rd_addr$D_OUT[20:18]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_rd_req &&
	  NOT_slave_xactor_f_rd_addr_first_BITS_31_TO_29_ETC___d18)
	$write(", ", "arburst: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_rd_req &&
	  NOT_slave_xactor_f_rd_addr_first_BITS_31_TO_29_ETC___d18)
	$write("'h%h", slave_xactor_f_rd_addr$D_OUT[17:16]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_rd_req &&
	  NOT_slave_xactor_f_rd_addr_first_BITS_31_TO_29_ETC___d18)
	$write(", ", "arlock: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_rd_req &&
	  NOT_slave_xactor_f_rd_addr_first_BITS_31_TO_29_ETC___d18)
	$write("'h%h", slave_xactor_f_rd_addr$D_OUT[15]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_rd_req &&
	  NOT_slave_xactor_f_rd_addr_first_BITS_31_TO_29_ETC___d18)
	$write(", ", "arcache: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_rd_req &&
	  NOT_slave_xactor_f_rd_addr_first_BITS_31_TO_29_ETC___d18)
	$write("'h%h", slave_xactor_f_rd_addr$D_OUT[14:11]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_rd_req &&
	  NOT_slave_xactor_f_rd_addr_first_BITS_31_TO_29_ETC___d18)
	$write(", ", "arprot: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_rd_req &&
	  NOT_slave_xactor_f_rd_addr_first_BITS_31_TO_29_ETC___d18)
	$write("'h%h", slave_xactor_f_rd_addr$D_OUT[10:8]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_rd_req &&
	  NOT_slave_xactor_f_rd_addr_first_BITS_31_TO_29_ETC___d18)
	$write(", ", "arqos: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_rd_req &&
	  NOT_slave_xactor_f_rd_addr_first_BITS_31_TO_29_ETC___d18)
	$write("'h%h", slave_xactor_f_rd_addr$D_OUT[7:4]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_rd_req &&
	  NOT_slave_xactor_f_rd_addr_first_BITS_31_TO_29_ETC___d18)
	$write(", ", "arregion: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_rd_req &&
	  NOT_slave_xactor_f_rd_addr_first_BITS_31_TO_29_ETC___d18)
	$write("'h%h", slave_xactor_f_rd_addr$D_OUT[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_rd_req &&
	  NOT_slave_xactor_f_rd_addr_first_BITS_31_TO_29_ETC___d18)
	$write(", ", "aruser: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_rd_req &&
	  NOT_slave_xactor_f_rd_addr_first_BITS_31_TO_29_ETC___d18)
	$write("'h%h", 1'd0, " }");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_rd_req &&
	  NOT_slave_xactor_f_rd_addr_first_BITS_31_TO_29_ETC___d18)
	$write("\n");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_wr_req &&
	  NOT_slave_xactor_f_wr_addr_first__208_BITS_31__ETC___d1218)
	begin
	  v__h8925 = $stime;
	  #0;
	end
    v__h8919 = v__h8925 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_wr_req &&
	  NOT_slave_xactor_f_wr_addr_first__208_BITS_31__ETC___d1218)
	$display("%0d: ERROR: Boot_ROM.rl_process_wr_req: unrecognized addr",
		 v__h8919);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_wr_req &&
	  NOT_slave_xactor_f_wr_addr_first__208_BITS_31__ETC___d1218)
	$write("    ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_wr_req &&
	  NOT_slave_xactor_f_wr_addr_first__208_BITS_31__ETC___d1218)
	$write("AXI4_Wr_Addr { ", "awid: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_wr_req &&
	  NOT_slave_xactor_f_wr_addr_first__208_BITS_31__ETC___d1218)
	$write("'h%h", slave_xactor_f_wr_addr$D_OUT[96:93]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_wr_req &&
	  NOT_slave_xactor_f_wr_addr_first__208_BITS_31__ETC___d1218)
	$write(", ", "awaddr: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_wr_req &&
	  NOT_slave_xactor_f_wr_addr_first__208_BITS_31__ETC___d1218)
	$write("'h%h", slave_xactor_f_wr_addr$D_OUT[92:29]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_wr_req &&
	  NOT_slave_xactor_f_wr_addr_first__208_BITS_31__ETC___d1218)
	$write(", ", "awlen: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_wr_req &&
	  NOT_slave_xactor_f_wr_addr_first__208_BITS_31__ETC___d1218)
	$write("'h%h", slave_xactor_f_wr_addr$D_OUT[28:21]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_wr_req &&
	  NOT_slave_xactor_f_wr_addr_first__208_BITS_31__ETC___d1218)
	$write(", ", "awsize: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_wr_req &&
	  NOT_slave_xactor_f_wr_addr_first__208_BITS_31__ETC___d1218)
	$write("'h%h", slave_xactor_f_wr_addr$D_OUT[20:18]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_wr_req &&
	  NOT_slave_xactor_f_wr_addr_first__208_BITS_31__ETC___d1218)
	$write(", ", "awburst: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_wr_req &&
	  NOT_slave_xactor_f_wr_addr_first__208_BITS_31__ETC___d1218)
	$write("'h%h", slave_xactor_f_wr_addr$D_OUT[17:16]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_wr_req &&
	  NOT_slave_xactor_f_wr_addr_first__208_BITS_31__ETC___d1218)
	$write(", ", "awlock: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_wr_req &&
	  NOT_slave_xactor_f_wr_addr_first__208_BITS_31__ETC___d1218)
	$write("'h%h", slave_xactor_f_wr_addr$D_OUT[15]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_wr_req &&
	  NOT_slave_xactor_f_wr_addr_first__208_BITS_31__ETC___d1218)
	$write(", ", "awcache: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_wr_req &&
	  NOT_slave_xactor_f_wr_addr_first__208_BITS_31__ETC___d1218)
	$write("'h%h", slave_xactor_f_wr_addr$D_OUT[14:11]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_wr_req &&
	  NOT_slave_xactor_f_wr_addr_first__208_BITS_31__ETC___d1218)
	$write(", ", "awprot: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_wr_req &&
	  NOT_slave_xactor_f_wr_addr_first__208_BITS_31__ETC___d1218)
	$write("'h%h", slave_xactor_f_wr_addr$D_OUT[10:8]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_wr_req &&
	  NOT_slave_xactor_f_wr_addr_first__208_BITS_31__ETC___d1218)
	$write(", ", "awqos: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_wr_req &&
	  NOT_slave_xactor_f_wr_addr_first__208_BITS_31__ETC___d1218)
	$write("'h%h", slave_xactor_f_wr_addr$D_OUT[7:4]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_wr_req &&
	  NOT_slave_xactor_f_wr_addr_first__208_BITS_31__ETC___d1218)
	$write(", ", "awregion: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_wr_req &&
	  NOT_slave_xactor_f_wr_addr_first__208_BITS_31__ETC___d1218)
	$write("'h%h", slave_xactor_f_wr_addr$D_OUT[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_wr_req &&
	  NOT_slave_xactor_f_wr_addr_first__208_BITS_31__ETC___d1218)
	$write(", ", "awuser: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_wr_req &&
	  NOT_slave_xactor_f_wr_addr_first__208_BITS_31__ETC___d1218)
	$write("'h%h", 1'd0, " }");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_wr_req &&
	  NOT_slave_xactor_f_wr_addr_first__208_BITS_31__ETC___d1218)
	$write("\n");
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_set_addr_map && set_addr_map_addr_base[2:0] != 3'd0)
	begin
	  v__h9218 = $stime;
	  #0;
	end
    v__h9212 = v__h9218 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_set_addr_map && set_addr_map_addr_base[2:0] != 3'd0)
	$display("%0d: WARNING: Boot_ROM.set_addr_map: addr_base 0x%0h is not 4-Byte-aligned",
		 v__h9212,
		 set_addr_map_addr_base);
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_set_addr_map && set_addr_map_addr_lim[2:0] != 3'd0)
	begin
	  v__h9328 = $stime;
	  #0;
	end
    v__h9322 = v__h9328 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_set_addr_map && set_addr_map_addr_lim[2:0] != 3'd0)
	$display("%0d: WARNING: Boot_ROM.set_addr_map: addr_lim 0x%0h is not 4-Byte-aligned",
		 v__h9322,
		 set_addr_map_addr_lim);
  end
  // synopsys translate_on
endmodule