module can be initiate
            init_flag <= 1;
            water_in_end_sign = 1'b0;
            water_out_end_sign = 1'b0;
            water_level = {3{1'b0}};
        end
    end
endmodule