module reset
    .pulse_out(start)
    );
endmodule