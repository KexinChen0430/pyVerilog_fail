module");
`endif
endmodule