module header
	// Internal signals
	// Generated Signal List
	// End of Generated Signal List
	// %COMPILER_OPTS%
	// Generated Signal Assignments
	// Generated Instances and Port Mappings
		// Generated Instance Port Map for inst_1
		inst_1_e	#(
			.FOO(16)
		) inst_1 (
		);
		// End of Generated Instance Port Map for inst_1
		// Generated Instance Port Map for inst_10
		inst_10_e	#(
			.FOO(32)
		) inst_10 (
		);
		// End of Generated Instance Port Map for inst_10
		// Generated Instance Port Map for inst_2
		inst_2_e	#(
			.FOO(16)
		) inst_2 (
		);
		// End of Generated Instance Port Map for inst_2
		// Generated Instance Port Map for inst_3
		inst_3_e	#(
			.FOO(16)
		) inst_3 (
		);
		// End of Generated Instance Port Map for inst_3
		// Generated Instance Port Map for inst_4
		inst_4_e	#(
			.FOO(16)
		) inst_4 (
		);
		// End of Generated Instance Port Map for inst_4
		// Generated Instance Port Map for inst_5
		inst_5_e inst_5 (
		);
		// End of Generated Instance Port Map for inst_5
		// Generated Instance Port Map for inst_6
		inst_6_e inst_6 (
		);
		// End of Generated Instance Port Map for inst_6
		// Generated Instance Port Map for inst_7
		inst_7_e	#(
			.FOO(32)
		) inst_7 (
		);
		// End of Generated Instance Port Map for inst_7
		// Generated Instance Port Map for inst_8
		inst_8_e	#(
			.FOO(32)
		) inst_8 (
		);
		// End of Generated Instance Port Map for inst_8
		// Generated Instance Port Map for inst_9
		inst_9_e	#(
			.FOO(32)
		) inst_9 (
		);
		// End of Generated Instance Port Map for inst_9
		// Generated Instance Port Map for inst_aa
		inst_aa_e	#(
			.NO_DEFAULT("nodefault"),
			.NO_NAME("noname"),
			.WIDTH(15)
		) inst_aa (
		);
		// End of Generated Instance Port Map for inst_aa
		// Generated Instance Port Map for inst_ab
		inst_ab_e	#(
			.WIDTH(31)
		) inst_ab (
		);
		// End of Generated Instance Port Map for inst_ab
		// Generated Instance Port Map for inst_ac
		inst_ac_e inst_ac (
		);
		// End of Generated Instance Port Map for inst_ac
		// Generated Instance Port Map for inst_ad
		inst_ad_e inst_ad (
		);
		// End of Generated Instance Port Map for inst_ad
		// Generated Instance Port Map for inst_ae
		inst_ae_e inst_ae (
		);
		// End of Generated Instance Port Map for inst_ae
		// Generated Instance Port Map for inst_m1
		inst_m_e	#(
			.FOO(15)
		) inst_m1 (
		);
		// End of Generated Instance Port Map for inst_m1
		// Generated Instance Port Map for inst_m10
		inst_m_e	#(
			.FOO(30)
		) inst_m10 (
		);
		// End of Generated Instance Port Map for inst_m10
		// Generated Instance Port Map for inst_m2
		inst_m_e	#(
			.FOO(15)
		) inst_m2 (
		);
		// End of Generated Instance Port Map for inst_m2
		// Generated Instance Port Map for inst_m3
		inst_m_e	#(
			.FOO(15)
		) inst_m3 (
		);
		// End of Generated Instance Port Map for inst_m3
		// Generated Instance Port Map for inst_m4
		inst_m_e	#(
			.FOO(15)
		) inst_m4 (
		);
		// End of Generated Instance Port Map for inst_m4
		// Generated Instance Port Map for inst_m5
		inst_m_e	#(
			.FOO(15)
		) inst_m5 (
		);
		// End of Generated Instance Port Map for inst_m5
		// Generated Instance Port Map for inst_m6
		inst_m_e	#(
			.FOO(30)
		) inst_m6 (
		);
		// End of Generated Instance Port Map for inst_m6
		// Generated Instance Port Map for inst_m7
		inst_m_e	#(
			.FOO(30)
		) inst_m7 (
		);
		// End of Generated Instance Port Map for inst_m7
		// Generated Instance Port Map for inst_m8
		inst_m_e	#(
			.FOO(30)
		) inst_m8 (
		);
		// End of Generated Instance Port Map for inst_m8
		// Generated Instance Port Map for inst_m9
		inst_m_e	#(
			.FOO(30)
		) inst_m9 (
		);
		// End of Generated Instance Port Map for inst_m9
endmodule