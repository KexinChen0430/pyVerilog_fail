module os4cb78 #(
   parameter FADDR    = 3,   parameter D_WIDTH  = 16 )
   (
   input wire                sys_clk ,
   input wire                rst_n ,
   input wire [(8*`NUM_VC)-1:0]    ofc3555,
   input wire [(8*`NUM_VC)-1:0]    mg1aaad,
   input wire [(8*`NUM_VC)-1:0]    jcd5569,
   input wire [(12*`NUM_VC)-1:0]   jraab4b,
   input wire [(12*`NUM_VC)-1:0]   vv55a5f,
   input wire [(12*`NUM_VC)-1:0]   vkad2fe,
   input wire [6:0]                lq697f3,
   input wire [10:0]               kd4bf9b,
   input wire [6:0]                jp5fcdc,
   input wire [10:0]               lqfe6e7,
   input wire [6:0]                thf373b,
   input wire [10:0]               bn9b9df,
   input wire [11:0]               nt8b8a0,
   input wire [`NUM_VC-1:0]        gb65b08,
   input wire [(`NUM_VC*16) -1:0]  pub7014,
   input wire [`NUM_VC-1:0]        uk10db8,
   input wire [`NUM_VC-1:0]        ng86dc0,
   input wire [`NUM_VC-1:0]        cb36e02,
   input wire                      ls35987,
   input wire [2:0]                phy_cfgln_sum,
   input wire [FADDR:0]            ba250d2,
   input wire                      thd20a8 ,
   input wire [15:0]               icd170d ,
   input wire                      bn8b869 ,
   input wire                      me5c34e ,
   input wire                      qgcbe8c,
   input wire                      fn5f460,
   input wire                      ayfa306,
   input wire [1:0]                sj397d1,
   input wire [2:0]                thec436,
   input wire [19:0]               ui621b7,
   input wire [`NUM_VC-1:0]        aaf45c ,
   input wire                      dmfe774,
   input wire [`NUM_VC -1:0]       ls1e282 ,
   input wire                      ym3bfe4,
   input wire                      rib82be,
   input wire                      icc15f2,
   input wire [`NUM_VC-1:0]        jpd27c8,
   input wire [`NUM_VC-1:0]        do93e46,
   input wire [`NUM_VC-1:0]        mt9f233,
   input wire [`NUM_VC-1:0]        mt18edf,
   input wire [`NUM_VC-1:0]        hbc76fc,
   input wire [`NUM_VC-1:0]        ie3b7e7,
   input wire [`NUM_VC-1:0]        sudbf39,
   input wire [`NUM_VC-1:0]        fadf9c9,
   input wire [`NUM_VC-1:0]        hbfce4b,
   input wire [`NUM_VC-1:0]        mre725f,
   input wire [`NUM_VC-1:0]        kf392fc,
   input wire [`NUM_VC-1:0]        gbc97e4,
   input wire [`NUM_VC-1:0]        cz4bf24,
   input wire [`NUM_VC-1:0]        xj5f924,
   input wire [`NUM_VC-1:0]        vvfc927,
   input wire [(8*`NUM_VC)-1:0]    tue493f,
   input wire [(8*`NUM_VC)-1:0]    mg249fa,
   input wire [(8*`NUM_VC)-1:0]    ie24fd0,
   `ifdef ECRC
      input wire                   ecrc_gen_enb ,
      input wire                   ecrc_chk_enb ,
   `endif
   input wire [2:0]                rtcdaa7 ,
   input wire                      zkd03c5 ,
   output wire                     fa79b01 ,
   output wire [15:0]              kf9ae61 ,
   output wire                     vvd730d ,
   output wire                     ukb986e ,
   output wire                     mrcc371 ,
   output wire                     xjcd80b ,
   output wire                     zk63316 ,
   output wire [`NUM_VC-1:0]       zx64b62,
   output wire [(`NUM_VC*9)-1:0]   qi1a518,
   output wire [(`NUM_VC*13)-1:0]  nrd28c0,
   output wire [(`NUM_VC*9)-1:0]   ph94607,
   output wire [(`NUM_VC*13)-1:0]  coa303f,
   output wire [(`NUM_VC*9)-1:0]   ir181f8,
   output wire [(`NUM_VC*13)-1:0]  dmc0fc5,
   output wire [(`NUM_VC*16)-1:0]  fadf3e5 ,
   output wire [`NUM_VC-1:0]       dzf9f2a ,
   output wire [`NUM_VC-1:0]       facf957 ,
   `ifdef ECRC
      output wire [`NUM_VC-1:0]    tu7caba ,
   `endif
   output wire [`NUM_VC-1:0]       cme55d3 ,
   output wire [`NUM_VC-1:0]       ls2ae99 ,
   output wire                     ftl_err_msg ,
   output wire                     nftl_err_msg ,
   output wire                     cor_err_msg ,
   output wire                     inta_n,
   output wire                     intb_n,
   output wire                     intc_n,
   output wire                     intd_n,
   output wire [`NUM_VC -1:0]      mgacc3b,
   output wire                     lf198b2,
   output wire [2:0]               yxcc596,
   output wire [1:0]               os62cb4,
   output wire                     fp165a1,
   output wire [2:0]               xyb2d0e,
   output wire [1:0]               ba96872,
   output wire [`NUM_VC -1:0]      wlb4393,
   output wire [`NUM_VC -1:0]      uxa1c9c,
   output wire [`NUM_VC -1:0]      vke4e4,
   output wire [(24*`NUM_VC)-1:0]  me6705e,
   output wire [(24*`NUM_VC)-1:0]  lf382f0,
   output wire [(24*`NUM_VC)-1:0]  mec1786
   ) ;
wire [D_WIDTH -1:0]         ksa79d ;
wire [D_WIDTH -1:0]         xwd08ab;
wire                        nt8455a ;
wire                        db22ad6 ;
wire                        sw156b7 ;
wire                        eaeab6b ;
wire                        hb55b59 ;
wire                        ngadace ;
wire                        ayfa03b ;
`ifdef CFG_REG
`endif
`ifdef ECRC
`endif
`ifdef CFG_REG
`endif
`ifdef CFG_VCAT
`endif
reg fn6b391 ;
reg ic59c8e ;
wire ykce470  = db22ad6 & ~fn6b391 ;
wire hd8e04e = sw156b7 & ~ic59c8e ;
`ifdef ECRC
`ifdef ECRC
`endif
`else
`endif
`ifdef ECRC
`endif
`ifdef ECRC
`endif
`ifdef AER
`endif
`ifdef AER
`endif
reg [(8 * `NUM_VC) - 1 : 0] hq83f1a;
reg [(8 * `NUM_VC) - 1 : 0] ec1f8d2;
reg [(8 * `NUM_VC) - 1 : 0] zxfc691;
reg [(12 * `NUM_VC) - 1 : 0] xje348e;
reg [(12 * `NUM_VC) - 1 : 0] sw1a476;
reg [(12 * `NUM_VC) - 1 : 0] dzd23b0;
reg [6 : 0] jr91d86;
reg [10 : 0] fp8ec36;
reg [6 : 0] tu761b6;
reg [10 : 0] bnb0db3;
reg [6 : 0] ls86d9f;
reg [10 : 0] mt36cfa;
reg [11 : 0] ir95972;
reg [`NUM_VC - 1 : 0] ym5efc;
reg [(`NUM_VC * 16) - 1 : 0] ks1f831;
reg [`NUM_VC - 1 : 0] ayce8fc;
reg [`NUM_VC - 1 : 0] hb747e0;
reg [`NUM_VC - 1 : 0] coa3f06;
reg bl64b01;
reg [2 : 0] ir9afed;
reg [FADDR : 0] gdbe052;
reg rtfc2b3;
reg [15 : 0] wl23286;
reg nt19434;
reg rgca1a7;
reg kf2c072;
reg cz60395;
reg ls1cad;
reg [1 : 0] pue56b;
reg [2 : 0] ld7b3a3;
reg [19 : 0] shd9d1f;
reg [`NUM_VC - 1 : 0] mgb992f;
reg wy8dd9b;
reg [`NUM_VC - 1 : 0] vv7e6c2;
reg an9f508;
reg ofc3f97;
reg ie1fcbc;
reg [`NUM_VC - 1 : 0] mefa844;
reg [`NUM_VC - 1 : 0] uid4220;
reg [`NUM_VC - 1 : 0] sja1101;
reg [`NUM_VC - 1 : 0] ri1b63;
reg [`NUM_VC - 1 : 0] mtdb1b;
reg [`NUM_VC - 1 : 0] ay6d8dd;
reg [`NUM_VC - 1 : 0] vi6c6e8;
reg [`NUM_VC - 1 : 0] lq63743;
reg [`NUM_VC - 1 : 0] ba1ba1a;
reg [`NUM_VC - 1 : 0] bldd0d3;
reg [`NUM_VC - 1 : 0] ale869f;
reg [`NUM_VC - 1 : 0] yk434fd;
reg [`NUM_VC - 1 : 0] ou1a7e9;
reg [`NUM_VC - 1 : 0] wjd3f48;
reg [`NUM_VC - 1 : 0] ir9fa45;
reg [(8 * `NUM_VC) - 1 : 0] enfd22d;
reg [(8 * `NUM_VC) - 1 : 0] lde916c;
reg [(8 * `NUM_VC) - 1 : 0] jc48b67;
reg [2 : 0] gd26aed;
reg wje877b;
reg [D_WIDTH - 1 : 0] fp197a6;
reg eacbd37;
reg mr5e9b8;
reg jcf4dc5;
reg jr2d704;
reg vv6b827;
reg kq5c13f;
reg ho6cefe;
reg fc4fc8;
reg vx27e43;
reg hq3f21f;
reg nrf90fb;
reg [2047:0] necf6c2;
wire [68:0] ld7b613;
`ifdef CFG_REG
`endif
`ifdef ECRC
`endif
`ifdef CFG_REG
`endif
`ifdef CFG_VCAT
`endif
`ifdef ECRC
`ifdef ECRC
`endif
`else
`endif
`ifdef ECRC
`endif
`ifdef ECRC
`endif
`ifdef AER
`endif
`ifdef AER
`endif
localparam qgdb09f = 69,nrd84f8 = 32'hfdffd30b;
localparam [31:0] thc27c7 = nrd84f8;
localparam mt9f1ff = nrd84f8 & 4'hf;
localparam [11:0] fnc7fe5 = 'h7ff;
wire  [(1 << mt9f1ff)  -1:0] suff972;
reg    [qgdb09f-1:0] cme5c87;
reg [mt9f1ff-1:0] qg721c0 [0:1];
reg [mt9f1ff-1:0] ym8700c;
reg rv38061;
integer jcc030e;
integer vk1872;
`ifdef CFG_REG
`endif
`ifdef ECRC
`endif
`ifdef CFG_REG
`endif
`ifdef CFG_VCAT
`endif
`ifdef ECRC
`ifdef ECRC
`endif
`else
`endif
`ifdef ECRC
`endif
`ifdef ECRC
`endif
`ifdef AER
`endif
`ifdef AER
`endif
gq9284a qge0915   (        .sys_clk              ( sys_clk ),    .rst_n                ( rst_n ),    .czcc9db         ( 3'd0 ),
    .ld4a3ee           ( 1'b0 ),    .uv51f77          ( 1'b0 ),    .oh8fbbc           ( 1'b0 ),
`ifdef CFG_REG
       .gb44cfd      ( 1'b0 ),       .zkeef21       ( 1'b0 ),       .qg7790b     ( 64'd0 ),       .kqce688     ( 1'b0 ),
`endif
`ifdef ECRC
       .cba14f3          ( ecrc_gen_enb ) ,
`endif
    .gb65b08               ( ym5efc ),    .pub7014              ( ks1f831 ),    .uk10db8                ( ayce8fc ),    .ng86dc0               ( hb747e0 ),    .cb36e02              ( coa3f06 ),    .thd20a8             ( rtfc2b3 ),    .ba250d2        ( gdbe052 ),    .ls1e282           ( vv7e6c2),        .en5b0c9     ( zk63316 ),    .cbab5b9       ( cbab5b9 ),
`ifdef CFG_REG
       .enc3267       (  ),
`endif
   .ux28d2           (  ),   .fc14694           (  ),   .twb80a3             (  ),   .zkc051a             (  ),
`ifdef CFG_VCAT
       .uxb10aa      (  ),
`endif
    .zx64b62               ( zx64b62 ),    .goefa4f           ( fa79b01 ),    .xwd08ab          ( xwd08ab ),    .nt8455a            ( nt8455a ),    .db22ad6           ( db22ad6 ),    .sw156b7          ( sw156b7 ),
    .by791cf       (  ),    .nrc8e7a      (  ),    .jc473d7        (  ),    .an39ebb         (  )    );
always @(posedge sys_clk, negedge rst_n) begin   if (!rst_n) begin      fn6b391  <= 1'b0 ;      ic59c8e <= 1'b0 ;   end   else if (vv6b827) begin      fn6b391  <= mr5e9b8 ;      ic59c8e <= jcf4dc5 ;   end
end
`ifdef ECRC
   ri20e84 tj8460b (            .sys_clk        ( sys_clk ) ,      .rst_n          ( rst_n ) ,            .xwd08ab    ( fp197a6 ) ,      .nt8455a      ( eacbd37 ) ,      .db22ad6     ( hq3f21f ) ,      .sw156b7    ( nrf90fb ) ,      .cbab5b9 ( cbab5b9 ) ,
`ifdef ECRC
         .cba14f3    ( ecrc_gen_enb ) ,
`endif
            .kf9ae61    ( kf9ae61 ) ,      .vvd730d      ( vvd730d ) ,      .ukb986e     ( ukb986e ) ,      .mrcc371    ( mrcc371 ) ,      .xjcd80b ( xjcd80b )      ) ;
`else
   assign kf9ae61    = fp197a6 ;   assign vvd730d      = eacbd37 ;   assign ukb986e     = hq3f21f ;   assign mrcc371    = nrf90fb ;   assign xjcd80b = cbab5b9 ;
`endif
ouacceb aa8dc71 (      .sys_clk            ( sys_clk ) ,   .rst_n              ( rst_n ) ,      .icd170d          ( wl23286 ) ,   .bn8b869            ( nt19434 ) ,   .me5c34e           ( rgca1a7 ) ,   .rtcdaa7        ( gd26aed ) ,   .aaf45c              ( mgb992f[0] ) ,
`ifdef ECRC
      .cba14f3        ( ecrc_chk_enb ) ,
`endif
      .ksa79d        ( fadf3e5 ) ,   .kq53ce9          ( dzf9f2a ) ,   .rv9e749         ( facf957 ) ,   .ayfa03b   ( ayfa03b ),
`ifdef ECRC
      .ks9d276 ( tu7caba ) ,
`endif
   .vve93b1    ( cme55d3 ) ,   .kq49d8f    ( ls2ae99 ),   .inta_n             ( inta_n ) ,   .intb_n             ( intb_n ) ,   .intc_n             ( intc_n ) ,   .intd_n             ( intd_n ) ,   .ftl_err_msg        ( ftl_err_msg ) ,   .nftl_err_msg       ( nftl_err_msg ) ,   .cor_err_msg        ( cor_err_msg )
   ) ;
bn1c004 pfc2dd1(      .sys_clk                  (sys_clk),   .rst_n                    (rst_n),   .dmfe774              (wy8dd9b),   .hb7e87f                    (1'b1),   .al4bbdd                     (3'd0),   .uk10db8                    (ayce8fc),   .ng86dc0                   (hb747e0),   .cb36e02                  (coa3f06),   .pub7014                  (ks1f831),   .twb80a3                (1'b0 ),   .zkc051a                (1'b0 ),   .ux28d2              (1'b0 ),   .fc14694              (1'b0 ),   .qgcbe8c            (kf2c072),   .fn5f460            (cz60395),   .ayfa306             (ls1cad),   .sj397d1            (pue56b),   .thec436            (ld7b3a3),   .ui621b7            (shd9d1f),      .aaa34a3          ( ),   .qi1a518                 (qi1a518),   .nrd28c0                 (nrd28c0),   .ph94607                (ph94607),   .coa303f                (coa303f),   .ir181f8               (ir181f8),   .dmc0fc5               (dmc0fc5)   ) ;
al7af2f pf55f78(         .sys_clk                  (sys_clk),   .rst_n                    (rst_n),      .ofc3555               (hq83f1a),   .mg1aaad              (ec1f8d2),   .jcd5569             (zxfc691),   .jraab4b               (xje348e),   .vv55a5f              (sw1a476),   .vkad2fe             (dzd23b0),   .lq697f3           (jr91d86),   .kd4bf9b           (fp8ec36),   .jp5fcdc          (tu761b6),   .lqfe6e7          (bnb0db3),   .thf373b         (ls86d9f),   .bn9b9df         (mt36cfa),   .nt8b8a0             (ir95972),
   .ls1e282               (vv7e6c2),   .yxe2831             (wje877b),   .ym3bfe4               (an9f508),   .rib82be               (ofc3f97),   .icc15f2               (ie1fcbc),   .jpd27c8              (mefa844),   .do93e46             (uid4220),   .mt9f233            (sja1101),   .mt18edf            (ri1b63),   .hbc76fc            (mtdb1b),   .ie3b7e7           (ay6d8dd),   .sudbf39           (vi6c6e8),   .fadf9c9          (lq63743),   .hbfce4b          (ba1ba1a),   .mre725f             (bldd0d3),   .kf392fc             (ale869f),   .gbc97e4            (yk434fd),   .cz4bf24            (ou1a7e9),   .xj5f924           (wjd3f48),   .vvfc927           (ir9fa45),   .fp27e80        (1'b0),   .je3f407        (1'b0),   .ayfa03b         (ho6cefe),
   .tue493f                   (enfd22d),   .mg249fa                  (lde916c),   .ie24fd0                 (jc48b67),
`ifdef AER
       .hod01d9                  ({(`NUM_VC){1'b0}}),   .sj80ecb                  (1'b0),   .ux765d                  (1'b0),   .ie3b2ed                 (1'b0),   .uvd9769                 (1'b0),   .uicbb4d             (9'd0),   .jc5da68              (1'b0),   .iped342              (1'b0),   .lq69a15             (1'b0),   .fa4d0aa             (1'b0),
`endif
      .lf198b2               (lf198b2),   .yxcc596                 (yxcc596),   .os62cb4                 (os62cb4),   .fp165a1               (fp165a1),   .xyb2d0e                 (xyb2d0e),   .ba96872                 (ba96872),   .wlb4393            (wlb4393),   .uxa1c9c           (uxa1c9c),   .vke4e4          (vke4e4),
`ifdef AER
      .kd54529           ( ),
`endif
   .me6705e                     (me6705e),   .lf382f0                    (lf382f0),   .mec1786                   (mec1786)   ) ;
always@* begin hq83f1a<={ofc3555>>1,ld7b613[0]};ec1f8d2<={mg1aaad>>1,ld7b613[1]};zxfc691<={jcd5569>>1,ld7b613[2]};xje348e<={jraab4b>>1,ld7b613[3]};sw1a476<={vv55a5f>>1,ld7b613[4]};dzd23b0<={vkad2fe>>1,ld7b613[5]};jr91d86<={lq697f3>>1,ld7b613[6]};fp8ec36<={kd4bf9b>>1,ld7b613[7]};tu761b6<={jp5fcdc>>1,ld7b613[8]};bnb0db3<={lqfe6e7>>1,ld7b613[9]};ls86d9f<={thf373b>>1,ld7b613[10]};mt36cfa<={bn9b9df>>1,ld7b613[11]};ir95972<={nt8b8a0>>1,ld7b613[12]};ym5efc<={gb65b08>>1,ld7b613[13]};ks1f831<={pub7014>>1,ld7b613[14]};ayce8fc<={uk10db8>>1,ld7b613[15]};hb747e0<={ng86dc0>>1,ld7b613[16]};coa3f06<={cb36e02>>1,ld7b613[17]};bl64b01<=ld7b613[18];ir9afed<={phy_cfgln_sum>>1,ld7b613[19]};gdbe052<={ba250d2>>1,ld7b613[20]};rtfc2b3<=ld7b613[21];wl23286<={icd170d>>1,ld7b613[22]};nt19434<=ld7b613[23];rgca1a7<=ld7b613[24];kf2c072<=ld7b613[25];cz60395<=ld7b613[26];ls1cad<=ld7b613[27];pue56b<={sj397d1>>1,ld7b613[28]};ld7b3a3<={thec436>>1,ld7b613[29]};shd9d1f<={ui621b7>>1,ld7b613[30]};mgb992f<={aaf45c>>1,ld7b613[31]};wy8dd9b<=ld7b613[32];vv7e6c2<={ls1e282>>1,ld7b613[33]};an9f508<=ld7b613[34];ofc3f97<=ld7b613[35];ie1fcbc<=ld7b613[36];mefa844<={jpd27c8>>1,ld7b613[37]};uid4220<={do93e46>>1,ld7b613[38]};sja1101<={mt9f233>>1,ld7b613[39]};ri1b63<={mt18edf>>1,ld7b613[40]};mtdb1b<={hbc76fc>>1,ld7b613[41]};ay6d8dd<={ie3b7e7>>1,ld7b613[42]};vi6c6e8<={sudbf39>>1,ld7b613[43]};lq63743<={fadf9c9>>1,ld7b613[44]};ba1ba1a<={hbfce4b>>1,ld7b613[45]};bldd0d3<={mre725f>>1,ld7b613[46]};ale869f<={kf392fc>>1,ld7b613[47]};yk434fd<={gbc97e4>>1,ld7b613[48]};ou1a7e9<={cz4bf24>>1,ld7b613[49]};wjd3f48<={xj5f924>>1,ld7b613[50]};ir9fa45<={vvfc927>>1,ld7b613[51]};enfd22d<={tue493f>>1,ld7b613[52]};lde916c<={mg249fa>>1,ld7b613[53]};jc48b67<={ie24fd0>>1,ld7b613[54]};gd26aed<={rtcdaa7>>1,ld7b613[55]};wje877b<=ld7b613[56];fp197a6<={xwd08ab>>1,ld7b613[57]};eacbd37<=ld7b613[58];mr5e9b8<=ld7b613[59];jcf4dc5<=ld7b613[60];jr2d704<=ld7b613[61];vv6b827<=ld7b613[62];kq5c13f<=ld7b613[63];ho6cefe<=ld7b613[64];fc4fc8<=ld7b613[65];vx27e43<=ld7b613[66];hq3f21f<=ld7b613[67];nrf90fb<=ld7b613[68];end
always@* begin necf6c2[2047]<=mg1aaad[0];necf6c2[2046]<=jcd5569[0];necf6c2[2044]<=jraab4b[0];necf6c2[2040]<=vv55a5f[0];necf6c2[2032]<=vkad2fe[0];necf6c2[2016]<=lq697f3[0];necf6c2[1985]<=kd4bf9b[0];necf6c2[1947]<=fn6b391;necf6c2[1922]<=jp5fcdc[0];necf6c2[1893]<=rtcdaa7[0];necf6c2[1847]<=ic59c8e;necf6c2[1796]<=lqfe6e7[0];necf6c2[1739]<=zkd03c5;necf6c2[1732]<=thec436[0];necf6c2[1646]<=ykce470;necf6c2[1630]<=db22ad6;necf6c2[1600]<=fadf9c9[0];necf6c2[1572]<=dmfe774;necf6c2[1544]<=thf373b[0];necf6c2[1510]<=ngadace;necf6c2[1457]<=ayfa306;necf6c2[1431]<=xwd08ab[0];necf6c2[1417]<=ui621b7[0];necf6c2[1302]<=thd20a8;necf6c2[1244]<=hd8e04e;necf6c2[1212]<=sw156b7;necf6c2[1164]<=jpd27c8[0];necf6c2[1153]<=hbfce4b[0];necf6c2[1124]<=mt18edf[0];necf6c2[1115]<=bn8b869;necf6c2[1105]<=cb36e02[0];necf6c2[1096]<=ls1e282[0];necf6c2[1041]<=bn9b9df[0];necf6c2[1038]<=gbc97e4[0];necf6c2[1023]<=ofc3555[0];necf6c2[973]<=ayfa03b;necf6c2[946]<=ie24fd0[0];necf6c2[866]<=sj397d1[0];necf6c2[815]<=nt8455a;necf6c2[800]<=sudbf39[0];necf6c2[786]<=aaf45c[0];necf6c2[755]<=hb55b59;necf6c2[728]<=fn5f460;necf6c2[651]<=ba250d2[0];necf6c2[582]<=icc15f2;necf6c2[562]<=mt9f233[0];necf6c2[557]<=icd170d[0];necf6c2[552]<=ng86dc0[0];necf6c2[519]<=kf392fc[0];necf6c2[473]<=mg249fa[0];necf6c2[400]<=ie3b7e7[0];necf6c2[377]<=eaeab6b;necf6c2[364]<=qgcbe8c;necf6c2[325]<=phy_cfgln_sum[0];necf6c2[291]<=rib82be;necf6c2[281]<=do93e46[0];necf6c2[276]<=uk10db8[0];necf6c2[259]<=mre725f[0];necf6c2[236]<=tue493f[0];necf6c2[200]<=hbc76fc[0];necf6c2[182]<=me5c34e;necf6c2[162]<=ls35987;necf6c2[145]<=ym3bfe4;necf6c2[138]<=pub7014[0];necf6c2[118]<=vvfc927[0];necf6c2[69]<=gb65b08[0];necf6c2[59]<=xj5f924[0];necf6c2[34]<=nt8b8a0[0];necf6c2[29]<=cz4bf24[0];end         assign suff972 = necf6c2,ld7b613 = cme5c87;   initial begin   jcc030e = $fopen(".fred");   $fdisplay( jcc030e, "%3h\n%3h", (thc27c7 >> 4) & fnc7fe5, (thc27c7 >> (mt9f1ff+4)) & fnc7fe5 );   $fclose(jcc030e);   $readmemh(".fred", qg721c0);   end   always @ (suff972) begin   ym8700c = qg721c0[1];       for (vk1872=0; vk1872<qgdb09f; vk1872=vk1872+1) begin           cme5c87[vk1872] = suff972[ym8700c];       rv38061  = ^(ym8700c & qg721c0[0]);       ym8700c =  {ym8700c, rv38061};       end   end
endmodule