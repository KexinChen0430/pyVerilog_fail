module biosrom (Address, OutClock, OutClockEn, Reset, Q)/* synthesis NGD_DRC_MASK=1 */;
    input wire [9:0] Address;
    input wire OutClock;
    input wire OutClockEn;
    input wire Reset;
    output wire [15:0] Q;
    wire scuba_vhi;
    wire scuba_vlo;
    VHI scuba_vhi_inst (.Z(scuba_vhi));
    VLO scuba_vlo_inst (.Z(scuba_vlo));
    defparam biosrom_0_0_0.INITVAL_3F = "0x0E500000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam biosrom_0_0_0.INITVAL_3E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam biosrom_0_0_0.INITVAL_3D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam biosrom_0_0_0.INITVAL_3C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam biosrom_0_0_0.INITVAL_3B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam biosrom_0_0_0.INITVAL_3A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam biosrom_0_0_0.INITVAL_39 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam biosrom_0_0_0.INITVAL_38 = "0x00000000000000000000000000000000000000000007406978045000202002020020200202002020" ;
    defparam biosrom_0_0_0.INITVAL_37 = "0x02020020200202002020020200202002020020200202002020020200202002020020200202002020" ;
    defparam biosrom_0_0_0.INITVAL_36 = "0x020200006C06F6306F7406F720500005D32031300303A0746C07561066650442002039039390392E" ;
    defparam biosrom_0_0_0.INITVAL_35 = "0x02E31030300305B02020020200202002020020200202002020020200202000070061470206506D61" ;
    defparam biosrom_0_0_0.INITVAL_34 = "0x07246020720657406E490005D038310353103A3702030038320313A03620034320303103A3502032" ;
    defparam biosrom_0_0_0.INITVAL_33 = "0x0313503A34020360353203A33020380323103A32020340363A0315B0202002020020200202002020" ;
    defparam biosrom_0_0_0.INITVAL_32 = "0x0202002020020200202002020020200006507A69053200746506B6306150000000047B0047800473" ;
    defparam biosrom_0_0_0.INITVAL_31 = "0x0070B004620045200441006D50041100401003D500698003C7003B7003AD006480006C0656306E61" ;
    defparam biosrom_0_0_0.INITVAL_30 = "0x0433A0637304520020730656706E6106863020640726106373069640206406E6102074069780453A" ;
    defparam biosrom_0_0_0.INITVAL_2F = "0x04E20073650676E061680632006576061730206406E6102074069780453A059000294E02F590283F" ;
    defparam biosrom_0_0_0.INITVAL_2E = "0x02073072650746506D61072610502006576061530006D06574049200656706E610684303A7206574" ;
    defparam biosrom_0_0_0.INITVAL_2D = "0x06E45020200736D0657404920074630656C0655303A1901800079740696C0697405520061720616B" ;
    defparam biosrom_0_0_0.INITVAL_2C = "0x075670614D0000A00D290756E0656D02065068740207007520074720617407320073690205A02D54" ;
    defparam biosrom_0_0_0.INITVAL_2B = "0x04C410280A00D0A00D2E0657506E690746E06F630206F074200796506B200796E061200737306572" ;
    defparam biosrom_0_0_0.INITVAL_2A = "0x0500A00D0A00D7006A2E0646102E65064690772E063660734007D6E06168063630616D02C610726F" ;
    defparam biosrom_0_0_0.INITVAL_29 = "0x0737B0202C034310303202D3203130032200746806769072790706F0430A00D300302E0302006E6F" ;
    defparam biosrom_0_0_0.INITVAL_28 = "0x069730726505620079740696C0697405520061720616B075670614D0C358059100CD20000B9001B4" ;
    defparam biosrom_0_0_0.INITVAL_27 = "0x051500C35805B59010CD0071100E8B001B4010CD002B40FF3205153050C30EAEB0465805B100CDFF" ;
    defparam biosrom_0_0_0.INITVAL_26 = "0x0320E0B453050900900F074C00840408A2E0C35A0585B059100CD090B4FF03251053500581F00450" ;
    defparam biosrom_0_0_0.INITVAL_25 = "0x016890D88E0C03301E50052C3058590EFEB0C2FE04600008E80909000A740C0840048A02E00001B9" ;
    defparam biosrom_0_0_0.INITVAL_24 = "0x051500C35805B5905A1F010CD000000B9070B706000B804A040843608A0404A1608AD808EC00331E" ;
    defparam biosrom_0_0_0.INITVAL_23 = "0x05251053500C3C30FFB40C346000040C6C305FF80E246047050880408A00010B90071A0BF570C3FD" ;
    defparam biosrom_0_0_0.INITVAL_22 = "0x0E6E80001000714006C70900000713006C60C35F0F8E204647004880058A000100B90701ABF057C3" ;
    defparam biosrom_0_0_0.INITVAL_21 = "0x00718016890DEEB0D00A004E20C12002C90090040721003C0702C900900C0720A03C3002C900901B" ;
    defparam biosrom_0_0_0.INITVAL_20 = "0x074C0084460048A0D2330909002A740003C080C30FE370E80000407014060C79000107013060C6C3" ;
    defparam biosrom_0_0_0.INITVAL_1F = "0x046040880700490090040723A03C30004040E2C1004E80C0C608AC305A00004C6000050E800008E8" ;
    defparam biosrom_0_0_0.INITVAL_1E = "0x0000B0E80000EE8007180168B052C3007170A23002C9009007074C00840408AC30FE810E80000107" ;
    defparam biosrom_0_0_0.INITVAL_1D = "0x014060C79000207013060C6C3004890E43203004007170A0C30CF030071400E8B0F4EB046C20FEFE" ;
    defparam biosrom_0_0_0.INITVAL_1C = "0x0B28400F0003C800FEB90E9F708BD002AC702BC608BFE0C4E905E5A0012D0E800001B9020B00011C" ;
    defparam biosrom_0_0_0.INITVAL_1B = "0x0E852056CA0FE4E05EF6075C0084460FF440880408A560FEE50840F0F73B090160EB5E0F6750C084" ;
    defparam biosrom_0_0_0.INITVAL_1A = "0x04604088010448A056FE0FA8400F0003C800FF010E94E0CAFE0FF070840F0F73B0FF0D0E9460C2FE" ;
    defparam biosrom_0_0_0.INITVAL_19 = "0x0FF130840F0003C080C30FF1B0E9C20FE01084E8000010B9240889009004075E408446004880248A" ;
    defparam biosrom_0_0_0.INITVAL_18 = "0x0FF330830F0F13B0008C0E8FF03CE905EFF040E90C2FE0465A05E01093E805652004880F6770F13B" ;
    defparam biosrom_0_0_0.INITVAL_17 = "0x04E24088FF0648A059900901C073F103BF3075E4084460248A09090029730F13B056000C1E809090" ;
    defparam biosrom_0_0_0.INITVAL_16 = "0x0377401F5808004017060F6D808EC00335001E820774603C860724103CDF0248C07490002070133E" ;
    defparam biosrom_0_0_0.INITVAL_15 = "0x08090090140763903C9A0723003C900901E07490000070133E080A80722003C000AB8400F530003D" ;
    defparam biosrom_0_0_0.INITVAL_14 = "0x0B3740520003D000FF8400F4F0003D000A50840F04D0003D000B98400F4B0003D000B20840F04800" ;
    defparam biosrom_0_0_0.INITVAL_13 = "0x03D010108400F470003D000C00840F0500003D000C78400F1C0FC80000CE0840F001FC0800100584" ;
    defparam biosrom_0_0_0.INITVAL_12 = "0x00F0803C160CD000B4100CD020B4FF0325E05A0204DE8052560FE8B0029F0E8F0000FF0F0EA0D7EB" ;
    defparam biosrom_0_0_0.INITVAL_11 = "0x0F8E204746005880048A000670BF0701ABE000100B900065A3007180A100064A2007170A0C3010CD" ;
    defparam biosrom_0_0_0.INITVAL_10 = "0x0007F025100CD0F0B4E90754E03C90090100745903CDF024FE0ED8400F010FC80016CD000B40029C" ;
    defparam biosrom_0_0_0.INITVAL_0F = "0x0E8050E7BE018000BA070B3020A7E8005D00BE14005BA070B30FF270E990006550FF2E0072A0BEFF" ;
    defparam biosrom_0_0_0.INITVAL_0E = "0x0328500F1C0FC8009090014740FFFC0805F0032C0E890004550FF2E057150B20702ABE09002055FF" ;
    defparam biosrom_0_0_0.INITVAL_0D = "0x02E0702ABE002E20E8070B3070163600202001BA090900358B02EF800306026BF0E4F6008B400716" ;
    defparam biosrom_0_0_0.INITVAL_0C = "0x0A0FF074E90900000716006C60FF7D0820F090040071603E8000716006FE08BEB0900300716006C6" ;
    defparam biosrom_0_0_0.INITVAL_0B = "0x093790071600EFE0E5EB090900297401CFC0809009019074500FC800909001274048FC080160CD00" ;
    defparam biosrom_0_0_0.INITVAL_0A = "0x0B4B90EBC60FE90008C708303047E80072A0BE150B290002550FF2E0072A0BE03070E80CA2A00015" ;
    defparam biosrom_0_0_0.INITVAL_09 = "0x0B9200B003061E8007B304603067E8070B3090900047500716006380022C0C68A007B30909003D74" ;
    defparam biosrom_0_0_0.INITVAL_08 = "0x0F685090900358B001B2006260BF020B60308BE8005AD0BE18000BA003940E80509CBE0D233007B3" ;
    defparam biosrom_0_0_0.INITVAL_07 = "0x0037C0E804001E80F8E204746005880048A0071A0BF00067BE000100B907018A3000650A107017A2" ;
    defparam biosrom_0_0_0.INITVAL_06 = "0x000640A0070110E089100CDFF032030B4CB004880FBE20460402AF6033C003249009E10C1CB00077" ;
    defparam biosrom_0_0_0.INITVAL_05 = "0x006C60000200E88009E90C1010FFC108100078B90CB00024E8090900057502C0003D160CD000B490" ;
    defparam biosrom_0_0_0.INITVAL_04 = "0x00FEB0E47504AEA0E2900900A075160CD010B4FA075100A8610E4FA074100A8610E482035B900008" ;
    defparam biosrom_0_0_0.INITVAL_03 = "0x0BA04053E80050A0BE1F00E20020200202002020020500445502F340565004900012010000000000" ;
    defparam biosrom_0_0_0.INITVAL_02 = "0x00000000040000000000000000000008000037760524904350000290204D04F52020540412F04350" ;
    defparam biosrom_0_0_0.INITVAL_01 = "0x0207206F6602028020650676106D490206D061720676F072500206506C7006D610532004D4F05220" ;
    defparam biosrom_0_0_0.INITVAL_00 = "0x06E6F069740704F0004C04D4F0526E06F690747004F20064720616F0424904350090720EB040AA55" ;
    defparam biosrom_0_0_0.CSDECODE_B = "0b111" ;
    defparam biosrom_0_0_0.CSDECODE_A = "0b000" ;
    defparam biosrom_0_0_0.WRITEMODE_B = "NORMAL" ;
    defparam biosrom_0_0_0.WRITEMODE_A = "NORMAL" ;
    defparam biosrom_0_0_0.GSR = "DISABLED" ;
    defparam biosrom_0_0_0.REGMODE_B = "NOREG" ;
    defparam biosrom_0_0_0.REGMODE_A = "NOREG" ;
    defparam biosrom_0_0_0.DATA_WIDTH_B = 18 ;
    defparam biosrom_0_0_0.DATA_WIDTH_A = 18 ;
    DP16KC biosrom_0_0_0 (.DIA0(scuba_vlo), .DIA1(scuba_vlo), .DIA2(scuba_vlo),
        .DIA3(scuba_vlo), .DIA4(scuba_vlo), .DIA5(scuba_vlo), .DIA6(scuba_vlo),
        .DIA7(scuba_vlo), .DIA8(scuba_vlo), .DIA9(scuba_vlo), .DIA10(scuba_vlo),
        .DIA11(scuba_vlo), .DIA12(scuba_vlo), .DIA13(scuba_vlo), .DIA14(scuba_vlo),
        .DIA15(scuba_vlo), .DIA16(scuba_vlo), .DIA17(scuba_vlo), .ADA0(scuba_vlo),
        .ADA1(scuba_vlo), .ADA2(scuba_vlo), .ADA3(scuba_vlo), .ADA4(Address[0]),
        .ADA5(Address[1]), .ADA6(Address[2]), .ADA7(Address[3]), .ADA8(Address[4]),
        .ADA9(Address[5]), .ADA10(Address[6]), .ADA11(Address[7]), .ADA12(Address[8]),
        .ADA13(Address[9]), .CEA(OutClockEn), .CLKA(OutClock), .OCEA(OutClockEn),
        .WEA(scuba_vlo), .CSA0(scuba_vlo), .CSA1(scuba_vlo), .CSA2(scuba_vlo),
        .RSTA(Reset), .DIB0(scuba_vlo), .DIB1(scuba_vlo), .DIB2(scuba_vlo),
        .DIB3(scuba_vlo), .DIB4(scuba_vlo), .DIB5(scuba_vlo), .DIB6(scuba_vlo),
        .DIB7(scuba_vlo), .DIB8(scuba_vlo), .DIB9(scuba_vlo), .DIB10(scuba_vlo),
        .DIB11(scuba_vlo), .DIB12(scuba_vlo), .DIB13(scuba_vlo), .DIB14(scuba_vlo),
        .DIB15(scuba_vlo), .DIB16(scuba_vlo), .DIB17(scuba_vlo), .ADB0(scuba_vlo),
        .ADB1(scuba_vlo), .ADB2(scuba_vlo), .ADB3(scuba_vlo), .ADB4(scuba_vlo),
        .ADB5(scuba_vlo), .ADB6(scuba_vlo), .ADB7(scuba_vlo), .ADB8(scuba_vlo),
        .ADB9(scuba_vlo), .ADB10(scuba_vlo), .ADB11(scuba_vlo), .ADB12(scuba_vlo),
        .ADB13(scuba_vlo), .CEB(scuba_vhi), .CLKB(scuba_vlo), .OCEB(scuba_vhi),
        .WEB(scuba_vlo), .CSB0(scuba_vlo), .CSB1(scuba_vlo), .CSB2(scuba_vlo),
        .RSTB(scuba_vlo), .DOA0(Q[0]), .DOA1(Q[1]), .DOA2(Q[2]), .DOA3(Q[3]),
        .DOA4(Q[4]), .DOA5(Q[5]), .DOA6(Q[6]), .DOA7(Q[7]), .DOA8(Q[8]),
        .DOA9(Q[9]), .DOA10(Q[10]), .DOA11(Q[11]), .DOA12(Q[12]), .DOA13(Q[13]),
        .DOA14(Q[14]), .DOA15(Q[15]), .DOA16(), .DOA17(), .DOB0(), .DOB1(),
        .DOB2(), .DOB3(), .DOB4(), .DOB5(), .DOB6(), .DOB7(), .DOB8(), .DOB9(),
        .DOB10(), .DOB11(), .DOB12(), .DOB13(), .DOB14(), .DOB15(), .DOB16(),
        .DOB17())
             /* synthesis MEM_LPC_FILE="biosrom.lpc" */
             /* synthesis MEM_INIT_FILE="biosrom.d16" */
             /* synthesis RESETMODE="SYNC" */;
    // exemplar begin
    // exemplar attribute biosrom_0_0_0 MEM_LPC_FILE biosrom.lpc
    // exemplar attribute biosrom_0_0_0 MEM_INIT_FILE biosrom.d16
    // exemplar attribute biosrom_0_0_0 RESETMODE SYNC
    // exemplar end
endmodule