module outputs
  wire [130 : 0] lookup;
  wire RDY_flush, RDY_insert, RDY_lookup;
  // register rg_flushing
  reg rg_flushing;
  wire rg_flushing$D_IN, rg_flushing$EN;
  // register tlb0_valids_0
  reg tlb0_valids_0;
  wire tlb0_valids_0$D_IN, tlb0_valids_0$EN;
  // register tlb0_valids_1
  reg tlb0_valids_1;
  wire tlb0_valids_1$D_IN, tlb0_valids_1$EN;
  // register tlb0_valids_10
  reg tlb0_valids_10;
  wire tlb0_valids_10$D_IN, tlb0_valids_10$EN;
  // register tlb0_valids_11
  reg tlb0_valids_11;
  wire tlb0_valids_11$D_IN, tlb0_valids_11$EN;
  // register tlb0_valids_12
  reg tlb0_valids_12;
  wire tlb0_valids_12$D_IN, tlb0_valids_12$EN;
  // register tlb0_valids_13
  reg tlb0_valids_13;
  wire tlb0_valids_13$D_IN, tlb0_valids_13$EN;
  // register tlb0_valids_14
  reg tlb0_valids_14;
  wire tlb0_valids_14$D_IN, tlb0_valids_14$EN;
  // register tlb0_valids_15
  reg tlb0_valids_15;
  wire tlb0_valids_15$D_IN, tlb0_valids_15$EN;
  // register tlb0_valids_2
  reg tlb0_valids_2;
  wire tlb0_valids_2$D_IN, tlb0_valids_2$EN;
  // register tlb0_valids_3
  reg tlb0_valids_3;
  wire tlb0_valids_3$D_IN, tlb0_valids_3$EN;
  // register tlb0_valids_4
  reg tlb0_valids_4;
  wire tlb0_valids_4$D_IN, tlb0_valids_4$EN;
  // register tlb0_valids_5
  reg tlb0_valids_5;
  wire tlb0_valids_5$D_IN, tlb0_valids_5$EN;
  // register tlb0_valids_6
  reg tlb0_valids_6;
  wire tlb0_valids_6$D_IN, tlb0_valids_6$EN;
  // register tlb0_valids_7
  reg tlb0_valids_7;
  wire tlb0_valids_7$D_IN, tlb0_valids_7$EN;
  // register tlb0_valids_8
  reg tlb0_valids_8;
  wire tlb0_valids_8$D_IN, tlb0_valids_8$EN;
  // register tlb0_valids_9
  reg tlb0_valids_9;
  wire tlb0_valids_9$D_IN, tlb0_valids_9$EN;
  // register tlb1_valids_0
  reg tlb1_valids_0;
  wire tlb1_valids_0$D_IN, tlb1_valids_0$EN;
  // register tlb1_valids_1
  reg tlb1_valids_1;
  wire tlb1_valids_1$D_IN, tlb1_valids_1$EN;
  // register tlb1_valids_2
  reg tlb1_valids_2;
  wire tlb1_valids_2$D_IN, tlb1_valids_2$EN;
  // register tlb1_valids_3
  reg tlb1_valids_3;
  wire tlb1_valids_3$D_IN, tlb1_valids_3$EN;
  // register tlb1_valids_4
  reg tlb1_valids_4;
  wire tlb1_valids_4$D_IN, tlb1_valids_4$EN;
  // register tlb1_valids_5
  reg tlb1_valids_5;
  wire tlb1_valids_5$D_IN, tlb1_valids_5$EN;
  // register tlb1_valids_6
  reg tlb1_valids_6;
  wire tlb1_valids_6$D_IN, tlb1_valids_6$EN;
  // register tlb1_valids_7
  reg tlb1_valids_7;
  wire tlb1_valids_7$D_IN, tlb1_valids_7$EN;
  // register tlb2_valids_0
  reg tlb2_valids_0;
  wire tlb2_valids_0$D_IN, tlb2_valids_0$EN;
  // register tlb2_valids_1
  reg tlb2_valids_1;
  wire tlb2_valids_1$D_IN, tlb2_valids_1$EN;
  // register tlb2_valids_2
  reg tlb2_valids_2;
  wire tlb2_valids_2$D_IN, tlb2_valids_2$EN;
  // register tlb2_valids_3
  reg tlb2_valids_3;
  wire tlb2_valids_3$D_IN, tlb2_valids_3$EN;
  // ports of submodule tlb0_entries
  wire [166 : 0] tlb0_entries$D_IN, tlb0_entries$D_OUT_1;
  wire [3 : 0] tlb0_entries$ADDR_1,
	       tlb0_entries$ADDR_2,
	       tlb0_entries$ADDR_3,
	       tlb0_entries$ADDR_4,
	       tlb0_entries$ADDR_5,
	       tlb0_entries$ADDR_IN;
  wire tlb0_entries$WE;
  // ports of submodule tlb1_entries
  wire [158 : 0] tlb1_entries$D_IN, tlb1_entries$D_OUT_1;
  wire [2 : 0] tlb1_entries$ADDR_1,
	       tlb1_entries$ADDR_2,
	       tlb1_entries$ADDR_3,
	       tlb1_entries$ADDR_4,
	       tlb1_entries$ADDR_5,
	       tlb1_entries$ADDR_IN;
  wire tlb1_entries$WE;
  // ports of submodule tlb2_entries
  wire [150 : 0] tlb2_entries$D_IN, tlb2_entries$D_OUT_1;
  wire [1 : 0] tlb2_entries$ADDR_1,
	       tlb2_entries$ADDR_2,
	       tlb2_entries$ADDR_3,
	       tlb2_entries$ADDR_4,
	       tlb2_entries$ADDR_5,
	       tlb2_entries$ADDR_IN;
  wire tlb2_entries$WE;
  // rule scheduling signals
  wire CAN_FIRE_RL_rl_initialize,
       CAN_FIRE_flush,
       CAN_FIRE_insert,
       WILL_FIRE_RL_rl_initialize,
       WILL_FIRE_flush,
       WILL_FIRE_insert;
  // inputs to muxes for submodule ports
  wire MUX_tlb0_valids_0$write_1__SEL_1,
       MUX_tlb0_valids_1$write_1__SEL_1,
       MUX_tlb0_valids_10$write_1__SEL_1,
       MUX_tlb0_valids_11$write_1__SEL_1,
       MUX_tlb0_valids_12$write_1__SEL_1,
       MUX_tlb0_valids_13$write_1__SEL_1,
       MUX_tlb0_valids_14$write_1__SEL_1,
       MUX_tlb0_valids_15$write_1__SEL_1,
       MUX_tlb0_valids_2$write_1__SEL_1,
       MUX_tlb0_valids_3$write_1__SEL_1,
       MUX_tlb0_valids_4$write_1__SEL_1,
       MUX_tlb0_valids_5$write_1__SEL_1,
       MUX_tlb0_valids_6$write_1__SEL_1,
       MUX_tlb0_valids_7$write_1__SEL_1,
       MUX_tlb0_valids_8$write_1__SEL_1,
       MUX_tlb0_valids_9$write_1__SEL_1,
       MUX_tlb1_valids_0$write_1__SEL_1,
       MUX_tlb1_valids_1$write_1__SEL_1,
       MUX_tlb1_valids_2$write_1__SEL_1,
       MUX_tlb1_valids_3$write_1__SEL_1,
       MUX_tlb1_valids_4$write_1__SEL_1,
       MUX_tlb1_valids_5$write_1__SEL_1,
       MUX_tlb1_valids_6$write_1__SEL_1,
       MUX_tlb1_valids_7$write_1__SEL_1,
       MUX_tlb2_valids_0$write_1__SEL_1,
       MUX_tlb2_valids_1$write_1__SEL_1,
       MUX_tlb2_valids_2$write_1__SEL_1,
       MUX_tlb2_valids_3$write_1__SEL_1;
  // remaining internal signals
  reg SEL_ARR_tlb0_valids_0_tlb0_valids_1_tlb0_valid_ETC___d20,
      SEL_ARR_tlb1_valids_0_1_tlb1_valids_1_2_tlb1_v_ETC___d41,
      SEL_ARR_tlb2_valids_0_3_tlb2_valids_1_4_tlb2_v_ETC___d59;
  wire [129 : 0] IF_SEL_ARR_tlb0_valids_0_tlb0_valids_1_tlb0_va_ETC___d85,
		 IF_SEL_ARR_tlb1_valids_0_1_tlb1_valids_1_2_tlb_ETC___d79,
		 IF_SEL_ARR_tlb2_valids_0_3_tlb2_valids_1_4_tlb_ETC___d84;
  wire [63 : 0] x__h6482, x__h6502;
  wire SEL_ARR_tlb0_valids_0_tlb0_valids_1_tlb0_valid_ETC___d26,
       SEL_ARR_tlb0_valids_0_tlb0_valids_1_tlb0_valid_ETC___d52,
       SEL_ARR_tlb0_valids_0_tlb0_valids_1_tlb0_valid_ETC___d70,
       SEL_ARR_tlb1_valids_0_1_tlb1_valids_1_2_tlb1_v_ETC___d47,
       SEL_ARR_tlb2_valids_0_3_tlb2_valids_1_4_tlb2_v_ETC___d65;
  // action method flush
  assign RDY_flush = 1'd1 ;
  assign CAN_FIRE_flush = 1'd1 ;
  assign WILL_FIRE_flush = EN_flush ;
  // value method lookup
  assign lookup =
	     { SEL_ARR_tlb0_valids_0_tlb0_valids_1_tlb0_valid_ETC___d70,
	       IF_SEL_ARR_tlb0_valids_0_tlb0_valids_1_tlb0_va_ETC___d85 } ;
  assign RDY_lookup = !rg_flushing ;
  // action method insert
  assign RDY_insert = !rg_flushing ;
  assign CAN_FIRE_insert = !rg_flushing ;
  assign WILL_FIRE_insert = EN_insert ;
  // submodule tlb0_entries
  RegFile #(.addr_width(32'd4),
	    .data_width(32'd167),
	    .lo(4'h0),
	    .hi(4'd15)) tlb0_entries(.CLK(CLK),
				     .ADDR_1(tlb0_entries$ADDR_1),
				     .ADDR_2(tlb0_entries$ADDR_2),
				     .ADDR_3(tlb0_entries$ADDR_3),
				     .ADDR_4(tlb0_entries$ADDR_4),
				     .ADDR_5(tlb0_entries$ADDR_5),
				     .ADDR_IN(tlb0_entries$ADDR_IN),
				     .D_IN(tlb0_entries$D_IN),
				     .WE(tlb0_entries$WE),
				     .D_OUT_1(tlb0_entries$D_OUT_1),
				     .D_OUT_2(),
				     .D_OUT_3(),
				     .D_OUT_4(),
				     .D_OUT_5());
  // submodule tlb1_entries
  RegFile #(.addr_width(32'd3),
	    .data_width(32'd159),
	    .lo(3'h0),
	    .hi(3'd7)) tlb1_entries(.CLK(CLK),
				    .ADDR_1(tlb1_entries$ADDR_1),
				    .ADDR_2(tlb1_entries$ADDR_2),
				    .ADDR_3(tlb1_entries$ADDR_3),
				    .ADDR_4(tlb1_entries$ADDR_4),
				    .ADDR_5(tlb1_entries$ADDR_5),
				    .ADDR_IN(tlb1_entries$ADDR_IN),
				    .D_IN(tlb1_entries$D_IN),
				    .WE(tlb1_entries$WE),
				    .D_OUT_1(tlb1_entries$D_OUT_1),
				    .D_OUT_2(),
				    .D_OUT_3(),
				    .D_OUT_4(),
				    .D_OUT_5());
  // submodule tlb2_entries
  RegFile #(.addr_width(32'd2),
	    .data_width(32'd151),
	    .lo(2'h0),
	    .hi(2'd3)) tlb2_entries(.CLK(CLK),
				    .ADDR_1(tlb2_entries$ADDR_1),
				    .ADDR_2(tlb2_entries$ADDR_2),
				    .ADDR_3(tlb2_entries$ADDR_3),
				    .ADDR_4(tlb2_entries$ADDR_4),
				    .ADDR_5(tlb2_entries$ADDR_5),
				    .ADDR_IN(tlb2_entries$ADDR_IN),
				    .D_IN(tlb2_entries$D_IN),
				    .WE(tlb2_entries$WE),
				    .D_OUT_1(tlb2_entries$D_OUT_1),
				    .D_OUT_2(),
				    .D_OUT_3(),
				    .D_OUT_4(),
				    .D_OUT_5());
  // rule RL_rl_initialize
  assign CAN_FIRE_RL_rl_initialize = rg_flushing ;
  assign WILL_FIRE_RL_rl_initialize = rg_flushing ;
  // inputs to muxes for submodule ports
  assign MUX_tlb0_valids_0$write_1__SEL_1 =
	     EN_insert && insert_vpn[3:0] == 4'd0 && insert_level == 2'd0 ;
  assign MUX_tlb0_valids_1$write_1__SEL_1 =
	     EN_insert && insert_vpn[3:0] == 4'd1 && insert_level == 2'd0 ;
  assign MUX_tlb0_valids_10$write_1__SEL_1 =
	     EN_insert && insert_vpn[3:0] == 4'd10 && insert_level == 2'd0 ;
  assign MUX_tlb0_valids_11$write_1__SEL_1 =
	     EN_insert && insert_vpn[3:0] == 4'd11 && insert_level == 2'd0 ;
  assign MUX_tlb0_valids_12$write_1__SEL_1 =
	     EN_insert && insert_vpn[3:0] == 4'd12 && insert_level == 2'd0 ;
  assign MUX_tlb0_valids_13$write_1__SEL_1 =
	     EN_insert && insert_vpn[3:0] == 4'd13 && insert_level == 2'd0 ;
  assign MUX_tlb0_valids_14$write_1__SEL_1 =
	     EN_insert && insert_vpn[3:0] == 4'd14 && insert_level == 2'd0 ;
  assign MUX_tlb0_valids_15$write_1__SEL_1 =
	     EN_insert && insert_vpn[3:0] == 4'd15 && insert_level == 2'd0 ;
  assign MUX_tlb0_valids_2$write_1__SEL_1 =
	     EN_insert && insert_vpn[3:0] == 4'd2 && insert_level == 2'd0 ;
  assign MUX_tlb0_valids_3$write_1__SEL_1 =
	     EN_insert && insert_vpn[3:0] == 4'd3 && insert_level == 2'd0 ;
  assign MUX_tlb0_valids_4$write_1__SEL_1 =
	     EN_insert && insert_vpn[3:0] == 4'd4 && insert_level == 2'd0 ;
  assign MUX_tlb0_valids_5$write_1__SEL_1 =
	     EN_insert && insert_vpn[3:0] == 4'd5 && insert_level == 2'd0 ;
  assign MUX_tlb0_valids_6$write_1__SEL_1 =
	     EN_insert && insert_vpn[3:0] == 4'd6 && insert_level == 2'd0 ;
  assign MUX_tlb0_valids_7$write_1__SEL_1 =
	     EN_insert && insert_vpn[3:0] == 4'd7 && insert_level == 2'd0 ;
  assign MUX_tlb0_valids_8$write_1__SEL_1 =
	     EN_insert && insert_vpn[3:0] == 4'd8 && insert_level == 2'd0 ;
  assign MUX_tlb0_valids_9$write_1__SEL_1 =
	     EN_insert && insert_vpn[3:0] == 4'd9 && insert_level == 2'd0 ;
  assign MUX_tlb1_valids_0$write_1__SEL_1 =
	     EN_insert && insert_vpn[11:9] == 3'd0 && insert_level == 2'd1 ;
  assign MUX_tlb1_valids_1$write_1__SEL_1 =
	     EN_insert && insert_vpn[11:9] == 3'd1 && insert_level == 2'd1 ;
  assign MUX_tlb1_valids_2$write_1__SEL_1 =
	     EN_insert && insert_vpn[11:9] == 3'd2 && insert_level == 2'd1 ;
  assign MUX_tlb1_valids_3$write_1__SEL_1 =
	     EN_insert && insert_vpn[11:9] == 3'd3 && insert_level == 2'd1 ;
  assign MUX_tlb1_valids_4$write_1__SEL_1 =
	     EN_insert && insert_vpn[11:9] == 3'd4 && insert_level == 2'd1 ;
  assign MUX_tlb1_valids_5$write_1__SEL_1 =
	     EN_insert && insert_vpn[11:9] == 3'd5 && insert_level == 2'd1 ;
  assign MUX_tlb1_valids_6$write_1__SEL_1 =
	     EN_insert && insert_vpn[11:9] == 3'd6 && insert_level == 2'd1 ;
  assign MUX_tlb1_valids_7$write_1__SEL_1 =
	     EN_insert && insert_vpn[11:9] == 3'd7 && insert_level == 2'd1 ;
  assign MUX_tlb2_valids_0$write_1__SEL_1 =
	     EN_insert && insert_vpn[19:18] == 2'd0 && insert_level != 2'd0 &&
	     insert_level != 2'd1 ;
  assign MUX_tlb2_valids_1$write_1__SEL_1 =
	     EN_insert && insert_vpn[19:18] == 2'd1 && insert_level != 2'd0 &&
	     insert_level != 2'd1 ;
  assign MUX_tlb2_valids_2$write_1__SEL_1 =
	     EN_insert && insert_vpn[19:18] == 2'd2 && insert_level != 2'd0 &&
	     insert_level != 2'd1 ;
  assign MUX_tlb2_valids_3$write_1__SEL_1 =
	     EN_insert && insert_vpn[19:18] == 2'd3 && insert_level != 2'd0 &&
	     insert_level != 2'd1 ;
  // register rg_flushing
  assign rg_flushing$D_IN = EN_flush ;
  assign rg_flushing$EN = rg_flushing || EN_flush ;
  // register tlb0_valids_0
  assign tlb0_valids_0$D_IN = MUX_tlb0_valids_0$write_1__SEL_1 ;
  assign tlb0_valids_0$EN =
	     EN_insert && insert_vpn[3:0] == 4'd0 && insert_level == 2'd0 ||
	     rg_flushing ;
  // register tlb0_valids_1
  assign tlb0_valids_1$D_IN = MUX_tlb0_valids_1$write_1__SEL_1 ;
  assign tlb0_valids_1$EN =
	     EN_insert && insert_vpn[3:0] == 4'd1 && insert_level == 2'd0 ||
	     rg_flushing ;
  // register tlb0_valids_10
  assign tlb0_valids_10$D_IN = MUX_tlb0_valids_10$write_1__SEL_1 ;
  assign tlb0_valids_10$EN =
	     EN_insert && insert_vpn[3:0] == 4'd10 && insert_level == 2'd0 ||
	     rg_flushing ;
  // register tlb0_valids_11
  assign tlb0_valids_11$D_IN = MUX_tlb0_valids_11$write_1__SEL_1 ;
  assign tlb0_valids_11$EN =
	     EN_insert && insert_vpn[3:0] == 4'd11 && insert_level == 2'd0 ||
	     rg_flushing ;
  // register tlb0_valids_12
  assign tlb0_valids_12$D_IN = MUX_tlb0_valids_12$write_1__SEL_1 ;
  assign tlb0_valids_12$EN =
	     EN_insert && insert_vpn[3:0] == 4'd12 && insert_level == 2'd0 ||
	     rg_flushing ;
  // register tlb0_valids_13
  assign tlb0_valids_13$D_IN = MUX_tlb0_valids_13$write_1__SEL_1 ;
  assign tlb0_valids_13$EN =
	     EN_insert && insert_vpn[3:0] == 4'd13 && insert_level == 2'd0 ||
	     rg_flushing ;
  // register tlb0_valids_14
  assign tlb0_valids_14$D_IN = MUX_tlb0_valids_14$write_1__SEL_1 ;
  assign tlb0_valids_14$EN =
	     EN_insert && insert_vpn[3:0] == 4'd14 && insert_level == 2'd0 ||
	     rg_flushing ;
  // register tlb0_valids_15
  assign tlb0_valids_15$D_IN = MUX_tlb0_valids_15$write_1__SEL_1 ;
  assign tlb0_valids_15$EN =
	     EN_insert && insert_vpn[3:0] == 4'd15 && insert_level == 2'd0 ||
	     rg_flushing ;
  // register tlb0_valids_2
  assign tlb0_valids_2$D_IN = MUX_tlb0_valids_2$write_1__SEL_1 ;
  assign tlb0_valids_2$EN =
	     EN_insert && insert_vpn[3:0] == 4'd2 && insert_level == 2'd0 ||
	     rg_flushing ;
  // register tlb0_valids_3
  assign tlb0_valids_3$D_IN = MUX_tlb0_valids_3$write_1__SEL_1 ;
  assign tlb0_valids_3$EN =
	     EN_insert && insert_vpn[3:0] == 4'd3 && insert_level == 2'd0 ||
	     rg_flushing ;
  // register tlb0_valids_4
  assign tlb0_valids_4$D_IN = MUX_tlb0_valids_4$write_1__SEL_1 ;
  assign tlb0_valids_4$EN =
	     EN_insert && insert_vpn[3:0] == 4'd4 && insert_level == 2'd0 ||
	     rg_flushing ;
  // register tlb0_valids_5
  assign tlb0_valids_5$D_IN = MUX_tlb0_valids_5$write_1__SEL_1 ;
  assign tlb0_valids_5$EN =
	     EN_insert && insert_vpn[3:0] == 4'd5 && insert_level == 2'd0 ||
	     rg_flushing ;
  // register tlb0_valids_6
  assign tlb0_valids_6$D_IN = MUX_tlb0_valids_6$write_1__SEL_1 ;
  assign tlb0_valids_6$EN =
	     EN_insert && insert_vpn[3:0] == 4'd6 && insert_level == 2'd0 ||
	     rg_flushing ;
  // register tlb0_valids_7
  assign tlb0_valids_7$D_IN = MUX_tlb0_valids_7$write_1__SEL_1 ;
  assign tlb0_valids_7$EN =
	     EN_insert && insert_vpn[3:0] == 4'd7 && insert_level == 2'd0 ||
	     rg_flushing ;
  // register tlb0_valids_8
  assign tlb0_valids_8$D_IN = MUX_tlb0_valids_8$write_1__SEL_1 ;
  assign tlb0_valids_8$EN =
	     EN_insert && insert_vpn[3:0] == 4'd8 && insert_level == 2'd0 ||
	     rg_flushing ;
  // register tlb0_valids_9
  assign tlb0_valids_9$D_IN = MUX_tlb0_valids_9$write_1__SEL_1 ;
  assign tlb0_valids_9$EN =
	     EN_insert && insert_vpn[3:0] == 4'd9 && insert_level == 2'd0 ||
	     rg_flushing ;
  // register tlb1_valids_0
  assign tlb1_valids_0$D_IN = MUX_tlb1_valids_0$write_1__SEL_1 ;
  assign tlb1_valids_0$EN =
	     EN_insert && insert_vpn[11:9] == 3'd0 && insert_level == 2'd1 ||
	     rg_flushing ;
  // register tlb1_valids_1
  assign tlb1_valids_1$D_IN = MUX_tlb1_valids_1$write_1__SEL_1 ;
  assign tlb1_valids_1$EN =
	     EN_insert && insert_vpn[11:9] == 3'd1 && insert_level == 2'd1 ||
	     rg_flushing ;
  // register tlb1_valids_2
  assign tlb1_valids_2$D_IN = MUX_tlb1_valids_2$write_1__SEL_1 ;
  assign tlb1_valids_2$EN =
	     EN_insert && insert_vpn[11:9] == 3'd2 && insert_level == 2'd1 ||
	     rg_flushing ;
  // register tlb1_valids_3
  assign tlb1_valids_3$D_IN = MUX_tlb1_valids_3$write_1__SEL_1 ;
  assign tlb1_valids_3$EN =
	     EN_insert && insert_vpn[11:9] == 3'd3 && insert_level == 2'd1 ||
	     rg_flushing ;
  // register tlb1_valids_4
  assign tlb1_valids_4$D_IN = MUX_tlb1_valids_4$write_1__SEL_1 ;
  assign tlb1_valids_4$EN =
	     EN_insert && insert_vpn[11:9] == 3'd4 && insert_level == 2'd1 ||
	     rg_flushing ;
  // register tlb1_valids_5
  assign tlb1_valids_5$D_IN = MUX_tlb1_valids_5$write_1__SEL_1 ;
  assign tlb1_valids_5$EN =
	     EN_insert && insert_vpn[11:9] == 3'd5 && insert_level == 2'd1 ||
	     rg_flushing ;
  // register tlb1_valids_6
  assign tlb1_valids_6$D_IN = MUX_tlb1_valids_6$write_1__SEL_1 ;
  assign tlb1_valids_6$EN =
	     EN_insert && insert_vpn[11:9] == 3'd6 && insert_level == 2'd1 ||
	     rg_flushing ;
  // register tlb1_valids_7
  assign tlb1_valids_7$D_IN = MUX_tlb1_valids_7$write_1__SEL_1 ;
  assign tlb1_valids_7$EN =
	     EN_insert && insert_vpn[11:9] == 3'd7 && insert_level == 2'd1 ||
	     rg_flushing ;
  // register tlb2_valids_0
  assign tlb2_valids_0$D_IN = MUX_tlb2_valids_0$write_1__SEL_1 ;
  assign tlb2_valids_0$EN =
	     EN_insert && insert_vpn[19:18] == 2'd0 && insert_level != 2'd0 &&
	     insert_level != 2'd1 ||
	     rg_flushing ;
  // register tlb2_valids_1
  assign tlb2_valids_1$D_IN = MUX_tlb2_valids_1$write_1__SEL_1 ;
  assign tlb2_valids_1$EN =
	     EN_insert && insert_vpn[19:18] == 2'd1 && insert_level != 2'd0 &&
	     insert_level != 2'd1 ||
	     rg_flushing ;
  // register tlb2_valids_2
  assign tlb2_valids_2$D_IN = MUX_tlb2_valids_2$write_1__SEL_1 ;
  assign tlb2_valids_2$EN =
	     EN_insert && insert_vpn[19:18] == 2'd2 && insert_level != 2'd0 &&
	     insert_level != 2'd1 ||
	     rg_flushing ;
  // register tlb2_valids_3
  assign tlb2_valids_3$D_IN = MUX_tlb2_valids_3$write_1__SEL_1 ;
  assign tlb2_valids_3$EN =
	     EN_insert && insert_vpn[19:18] == 2'd3 && insert_level != 2'd0 &&
	     insert_level != 2'd1 ||
	     rg_flushing ;
  // submodule tlb0_entries
  assign tlb0_entries$ADDR_1 = lookup_vpn[3:0] ;
  assign tlb0_entries$ADDR_2 = 4'h0 ;
  assign tlb0_entries$ADDR_3 = 4'h0 ;
  assign tlb0_entries$ADDR_4 = 4'h0 ;
  assign tlb0_entries$ADDR_5 = 4'h0 ;
  assign tlb0_entries$ADDR_IN = insert_vpn[3:0] ;
  assign tlb0_entries$D_IN =
	     { insert_asid, insert_vpn[26:4], insert_pte, insert_pte_pa } ;
  assign tlb0_entries$WE = EN_insert && insert_level == 2'd0 ;
  // submodule tlb1_entries
  assign tlb1_entries$ADDR_1 = lookup_vpn[11:9] ;
  assign tlb1_entries$ADDR_2 = 3'h0 ;
  assign tlb1_entries$ADDR_3 = 3'h0 ;
  assign tlb1_entries$ADDR_4 = 3'h0 ;
  assign tlb1_entries$ADDR_5 = 3'h0 ;
  assign tlb1_entries$ADDR_IN = insert_vpn[11:9] ;
  assign tlb1_entries$D_IN =
	     { insert_asid, insert_vpn[26:12], insert_pte, insert_pte_pa } ;
  assign tlb1_entries$WE = EN_insert && insert_level == 2'd1 ;
  // submodule tlb2_entries
  assign tlb2_entries$ADDR_1 = lookup_vpn[19:18] ;
  assign tlb2_entries$ADDR_2 = 2'h0 ;
  assign tlb2_entries$ADDR_3 = 2'h0 ;
  assign tlb2_entries$ADDR_4 = 2'h0 ;
  assign tlb2_entries$ADDR_5 = 2'h0 ;
  assign tlb2_entries$ADDR_IN = insert_vpn[19:18] ;
  assign tlb2_entries$D_IN =
	     { insert_asid, insert_vpn[26:20], insert_pte, insert_pte_pa } ;
  assign tlb2_entries$WE =
	     EN_insert && insert_level != 2'd0 && insert_level != 2'd1 ;
  // remaining internal signals
  assign IF_SEL_ARR_tlb0_valids_0_tlb0_valids_1_tlb0_va_ETC___d85 =
	     { x__h6482, 2'd0, x__h6502 } |
	     IF_SEL_ARR_tlb1_valids_0_1_tlb1_valids_1_2_tlb_ETC___d79 |
	     IF_SEL_ARR_tlb2_valids_0_3_tlb2_valids_1_4_tlb_ETC___d84 ;
  assign IF_SEL_ARR_tlb1_valids_0_1_tlb1_valids_1_2_tlb_ETC___d79 =
	     (SEL_ARR_tlb1_valids_0_1_tlb1_valids_1_2_tlb1_v_ETC___d47 &&
	      tlb1_entries$D_OUT_1[142:128] == lookup_vpn[26:12]) ?
	       { tlb1_entries$D_OUT_1[127:64],
		 2'd1,
		 tlb1_entries$D_OUT_1[63:0] } :
	       130'd0 ;
  assign IF_SEL_ARR_tlb2_valids_0_3_tlb2_valids_1_4_tlb_ETC___d84 =
	     (SEL_ARR_tlb2_valids_0_3_tlb2_valids_1_4_tlb2_v_ETC___d65 &&
	      tlb2_entries$D_OUT_1[134:128] == lookup_vpn[26:20]) ?
	       { tlb2_entries$D_OUT_1[127:64],
		 2'd2,
		 tlb2_entries$D_OUT_1[63:0] } :
	       130'd0 ;
  assign SEL_ARR_tlb0_valids_0_tlb0_valids_1_tlb0_valid_ETC___d26 =
	     SEL_ARR_tlb0_valids_0_tlb0_valids_1_tlb0_valid_ETC___d20 &&
	     (tlb0_entries$D_OUT_1[166:151] == lookup_asid ||
	      tlb0_entries$D_OUT_1[69]) ;
  assign SEL_ARR_tlb0_valids_0_tlb0_valids_1_tlb0_valid_ETC___d52 =
	     (SEL_ARR_tlb0_valids_0_tlb0_valids_1_tlb0_valid_ETC___d26 &&
	      tlb0_entries$D_OUT_1[150:128] == lookup_vpn[26:4]) |
	     (SEL_ARR_tlb1_valids_0_1_tlb1_valids_1_2_tlb1_v_ETC___d47 &&
	      tlb1_entries$D_OUT_1[142:128] == lookup_vpn[26:12]) ;
  assign SEL_ARR_tlb0_valids_0_tlb0_valids_1_tlb0_valid_ETC___d70 =
	     SEL_ARR_tlb0_valids_0_tlb0_valids_1_tlb0_valid_ETC___d52 |
	     (SEL_ARR_tlb2_valids_0_3_tlb2_valids_1_4_tlb2_v_ETC___d65 &&
	      tlb2_entries$D_OUT_1[134:128] == lookup_vpn[26:20]) ;
  assign SEL_ARR_tlb1_valids_0_1_tlb1_valids_1_2_tlb1_v_ETC___d47 =
	     SEL_ARR_tlb1_valids_0_1_tlb1_valids_1_2_tlb1_v_ETC___d41 &&
	     (tlb1_entries$D_OUT_1[158:143] == lookup_asid ||
	      tlb1_entries$D_OUT_1[69]) ;
  assign SEL_ARR_tlb2_valids_0_3_tlb2_valids_1_4_tlb2_v_ETC___d65 =
	     SEL_ARR_tlb2_valids_0_3_tlb2_valids_1_4_tlb2_v_ETC___d59 &&
	     (tlb2_entries$D_OUT_1[150:135] == lookup_asid ||
	      tlb2_entries$D_OUT_1[69]) ;
  assign x__h6482 =
	     (SEL_ARR_tlb0_valids_0_tlb0_valids_1_tlb0_valid_ETC___d26 &&
	      tlb0_entries$D_OUT_1[150:128] == lookup_vpn[26:4]) ?
	       tlb0_entries$D_OUT_1[127:64] :
	       64'd0 ;
  assign x__h6502 =
	     (SEL_ARR_tlb0_valids_0_tlb0_valids_1_tlb0_valid_ETC___d26 &&
	      tlb0_entries$D_OUT_1[150:128] == lookup_vpn[26:4]) ?
	       tlb0_entries$D_OUT_1[63:0] :
	       64'd0 ;
  always@(lookup_vpn or
	  tlb0_valids_0 or
	  tlb0_valids_1 or
	  tlb0_valids_2 or
	  tlb0_valids_3 or
	  tlb0_valids_4 or
	  tlb0_valids_5 or
	  tlb0_valids_6 or
	  tlb0_valids_7 or
	  tlb0_valids_8 or
	  tlb0_valids_9 or
	  tlb0_valids_10 or
	  tlb0_valids_11 or
	  tlb0_valids_12 or
	  tlb0_valids_13 or tlb0_valids_14 or tlb0_valids_15)
  begin
    case (lookup_vpn[3:0])
      4'd0:
	  SEL_ARR_tlb0_valids_0_tlb0_valids_1_tlb0_valid_ETC___d20 =
	      tlb0_valids_0;
      4'd1:
	  SEL_ARR_tlb0_valids_0_tlb0_valids_1_tlb0_valid_ETC___d20 =
	      tlb0_valids_1;
      4'd2:
	  SEL_ARR_tlb0_valids_0_tlb0_valids_1_tlb0_valid_ETC___d20 =
	      tlb0_valids_2;
      4'd3:
	  SEL_ARR_tlb0_valids_0_tlb0_valids_1_tlb0_valid_ETC___d20 =
	      tlb0_valids_3;
      4'd4:
	  SEL_ARR_tlb0_valids_0_tlb0_valids_1_tlb0_valid_ETC___d20 =
	      tlb0_valids_4;
      4'd5:
	  SEL_ARR_tlb0_valids_0_tlb0_valids_1_tlb0_valid_ETC___d20 =
	      tlb0_valids_5;
      4'd6:
	  SEL_ARR_tlb0_valids_0_tlb0_valids_1_tlb0_valid_ETC___d20 =
	      tlb0_valids_6;
      4'd7:
	  SEL_ARR_tlb0_valids_0_tlb0_valids_1_tlb0_valid_ETC___d20 =
	      tlb0_valids_7;
      4'd8:
	  SEL_ARR_tlb0_valids_0_tlb0_valids_1_tlb0_valid_ETC___d20 =
	      tlb0_valids_8;
      4'd9:
	  SEL_ARR_tlb0_valids_0_tlb0_valids_1_tlb0_valid_ETC___d20 =
	      tlb0_valids_9;
      4'd10:
	  SEL_ARR_tlb0_valids_0_tlb0_valids_1_tlb0_valid_ETC___d20 =
	      tlb0_valids_10;
      4'd11:
	  SEL_ARR_tlb0_valids_0_tlb0_valids_1_tlb0_valid_ETC___d20 =
	      tlb0_valids_11;
      4'd12:
	  SEL_ARR_tlb0_valids_0_tlb0_valids_1_tlb0_valid_ETC___d20 =
	      tlb0_valids_12;
      4'd13:
	  SEL_ARR_tlb0_valids_0_tlb0_valids_1_tlb0_valid_ETC___d20 =
	      tlb0_valids_13;
      4'd14:
	  SEL_ARR_tlb0_valids_0_tlb0_valids_1_tlb0_valid_ETC___d20 =
	      tlb0_valids_14;
      4'd15:
	  SEL_ARR_tlb0_valids_0_tlb0_valids_1_tlb0_valid_ETC___d20 =
	      tlb0_valids_15;
    endcase
  end
  always@(lookup_vpn or
	  tlb1_valids_0 or
	  tlb1_valids_1 or
	  tlb1_valids_2 or
	  tlb1_valids_3 or
	  tlb1_valids_4 or tlb1_valids_5 or tlb1_valids_6 or tlb1_valids_7)
  begin
    case (lookup_vpn[11:9])
      3'd0:
	  SEL_ARR_tlb1_valids_0_1_tlb1_valids_1_2_tlb1_v_ETC___d41 =
	      tlb1_valids_0;
      3'd1:
	  SEL_ARR_tlb1_valids_0_1_tlb1_valids_1_2_tlb1_v_ETC___d41 =
	      tlb1_valids_1;
      3'd2:
	  SEL_ARR_tlb1_valids_0_1_tlb1_valids_1_2_tlb1_v_ETC___d41 =
	      tlb1_valids_2;
      3'd3:
	  SEL_ARR_tlb1_valids_0_1_tlb1_valids_1_2_tlb1_v_ETC___d41 =
	      tlb1_valids_3;
      3'd4:
	  SEL_ARR_tlb1_valids_0_1_tlb1_valids_1_2_tlb1_v_ETC___d41 =
	      tlb1_valids_4;
      3'd5:
	  SEL_ARR_tlb1_valids_0_1_tlb1_valids_1_2_tlb1_v_ETC___d41 =
	      tlb1_valids_5;
      3'd6:
	  SEL_ARR_tlb1_valids_0_1_tlb1_valids_1_2_tlb1_v_ETC___d41 =
	      tlb1_valids_6;
      3'd7:
	  SEL_ARR_tlb1_valids_0_1_tlb1_valids_1_2_tlb1_v_ETC___d41 =
	      tlb1_valids_7;
    endcase
  end
  always@(lookup_vpn or
	  tlb2_valids_0 or tlb2_valids_1 or tlb2_valids_2 or tlb2_valids_3)
  begin
    case (lookup_vpn[19:18])
      2'd0:
	  SEL_ARR_tlb2_valids_0_3_tlb2_valids_1_4_tlb2_v_ETC___d59 =
	      tlb2_valids_0;
      2'd1:
	  SEL_ARR_tlb2_valids_0_3_tlb2_valids_1_4_tlb2_v_ETC___d59 =
	      tlb2_valids_1;
      2'd2:
	  SEL_ARR_tlb2_valids_0_3_tlb2_valids_1_4_tlb2_v_ETC___d59 =
	      tlb2_valids_2;
      2'd3:
	  SEL_ARR_tlb2_valids_0_3_tlb2_valids_1_4_tlb2_v_ETC___d59 =
	      tlb2_valids_3;
    endcase
  end
  // handling of inlined registers
  always@(posedge CLK)
  begin
    if (RST_N == `BSV_RESET_VALUE)
      begin
        rg_flushing <= `BSV_ASSIGNMENT_DELAY 1'd1;
      end
    else
      begin
        if (rg_flushing$EN)
	  rg_flushing <= `BSV_ASSIGNMENT_DELAY rg_flushing$D_IN;
      end
    if (tlb0_valids_0$EN)
      tlb0_valids_0 <= `BSV_ASSIGNMENT_DELAY tlb0_valids_0$D_IN;
    if (tlb0_valids_1$EN)
      tlb0_valids_1 <= `BSV_ASSIGNMENT_DELAY tlb0_valids_1$D_IN;
    if (tlb0_valids_10$EN)
      tlb0_valids_10 <= `BSV_ASSIGNMENT_DELAY tlb0_valids_10$D_IN;
    if (tlb0_valids_11$EN)
      tlb0_valids_11 <= `BSV_ASSIGNMENT_DELAY tlb0_valids_11$D_IN;
    if (tlb0_valids_12$EN)
      tlb0_valids_12 <= `BSV_ASSIGNMENT_DELAY tlb0_valids_12$D_IN;
    if (tlb0_valids_13$EN)
      tlb0_valids_13 <= `BSV_ASSIGNMENT_DELAY tlb0_valids_13$D_IN;
    if (tlb0_valids_14$EN)
      tlb0_valids_14 <= `BSV_ASSIGNMENT_DELAY tlb0_valids_14$D_IN;
    if (tlb0_valids_15$EN)
      tlb0_valids_15 <= `BSV_ASSIGNMENT_DELAY tlb0_valids_15$D_IN;
    if (tlb0_valids_2$EN)
      tlb0_valids_2 <= `BSV_ASSIGNMENT_DELAY tlb0_valids_2$D_IN;
    if (tlb0_valids_3$EN)
      tlb0_valids_3 <= `BSV_ASSIGNMENT_DELAY tlb0_valids_3$D_IN;
    if (tlb0_valids_4$EN)
      tlb0_valids_4 <= `BSV_ASSIGNMENT_DELAY tlb0_valids_4$D_IN;
    if (tlb0_valids_5$EN)
      tlb0_valids_5 <= `BSV_ASSIGNMENT_DELAY tlb0_valids_5$D_IN;
    if (tlb0_valids_6$EN)
      tlb0_valids_6 <= `BSV_ASSIGNMENT_DELAY tlb0_valids_6$D_IN;
    if (tlb0_valids_7$EN)
      tlb0_valids_7 <= `BSV_ASSIGNMENT_DELAY tlb0_valids_7$D_IN;
    if (tlb0_valids_8$EN)
      tlb0_valids_8 <= `BSV_ASSIGNMENT_DELAY tlb0_valids_8$D_IN;
    if (tlb0_valids_9$EN)
      tlb0_valids_9 <= `BSV_ASSIGNMENT_DELAY tlb0_valids_9$D_IN;
    if (tlb1_valids_0$EN)
      tlb1_valids_0 <= `BSV_ASSIGNMENT_DELAY tlb1_valids_0$D_IN;
    if (tlb1_valids_1$EN)
      tlb1_valids_1 <= `BSV_ASSIGNMENT_DELAY tlb1_valids_1$D_IN;
    if (tlb1_valids_2$EN)
      tlb1_valids_2 <= `BSV_ASSIGNMENT_DELAY tlb1_valids_2$D_IN;
    if (tlb1_valids_3$EN)
      tlb1_valids_3 <= `BSV_ASSIGNMENT_DELAY tlb1_valids_3$D_IN;
    if (tlb1_valids_4$EN)
      tlb1_valids_4 <= `BSV_ASSIGNMENT_DELAY tlb1_valids_4$D_IN;
    if (tlb1_valids_5$EN)
      tlb1_valids_5 <= `BSV_ASSIGNMENT_DELAY tlb1_valids_5$D_IN;
    if (tlb1_valids_6$EN)
      tlb1_valids_6 <= `BSV_ASSIGNMENT_DELAY tlb1_valids_6$D_IN;
    if (tlb1_valids_7$EN)
      tlb1_valids_7 <= `BSV_ASSIGNMENT_DELAY tlb1_valids_7$D_IN;
    if (tlb2_valids_0$EN)
      tlb2_valids_0 <= `BSV_ASSIGNMENT_DELAY tlb2_valids_0$D_IN;
    if (tlb2_valids_1$EN)
      tlb2_valids_1 <= `BSV_ASSIGNMENT_DELAY tlb2_valids_1$D_IN;
    if (tlb2_valids_2$EN)
      tlb2_valids_2 <= `BSV_ASSIGNMENT_DELAY tlb2_valids_2$D_IN;
    if (tlb2_valids_3$EN)
      tlb2_valids_3 <= `BSV_ASSIGNMENT_DELAY tlb2_valids_3$D_IN;
  end
  // synopsys translate_off
  `ifdef BSV_NO_INITIAL_BLOCKS
  `else // not BSV_NO_INITIAL_BLOCKS
  initial
  begin
    rg_flushing = 1'h0;
    tlb0_valids_0 = 1'h0;
    tlb0_valids_1 = 1'h0;
    tlb0_valids_10 = 1'h0;
    tlb0_valids_11 = 1'h0;
    tlb0_valids_12 = 1'h0;
    tlb0_valids_13 = 1'h0;
    tlb0_valids_14 = 1'h0;
    tlb0_valids_15 = 1'h0;
    tlb0_valids_2 = 1'h0;
    tlb0_valids_3 = 1'h0;
    tlb0_valids_4 = 1'h0;
    tlb0_valids_5 = 1'h0;
    tlb0_valids_6 = 1'h0;
    tlb0_valids_7 = 1'h0;
    tlb0_valids_8 = 1'h0;
    tlb0_valids_9 = 1'h0;
    tlb1_valids_0 = 1'h0;
    tlb1_valids_1 = 1'h0;
    tlb1_valids_2 = 1'h0;
    tlb1_valids_3 = 1'h0;
    tlb1_valids_4 = 1'h0;
    tlb1_valids_5 = 1'h0;
    tlb1_valids_6 = 1'h0;
    tlb1_valids_7 = 1'h0;
    tlb2_valids_0 = 1'h0;
    tlb2_valids_1 = 1'h0;
    tlb2_valids_2 = 1'h0;
    tlb2_valids_3 = 1'h0;
  end
  `endif // BSV_NO_INITIAL_BLOCKS
  // synopsys translate_on
endmodule