module SCB_P4_v1_10_2 (
    sclk,
    interrupt,
    clock);
    output      sclk;
    output      interrupt;
    input       clock;
          wire [3:0] ss;
          wire  Net_88;
          wire  Net_84;
          wire  Net_149;
          wire  Net_150;
          wire  Net_152;
          wire  Net_453;
          wire  uncfg_rx_irq;
          wire  Net_427;
          wire  Net_436;
          wire  Net_449;
          wire  Net_433;
          wire  Net_373;
          wire  Net_452;
          wire  Net_459;
          wire  Net_458;
          wire  Net_430;
          wire  Net_237;
          wire  Net_413;
          wire  Net_244;
          wire  Net_422;
          wire  rx_irq;
          wire  Net_379;
          wire  Net_409;
          wire  Net_246;
          wire  Net_252;
          wire  Net_245;
          wire  Net_243;
          wire  Net_89;
          wire  Net_284;
          wire  Net_416;
          wire  Net_387;
          wire  Net_151;
          wire  Net_410;
    cy_m0s8_scb_v1_0 SCB (
        .rx(Net_244),
        .miso_m(Net_410),
        .clock(Net_237),
        .select_m(ss[3:0]),
        .sclk_m(Net_88),
        .mosi_s(Net_89),
        .select_s(Net_430),
        .sclk_s(Net_413),
        .mosi_m(Net_84),
        .scl(Net_149),
        .sda(Net_150),
        .tx(Net_151),
        .miso_s(Net_152),
        .interrupt(interrupt));
    defparam SCB.scb_mode = 2;
	wire [0:0] tmpOE__rx_net;
	wire [0:0] tmpIO_0__rx_net;
	wire [0:0] tmpINTERRUPT_0__rx_net;
	electrical [0:0] tmpSIOVREF__rx_net;
	cy_psoc3_pins_v1_10
		#(.id("43ec2fa1-bf22-4b71-9477-b6ca7b97f0b0/78e33e5d-45ea-4b75-88d5-73274e8a7ce4"),
		  .drive_mode(3'b001),
		  .ibuf_enabled(1'b1),
		  .init_dr_st(1'b0),
		  .input_clk_en(0),
		  .input_sync(1'b0),
		  .input_sync_mode(1'b0),
		  .intr_mode(2'b00),
		  .invert_in_clock(0),
		  .invert_in_clock_en(0),
		  .invert_in_reset(0),
		  .invert_out_clock(0),
		  .invert_out_clock_en(0),
		  .invert_out_reset(0),
		  .io_voltage(""),
		  .layout_mode("CONTIGUOUS"),
		  .oe_conn(1'b0),
		  .oe_reset(0),
		  .oe_sync(1'b0),
		  .output_clk_en(0),
		  .output_clock_mode(1'b0),
		  .output_conn(1'b0),
		  .output_mode(1'b0),
		  .output_reset(0),
		  .output_sync(1'b0),
		  .pa_in_clock(-1),
		  .pa_in_clock_en(-1),
		  .pa_in_reset(-1),
		  .pa_out_clock(-1),
		  .pa_out_clock_en(-1),
		  .pa_out_reset(-1),
		  .pin_aliases(""),
		  .pin_mode("I"),
		  .por_state(4),
		  .use_annotation(1'b0),
		  .sio_group_cnt(0),
		  .sio_hyst(1'b0),
		  .sio_ibuf(""),
		  .sio_info(2'b00),
		  .sio_obuf(""),
		  .sio_refsel(""),
		  .sio_vtrip(""),
		  .slew_rate(1'b0),
		  .spanning(0),
		  .vtrip(2'b00),
		  .width(1))
		rx
		 (.oe(tmpOE__rx_net),
		  .y({1'b0}),
		  .fb({Net_379}),
		  .io({tmpIO_0__rx_net[0:0]}),
		  .siovref(tmpSIOVREF__rx_net),
		  .interrupt({tmpINTERRUPT_0__rx_net[0:0]}),
		  .in_clock({1'b0}),
		  .in_clock_en({1'b1}),
		  .in_reset({1'b0}),
		  .out_clock({1'b0}),
		  .out_clock_en({1'b1}),
		  .out_reset({1'b0}));
	assign tmpOE__rx_net = (`CYDEV_CHIP_MEMBER_USED == `CYDEV_CHIP_MEMBER_3A && `CYDEV_CHIP_REVISION_USED < `CYDEV_CHIP_REVISION_3A_ES3) ? ~{1'b1} : {1'b1};
	cy_clock_v1_0
		#(.id("43ec2fa1-bf22-4b71-9477-b6ca7b97f0b0/29084e80-7594-46a9-94af-639e276dfc5f"),
		  .source_clock_id(""),
		  .divisor(0),
		  .period("8680555555.55556"),
		  .is_direct(0),
		  .is_digital(0))
		SCBCLK
		 (.clock_out(Net_284));
    assign sclk = Net_284 | Net_427;
    ZeroTerminal ZeroTerminal_7 (
        .z(Net_427));
	wire [0:0] tmpOE__tx_net;
	wire [0:0] tmpFB_0__tx_net;
	wire [0:0] tmpIO_0__tx_net;
	wire [0:0] tmpINTERRUPT_0__tx_net;
	electrical [0:0] tmpSIOVREF__tx_net;
	cy_psoc3_pins_v1_10
		#(.id("43ec2fa1-bf22-4b71-9477-b6ca7b97f0b0/23b8206d-1c77-4e61-be4a-b4037d5de5fc"),
		  .drive_mode(3'b110),
		  .ibuf_enabled(1'b1),
		  .init_dr_st(1'b1),
		  .input_clk_en(0),
		  .input_sync(1'b1),
		  .input_sync_mode(1'b0),
		  .intr_mode(2'b00),
		  .invert_in_clock(0),
		  .invert_in_clock_en(0),
		  .invert_in_reset(0),
		  .invert_out_clock(0),
		  .invert_out_clock_en(0),
		  .invert_out_reset(0),
		  .io_voltage(""),
		  .layout_mode("CONTIGUOUS"),
		  .oe_conn(1'b0),
		  .oe_reset(0),
		  .oe_sync(1'b0),
		  .output_clk_en(0),
		  .output_clock_mode(1'b0),
		  .output_conn(1'b1),
		  .output_mode(1'b0),
		  .output_reset(0),
		  .output_sync(1'b0),
		  .pa_in_clock(-1),
		  .pa_in_clock_en(-1),
		  .pa_in_reset(-1),
		  .pa_out_clock(-1),
		  .pa_out_clock_en(-1),
		  .pa_out_reset(-1),
		  .pin_aliases(""),
		  .pin_mode("O"),
		  .por_state(4),
		  .use_annotation(1'b0),
		  .sio_group_cnt(0),
		  .sio_hyst(1'b0),
		  .sio_ibuf(""),
		  .sio_info(2'b00),
		  .sio_obuf(""),
		  .sio_refsel(""),
		  .sio_vtrip(""),
		  .slew_rate(1'b0),
		  .spanning(0),
		  .vtrip(2'b10),
		  .width(1))
		tx
		 (.oe(tmpOE__tx_net),
		  .y({Net_151}),
		  .fb({tmpFB_0__tx_net[0:0]}),
		  .io({tmpIO_0__tx_net[0:0]}),
		  .siovref(tmpSIOVREF__tx_net),
		  .interrupt({tmpINTERRUPT_0__tx_net[0:0]}),
		  .in_clock({1'b0}),
		  .in_clock_en({1'b1}),
		  .in_reset({1'b0}),
		  .out_clock({1'b0}),
		  .out_clock_en({1'b1}),
		  .out_reset({1'b0}));
	assign tmpOE__tx_net = (`CYDEV_CHIP_MEMBER_USED == `CYDEV_CHIP_MEMBER_3A && `CYDEV_CHIP_REVISION_USED < `CYDEV_CHIP_REVISION_3A_ES3) ? ~{1'b1} : {1'b1};
	// miso_m_VM (cy_virtualmux_v1_0)
	assign Net_410 = Net_436;
	// mosi_s_VM (cy_virtualmux_v1_0)
	assign Net_89 = Net_449;
	// sclk_s_VM (cy_virtualmux_v1_0)
	assign Net_413 = Net_433;
	// clock_VM (cy_virtualmux_v1_0)
	assign Net_237 = Net_284;
	// rx_wake_VM (cy_virtualmux_v1_0)
	assign Net_373 = uncfg_rx_irq;
	// rx_VM (cy_virtualmux_v1_0)
	assign Net_244 = Net_379;
    ZeroTerminal ZeroTerminal_1 (
        .z(Net_433));
    ZeroTerminal ZeroTerminal_2 (
        .z(Net_436));
    ZeroTerminal ZeroTerminal_3 (
        .z(Net_449));
    ZeroTerminal ZeroTerminal_4 (
        .z(Net_452));
	// select_s_VM (cy_virtualmux_v1_0)
	assign Net_430 = Net_459;
    ZeroTerminal ZeroTerminal_5 (
        .z(Net_459));
endmodule