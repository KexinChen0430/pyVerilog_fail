module parse_instr (input [31:0] instr,
                    output      `ALL_SUPPORT_INSTR);
   wire                         rtype,regimm,cop0;
   wire [5:0]                  OpCode;
   wire [5:0]                  Funct;
   assign OpCode=instr[`OP];
   assign Funct=instr[`FUNCT];
   assign rtype=(OpCode==`RTYPE);
   assign add=rtype&(Funct==`ADD_R);
   assign addu=rtype&(Funct==`ADDU_R);
   assign sub=rtype&(Funct==`SUB_R);
   assign subu=rtype&(Funct==`SUBU_R);
   assign mult=rtype&(Funct==`MULT_R);
   assign multu=rtype&(Funct==`MULTU_R);
   assign div=rtype&(Funct==`DIV_R);
   assign divu=rtype&(Funct==`DIVU_R);
   assign slt=rtype&(Funct==`SLT_R);
   assign sltu=rtype&(Funct==`SLTU_R);
   assign sll=rtype&(Funct==`SLL_R);
   assign srl=rtype&(Funct==`SRL_R);
   assign sra=rtype&(Funct==`SRA_R);
   assign sllv=rtype&(Funct==`SLLV_R);
   assign srlv=rtype&(Funct==`SRLV_R);
   assign srav=rtype&(Funct==`SRAV_R);
   assign and_r=rtype&(Funct==`AND_R);
   assign or_r=rtype&(Funct==`OR_R);
   assign nor_r=rtype&(Funct==`NOR_R);
   assign xor_r=rtype&(Funct==`XOR_R);
   assign andi=(OpCode==`ANDI);
   assign ori=(OpCode==`ORI);
   assign lui=(OpCode==`LUI);
   assign xori=(OpCode==`XORI);
   assign lb=(OpCode==`LB);
   assign lbu=(OpCode==`LBU);
   assign lh=(OpCode==`LH);
   assign lhu=(OpCode==`LHU);
   assign lw=(OpCode==`LW);
   assign sb=(OpCode==`SB);
   assign sh=(OpCode==`SH);
   assign sw=(OpCode==`SW);
   assign slti=(OpCode==`SLTI);
   assign sltiu=(OpCode==`SLTIU);
   assign beq=(OpCode==`BEQ);
   assign bne=(OpCode==`BNE);
   assign blez=(OpCode==`BLEZ);
   assign bgtz=(OpCode==`BGTZ);
   assign regimm=(OpCode==`REGIMM);
   assign bltz=regimm&(instr[`RT]==`BLTZ);
   assign bgez=regimm&(instr[`RT]==`BGEZ);
   assign addi=(OpCode==`ADDI);
   assign addiu=(OpCode==`ADDIU);
   assign j=(OpCode==`J);
   assign jal=(OpCode==`JAL);
   assign jr=rtype&(Funct==`JR_R);
   assign jalr=rtype&(Funct==`JALR_R);
   assign mtlo=rtype&(Funct==`MTLO_R);
   assign mthi=rtype&(Funct==`MTHI_R);
   assign mflo=rtype&(Funct==`MFLO_R);
   assign mfhi=rtype&(Funct==`MFHI_R);
   assign cop0=(OpCode==`COP0);
   assign mtc0=cop0&(instr[`RS]==`MT);
   assign mfc0=cop0&(instr[`RS]==`MF);
   assign eret=cop0&(Funct==`ERET_R);
endmodule