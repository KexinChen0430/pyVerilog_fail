module mac_fixpt_tb
          (
          );
  reg  clk;
  reg  reset;
  wire enb;
  wire M_out_0_addr;  // ufix1
  wire M_out_0_lastAddr;  // ufix1
  reg  check1_done;  // ufix1
  wire snkDonen;
  wire resetn;
  wire tb_enb;
  wire rdEnb;
  wire M_out_0_done;  // ufix1
  wire M_out_0_done_enb;  // ufix1
  wire ce_out;
  wire rawData_M_0;  // ufix1
  reg  holdData_M_0;  // ufix1
  wire rawData_M_1;  // ufix1
  reg  holdData_M_1;  // ufix1
  wire rawData_M_2;  // ufix1
  reg  holdData_M_2;  // ufix1
  wire rawData_M_3;  // ufix1
  reg  holdData_M_3;  // ufix1
  wire rawData_M_4;  // ufix1
  reg  holdData_M_4;  // ufix1
  wire rawData_M_5;  // ufix1
  reg  holdData_M_5;  // ufix1
  wire rawData_M_6;  // ufix1
  reg  holdData_M_6;  // ufix1
  wire rawData_M_7;  // ufix1
  reg  holdData_M_7;  // ufix1
  wire rawData_M_8;  // ufix1
  reg  holdData_M_8;  // ufix1
  wire rawData_M_9;  // ufix1
  reg  holdData_M_9;  // ufix1
  wire rawData_M_10;  // ufix1
  reg  holdData_M_10;  // ufix1
  wire rawData_M_11;  // ufix1
  reg  holdData_M_11;  // ufix1
  wire rawData_M_12;  // ufix1
  reg  holdData_M_12;  // ufix1
  wire rawData_M_13;  // ufix1
  reg  holdData_M_13;  // ufix1
  wire rawData_M_14;  // ufix1
  reg  holdData_M_14;  // ufix1
  wire rawData_M_15;  // ufix1
  reg  holdData_M_15;  // ufix1
  wire rawData_M_16;  // ufix1
  reg  holdData_M_16;  // ufix1
  wire rawData_M_17;  // ufix1
  reg  holdData_M_17;  // ufix1
  wire rawData_M_18;  // ufix1
  reg  holdData_M_18;  // ufix1
  wire rawData_M_19;  // ufix1
  reg  holdData_M_19;  // ufix1
  wire rawData_M_20;  // ufix1
  reg  holdData_M_20;  // ufix1
  wire rawData_M_21;  // ufix1
  reg  holdData_M_21;  // ufix1
  wire rawData_M_22;  // ufix1
  reg  holdData_M_22;  // ufix1
  wire rawData_M_23;  // ufix1
  reg  holdData_M_23;  // ufix1
  wire rawData_M_24;  // ufix1
  reg  holdData_M_24;  // ufix1
  wire rawData_M_25;  // ufix1
  reg  holdData_M_25;  // ufix1
  wire rawData_M_26;  // ufix1
  reg  holdData_M_26;  // ufix1
  wire rawData_M_27;  // ufix1
  reg  holdData_M_27;  // ufix1
  wire rawData_M_28;  // ufix1
  reg  holdData_M_28;  // ufix1
  wire rawData_M_29;  // ufix1
  reg  holdData_M_29;  // ufix1
  wire rawData_M_30;  // ufix1
  reg  holdData_M_30;  // ufix1
  wire rawData_M_31;  // ufix1
  reg  holdData_M_31;  // ufix1
  wire rawData_M_32;  // ufix1
  reg  holdData_M_32;  // ufix1
  wire rawData_M_33;  // ufix1
  reg  holdData_M_33;  // ufix1
  wire rawData_M_34;  // ufix1
  reg  holdData_M_34;  // ufix1
  wire rawData_M_35;  // ufix1
  reg  holdData_M_35;  // ufix1
  wire rawData_M_36;  // ufix1
  reg  holdData_M_36;  // ufix1
  wire rawData_M_37;  // ufix1
  reg  holdData_M_37;  // ufix1
  wire rawData_M_38;  // ufix1
  reg  holdData_M_38;  // ufix1
  wire rawData_M_39;  // ufix1
  reg  holdData_M_39;  // ufix1
  wire rawData_M_40;  // ufix1
  reg  holdData_M_40;  // ufix1
  wire rawData_M_41;  // ufix1
  reg  holdData_M_41;  // ufix1
  wire rawData_M_42;  // ufix1
  reg  holdData_M_42;  // ufix1
  wire rawData_M_43;  // ufix1
  reg  holdData_M_43;  // ufix1
  wire rawData_M_44;  // ufix1
  reg  holdData_M_44;  // ufix1
  wire rawData_M_45;  // ufix1
  reg  holdData_M_45;  // ufix1
  wire rawData_M_46;  // ufix1
  reg  holdData_M_46;  // ufix1
  wire rawData_M_47;  // ufix1
  reg  holdData_M_47;  // ufix1
  wire rawData_M_48;  // ufix1
  reg  holdData_M_48;  // ufix1
  wire rawData_M_49;  // ufix1
  reg  holdData_M_49;  // ufix1
  wire rawData_M_50;  // ufix1
  reg  holdData_M_50;  // ufix1
  wire rawData_M_51;  // ufix1
  reg  holdData_M_51;  // ufix1
  wire rawData_M_52;  // ufix1
  reg  holdData_M_52;  // ufix1
  wire rawData_M_53;  // ufix1
  reg  holdData_M_53;  // ufix1
  wire rawData_M_54;  // ufix1
  reg  holdData_M_54;  // ufix1
  wire rawData_M_55;  // ufix1
  reg  holdData_M_55;  // ufix1
  wire rawData_M_56;  // ufix1
  reg  holdData_M_56;  // ufix1
  wire rawData_M_57;  // ufix1
  reg  holdData_M_57;  // ufix1
  wire rawData_M_58;  // ufix1
  reg  holdData_M_58;  // ufix1
  wire rawData_M_59;  // ufix1
  reg  holdData_M_59;  // ufix1
  wire rawData_M_60;  // ufix1
  reg  holdData_M_60;  // ufix1
  wire rawData_M_61;  // ufix1
  reg  holdData_M_61;  // ufix1
  wire rawData_M_62;  // ufix1
  reg  holdData_M_62;  // ufix1
  wire rawData_M_63;  // ufix1
  reg  holdData_M_63;  // ufix1
  wire rawData_N_0;  // ufix1
  reg  holdData_N_0;  // ufix1
  wire rawData_N_1;  // ufix1
  reg  holdData_N_1;  // ufix1
  wire rawData_N_2;  // ufix1
  reg  holdData_N_2;  // ufix1
  wire rawData_N_3;  // ufix1
  reg  holdData_N_3;  // ufix1
  wire rawData_N_4;  // ufix1
  reg  holdData_N_4;  // ufix1
  wire rawData_N_5;  // ufix1
  reg  holdData_N_5;  // ufix1
  wire rawData_N_6;  // ufix1
  reg  holdData_N_6;  // ufix1
  wire [13:0] rawData_W_0;  // ufix14_En13
  reg [13:0] holdData_W_0;  // ufix14_En13
  wire [13:0] rawData_W_1;  // ufix14_En13
  reg [13:0] holdData_W_1;  // ufix14_En13
  wire [13:0] rawData_W_2;  // ufix14_En13
  reg [13:0] holdData_W_2;  // ufix14_En13
  wire [13:0] rawData_W_3;  // ufix14_En13
  reg [13:0] holdData_W_3;  // ufix14_En13
  wire [13:0] rawData_W_4;  // ufix14_En13
  reg [13:0] holdData_W_4;  // ufix14_En13
  wire [13:0] rawData_W_5;  // ufix14_En13
  reg [13:0] holdData_W_5;  // ufix14_En13
  wire [13:0] rawData_W_6;  // ufix14_En13
  reg [13:0] holdData_W_6;  // ufix14_En13
  wire [6:0] rawData_Tm;  // ufix7
  reg [6:0] holdData_Tm;  // ufix7
  wire [2:0] rawData_Tn;  // ufix3
  reg [2:0] holdData_Tn;  // ufix3
  reg  M_0_offset;  // ufix1
  wire M_0_1;  // ufix1
  reg  M_1_offset;  // ufix1
  wire M_1_1;  // ufix1
  reg  M_2_offset;  // ufix1
  wire M_2_1;  // ufix1
  reg  M_3_offset;  // ufix1
  wire M_3_1;  // ufix1
  reg  M_4_offset;  // ufix1
  wire M_4_1;  // ufix1
  reg  M_5_offset;  // ufix1
  wire M_5_1;  // ufix1
  reg  M_6_offset;  // ufix1
  wire M_6_1;  // ufix1
  reg  M_7_offset;  // ufix1
  wire M_7_1;  // ufix1
  reg  M_8_offset;  // ufix1
  wire M_8_1;  // ufix1
  reg  M_9_offset;  // ufix1
  wire M_9_1;  // ufix1
  reg  M_10_offset;  // ufix1
  wire M_10_1;  // ufix1
  reg  M_11_offset;  // ufix1
  wire M_11_1;  // ufix1
  reg  M_12_offset;  // ufix1
  wire M_12_1;  // ufix1
  reg  M_13_offset;  // ufix1
  wire M_13_1;  // ufix1
  reg  M_14_offset;  // ufix1
  wire M_14_1;  // ufix1
  reg  M_15_offset;  // ufix1
  wire M_15_1;  // ufix1
  reg  M_16_offset;  // ufix1
  wire M_16_1;  // ufix1
  reg  M_17_offset;  // ufix1
  wire M_17_1;  // ufix1
  reg  M_18_offset;  // ufix1
  wire M_18_1;  // ufix1
  reg  M_19_offset;  // ufix1
  wire M_19_1;  // ufix1
  reg  M_20_offset;  // ufix1
  wire M_20_1;  // ufix1
  reg  M_21_offset;  // ufix1
  wire M_21_1;  // ufix1
  reg  M_22_offset;  // ufix1
  wire M_22_1;  // ufix1
  reg  M_23_offset;  // ufix1
  wire M_23_1;  // ufix1
  reg  M_24_offset;  // ufix1
  wire M_24_1;  // ufix1
  reg  M_25_offset;  // ufix1
  wire M_25_1;  // ufix1
  reg  M_26_offset;  // ufix1
  wire M_26_1;  // ufix1
  reg  M_27_offset;  // ufix1
  wire M_27_1;  // ufix1
  reg  M_28_offset;  // ufix1
  wire M_28_1;  // ufix1
  reg  M_29_offset;  // ufix1
  wire M_29_1;  // ufix1
  reg  M_30_offset;  // ufix1
  wire M_30_1;  // ufix1
  reg  M_31_offset;  // ufix1
  wire M_31_1;  // ufix1
  reg  M_32_offset;  // ufix1
  wire M_32_1;  // ufix1
  reg  M_33_offset;  // ufix1
  wire M_33_1;  // ufix1
  reg  M_34_offset;  // ufix1
  wire M_34_1;  // ufix1
  reg  M_35_offset;  // ufix1
  wire M_35_1;  // ufix1
  reg  M_36_offset;  // ufix1
  wire M_36_1;  // ufix1
  reg  M_37_offset;  // ufix1
  wire M_37_1;  // ufix1
  reg  M_38_offset;  // ufix1
  wire M_38_1;  // ufix1
  reg  M_39_offset;  // ufix1
  wire M_39_1;  // ufix1
  reg  M_40_offset;  // ufix1
  wire M_40_1;  // ufix1
  reg  M_41_offset;  // ufix1
  wire M_41_1;  // ufix1
  reg  M_42_offset;  // ufix1
  wire M_42_1;  // ufix1
  reg  M_43_offset;  // ufix1
  wire M_43_1;  // ufix1
  reg  M_44_offset;  // ufix1
  wire M_44_1;  // ufix1
  reg  M_45_offset;  // ufix1
  wire M_45_1;  // ufix1
  reg  M_46_offset;  // ufix1
  wire M_46_1;  // ufix1
  reg  M_47_offset;  // ufix1
  wire M_47_1;  // ufix1
  reg  M_48_offset;  // ufix1
  wire M_48_1;  // ufix1
  reg  M_49_offset;  // ufix1
  wire M_49_1;  // ufix1
  reg  M_50_offset;  // ufix1
  wire M_50_1;  // ufix1
  reg  M_51_offset;  // ufix1
  wire M_51_1;  // ufix1
  reg  M_52_offset;  // ufix1
  wire M_52_1;  // ufix1
  reg  M_53_offset;  // ufix1
  wire M_53_1;  // ufix1
  reg  M_54_offset;  // ufix1
  wire M_54_1;  // ufix1
  reg  M_55_offset;  // ufix1
  wire M_55_1;  // ufix1
  reg  M_56_offset;  // ufix1
  wire M_56_1;  // ufix1
  reg  M_57_offset;  // ufix1
  wire M_57_1;  // ufix1
  reg  M_58_offset;  // ufix1
  wire M_58_1;  // ufix1
  reg  M_59_offset;  // ufix1
  wire M_59_1;  // ufix1
  reg  M_60_offset;  // ufix1
  wire M_60_1;  // ufix1
  reg  M_61_offset;  // ufix1
  wire M_61_1;  // ufix1
  reg  M_62_offset;  // ufix1
  wire M_62_1;  // ufix1
  reg  M_63_offset;  // ufix1
  wire M_63_1;  // ufix1
  reg  N_0_offset;  // ufix1
  wire N_0_1;  // ufix1
  reg  N_1_offset;  // ufix1
  wire N_1_1;  // ufix1
  reg  N_2_offset;  // ufix1
  wire N_2_1;  // ufix1
  reg  N_3_offset;  // ufix1
  wire N_3_1;  // ufix1
  reg  N_4_offset;  // ufix1
  wire N_4_1;  // ufix1
  reg  N_5_offset;  // ufix1
  wire N_5_1;  // ufix1
  reg  N_6_offset;  // ufix1
  wire N_6_1;  // ufix1
  reg [13:0] W_0_offset;  // ufix14_En13
  wire [13:0] W_0_1;  // ufix14_En13
  reg [13:0] W_1_offset;  // ufix14_En13
  wire [13:0] W_1_1;  // ufix14_En13
  reg [13:0] W_2_offset;  // ufix14_En13
  wire [13:0] W_2_1;  // ufix14_En13
  reg [13:0] W_3_offset;  // ufix14_En13
  wire [13:0] W_3_1;  // ufix14_En13
  reg [13:0] W_4_offset;  // ufix14_En13
  wire [13:0] W_4_1;  // ufix14_En13
  reg [13:0] W_5_offset;  // ufix14_En13
  wire [13:0] W_5_1;  // ufix14_En13
  reg [13:0] W_6_offset;  // ufix14_En13
  wire [13:0] W_6_1;  // ufix14_En13
  reg [6:0] Tm_offset;  // ufix7
  wire [6:0] Tm_1;  // ufix7
  reg [2:0] Tn_offset;  // ufix3
  wire [2:0] Tn_1;  // ufix3
  wire [13:0] M_out_0;  // ufix14_En12
  wire [13:0] M_out_1;  // ufix14_En12
  wire [13:0] M_out_2;  // ufix14_En12
  wire [13:0] M_out_3;  // ufix14_En12
  wire [13:0] M_out_4;  // ufix14_En12
  wire [13:0] M_out_5;  // ufix14_En12
  wire [13:0] M_out_6;  // ufix14_En12
  wire [13:0] M_out_7;  // ufix14_En12
  wire [13:0] M_out_8;  // ufix14_En12
  wire [13:0] M_out_9;  // ufix14_En12
  wire [13:0] M_out_10;  // ufix14_En12
  wire [13:0] M_out_11;  // ufix14_En12
  wire [13:0] M_out_12;  // ufix14_En12
  wire [13:0] M_out_13;  // ufix14_En12
  wire [13:0] M_out_14;  // ufix14_En12
  wire [13:0] M_out_15;  // ufix14_En12
  wire [13:0] M_out_16;  // ufix14_En12
  wire [13:0] M_out_17;  // ufix14_En12
  wire [13:0] M_out_18;  // ufix14_En12
  wire [13:0] M_out_19;  // ufix14_En12
  wire [13:0] M_out_20;  // ufix14_En12
  wire [13:0] M_out_21;  // ufix14_En12
  wire [13:0] M_out_22;  // ufix14_En12
  wire [13:0] M_out_23;  // ufix14_En12
  wire [13:0] M_out_24;  // ufix14_En12
  wire [13:0] M_out_25;  // ufix14_En12
  wire [13:0] M_out_26;  // ufix14_En12
  wire [13:0] M_out_27;  // ufix14_En12
  wire [13:0] M_out_28;  // ufix14_En12
  wire [13:0] M_out_29;  // ufix14_En12
  wire [13:0] M_out_30;  // ufix14_En12
  wire [13:0] M_out_31;  // ufix14_En12
  wire [13:0] M_out_32;  // ufix14_En12
  wire [13:0] M_out_33;  // ufix14_En12
  wire [13:0] M_out_34;  // ufix14_En12
  wire [13:0] M_out_35;  // ufix14_En12
  wire [13:0] M_out_36;  // ufix14_En12
  wire [13:0] M_out_37;  // ufix14_En12
  wire [13:0] M_out_38;  // ufix14_En12
  wire [13:0] M_out_39;  // ufix14_En12
  wire [13:0] M_out_40;  // ufix14_En12
  wire [13:0] M_out_41;  // ufix14_En12
  wire [13:0] M_out_42;  // ufix14_En12
  wire [13:0] M_out_43;  // ufix14_En12
  wire [13:0] M_out_44;  // ufix14_En12
  wire [13:0] M_out_45;  // ufix14_En12
  wire [13:0] M_out_46;  // ufix14_En12
  wire [13:0] M_out_47;  // ufix14_En12
  wire [13:0] M_out_48;  // ufix14_En12
  wire [13:0] M_out_49;  // ufix14_En12
  wire [13:0] M_out_50;  // ufix14_En12
  wire [13:0] M_out_51;  // ufix14_En12
  wire [13:0] M_out_52;  // ufix14_En12
  wire [13:0] M_out_53;  // ufix14_En12
  wire [13:0] M_out_54;  // ufix14_En12
  wire [13:0] M_out_55;  // ufix14_En12
  wire [13:0] M_out_56;  // ufix14_En12
  wire [13:0] M_out_57;  // ufix14_En12
  wire [13:0] M_out_58;  // ufix14_En12
  wire [13:0] M_out_59;  // ufix14_En12
  wire [13:0] M_out_60;  // ufix14_En12
  wire [13:0] M_out_61;  // ufix14_En12
  wire [13:0] M_out_62;  // ufix14_En12
  wire [13:0] M_out_63;  // ufix14_En12
  wire [13:0] M_out_0_0_expected_1;  // ufix14_En12
  wire [13:0] M_out_0_ref;  // ufix14_En12
  reg  M_out_0_testFailure;  // ufix1
  wire [13:0] M_out_0_1_expected_1;  // ufix14_En12
  wire [13:0] M_out_1_ref;  // ufix14_En12
  reg  M_out_1_testFailure;  // ufix1
  wire [13:0] M_out_0_2_expected_1;  // ufix14_En12
  wire [13:0] M_out_2_ref;  // ufix14_En12
  reg  M_out_2_testFailure;  // ufix1
  wire [13:0] M_out_0_3_expected_1;  // ufix14_En12
  wire [13:0] M_out_3_ref;  // ufix14_En12
  reg  M_out_3_testFailure;  // ufix1
  wire [13:0] M_out_0_4_expected_1;  // ufix14_En12
  wire [13:0] M_out_4_ref;  // ufix14_En12
  reg  M_out_4_testFailure;  // ufix1
  wire [13:0] M_out_0_5_expected_1;  // ufix14_En12
  wire [13:0] M_out_5_ref;  // ufix14_En12
  reg  M_out_5_testFailure;  // ufix1
  wire [13:0] M_out_0_6_expected_1;  // ufix14_En12
  wire [13:0] M_out_6_ref;  // ufix14_En12
  reg  M_out_6_testFailure;  // ufix1
  wire [13:0] M_out_0_7_expected_1;  // ufix14_En12
  wire [13:0] M_out_7_ref;  // ufix14_En12
  reg  M_out_7_testFailure;  // ufix1
  wire [13:0] M_out_0_8_expected_1;  // ufix14_En12
  wire [13:0] M_out_8_ref;  // ufix14_En12
  reg  M_out_8_testFailure;  // ufix1
  wire [13:0] M_out_0_9_expected_1;  // ufix14_En12
  wire [13:0] M_out_9_ref;  // ufix14_En12
  reg  M_out_9_testFailure;  // ufix1
  wire [13:0] M_out_0_10_expected_1;  // ufix14_En12
  wire [13:0] M_out_10_ref;  // ufix14_En12
  reg  M_out_10_testFailure;  // ufix1
  wire [13:0] M_out_0_11_expected_1;  // ufix14_En12
  wire [13:0] M_out_11_ref;  // ufix14_En12
  reg  M_out_11_testFailure;  // ufix1
  wire [13:0] M_out_0_12_expected_1;  // ufix14_En12
  wire [13:0] M_out_12_ref;  // ufix14_En12
  reg  M_out_12_testFailure;  // ufix1
  wire [13:0] M_out_0_13_expected_1;  // ufix14_En12
  wire [13:0] M_out_13_ref;  // ufix14_En12
  reg  M_out_13_testFailure;  // ufix1
  wire [13:0] M_out_0_14_expected_1;  // ufix14_En12
  wire [13:0] M_out_14_ref;  // ufix14_En12
  reg  M_out_14_testFailure;  // ufix1
  wire [13:0] M_out_0_15_expected_1;  // ufix14_En12
  wire [13:0] M_out_15_ref;  // ufix14_En12
  reg  M_out_15_testFailure;  // ufix1
  wire [13:0] M_out_0_16_expected_1;  // ufix14_En12
  wire [13:0] M_out_16_ref;  // ufix14_En12
  reg  M_out_16_testFailure;  // ufix1
  wire [13:0] M_out_0_17_expected_1;  // ufix14_En12
  wire [13:0] M_out_17_ref;  // ufix14_En12
  reg  M_out_17_testFailure;  // ufix1
  wire [13:0] M_out_0_18_expected_1;  // ufix14_En12
  wire [13:0] M_out_18_ref;  // ufix14_En12
  reg  M_out_18_testFailure;  // ufix1
  wire [13:0] M_out_0_19_expected_1;  // ufix14_En12
  wire [13:0] M_out_19_ref;  // ufix14_En12
  reg  M_out_19_testFailure;  // ufix1
  wire [13:0] M_out_0_20_expected_1;  // ufix14_En12
  wire [13:0] M_out_20_ref;  // ufix14_En12
  reg  M_out_20_testFailure;  // ufix1
  wire [13:0] M_out_0_21_expected_1;  // ufix14_En12
  wire [13:0] M_out_21_ref;  // ufix14_En12
  reg  M_out_21_testFailure;  // ufix1
  wire [13:0] M_out_0_22_expected_1;  // ufix14_En12
  wire [13:0] M_out_22_ref;  // ufix14_En12
  reg  M_out_22_testFailure;  // ufix1
  wire [13:0] M_out_0_23_expected_1;  // ufix14_En12
  wire [13:0] M_out_23_ref;  // ufix14_En12
  reg  M_out_23_testFailure;  // ufix1
  wire [13:0] M_out_0_24_expected_1;  // ufix14_En12
  wire [13:0] M_out_24_ref;  // ufix14_En12
  reg  M_out_24_testFailure;  // ufix1
  wire [13:0] M_out_0_25_expected_1;  // ufix14_En12
  wire [13:0] M_out_25_ref;  // ufix14_En12
  reg  M_out_25_testFailure;  // ufix1
  wire [13:0] M_out_0_26_expected_1;  // ufix14_En12
  wire [13:0] M_out_26_ref;  // ufix14_En12
  reg  M_out_26_testFailure;  // ufix1
  wire [13:0] M_out_0_27_expected_1;  // ufix14_En12
  wire [13:0] M_out_27_ref;  // ufix14_En12
  reg  M_out_27_testFailure;  // ufix1
  wire [13:0] M_out_0_28_expected_1;  // ufix14_En12
  wire [13:0] M_out_28_ref;  // ufix14_En12
  reg  M_out_28_testFailure;  // ufix1
  wire [13:0] M_out_0_29_expected_1;  // ufix14_En12
  wire [13:0] M_out_29_ref;  // ufix14_En12
  reg  M_out_29_testFailure;  // ufix1
  wire [13:0] M_out_0_30_expected_1;  // ufix14_En12
  wire [13:0] M_out_30_ref;  // ufix14_En12
  reg  M_out_30_testFailure;  // ufix1
  wire [13:0] M_out_0_31_expected_1;  // ufix14_En12
  wire [13:0] M_out_31_ref;  // ufix14_En12
  reg  M_out_31_testFailure;  // ufix1
  wire [13:0] M_out_0_32_expected_1;  // ufix14_En12
  wire [13:0] M_out_32_ref;  // ufix14_En12
  reg  M_out_32_testFailure;  // ufix1
  wire [13:0] M_out_0_33_expected_1;  // ufix14_En12
  wire [13:0] M_out_33_ref;  // ufix14_En12
  reg  M_out_33_testFailure;  // ufix1
  wire [13:0] M_out_0_34_expected_1;  // ufix14_En12
  wire [13:0] M_out_34_ref;  // ufix14_En12
  reg  M_out_34_testFailure;  // ufix1
  wire [13:0] M_out_0_35_expected_1;  // ufix14_En12
  wire [13:0] M_out_35_ref;  // ufix14_En12
  reg  M_out_35_testFailure;  // ufix1
  wire [13:0] M_out_0_36_expected_1;  // ufix14_En12
  wire [13:0] M_out_36_ref;  // ufix14_En12
  reg  M_out_36_testFailure;  // ufix1
  wire [13:0] M_out_0_37_expected_1;  // ufix14_En12
  wire [13:0] M_out_37_ref;  // ufix14_En12
  reg  M_out_37_testFailure;  // ufix1
  wire [13:0] M_out_0_38_expected_1;  // ufix14_En12
  wire [13:0] M_out_38_ref;  // ufix14_En12
  reg  M_out_38_testFailure;  // ufix1
  wire [13:0] M_out_0_39_expected_1;  // ufix14_En12
  wire [13:0] M_out_39_ref;  // ufix14_En12
  reg  M_out_39_testFailure;  // ufix1
  wire [13:0] M_out_0_40_expected_1;  // ufix14_En12
  wire [13:0] M_out_40_ref;  // ufix14_En12
  reg  M_out_40_testFailure;  // ufix1
  wire [13:0] M_out_0_41_expected_1;  // ufix14_En12
  wire [13:0] M_out_41_ref;  // ufix14_En12
  reg  M_out_41_testFailure;  // ufix1
  wire [13:0] M_out_0_42_expected_1;  // ufix14_En12
  wire [13:0] M_out_42_ref;  // ufix14_En12
  reg  M_out_42_testFailure;  // ufix1
  wire [13:0] M_out_0_43_expected_1;  // ufix14_En12
  wire [13:0] M_out_43_ref;  // ufix14_En12
  reg  M_out_43_testFailure;  // ufix1
  wire [13:0] M_out_0_44_expected_1;  // ufix14_En12
  wire [13:0] M_out_44_ref;  // ufix14_En12
  reg  M_out_44_testFailure;  // ufix1
  wire [13:0] M_out_0_45_expected_1;  // ufix14_En12
  wire [13:0] M_out_45_ref;  // ufix14_En12
  reg  M_out_45_testFailure;  // ufix1
  wire [13:0] M_out_0_46_expected_1;  // ufix14_En12
  wire [13:0] M_out_46_ref;  // ufix14_En12
  reg  M_out_46_testFailure;  // ufix1
  wire [13:0] M_out_0_47_expected_1;  // ufix14_En12
  wire [13:0] M_out_47_ref;  // ufix14_En12
  reg  M_out_47_testFailure;  // ufix1
  wire [13:0] M_out_0_48_expected_1;  // ufix14_En12
  wire [13:0] M_out_48_ref;  // ufix14_En12
  reg  M_out_48_testFailure;  // ufix1
  wire [13:0] M_out_0_49_expected_1;  // ufix14_En12
  wire [13:0] M_out_49_ref;  // ufix14_En12
  reg  M_out_49_testFailure;  // ufix1
  wire [13:0] M_out_0_50_expected_1;  // ufix14_En12
  wire [13:0] M_out_50_ref;  // ufix14_En12
  reg  M_out_50_testFailure;  // ufix1
  wire [13:0] M_out_0_51_expected_1;  // ufix14_En12
  wire [13:0] M_out_51_ref;  // ufix14_En12
  reg  M_out_51_testFailure;  // ufix1
  wire [13:0] M_out_0_52_expected_1;  // ufix14_En12
  wire [13:0] M_out_52_ref;  // ufix14_En12
  reg  M_out_52_testFailure;  // ufix1
  wire [13:0] M_out_0_53_expected_1;  // ufix14_En12
  wire [13:0] M_out_53_ref;  // ufix14_En12
  reg  M_out_53_testFailure;  // ufix1
  wire [13:0] M_out_0_54_expected_1;  // ufix14_En12
  wire [13:0] M_out_54_ref;  // ufix14_En12
  reg  M_out_54_testFailure;  // ufix1
  wire [13:0] M_out_0_55_expected_1;  // ufix14_En12
  wire [13:0] M_out_55_ref;  // ufix14_En12
  reg  M_out_55_testFailure;  // ufix1
  wire [13:0] M_out_0_56_expected_1;  // ufix14_En12
  wire [13:0] M_out_56_ref;  // ufix14_En12
  reg  M_out_56_testFailure;  // ufix1
  wire [13:0] M_out_0_57_expected_1;  // ufix14_En12
  wire [13:0] M_out_57_ref;  // ufix14_En12
  reg  M_out_57_testFailure;  // ufix1
  wire [13:0] M_out_0_58_expected_1;  // ufix14_En12
  wire [13:0] M_out_58_ref;  // ufix14_En12
  reg  M_out_58_testFailure;  // ufix1
  wire [13:0] M_out_0_59_expected_1;  // ufix14_En12
  wire [13:0] M_out_59_ref;  // ufix14_En12
  reg  M_out_59_testFailure;  // ufix1
  wire [13:0] M_out_0_60_expected_1;  // ufix14_En12
  wire [13:0] M_out_60_ref;  // ufix14_En12
  reg  M_out_60_testFailure;  // ufix1
  wire [13:0] M_out_0_61_expected_1;  // ufix14_En12
  wire [13:0] M_out_61_ref;  // ufix14_En12
  reg  M_out_61_testFailure;  // ufix1
  wire [13:0] M_out_0_62_expected_1;  // ufix14_En12
  wire [13:0] M_out_62_ref;  // ufix14_En12
  reg  M_out_62_testFailure;  // ufix1
  wire [13:0] M_out_0_63_expected_1;  // ufix14_En12
  wire [13:0] M_out_63_ref;  // ufix14_En12
  reg  M_out_63_testFailure;  // ufix1
  reg  testFailure;  // ufix1
  reg  or_t;  // ufix1
  assign M_out_0_lastAddr = 1'b1;
  assign snkDonen =  ~ check1_done;
  assign tb_enb = resetn & snkDonen;
  assign rdEnb = (check1_done == 1'b0 ? tb_enb :
              1'b0);
  assign M_out_0_done_enb = M_out_0_done & rdEnb;
  always
    begin : clk_gen
      clk <= 1'b1;
      # (5);
      clk <= 1'b0;
      # (5);
      if (check1_done == 1'b1) begin
        clk <= 1'b1;
        # (5);
        clk <= 1'b0;
        # (5);
        $stop;
      end
    end
  initial
    begin : reset_gen
      reset <= 1'b1;
      # (20);
      @ (posedge clk)
      # (2);
      reset <= 1'b0;
    end
  assign resetn =  ~ reset;
  assign M_out_0_done = M_out_0_lastAddr & resetn;
  // Delay to allow last sim cycle to complete
  always @(posedge clk or posedge reset)
    begin : checkDone_1
      if (reset) begin
        check1_done <= 0;
      end
      else begin
        if (M_out_0_done_enb) begin
          check1_done <= M_out_0_done;
        end
      end
    end
  assign #2 enb = rdEnb;
  assign ce_out = enb & (rdEnb & tb_enb);
  // Data source for M_0
  assign rawData_M_0 = 1'b0;
  // holdData reg for M
  always @(posedge clk or posedge reset)
    begin : stimuli_M
      if (reset) begin
        holdData_M_0 <= 1'bx;
      end
      else begin
        holdData_M_0 <= rawData_M_0;
      end
    end
  // Data source for M_1
  assign rawData_M_1 = 1'b0;
  // holdData reg for M
  always @(posedge clk or posedge reset)
    begin : stimuli_M_1
      if (reset) begin
        holdData_M_1 <= 1'bx;
      end
      else begin
        holdData_M_1 <= rawData_M_1;
      end
    end
  // Data source for M_2
  assign rawData_M_2 = 1'b0;
  // holdData reg for M
  always @(posedge clk or posedge reset)
    begin : stimuli_M_2
      if (reset) begin
        holdData_M_2 <= 1'bx;
      end
      else begin
        holdData_M_2 <= rawData_M_2;
      end
    end
  // Data source for M_3
  assign rawData_M_3 = 1'b0;
  // holdData reg for M
  always @(posedge clk or posedge reset)
    begin : stimuli_M_3
      if (reset) begin
        holdData_M_3 <= 1'bx;
      end
      else begin
        holdData_M_3 <= rawData_M_3;
      end
    end
  // Data source for M_4
  assign rawData_M_4 = 1'b0;
  // holdData reg for M
  always @(posedge clk or posedge reset)
    begin : stimuli_M_4
      if (reset) begin
        holdData_M_4 <= 1'bx;
      end
      else begin
        holdData_M_4 <= rawData_M_4;
      end
    end
  // Data source for M_5
  assign rawData_M_5 = 1'b0;
  // holdData reg for M
  always @(posedge clk or posedge reset)
    begin : stimuli_M_5
      if (reset) begin
        holdData_M_5 <= 1'bx;
      end
      else begin
        holdData_M_5 <= rawData_M_5;
      end
    end
  // Data source for M_6
  assign rawData_M_6 = 1'b0;
  // holdData reg for M
  always @(posedge clk or posedge reset)
    begin : stimuli_M_6
      if (reset) begin
        holdData_M_6 <= 1'bx;
      end
      else begin
        holdData_M_6 <= rawData_M_6;
      end
    end
  // Data source for M_7
  assign rawData_M_7 = 1'b0;
  // holdData reg for M
  always @(posedge clk or posedge reset)
    begin : stimuli_M_7
      if (reset) begin
        holdData_M_7 <= 1'bx;
      end
      else begin
        holdData_M_7 <= rawData_M_7;
      end
    end
  // Data source for M_8
  assign rawData_M_8 = 1'b0;
  // holdData reg for M
  always @(posedge clk or posedge reset)
    begin : stimuli_M_8
      if (reset) begin
        holdData_M_8 <= 1'bx;
      end
      else begin
        holdData_M_8 <= rawData_M_8;
      end
    end
  // Data source for M_9
  assign rawData_M_9 = 1'b0;
  // holdData reg for M
  always @(posedge clk or posedge reset)
    begin : stimuli_M_9
      if (reset) begin
        holdData_M_9 <= 1'bx;
      end
      else begin
        holdData_M_9 <= rawData_M_9;
      end
    end
  // Data source for M_10
  assign rawData_M_10 = 1'b0;
  // holdData reg for M
  always @(posedge clk or posedge reset)
    begin : stimuli_M_10
      if (reset) begin
        holdData_M_10 <= 1'bx;
      end
      else begin
        holdData_M_10 <= rawData_M_10;
      end
    end
  // Data source for M_11
  assign rawData_M_11 = 1'b0;
  // holdData reg for M
  always @(posedge clk or posedge reset)
    begin : stimuli_M_11
      if (reset) begin
        holdData_M_11 <= 1'bx;
      end
      else begin
        holdData_M_11 <= rawData_M_11;
      end
    end
  // Data source for M_12
  assign rawData_M_12 = 1'b0;
  // holdData reg for M
  always @(posedge clk or posedge reset)
    begin : stimuli_M_12
      if (reset) begin
        holdData_M_12 <= 1'bx;
      end
      else begin
        holdData_M_12 <= rawData_M_12;
      end
    end
  // Data source for M_13
  assign rawData_M_13 = 1'b0;
  // holdData reg for M
  always @(posedge clk or posedge reset)
    begin : stimuli_M_13
      if (reset) begin
        holdData_M_13 <= 1'bx;
      end
      else begin
        holdData_M_13 <= rawData_M_13;
      end
    end
  // Data source for M_14
  assign rawData_M_14 = 1'b0;
  // holdData reg for M
  always @(posedge clk or posedge reset)
    begin : stimuli_M_14
      if (reset) begin
        holdData_M_14 <= 1'bx;
      end
      else begin
        holdData_M_14 <= rawData_M_14;
      end
    end
  // Data source for M_15
  assign rawData_M_15 = 1'b0;
  // holdData reg for M
  always @(posedge clk or posedge reset)
    begin : stimuli_M_15
      if (reset) begin
        holdData_M_15 <= 1'bx;
      end
      else begin
        holdData_M_15 <= rawData_M_15;
      end
    end
  // Data source for M_16
  assign rawData_M_16 = 1'b0;
  // holdData reg for M
  always @(posedge clk or posedge reset)
    begin : stimuli_M_16
      if (reset) begin
        holdData_M_16 <= 1'bx;
      end
      else begin
        holdData_M_16 <= rawData_M_16;
      end
    end
  // Data source for M_17
  assign rawData_M_17 = 1'b0;
  // holdData reg for M
  always @(posedge clk or posedge reset)
    begin : stimuli_M_17
      if (reset) begin
        holdData_M_17 <= 1'bx;
      end
      else begin
        holdData_M_17 <= rawData_M_17;
      end
    end
  // Data source for M_18
  assign rawData_M_18 = 1'b0;
  // holdData reg for M
  always @(posedge clk or posedge reset)
    begin : stimuli_M_18
      if (reset) begin
        holdData_M_18 <= 1'bx;
      end
      else begin
        holdData_M_18 <= rawData_M_18;
      end
    end
  // Data source for M_19
  assign rawData_M_19 = 1'b0;
  // holdData reg for M
  always @(posedge clk or posedge reset)
    begin : stimuli_M_19
      if (reset) begin
        holdData_M_19 <= 1'bx;
      end
      else begin
        holdData_M_19 <= rawData_M_19;
      end
    end
  // Data source for M_20
  assign rawData_M_20 = 1'b0;
  // holdData reg for M
  always @(posedge clk or posedge reset)
    begin : stimuli_M_20
      if (reset) begin
        holdData_M_20 <= 1'bx;
      end
      else begin
        holdData_M_20 <= rawData_M_20;
      end
    end
  // Data source for M_21
  assign rawData_M_21 = 1'b0;
  // holdData reg for M
  always @(posedge clk or posedge reset)
    begin : stimuli_M_21
      if (reset) begin
        holdData_M_21 <= 1'bx;
      end
      else begin
        holdData_M_21 <= rawData_M_21;
      end
    end
  // Data source for M_22
  assign rawData_M_22 = 1'b0;
  // holdData reg for M
  always @(posedge clk or posedge reset)
    begin : stimuli_M_22
      if (reset) begin
        holdData_M_22 <= 1'bx;
      end
      else begin
        holdData_M_22 <= rawData_M_22;
      end
    end
  // Data source for M_23
  assign rawData_M_23 = 1'b0;
  // holdData reg for M
  always @(posedge clk or posedge reset)
    begin : stimuli_M_23
      if (reset) begin
        holdData_M_23 <= 1'bx;
      end
      else begin
        holdData_M_23 <= rawData_M_23;
      end
    end
  // Data source for M_24
  assign rawData_M_24 = 1'b0;
  // holdData reg for M
  always @(posedge clk or posedge reset)
    begin : stimuli_M_24
      if (reset) begin
        holdData_M_24 <= 1'bx;
      end
      else begin
        holdData_M_24 <= rawData_M_24;
      end
    end
  // Data source for M_25
  assign rawData_M_25 = 1'b0;
  // holdData reg for M
  always @(posedge clk or posedge reset)
    begin : stimuli_M_25
      if (reset) begin
        holdData_M_25 <= 1'bx;
      end
      else begin
        holdData_M_25 <= rawData_M_25;
      end
    end
  // Data source for M_26
  assign rawData_M_26 = 1'b0;
  // holdData reg for M
  always @(posedge clk or posedge reset)
    begin : stimuli_M_26
      if (reset) begin
        holdData_M_26 <= 1'bx;
      end
      else begin
        holdData_M_26 <= rawData_M_26;
      end
    end
  // Data source for M_27
  assign rawData_M_27 = 1'b0;
  // holdData reg for M
  always @(posedge clk or posedge reset)
    begin : stimuli_M_27
      if (reset) begin
        holdData_M_27 <= 1'bx;
      end
      else begin
        holdData_M_27 <= rawData_M_27;
      end
    end
  // Data source for M_28
  assign rawData_M_28 = 1'b0;
  // holdData reg for M
  always @(posedge clk or posedge reset)
    begin : stimuli_M_28
      if (reset) begin
        holdData_M_28 <= 1'bx;
      end
      else begin
        holdData_M_28 <= rawData_M_28;
      end
    end
  // Data source for M_29
  assign rawData_M_29 = 1'b0;
  // holdData reg for M
  always @(posedge clk or posedge reset)
    begin : stimuli_M_29
      if (reset) begin
        holdData_M_29 <= 1'bx;
      end
      else begin
        holdData_M_29 <= rawData_M_29;
      end
    end
  // Data source for M_30
  assign rawData_M_30 = 1'b0;
  // holdData reg for M
  always @(posedge clk or posedge reset)
    begin : stimuli_M_30
      if (reset) begin
        holdData_M_30 <= 1'bx;
      end
      else begin
        holdData_M_30 <= rawData_M_30;
      end
    end
  // Data source for M_31
  assign rawData_M_31 = 1'b0;
  // holdData reg for M
  always @(posedge clk or posedge reset)
    begin : stimuli_M_31
      if (reset) begin
        holdData_M_31 <= 1'bx;
      end
      else begin
        holdData_M_31 <= rawData_M_31;
      end
    end
  // Data source for M_32
  assign rawData_M_32 = 1'b0;
  // holdData reg for M
  always @(posedge clk or posedge reset)
    begin : stimuli_M_32
      if (reset) begin
        holdData_M_32 <= 1'bx;
      end
      else begin
        holdData_M_32 <= rawData_M_32;
      end
    end
  // Data source for M_33
  assign rawData_M_33 = 1'b0;
  // holdData reg for M
  always @(posedge clk or posedge reset)
    begin : stimuli_M_33
      if (reset) begin
        holdData_M_33 <= 1'bx;
      end
      else begin
        holdData_M_33 <= rawData_M_33;
      end
    end
  // Data source for M_34
  assign rawData_M_34 = 1'b0;
  // holdData reg for M
  always @(posedge clk or posedge reset)
    begin : stimuli_M_34
      if (reset) begin
        holdData_M_34 <= 1'bx;
      end
      else begin
        holdData_M_34 <= rawData_M_34;
      end
    end
  // Data source for M_35
  assign rawData_M_35 = 1'b0;
  // holdData reg for M
  always @(posedge clk or posedge reset)
    begin : stimuli_M_35
      if (reset) begin
        holdData_M_35 <= 1'bx;
      end
      else begin
        holdData_M_35 <= rawData_M_35;
      end
    end
  // Data source for M_36
  assign rawData_M_36 = 1'b0;
  // holdData reg for M
  always @(posedge clk or posedge reset)
    begin : stimuli_M_36
      if (reset) begin
        holdData_M_36 <= 1'bx;
      end
      else begin
        holdData_M_36 <= rawData_M_36;
      end
    end
  // Data source for M_37
  assign rawData_M_37 = 1'b0;
  // holdData reg for M
  always @(posedge clk or posedge reset)
    begin : stimuli_M_37
      if (reset) begin
        holdData_M_37 <= 1'bx;
      end
      else begin
        holdData_M_37 <= rawData_M_37;
      end
    end
  // Data source for M_38
  assign rawData_M_38 = 1'b0;
  // holdData reg for M
  always @(posedge clk or posedge reset)
    begin : stimuli_M_38
      if (reset) begin
        holdData_M_38 <= 1'bx;
      end
      else begin
        holdData_M_38 <= rawData_M_38;
      end
    end
  // Data source for M_39
  assign rawData_M_39 = 1'b0;
  // holdData reg for M
  always @(posedge clk or posedge reset)
    begin : stimuli_M_39
      if (reset) begin
        holdData_M_39 <= 1'bx;
      end
      else begin
        holdData_M_39 <= rawData_M_39;
      end
    end
  // Data source for M_40
  assign rawData_M_40 = 1'b0;
  // holdData reg for M
  always @(posedge clk or posedge reset)
    begin : stimuli_M_40
      if (reset) begin
        holdData_M_40 <= 1'bx;
      end
      else begin
        holdData_M_40 <= rawData_M_40;
      end
    end
  // Data source for M_41
  assign rawData_M_41 = 1'b0;
  // holdData reg for M
  always @(posedge clk or posedge reset)
    begin : stimuli_M_41
      if (reset) begin
        holdData_M_41 <= 1'bx;
      end
      else begin
        holdData_M_41 <= rawData_M_41;
      end
    end
  // Data source for M_42
  assign rawData_M_42 = 1'b0;
  // holdData reg for M
  always @(posedge clk or posedge reset)
    begin : stimuli_M_42
      if (reset) begin
        holdData_M_42 <= 1'bx;
      end
      else begin
        holdData_M_42 <= rawData_M_42;
      end
    end
  // Data source for M_43
  assign rawData_M_43 = 1'b0;
  // holdData reg for M
  always @(posedge clk or posedge reset)
    begin : stimuli_M_43
      if (reset) begin
        holdData_M_43 <= 1'bx;
      end
      else begin
        holdData_M_43 <= rawData_M_43;
      end
    end
  // Data source for M_44
  assign rawData_M_44 = 1'b0;
  // holdData reg for M
  always @(posedge clk or posedge reset)
    begin : stimuli_M_44
      if (reset) begin
        holdData_M_44 <= 1'bx;
      end
      else begin
        holdData_M_44 <= rawData_M_44;
      end
    end
  // Data source for M_45
  assign rawData_M_45 = 1'b0;
  // holdData reg for M
  always @(posedge clk or posedge reset)
    begin : stimuli_M_45
      if (reset) begin
        holdData_M_45 <= 1'bx;
      end
      else begin
        holdData_M_45 <= rawData_M_45;
      end
    end
  // Data source for M_46
  assign rawData_M_46 = 1'b0;
  // holdData reg for M
  always @(posedge clk or posedge reset)
    begin : stimuli_M_46
      if (reset) begin
        holdData_M_46 <= 1'bx;
      end
      else begin
        holdData_M_46 <= rawData_M_46;
      end
    end
  // Data source for M_47
  assign rawData_M_47 = 1'b0;
  // holdData reg for M
  always @(posedge clk or posedge reset)
    begin : stimuli_M_47
      if (reset) begin
        holdData_M_47 <= 1'bx;
      end
      else begin
        holdData_M_47 <= rawData_M_47;
      end
    end
  // Data source for M_48
  assign rawData_M_48 = 1'b0;
  // holdData reg for M
  always @(posedge clk or posedge reset)
    begin : stimuli_M_48
      if (reset) begin
        holdData_M_48 <= 1'bx;
      end
      else begin
        holdData_M_48 <= rawData_M_48;
      end
    end
  // Data source for M_49
  assign rawData_M_49 = 1'b0;
  // holdData reg for M
  always @(posedge clk or posedge reset)
    begin : stimuli_M_49
      if (reset) begin
        holdData_M_49 <= 1'bx;
      end
      else begin
        holdData_M_49 <= rawData_M_49;
      end
    end
  // Data source for M_50
  assign rawData_M_50 = 1'b0;
  // holdData reg for M
  always @(posedge clk or posedge reset)
    begin : stimuli_M_50
      if (reset) begin
        holdData_M_50 <= 1'bx;
      end
      else begin
        holdData_M_50 <= rawData_M_50;
      end
    end
  // Data source for M_51
  assign rawData_M_51 = 1'b0;
  // holdData reg for M
  always @(posedge clk or posedge reset)
    begin : stimuli_M_51
      if (reset) begin
        holdData_M_51 <= 1'bx;
      end
      else begin
        holdData_M_51 <= rawData_M_51;
      end
    end
  // Data source for M_52
  assign rawData_M_52 = 1'b0;
  // holdData reg for M
  always @(posedge clk or posedge reset)
    begin : stimuli_M_52
      if (reset) begin
        holdData_M_52 <= 1'bx;
      end
      else begin
        holdData_M_52 <= rawData_M_52;
      end
    end
  // Data source for M_53
  assign rawData_M_53 = 1'b0;
  // holdData reg for M
  always @(posedge clk or posedge reset)
    begin : stimuli_M_53
      if (reset) begin
        holdData_M_53 <= 1'bx;
      end
      else begin
        holdData_M_53 <= rawData_M_53;
      end
    end
  // Data source for M_54
  assign rawData_M_54 = 1'b0;
  // holdData reg for M
  always @(posedge clk or posedge reset)
    begin : stimuli_M_54
      if (reset) begin
        holdData_M_54 <= 1'bx;
      end
      else begin
        holdData_M_54 <= rawData_M_54;
      end
    end
  // Data source for M_55
  assign rawData_M_55 = 1'b0;
  // holdData reg for M
  always @(posedge clk or posedge reset)
    begin : stimuli_M_55
      if (reset) begin
        holdData_M_55 <= 1'bx;
      end
      else begin
        holdData_M_55 <= rawData_M_55;
      end
    end
  // Data source for M_56
  assign rawData_M_56 = 1'b0;
  // holdData reg for M
  always @(posedge clk or posedge reset)
    begin : stimuli_M_56
      if (reset) begin
        holdData_M_56 <= 1'bx;
      end
      else begin
        holdData_M_56 <= rawData_M_56;
      end
    end
  // Data source for M_57
  assign rawData_M_57 = 1'b0;
  // holdData reg for M
  always @(posedge clk or posedge reset)
    begin : stimuli_M_57
      if (reset) begin
        holdData_M_57 <= 1'bx;
      end
      else begin
        holdData_M_57 <= rawData_M_57;
      end
    end
  // Data source for M_58
  assign rawData_M_58 = 1'b0;
  // holdData reg for M
  always @(posedge clk or posedge reset)
    begin : stimuli_M_58
      if (reset) begin
        holdData_M_58 <= 1'bx;
      end
      else begin
        holdData_M_58 <= rawData_M_58;
      end
    end
  // Data source for M_59
  assign rawData_M_59 = 1'b0;
  // holdData reg for M
  always @(posedge clk or posedge reset)
    begin : stimuli_M_59
      if (reset) begin
        holdData_M_59 <= 1'bx;
      end
      else begin
        holdData_M_59 <= rawData_M_59;
      end
    end
  // Data source for M_60
  assign rawData_M_60 = 1'b0;
  // holdData reg for M
  always @(posedge clk or posedge reset)
    begin : stimuli_M_60
      if (reset) begin
        holdData_M_60 <= 1'bx;
      end
      else begin
        holdData_M_60 <= rawData_M_60;
      end
    end
  // Data source for M_61
  assign rawData_M_61 = 1'b0;
  // holdData reg for M
  always @(posedge clk or posedge reset)
    begin : stimuli_M_61
      if (reset) begin
        holdData_M_61 <= 1'bx;
      end
      else begin
        holdData_M_61 <= rawData_M_61;
      end
    end
  // Data source for M_62
  assign rawData_M_62 = 1'b0;
  // holdData reg for M
  always @(posedge clk or posedge reset)
    begin : stimuli_M_62
      if (reset) begin
        holdData_M_62 <= 1'bx;
      end
      else begin
        holdData_M_62 <= rawData_M_62;
      end
    end
  // Data source for M_63
  assign rawData_M_63 = 1'b0;
  // holdData reg for M
  always @(posedge clk or posedge reset)
    begin : stimuli_M_63
      if (reset) begin
        holdData_M_63 <= 1'bx;
      end
      else begin
        holdData_M_63 <= rawData_M_63;
      end
    end
  // Data source for N_0
  assign rawData_N_0 = 1'b1;
  // holdData reg for N
  always @(posedge clk or posedge reset)
    begin : stimuli_N
      if (reset) begin
        holdData_N_0 <= 1'bx;
      end
      else begin
        holdData_N_0 <= rawData_N_0;
      end
    end
  // Data source for N_1
  assign rawData_N_1 = 1'b1;
  // holdData reg for N
  always @(posedge clk or posedge reset)
    begin : stimuli_N_1
      if (reset) begin
        holdData_N_1 <= 1'bx;
      end
      else begin
        holdData_N_1 <= rawData_N_1;
      end
    end
  // Data source for N_2
  assign rawData_N_2 = 1'b1;
  // holdData reg for N
  always @(posedge clk or posedge reset)
    begin : stimuli_N_2
      if (reset) begin
        holdData_N_2 <= 1'bx;
      end
      else begin
        holdData_N_2 <= rawData_N_2;
      end
    end
  // Data source for N_3
  assign rawData_N_3 = 1'b1;
  // holdData reg for N
  always @(posedge clk or posedge reset)
    begin : stimuli_N_3
      if (reset) begin
        holdData_N_3 <= 1'bx;
      end
      else begin
        holdData_N_3 <= rawData_N_3;
      end
    end
  // Data source for N_4
  assign rawData_N_4 = 1'b1;
  // holdData reg for N
  always @(posedge clk or posedge reset)
    begin : stimuli_N_4
      if (reset) begin
        holdData_N_4 <= 1'bx;
      end
      else begin
        holdData_N_4 <= rawData_N_4;
      end
    end
  // Data source for N_5
  assign rawData_N_5 = 1'b1;
  // holdData reg for N
  always @(posedge clk or posedge reset)
    begin : stimuli_N_5
      if (reset) begin
        holdData_N_5 <= 1'bx;
      end
      else begin
        holdData_N_5 <= rawData_N_5;
      end
    end
  // Data source for N_6
  assign rawData_N_6 = 1'b1;
  // holdData reg for N
  always @(posedge clk or posedge reset)
    begin : stimuli_N_6
      if (reset) begin
        holdData_N_6 <= 1'bx;
      end
      else begin
        holdData_N_6 <= rawData_N_6;
      end
    end
  // Data source for W_0
  assign rawData_W_0 = 14'b10000000000000;
  // holdData reg for W
  always @(posedge clk or posedge reset)
    begin : stimuli_W
      if (reset) begin
        holdData_W_0 <= 14'bx;
      end
      else begin
        holdData_W_0 <= rawData_W_0;
      end
    end
  // Data source for W_1
  assign rawData_W_1 = 14'b01111001100110;
  // holdData reg for W
  always @(posedge clk or posedge reset)
    begin : stimuli_W_1
      if (reset) begin
        holdData_W_1 <= 14'bx;
      end
      else begin
        holdData_W_1 <= rawData_W_1;
      end
    end
  // Data source for W_2
  assign rawData_W_2 = 14'b01101100110011;
  // holdData reg for W
  always @(posedge clk or posedge reset)
    begin : stimuli_W_2
      if (reset) begin
        holdData_W_2 <= 14'bx;
      end
      else begin
        holdData_W_2 <= rawData_W_2;
      end
    end
  // Data source for W_3
  assign rawData_W_3 = 14'b00100000000000;
  // holdData reg for W
  always @(posedge clk or posedge reset)
    begin : stimuli_W_3
      if (reset) begin
        holdData_W_3 <= 14'bx;
      end
      else begin
        holdData_W_3 <= rawData_W_3;
      end
    end
  // Data source for W_4
  assign rawData_W_4 = 14'b00000000000000;
  // holdData reg for W
  always @(posedge clk or posedge reset)
    begin : stimuli_W_4
      if (reset) begin
        holdData_W_4 <= 14'bx;
      end
      else begin
        holdData_W_4 <= rawData_W_4;
      end
    end
  // Data source for W_5
  assign rawData_W_5 = 14'b00000000000000;
  // holdData reg for W
  always @(posedge clk or posedge reset)
    begin : stimuli_W_5
      if (reset) begin
        holdData_W_5 <= 14'bx;
      end
      else begin
        holdData_W_5 <= rawData_W_5;
      end
    end
  // Data source for W_6
  assign rawData_W_6 = 14'b00111001100110;
  // holdData reg for W
  always @(posedge clk or posedge reset)
    begin : stimuli_W_6
      if (reset) begin
        holdData_W_6 <= 14'bx;
      end
      else begin
        holdData_W_6 <= rawData_W_6;
      end
    end
  // Data source for Tm
  assign rawData_Tm = 7'b1000000;
  // holdData reg for Tm
  always @(posedge clk or posedge reset)
    begin : stimuli_Tm
      if (reset) begin
        holdData_Tm <= 7'bx;
      end
      else begin
        holdData_Tm <= rawData_Tm;
      end
    end
  // Data source for Tn
  assign rawData_Tn = 3'b111;
  // holdData reg for Tn
  always @(posedge clk or posedge reset)
    begin : stimuli_Tn
      if (reset) begin
        holdData_Tn <= 3'bx;
      end
      else begin
        holdData_Tn <= rawData_Tn;
      end
    end
  always @(rawData_M_0 or rdEnb)
    begin : stimuli_M_64
      if (rdEnb == 1'b0) begin
        M_0_offset <= holdData_M_0;
      end
      else begin
        M_0_offset <= rawData_M_0;
      end
    end
  assign #2 M_0_1 = M_0_offset;
  always @(rawData_M_1 or rdEnb)
    begin : stimuli_M_65
      if (rdEnb == 1'b0) begin
        M_1_offset <= holdData_M_1;
      end
      else begin
        M_1_offset <= rawData_M_1;
      end
    end
  assign #2 M_1_1 = M_1_offset;
  always @(rawData_M_2 or rdEnb)
    begin : stimuli_M_66
      if (rdEnb == 1'b0) begin
        M_2_offset <= holdData_M_2;
      end
      else begin
        M_2_offset <= rawData_M_2;
      end
    end
  assign #2 M_2_1 = M_2_offset;
  always @(rawData_M_3 or rdEnb)
    begin : stimuli_M_67
      if (rdEnb == 1'b0) begin
        M_3_offset <= holdData_M_3;
      end
      else begin
        M_3_offset <= rawData_M_3;
      end
    end
  assign #2 M_3_1 = M_3_offset;
  always @(rawData_M_4 or rdEnb)
    begin : stimuli_M_68
      if (rdEnb == 1'b0) begin
        M_4_offset <= holdData_M_4;
      end
      else begin
        M_4_offset <= rawData_M_4;
      end
    end
  assign #2 M_4_1 = M_4_offset;
  always @(rawData_M_5 or rdEnb)
    begin : stimuli_M_69
      if (rdEnb == 1'b0) begin
        M_5_offset <= holdData_M_5;
      end
      else begin
        M_5_offset <= rawData_M_5;
      end
    end
  assign #2 M_5_1 = M_5_offset;
  always @(rawData_M_6 or rdEnb)
    begin : stimuli_M_70
      if (rdEnb == 1'b0) begin
        M_6_offset <= holdData_M_6;
      end
      else begin
        M_6_offset <= rawData_M_6;
      end
    end
  assign #2 M_6_1 = M_6_offset;
  always @(rawData_M_7 or rdEnb)
    begin : stimuli_M_71
      if (rdEnb == 1'b0) begin
        M_7_offset <= holdData_M_7;
      end
      else begin
        M_7_offset <= rawData_M_7;
      end
    end
  assign #2 M_7_1 = M_7_offset;
  always @(rawData_M_8 or rdEnb)
    begin : stimuli_M_72
      if (rdEnb == 1'b0) begin
        M_8_offset <= holdData_M_8;
      end
      else begin
        M_8_offset <= rawData_M_8;
      end
    end
  assign #2 M_8_1 = M_8_offset;
  always @(rawData_M_9 or rdEnb)
    begin : stimuli_M_73
      if (rdEnb == 1'b0) begin
        M_9_offset <= holdData_M_9;
      end
      else begin
        M_9_offset <= rawData_M_9;
      end
    end
  assign #2 M_9_1 = M_9_offset;
  always @(rawData_M_10 or rdEnb)
    begin : stimuli_M_74
      if (rdEnb == 1'b0) begin
        M_10_offset <= holdData_M_10;
      end
      else begin
        M_10_offset <= rawData_M_10;
      end
    end
  assign #2 M_10_1 = M_10_offset;
  always @(rawData_M_11 or rdEnb)
    begin : stimuli_M_75
      if (rdEnb == 1'b0) begin
        M_11_offset <= holdData_M_11;
      end
      else begin
        M_11_offset <= rawData_M_11;
      end
    end
  assign #2 M_11_1 = M_11_offset;
  always @(rawData_M_12 or rdEnb)
    begin : stimuli_M_76
      if (rdEnb == 1'b0) begin
        M_12_offset <= holdData_M_12;
      end
      else begin
        M_12_offset <= rawData_M_12;
      end
    end
  assign #2 M_12_1 = M_12_offset;
  always @(rawData_M_13 or rdEnb)
    begin : stimuli_M_77
      if (rdEnb == 1'b0) begin
        M_13_offset <= holdData_M_13;
      end
      else begin
        M_13_offset <= rawData_M_13;
      end
    end
  assign #2 M_13_1 = M_13_offset;
  always @(rawData_M_14 or rdEnb)
    begin : stimuli_M_78
      if (rdEnb == 1'b0) begin
        M_14_offset <= holdData_M_14;
      end
      else begin
        M_14_offset <= rawData_M_14;
      end
    end
  assign #2 M_14_1 = M_14_offset;
  always @(rawData_M_15 or rdEnb)
    begin : stimuli_M_79
      if (rdEnb == 1'b0) begin
        M_15_offset <= holdData_M_15;
      end
      else begin
        M_15_offset <= rawData_M_15;
      end
    end
  assign #2 M_15_1 = M_15_offset;
  always @(rawData_M_16 or rdEnb)
    begin : stimuli_M_80
      if (rdEnb == 1'b0) begin
        M_16_offset <= holdData_M_16;
      end
      else begin
        M_16_offset <= rawData_M_16;
      end
    end
  assign #2 M_16_1 = M_16_offset;
  always @(rawData_M_17 or rdEnb)
    begin : stimuli_M_81
      if (rdEnb == 1'b0) begin
        M_17_offset <= holdData_M_17;
      end
      else begin
        M_17_offset <= rawData_M_17;
      end
    end
  assign #2 M_17_1 = M_17_offset;
  always @(rawData_M_18 or rdEnb)
    begin : stimuli_M_82
      if (rdEnb == 1'b0) begin
        M_18_offset <= holdData_M_18;
      end
      else begin
        M_18_offset <= rawData_M_18;
      end
    end
  assign #2 M_18_1 = M_18_offset;
  always @(rawData_M_19 or rdEnb)
    begin : stimuli_M_83
      if (rdEnb == 1'b0) begin
        M_19_offset <= holdData_M_19;
      end
      else begin
        M_19_offset <= rawData_M_19;
      end
    end
  assign #2 M_19_1 = M_19_offset;
  always @(rawData_M_20 or rdEnb)
    begin : stimuli_M_84
      if (rdEnb == 1'b0) begin
        M_20_offset <= holdData_M_20;
      end
      else begin
        M_20_offset <= rawData_M_20;
      end
    end
  assign #2 M_20_1 = M_20_offset;
  always @(rawData_M_21 or rdEnb)
    begin : stimuli_M_85
      if (rdEnb == 1'b0) begin
        M_21_offset <= holdData_M_21;
      end
      else begin
        M_21_offset <= rawData_M_21;
      end
    end
  assign #2 M_21_1 = M_21_offset;
  always @(rawData_M_22 or rdEnb)
    begin : stimuli_M_86
      if (rdEnb == 1'b0) begin
        M_22_offset <= holdData_M_22;
      end
      else begin
        M_22_offset <= rawData_M_22;
      end
    end
  assign #2 M_22_1 = M_22_offset;
  always @(rawData_M_23 or rdEnb)
    begin : stimuli_M_87
      if (rdEnb == 1'b0) begin
        M_23_offset <= holdData_M_23;
      end
      else begin
        M_23_offset <= rawData_M_23;
      end
    end
  assign #2 M_23_1 = M_23_offset;
  always @(rawData_M_24 or rdEnb)
    begin : stimuli_M_88
      if (rdEnb == 1'b0) begin
        M_24_offset <= holdData_M_24;
      end
      else begin
        M_24_offset <= rawData_M_24;
      end
    end
  assign #2 M_24_1 = M_24_offset;
  always @(rawData_M_25 or rdEnb)
    begin : stimuli_M_89
      if (rdEnb == 1'b0) begin
        M_25_offset <= holdData_M_25;
      end
      else begin
        M_25_offset <= rawData_M_25;
      end
    end
  assign #2 M_25_1 = M_25_offset;
  always @(rawData_M_26 or rdEnb)
    begin : stimuli_M_90
      if (rdEnb == 1'b0) begin
        M_26_offset <= holdData_M_26;
      end
      else begin
        M_26_offset <= rawData_M_26;
      end
    end
  assign #2 M_26_1 = M_26_offset;
  always @(rawData_M_27 or rdEnb)
    begin : stimuli_M_91
      if (rdEnb == 1'b0) begin
        M_27_offset <= holdData_M_27;
      end
      else begin
        M_27_offset <= rawData_M_27;
      end
    end
  assign #2 M_27_1 = M_27_offset;
  always @(rawData_M_28 or rdEnb)
    begin : stimuli_M_92
      if (rdEnb == 1'b0) begin
        M_28_offset <= holdData_M_28;
      end
      else begin
        M_28_offset <= rawData_M_28;
      end
    end
  assign #2 M_28_1 = M_28_offset;
  always @(rawData_M_29 or rdEnb)
    begin : stimuli_M_93
      if (rdEnb == 1'b0) begin
        M_29_offset <= holdData_M_29;
      end
      else begin
        M_29_offset <= rawData_M_29;
      end
    end
  assign #2 M_29_1 = M_29_offset;
  always @(rawData_M_30 or rdEnb)
    begin : stimuli_M_94
      if (rdEnb == 1'b0) begin
        M_30_offset <= holdData_M_30;
      end
      else begin
        M_30_offset <= rawData_M_30;
      end
    end
  assign #2 M_30_1 = M_30_offset;
  always @(rawData_M_31 or rdEnb)
    begin : stimuli_M_95
      if (rdEnb == 1'b0) begin
        M_31_offset <= holdData_M_31;
      end
      else begin
        M_31_offset <= rawData_M_31;
      end
    end
  assign #2 M_31_1 = M_31_offset;
  always @(rawData_M_32 or rdEnb)
    begin : stimuli_M_96
      if (rdEnb == 1'b0) begin
        M_32_offset <= holdData_M_32;
      end
      else begin
        M_32_offset <= rawData_M_32;
      end
    end
  assign #2 M_32_1 = M_32_offset;
  always @(rawData_M_33 or rdEnb)
    begin : stimuli_M_97
      if (rdEnb == 1'b0) begin
        M_33_offset <= holdData_M_33;
      end
      else begin
        M_33_offset <= rawData_M_33;
      end
    end
  assign #2 M_33_1 = M_33_offset;
  always @(rawData_M_34 or rdEnb)
    begin : stimuli_M_98
      if (rdEnb == 1'b0) begin
        M_34_offset <= holdData_M_34;
      end
      else begin
        M_34_offset <= rawData_M_34;
      end
    end
  assign #2 M_34_1 = M_34_offset;
  always @(rawData_M_35 or rdEnb)
    begin : stimuli_M_99
      if (rdEnb == 1'b0) begin
        M_35_offset <= holdData_M_35;
      end
      else begin
        M_35_offset <= rawData_M_35;
      end
    end
  assign #2 M_35_1 = M_35_offset;
  always @(rawData_M_36 or rdEnb)
    begin : stimuli_M_100
      if (rdEnb == 1'b0) begin
        M_36_offset <= holdData_M_36;
      end
      else begin
        M_36_offset <= rawData_M_36;
      end
    end
  assign #2 M_36_1 = M_36_offset;
  always @(rawData_M_37 or rdEnb)
    begin : stimuli_M_101
      if (rdEnb == 1'b0) begin
        M_37_offset <= holdData_M_37;
      end
      else begin
        M_37_offset <= rawData_M_37;
      end
    end
  assign #2 M_37_1 = M_37_offset;
  always @(rawData_M_38 or rdEnb)
    begin : stimuli_M_102
      if (rdEnb == 1'b0) begin
        M_38_offset <= holdData_M_38;
      end
      else begin
        M_38_offset <= rawData_M_38;
      end
    end
  assign #2 M_38_1 = M_38_offset;
  always @(rawData_M_39 or rdEnb)
    begin : stimuli_M_103
      if (rdEnb == 1'b0) begin
        M_39_offset <= holdData_M_39;
      end
      else begin
        M_39_offset <= rawData_M_39;
      end
    end
  assign #2 M_39_1 = M_39_offset;
  always @(rawData_M_40 or rdEnb)
    begin : stimuli_M_104
      if (rdEnb == 1'b0) begin
        M_40_offset <= holdData_M_40;
      end
      else begin
        M_40_offset <= rawData_M_40;
      end
    end
  assign #2 M_40_1 = M_40_offset;
  always @(rawData_M_41 or rdEnb)
    begin : stimuli_M_105
      if (rdEnb == 1'b0) begin
        M_41_offset <= holdData_M_41;
      end
      else begin
        M_41_offset <= rawData_M_41;
      end
    end
  assign #2 M_41_1 = M_41_offset;
  always @(rawData_M_42 or rdEnb)
    begin : stimuli_M_106
      if (rdEnb == 1'b0) begin
        M_42_offset <= holdData_M_42;
      end
      else begin
        M_42_offset <= rawData_M_42;
      end
    end
  assign #2 M_42_1 = M_42_offset;
  always @(rawData_M_43 or rdEnb)
    begin : stimuli_M_107
      if (rdEnb == 1'b0) begin
        M_43_offset <= holdData_M_43;
      end
      else begin
        M_43_offset <= rawData_M_43;
      end
    end
  assign #2 M_43_1 = M_43_offset;
  always @(rawData_M_44 or rdEnb)
    begin : stimuli_M_108
      if (rdEnb == 1'b0) begin
        M_44_offset <= holdData_M_44;
      end
      else begin
        M_44_offset <= rawData_M_44;
      end
    end
  assign #2 M_44_1 = M_44_offset;
  always @(rawData_M_45 or rdEnb)
    begin : stimuli_M_109
      if (rdEnb == 1'b0) begin
        M_45_offset <= holdData_M_45;
      end
      else begin
        M_45_offset <= rawData_M_45;
      end
    end
  assign #2 M_45_1 = M_45_offset;
  always @(rawData_M_46 or rdEnb)
    begin : stimuli_M_110
      if (rdEnb == 1'b0) begin
        M_46_offset <= holdData_M_46;
      end
      else begin
        M_46_offset <= rawData_M_46;
      end
    end
  assign #2 M_46_1 = M_46_offset;
  always @(rawData_M_47 or rdEnb)
    begin : stimuli_M_111
      if (rdEnb == 1'b0) begin
        M_47_offset <= holdData_M_47;
      end
      else begin
        M_47_offset <= rawData_M_47;
      end
    end
  assign #2 M_47_1 = M_47_offset;
  always @(rawData_M_48 or rdEnb)
    begin : stimuli_M_112
      if (rdEnb == 1'b0) begin
        M_48_offset <= holdData_M_48;
      end
      else begin
        M_48_offset <= rawData_M_48;
      end
    end
  assign #2 M_48_1 = M_48_offset;
  always @(rawData_M_49 or rdEnb)
    begin : stimuli_M_113
      if (rdEnb == 1'b0) begin
        M_49_offset <= holdData_M_49;
      end
      else begin
        M_49_offset <= rawData_M_49;
      end
    end
  assign #2 M_49_1 = M_49_offset;
  always @(rawData_M_50 or rdEnb)
    begin : stimuli_M_114
      if (rdEnb == 1'b0) begin
        M_50_offset <= holdData_M_50;
      end
      else begin
        M_50_offset <= rawData_M_50;
      end
    end
  assign #2 M_50_1 = M_50_offset;
  always @(rawData_M_51 or rdEnb)
    begin : stimuli_M_115
      if (rdEnb == 1'b0) begin
        M_51_offset <= holdData_M_51;
      end
      else begin
        M_51_offset <= rawData_M_51;
      end
    end
  assign #2 M_51_1 = M_51_offset;
  always @(rawData_M_52 or rdEnb)
    begin : stimuli_M_116
      if (rdEnb == 1'b0) begin
        M_52_offset <= holdData_M_52;
      end
      else begin
        M_52_offset <= rawData_M_52;
      end
    end
  assign #2 M_52_1 = M_52_offset;
  always @(rawData_M_53 or rdEnb)
    begin : stimuli_M_117
      if (rdEnb == 1'b0) begin
        M_53_offset <= holdData_M_53;
      end
      else begin
        M_53_offset <= rawData_M_53;
      end
    end
  assign #2 M_53_1 = M_53_offset;
  always @(rawData_M_54 or rdEnb)
    begin : stimuli_M_118
      if (rdEnb == 1'b0) begin
        M_54_offset <= holdData_M_54;
      end
      else begin
        M_54_offset <= rawData_M_54;
      end
    end
  assign #2 M_54_1 = M_54_offset;
  always @(rawData_M_55 or rdEnb)
    begin : stimuli_M_119
      if (rdEnb == 1'b0) begin
        M_55_offset <= holdData_M_55;
      end
      else begin
        M_55_offset <= rawData_M_55;
      end
    end
  assign #2 M_55_1 = M_55_offset;
  always @(rawData_M_56 or rdEnb)
    begin : stimuli_M_120
      if (rdEnb == 1'b0) begin
        M_56_offset <= holdData_M_56;
      end
      else begin
        M_56_offset <= rawData_M_56;
      end
    end
  assign #2 M_56_1 = M_56_offset;
  always @(rawData_M_57 or rdEnb)
    begin : stimuli_M_121
      if (rdEnb == 1'b0) begin
        M_57_offset <= holdData_M_57;
      end
      else begin
        M_57_offset <= rawData_M_57;
      end
    end
  assign #2 M_57_1 = M_57_offset;
  always @(rawData_M_58 or rdEnb)
    begin : stimuli_M_122
      if (rdEnb == 1'b0) begin
        M_58_offset <= holdData_M_58;
      end
      else begin
        M_58_offset <= rawData_M_58;
      end
    end
  assign #2 M_58_1 = M_58_offset;
  always @(rawData_M_59 or rdEnb)
    begin : stimuli_M_123
      if (rdEnb == 1'b0) begin
        M_59_offset <= holdData_M_59;
      end
      else begin
        M_59_offset <= rawData_M_59;
      end
    end
  assign #2 M_59_1 = M_59_offset;
  always @(rawData_M_60 or rdEnb)
    begin : stimuli_M_124
      if (rdEnb == 1'b0) begin
        M_60_offset <= holdData_M_60;
      end
      else begin
        M_60_offset <= rawData_M_60;
      end
    end
  assign #2 M_60_1 = M_60_offset;
  always @(rawData_M_61 or rdEnb)
    begin : stimuli_M_125
      if (rdEnb == 1'b0) begin
        M_61_offset <= holdData_M_61;
      end
      else begin
        M_61_offset <= rawData_M_61;
      end
    end
  assign #2 M_61_1 = M_61_offset;
  always @(rawData_M_62 or rdEnb)
    begin : stimuli_M_126
      if (rdEnb == 1'b0) begin
        M_62_offset <= holdData_M_62;
      end
      else begin
        M_62_offset <= rawData_M_62;
      end
    end
  assign #2 M_62_1 = M_62_offset;
  always @(rawData_M_63 or rdEnb)
    begin : stimuli_M_127
      if (rdEnb == 1'b0) begin
        M_63_offset <= holdData_M_63;
      end
      else begin
        M_63_offset <= rawData_M_63;
      end
    end
  assign #2 M_63_1 = M_63_offset;
  always @(rawData_N_0 or rdEnb)
    begin : stimuli_N_7
      if (rdEnb == 1'b0) begin
        N_0_offset <= holdData_N_0;
      end
      else begin
        N_0_offset <= rawData_N_0;
      end
    end
  assign #2 N_0_1 = N_0_offset;
  always @(rawData_N_1 or rdEnb)
    begin : stimuli_N_8
      if (rdEnb == 1'b0) begin
        N_1_offset <= holdData_N_1;
      end
      else begin
        N_1_offset <= rawData_N_1;
      end
    end
  assign #2 N_1_1 = N_1_offset;
  always @(rawData_N_2 or rdEnb)
    begin : stimuli_N_9
      if (rdEnb == 1'b0) begin
        N_2_offset <= holdData_N_2;
      end
      else begin
        N_2_offset <= rawData_N_2;
      end
    end
  assign #2 N_2_1 = N_2_offset;
  always @(rawData_N_3 or rdEnb)
    begin : stimuli_N_10
      if (rdEnb == 1'b0) begin
        N_3_offset <= holdData_N_3;
      end
      else begin
        N_3_offset <= rawData_N_3;
      end
    end
  assign #2 N_3_1 = N_3_offset;
  always @(rawData_N_4 or rdEnb)
    begin : stimuli_N_11
      if (rdEnb == 1'b0) begin
        N_4_offset <= holdData_N_4;
      end
      else begin
        N_4_offset <= rawData_N_4;
      end
    end
  assign #2 N_4_1 = N_4_offset;
  always @(rawData_N_5 or rdEnb)
    begin : stimuli_N_12
      if (rdEnb == 1'b0) begin
        N_5_offset <= holdData_N_5;
      end
      else begin
        N_5_offset <= rawData_N_5;
      end
    end
  assign #2 N_5_1 = N_5_offset;
  always @(rawData_N_6 or rdEnb)
    begin : stimuli_N_13
      if (rdEnb == 1'b0) begin
        N_6_offset <= holdData_N_6;
      end
      else begin
        N_6_offset <= rawData_N_6;
      end
    end
  assign #2 N_6_1 = N_6_offset;
  always @(rawData_W_0 or rdEnb)
    begin : stimuli_W_7
      if (rdEnb == 1'b0) begin
        W_0_offset <= holdData_W_0;
      end
      else begin
        W_0_offset <= rawData_W_0;
      end
    end
  assign #2 W_0_1 = W_0_offset;
  always @(rawData_W_1 or rdEnb)
    begin : stimuli_W_8
      if (rdEnb == 1'b0) begin
        W_1_offset <= holdData_W_1;
      end
      else begin
        W_1_offset <= rawData_W_1;
      end
    end
  assign #2 W_1_1 = W_1_offset;
  always @(rawData_W_2 or rdEnb)
    begin : stimuli_W_9
      if (rdEnb == 1'b0) begin
        W_2_offset <= holdData_W_2;
      end
      else begin
        W_2_offset <= rawData_W_2;
      end
    end
  assign #2 W_2_1 = W_2_offset;
  always @(rawData_W_3 or rdEnb)
    begin : stimuli_W_10
      if (rdEnb == 1'b0) begin
        W_3_offset <= holdData_W_3;
      end
      else begin
        W_3_offset <= rawData_W_3;
      end
    end
  assign #2 W_3_1 = W_3_offset;
  always @(rawData_W_4 or rdEnb)
    begin : stimuli_W_11
      if (rdEnb == 1'b0) begin
        W_4_offset <= holdData_W_4;
      end
      else begin
        W_4_offset <= rawData_W_4;
      end
    end
  assign #2 W_4_1 = W_4_offset;
  always @(rawData_W_5 or rdEnb)
    begin : stimuli_W_12
      if (rdEnb == 1'b0) begin
        W_5_offset <= holdData_W_5;
      end
      else begin
        W_5_offset <= rawData_W_5;
      end
    end
  assign #2 W_5_1 = W_5_offset;
  always @(rawData_W_6 or rdEnb)
    begin : stimuli_W_13
      if (rdEnb == 1'b0) begin
        W_6_offset <= holdData_W_6;
      end
      else begin
        W_6_offset <= rawData_W_6;
      end
    end
  assign #2 W_6_1 = W_6_offset;
  always @(rawData_Tm or rdEnb)
    begin : stimuli_Tm_1
      if (rdEnb == 1'b0) begin
        Tm_offset <= holdData_Tm;
      end
      else begin
        Tm_offset <= rawData_Tm;
      end
    end
  assign #2 Tm_1 = Tm_offset;
  always @(rawData_Tn or rdEnb)
    begin : stimuli_Tn_1
      if (rdEnb == 1'b0) begin
        Tn_offset <= holdData_Tn;
      end
      else begin
        Tn_offset <= rawData_Tn;
      end
    end
  assign #2 Tn_1 = Tn_offset;
  mac_fixpt   u_mac_fixpt   (.M_0(M_0_1),  // ufix1
                             .M_1(M_1_1),  // ufix1
                             .M_2(M_2_1),  // ufix1
                             .M_3(M_3_1),  // ufix1
                             .M_4(M_4_1),  // ufix1
                             .M_5(M_5_1),  // ufix1
                             .M_6(M_6_1),  // ufix1
                             .M_7(M_7_1),  // ufix1
                             .M_8(M_8_1),  // ufix1
                             .M_9(M_9_1),  // ufix1
                             .M_10(M_10_1),  // ufix1
                             .M_11(M_11_1),  // ufix1
                             .M_12(M_12_1),  // ufix1
                             .M_13(M_13_1),  // ufix1
                             .M_14(M_14_1),  // ufix1
                             .M_15(M_15_1),  // ufix1
                             .M_16(M_16_1),  // ufix1
                             .M_17(M_17_1),  // ufix1
                             .M_18(M_18_1),  // ufix1
                             .M_19(M_19_1),  // ufix1
                             .M_20(M_20_1),  // ufix1
                             .M_21(M_21_1),  // ufix1
                             .M_22(M_22_1),  // ufix1
                             .M_23(M_23_1),  // ufix1
                             .M_24(M_24_1),  // ufix1
                             .M_25(M_25_1),  // ufix1
                             .M_26(M_26_1),  // ufix1
                             .M_27(M_27_1),  // ufix1
                             .M_28(M_28_1),  // ufix1
                             .M_29(M_29_1),  // ufix1
                             .M_30(M_30_1),  // ufix1
                             .M_31(M_31_1),  // ufix1
                             .M_32(M_32_1),  // ufix1
                             .M_33(M_33_1),  // ufix1
                             .M_34(M_34_1),  // ufix1
                             .M_35(M_35_1),  // ufix1
                             .M_36(M_36_1),  // ufix1
                             .M_37(M_37_1),  // ufix1
                             .M_38(M_38_1),  // ufix1
                             .M_39(M_39_1),  // ufix1
                             .M_40(M_40_1),  // ufix1
                             .M_41(M_41_1),  // ufix1
                             .M_42(M_42_1),  // ufix1
                             .M_43(M_43_1),  // ufix1
                             .M_44(M_44_1),  // ufix1
                             .M_45(M_45_1),  // ufix1
                             .M_46(M_46_1),  // ufix1
                             .M_47(M_47_1),  // ufix1
                             .M_48(M_48_1),  // ufix1
                             .M_49(M_49_1),  // ufix1
                             .M_50(M_50_1),  // ufix1
                             .M_51(M_51_1),  // ufix1
                             .M_52(M_52_1),  // ufix1
                             .M_53(M_53_1),  // ufix1
                             .M_54(M_54_1),  // ufix1
                             .M_55(M_55_1),  // ufix1
                             .M_56(M_56_1),  // ufix1
                             .M_57(M_57_1),  // ufix1
                             .M_58(M_58_1),  // ufix1
                             .M_59(M_59_1),  // ufix1
                             .M_60(M_60_1),  // ufix1
                             .M_61(M_61_1),  // ufix1
                             .M_62(M_62_1),  // ufix1
                             .M_63(M_63_1),  // ufix1
                             .N_0(N_0_1),  // ufix1
                             .N_1(N_1_1),  // ufix1
                             .N_2(N_2_1),  // ufix1
                             .N_3(N_3_1),  // ufix1
                             .N_4(N_4_1),  // ufix1
                             .N_5(N_5_1),  // ufix1
                             .N_6(N_6_1),  // ufix1
                             .W_0(W_0_1),  // ufix14_En13
                             .W_1(W_1_1),  // ufix14_En13
                             .W_2(W_2_1),  // ufix14_En13
                             .W_3(W_3_1),  // ufix14_En13
                             .W_4(W_4_1),  // ufix14_En13
                             .W_5(W_5_1),  // ufix14_En13
                             .W_6(W_6_1),  // ufix14_En13
                             .Tm(Tm_1),  // ufix7
                             .Tn(Tn_1),  // ufix3
                             .M_out_0(M_out_0),  // ufix14_En12
                             .M_out_1(M_out_1),  // ufix14_En12
                             .M_out_2(M_out_2),  // ufix14_En12
                             .M_out_3(M_out_3),  // ufix14_En12
                             .M_out_4(M_out_4),  // ufix14_En12
                             .M_out_5(M_out_5),  // ufix14_En12
                             .M_out_6(M_out_6),  // ufix14_En12
                             .M_out_7(M_out_7),  // ufix14_En12
                             .M_out_8(M_out_8),  // ufix14_En12
                             .M_out_9(M_out_9),  // ufix14_En12
                             .M_out_10(M_out_10),  // ufix14_En12
                             .M_out_11(M_out_11),  // ufix14_En12
                             .M_out_12(M_out_12),  // ufix14_En12
                             .M_out_13(M_out_13),  // ufix14_En12
                             .M_out_14(M_out_14),  // ufix14_En12
                             .M_out_15(M_out_15),  // ufix14_En12
                             .M_out_16(M_out_16),  // ufix14_En12
                             .M_out_17(M_out_17),  // ufix14_En12
                             .M_out_18(M_out_18),  // ufix14_En12
                             .M_out_19(M_out_19),  // ufix14_En12
                             .M_out_20(M_out_20),  // ufix14_En12
                             .M_out_21(M_out_21),  // ufix14_En12
                             .M_out_22(M_out_22),  // ufix14_En12
                             .M_out_23(M_out_23),  // ufix14_En12
                             .M_out_24(M_out_24),  // ufix14_En12
                             .M_out_25(M_out_25),  // ufix14_En12
                             .M_out_26(M_out_26),  // ufix14_En12
                             .M_out_27(M_out_27),  // ufix14_En12
                             .M_out_28(M_out_28),  // ufix14_En12
                             .M_out_29(M_out_29),  // ufix14_En12
                             .M_out_30(M_out_30),  // ufix14_En12
                             .M_out_31(M_out_31),  // ufix14_En12
                             .M_out_32(M_out_32),  // ufix14_En12
                             .M_out_33(M_out_33),  // ufix14_En12
                             .M_out_34(M_out_34),  // ufix14_En12
                             .M_out_35(M_out_35),  // ufix14_En12
                             .M_out_36(M_out_36),  // ufix14_En12
                             .M_out_37(M_out_37),  // ufix14_En12
                             .M_out_38(M_out_38),  // ufix14_En12
                             .M_out_39(M_out_39),  // ufix14_En12
                             .M_out_40(M_out_40),  // ufix14_En12
                             .M_out_41(M_out_41),  // ufix14_En12
                             .M_out_42(M_out_42),  // ufix14_En12
                             .M_out_43(M_out_43),  // ufix14_En12
                             .M_out_44(M_out_44),  // ufix14_En12
                             .M_out_45(M_out_45),  // ufix14_En12
                             .M_out_46(M_out_46),  // ufix14_En12
                             .M_out_47(M_out_47),  // ufix14_En12
                             .M_out_48(M_out_48),  // ufix14_En12
                             .M_out_49(M_out_49),  // ufix14_En12
                             .M_out_50(M_out_50),  // ufix14_En12
                             .M_out_51(M_out_51),  // ufix14_En12
                             .M_out_52(M_out_52),  // ufix14_En12
                             .M_out_53(M_out_53),  // ufix14_En12
                             .M_out_54(M_out_54),  // ufix14_En12
                             .M_out_55(M_out_55),  // ufix14_En12
                             .M_out_56(M_out_56),  // ufix14_En12
                             .M_out_57(M_out_57),  // ufix14_En12
                             .M_out_58(M_out_58),  // ufix14_En12
                             .M_out_59(M_out_59),  // ufix14_En12
                             .M_out_60(M_out_60),  // ufix14_En12
                             .M_out_61(M_out_61),  // ufix14_En12
                             .M_out_62(M_out_62),  // ufix14_En12
                             .M_out_63(M_out_63)  // ufix14_En12
                             );
  // Data source for M_out_0_0_expected
  assign M_out_0_0_expected_1 = 14'b11011111111111;
  assign M_out_0_ref = M_out_0_0_expected_1;
  always @(posedge clk or posedge reset)
    begin : M_out_0_checker
      if (reset == 1'b1) begin
        M_out_0_testFailure <= 1'b0;
      end
      else begin
        if (ce_out == 1'b1 && M_out_0 !== M_out_0_ref) begin
          M_out_0_testFailure <= 1'b1;
          $display("ERROR in M_out_0 at time %t : Expected '%h' Actual '%h'", $time, M_out_0_ref, M_out_0);
        end
      end
    end
  // Data source for M_out_0_1_expected
  assign M_out_0_1_expected_1 = 14'b11011111111111;
  assign M_out_1_ref = M_out_0_1_expected_1;
  always @(posedge clk or posedge reset)
    begin : M_out_1_checker
      if (reset == 1'b1) begin
        M_out_1_testFailure <= 1'b0;
      end
      else begin
        if (ce_out == 1'b1 && M_out_1 !== M_out_1_ref) begin
          M_out_1_testFailure <= 1'b1;
          $display("ERROR in M_out_1 at time %t : Expected '%h' Actual '%h'", $time, M_out_1_ref, M_out_1);
        end
      end
    end
  // Data source for M_out_0_2_expected
  assign M_out_0_2_expected_1 = 14'b11011111111111;
  assign M_out_2_ref = M_out_0_2_expected_1;
  always @(posedge clk or posedge reset)
    begin : M_out_2_checker
      if (reset == 1'b1) begin
        M_out_2_testFailure <= 1'b0;
      end
      else begin
        if (ce_out == 1'b1 && M_out_2 !== M_out_2_ref) begin
          M_out_2_testFailure <= 1'b1;
          $display("ERROR in M_out_2 at time %t : Expected '%h' Actual '%h'", $time, M_out_2_ref, M_out_2);
        end
      end
    end
  // Data source for M_out_0_3_expected
  assign M_out_0_3_expected_1 = 14'b11011111111111;
  assign M_out_3_ref = M_out_0_3_expected_1;
  always @(posedge clk or posedge reset)
    begin : M_out_3_checker
      if (reset == 1'b1) begin
        M_out_3_testFailure <= 1'b0;
      end
      else begin
        if (ce_out == 1'b1 && M_out_3 !== M_out_3_ref) begin
          M_out_3_testFailure <= 1'b1;
          $display("ERROR in M_out_3 at time %t : Expected '%h' Actual '%h'", $time, M_out_3_ref, M_out_3);
        end
      end
    end
  // Data source for M_out_0_4_expected
  assign M_out_0_4_expected_1 = 14'b11011111111111;
  assign M_out_4_ref = M_out_0_4_expected_1;
  always @(posedge clk or posedge reset)
    begin : M_out_4_checker
      if (reset == 1'b1) begin
        M_out_4_testFailure <= 1'b0;
      end
      else begin
        if (ce_out == 1'b1 && M_out_4 !== M_out_4_ref) begin
          M_out_4_testFailure <= 1'b1;
          $display("ERROR in M_out_4 at time %t : Expected '%h' Actual '%h'", $time, M_out_4_ref, M_out_4);
        end
      end
    end
  // Data source for M_out_0_5_expected
  assign M_out_0_5_expected_1 = 14'b11011111111111;
  assign M_out_5_ref = M_out_0_5_expected_1;
  always @(posedge clk or posedge reset)
    begin : M_out_5_checker
      if (reset == 1'b1) begin
        M_out_5_testFailure <= 1'b0;
      end
      else begin
        if (ce_out == 1'b1 && M_out_5 !== M_out_5_ref) begin
          M_out_5_testFailure <= 1'b1;
          $display("ERROR in M_out_5 at time %t : Expected '%h' Actual '%h'", $time, M_out_5_ref, M_out_5);
        end
      end
    end
  // Data source for M_out_0_6_expected
  assign M_out_0_6_expected_1 = 14'b11011111111111;
  assign M_out_6_ref = M_out_0_6_expected_1;
  always @(posedge clk or posedge reset)
    begin : M_out_6_checker
      if (reset == 1'b1) begin
        M_out_6_testFailure <= 1'b0;
      end
      else begin
        if (ce_out == 1'b1 && M_out_6 !== M_out_6_ref) begin
          M_out_6_testFailure <= 1'b1;
          $display("ERROR in M_out_6 at time %t : Expected '%h' Actual '%h'", $time, M_out_6_ref, M_out_6);
        end
      end
    end
  // Data source for M_out_0_7_expected
  assign M_out_0_7_expected_1 = 14'b11011111111111;
  assign M_out_7_ref = M_out_0_7_expected_1;
  always @(posedge clk or posedge reset)
    begin : M_out_7_checker
      if (reset == 1'b1) begin
        M_out_7_testFailure <= 1'b0;
      end
      else begin
        if (ce_out == 1'b1 && M_out_7 !== M_out_7_ref) begin
          M_out_7_testFailure <= 1'b1;
          $display("ERROR in M_out_7 at time %t : Expected '%h' Actual '%h'", $time, M_out_7_ref, M_out_7);
        end
      end
    end
  // Data source for M_out_0_8_expected
  assign M_out_0_8_expected_1 = 14'b11011111111111;
  assign M_out_8_ref = M_out_0_8_expected_1;
  always @(posedge clk or posedge reset)
    begin : M_out_8_checker
      if (reset == 1'b1) begin
        M_out_8_testFailure <= 1'b0;
      end
      else begin
        if (ce_out == 1'b1 && M_out_8 !== M_out_8_ref) begin
          M_out_8_testFailure <= 1'b1;
          $display("ERROR in M_out_8 at time %t : Expected '%h' Actual '%h'", $time, M_out_8_ref, M_out_8);
        end
      end
    end
  // Data source for M_out_0_9_expected
  assign M_out_0_9_expected_1 = 14'b11011111111111;
  assign M_out_9_ref = M_out_0_9_expected_1;
  always @(posedge clk or posedge reset)
    begin : M_out_9_checker
      if (reset == 1'b1) begin
        M_out_9_testFailure <= 1'b0;
      end
      else begin
        if (ce_out == 1'b1 && M_out_9 !== M_out_9_ref) begin
          M_out_9_testFailure <= 1'b1;
          $display("ERROR in M_out_9 at time %t : Expected '%h' Actual '%h'", $time, M_out_9_ref, M_out_9);
        end
      end
    end
  // Data source for M_out_0_10_expected
  assign M_out_0_10_expected_1 = 14'b11011111111111;
  assign M_out_10_ref = M_out_0_10_expected_1;
  always @(posedge clk or posedge reset)
    begin : M_out_10_checker
      if (reset == 1'b1) begin
        M_out_10_testFailure <= 1'b0;
      end
      else begin
        if (ce_out == 1'b1 && M_out_10 !== M_out_10_ref) begin
          M_out_10_testFailure <= 1'b1;
          $display("ERROR in M_out_10 at time %t : Expected '%h' Actual '%h'", $time, M_out_10_ref, M_out_10);
        end
      end
    end
  // Data source for M_out_0_11_expected
  assign M_out_0_11_expected_1 = 14'b11011111111111;
  assign M_out_11_ref = M_out_0_11_expected_1;
  always @(posedge clk or posedge reset)
    begin : M_out_11_checker
      if (reset == 1'b1) begin
        M_out_11_testFailure <= 1'b0;
      end
      else begin
        if (ce_out == 1'b1 && M_out_11 !== M_out_11_ref) begin
          M_out_11_testFailure <= 1'b1;
          $display("ERROR in M_out_11 at time %t : Expected '%h' Actual '%h'", $time, M_out_11_ref, M_out_11);
        end
      end
    end
  // Data source for M_out_0_12_expected
  assign M_out_0_12_expected_1 = 14'b11011111111111;
  assign M_out_12_ref = M_out_0_12_expected_1;
  always @(posedge clk or posedge reset)
    begin : M_out_12_checker
      if (reset == 1'b1) begin
        M_out_12_testFailure <= 1'b0;
      end
      else begin
        if (ce_out == 1'b1 && M_out_12 !== M_out_12_ref) begin
          M_out_12_testFailure <= 1'b1;
          $display("ERROR in M_out_12 at time %t : Expected '%h' Actual '%h'", $time, M_out_12_ref, M_out_12);
        end
      end
    end
  // Data source for M_out_0_13_expected
  assign M_out_0_13_expected_1 = 14'b11011111111111;
  assign M_out_13_ref = M_out_0_13_expected_1;
  always @(posedge clk or posedge reset)
    begin : M_out_13_checker
      if (reset == 1'b1) begin
        M_out_13_testFailure <= 1'b0;
      end
      else begin
        if (ce_out == 1'b1 && M_out_13 !== M_out_13_ref) begin
          M_out_13_testFailure <= 1'b1;
          $display("ERROR in M_out_13 at time %t : Expected '%h' Actual '%h'", $time, M_out_13_ref, M_out_13);
        end
      end
    end
  // Data source for M_out_0_14_expected
  assign M_out_0_14_expected_1 = 14'b11011111111111;
  assign M_out_14_ref = M_out_0_14_expected_1;
  always @(posedge clk or posedge reset)
    begin : M_out_14_checker
      if (reset == 1'b1) begin
        M_out_14_testFailure <= 1'b0;
      end
      else begin
        if (ce_out == 1'b1 && M_out_14 !== M_out_14_ref) begin
          M_out_14_testFailure <= 1'b1;
          $display("ERROR in M_out_14 at time %t : Expected '%h' Actual '%h'", $time, M_out_14_ref, M_out_14);
        end
      end
    end
  // Data source for M_out_0_15_expected
  assign M_out_0_15_expected_1 = 14'b11011111111111;
  assign M_out_15_ref = M_out_0_15_expected_1;
  always @(posedge clk or posedge reset)
    begin : M_out_15_checker
      if (reset == 1'b1) begin
        M_out_15_testFailure <= 1'b0;
      end
      else begin
        if (ce_out == 1'b1 && M_out_15 !== M_out_15_ref) begin
          M_out_15_testFailure <= 1'b1;
          $display("ERROR in M_out_15 at time %t : Expected '%h' Actual '%h'", $time, M_out_15_ref, M_out_15);
        end
      end
    end
  // Data source for M_out_0_16_expected
  assign M_out_0_16_expected_1 = 14'b11011111111111;
  assign M_out_16_ref = M_out_0_16_expected_1;
  always @(posedge clk or posedge reset)
    begin : M_out_16_checker
      if (reset == 1'b1) begin
        M_out_16_testFailure <= 1'b0;
      end
      else begin
        if (ce_out == 1'b1 && M_out_16 !== M_out_16_ref) begin
          M_out_16_testFailure <= 1'b1;
          $display("ERROR in M_out_16 at time %t : Expected '%h' Actual '%h'", $time, M_out_16_ref, M_out_16);
        end
      end
    end
  // Data source for M_out_0_17_expected
  assign M_out_0_17_expected_1 = 14'b11011111111111;
  assign M_out_17_ref = M_out_0_17_expected_1;
  always @(posedge clk or posedge reset)
    begin : M_out_17_checker
      if (reset == 1'b1) begin
        M_out_17_testFailure <= 1'b0;
      end
      else begin
        if (ce_out == 1'b1 && M_out_17 !== M_out_17_ref) begin
          M_out_17_testFailure <= 1'b1;
          $display("ERROR in M_out_17 at time %t : Expected '%h' Actual '%h'", $time, M_out_17_ref, M_out_17);
        end
      end
    end
  // Data source for M_out_0_18_expected
  assign M_out_0_18_expected_1 = 14'b11011111111111;
  assign M_out_18_ref = M_out_0_18_expected_1;
  always @(posedge clk or posedge reset)
    begin : M_out_18_checker
      if (reset == 1'b1) begin
        M_out_18_testFailure <= 1'b0;
      end
      else begin
        if (ce_out == 1'b1 && M_out_18 !== M_out_18_ref) begin
          M_out_18_testFailure <= 1'b1;
          $display("ERROR in M_out_18 at time %t : Expected '%h' Actual '%h'", $time, M_out_18_ref, M_out_18);
        end
      end
    end
  // Data source for M_out_0_19_expected
  assign M_out_0_19_expected_1 = 14'b11011111111111;
  assign M_out_19_ref = M_out_0_19_expected_1;
  always @(posedge clk or posedge reset)
    begin : M_out_19_checker
      if (reset == 1'b1) begin
        M_out_19_testFailure <= 1'b0;
      end
      else begin
        if (ce_out == 1'b1 && M_out_19 !== M_out_19_ref) begin
          M_out_19_testFailure <= 1'b1;
          $display("ERROR in M_out_19 at time %t : Expected '%h' Actual '%h'", $time, M_out_19_ref, M_out_19);
        end
      end
    end
  // Data source for M_out_0_20_expected
  assign M_out_0_20_expected_1 = 14'b11011111111111;
  assign M_out_20_ref = M_out_0_20_expected_1;
  always @(posedge clk or posedge reset)
    begin : M_out_20_checker
      if (reset == 1'b1) begin
        M_out_20_testFailure <= 1'b0;
      end
      else begin
        if (ce_out == 1'b1 && M_out_20 !== M_out_20_ref) begin
          M_out_20_testFailure <= 1'b1;
          $display("ERROR in M_out_20 at time %t : Expected '%h' Actual '%h'", $time, M_out_20_ref, M_out_20);
        end
      end
    end
  // Data source for M_out_0_21_expected
  assign M_out_0_21_expected_1 = 14'b11011111111111;
  assign M_out_21_ref = M_out_0_21_expected_1;
  always @(posedge clk or posedge reset)
    begin : M_out_21_checker
      if (reset == 1'b1) begin
        M_out_21_testFailure <= 1'b0;
      end
      else begin
        if (ce_out == 1'b1 && M_out_21 !== M_out_21_ref) begin
          M_out_21_testFailure <= 1'b1;
          $display("ERROR in M_out_21 at time %t : Expected '%h' Actual '%h'", $time, M_out_21_ref, M_out_21);
        end
      end
    end
  // Data source for M_out_0_22_expected
  assign M_out_0_22_expected_1 = 14'b11011111111111;
  assign M_out_22_ref = M_out_0_22_expected_1;
  always @(posedge clk or posedge reset)
    begin : M_out_22_checker
      if (reset == 1'b1) begin
        M_out_22_testFailure <= 1'b0;
      end
      else begin
        if (ce_out == 1'b1 && M_out_22 !== M_out_22_ref) begin
          M_out_22_testFailure <= 1'b1;
          $display("ERROR in M_out_22 at time %t : Expected '%h' Actual '%h'", $time, M_out_22_ref, M_out_22);
        end
      end
    end
  // Data source for M_out_0_23_expected
  assign M_out_0_23_expected_1 = 14'b11011111111111;
  assign M_out_23_ref = M_out_0_23_expected_1;
  always @(posedge clk or posedge reset)
    begin : M_out_23_checker
      if (reset == 1'b1) begin
        M_out_23_testFailure <= 1'b0;
      end
      else begin
        if (ce_out == 1'b1 && M_out_23 !== M_out_23_ref) begin
          M_out_23_testFailure <= 1'b1;
          $display("ERROR in M_out_23 at time %t : Expected '%h' Actual '%h'", $time, M_out_23_ref, M_out_23);
        end
      end
    end
  // Data source for M_out_0_24_expected
  assign M_out_0_24_expected_1 = 14'b11011111111111;
  assign M_out_24_ref = M_out_0_24_expected_1;
  always @(posedge clk or posedge reset)
    begin : M_out_24_checker
      if (reset == 1'b1) begin
        M_out_24_testFailure <= 1'b0;
      end
      else begin
        if (ce_out == 1'b1 && M_out_24 !== M_out_24_ref) begin
          M_out_24_testFailure <= 1'b1;
          $display("ERROR in M_out_24 at time %t : Expected '%h' Actual '%h'", $time, M_out_24_ref, M_out_24);
        end
      end
    end
  // Data source for M_out_0_25_expected
  assign M_out_0_25_expected_1 = 14'b11011111111111;
  assign M_out_25_ref = M_out_0_25_expected_1;
  always @(posedge clk or posedge reset)
    begin : M_out_25_checker
      if (reset == 1'b1) begin
        M_out_25_testFailure <= 1'b0;
      end
      else begin
        if (ce_out == 1'b1 && M_out_25 !== M_out_25_ref) begin
          M_out_25_testFailure <= 1'b1;
          $display("ERROR in M_out_25 at time %t : Expected '%h' Actual '%h'", $time, M_out_25_ref, M_out_25);
        end
      end
    end
  // Data source for M_out_0_26_expected
  assign M_out_0_26_expected_1 = 14'b11011111111111;
  assign M_out_26_ref = M_out_0_26_expected_1;
  always @(posedge clk or posedge reset)
    begin : M_out_26_checker
      if (reset == 1'b1) begin
        M_out_26_testFailure <= 1'b0;
      end
      else begin
        if (ce_out == 1'b1 && M_out_26 !== M_out_26_ref) begin
          M_out_26_testFailure <= 1'b1;
          $display("ERROR in M_out_26 at time %t : Expected '%h' Actual '%h'", $time, M_out_26_ref, M_out_26);
        end
      end
    end
  // Data source for M_out_0_27_expected
  assign M_out_0_27_expected_1 = 14'b11011111111111;
  assign M_out_27_ref = M_out_0_27_expected_1;
  always @(posedge clk or posedge reset)
    begin : M_out_27_checker
      if (reset == 1'b1) begin
        M_out_27_testFailure <= 1'b0;
      end
      else begin
        if (ce_out == 1'b1 && M_out_27 !== M_out_27_ref) begin
          M_out_27_testFailure <= 1'b1;
          $display("ERROR in M_out_27 at time %t : Expected '%h' Actual '%h'", $time, M_out_27_ref, M_out_27);
        end
      end
    end
  // Data source for M_out_0_28_expected
  assign M_out_0_28_expected_1 = 14'b11011111111111;
  assign M_out_28_ref = M_out_0_28_expected_1;
  always @(posedge clk or posedge reset)
    begin : M_out_28_checker
      if (reset == 1'b1) begin
        M_out_28_testFailure <= 1'b0;
      end
      else begin
        if (ce_out == 1'b1 && M_out_28 !== M_out_28_ref) begin
          M_out_28_testFailure <= 1'b1;
          $display("ERROR in M_out_28 at time %t : Expected '%h' Actual '%h'", $time, M_out_28_ref, M_out_28);
        end
      end
    end
  // Data source for M_out_0_29_expected
  assign M_out_0_29_expected_1 = 14'b11011111111111;
  assign M_out_29_ref = M_out_0_29_expected_1;
  always @(posedge clk or posedge reset)
    begin : M_out_29_checker
      if (reset == 1'b1) begin
        M_out_29_testFailure <= 1'b0;
      end
      else begin
        if (ce_out == 1'b1 && M_out_29 !== M_out_29_ref) begin
          M_out_29_testFailure <= 1'b1;
          $display("ERROR in M_out_29 at time %t : Expected '%h' Actual '%h'", $time, M_out_29_ref, M_out_29);
        end
      end
    end
  // Data source for M_out_0_30_expected
  assign M_out_0_30_expected_1 = 14'b11011111111111;
  assign M_out_30_ref = M_out_0_30_expected_1;
  always @(posedge clk or posedge reset)
    begin : M_out_30_checker
      if (reset == 1'b1) begin
        M_out_30_testFailure <= 1'b0;
      end
      else begin
        if (ce_out == 1'b1 && M_out_30 !== M_out_30_ref) begin
          M_out_30_testFailure <= 1'b1;
          $display("ERROR in M_out_30 at time %t : Expected '%h' Actual '%h'", $time, M_out_30_ref, M_out_30);
        end
      end
    end
  // Data source for M_out_0_31_expected
  assign M_out_0_31_expected_1 = 14'b11011111111111;
  assign M_out_31_ref = M_out_0_31_expected_1;
  always @(posedge clk or posedge reset)
    begin : M_out_31_checker
      if (reset == 1'b1) begin
        M_out_31_testFailure <= 1'b0;
      end
      else begin
        if (ce_out == 1'b1 && M_out_31 !== M_out_31_ref) begin
          M_out_31_testFailure <= 1'b1;
          $display("ERROR in M_out_31 at time %t : Expected '%h' Actual '%h'", $time, M_out_31_ref, M_out_31);
        end
      end
    end
  // Data source for M_out_0_32_expected
  assign M_out_0_32_expected_1 = 14'b11011111111111;
  assign M_out_32_ref = M_out_0_32_expected_1;
  always @(posedge clk or posedge reset)
    begin : M_out_32_checker
      if (reset == 1'b1) begin
        M_out_32_testFailure <= 1'b0;
      end
      else begin
        if (ce_out == 1'b1 && M_out_32 !== M_out_32_ref) begin
          M_out_32_testFailure <= 1'b1;
          $display("ERROR in M_out_32 at time %t : Expected '%h' Actual '%h'", $time, M_out_32_ref, M_out_32);
        end
      end
    end
  // Data source for M_out_0_33_expected
  assign M_out_0_33_expected_1 = 14'b11011111111111;
  assign M_out_33_ref = M_out_0_33_expected_1;
  always @(posedge clk or posedge reset)
    begin : M_out_33_checker
      if (reset == 1'b1) begin
        M_out_33_testFailure <= 1'b0;
      end
      else begin
        if (ce_out == 1'b1 && M_out_33 !== M_out_33_ref) begin
          M_out_33_testFailure <= 1'b1;
          $display("ERROR in M_out_33 at time %t : Expected '%h' Actual '%h'", $time, M_out_33_ref, M_out_33);
        end
      end
    end
  // Data source for M_out_0_34_expected
  assign M_out_0_34_expected_1 = 14'b11011111111111;
  assign M_out_34_ref = M_out_0_34_expected_1;
  always @(posedge clk or posedge reset)
    begin : M_out_34_checker
      if (reset == 1'b1) begin
        M_out_34_testFailure <= 1'b0;
      end
      else begin
        if (ce_out == 1'b1 && M_out_34 !== M_out_34_ref) begin
          M_out_34_testFailure <= 1'b1;
          $display("ERROR in M_out_34 at time %t : Expected '%h' Actual '%h'", $time, M_out_34_ref, M_out_34);
        end
      end
    end
  // Data source for M_out_0_35_expected
  assign M_out_0_35_expected_1 = 14'b11011111111111;
  assign M_out_35_ref = M_out_0_35_expected_1;
  always @(posedge clk or posedge reset)
    begin : M_out_35_checker
      if (reset == 1'b1) begin
        M_out_35_testFailure <= 1'b0;
      end
      else begin
        if (ce_out == 1'b1 && M_out_35 !== M_out_35_ref) begin
          M_out_35_testFailure <= 1'b1;
          $display("ERROR in M_out_35 at time %t : Expected '%h' Actual '%h'", $time, M_out_35_ref, M_out_35);
        end
      end
    end
  // Data source for M_out_0_36_expected
  assign M_out_0_36_expected_1 = 14'b11011111111111;
  assign M_out_36_ref = M_out_0_36_expected_1;
  always @(posedge clk or posedge reset)
    begin : M_out_36_checker
      if (reset == 1'b1) begin
        M_out_36_testFailure <= 1'b0;
      end
      else begin
        if (ce_out == 1'b1 && M_out_36 !== M_out_36_ref) begin
          M_out_36_testFailure <= 1'b1;
          $display("ERROR in M_out_36 at time %t : Expected '%h' Actual '%h'", $time, M_out_36_ref, M_out_36);
        end
      end
    end
  // Data source for M_out_0_37_expected
  assign M_out_0_37_expected_1 = 14'b11011111111111;
  assign M_out_37_ref = M_out_0_37_expected_1;
  always @(posedge clk or posedge reset)
    begin : M_out_37_checker
      if (reset == 1'b1) begin
        M_out_37_testFailure <= 1'b0;
      end
      else begin
        if (ce_out == 1'b1 && M_out_37 !== M_out_37_ref) begin
          M_out_37_testFailure <= 1'b1;
          $display("ERROR in M_out_37 at time %t : Expected '%h' Actual '%h'", $time, M_out_37_ref, M_out_37);
        end
      end
    end
  // Data source for M_out_0_38_expected
  assign M_out_0_38_expected_1 = 14'b11011111111111;
  assign M_out_38_ref = M_out_0_38_expected_1;
  always @(posedge clk or posedge reset)
    begin : M_out_38_checker
      if (reset == 1'b1) begin
        M_out_38_testFailure <= 1'b0;
      end
      else begin
        if (ce_out == 1'b1 && M_out_38 !== M_out_38_ref) begin
          M_out_38_testFailure <= 1'b1;
          $display("ERROR in M_out_38 at time %t : Expected '%h' Actual '%h'", $time, M_out_38_ref, M_out_38);
        end
      end
    end
  // Data source for M_out_0_39_expected
  assign M_out_0_39_expected_1 = 14'b11011111111111;
  assign M_out_39_ref = M_out_0_39_expected_1;
  always @(posedge clk or posedge reset)
    begin : M_out_39_checker
      if (reset == 1'b1) begin
        M_out_39_testFailure <= 1'b0;
      end
      else begin
        if (ce_out == 1'b1 && M_out_39 !== M_out_39_ref) begin
          M_out_39_testFailure <= 1'b1;
          $display("ERROR in M_out_39 at time %t : Expected '%h' Actual '%h'", $time, M_out_39_ref, M_out_39);
        end
      end
    end
  // Data source for M_out_0_40_expected
  assign M_out_0_40_expected_1 = 14'b11011111111111;
  assign M_out_40_ref = M_out_0_40_expected_1;
  always @(posedge clk or posedge reset)
    begin : M_out_40_checker
      if (reset == 1'b1) begin
        M_out_40_testFailure <= 1'b0;
      end
      else begin
        if (ce_out == 1'b1 && M_out_40 !== M_out_40_ref) begin
          M_out_40_testFailure <= 1'b1;
          $display("ERROR in M_out_40 at time %t : Expected '%h' Actual '%h'", $time, M_out_40_ref, M_out_40);
        end
      end
    end
  // Data source for M_out_0_41_expected
  assign M_out_0_41_expected_1 = 14'b11011111111111;
  assign M_out_41_ref = M_out_0_41_expected_1;
  always @(posedge clk or posedge reset)
    begin : M_out_41_checker
      if (reset == 1'b1) begin
        M_out_41_testFailure <= 1'b0;
      end
      else begin
        if (ce_out == 1'b1 && M_out_41 !== M_out_41_ref) begin
          M_out_41_testFailure <= 1'b1;
          $display("ERROR in M_out_41 at time %t : Expected '%h' Actual '%h'", $time, M_out_41_ref, M_out_41);
        end
      end
    end
  // Data source for M_out_0_42_expected
  assign M_out_0_42_expected_1 = 14'b11011111111111;
  assign M_out_42_ref = M_out_0_42_expected_1;
  always @(posedge clk or posedge reset)
    begin : M_out_42_checker
      if (reset == 1'b1) begin
        M_out_42_testFailure <= 1'b0;
      end
      else begin
        if (ce_out == 1'b1 && M_out_42 !== M_out_42_ref) begin
          M_out_42_testFailure <= 1'b1;
          $display("ERROR in M_out_42 at time %t : Expected '%h' Actual '%h'", $time, M_out_42_ref, M_out_42);
        end
      end
    end
  // Data source for M_out_0_43_expected
  assign M_out_0_43_expected_1 = 14'b11011111111111;
  assign M_out_43_ref = M_out_0_43_expected_1;
  always @(posedge clk or posedge reset)
    begin : M_out_43_checker
      if (reset == 1'b1) begin
        M_out_43_testFailure <= 1'b0;
      end
      else begin
        if (ce_out == 1'b1 && M_out_43 !== M_out_43_ref) begin
          M_out_43_testFailure <= 1'b1;
          $display("ERROR in M_out_43 at time %t : Expected '%h' Actual '%h'", $time, M_out_43_ref, M_out_43);
        end
      end
    end
  // Data source for M_out_0_44_expected
  assign M_out_0_44_expected_1 = 14'b11011111111111;
  assign M_out_44_ref = M_out_0_44_expected_1;
  always @(posedge clk or posedge reset)
    begin : M_out_44_checker
      if (reset == 1'b1) begin
        M_out_44_testFailure <= 1'b0;
      end
      else begin
        if (ce_out == 1'b1 && M_out_44 !== M_out_44_ref) begin
          M_out_44_testFailure <= 1'b1;
          $display("ERROR in M_out_44 at time %t : Expected '%h' Actual '%h'", $time, M_out_44_ref, M_out_44);
        end
      end
    end
  // Data source for M_out_0_45_expected
  assign M_out_0_45_expected_1 = 14'b11011111111111;
  assign M_out_45_ref = M_out_0_45_expected_1;
  always @(posedge clk or posedge reset)
    begin : M_out_45_checker
      if (reset == 1'b1) begin
        M_out_45_testFailure <= 1'b0;
      end
      else begin
        if (ce_out == 1'b1 && M_out_45 !== M_out_45_ref) begin
          M_out_45_testFailure <= 1'b1;
          $display("ERROR in M_out_45 at time %t : Expected '%h' Actual '%h'", $time, M_out_45_ref, M_out_45);
        end
      end
    end
  // Data source for M_out_0_46_expected
  assign M_out_0_46_expected_1 = 14'b11011111111111;
  assign M_out_46_ref = M_out_0_46_expected_1;
  always @(posedge clk or posedge reset)
    begin : M_out_46_checker
      if (reset == 1'b1) begin
        M_out_46_testFailure <= 1'b0;
      end
      else begin
        if (ce_out == 1'b1 && M_out_46 !== M_out_46_ref) begin
          M_out_46_testFailure <= 1'b1;
          $display("ERROR in M_out_46 at time %t : Expected '%h' Actual '%h'", $time, M_out_46_ref, M_out_46);
        end
      end
    end
  // Data source for M_out_0_47_expected
  assign M_out_0_47_expected_1 = 14'b11011111111111;
  assign M_out_47_ref = M_out_0_47_expected_1;
  always @(posedge clk or posedge reset)
    begin : M_out_47_checker
      if (reset == 1'b1) begin
        M_out_47_testFailure <= 1'b0;
      end
      else begin
        if (ce_out == 1'b1 && M_out_47 !== M_out_47_ref) begin
          M_out_47_testFailure <= 1'b1;
          $display("ERROR in M_out_47 at time %t : Expected '%h' Actual '%h'", $time, M_out_47_ref, M_out_47);
        end
      end
    end
  // Data source for M_out_0_48_expected
  assign M_out_0_48_expected_1 = 14'b11011111111111;
  assign M_out_48_ref = M_out_0_48_expected_1;
  always @(posedge clk or posedge reset)
    begin : M_out_48_checker
      if (reset == 1'b1) begin
        M_out_48_testFailure <= 1'b0;
      end
      else begin
        if (ce_out == 1'b1 && M_out_48 !== M_out_48_ref) begin
          M_out_48_testFailure <= 1'b1;
          $display("ERROR in M_out_48 at time %t : Expected '%h' Actual '%h'", $time, M_out_48_ref, M_out_48);
        end
      end
    end
  // Data source for M_out_0_49_expected
  assign M_out_0_49_expected_1 = 14'b11011111111111;
  assign M_out_49_ref = M_out_0_49_expected_1;
  always @(posedge clk or posedge reset)
    begin : M_out_49_checker
      if (reset == 1'b1) begin
        M_out_49_testFailure <= 1'b0;
      end
      else begin
        if (ce_out == 1'b1 && M_out_49 !== M_out_49_ref) begin
          M_out_49_testFailure <= 1'b1;
          $display("ERROR in M_out_49 at time %t : Expected '%h' Actual '%h'", $time, M_out_49_ref, M_out_49);
        end
      end
    end
  // Data source for M_out_0_50_expected
  assign M_out_0_50_expected_1 = 14'b11011111111111;
  assign M_out_50_ref = M_out_0_50_expected_1;
  always @(posedge clk or posedge reset)
    begin : M_out_50_checker
      if (reset == 1'b1) begin
        M_out_50_testFailure <= 1'b0;
      end
      else begin
        if (ce_out == 1'b1 && M_out_50 !== M_out_50_ref) begin
          M_out_50_testFailure <= 1'b1;
          $display("ERROR in M_out_50 at time %t : Expected '%h' Actual '%h'", $time, M_out_50_ref, M_out_50);
        end
      end
    end
  // Data source for M_out_0_51_expected
  assign M_out_0_51_expected_1 = 14'b11011111111111;
  assign M_out_51_ref = M_out_0_51_expected_1;
  always @(posedge clk or posedge reset)
    begin : M_out_51_checker
      if (reset == 1'b1) begin
        M_out_51_testFailure <= 1'b0;
      end
      else begin
        if (ce_out == 1'b1 && M_out_51 !== M_out_51_ref) begin
          M_out_51_testFailure <= 1'b1;
          $display("ERROR in M_out_51 at time %t : Expected '%h' Actual '%h'", $time, M_out_51_ref, M_out_51);
        end
      end
    end
  // Data source for M_out_0_52_expected
  assign M_out_0_52_expected_1 = 14'b11011111111111;
  assign M_out_52_ref = M_out_0_52_expected_1;
  always @(posedge clk or posedge reset)
    begin : M_out_52_checker
      if (reset == 1'b1) begin
        M_out_52_testFailure <= 1'b0;
      end
      else begin
        if (ce_out == 1'b1 && M_out_52 !== M_out_52_ref) begin
          M_out_52_testFailure <= 1'b1;
          $display("ERROR in M_out_52 at time %t : Expected '%h' Actual '%h'", $time, M_out_52_ref, M_out_52);
        end
      end
    end
  // Data source for M_out_0_53_expected
  assign M_out_0_53_expected_1 = 14'b11011111111111;
  assign M_out_53_ref = M_out_0_53_expected_1;
  always @(posedge clk or posedge reset)
    begin : M_out_53_checker
      if (reset == 1'b1) begin
        M_out_53_testFailure <= 1'b0;
      end
      else begin
        if (ce_out == 1'b1 && M_out_53 !== M_out_53_ref) begin
          M_out_53_testFailure <= 1'b1;
          $display("ERROR in M_out_53 at time %t : Expected '%h' Actual '%h'", $time, M_out_53_ref, M_out_53);
        end
      end
    end
  // Data source for M_out_0_54_expected
  assign M_out_0_54_expected_1 = 14'b11011111111111;
  assign M_out_54_ref = M_out_0_54_expected_1;
  always @(posedge clk or posedge reset)
    begin : M_out_54_checker
      if (reset == 1'b1) begin
        M_out_54_testFailure <= 1'b0;
      end
      else begin
        if (ce_out == 1'b1 && M_out_54 !== M_out_54_ref) begin
          M_out_54_testFailure <= 1'b1;
          $display("ERROR in M_out_54 at time %t : Expected '%h' Actual '%h'", $time, M_out_54_ref, M_out_54);
        end
      end
    end
  // Data source for M_out_0_55_expected
  assign M_out_0_55_expected_1 = 14'b11011111111111;
  assign M_out_55_ref = M_out_0_55_expected_1;
  always @(posedge clk or posedge reset)
    begin : M_out_55_checker
      if (reset == 1'b1) begin
        M_out_55_testFailure <= 1'b0;
      end
      else begin
        if (ce_out == 1'b1 && M_out_55 !== M_out_55_ref) begin
          M_out_55_testFailure <= 1'b1;
          $display("ERROR in M_out_55 at time %t : Expected '%h' Actual '%h'", $time, M_out_55_ref, M_out_55);
        end
      end
    end
  // Data source for M_out_0_56_expected
  assign M_out_0_56_expected_1 = 14'b11011111111111;
  assign M_out_56_ref = M_out_0_56_expected_1;
  always @(posedge clk or posedge reset)
    begin : M_out_56_checker
      if (reset == 1'b1) begin
        M_out_56_testFailure <= 1'b0;
      end
      else begin
        if (ce_out == 1'b1 && M_out_56 !== M_out_56_ref) begin
          M_out_56_testFailure <= 1'b1;
          $display("ERROR in M_out_56 at time %t : Expected '%h' Actual '%h'", $time, M_out_56_ref, M_out_56);
        end
      end
    end
  // Data source for M_out_0_57_expected
  assign M_out_0_57_expected_1 = 14'b11011111111111;
  assign M_out_57_ref = M_out_0_57_expected_1;
  always @(posedge clk or posedge reset)
    begin : M_out_57_checker
      if (reset == 1'b1) begin
        M_out_57_testFailure <= 1'b0;
      end
      else begin
        if (ce_out == 1'b1 && M_out_57 !== M_out_57_ref) begin
          M_out_57_testFailure <= 1'b1;
          $display("ERROR in M_out_57 at time %t : Expected '%h' Actual '%h'", $time, M_out_57_ref, M_out_57);
        end
      end
    end
  // Data source for M_out_0_58_expected
  assign M_out_0_58_expected_1 = 14'b11011111111111;
  assign M_out_58_ref = M_out_0_58_expected_1;
  always @(posedge clk or posedge reset)
    begin : M_out_58_checker
      if (reset == 1'b1) begin
        M_out_58_testFailure <= 1'b0;
      end
      else begin
        if (ce_out == 1'b1 && M_out_58 !== M_out_58_ref) begin
          M_out_58_testFailure <= 1'b1;
          $display("ERROR in M_out_58 at time %t : Expected '%h' Actual '%h'", $time, M_out_58_ref, M_out_58);
        end
      end
    end
  // Data source for M_out_0_59_expected
  assign M_out_0_59_expected_1 = 14'b11011111111111;
  assign M_out_59_ref = M_out_0_59_expected_1;
  always @(posedge clk or posedge reset)
    begin : M_out_59_checker
      if (reset == 1'b1) begin
        M_out_59_testFailure <= 1'b0;
      end
      else begin
        if (ce_out == 1'b1 && M_out_59 !== M_out_59_ref) begin
          M_out_59_testFailure <= 1'b1;
          $display("ERROR in M_out_59 at time %t : Expected '%h' Actual '%h'", $time, M_out_59_ref, M_out_59);
        end
      end
    end
  // Data source for M_out_0_60_expected
  assign M_out_0_60_expected_1 = 14'b11011111111111;
  assign M_out_60_ref = M_out_0_60_expected_1;
  always @(posedge clk or posedge reset)
    begin : M_out_60_checker
      if (reset == 1'b1) begin
        M_out_60_testFailure <= 1'b0;
      end
      else begin
        if (ce_out == 1'b1 && M_out_60 !== M_out_60_ref) begin
          M_out_60_testFailure <= 1'b1;
          $display("ERROR in M_out_60 at time %t : Expected '%h' Actual '%h'", $time, M_out_60_ref, M_out_60);
        end
      end
    end
  // Data source for M_out_0_61_expected
  assign M_out_0_61_expected_1 = 14'b11011111111111;
  assign M_out_61_ref = M_out_0_61_expected_1;
  always @(posedge clk or posedge reset)
    begin : M_out_61_checker
      if (reset == 1'b1) begin
        M_out_61_testFailure <= 1'b0;
      end
      else begin
        if (ce_out == 1'b1 && M_out_61 !== M_out_61_ref) begin
          M_out_61_testFailure <= 1'b1;
          $display("ERROR in M_out_61 at time %t : Expected '%h' Actual '%h'", $time, M_out_61_ref, M_out_61);
        end
      end
    end
  // Data source for M_out_0_62_expected
  assign M_out_0_62_expected_1 = 14'b11011111111111;
  assign M_out_62_ref = M_out_0_62_expected_1;
  always @(posedge clk or posedge reset)
    begin : M_out_62_checker
      if (reset == 1'b1) begin
        M_out_62_testFailure <= 1'b0;
      end
      else begin
        if (ce_out == 1'b1 && M_out_62 !== M_out_62_ref) begin
          M_out_62_testFailure <= 1'b1;
          $display("ERROR in M_out_62 at time %t : Expected '%h' Actual '%h'", $time, M_out_62_ref, M_out_62);
        end
      end
    end
  // Data source for M_out_0_63_expected
  assign M_out_0_63_expected_1 = 14'b11011111111111;
  assign M_out_63_ref = M_out_0_63_expected_1;
  always @(posedge clk or posedge reset)
    begin : M_out_63_checker
      if (reset == 1'b1) begin
        M_out_63_testFailure <= 1'b0;
      end
      else begin
        if (ce_out == 1'b1 && M_out_63 !== M_out_63_ref) begin
          M_out_63_testFailure <= 1'b1;
          $display("ERROR in M_out_63 at time %t : Expected '%h' Actual '%h'", $time, M_out_63_ref, M_out_63);
        end
      end
    end
  always @(M_out_0_testFailure, M_out_1_testFailure, M_out_2_testFailure,
       M_out_3_testFailure, M_out_4_testFailure, M_out_5_testFailure,
       M_out_6_testFailure, M_out_7_testFailure, M_out_8_testFailure,
       M_out_9_testFailure, M_out_10_testFailure, M_out_11_testFailure,
       M_out_12_testFailure, M_out_13_testFailure, M_out_14_testFailure,
       M_out_15_testFailure, M_out_16_testFailure, M_out_17_testFailure,
       M_out_18_testFailure, M_out_19_testFailure, M_out_20_testFailure,
       M_out_21_testFailure, M_out_22_testFailure, M_out_23_testFailure,
       M_out_24_testFailure, M_out_25_testFailure, M_out_26_testFailure,
       M_out_27_testFailure, M_out_28_testFailure, M_out_29_testFailure,
       M_out_30_testFailure, M_out_31_testFailure, M_out_32_testFailure,
       M_out_33_testFailure, M_out_34_testFailure, M_out_35_testFailure,
       M_out_36_testFailure, M_out_37_testFailure, M_out_38_testFailure,
       M_out_39_testFailure, M_out_40_testFailure, M_out_41_testFailure,
       M_out_42_testFailure, M_out_43_testFailure, M_out_44_testFailure,
       M_out_45_testFailure, M_out_46_testFailure, M_out_47_testFailure,
       M_out_48_testFailure, M_out_49_testFailure, M_out_50_testFailure,
       M_out_51_testFailure, M_out_52_testFailure, M_out_53_testFailure,
       M_out_54_testFailure, M_out_55_testFailure, M_out_56_testFailure,
       M_out_57_testFailure, M_out_58_testFailure, M_out_59_testFailure,
       M_out_60_testFailure, M_out_61_testFailure, M_out_62_testFailure,
       M_out_63_testFailure) begin
    or_t = M_out_21_testFailure | (M_out_20_testFailure | (M_out_19_testFailure | (M_out_18_testFailure | (M_out_17_testFailure | (M_out_16_testFailure | (M_out_15_testFailure | (M_out_14_testFailure | (M_out_13_testFailure | (M_out_12_testFailure | (M_out_11_testFailure | (M_out_10_testFailure | (M_out_9_testFailure | (M_out_8_testFailure | (M_out_7_testFailure | (M_out_6_testFailure | (M_out_5_testFailure | (M_out_4_testFailure | (M_out_3_testFailure | (M_out_2_testFailure | (M_out_0_testFailure | M_out_1_testFailure))))))))))))))))))));
    or_t = M_out_22_testFailure | or_t;
    or_t = M_out_23_testFailure | or_t;
    or_t = M_out_24_testFailure | or_t;
    or_t = M_out_25_testFailure | or_t;
    or_t = M_out_26_testFailure | or_t;
    or_t = M_out_27_testFailure | or_t;
    or_t = M_out_28_testFailure | or_t;
    or_t = M_out_29_testFailure | or_t;
    or_t = M_out_30_testFailure | or_t;
    or_t = M_out_31_testFailure | or_t;
    or_t = M_out_32_testFailure | or_t;
    or_t = M_out_33_testFailure | or_t;
    or_t = M_out_34_testFailure | or_t;
    or_t = M_out_35_testFailure | or_t;
    or_t = M_out_36_testFailure | or_t;
    or_t = M_out_37_testFailure | or_t;
    or_t = M_out_38_testFailure | or_t;
    or_t = M_out_39_testFailure | or_t;
    or_t = M_out_40_testFailure | or_t;
    or_t = M_out_41_testFailure | or_t;
    or_t = M_out_42_testFailure | or_t;
    or_t = M_out_43_testFailure | or_t;
    or_t = M_out_44_testFailure | or_t;
    or_t = M_out_45_testFailure | or_t;
    or_t = M_out_46_testFailure | or_t;
    or_t = M_out_47_testFailure | or_t;
    or_t = M_out_48_testFailure | or_t;
    or_t = M_out_49_testFailure | or_t;
    or_t = M_out_50_testFailure | or_t;
    or_t = M_out_51_testFailure | or_t;
    or_t = M_out_52_testFailure | or_t;
    or_t = M_out_53_testFailure | or_t;
    or_t = M_out_54_testFailure | or_t;
    or_t = M_out_55_testFailure | or_t;
    or_t = M_out_56_testFailure | or_t;
    or_t = M_out_57_testFailure | or_t;
    or_t = M_out_58_testFailure | or_t;
    or_t = M_out_59_testFailure | or_t;
    or_t = M_out_60_testFailure | or_t;
    or_t = M_out_61_testFailure | or_t;
    or_t = M_out_62_testFailure | or_t;
    or_t = M_out_63_testFailure | or_t;
    testFailure = or_t;
  end
  always @(posedge clk)
    begin : completed_msg
      if (check1_done == 1'b1) begin
        if (testFailure == 1'b0) begin
          $display("**************TEST COMPLETED (PASSED)**************");
        end
        else begin
          $display("**************TEST COMPLETED (FAILED)**************");
        end
      end
    end
endmodule