module outputs
  wire [69 : 0] server_core_response_get;
  wire RDY_server_core_request_put,
       RDY_server_core_response_get,
       RDY_server_reset_request_put,
       RDY_server_reset_response_get;
  // inlined wires
  reg [68 : 0] resWire$wget;
  wire crg_done$EN_port0__write,
       crg_done$EN_port1__write,
       crg_done$port1__read,
       crg_done$port2__read,
       crg_done_1$EN_port0__write,
       crg_done_1$EN_port1__write,
       crg_done_1$port1__read,
       crg_done_1$port2__read,
       resWire$whas;
  // register crg_done
  reg crg_done;
  wire crg_done$D_IN, crg_done$EN;
  // register crg_done_1
  reg crg_done_1;
  wire crg_done_1$D_IN, crg_done_1$EN;
  // register rg_b
  reg [115 : 0] rg_b;
  wire [115 : 0] rg_b$D_IN;
  wire rg_b$EN;
  // register rg_busy
  reg rg_busy;
  wire rg_busy$D_IN, rg_busy$EN;
  // register rg_busy_1
  reg rg_busy_1;
  wire rg_busy_1$D_IN, rg_busy_1$EN;
  // register rg_d
  reg [57 : 0] rg_d;
  wire [57 : 0] rg_d$D_IN;
  wire rg_d$EN;
  // register rg_index
  reg [5 : 0] rg_index;
  wire [5 : 0] rg_index$D_IN;
  wire rg_index$EN;
  // register rg_index_1
  reg [5 : 0] rg_index_1;
  wire [5 : 0] rg_index_1$D_IN;
  wire rg_index_1$EN;
  // register rg_q
  reg [57 : 0] rg_q;
  wire [57 : 0] rg_q$D_IN;
  wire rg_q$EN;
  // register rg_r
  reg [115 : 0] rg_r;
  wire [115 : 0] rg_r$D_IN;
  wire rg_r$EN;
  // register rg_r_1
  reg [115 : 0] rg_r_1;
  wire [115 : 0] rg_r_1$D_IN;
  wire rg_r_1$EN;
  // register rg_res
  reg [116 : 0] rg_res;
  wire [116 : 0] rg_res$D_IN;
  wire rg_res$EN;
  // register rg_s
  reg [115 : 0] rg_s;
  wire [115 : 0] rg_s$D_IN;
  wire rg_s$EN;
  // ports of submodule fpu_div_fOperands_S0
  wire [130 : 0] fpu_div_fOperands_S0$D_IN, fpu_div_fOperands_S0$D_OUT;
  wire fpu_div_fOperands_S0$CLR,
       fpu_div_fOperands_S0$DEQ,
       fpu_div_fOperands_S0$EMPTY_N,
       fpu_div_fOperands_S0$ENQ,
       fpu_div_fOperands_S0$FULL_N;
  // ports of submodule fpu_div_fResult_S5
  wire [68 : 0] fpu_div_fResult_S5$D_IN, fpu_div_fResult_S5$D_OUT;
  wire fpu_div_fResult_S5$CLR,
       fpu_div_fResult_S5$DEQ,
       fpu_div_fResult_S5$EMPTY_N,
       fpu_div_fResult_S5$ENQ,
       fpu_div_fResult_S5$FULL_N;
  // ports of submodule fpu_div_fState_S1
  wire [318 : 0] fpu_div_fState_S1$D_IN, fpu_div_fState_S1$D_OUT;
  wire fpu_div_fState_S1$CLR,
       fpu_div_fState_S1$DEQ,
       fpu_div_fState_S1$EMPTY_N,
       fpu_div_fState_S1$ENQ,
       fpu_div_fState_S1$FULL_N;
  // ports of submodule fpu_div_fState_S2
  wire [147 : 0] fpu_div_fState_S2$D_IN, fpu_div_fState_S2$D_OUT;
  wire fpu_div_fState_S2$CLR,
       fpu_div_fState_S2$DEQ,
       fpu_div_fState_S2$EMPTY_N,
       fpu_div_fState_S2$ENQ,
       fpu_div_fState_S2$FULL_N;
  // ports of submodule fpu_div_fState_S3
  wire [194 : 0] fpu_div_fState_S3$D_IN, fpu_div_fState_S3$D_OUT;
  wire fpu_div_fState_S3$CLR,
       fpu_div_fState_S3$DEQ,
       fpu_div_fState_S3$EMPTY_N,
       fpu_div_fState_S3$ENQ,
       fpu_div_fState_S3$FULL_N;
  // ports of submodule fpu_div_fState_S4
  wire [138 : 0] fpu_div_fState_S4$D_IN, fpu_div_fState_S4$D_OUT;
  wire fpu_div_fState_S4$CLR,
       fpu_div_fState_S4$DEQ,
       fpu_div_fState_S4$EMPTY_N,
       fpu_div_fState_S4$ENQ,
       fpu_div_fState_S4$FULL_N;
  // ports of submodule fpu_madd_fOperand_S0
  wire [195 : 0] fpu_madd_fOperand_S0$D_IN, fpu_madd_fOperand_S0$D_OUT;
  wire fpu_madd_fOperand_S0$CLR,
       fpu_madd_fOperand_S0$DEQ,
       fpu_madd_fOperand_S0$EMPTY_N,
       fpu_madd_fOperand_S0$ENQ,
       fpu_madd_fOperand_S0$FULL_N;
  // ports of submodule fpu_madd_fProd_S2
  wire [105 : 0] fpu_madd_fProd_S2$D_IN, fpu_madd_fProd_S2$D_OUT;
  wire fpu_madd_fProd_S2$CLR,
       fpu_madd_fProd_S2$DEQ,
       fpu_madd_fProd_S2$EMPTY_N,
       fpu_madd_fProd_S2$ENQ,
       fpu_madd_fProd_S2$FULL_N;
  // ports of submodule fpu_madd_fProd_S3
  wire [105 : 0] fpu_madd_fProd_S3$D_IN, fpu_madd_fProd_S3$D_OUT;
  wire fpu_madd_fProd_S3$CLR,
       fpu_madd_fProd_S3$DEQ,
       fpu_madd_fProd_S3$EMPTY_N,
       fpu_madd_fProd_S3$ENQ,
       fpu_madd_fProd_S3$FULL_N;
  // ports of submodule fpu_madd_fResult_S9
  wire [68 : 0] fpu_madd_fResult_S9$D_IN, fpu_madd_fResult_S9$D_OUT;
  wire fpu_madd_fResult_S9$CLR,
       fpu_madd_fResult_S9$DEQ,
       fpu_madd_fResult_S9$EMPTY_N,
       fpu_madd_fResult_S9$ENQ,
       fpu_madd_fResult_S9$FULL_N;
  // ports of submodule fpu_madd_fState_S1
  wire [257 : 0] fpu_madd_fState_S1$D_IN, fpu_madd_fState_S1$D_OUT;
  wire fpu_madd_fState_S1$CLR,
       fpu_madd_fState_S1$DEQ,
       fpu_madd_fState_S1$EMPTY_N,
       fpu_madd_fState_S1$ENQ,
       fpu_madd_fState_S1$FULL_N;
  // ports of submodule fpu_madd_fState_S2
  wire [151 : 0] fpu_madd_fState_S2$D_IN, fpu_madd_fState_S2$D_OUT;
  wire fpu_madd_fState_S2$CLR,
       fpu_madd_fState_S2$DEQ,
       fpu_madd_fState_S2$EMPTY_N,
       fpu_madd_fState_S2$ENQ,
       fpu_madd_fState_S2$FULL_N;
  // ports of submodule fpu_madd_fState_S3
  wire [151 : 0] fpu_madd_fState_S3$D_IN, fpu_madd_fState_S3$D_OUT;
  wire fpu_madd_fState_S3$CLR,
       fpu_madd_fState_S3$DEQ,
       fpu_madd_fState_S3$EMPTY_N,
       fpu_madd_fState_S3$ENQ,
       fpu_madd_fState_S3$FULL_N;
  // ports of submodule fpu_madd_fState_S4
  wire [203 : 0] fpu_madd_fState_S4$D_IN, fpu_madd_fState_S4$D_OUT;
  wire fpu_madd_fState_S4$CLR,
       fpu_madd_fState_S4$DEQ,
       fpu_madd_fState_S4$EMPTY_N,
       fpu_madd_fState_S4$ENQ,
       fpu_madd_fState_S4$FULL_N;
  // ports of submodule fpu_madd_fState_S5
  wire [215 : 0] fpu_madd_fState_S5$D_IN, fpu_madd_fState_S5$D_OUT;
  wire fpu_madd_fState_S5$CLR,
       fpu_madd_fState_S5$DEQ,
       fpu_madd_fState_S5$EMPTY_N,
       fpu_madd_fState_S5$ENQ,
       fpu_madd_fState_S5$FULL_N;
  // ports of submodule fpu_madd_fState_S6
  wire [202 : 0] fpu_madd_fState_S6$D_IN, fpu_madd_fState_S6$D_OUT;
  wire fpu_madd_fState_S6$CLR,
       fpu_madd_fState_S6$DEQ,
       fpu_madd_fState_S6$EMPTY_N,
       fpu_madd_fState_S6$ENQ,
       fpu_madd_fState_S6$FULL_N;
  // ports of submodule fpu_madd_fState_S7
  wire [202 : 0] fpu_madd_fState_S7$D_IN, fpu_madd_fState_S7$D_OUT;
  wire fpu_madd_fState_S7$CLR,
       fpu_madd_fState_S7$DEQ,
       fpu_madd_fState_S7$EMPTY_N,
       fpu_madd_fState_S7$ENQ,
       fpu_madd_fState_S7$FULL_N;
  // ports of submodule fpu_madd_fState_S8
  wire [140 : 0] fpu_madd_fState_S8$D_IN, fpu_madd_fState_S8$D_OUT;
  wire fpu_madd_fState_S8$CLR,
       fpu_madd_fState_S8$DEQ,
       fpu_madd_fState_S8$EMPTY_N,
       fpu_madd_fState_S8$ENQ,
       fpu_madd_fState_S8$FULL_N;
  // ports of submodule fpu_sqr_fOperand_S0
  wire [66 : 0] fpu_sqr_fOperand_S0$D_IN, fpu_sqr_fOperand_S0$D_OUT;
  wire fpu_sqr_fOperand_S0$CLR,
       fpu_sqr_fOperand_S0$DEQ,
       fpu_sqr_fOperand_S0$EMPTY_N,
       fpu_sqr_fOperand_S0$ENQ,
       fpu_sqr_fOperand_S0$FULL_N;
  // ports of submodule fpu_sqr_fResult_S5
  wire [68 : 0] fpu_sqr_fResult_S5$D_IN, fpu_sqr_fResult_S5$D_OUT;
  wire fpu_sqr_fResult_S5$CLR,
       fpu_sqr_fResult_S5$DEQ,
       fpu_sqr_fResult_S5$EMPTY_N,
       fpu_sqr_fResult_S5$ENQ,
       fpu_sqr_fResult_S5$FULL_N;
  // ports of submodule fpu_sqr_fState_S1
  wire [194 : 0] fpu_sqr_fState_S1$D_IN, fpu_sqr_fState_S1$D_OUT;
  wire fpu_sqr_fState_S1$CLR,
       fpu_sqr_fState_S1$DEQ,
       fpu_sqr_fState_S1$EMPTY_N,
       fpu_sqr_fState_S1$ENQ,
       fpu_sqr_fState_S1$FULL_N;
  // ports of submodule fpu_sqr_fState_S2
  wire [136 : 0] fpu_sqr_fState_S2$D_IN, fpu_sqr_fState_S2$D_OUT;
  wire fpu_sqr_fState_S2$CLR,
       fpu_sqr_fState_S2$DEQ,
       fpu_sqr_fState_S2$EMPTY_N,
       fpu_sqr_fState_S2$ENQ,
       fpu_sqr_fState_S2$FULL_N;
  // ports of submodule fpu_sqr_fState_S3
  wire [195 : 0] fpu_sqr_fState_S3$D_IN, fpu_sqr_fState_S3$D_OUT;
  wire fpu_sqr_fState_S3$CLR,
       fpu_sqr_fState_S3$DEQ,
       fpu_sqr_fState_S3$EMPTY_N,
       fpu_sqr_fState_S3$ENQ,
       fpu_sqr_fState_S3$FULL_N;
  // ports of submodule fpu_sqr_fState_S4
  wire [138 : 0] fpu_sqr_fState_S4$D_IN, fpu_sqr_fState_S4$D_OUT;
  wire fpu_sqr_fState_S4$CLR,
       fpu_sqr_fState_S4$DEQ,
       fpu_sqr_fState_S4$EMPTY_N,
       fpu_sqr_fState_S4$ENQ,
       fpu_sqr_fState_S4$FULL_N;
  // ports of submodule iFifo
  wire [201 : 0] iFifo$D_IN, iFifo$D_OUT;
  wire iFifo$CLR, iFifo$DEQ, iFifo$EMPTY_N, iFifo$ENQ, iFifo$FULL_N;
  // ports of submodule isDoubleFifo
  wire isDoubleFifo$CLR,
       isDoubleFifo$DEQ,
       isDoubleFifo$D_IN,
       isDoubleFifo$D_OUT,
       isDoubleFifo$EMPTY_N,
       isDoubleFifo$ENQ,
       isDoubleFifo$FULL_N;
  // ports of submodule isNegateFifo
  wire isNegateFifo$CLR,
       isNegateFifo$DEQ,
       isNegateFifo$D_IN,
       isNegateFifo$D_OUT,
       isNegateFifo$EMPTY_N,
       isNegateFifo$ENQ,
       isNegateFifo$FULL_N;
  // ports of submodule oFifo
  wire [69 : 0] oFifo$D_IN, oFifo$D_OUT;
  wire oFifo$CLR, oFifo$DEQ, oFifo$EMPTY_N, oFifo$ENQ, oFifo$FULL_N;
  // ports of submodule resetReqsF
  wire resetReqsF$CLR,
       resetReqsF$DEQ,
       resetReqsF$EMPTY_N,
       resetReqsF$ENQ,
       resetReqsF$FULL_N;
  // ports of submodule resetRspsF
  wire resetRspsF$CLR,
       resetRspsF$DEQ,
       resetRspsF$EMPTY_N,
       resetRspsF$ENQ,
       resetRspsF$FULL_N;
  // ports of submodule rmdFifo
  wire [2 : 0] rmdFifo$D_IN, rmdFifo$D_OUT;
  wire rmdFifo$CLR, rmdFifo$DEQ, rmdFifo$EMPTY_N, rmdFifo$ENQ, rmdFifo$FULL_N;
  // rule scheduling signals
  wire CAN_FIRE_RL_fpu_div_s1_stage,
       CAN_FIRE_RL_fpu_div_s2_stage,
       CAN_FIRE_RL_fpu_div_s3_stage,
       CAN_FIRE_RL_fpu_div_s4_stage,
       CAN_FIRE_RL_fpu_div_s5_stage,
       CAN_FIRE_RL_fpu_madd_s1_stage,
       CAN_FIRE_RL_fpu_madd_s2_stage,
       CAN_FIRE_RL_fpu_madd_s3_stage,
       CAN_FIRE_RL_fpu_madd_s4_stage,
       CAN_FIRE_RL_fpu_madd_s5_stage,
       CAN_FIRE_RL_fpu_madd_s6_stage,
       CAN_FIRE_RL_fpu_madd_s7_stage,
       CAN_FIRE_RL_fpu_madd_s8_stage,
       CAN_FIRE_RL_fpu_madd_s9_stage,
       CAN_FIRE_RL_fpu_sqr_s1_stage,
       CAN_FIRE_RL_fpu_sqr_s2_stage,
       CAN_FIRE_RL_fpu_sqr_s3_stage,
       CAN_FIRE_RL_fpu_sqr_s4_stage,
       CAN_FIRE_RL_fpu_sqr_s5_stage,
       CAN_FIRE_RL_getResFromPipe,
       CAN_FIRE_RL_getResFromPipe_1,
       CAN_FIRE_RL_getResFromPipe_2,
       CAN_FIRE_RL_passResult,
       CAN_FIRE_RL_rl_reset,
       CAN_FIRE_RL_start_op,
       CAN_FIRE_RL_work,
       CAN_FIRE_RL_work_1,
       CAN_FIRE___me_check_22,
       CAN_FIRE_server_core_request_put,
       CAN_FIRE_server_core_response_get,
       CAN_FIRE_server_reset_request_put,
       CAN_FIRE_server_reset_response_get,
       WILL_FIRE_RL_fpu_div_s1_stage,
       WILL_FIRE_RL_fpu_div_s2_stage,
       WILL_FIRE_RL_fpu_div_s3_stage,
       WILL_FIRE_RL_fpu_div_s4_stage,
       WILL_FIRE_RL_fpu_div_s5_stage,
       WILL_FIRE_RL_fpu_madd_s1_stage,
       WILL_FIRE_RL_fpu_madd_s2_stage,
       WILL_FIRE_RL_fpu_madd_s3_stage,
       WILL_FIRE_RL_fpu_madd_s4_stage,
       WILL_FIRE_RL_fpu_madd_s5_stage,
       WILL_FIRE_RL_fpu_madd_s6_stage,
       WILL_FIRE_RL_fpu_madd_s7_stage,
       WILL_FIRE_RL_fpu_madd_s8_stage,
       WILL_FIRE_RL_fpu_madd_s9_stage,
       WILL_FIRE_RL_fpu_sqr_s1_stage,
       WILL_FIRE_RL_fpu_sqr_s2_stage,
       WILL_FIRE_RL_fpu_sqr_s3_stage,
       WILL_FIRE_RL_fpu_sqr_s4_stage,
       WILL_FIRE_RL_fpu_sqr_s5_stage,
       WILL_FIRE_RL_getResFromPipe,
       WILL_FIRE_RL_getResFromPipe_1,
       WILL_FIRE_RL_getResFromPipe_2,
       WILL_FIRE_RL_passResult,
       WILL_FIRE_RL_rl_reset,
       WILL_FIRE_RL_start_op,
       WILL_FIRE_RL_work,
       WILL_FIRE_RL_work_1,
       WILL_FIRE___me_check_22,
       WILL_FIRE_server_core_request_put,
       WILL_FIRE_server_core_response_get,
       WILL_FIRE_server_reset_request_put,
       WILL_FIRE_server_reset_response_get;
  // inputs to muxes for submodule ports
  wire [116 : 0] MUX_rg_res$write_1__VAL_2;
  wire [115 : 0] MUX_rg_b$write_1__VAL_1,
		 MUX_rg_b$write_1__VAL_2,
		 MUX_rg_r$write_1__VAL_1,
		 MUX_rg_r$write_1__VAL_2,
		 MUX_rg_r_1$write_1__VAL_2,
		 MUX_rg_s$write_1__VAL_1,
		 MUX_rg_s$write_1__VAL_2;
  wire [57 : 0] MUX_rg_d$write_1__VAL_1, MUX_rg_q$write_1__VAL_2;
  wire [5 : 0] MUX_rg_index$write_1__VAL_2, MUX_rg_index_1$write_1__VAL_2;
  wire MUX_crg_done$port1__write_1__SEL_1,
       MUX_crg_done_1$port1__write_1__SEL_1,
       MUX_crg_done_1$port1__write_1__SEL_2,
       MUX_rg_index$write_1__SEL_1;
  // remaining internal signals
  reg [63 : 0] CASE_fpu_div_fState_S4D_OUT_BITS_68_TO_66_0_C_ETC__q173,
	       CASE_fpu_sqr_fState_S4D_OUT_BITS_68_TO_66_0_C_ETC__q183,
	       CASE_iFifoD_OUT_BITS_3_TO_0_0_460718241880001_ETC__q177,
	       CASE_iFifoD_OUT_BITS_3_TO_0_0_IF_iFifo_first__ETC__q176,
	       IF_iFifo_first__087_BITS_3_TO_0_088_EQ_0_089_O_ETC___d4623;
  reg [62 : 0] CASE_fpu_div_fState_S3D_OUT_BITS_124_TO_122_0_ETC__q175,
	       CASE_fpu_div_fState_S4D_OUT_BITS_1_TO_0_0_0_0_ETC__q172,
	       CASE_fpu_div_fState_S4D_OUT_BITS_1_TO_0_0b0_f_ETC__q171,
	       CASE_fpu_div_fState_S4D_OUT_BITS_68_TO_66_2_I_ETC__q169,
	       CASE_fpu_madd_fState_S8D_OUT_BITS_2_TO_1_0b0__ETC__q130,
	       CASE_fpu_madd_fState_S8D_OUT_BITS_2_TO_1_0b0__ETC__q131,
	       CASE_fpu_madd_fState_S8D_OUT_BITS_70_TO_68_0__ETC__q132,
	       CASE_fpu_sqr_fState_S4D_OUT_BITS_1_TO_0_0_0_0_ETC__q182,
	       CASE_fpu_sqr_fState_S4D_OUT_BITS_1_TO_0_0b0_f_ETC__q181,
	       CASE_fpu_sqr_fState_S4D_OUT_BITS_68_TO_66_2_I_ETC__q179;
  reg [51 : 0] CASE_fpu_div_fState_S4D_OUT_BITS_1_TO_0_0b0_f_ETC__q1,
	       CASE_fpu_div_fState_S4D_OUT_BITS_1_TO_0_0b0_f_ETC__q2,
	       CASE_fpu_madd_fState_S8D_OUT_BITS_2_TO_1_0b0__ETC__q5,
	       CASE_fpu_madd_fState_S8D_OUT_BITS_2_TO_1_0b0__ETC__q6,
	       CASE_fpu_sqr_fState_S4D_OUT_BITS_1_TO_0_0b0_f_ETC__q3,
	       CASE_fpu_sqr_fState_S4D_OUT_BITS_1_TO_0_0b0_f_ETC__q4,
	       CASE_guard03260_0b0_sfdin11482_BITS_56_TO_5_0b_ETC__q110,
	       CASE_guard03260_0b0_sfdin11482_BITS_56_TO_5_0b_ETC__q111,
	       CASE_guard12299_0b0_theResult___snd20235_BITS__ETC__q112,
	       CASE_guard12299_0b0_theResult___snd20235_BITS__ETC__q113,
	       CASE_guard32950_0b0_theResult___snd40862_BITS__ETC__q75,
	       CASE_guard32950_0b0_theResult___snd40862_BITS__ETC__q76,
	       CASE_guard42199_0b0_sfdin50421_BITS_56_TO_5_0b_ETC__q77,
	       CASE_guard42199_0b0_sfdin50421_BITS_56_TO_5_0b_ETC__q78,
	       CASE_guard51238_0b0_theResult___snd59174_BITS__ETC__q81,
	       CASE_guard51238_0b0_theResult___snd59174_BITS__ETC__q82,
	       CASE_guard55373_0b0_theResult___snd63285_BITS__ETC__q48,
	       CASE_guard55373_0b0_theResult___snd63285_BITS__ETC__q49,
	       CASE_guard64622_0b0_sfdin72844_BITS_56_TO_5_0b_ETC__q50,
	       CASE_guard64622_0b0_sfdin72844_BITS_56_TO_5_0b_ETC__q51,
	       CASE_guard73661_0b0_theResult___snd81597_BITS__ETC__q52,
	       CASE_guard73661_0b0_theResult___snd81597_BITS__ETC__q53,
	       CASE_guard94011_0b0_theResult___snd01923_BITS__ETC__q108,
	       CASE_guard94011_0b0_theResult___snd01923_BITS__ETC__q109,
	       _theResult___fst_sfd__h142620,
	       _theResult___fst_sfd__h148290,
	       _theResult___fst_sfd__h164058,
	       _theResult___fst_sfd__h173648,
	       _theResult___fst_sfd__h182400,
	       _theResult___fst_sfd__h18519,
	       _theResult___fst_sfd__h186930,
	       _theResult___fst_sfd__h19008,
	       _theResult___fst_sfd__h202696,
	       _theResult___fst_sfd__h212286,
	       _theResult___fst_sfd__h221038,
	       _theResult___fst_sfd__h225869,
	       _theResult___fst_sfd__h241635,
	       _theResult___fst_sfd__h251225,
	       _theResult___fst_sfd__h259977,
	       _theResult___fst_sfd__h42605,
	       _theResult___fst_sfd__h95988;
  reg [22 : 0] CASE_guard69623_0b0_sfdin77716_BITS_56_TO_34_0_ETC__q162,
	       CASE_guard69623_0b0_sfdin77716_BITS_56_TO_34_0_ETC__q163,
	       CASE_guard78330_0b0_theResult___snd86329_BITS__ETC__q160,
	       CASE_guard78330_0b0_theResult___snd86329_BITS__ETC__q161,
	       CASE_guard87260_0b0_sfdin95482_BITS_56_TO_34_0_ETC__q164,
	       CASE_guard87260_0b0_sfdin95482_BITS_56_TO_34_0_ETC__q165,
	       CASE_guard96096_0b0_theResult___snd04119_BITS__ETC__q166,
	       CASE_guard96096_0b0_theResult___snd04119_BITS__ETC__q167,
	       _theResult___fst_sfd__h269596,
	       _theResult___fst_sfd__h278317,
	       _theResult___fst_sfd__h286899,
	       _theResult___fst_sfd__h296083,
	       _theResult___fst_sfd__h304719;
  reg [10 : 0] CASE_fpu_div_fState_S4D_OUT_BITS_1_TO_0_0b0_f_ETC__q14,
	       CASE_fpu_div_fState_S4D_OUT_BITS_1_TO_0_0b0_f_ETC__q15,
	       CASE_fpu_madd_fState_S8D_OUT_BITS_2_TO_1_0b0__ETC__q31,
	       CASE_fpu_madd_fState_S8D_OUT_BITS_2_TO_1_0b0__ETC__q32,
	       CASE_fpu_sqr_fState_S4D_OUT_BITS_1_TO_0_0b0_f_ETC__q21,
	       CASE_fpu_sqr_fState_S4D_OUT_BITS_1_TO_0_0b0_f_ETC__q22,
	       CASE_guard03260_0b0_theResult___fst_exp11488_0_ETC__q104,
	       CASE_guard03260_0b0_theResult___fst_exp11488_0_ETC__q105,
	       CASE_guard12299_0b0_theResult___fst_exp20289_0_ETC__q106,
	       CASE_guard12299_0b0_theResult___fst_exp20289_0_ETC__q107,
	       CASE_guard32950_0b0_theResult___fst_exp40911_0_ETC__q69,
	       CASE_guard32950_0b0_theResult___fst_exp40911_0_ETC__q70,
	       CASE_guard42199_0b0_theResult___fst_exp50427_0_ETC__q71,
	       CASE_guard42199_0b0_theResult___fst_exp50427_0_ETC__q72,
	       CASE_guard51238_0b0_theResult___fst_exp59228_0_ETC__q73,
	       CASE_guard51238_0b0_theResult___fst_exp59228_0_ETC__q74,
	       CASE_guard55373_0b0_theResult___fst_exp63334_0_ETC__q42,
	       CASE_guard55373_0b0_theResult___fst_exp63334_0_ETC__q43,
	       CASE_guard64622_0b0_theResult___fst_exp72850_0_ETC__q44,
	       CASE_guard64622_0b0_theResult___fst_exp72850_0_ETC__q45,
	       CASE_guard73661_0b0_theResult___fst_exp81651_0_ETC__q46,
	       CASE_guard73661_0b0_theResult___fst_exp81651_0_ETC__q47,
	       CASE_guard94011_0b0_theResult___fst_exp01972_0_ETC__q102,
	       CASE_guard94011_0b0_theResult___fst_exp01972_0_ETC__q103,
	       _theResult___fst_exp__h142619,
	       _theResult___fst_exp__h148289,
	       _theResult___fst_exp__h164057,
	       _theResult___fst_exp__h173647,
	       _theResult___fst_exp__h182399,
	       _theResult___fst_exp__h18518,
	       _theResult___fst_exp__h186929,
	       _theResult___fst_exp__h202695,
	       _theResult___fst_exp__h212285,
	       _theResult___fst_exp__h221037,
	       _theResult___fst_exp__h225868,
	       _theResult___fst_exp__h241634,
	       _theResult___fst_exp__h251224,
	       _theResult___fst_exp__h259976,
	       _theResult___fst_exp__h42604,
	       _theResult___fst_exp__h95987;
  reg [7 : 0] CASE_guard69623_0b0_theResult___fst_exp77722_0_ETC__q154,
	      CASE_guard69623_0b0_theResult___fst_exp77722_0_ETC__q155,
	      CASE_guard78330_0b0_theResult___fst_exp86378_0_ETC__q152,
	      CASE_guard78330_0b0_theResult___fst_exp86378_0_ETC__q153,
	      CASE_guard87260_0b0_theResult___fst_exp95488_0_ETC__q156,
	      CASE_guard87260_0b0_theResult___fst_exp95488_0_ETC__q157,
	      CASE_guard96096_0b0_theResult___fst_exp04173_0_ETC__q158,
	      CASE_guard96096_0b0_theResult___fst_exp04173_0_ETC__q159,
	      _theResult___fst_exp__h269595,
	      _theResult___fst_exp__h278316,
	      _theResult___fst_exp__h286898,
	      _theResult___fst_exp__h296082,
	      _theResult___fst_exp__h304718;
  reg CASE_fpu_div_fOperands_S0D_OUT_BITS_2_TO_0_0__ETC__q9,
      CASE_fpu_div_fState_S3D_OUT_BITS_124_TO_122_0_ETC__q174,
      CASE_fpu_div_fState_S4D_OUT_BITS_1_TO_0_0b0_f_ETC__q170,
      CASE_fpu_div_fState_S4D_OUT_BITS_68_TO_66_2_f_ETC__q168,
      CASE_fpu_madd_fState_S8D_OUT_BITS_2_TO_1_0b0__ETC__q126,
      CASE_fpu_madd_fState_S8D_OUT_BITS_70_TO_68_0__ETC__q127,
      CASE_fpu_sqr_fState_S4D_OUT_BITS_1_TO_0_0b0_f_ETC__q180,
      CASE_fpu_sqr_fState_S4D_OUT_BITS_68_TO_66_2_f_ETC__q178,
      CASE_guard03260_0b0_NOT_iFifoD_OUT_BIT_103_0b_ETC__q122,
      CASE_guard03260_0b0_iFifoD_OUT_BIT_103_0b1_iF_ETC__q116,
      CASE_guard12299_0b0_NOT_iFifoD_OUT_BIT_103_0b_ETC__q124,
      CASE_guard12299_0b0_iFifoD_OUT_BIT_103_0b1_iF_ETC__q118,
      CASE_guard32950_0b0_NOT_iFifoD_OUT_BIT_38_0b1_ETC__q87,
      CASE_guard32950_0b0_iFifoD_OUT_BIT_38_0b1_iFi_ETC__q79,
      CASE_guard42199_0b0_NOT_iFifoD_OUT_BIT_38_0b1_ETC__q89,
      CASE_guard42199_0b0_iFifoD_OUT_BIT_38_0b1_iFi_ETC__q83,
      CASE_guard51238_0b0_NOT_iFifoD_OUT_BIT_38_0b1_ETC__q91,
      CASE_guard51238_0b0_iFifoD_OUT_BIT_38_0b1_iFi_ETC__q85,
      CASE_guard55373_0b0_iFifoD_OUT_BIT_168_0b1_iF_ETC__q54,
      CASE_guard64622_0b0_iFifoD_OUT_BIT_168_0b1_iF_ETC__q56,
      CASE_guard69623_0b0_NOT_resWirewget_BIT_68_0b_ETC__q145,
      CASE_guard69623_0b0_resWirewget_BIT_68_0b1_re_ETC__q144,
      CASE_guard73661_0b0_iFifoD_OUT_BIT_168_0b1_iF_ETC__q58,
      CASE_guard78330_0b0_NOT_resWirewget_BIT_68_0b_ETC__q147,
      CASE_guard78330_0b0_resWirewget_BIT_68_0b1_re_ETC__q146,
      CASE_guard87260_0b0_NOT_resWirewget_BIT_68_0b_ETC__q149,
      CASE_guard87260_0b0_resWirewget_BIT_68_0b1_re_ETC__q148,
      CASE_guard94011_0b0_NOT_iFifoD_OUT_BIT_103_0b_ETC__q120,
      CASE_guard94011_0b0_iFifoD_OUT_BIT_103_0b1_iF_ETC__q114,
      CASE_guard96096_0b0_NOT_resWirewget_BIT_68_0b_ETC__q151,
      CASE_guard96096_0b0_resWirewget_BIT_68_0b1_re_ETC__q150,
      CASE_iFifoD_OUT_BITS_6_TO_4_0_CASE_guard03260_ETC__q117,
      CASE_iFifoD_OUT_BITS_6_TO_4_0_CASE_guard03260_ETC__q123,
      CASE_iFifoD_OUT_BITS_6_TO_4_0_CASE_guard12299_ETC__q119,
      CASE_iFifoD_OUT_BITS_6_TO_4_0_CASE_guard12299_ETC__q125,
      CASE_iFifoD_OUT_BITS_6_TO_4_0_CASE_guard32950_ETC__q80,
      CASE_iFifoD_OUT_BITS_6_TO_4_0_CASE_guard32950_ETC__q88,
      CASE_iFifoD_OUT_BITS_6_TO_4_0_CASE_guard42199_ETC__q84,
      CASE_iFifoD_OUT_BITS_6_TO_4_0_CASE_guard42199_ETC__q90,
      CASE_iFifoD_OUT_BITS_6_TO_4_0_CASE_guard51238_ETC__q86,
      CASE_iFifoD_OUT_BITS_6_TO_4_0_CASE_guard51238_ETC__q92,
      CASE_iFifoD_OUT_BITS_6_TO_4_0_CASE_guard55373_ETC__q55,
      CASE_iFifoD_OUT_BITS_6_TO_4_0_CASE_guard64622_ETC__q57,
      CASE_iFifoD_OUT_BITS_6_TO_4_0_CASE_guard73661_ETC__q59,
      CASE_iFifoD_OUT_BITS_6_TO_4_0_CASE_guard94011_ETC__q115,
      CASE_iFifoD_OUT_BITS_6_TO_4_0_CASE_guard94011_ETC__q121,
      IF_iFifo_first__087_BITS_3_TO_0_088_EQ_0_089_O_ETC___d3110,
      IF_iFifo_first__087_BITS_6_TO_4_118_EQ_0_191_O_ETC___d3320,
      IF_iFifo_first__087_BITS_6_TO_4_118_EQ_0_191_O_ETC___d4028,
      IF_iFifo_first__087_BITS_6_TO_4_118_EQ_0_191_O_ETC___d4582,
      IF_iFifo_first__087_BITS_6_TO_4_118_EQ_0_191_O_ETC___d4803,
      IF_iFifo_first__087_BITS_6_TO_4_118_EQ_0_191_O_ETC___d5348,
      IF_rmdFifo_first__778_EQ_0_779_OR_rmdFifo_firs_ETC___d6028,
      IF_rmdFifo_first__778_EQ_0_779_OR_rmdFifo_firs_ETC___d6400,
      IF_rmdFifo_first__778_EQ_0_779_THEN_IF_IF_IF_I_ETC___d5823,
      IF_rmdFifo_first__778_EQ_0_779_THEN_IF_IF_IF_I_ETC___d6324,
      IF_rmdFifo_first__778_EQ_0_779_THEN_IF_IF_IF_I_ETC___d6388,
      IF_rmdFifo_first__778_EQ_0_779_THEN_IF_IF_IF_I_ETC___d6409,
      IF_rmdFifo_first__778_EQ_0_779_THEN_IF_IF_IF_r_ETC___d6023,
      IF_rmdFifo_first__778_EQ_0_779_THEN_IF_IF_IF_r_ETC___d6373,
      IF_rmdFifo_first__778_EQ_0_779_THEN_IF_IF_IF_r_ETC___d6397,
      IF_rmdFifo_first__778_EQ_0_779_THEN_IF_IF_IF_r_ETC___d6418;
  wire [194 : 0] IF_fpu_sqr_fOperand_S0_first__059_BITS_65_TO_5_ETC___d1212;
  wire [139 : 0] IF_NOT_fpu_madd_fState_S4_first__547_BIT_130_5_ETC___d2595;
  wire [118 : 0] IF_fpu_madd_fOperand_S0_first__803_BITS_129_TO_ETC___d1959;
  wire [115 : 0] IF_IF_rg_index_1_87_ULE_58_91_THEN_NOT_rg_b_92_ETC___d1028,
		 IF_rg_index_1_87_ULE_58_91_THEN_IF_rg_res_94_B_ETC___d1002,
		 IF_rg_index_1_87_ULE_58_91_THEN_IF_rg_res_94_B_ETC___d1022,
		 IF_rg_index_1_87_ULE_58_91_THEN_IF_rg_res_94_B_ETC___d1026,
		 IF_rg_index_1_87_ULE_58_91_THEN_IF_rg_res_94_B_ETC___d1036,
		 IF_rg_index_ULE_57_THEN_IF_rg_r_0_BIT_115_1_TH_ETC___d22,
		 IF_rg_res_94_BIT_116_95_THEN_rg_res_94_BITS_11_ETC___d1025,
		 _theResult___fst__h43498,
		 _theResult___fst__h43537,
		 _theResult___fst__h43622,
		 _theResult___snd_fst__h43500,
		 _theResult___snd_fst__h43539,
		 _theResult___snd_fst__h43624,
		 _theResult___snd_snd__h43671,
		 _theResult___snd_snd__h43737,
		 _theResult___snd_snd_snd__h43503,
		 _theResult___snd_snd_snd__h43542,
		 _theResult___snd_snd_snd__h43627,
		 b___1__h77160,
		 b__h31634,
		 b__h43630,
		 b__h43734,
		 r__h43681,
		 r__h43685,
		 r__h43746,
		 r__h43775,
		 s__h43680,
		 s__h43745,
		 sum__h43628,
		 sum__h43732,
		 value__h31592,
		 x__h85931;
  wire [113 : 0] x__h30477;
  wire [105 : 0] IF_0_CONCAT_IF_IF_7170_MINUS_fpu_madd_fState_S_ETC__q24,
		 _theResult___fst__h116827,
		 _theResult___snd__h130966,
		 _theResult___snd__h130980,
		 _theResult___snd__h130982,
		 _theResult___snd__h130994,
		 _theResult___snd__h131000,
		 _theResult___snd__h131018,
		 _theResult___snd__h131023,
		 fpu_madd_fProd_S3_first__009_SRL_IF_7170_MINUS_ETC___d2012,
		 sfdBC__h115662,
		 sfdin__h130943,
		 x__h116896;
  wire [68 : 0] IF_fpu_madd_fState_S8_first__960_BIT_67_963_AN_ETC___d3081;
  wire [63 : 0] IF_IF_fpu_madd_fOperand_S0_first__803_BIT_195__ETC___d1936,
		IF_IF_fpu_madd_fOperand_S0_first__803_BIT_195__ETC___d1939,
		IF_fpu_div_fOperands_S0_first__6_BITS_65_TO_55_ETC___d385,
		IF_fpu_madd_fOperand_S0_first__803_BITS_129_TO_ETC___d1938,
		IF_iFifo_first__087_BITS_102_TO_95_625_EQ_255__ETC___d5328,
		IF_iFifo_first__087_BITS_102_TO_95_625_EQ_255__ETC___d5378,
		IF_iFifo_first__087_BITS_167_TO_160_130_EQ_255_ETC___d3846,
		IF_iFifo_first__087_BITS_37_TO_30_850_EQ_255_8_ETC___d4553,
		IF_iFifo_first__087_BITS_37_TO_30_850_EQ_255_8_ETC___d4612,
		IF_iFifo_first__087_BIT_136_624_THEN_IF_iFifo__ETC___d5330,
		IF_iFifo_first__087_BIT_201_115_THEN_IF_iFifo__ETC___d3848,
		IF_iFifo_first__087_BIT_71_849_THEN_IF_iFifo_f_ETC___d4555,
		IF_iFifo_first__087_BIT_71_849_THEN_IF_iFifo_f_ETC___d4618,
		IF_isDoubleFifo_first__407_THEN_IF_isNegateFif_ETC___d6657,
		NOT_fpu_div_fOperands_S0_first__6_BITS_129_TO__ETC___d382,
		fpu_div_fState_S3_first__16_BIT_121_37_CONCAT__ETC___d866;
  wire [62 : 0] IF_0b0_CONCAT_NOT_fpu_div_fState_S4_first__73__ETC___d910,
		IF_0b0_CONCAT_NOT_fpu_madd_fState_S8_first__96_ETC___d3065,
		IF_0b0_CONCAT_NOT_fpu_sqr_fState_S4_first__687_ETC___d1724,
		IF_IF_7170_MINUS_fpu_madd_fState_S3_first__995_ETC___d2534,
		IF_IF_fpu_div_fState_S3_first__16_BITS_120_TO__ETC___d859,
		IF_IF_fpu_madd_fOperand_S0_first__803_BIT_195__ETC___d1931,
		IF_IF_fpu_madd_fState_S7_first__651_BIT_128_65_ETC___d2952,
		IF_fpu_madd_fOperand_S0_first__803_BITS_129_TO_ETC___d1932,
		IF_fpu_madd_fOperand_S0_first__803_BIT_195_804_ETC___d1911,
		IF_fpu_madd_fState_S3_first__995_BITS_12_TO_0__ETC___d2536,
		IF_fpu_sqr_fState_S3_first__375_BIT_58_384_AND_ETC___d1678,
		IF_iFifo_first__087_BITS_102_TO_95_625_EQ_255__ETC___d5327,
		IF_iFifo_first__087_BITS_37_TO_30_850_EQ_255_8_ETC___d4552;
  wire [58 : 0] IF_0_CONCAT_IF_fpu_sqr_fState_S3_first__375_BI_ETC__q19,
		_theResult___snd__h94767,
		_theResult___snd__h94782,
		_theResult___snd__h94784,
		_theResult___snd__h94797,
		_theResult___snd__h94803,
		_theResult___snd__h94821,
		_theResult___snd__h94826,
		result__h85925,
		sfdin__h94744,
		x__h86149;
  wire [57 : 0] IF_0_CONCAT_IF_IF_fpu_div_fState_S3_first__16__ETC__q12,
		IF_rg_index_ULE_57_THEN_rg_q_BITS_56_TO_0_CONC_ETC___d14,
		IF_rg_r_BIT_115_THEN_rg_q_PLUS_NEG_INV_rg_q_89_ETC__q10,
		_theResult____h31574,
		_theResult___snd__h33766,
		_theResult___snd__h41401,
		_theResult___snd__h41416,
		_theResult___snd__h41418,
		_theResult___snd__h41431,
		_theResult___snd__h41437,
		_theResult___snd__h41455,
		_theResult___snd__h41460,
		_theResult___snd_snd_snd__h33014,
		result__h31668,
		result__h31699,
		result__h31874,
		rg_q_PLUS_NEG_INV_rg_q_89_90___d491,
		sfd___1__h60702,
		sfd__h44951,
		sfd__h44953,
		sfdin__h33169,
		sfdin__h41378,
		x__h31813,
		x__h32103,
		x__h60693;
  wire [56 : 0] IF_0_CONCAT_IF_IF_0b0_CONCAT_NOT_resWire_wget__ETC__q133,
		IF_0_CONCAT_IF_IF_3074_MINUS_SEXT_iFifo_first__ETC__q37,
		IF_0_CONCAT_IF_IF_3074_MINUS_SEXT_iFifo_first__ETC__q64,
		IF_0_CONCAT_IF_IF_3074_MINUS_SEXT_iFifo_first__ETC__q97,
		IF_0_CONCAT_IF_IF_3970_MINUS_SEXT_resWire_wget_ETC__q139,
		IF_0_CONCAT_IF_IF_fpu_madd_fState_S7_first__65_ETC__q29,
		IF_0_CONCAT_IF_iFifo_first__087_BITS_102_TO_95_ETC__q100,
		IF_0_CONCAT_IF_iFifo_first__087_BITS_102_TO_95_ETC__q93,
		IF_0_CONCAT_IF_iFifo_first__087_BITS_167_TO_16_ETC__q33,
		IF_0_CONCAT_IF_iFifo_first__087_BITS_167_TO_16_ETC__q40,
		IF_0_CONCAT_IF_iFifo_first__087_BITS_37_TO_30__ETC__q60,
		IF_0_CONCAT_IF_iFifo_first__087_BITS_37_TO_30__ETC__q67,
		IF_0_CONCAT_IF_resWire_wget__410_BITS_67_TO_57_ETC__q135,
		IF_0_CONCAT_IF_resWire_wget__410_BITS_67_TO_57_ETC__q142,
		_0b0_CONCAT_NOT_iFifo_first__087_BITS_102_TO_95_ETC___d4813,
		_0b0_CONCAT_NOT_iFifo_first__087_BITS_167_TO_16_ETC___d3330,
		_0b0_CONCAT_NOT_iFifo_first__087_BITS_37_TO_30__ETC___d4038,
		_0b0_CONCAT_NOT_resWire_wget__410_BITS_67_TO_57_ETC___d6038,
		_theResult____h164612,
		_theResult____h203250,
		_theResult____h242189,
		_theResult____h269613,
		_theResult____h287250,
		_theResult___snd__h141392,
		_theResult___snd__h141406,
		_theResult___snd__h141408,
		_theResult___snd__h141420,
		_theResult___snd__h141426,
		_theResult___snd__h141444,
		_theResult___snd__h141449,
		_theResult___snd__h163285,
		_theResult___snd__h163287,
		_theResult___snd__h163294,
		_theResult___snd__h163300,
		_theResult___snd__h163323,
		_theResult___snd__h172861,
		_theResult___snd__h172872,
		_theResult___snd__h172874,
		_theResult___snd__h172884,
		_theResult___snd__h172890,
		_theResult___snd__h172913,
		_theResult___snd__h181597,
		_theResult___snd__h181611,
		_theResult___snd__h181617,
		_theResult___snd__h181635,
		_theResult___snd__h201923,
		_theResult___snd__h201925,
		_theResult___snd__h201932,
		_theResult___snd__h201938,
		_theResult___snd__h201961,
		_theResult___snd__h211499,
		_theResult___snd__h211510,
		_theResult___snd__h211512,
		_theResult___snd__h211522,
		_theResult___snd__h211528,
		_theResult___snd__h211551,
		_theResult___snd__h220235,
		_theResult___snd__h220249,
		_theResult___snd__h220255,
		_theResult___snd__h220273,
		_theResult___snd__h240862,
		_theResult___snd__h240864,
		_theResult___snd__h240871,
		_theResult___snd__h240877,
		_theResult___snd__h240900,
		_theResult___snd__h250438,
		_theResult___snd__h250449,
		_theResult___snd__h250451,
		_theResult___snd__h250461,
		_theResult___snd__h250467,
		_theResult___snd__h250490,
		_theResult___snd__h259174,
		_theResult___snd__h259188,
		_theResult___snd__h259194,
		_theResult___snd__h259212,
		_theResult___snd__h277733,
		_theResult___snd__h277744,
		_theResult___snd__h277746,
		_theResult___snd__h277756,
		_theResult___snd__h277762,
		_theResult___snd__h277785,
		_theResult___snd__h286329,
		_theResult___snd__h286331,
		_theResult___snd__h286338,
		_theResult___snd__h286344,
		_theResult___snd__h286367,
		_theResult___snd__h295499,
		_theResult___snd__h295510,
		_theResult___snd__h295512,
		_theResult___snd__h295522,
		_theResult___snd__h295528,
		_theResult___snd__h295551,
		_theResult___snd__h304119,
		_theResult___snd__h304133,
		_theResult___snd__h304139,
		_theResult___snd__h304157,
		fpu_madd_fState_S5_first__601_BITS_56_TO_0_610_ETC___d2615,
		guard__h132367,
		result__h132372,
		result__h165225,
		result__h203863,
		result__h242802,
		result__h287863,
		sfdA__h131577,
		sfdBC__h131578,
		sfd__h133119,
		sfd__h144534,
		sfd__h183174,
		sfd__h222113,
		sfd__h262011,
		sfdin__h141369,
		sfdin__h172844,
		sfdin__h211482,
		sfdin__h250421,
		sfdin__h277716,
		sfdin__h295482,
		value__h31712,
		x__h131940,
		x__h131944,
		x__h132359,
		x__h132871,
		x__h132880,
		x__h165322,
		x__h203960,
		x__h242899,
		x__h287960,
		x__h30538;
  wire [53 : 0] sfd__h142040,
		sfd__h163352,
		sfd__h172942,
		sfd__h181670,
		sfd__h201990,
		sfd__h211580,
		sfd__h220308,
		sfd__h240929,
		sfd__h250519,
		sfd__h259247,
		sfd__h42033,
		sfd__h95416,
		value__h270233,
		value__h30480,
		value__h53174;
  wire [52 : 0] sfdA__h1086,
		sfdA__h1090,
		sfdB__h1087,
		sfdB__h1092,
		x__h114243,
		x__h114255;
  wire [51 : 0] IF_IF_IF_IF_3074_MINUS_SEXT_iFifo_first__087_B_ETC___d3813,
		IF_IF_IF_IF_3074_MINUS_SEXT_iFifo_first__087_B_ETC___d3815,
		IF_IF_IF_IF_3074_MINUS_SEXT_iFifo_first__087_B_ETC___d4519,
		IF_IF_IF_IF_3074_MINUS_SEXT_iFifo_first__087_B_ETC___d4521,
		IF_IF_IF_IF_3074_MINUS_SEXT_iFifo_first__087_B_ETC___d5294,
		IF_IF_IF_IF_3074_MINUS_SEXT_iFifo_first__087_B_ETC___d5296,
		IF_IF_IF_iFifo_first__087_BITS_102_TO_95_625_E_ETC___d5268,
		IF_IF_IF_iFifo_first__087_BITS_102_TO_95_625_E_ETC___d5270,
		IF_IF_IF_iFifo_first__087_BITS_102_TO_95_625_E_ETC___d5313,
		IF_IF_IF_iFifo_first__087_BITS_102_TO_95_625_E_ETC___d5315,
		IF_IF_IF_iFifo_first__087_BITS_167_TO_160_130__ETC___d3786,
		IF_IF_IF_iFifo_first__087_BITS_167_TO_160_130__ETC___d3788,
		IF_IF_IF_iFifo_first__087_BITS_167_TO_160_130__ETC___d3832,
		IF_IF_IF_iFifo_first__087_BITS_167_TO_160_130__ETC___d3834,
		IF_IF_IF_iFifo_first__087_BITS_37_TO_30_850_EQ_ETC___d4493,
		IF_IF_IF_iFifo_first__087_BITS_37_TO_30_850_EQ_ETC___d4495,
		IF_IF_IF_iFifo_first__087_BITS_37_TO_30_850_EQ_ETC___d4538,
		IF_IF_IF_iFifo_first__087_BITS_37_TO_30_850_EQ_ETC___d4540,
		IF_fpu_div_fOperands_S0_first__6_BITS_65_TO_55_ETC___d380,
		_theResult___fst_sfd__h164061,
		_theResult___fst_sfd__h173651,
		_theResult___fst_sfd__h182403,
		_theResult___fst_sfd__h182412,
		_theResult___fst_sfd__h182418,
		_theResult___fst_sfd__h202699,
		_theResult___fst_sfd__h212289,
		_theResult___fst_sfd__h221041,
		_theResult___fst_sfd__h221050,
		_theResult___fst_sfd__h221056,
		_theResult___fst_sfd__h241638,
		_theResult___fst_sfd__h251228,
		_theResult___fst_sfd__h259980,
		_theResult___fst_sfd__h259989,
		_theResult___fst_sfd__h259995,
		_theResult___fst_sfd__h42608,
		_theResult___fst_sfd__h95991,
		_theResult___fst_sfd__h96608,
		_theResult___sfd__h142542,
		_theResult___sfd__h163980,
		_theResult___sfd__h173570,
		_theResult___sfd__h182322,
		_theResult___sfd__h202618,
		_theResult___sfd__h212208,
		_theResult___sfd__h220960,
		_theResult___sfd__h241557,
		_theResult___sfd__h251147,
		_theResult___sfd__h259899,
		_theResult___sfd__h42527,
		_theResult___sfd__h95910,
		_theResult___snd_fst_sfd__h144484,
		_theResult___snd_fst_sfd__h164064,
		_theResult___snd_fst_sfd__h182406,
		_theResult___snd_fst_sfd__h183124,
		_theResult___snd_fst_sfd__h202702,
		_theResult___snd_fst_sfd__h221044,
		_theResult___snd_fst_sfd__h222063,
		_theResult___snd_fst_sfd__h241641,
		_theResult___snd_fst_sfd__h259983,
		_theResult___snd_fst_sfd__h30413,
		out___1_sfd__h144233,
		out___1_sfd__h182873,
		out___1_sfd__h221812,
		out_sfd__h142545,
		out_sfd__h163983,
		out_sfd__h173573,
		out_sfd__h182325,
		out_sfd__h202621,
		out_sfd__h212211,
		out_sfd__h220963,
		out_sfd__h241560,
		out_sfd__h251150,
		out_sfd__h259902,
		out_sfd__h42530,
		out_sfd__h95913,
		sfd__h17985,
		sfd__h17988,
		sfd__h45004,
		sfd__h99402,
		sfd__h99405,
		sfd__h99408;
  wire [24 : 0] sfd__h277814,
		sfd__h286396,
		sfd__h295580,
		sfd__h304192,
		value__h148921,
		value__h187559,
		value__h226498;
  wire [22 : 0] IF_IF_IF_IF_0b0_CONCAT_NOT_resWire_wget__410_B_ETC___d6576,
		IF_IF_IF_IF_0b0_CONCAT_NOT_resWire_wget__410_B_ETC___d6578,
		IF_IF_IF_IF_3970_MINUS_SEXT_resWire_wget__410__ETC___d6622,
		IF_IF_IF_IF_3970_MINUS_SEXT_resWire_wget__410__ETC___d6624,
		IF_IF_IF_resWire_wget__410_BITS_67_TO_57_416_E_ETC___d6595,
		IF_IF_IF_resWire_wget__410_BITS_67_TO_57_416_E_ETC___d6597,
		IF_IF_IF_resWire_wget__410_BITS_67_TO_57_416_E_ETC___d6641,
		IF_IF_IF_resWire_wget__410_BITS_67_TO_57_416_E_ETC___d6643,
		_theResult___fst_sfd__h278320,
		_theResult___fst_sfd__h286902,
		_theResult___fst_sfd__h296086,
		_theResult___fst_sfd__h304722,
		_theResult___fst_sfd__h304731,
		_theResult___fst_sfd__h304737,
		_theResult___sfd__h278239,
		_theResult___sfd__h286821,
		_theResult___sfd__h296005,
		_theResult___sfd__h304641,
		_theResult___snd_fst_sfd__h261961,
		_theResult___snd_fst_sfd__h286905,
		_theResult___snd_fst_sfd__h304725,
		out_sfd__h278242,
		out_sfd__h286824,
		out_sfd__h296008,
		out_sfd__h304644,
		sfd__h304743;
  wire [12 : 0] IF_fpu_div_fOperands_S0_first__6_BITS_129_TO_1_ETC___d282,
		IF_fpu_madd_fState_S4_first__547_BITS_128_TO_1_ETC___d2568,
		IF_fpu_madd_fState_S4_first__547_BITS_64_TO_54_ETC___d2563,
		IF_fpu_sqr_fOperand_S0_first__059_BITS_65_TO_5_ETC___d1195,
		_7170_MINUS_fpu_madd_fState_S3_first__995_BITS__ETC___d2007,
		value__h130883,
		value__h141307,
		value__h30425,
		value__h30601,
		x__h116929,
		x__h132471,
		x__h52551,
		x__h52569;
  wire [11 : 0] IF_IF_7170_MINUS_fpu_madd_fState_S3_first__995_ETC___d2031,
		IF_IF_7170_MINUS_fpu_madd_fState_S3_first__995_ETC___d2462,
		IF_IF_fpu_div_fState_S3_first__16_BITS_120_TO__ETC___d573,
		IF_IF_fpu_div_fState_S3_first__16_BITS_120_TO__ETC___d812,
		IF_SEXT_iFifo_first__087_BITS_102_TO_95_625_MI_ETC___d5106,
		IF_SEXT_iFifo_first__087_BITS_167_TO_160_130_M_ETC___d3623,
		IF_SEXT_iFifo_first__087_BITS_37_TO_30_850_MIN_ETC___d4331,
		IF_fpu_madd_fState_S7_first__651_BITS_126_TO_1_ETC___d2668,
		IF_fpu_madd_fState_S7_first__651_BITS_126_TO_1_ETC___d2903,
		IF_fpu_sqr_fOperand_S0_first__059_BITS_65_TO_5_ETC__q17,
		IF_fpu_sqr_fState_S3_first__375_BITS_121_TO_11_ETC___d1389,
		IF_fpu_sqr_fState_S3_first__375_BITS_121_TO_11_ETC___d1632,
		SEXT_iFifo_first__087_BITS_102_TO_95_625_MINUS_ETC___d4806,
		SEXT_iFifo_first__087_BITS_102_TO_95_625_MINUS_ETC__q96,
		SEXT_iFifo_first__087_BITS_167_TO_160_130_MINU_ETC___d3323,
		SEXT_iFifo_first__087_BITS_167_TO_160_130_MINU_ETC__q36,
		SEXT_iFifo_first__087_BITS_37_TO_30_850_MINUS__ETC___d4031,
		SEXT_iFifo_first__087_BITS_37_TO_30_850_MINUS__ETC__q63,
		SEXT_resWire_wget__410_BITS_67_TO_57_416_MINUS_ETC___d6031,
		SEXT_resWire_wget__410_BITS_67_TO_57_416_MINUS_ETC__q138,
		_3074_MINUS_0_CONCAT_IF_resWire_wget__410_BIT_5_ETC___d5531,
		_3074_MINUS_SEXT_iFifo_first__087_BITS_102_TO_9_ETC___d4809,
		_3074_MINUS_SEXT_iFifo_first__087_BITS_167_TO_1_ETC___d3326,
		_3074_MINUS_SEXT_iFifo_first__087_BITS_37_TO_30_ETC___d4034,
		_3970_MINUS_0_CONCAT_IF_iFifo_first__087_BIT_15_ETC___d3188,
		_3970_MINUS_0_CONCAT_IF_iFifo_first__087_BIT_29_ETC___d3908,
		_3970_MINUS_0_CONCAT_IF_iFifo_first__087_BIT_94_ETC___d4683,
		_3970_MINUS_SEXT_resWire_wget__410_BITS_67_TO_5_ETC___d6034,
		x__h165355,
		x__h203993,
		x__h242932,
		x__h287993;
  wire [10 : 0] IF_IF_IF_IF_3074_MINUS_SEXT_iFifo_first__087_B_ETC___d3729,
		IF_IF_IF_IF_3074_MINUS_SEXT_iFifo_first__087_B_ETC___d3731,
		IF_IF_IF_IF_3074_MINUS_SEXT_iFifo_first__087_B_ETC___d4436,
		IF_IF_IF_IF_3074_MINUS_SEXT_iFifo_first__087_B_ETC___d4438,
		IF_IF_IF_IF_3074_MINUS_SEXT_iFifo_first__087_B_ETC___d5211,
		IF_IF_IF_IF_3074_MINUS_SEXT_iFifo_first__087_B_ETC___d5213,
		IF_IF_IF_iFifo_first__087_BITS_102_TO_95_625_E_ETC___d5173,
		IF_IF_IF_iFifo_first__087_BITS_102_TO_95_625_E_ETC___d5175,
		IF_IF_IF_iFifo_first__087_BITS_102_TO_95_625_E_ETC___d5242,
		IF_IF_IF_iFifo_first__087_BITS_102_TO_95_625_E_ETC___d5244,
		IF_IF_IF_iFifo_first__087_BITS_167_TO_160_130__ETC___d3690,
		IF_IF_IF_iFifo_first__087_BITS_167_TO_160_130__ETC___d3692,
		IF_IF_IF_iFifo_first__087_BITS_167_TO_160_130__ETC___d3760,
		IF_IF_IF_iFifo_first__087_BITS_167_TO_160_130__ETC___d3762,
		IF_IF_IF_iFifo_first__087_BITS_37_TO_30_850_EQ_ETC___d4398,
		IF_IF_IF_iFifo_first__087_BITS_37_TO_30_850_EQ_ETC___d4400,
		IF_IF_IF_iFifo_first__087_BITS_37_TO_30_850_EQ_ETC___d4467,
		IF_IF_IF_iFifo_first__087_BITS_37_TO_30_850_EQ_ETC___d4469,
		IF_fpu_div_fOperands_S0_first__6_BITS_65_TO_55_ETC___d363,
		IF_fpu_div_fState_S4_first__73_BITS_64_TO_54_7_ETC___d907,
		IF_fpu_madd_fState_S8_first__960_BITS_65_TO_55_ETC___d2986,
		IF_fpu_madd_fState_S8_first__960_BITS_65_TO_55_ETC___d3011,
		IF_fpu_sqr_fState_S4_first__687_BITS_64_TO_54__ETC___d1721,
		SEXT_iFifo_first__087_BITS_102_TO_95_625_MINUS_ETC__q99,
		SEXT_iFifo_first__087_BITS_167_TO_160_130_MINU_ETC__q39,
		SEXT_iFifo_first__087_BITS_37_TO_30_850_MINUS__ETC__q66,
		_theResult___exp__h142541,
		_theResult___exp__h163979,
		_theResult___exp__h173569,
		_theResult___exp__h182321,
		_theResult___exp__h202617,
		_theResult___exp__h212207,
		_theResult___exp__h220959,
		_theResult___exp__h241556,
		_theResult___exp__h251146,
		_theResult___exp__h259898,
		_theResult___exp__h42526,
		_theResult___exp__h95909,
		_theResult___fst__h30373,
		_theResult___fst_exp__h130949,
		_theResult___fst_exp__h130952,
		_theResult___fst_exp__h130971,
		_theResult___fst_exp__h130986,
		_theResult___fst_exp__h131025,
		_theResult___fst_exp__h131031,
		_theResult___fst_exp__h131034,
		_theResult___fst_exp__h141375,
		_theResult___fst_exp__h141378,
		_theResult___fst_exp__h141397,
		_theResult___fst_exp__h141412,
		_theResult___fst_exp__h141451,
		_theResult___fst_exp__h141457,
		_theResult___fst_exp__h141460,
		_theResult___fst_exp__h163325,
		_theResult___fst_exp__h163331,
		_theResult___fst_exp__h163334,
		_theResult___fst_exp__h164060,
		_theResult___fst_exp__h172850,
		_theResult___fst_exp__h172915,
		_theResult___fst_exp__h172921,
		_theResult___fst_exp__h172924,
		_theResult___fst_exp__h173650,
		_theResult___fst_exp__h181603,
		_theResult___fst_exp__h181642,
		_theResult___fst_exp__h181648,
		_theResult___fst_exp__h181651,
		_theResult___fst_exp__h182402,
		_theResult___fst_exp__h182411,
		_theResult___fst_exp__h182414,
		_theResult___fst_exp__h201963,
		_theResult___fst_exp__h201969,
		_theResult___fst_exp__h201972,
		_theResult___fst_exp__h202698,
		_theResult___fst_exp__h211488,
		_theResult___fst_exp__h211553,
		_theResult___fst_exp__h211559,
		_theResult___fst_exp__h211562,
		_theResult___fst_exp__h212288,
		_theResult___fst_exp__h220241,
		_theResult___fst_exp__h220280,
		_theResult___fst_exp__h220286,
		_theResult___fst_exp__h220289,
		_theResult___fst_exp__h221040,
		_theResult___fst_exp__h221049,
		_theResult___fst_exp__h221052,
		_theResult___fst_exp__h240902,
		_theResult___fst_exp__h240908,
		_theResult___fst_exp__h240911,
		_theResult___fst_exp__h241637,
		_theResult___fst_exp__h250427,
		_theResult___fst_exp__h250492,
		_theResult___fst_exp__h250498,
		_theResult___fst_exp__h250501,
		_theResult___fst_exp__h251227,
		_theResult___fst_exp__h259180,
		_theResult___fst_exp__h259219,
		_theResult___fst_exp__h259225,
		_theResult___fst_exp__h259228,
		_theResult___fst_exp__h259979,
		_theResult___fst_exp__h259988,
		_theResult___fst_exp__h259991,
		_theResult___fst_exp__h41335,
		_theResult___fst_exp__h41338,
		_theResult___fst_exp__h41341,
		_theResult___fst_exp__h41384,
		_theResult___fst_exp__h41387,
		_theResult___fst_exp__h41407,
		_theResult___fst_exp__h41423,
		_theResult___fst_exp__h41462,
		_theResult___fst_exp__h41468,
		_theResult___fst_exp__h41471,
		_theResult___fst_exp__h42607,
		_theResult___fst_exp__h94750,
		_theResult___fst_exp__h94753,
		_theResult___fst_exp__h94773,
		_theResult___fst_exp__h94789,
		_theResult___fst_exp__h94828,
		_theResult___fst_exp__h94834,
		_theResult___fst_exp__h94837,
		_theResult___fst_exp__h95990,
		_theResult___snd_fst_exp__h164063,
		_theResult___snd_fst_exp__h182405,
		_theResult___snd_fst_exp__h202701,
		_theResult___snd_fst_exp__h221043,
		_theResult___snd_fst_exp__h241640,
		_theResult___snd_fst_exp__h259982,
		_theResult___snd_fst_exp__h30385,
		_theResult___snd_fst_exp__h30388,
		_theResult___snd_fst_exp__h30412,
		din_exp30866_MINUS_1023__q23,
		din_exp__h130866,
		din_inc___2_exp__h142626,
		din_inc___2_exp__h182467,
		din_inc___2_exp__h182502,
		din_inc___2_exp__h182528,
		din_inc___2_exp__h221105,
		din_inc___2_exp__h221140,
		din_inc___2_exp__h221166,
		din_inc___2_exp__h260044,
		din_inc___2_exp__h260079,
		din_inc___2_exp__h260105,
		din_inc___2_exp__h42617,
		din_inc___2_exp__h96000,
		fpu_div_fOperands_S0D_OUT_BITS_129_TO_119_MIN_ETC__q7,
		fpu_div_fOperands_S0D_OUT_BITS_65_TO_55_MINUS_ETC__q8,
		fpu_madd_fOperand_S0D_OUT_BITS_129_TO_119_MIN_ETC__q128,
		fpu_madd_fOperand_S0D_OUT_BITS_65_TO_55_MINUS_ETC__q129,
		fpu_madd_fState_S4D_OUT_BITS_128_TO_118_MINUS_ETC__q26,
		fpu_madd_fState_S4D_OUT_BITS_64_TO_54_MINUS_1023__q27,
		fpu_sqr_fOperand_S0D_OUT_BITS_65_TO_55_MINUS__ETC__q16,
		fpu_sqr_fState_S3D_OUT_BITS_121_TO_111_MINUS__ETC__q18,
		out_exp__h142544,
		out_exp__h163982,
		out_exp__h173572,
		out_exp__h182324,
		out_exp__h202620,
		out_exp__h212210,
		out_exp__h220962,
		out_exp__h241559,
		out_exp__h251149,
		out_exp__h259901,
		out_exp__h42529,
		out_exp__h95912,
		resWirewget_BITS_67_TO_57_MINUS_1023__q137,
		theResult___fst_exp1341_MINUS_1023__q11,
		value41307_BITS_10_TO_0_MINUS_1023__q28,
		x__h30592,
		x__h31820,
		x__h96539;
  wire [8 : 0] IF_SEXT_resWire_wget__410_BITS_67_TO_57_416_MI_ETC___d6332;
  wire [7 : 0] IF_IF_IF_IF_0b0_CONCAT_NOT_resWire_wget__410_B_ETC___d6448,
	       IF_IF_IF_IF_0b0_CONCAT_NOT_resWire_wget__410_B_ETC___d6450,
	       IF_IF_IF_IF_3970_MINUS_SEXT_resWire_wget__410__ETC___d6518,
	       IF_IF_IF_IF_3970_MINUS_SEXT_resWire_wget__410__ETC___d6520,
	       IF_IF_IF_resWire_wget__410_BITS_67_TO_57_416_E_ETC___d6479,
	       IF_IF_IF_resWire_wget__410_BITS_67_TO_57_416_E_ETC___d6481,
	       IF_IF_IF_resWire_wget__410_BITS_67_TO_57_416_E_ETC___d6549,
	       IF_IF_IF_resWire_wget__410_BITS_67_TO_57_416_E_ETC___d6551,
	       SEXT_resWire_wget__410_BITS_67_TO_57_416_MINUS_ETC__q141,
	       _theResult___exp__h278238,
	       _theResult___exp__h286820,
	       _theResult___exp__h296004,
	       _theResult___exp__h304640,
	       _theResult___fst_exp__h277722,
	       _theResult___fst_exp__h277787,
	       _theResult___fst_exp__h277793,
	       _theResult___fst_exp__h277796,
	       _theResult___fst_exp__h278319,
	       _theResult___fst_exp__h286369,
	       _theResult___fst_exp__h286375,
	       _theResult___fst_exp__h286378,
	       _theResult___fst_exp__h286901,
	       _theResult___fst_exp__h295488,
	       _theResult___fst_exp__h295553,
	       _theResult___fst_exp__h295559,
	       _theResult___fst_exp__h295562,
	       _theResult___fst_exp__h296085,
	       _theResult___fst_exp__h304125,
	       _theResult___fst_exp__h304164,
	       _theResult___fst_exp__h304170,
	       _theResult___fst_exp__h304173,
	       _theResult___fst_exp__h304721,
	       _theResult___fst_exp__h304730,
	       _theResult___fst_exp__h304733,
	       _theResult___snd_fst_exp__h286904,
	       _theResult___snd_fst_exp__h304724,
	       din_inc___2_exp__h304759,
	       din_inc___2_exp__h304785,
	       din_inc___2_exp__h304820,
	       din_inc___2_exp__h304846,
	       exp__h304742,
	       iFifoD_OUT_BITS_102_TO_95_MINUS_127__q95,
	       iFifoD_OUT_BITS_167_TO_160_MINUS_127__q35,
	       iFifoD_OUT_BITS_37_TO_30_MINUS_127__q62,
	       out_exp__h278241,
	       out_exp__h286823,
	       out_exp__h296007,
	       out_exp__h304643;
  wire [6 : 0] IF_IF_7170_MINUS_fpu_madd_fState_S3_first__995_ETC___d2460,
	       IF_fpu_sqr_fState_S1_first__216_BIT_57_226_THE_ETC___d1342,
	       x__h85465;
  wire [5 : 0] IF_IF_0b0_CONCAT_NOT_resWire_wget__410_BITS_67_ETC___d5767,
	       IF_IF_3074_MINUS_SEXT_iFifo_first__087_BITS_10_ETC___d5055,
	       IF_IF_3074_MINUS_SEXT_iFifo_first__087_BITS_16_ETC___d3572,
	       IF_IF_3074_MINUS_SEXT_iFifo_first__087_BITS_37_ETC___d4280,
	       IF_IF_3970_MINUS_SEXT_resWire_wget__410_BITS_6_ETC___d6278,
	       IF_IF_fpu_div_fState_S3_first__16_BITS_120_TO__ETC___d810,
	       IF_IF_fpu_madd_fState_S7_first__651_BIT_128_65_ETC___d2901,
	       IF_fpu_sqr_fOperand_S0_first__059_BITS_65_TO_5_ETC___d1193,
	       IF_fpu_sqr_fState_S3_first__375_BIT_58_384_THE_ETC___d1630,
	       IF_iFifo_first__087_BITS_102_TO_95_625_EQ_0_63_ETC___d4757,
	       IF_iFifo_first__087_BITS_167_TO_160_130_EQ_0_1_ETC___d3271,
	       IF_iFifo_first__087_BITS_37_TO_30_850_EQ_0_856_ETC___d3982,
	       IF_resWire_wget__410_BITS_67_TO_57_416_EQ_0_42_ETC___d5982,
	       b__h10508,
	       b__h3090,
	       x__h60732;
  wire [4 : 0] IF_IF_fpu_div_fState_S3_first__16_BITS_120_TO__ETC___d856,
	       IF_fpu_div_fState_S3_first__16_BITS_120_TO_110_ETC___d851,
	       IF_fpu_madd_fState_S3_first__995_BIT_151_996_T_ETC___d2525,
	       _0_CONCAT_IF_IF_0b0_CONCAT_NOT_resWire_wget__41_ETC___d6676,
	       _0_CONCAT_IF_IF_3970_MINUS_SEXT_resWire_wget__4_ETC___d6705,
	       _0_CONCAT_IF_resWire_wget__410_BITS_67_TO_57_41_ETC___d6688,
	       fpu_madd_fState_S3_first__995_BITS_86_TO_82_00_ETC___d2501,
	       fpu_madd_fState_S7_first__651_BITS_137_TO_133__ETC___d2942,
	       fpu_madd_fState_S8_first__960_BITS_75_TO_71_03_ETC___d3043,
	       resWire_wget__410_BITS_4_TO_0_658_OR_NOT_resWi_ETC___d6768;
  wire [2 : 0] IF_fpu_sqr_fState_S3_first__375_BIT_195_376_TH_ETC___d1671,
	       NOT_fpu_madd_fState_S3_first__995_BITS_12_TO_0_ETC___d2523;
  wire [1 : 0] IF_sfdin11482_BIT_4_THEN_2_ELSE_0__q98,
	       IF_sfdin1378_BIT_5_THEN_2_ELSE_0__q13,
	       IF_sfdin30943_BIT_53_THEN_2_ELSE_0__q25,
	       IF_sfdin41369_BIT_4_THEN_2_ELSE_0__q30,
	       IF_sfdin4744_BIT_6_THEN_2_ELSE_0__q20,
	       IF_sfdin50421_BIT_4_THEN_2_ELSE_0__q65,
	       IF_sfdin72844_BIT_4_THEN_2_ELSE_0__q38,
	       IF_sfdin77716_BIT_33_THEN_2_ELSE_0__q134,
	       IF_sfdin95482_BIT_33_THEN_2_ELSE_0__q140,
	       IF_theResult___snd01923_BIT_4_THEN_2_ELSE_0__q94,
	       IF_theResult___snd04119_BIT_33_THEN_2_ELSE_0__q143,
	       IF_theResult___snd20235_BIT_4_THEN_2_ELSE_0__q101,
	       IF_theResult___snd40862_BIT_4_THEN_2_ELSE_0__q61,
	       IF_theResult___snd59174_BIT_4_THEN_2_ELSE_0__q68,
	       IF_theResult___snd63285_BIT_4_THEN_2_ELSE_0__q34,
	       IF_theResult___snd81597_BIT_4_THEN_2_ELSE_0__q41,
	       IF_theResult___snd86329_BIT_33_THEN_2_ELSE_0__q136,
	       _theResult___snd_fst__h131051,
	       _theResult___snd_fst__h141477,
	       _theResult___snd_fst__h41490,
	       _theResult___snd_fst__h94856,
	       _theResult___snd_snd__h131371,
	       _theResult___snd_snd_snd__h131369,
	       guardBC__h115666,
	       guard__h133123,
	       guard__h155373,
	       guard__h164622,
	       guard__h173661,
	       guard__h194011,
	       guard__h203260,
	       guard__h212299,
	       guard__h232950,
	       guard__h242199,
	       guard__h251238,
	       guard__h269623,
	       guard__h278330,
	       guard__h287260,
	       guard__h296096,
	       guard__h32997,
	       guard__h86435,
	       x__h131406,
	       x__h141760,
	       x__h41756,
	       x__h95138;
  wire IF_3074_MINUS_0_CONCAT_IF_resWire_wget__410_BI_ETC___d6025,
       IF_3074_MINUS_0_CONCAT_IF_resWire_wget__410_BI_ETC___d6399,
       IF_3970_MINUS_0_CONCAT_IF_iFifo_first__087_BIT_ETC___d3317,
       IF_3970_MINUS_0_CONCAT_IF_iFifo_first__087_BIT_ETC___d4027,
       IF_3970_MINUS_0_CONCAT_IF_iFifo_first__087_BIT_ETC___d4581,
       IF_3970_MINUS_0_CONCAT_IF_iFifo_first__087_BIT_ETC___d4802,
       IF_3970_MINUS_0_CONCAT_IF_iFifo_first__087_BIT_ETC___d5347,
       IF_IF_fpu_madd_fOperand_S0_first__803_BIT_195__ETC___d1922,
       IF_NOT_fpu_madd_fState_S3_first__995_BITS_12_T_ETC___d2503,
       IF_NOT_fpu_madd_fState_S3_first__995_BITS_12_T_ETC___d2506,
       IF_SEXT_iFifo_first__087_BITS_102_TO_95_625_MI_ETC___d5146,
       IF_SEXT_iFifo_first__087_BITS_102_TO_95_625_MI_ETC___d5374,
       IF_SEXT_iFifo_first__087_BITS_167_TO_160_130_M_ETC___d3663,
       IF_SEXT_iFifo_first__087_BITS_37_TO_30_850_MIN_ETC___d4371,
       IF_SEXT_iFifo_first__087_BITS_37_TO_30_850_MIN_ETC___d4608,
       IF_SEXT_resWire_wget__410_BITS_67_TO_57_416_MI_ETC___d6375,
       IF_SEXT_resWire_wget__410_BITS_67_TO_57_416_MI_ETC___d6420,
       IF_SEXT_resWire_wget__410_BITS_67_TO_57_416_MI_ETC___d6734,
       IF_SEXT_resWire_wget__410_BITS_67_TO_57_416_MI_ETC___d6747,
       IF_SEXT_resWire_wget__410_BITS_67_TO_57_416_MI_ETC___d6760,
       IF_fpu_div_fOperands_S0_first__6_BITS_129_TO_1_ETC___d283,
       IF_fpu_div_fOperands_S0_first__6_BITS_129_TO_1_ETC___d285,
       IF_fpu_div_fOperands_S0_first__6_BITS_129_TO_1_ETC___d429,
       IF_fpu_div_fOperands_S0_first__6_BITS_65_TO_55_ETC___d352,
       IF_fpu_div_fState_S3_first__16_BITS_120_TO_110_ETC___d527,
       IF_fpu_madd_fOperand_S0_first__803_BIT_195_804_ETC___d1861,
       IF_fpu_madd_fOperand_S0_first__803_BIT_195_804_ETC___d1927,
       IF_fpu_madd_fOperand_S0_first__803_BIT_195_804_ETC___d1947,
       IF_fpu_madd_fState_S3_first__995_BITS_12_TO_0__ETC___d2516,
       IF_fpu_madd_fState_S3_first__995_BITS_12_TO_0__ETC___d2521,
       IF_fpu_madd_fState_S8_first__960_BIT_67_963_AN_ETC___d3060,
       IF_iFifo_first__087_BITS_102_TO_95_625_EQ_0_63_ETC___d5148,
       IF_iFifo_first__087_BITS_102_TO_95_625_EQ_0_63_ETC___d5376,
       IF_iFifo_first__087_BITS_167_TO_160_130_EQ_0_1_ETC___d3665,
       IF_iFifo_first__087_BITS_37_TO_30_850_EQ_0_856_ETC___d4373,
       IF_iFifo_first__087_BITS_37_TO_30_850_EQ_0_856_ETC___d4610,
       IF_isNegateFifo_first__409_THEN_IF_resWire_wge_ETC___d6424,
       IF_resWire_wget__410_BITS_67_TO_57_416_EQ_0_42_ETC___d6377,
       IF_resWire_wget__410_BITS_67_TO_57_416_EQ_0_42_ETC___d6422,
       IF_resWire_wget__410_BITS_67_TO_57_416_EQ_0_42_ETC___d6709,
       IF_resWire_wget__410_BITS_67_TO_57_416_EQ_0_42_ETC___d6720,
       IF_resWire_wget__410_BITS_67_TO_57_416_EQ_0_42_ETC___d6736,
       IF_resWire_wget__410_BITS_67_TO_57_416_EQ_0_42_ETC___d6749,
       IF_resWire_wget__410_BITS_67_TO_57_416_EQ_0_42_ETC___d6762,
       IF_rg_index_1_87_ULE_58_91_THEN_IF_rg_res_94_B_ETC___d1038,
       IF_rg_index_1_87_ULE_58_91_THEN_NOT_rg_b_92_EQ_ETC___d1009,
       IF_rg_index_1_87_ULE_58_91_THEN_rg_b_92_EQ_0_9_ETC___d997,
       NOT_3074_MINUS_0_CONCAT_IF_resWire_wget__410_B_ETC___d6728,
       NOT_3074_MINUS_0_CONCAT_IF_resWire_wget__410_B_ETC___d6756,
       NOT_IF_fpu_madd_fOperand_S0_first__803_BIT_195_ETC___d1946,
       NOT_fpu_div_fOperands_S0_first__6_BITS_129_TO__ETC___d330,
       NOT_fpu_div_fOperands_S0_first__6_BITS_65_TO_5_ETC___d411,
       NOT_fpu_div_fOperands_S0_first__6_BITS_65_TO_5_ETC___d418,
       NOT_fpu_madd_fOperand_S0_first__803_BITS_129_T_ETC___d1923,
       NOT_fpu_madd_fOperand_S0_first__803_BIT_130_85_ETC___d1854,
       NOT_fpu_madd_fState_S3_first__995_BITS_12_TO_0_ETC___d2510,
       NOT_fpu_madd_fState_S4_first__547_BIT_130_553__ETC___d2584,
       NOT_iFifo_first__087_BIT_158_142_202_AND_NOT_i_ETC___d3244,
       NOT_iFifo_first__087_BIT_28_862_913_AND_NOT_iF_ETC___d3955,
       NOT_iFifo_first__087_BIT_93_637_688_AND_NOT_iF_ETC___d4730,
       NOT_resWire_wget__410_BIT_56_426_825_AND_NOT_r_ETC___d5927,
       SEXT_iFifo_first__087_BITS_102_TO_95_625_MINUS_ETC___d4807,
       SEXT_iFifo_first__087_BITS_102_TO_95_625_MINUS_ETC___d4808,
       SEXT_iFifo_first__087_BITS_167_TO_160_130_MINU_ETC___d3324,
       SEXT_iFifo_first__087_BITS_167_TO_160_130_MINU_ETC___d3325,
       SEXT_iFifo_first__087_BITS_37_TO_30_850_MINUS__ETC___d4032,
       SEXT_iFifo_first__087_BITS_37_TO_30_850_MINUS__ETC___d4033,
       SEXT_resWire_wget__410_BITS_67_TO_57_416_MINUS_ETC___d6032,
       SEXT_resWire_wget__410_BITS_67_TO_57_416_MINUS_ETC___d6033,
       _0_CONCAT_IF_IF_0b0_CONCAT_NOT_resWire_wget__41_ETC___d5769,
       _0_CONCAT_IF_IF_3074_MINUS_SEXT_iFifo_first__08_ETC___d3574,
       _0_CONCAT_IF_IF_3074_MINUS_SEXT_iFifo_first__08_ETC___d4282,
       _0_CONCAT_IF_IF_3074_MINUS_SEXT_iFifo_first__08_ETC___d5057,
       _0_CONCAT_IF_IF_3970_MINUS_SEXT_resWire_wget__4_ETC___d6280,
       _0_CONCAT_IF_IF_7170_MINUS_fpu_madd_fState_S3_f_ETC___d2463,
       _0_CONCAT_IF_IF_fpu_div_fState_S3_first__16_BIT_ETC___d813,
       _0_CONCAT_IF_IF_fpu_madd_fState_S7_first__651_B_ETC___d2904,
       _0_CONCAT_IF_fpu_sqr_fState_S3_first__375_BIT_5_ETC___d1633,
       _0_CONCAT_IF_iFifo_first__087_BITS_102_TO_95_62_ETC___d4759,
       _0_CONCAT_IF_iFifo_first__087_BITS_102_TO_95_62_ETC___d5107,
       _0_CONCAT_IF_iFifo_first__087_BITS_167_TO_160_1_ETC___d3273,
       _0_CONCAT_IF_iFifo_first__087_BITS_167_TO_160_1_ETC___d3624,
       _0_CONCAT_IF_iFifo_first__087_BITS_37_TO_30_850_ETC___d3984,
       _0_CONCAT_IF_iFifo_first__087_BITS_37_TO_30_850_ETC___d4332,
       _0_CONCAT_IF_resWire_wget__410_BITS_67_TO_57_41_ETC___d5984,
       _0_CONCAT_IF_resWire_wget__410_BITS_67_TO_57_41_ETC___d6333,
       _3074_MINUS_0_CONCAT_IF_resWire_wget__410_BIT_5_ETC___d5532,
       _3074_MINUS_0_CONCAT_IF_resWire_wget__410_BIT_5_ETC___d5533,
       _3074_MINUS_0_CONCAT_IF_resWire_wget__410_BIT_5_ETC___d6691,
       _3074_MINUS_0_CONCAT_IF_resWire_wget__410_BIT_5_ETC___d6716,
       _3074_MINUS_0_CONCAT_IF_resWire_wget__410_BIT_5_ETC___d6743,
       _3970_MINUS_0_CONCAT_IF_iFifo_first__087_BIT_15_ETC___d3189,
       _3970_MINUS_0_CONCAT_IF_iFifo_first__087_BIT_15_ETC___d3190,
       _3970_MINUS_0_CONCAT_IF_iFifo_first__087_BIT_29_ETC___d3909,
       _3970_MINUS_0_CONCAT_IF_iFifo_first__087_BIT_29_ETC___d3910,
       _3970_MINUS_0_CONCAT_IF_iFifo_first__087_BIT_94_ETC___d4684,
       _3970_MINUS_0_CONCAT_IF_iFifo_first__087_BIT_94_ETC___d4685,
       _7170_MINUS_fpu_madd_fState_S3_first__995_BITS__ETC___d2008,
       fpu_div_fOperands_S0_first__6_BITS_129_TO_119__ETC___d293,
       fpu_div_fOperands_S0_first__6_BITS_129_TO_119__ETC___d331,
       fpu_div_fOperands_S0_first__6_BITS_129_TO_119__ETC___d366,
       fpu_div_fOperands_S0_first__6_BITS_129_TO_119__ETC___d428,
       fpu_div_fOperands_S0_first__6_BITS_65_TO_55_6__ETC___d289,
       fpu_div_fOperands_S0_first__6_BIT_130_33_EQ_fp_ETC___d335,
       fpu_madd_fOperand_S0_first__803_BITS_129_TO_11_ETC___d1857,
       fpu_madd_fOperand_S0_first__803_BITS_129_TO_11_ETC___d1926,
       fpu_madd_fOperand_S0_first__803_BIT_195_804_AN_ETC___d1855,
       fpu_madd_fState_S3_first__995_BITS_12_TO_0_001_ETC___d2002,
       fpu_madd_fState_S3_first__995_BITS_12_TO_0_001_ETC___d2004,
       guard__h165220,
       guard__h203858,
       guard__h242797,
       guard__h287858,
       rg_index_1_87_PLUS_1_89_ULE_58___d990,
       rg_index_1_87_ULE_58___d991,
       rg_index_PLUS_1_ULE_57___d6,
       rg_index_ULE_57___d7,
       rg_s_014_ULT_rg_r_1_013_PLUS_rg_b_92_015___d1016,
       sfdlsb__h116825,
       sfdlsb__h31694,
       value_BIT_52___h53270;
  // action method server_core_request_put
  assign RDY_server_core_request_put = iFifo$FULL_N ;
  assign CAN_FIRE_server_core_request_put = iFifo$FULL_N ;
  assign WILL_FIRE_server_core_request_put = EN_server_core_request_put ;
  // actionvalue method server_core_response_get
  assign server_core_response_get = oFifo$D_OUT ;
  assign RDY_server_core_response_get = oFifo$EMPTY_N ;
  assign CAN_FIRE_server_core_response_get = oFifo$EMPTY_N ;
  assign WILL_FIRE_server_core_response_get = EN_server_core_response_get ;
  // action method server_reset_request_put
  assign RDY_server_reset_request_put = resetReqsF$FULL_N ;
  assign CAN_FIRE_server_reset_request_put = resetReqsF$FULL_N ;
  assign WILL_FIRE_server_reset_request_put = EN_server_reset_request_put ;
  // action method server_reset_response_get
  assign RDY_server_reset_response_get = resetRspsF$EMPTY_N ;
  assign CAN_FIRE_server_reset_response_get = resetRspsF$EMPTY_N ;
  assign WILL_FIRE_server_reset_response_get = EN_server_reset_response_get ;
  // submodule fpu_div_fOperands_S0
  FIFOL1 #(.width(32'd131)) fpu_div_fOperands_S0(.RST(RST_N),
						 .CLK(CLK),
						 .D_IN(fpu_div_fOperands_S0$D_IN),
						 .ENQ(fpu_div_fOperands_S0$ENQ),
						 .DEQ(fpu_div_fOperands_S0$DEQ),
						 .CLR(fpu_div_fOperands_S0$CLR),
						 .D_OUT(fpu_div_fOperands_S0$D_OUT),
						 .FULL_N(fpu_div_fOperands_S0$FULL_N),
						 .EMPTY_N(fpu_div_fOperands_S0$EMPTY_N));
  // submodule fpu_div_fResult_S5
  FIFOL1 #(.width(32'd69)) fpu_div_fResult_S5(.RST(RST_N),
					      .CLK(CLK),
					      .D_IN(fpu_div_fResult_S5$D_IN),
					      .ENQ(fpu_div_fResult_S5$ENQ),
					      .DEQ(fpu_div_fResult_S5$DEQ),
					      .CLR(fpu_div_fResult_S5$CLR),
					      .D_OUT(fpu_div_fResult_S5$D_OUT),
					      .FULL_N(fpu_div_fResult_S5$FULL_N),
					      .EMPTY_N(fpu_div_fResult_S5$EMPTY_N));
  // submodule fpu_div_fState_S1
  FIFOL1 #(.width(32'd319)) fpu_div_fState_S1(.RST(RST_N),
					      .CLK(CLK),
					      .D_IN(fpu_div_fState_S1$D_IN),
					      .ENQ(fpu_div_fState_S1$ENQ),
					      .DEQ(fpu_div_fState_S1$DEQ),
					      .CLR(fpu_div_fState_S1$CLR),
					      .D_OUT(fpu_div_fState_S1$D_OUT),
					      .FULL_N(fpu_div_fState_S1$FULL_N),
					      .EMPTY_N(fpu_div_fState_S1$EMPTY_N));
  // submodule fpu_div_fState_S2
  FIFOL1 #(.width(32'd148)) fpu_div_fState_S2(.RST(RST_N),
					      .CLK(CLK),
					      .D_IN(fpu_div_fState_S2$D_IN),
					      .ENQ(fpu_div_fState_S2$ENQ),
					      .DEQ(fpu_div_fState_S2$DEQ),
					      .CLR(fpu_div_fState_S2$CLR),
					      .D_OUT(fpu_div_fState_S2$D_OUT),
					      .FULL_N(fpu_div_fState_S2$FULL_N),
					      .EMPTY_N(fpu_div_fState_S2$EMPTY_N));
  // submodule fpu_div_fState_S3
  FIFOL1 #(.width(32'd195)) fpu_div_fState_S3(.RST(RST_N),
					      .CLK(CLK),
					      .D_IN(fpu_div_fState_S3$D_IN),
					      .ENQ(fpu_div_fState_S3$ENQ),
					      .DEQ(fpu_div_fState_S3$DEQ),
					      .CLR(fpu_div_fState_S3$CLR),
					      .D_OUT(fpu_div_fState_S3$D_OUT),
					      .FULL_N(fpu_div_fState_S3$FULL_N),
					      .EMPTY_N(fpu_div_fState_S3$EMPTY_N));
  // submodule fpu_div_fState_S4
  FIFOL1 #(.width(32'd139)) fpu_div_fState_S4(.RST(RST_N),
					      .CLK(CLK),
					      .D_IN(fpu_div_fState_S4$D_IN),
					      .ENQ(fpu_div_fState_S4$ENQ),
					      .DEQ(fpu_div_fState_S4$DEQ),
					      .CLR(fpu_div_fState_S4$CLR),
					      .D_OUT(fpu_div_fState_S4$D_OUT),
					      .FULL_N(fpu_div_fState_S4$FULL_N),
					      .EMPTY_N(fpu_div_fState_S4$EMPTY_N));
  // submodule fpu_madd_fOperand_S0
  FIFOL1 #(.width(32'd196)) fpu_madd_fOperand_S0(.RST(RST_N),
						 .CLK(CLK),
						 .D_IN(fpu_madd_fOperand_S0$D_IN),
						 .ENQ(fpu_madd_fOperand_S0$ENQ),
						 .DEQ(fpu_madd_fOperand_S0$DEQ),
						 .CLR(fpu_madd_fOperand_S0$CLR),
						 .D_OUT(fpu_madd_fOperand_S0$D_OUT),
						 .FULL_N(fpu_madd_fOperand_S0$FULL_N),
						 .EMPTY_N(fpu_madd_fOperand_S0$EMPTY_N));
  // submodule fpu_madd_fProd_S2
  FIFOL1 #(.width(32'd106)) fpu_madd_fProd_S2(.RST(RST_N),
					      .CLK(CLK),
					      .D_IN(fpu_madd_fProd_S2$D_IN),
					      .ENQ(fpu_madd_fProd_S2$ENQ),
					      .DEQ(fpu_madd_fProd_S2$DEQ),
					      .CLR(fpu_madd_fProd_S2$CLR),
					      .D_OUT(fpu_madd_fProd_S2$D_OUT),
					      .FULL_N(fpu_madd_fProd_S2$FULL_N),
					      .EMPTY_N(fpu_madd_fProd_S2$EMPTY_N));
  // submodule fpu_madd_fProd_S3
  FIFOL1 #(.width(32'd106)) fpu_madd_fProd_S3(.RST(RST_N),
					      .CLK(CLK),
					      .D_IN(fpu_madd_fProd_S3$D_IN),
					      .ENQ(fpu_madd_fProd_S3$ENQ),
					      .DEQ(fpu_madd_fProd_S3$DEQ),
					      .CLR(fpu_madd_fProd_S3$CLR),
					      .D_OUT(fpu_madd_fProd_S3$D_OUT),
					      .FULL_N(fpu_madd_fProd_S3$FULL_N),
					      .EMPTY_N(fpu_madd_fProd_S3$EMPTY_N));
  // submodule fpu_madd_fResult_S9
  FIFOL1 #(.width(32'd69)) fpu_madd_fResult_S9(.RST(RST_N),
					       .CLK(CLK),
					       .D_IN(fpu_madd_fResult_S9$D_IN),
					       .ENQ(fpu_madd_fResult_S9$ENQ),
					       .DEQ(fpu_madd_fResult_S9$DEQ),
					       .CLR(fpu_madd_fResult_S9$CLR),
					       .D_OUT(fpu_madd_fResult_S9$D_OUT),
					       .FULL_N(fpu_madd_fResult_S9$FULL_N),
					       .EMPTY_N(fpu_madd_fResult_S9$EMPTY_N));
  // submodule fpu_madd_fState_S1
  FIFOL1 #(.width(32'd258)) fpu_madd_fState_S1(.RST(RST_N),
					       .CLK(CLK),
					       .D_IN(fpu_madd_fState_S1$D_IN),
					       .ENQ(fpu_madd_fState_S1$ENQ),
					       .DEQ(fpu_madd_fState_S1$DEQ),
					       .CLR(fpu_madd_fState_S1$CLR),
					       .D_OUT(fpu_madd_fState_S1$D_OUT),
					       .FULL_N(fpu_madd_fState_S1$FULL_N),
					       .EMPTY_N(fpu_madd_fState_S1$EMPTY_N));
  // submodule fpu_madd_fState_S2
  FIFOL1 #(.width(32'd152)) fpu_madd_fState_S2(.RST(RST_N),
					       .CLK(CLK),
					       .D_IN(fpu_madd_fState_S2$D_IN),
					       .ENQ(fpu_madd_fState_S2$ENQ),
					       .DEQ(fpu_madd_fState_S2$DEQ),
					       .CLR(fpu_madd_fState_S2$CLR),
					       .D_OUT(fpu_madd_fState_S2$D_OUT),
					       .FULL_N(fpu_madd_fState_S2$FULL_N),
					       .EMPTY_N(fpu_madd_fState_S2$EMPTY_N));
  // submodule fpu_madd_fState_S3
  FIFOL1 #(.width(32'd152)) fpu_madd_fState_S3(.RST(RST_N),
					       .CLK(CLK),
					       .D_IN(fpu_madd_fState_S3$D_IN),
					       .ENQ(fpu_madd_fState_S3$ENQ),
					       .DEQ(fpu_madd_fState_S3$DEQ),
					       .CLR(fpu_madd_fState_S3$CLR),
					       .D_OUT(fpu_madd_fState_S3$D_OUT),
					       .FULL_N(fpu_madd_fState_S3$FULL_N),
					       .EMPTY_N(fpu_madd_fState_S3$EMPTY_N));
  // submodule fpu_madd_fState_S4
  FIFOL1 #(.width(32'd204)) fpu_madd_fState_S4(.RST(RST_N),
					       .CLK(CLK),
					       .D_IN(fpu_madd_fState_S4$D_IN),
					       .ENQ(fpu_madd_fState_S4$ENQ),
					       .DEQ(fpu_madd_fState_S4$DEQ),
					       .CLR(fpu_madd_fState_S4$CLR),
					       .D_OUT(fpu_madd_fState_S4$D_OUT),
					       .FULL_N(fpu_madd_fState_S4$FULL_N),
					       .EMPTY_N(fpu_madd_fState_S4$EMPTY_N));
  // submodule fpu_madd_fState_S5
  FIFOL1 #(.width(32'd216)) fpu_madd_fState_S5(.RST(RST_N),
					       .CLK(CLK),
					       .D_IN(fpu_madd_fState_S5$D_IN),
					       .ENQ(fpu_madd_fState_S5$ENQ),
					       .DEQ(fpu_madd_fState_S5$DEQ),
					       .CLR(fpu_madd_fState_S5$CLR),
					       .D_OUT(fpu_madd_fState_S5$D_OUT),
					       .FULL_N(fpu_madd_fState_S5$FULL_N),
					       .EMPTY_N(fpu_madd_fState_S5$EMPTY_N));
  // submodule fpu_madd_fState_S6
  FIFOL1 #(.width(32'd203)) fpu_madd_fState_S6(.RST(RST_N),
					       .CLK(CLK),
					       .D_IN(fpu_madd_fState_S6$D_IN),
					       .ENQ(fpu_madd_fState_S6$ENQ),
					       .DEQ(fpu_madd_fState_S6$DEQ),
					       .CLR(fpu_madd_fState_S6$CLR),
					       .D_OUT(fpu_madd_fState_S6$D_OUT),
					       .FULL_N(fpu_madd_fState_S6$FULL_N),
					       .EMPTY_N(fpu_madd_fState_S6$EMPTY_N));
  // submodule fpu_madd_fState_S7
  FIFOL1 #(.width(32'd203)) fpu_madd_fState_S7(.RST(RST_N),
					       .CLK(CLK),
					       .D_IN(fpu_madd_fState_S7$D_IN),
					       .ENQ(fpu_madd_fState_S7$ENQ),
					       .DEQ(fpu_madd_fState_S7$DEQ),
					       .CLR(fpu_madd_fState_S7$CLR),
					       .D_OUT(fpu_madd_fState_S7$D_OUT),
					       .FULL_N(fpu_madd_fState_S7$FULL_N),
					       .EMPTY_N(fpu_madd_fState_S7$EMPTY_N));
  // submodule fpu_madd_fState_S8
  FIFOL1 #(.width(32'd141)) fpu_madd_fState_S8(.RST(RST_N),
					       .CLK(CLK),
					       .D_IN(fpu_madd_fState_S8$D_IN),
					       .ENQ(fpu_madd_fState_S8$ENQ),
					       .DEQ(fpu_madd_fState_S8$DEQ),
					       .CLR(fpu_madd_fState_S8$CLR),
					       .D_OUT(fpu_madd_fState_S8$D_OUT),
					       .FULL_N(fpu_madd_fState_S8$FULL_N),
					       .EMPTY_N(fpu_madd_fState_S8$EMPTY_N));
  // submodule fpu_sqr_fOperand_S0
  FIFOL1 #(.width(32'd67)) fpu_sqr_fOperand_S0(.RST(RST_N),
					       .CLK(CLK),
					       .D_IN(fpu_sqr_fOperand_S0$D_IN),
					       .ENQ(fpu_sqr_fOperand_S0$ENQ),
					       .DEQ(fpu_sqr_fOperand_S0$DEQ),
					       .CLR(fpu_sqr_fOperand_S0$CLR),
					       .D_OUT(fpu_sqr_fOperand_S0$D_OUT),
					       .FULL_N(fpu_sqr_fOperand_S0$FULL_N),
					       .EMPTY_N(fpu_sqr_fOperand_S0$EMPTY_N));
  // submodule fpu_sqr_fResult_S5
  FIFOL1 #(.width(32'd69)) fpu_sqr_fResult_S5(.RST(RST_N),
					      .CLK(CLK),
					      .D_IN(fpu_sqr_fResult_S5$D_IN),
					      .ENQ(fpu_sqr_fResult_S5$ENQ),
					      .DEQ(fpu_sqr_fResult_S5$DEQ),
					      .CLR(fpu_sqr_fResult_S5$CLR),
					      .D_OUT(fpu_sqr_fResult_S5$D_OUT),
					      .FULL_N(fpu_sqr_fResult_S5$FULL_N),
					      .EMPTY_N(fpu_sqr_fResult_S5$EMPTY_N));
  // submodule fpu_sqr_fState_S1
  FIFOL1 #(.width(32'd195)) fpu_sqr_fState_S1(.RST(RST_N),
					      .CLK(CLK),
					      .D_IN(fpu_sqr_fState_S1$D_IN),
					      .ENQ(fpu_sqr_fState_S1$ENQ),
					      .DEQ(fpu_sqr_fState_S1$DEQ),
					      .CLR(fpu_sqr_fState_S1$CLR),
					      .D_OUT(fpu_sqr_fState_S1$D_OUT),
					      .FULL_N(fpu_sqr_fState_S1$FULL_N),
					      .EMPTY_N(fpu_sqr_fState_S1$EMPTY_N));
  // submodule fpu_sqr_fState_S2
  FIFOL1 #(.width(32'd137)) fpu_sqr_fState_S2(.RST(RST_N),
					      .CLK(CLK),
					      .D_IN(fpu_sqr_fState_S2$D_IN),
					      .ENQ(fpu_sqr_fState_S2$ENQ),
					      .DEQ(fpu_sqr_fState_S2$DEQ),
					      .CLR(fpu_sqr_fState_S2$CLR),
					      .D_OUT(fpu_sqr_fState_S2$D_OUT),
					      .FULL_N(fpu_sqr_fState_S2$FULL_N),
					      .EMPTY_N(fpu_sqr_fState_S2$EMPTY_N));
  // submodule fpu_sqr_fState_S3
  FIFOL1 #(.width(32'd196)) fpu_sqr_fState_S3(.RST(RST_N),
					      .CLK(CLK),
					      .D_IN(fpu_sqr_fState_S3$D_IN),
					      .ENQ(fpu_sqr_fState_S3$ENQ),
					      .DEQ(fpu_sqr_fState_S3$DEQ),
					      .CLR(fpu_sqr_fState_S3$CLR),
					      .D_OUT(fpu_sqr_fState_S3$D_OUT),
					      .FULL_N(fpu_sqr_fState_S3$FULL_N),
					      .EMPTY_N(fpu_sqr_fState_S3$EMPTY_N));
  // submodule fpu_sqr_fState_S4
  FIFOL1 #(.width(32'd139)) fpu_sqr_fState_S4(.RST(RST_N),
					      .CLK(CLK),
					      .D_IN(fpu_sqr_fState_S4$D_IN),
					      .ENQ(fpu_sqr_fState_S4$ENQ),
					      .DEQ(fpu_sqr_fState_S4$DEQ),
					      .CLR(fpu_sqr_fState_S4$CLR),
					      .D_OUT(fpu_sqr_fState_S4$D_OUT),
					      .FULL_N(fpu_sqr_fState_S4$FULL_N),
					      .EMPTY_N(fpu_sqr_fState_S4$EMPTY_N));
  // submodule iFifo
  FIFO2 #(.width(32'd202), .guarded(32'd1)) iFifo(.RST(RST_N),
						  .CLK(CLK),
						  .D_IN(iFifo$D_IN),
						  .ENQ(iFifo$ENQ),
						  .DEQ(iFifo$DEQ),
						  .CLR(iFifo$CLR),
						  .D_OUT(iFifo$D_OUT),
						  .FULL_N(iFifo$FULL_N),
						  .EMPTY_N(iFifo$EMPTY_N));
  // submodule isDoubleFifo
  FIFO2 #(.width(32'd1), .guarded(32'd1)) isDoubleFifo(.RST(RST_N),
						       .CLK(CLK),
						       .D_IN(isDoubleFifo$D_IN),
						       .ENQ(isDoubleFifo$ENQ),
						       .DEQ(isDoubleFifo$DEQ),
						       .CLR(isDoubleFifo$CLR),
						       .D_OUT(isDoubleFifo$D_OUT),
						       .FULL_N(isDoubleFifo$FULL_N),
						       .EMPTY_N(isDoubleFifo$EMPTY_N));
  // submodule isNegateFifo
  FIFO2 #(.width(32'd1), .guarded(32'd1)) isNegateFifo(.RST(RST_N),
						       .CLK(CLK),
						       .D_IN(isNegateFifo$D_IN),
						       .ENQ(isNegateFifo$ENQ),
						       .DEQ(isNegateFifo$DEQ),
						       .CLR(isNegateFifo$CLR),
						       .D_OUT(isNegateFifo$D_OUT),
						       .FULL_N(isNegateFifo$FULL_N),
						       .EMPTY_N(isNegateFifo$EMPTY_N));
  // submodule oFifo
  FIFO2 #(.width(32'd70), .guarded(32'd1)) oFifo(.RST(RST_N),
						 .CLK(CLK),
						 .D_IN(oFifo$D_IN),
						 .ENQ(oFifo$ENQ),
						 .DEQ(oFifo$DEQ),
						 .CLR(oFifo$CLR),
						 .D_OUT(oFifo$D_OUT),
						 .FULL_N(oFifo$FULL_N),
						 .EMPTY_N(oFifo$EMPTY_N));
  // submodule resetReqsF
  FIFO20 #(.guarded(32'd1)) resetReqsF(.RST(RST_N),
				       .CLK(CLK),
				       .ENQ(resetReqsF$ENQ),
				       .DEQ(resetReqsF$DEQ),
				       .CLR(resetReqsF$CLR),
				       .FULL_N(resetReqsF$FULL_N),
				       .EMPTY_N(resetReqsF$EMPTY_N));
  // submodule resetRspsF
  FIFO20 #(.guarded(32'd1)) resetRspsF(.RST(RST_N),
				       .CLK(CLK),
				       .ENQ(resetRspsF$ENQ),
				       .DEQ(resetRspsF$DEQ),
				       .CLR(resetRspsF$CLR),
				       .FULL_N(resetRspsF$FULL_N),
				       .EMPTY_N(resetRspsF$EMPTY_N));
  // submodule rmdFifo
  FIFO2 #(.width(32'd3), .guarded(32'd1)) rmdFifo(.RST(RST_N),
						  .CLK(CLK),
						  .D_IN(rmdFifo$D_IN),
						  .ENQ(rmdFifo$ENQ),
						  .DEQ(rmdFifo$DEQ),
						  .CLR(rmdFifo$CLR),
						  .D_OUT(rmdFifo$D_OUT),
						  .FULL_N(rmdFifo$FULL_N),
						  .EMPTY_N(rmdFifo$EMPTY_N));
  // rule RL_getResFromPipe
  assign CAN_FIRE_RL_getResFromPipe = fpu_madd_fResult_S9$EMPTY_N ;
  assign WILL_FIRE_RL_getResFromPipe = fpu_madd_fResult_S9$EMPTY_N ;
  // rule RL_getResFromPipe_1
  assign CAN_FIRE_RL_getResFromPipe_1 = fpu_div_fResult_S5$EMPTY_N ;
  assign WILL_FIRE_RL_getResFromPipe_1 = fpu_div_fResult_S5$EMPTY_N ;
  // rule RL_getResFromPipe_2
  assign CAN_FIRE_RL_getResFromPipe_2 = fpu_sqr_fResult_S5$EMPTY_N ;
  assign WILL_FIRE_RL_getResFromPipe_2 = fpu_sqr_fResult_S5$EMPTY_N ;
  // rule __me_check_22
  assign CAN_FIRE___me_check_22 = 1'b1 ;
  assign WILL_FIRE___me_check_22 = 1'b1 ;
  // rule RL_passResult
  assign CAN_FIRE_RL_passResult =
	     isDoubleFifo$EMPTY_N && isNegateFifo$EMPTY_N &&
	     rmdFifo$EMPTY_N &&
	     oFifo$FULL_N &&
	     resWire$whas ;
  assign WILL_FIRE_RL_passResult = CAN_FIRE_RL_passResult ;
  // rule RL_fpu_div_s5_stage
  assign CAN_FIRE_RL_fpu_div_s5_stage =
	     fpu_div_fState_S4$EMPTY_N && fpu_div_fResult_S5$FULL_N ;
  assign WILL_FIRE_RL_fpu_div_s5_stage = CAN_FIRE_RL_fpu_div_s5_stage ;
  // rule RL_fpu_div_s4_stage
  assign CAN_FIRE_RL_fpu_div_s4_stage =
	     fpu_div_fState_S3$EMPTY_N && fpu_div_fState_S4$FULL_N ;
  assign WILL_FIRE_RL_fpu_div_s4_stage = CAN_FIRE_RL_fpu_div_s4_stage ;
  // rule RL_fpu_div_s3_stage
  assign CAN_FIRE_RL_fpu_div_s3_stage =
	     fpu_div_fState_S2$EMPTY_N && fpu_div_fState_S3$FULL_N &&
	     (fpu_div_fState_S2$D_OUT[147] || crg_done) ;
  assign WILL_FIRE_RL_fpu_div_s3_stage = CAN_FIRE_RL_fpu_div_s3_stage ;
  // rule RL_work
  assign CAN_FIRE_RL_work = rg_busy ;
  assign WILL_FIRE_RL_work = rg_busy ;
  // rule RL_fpu_div_s2_stage
  assign CAN_FIRE_RL_fpu_div_s2_stage =
	     fpu_div_fState_S1$EMPTY_N && fpu_div_fState_S2$FULL_N &&
	     (fpu_div_fState_S1$D_OUT[318] || !rg_busy) ;
  assign WILL_FIRE_RL_fpu_div_s2_stage =
	     CAN_FIRE_RL_fpu_div_s2_stage && !rg_busy ;
  // rule RL_fpu_div_s1_stage
  assign CAN_FIRE_RL_fpu_div_s1_stage =
	     fpu_div_fOperands_S0$EMPTY_N && fpu_div_fState_S1$FULL_N ;
  assign WILL_FIRE_RL_fpu_div_s1_stage = CAN_FIRE_RL_fpu_div_s1_stage ;
  // rule RL_fpu_sqr_s5_stage
  assign CAN_FIRE_RL_fpu_sqr_s5_stage =
	     fpu_sqr_fState_S4$EMPTY_N && fpu_sqr_fResult_S5$FULL_N ;
  assign WILL_FIRE_RL_fpu_sqr_s5_stage = CAN_FIRE_RL_fpu_sqr_s5_stage ;
  // rule RL_fpu_sqr_s4_stage
  assign CAN_FIRE_RL_fpu_sqr_s4_stage =
	     fpu_sqr_fState_S3$EMPTY_N && fpu_sqr_fState_S4$FULL_N ;
  assign WILL_FIRE_RL_fpu_sqr_s4_stage = CAN_FIRE_RL_fpu_sqr_s4_stage ;
  // rule RL_fpu_sqr_s3_stage
  assign CAN_FIRE_RL_fpu_sqr_s3_stage =
	     fpu_sqr_fState_S2$EMPTY_N && fpu_sqr_fState_S3$FULL_N &&
	     (fpu_sqr_fState_S2$D_OUT[136] || crg_done_1) ;
  assign WILL_FIRE_RL_fpu_sqr_s3_stage = CAN_FIRE_RL_fpu_sqr_s3_stage ;
  // rule RL_work_1
  assign CAN_FIRE_RL_work_1 = rg_busy_1 ;
  assign WILL_FIRE_RL_work_1 = rg_busy_1 ;
  // rule RL_fpu_sqr_s2_stage
  assign CAN_FIRE_RL_fpu_sqr_s2_stage =
	     fpu_sqr_fState_S1$EMPTY_N && fpu_sqr_fState_S2$FULL_N &&
	     (fpu_sqr_fState_S1$D_OUT[194] || !rg_busy_1) ;
  assign WILL_FIRE_RL_fpu_sqr_s2_stage =
	     CAN_FIRE_RL_fpu_sqr_s2_stage && !rg_busy_1 ;
  // rule RL_fpu_sqr_s1_stage
  assign CAN_FIRE_RL_fpu_sqr_s1_stage =
	     fpu_sqr_fOperand_S0$EMPTY_N && fpu_sqr_fState_S1$FULL_N ;
  assign WILL_FIRE_RL_fpu_sqr_s1_stage = CAN_FIRE_RL_fpu_sqr_s1_stage ;
  // rule RL_fpu_madd_s9_stage
  assign CAN_FIRE_RL_fpu_madd_s9_stage =
	     fpu_madd_fState_S8$EMPTY_N && fpu_madd_fResult_S9$FULL_N ;
  assign WILL_FIRE_RL_fpu_madd_s9_stage = CAN_FIRE_RL_fpu_madd_s9_stage ;
  // rule RL_fpu_madd_s8_stage
  assign CAN_FIRE_RL_fpu_madd_s8_stage =
	     fpu_madd_fState_S7$EMPTY_N && fpu_madd_fState_S8$FULL_N ;
  assign WILL_FIRE_RL_fpu_madd_s8_stage = CAN_FIRE_RL_fpu_madd_s8_stage ;
  // rule RL_fpu_madd_s7_stage
  assign CAN_FIRE_RL_fpu_madd_s7_stage =
	     fpu_madd_fState_S6$EMPTY_N && fpu_madd_fState_S7$FULL_N ;
  assign WILL_FIRE_RL_fpu_madd_s7_stage = CAN_FIRE_RL_fpu_madd_s7_stage ;
  // rule RL_fpu_madd_s6_stage
  assign CAN_FIRE_RL_fpu_madd_s6_stage =
	     fpu_madd_fState_S5$EMPTY_N && fpu_madd_fState_S6$FULL_N ;
  assign WILL_FIRE_RL_fpu_madd_s6_stage = CAN_FIRE_RL_fpu_madd_s6_stage ;
  // rule RL_fpu_madd_s5_stage
  assign CAN_FIRE_RL_fpu_madd_s5_stage =
	     fpu_madd_fState_S4$EMPTY_N && fpu_madd_fState_S5$FULL_N ;
  assign WILL_FIRE_RL_fpu_madd_s5_stage = CAN_FIRE_RL_fpu_madd_s5_stage ;
  // rule RL_fpu_madd_s4_stage
  assign CAN_FIRE_RL_fpu_madd_s4_stage =
	     fpu_madd_fState_S3$EMPTY_N && fpu_madd_fProd_S3$EMPTY_N &&
	     fpu_madd_fState_S4$FULL_N ;
  assign WILL_FIRE_RL_fpu_madd_s4_stage = CAN_FIRE_RL_fpu_madd_s4_stage ;
  // rule RL_fpu_madd_s3_stage
  assign CAN_FIRE_RL_fpu_madd_s3_stage =
	     fpu_madd_fState_S2$EMPTY_N && fpu_madd_fProd_S2$EMPTY_N &&
	     fpu_madd_fProd_S3$FULL_N &&
	     fpu_madd_fState_S3$FULL_N ;
  assign WILL_FIRE_RL_fpu_madd_s3_stage = CAN_FIRE_RL_fpu_madd_s3_stage ;
  // rule RL_fpu_madd_s2_stage
  assign CAN_FIRE_RL_fpu_madd_s2_stage =
	     fpu_madd_fState_S1$EMPTY_N && fpu_madd_fProd_S2$FULL_N &&
	     fpu_madd_fState_S2$FULL_N ;
  assign WILL_FIRE_RL_fpu_madd_s2_stage = CAN_FIRE_RL_fpu_madd_s2_stage ;
  // rule RL_fpu_madd_s1_stage
  assign CAN_FIRE_RL_fpu_madd_s1_stage =
	     fpu_madd_fOperand_S0$EMPTY_N && fpu_madd_fState_S1$FULL_N ;
  assign WILL_FIRE_RL_fpu_madd_s1_stage = CAN_FIRE_RL_fpu_madd_s1_stage ;
  // rule RL_start_op
  assign CAN_FIRE_RL_start_op =
	     iFifo$EMPTY_N && isDoubleFifo$FULL_N && isNegateFifo$FULL_N &&
	     rmdFifo$FULL_N &&
	     IF_iFifo_first__087_BITS_3_TO_0_088_EQ_0_089_O_ETC___d3110 ;
  assign WILL_FIRE_RL_start_op = CAN_FIRE_RL_start_op ;
  // rule RL_rl_reset
  assign CAN_FIRE_RL_rl_reset = resetReqsF$EMPTY_N && resetRspsF$FULL_N ;
  assign WILL_FIRE_RL_rl_reset = CAN_FIRE_RL_rl_reset ;
  // inputs to muxes for submodule ports
  assign MUX_crg_done$port1__write_1__SEL_1 = rg_busy && rg_index == 6'd28 ;
  assign MUX_crg_done_1$port1__write_1__SEL_1 =
	     rg_busy_1 && rg_index_1 == 6'd29 ;
  assign MUX_crg_done_1$port1__write_1__SEL_2 =
	     WILL_FIRE_RL_fpu_sqr_s2_stage && !fpu_sqr_fState_S1$D_OUT[194] ;
  assign MUX_rg_index$write_1__SEL_1 =
	     WILL_FIRE_RL_fpu_div_s2_stage && !fpu_div_fState_S1$D_OUT[318] ;
  assign MUX_rg_b$write_1__VAL_1 =
	     fpu_sqr_fState_S1$D_OUT[57] ?
	       116'h40000000000000000000000000000 :
	       b___1__h77160 ;
  assign MUX_rg_b$write_1__VAL_2 =
	     rg_index_1_87_PLUS_1_89_ULE_58___d990 ?
	       _theResult___fst__h43498 :
	       IF_rg_index_1_87_ULE_58_91_THEN_IF_rg_res_94_B_ETC___d1002 ;
  assign MUX_rg_d$write_1__VAL_1 = { 1'd0, fpu_div_fState_S1$D_OUT[67:11] } ;
  assign MUX_rg_index$write_1__VAL_2 = rg_index + 6'd1 ;
  assign MUX_rg_index_1$write_1__VAL_2 = rg_index_1 + 6'd1 ;
  assign MUX_rg_q$write_1__VAL_2 =
	     rg_index_PLUS_1_ULE_57___d6 ?
	       { IF_rg_index_ULE_57_THEN_rg_q_BITS_56_TO_0_CONC_ETC___d14[56:0],
		 !IF_rg_index_ULE_57_THEN_IF_rg_r_0_BIT_115_1_TH_ETC___d22[115] } :
	       IF_rg_index_ULE_57_THEN_rg_q_BITS_56_TO_0_CONC_ETC___d14 ;
  assign MUX_rg_r$write_1__VAL_1 = { 2'd0, fpu_div_fState_S1$D_OUT[181:68] } ;
  assign MUX_rg_r$write_1__VAL_2 =
	     rg_index_PLUS_1_ULE_57___d6 ?
	       (IF_rg_index_ULE_57_THEN_IF_rg_r_0_BIT_115_1_TH_ETC___d22[115] ?
		  { IF_rg_index_ULE_57_THEN_IF_rg_r_0_BIT_115_1_TH_ETC___d22[114:0],
		    1'd0 } +
		  b__h31634 :
		  { IF_rg_index_ULE_57_THEN_IF_rg_r_0_BIT_115_1_TH_ETC___d22[114:0],
		    1'd0 } -
		  b__h31634) :
	       IF_rg_index_ULE_57_THEN_IF_rg_r_0_BIT_115_1_TH_ETC___d22 ;
  assign MUX_rg_r_1$write_1__VAL_2 =
	     rg_index_1_87_PLUS_1_89_ULE_58___d990 ?
	       _theResult___snd_snd_snd__h43503 :
	       IF_rg_index_1_87_ULE_58_91_THEN_IF_rg_res_94_B_ETC___d1022 ;
  assign MUX_rg_res$write_1__VAL_2 =
	     { rg_index_1_87_PLUS_1_89_ULE_58___d990 ?
		 IF_rg_index_1_87_ULE_58_91_THEN_rg_b_92_EQ_0_9_ETC___d997 ||
		 IF_rg_index_1_87_ULE_58_91_THEN_IF_rg_res_94_B_ETC___d1002 ==
		 116'd0 :
		 IF_rg_index_1_87_ULE_58_91_THEN_rg_b_92_EQ_0_9_ETC___d997,
	       rg_index_1_87_PLUS_1_89_ULE_58___d990 ?
		 IF_IF_rg_index_1_87_ULE_58_91_THEN_NOT_rg_b_92_ETC___d1028 :
		 IF_rg_index_1_87_ULE_58_91_THEN_IF_rg_res_94_B_ETC___d1026 } ;
  assign MUX_rg_s$write_1__VAL_1 = { fpu_sqr_fState_S1$D_OUT[57:0], 58'd0 } ;
  assign MUX_rg_s$write_1__VAL_2 =
	     rg_index_1_87_PLUS_1_89_ULE_58___d990 ?
	       _theResult___snd_fst__h43500 :
	       IF_rg_index_1_87_ULE_58_91_THEN_IF_rg_res_94_B_ETC___d1036 ;
  // inlined wires
  always@(fpu_madd_fResult_S9$EMPTY_N or
	  fpu_madd_fResult_S9$D_OUT or
	  fpu_div_fResult_S5$EMPTY_N or
	  fpu_div_fResult_S5$D_OUT or
	  fpu_sqr_fResult_S5$EMPTY_N or fpu_sqr_fResult_S5$D_OUT)
  begin
    case (1'b1) // synopsys parallel_case
      fpu_madd_fResult_S9$EMPTY_N: resWire$wget = fpu_madd_fResult_S9$D_OUT;
      fpu_div_fResult_S5$EMPTY_N: resWire$wget = fpu_div_fResult_S5$D_OUT;
      fpu_sqr_fResult_S5$EMPTY_N: resWire$wget = fpu_sqr_fResult_S5$D_OUT;
      default: resWire$wget = 69'h0AAAAAAAAAAAAAAAAA /* unspecified value */ ;
    endcase
  end
  assign resWire$whas =
	     fpu_madd_fResult_S9$EMPTY_N || fpu_div_fResult_S5$EMPTY_N ||
	     fpu_sqr_fResult_S5$EMPTY_N ;
  assign crg_done$EN_port0__write =
	     WILL_FIRE_RL_fpu_div_s3_stage && !fpu_div_fState_S2$D_OUT[147] ;
  assign crg_done$port1__read = !crg_done$EN_port0__write && crg_done ;
  assign crg_done$EN_port1__write =
	     rg_busy && rg_index == 6'd28 ||
	     WILL_FIRE_RL_fpu_div_s2_stage && !fpu_div_fState_S1$D_OUT[318] ;
  assign crg_done$port2__read =
	     crg_done$EN_port1__write ?
	       MUX_crg_done$port1__write_1__SEL_1 :
	       crg_done$port1__read ;
  assign crg_done_1$EN_port0__write =
	     WILL_FIRE_RL_fpu_sqr_s3_stage && !fpu_sqr_fState_S2$D_OUT[136] ;
  assign crg_done_1$port1__read = !crg_done_1$EN_port0__write && crg_done_1 ;
  assign crg_done_1$EN_port1__write =
	     rg_busy_1 && rg_index_1 == 6'd29 ||
	     WILL_FIRE_RL_fpu_sqr_s2_stage && !fpu_sqr_fState_S1$D_OUT[194] ;
  assign crg_done_1$port2__read =
	     crg_done_1$EN_port1__write ?
	       MUX_crg_done_1$port1__write_1__SEL_1 :
	       crg_done_1$port1__read ;
  // register crg_done
  assign crg_done$D_IN = crg_done$port2__read ;
  assign crg_done$EN = 1'b1 ;
  // register crg_done_1
  assign crg_done_1$D_IN = crg_done_1$port2__read ;
  assign crg_done_1$EN = 1'b1 ;
  // register rg_b
  assign rg_b$D_IN =
	     MUX_crg_done_1$port1__write_1__SEL_2 ?
	       MUX_rg_b$write_1__VAL_1 :
	       MUX_rg_b$write_1__VAL_2 ;
  assign rg_b$EN =
	     WILL_FIRE_RL_fpu_sqr_s2_stage && !fpu_sqr_fState_S1$D_OUT[194] ||
	     rg_busy_1 ;
  // register rg_busy
  assign rg_busy$D_IN = !MUX_crg_done$port1__write_1__SEL_1 ;
  assign rg_busy$EN =
	     rg_busy && rg_index == 6'd28 ||
	     WILL_FIRE_RL_fpu_div_s2_stage && !fpu_div_fState_S1$D_OUT[318] ;
  // register rg_busy_1
  assign rg_busy_1$D_IN = !MUX_crg_done_1$port1__write_1__SEL_1 ;
  assign rg_busy_1$EN =
	     rg_busy_1 && rg_index_1 == 6'd29 ||
	     WILL_FIRE_RL_fpu_sqr_s2_stage && !fpu_sqr_fState_S1$D_OUT[194] ;
  // register rg_d
  assign rg_d$D_IN =
	     MUX_rg_index$write_1__SEL_1 ? MUX_rg_d$write_1__VAL_1 : rg_d ;
  assign rg_d$EN =
	     WILL_FIRE_RL_fpu_div_s2_stage && !fpu_div_fState_S1$D_OUT[318] ||
	     rg_busy ;
  // register rg_index
  assign rg_index$D_IN =
	     MUX_rg_index$write_1__SEL_1 ?
	       6'd0 :
	       MUX_rg_index$write_1__VAL_2 ;
  assign rg_index$EN =
	     WILL_FIRE_RL_fpu_div_s2_stage && !fpu_div_fState_S1$D_OUT[318] ||
	     rg_busy ;
  // register rg_index_1
  assign rg_index_1$D_IN =
	     MUX_crg_done_1$port1__write_1__SEL_2 ?
	       6'd0 :
	       MUX_rg_index_1$write_1__VAL_2 ;
  assign rg_index_1$EN =
	     WILL_FIRE_RL_fpu_sqr_s2_stage && !fpu_sqr_fState_S1$D_OUT[194] ||
	     rg_busy_1 ;
  // register rg_q
  assign rg_q$D_IN =
	     MUX_rg_index$write_1__SEL_1 ? 58'd0 : MUX_rg_q$write_1__VAL_2 ;
  assign rg_q$EN =
	     WILL_FIRE_RL_fpu_div_s2_stage && !fpu_div_fState_S1$D_OUT[318] ||
	     rg_busy ;
  // register rg_r
  assign rg_r$D_IN =
	     MUX_rg_index$write_1__SEL_1 ?
	       MUX_rg_r$write_1__VAL_1 :
	       MUX_rg_r$write_1__VAL_2 ;
  assign rg_r$EN =
	     WILL_FIRE_RL_fpu_div_s2_stage && !fpu_div_fState_S1$D_OUT[318] ||
	     rg_busy ;
  // register rg_r_1
  assign rg_r_1$D_IN =
	     MUX_crg_done_1$port1__write_1__SEL_2 ?
	       116'd0 :
	       MUX_rg_r_1$write_1__VAL_2 ;
  assign rg_r_1$EN =
	     WILL_FIRE_RL_fpu_sqr_s2_stage && !fpu_sqr_fState_S1$D_OUT[194] ||
	     rg_busy_1 ;
  // register rg_res
  assign rg_res$D_IN =
	     MUX_crg_done_1$port1__write_1__SEL_2 ?
	       117'h0AAAAAAAAAAAAAAAAAAAAAAAAAAAAA :
	       MUX_rg_res$write_1__VAL_2 ;
  assign rg_res$EN =
	     WILL_FIRE_RL_fpu_sqr_s2_stage && !fpu_sqr_fState_S1$D_OUT[194] ||
	     rg_busy_1 ;
  // register rg_s
  assign rg_s$D_IN =
	     MUX_crg_done_1$port1__write_1__SEL_2 ?
	       MUX_rg_s$write_1__VAL_1 :
	       MUX_rg_s$write_1__VAL_2 ;
  assign rg_s$EN =
	     WILL_FIRE_RL_fpu_sqr_s2_stage && !fpu_sqr_fState_S1$D_OUT[194] ||
	     rg_busy_1 ;
  // submodule fpu_div_fOperands_S0
  assign fpu_div_fOperands_S0$D_IN =
	     { IF_iFifo_first__087_BIT_201_115_THEN_IF_iFifo__ETC___d3848,
	       IF_iFifo_first__087_BIT_136_624_THEN_IF_iFifo__ETC___d5330,
	       iFifo$D_OUT[6:4] } ;
  assign fpu_div_fOperands_S0$ENQ =
	     WILL_FIRE_RL_start_op && iFifo$D_OUT[3:0] == 4'd3 ;
  assign fpu_div_fOperands_S0$DEQ = CAN_FIRE_RL_fpu_div_s1_stage ;
  assign fpu_div_fOperands_S0$CLR = 1'b0 ;
  // submodule fpu_div_fResult_S5
  assign fpu_div_fResult_S5$D_IN =
	     fpu_div_fState_S4$D_OUT[138] ?
	       fpu_div_fState_S4$D_OUT[137:69] :
	       { (fpu_div_fState_S4$D_OUT[64:54] == 11'd2047) ?
		   fpu_div_fState_S4$D_OUT[65:2] :
		   CASE_fpu_div_fState_S4D_OUT_BITS_68_TO_66_0_C_ETC__q173,
		 fpu_div_fState_S4$D_OUT[73:69] |
		 { 2'd0,
		   _theResult___fst_exp__h42607 == 11'd2047 &&
		   _theResult___fst_sfd__h42608 == 52'd0,
		   1'd0,
		   fpu_div_fState_S4$D_OUT[64:54] != 11'd2047 &&
		   fpu_div_fState_S4$D_OUT[1:0] != 2'b0 } } ;
  assign fpu_div_fResult_S5$ENQ = CAN_FIRE_RL_fpu_div_s5_stage ;
  assign fpu_div_fResult_S5$DEQ = fpu_div_fResult_S5$EMPTY_N ;
  assign fpu_div_fResult_S5$CLR = 1'b0 ;
  // submodule fpu_div_fState_S1
  assign fpu_div_fState_S1$D_IN =
	     { fpu_div_fOperands_S0_first__6_BITS_129_TO_119__ETC___d293,
	       (fpu_div_fOperands_S0$D_OUT[129:119] == 11'd2047 &&
		fpu_div_fOperands_S0$D_OUT[118:67] != 52'd0 &&
		!fpu_div_fOperands_S0$D_OUT[118]) ?
		 { fpu_div_fOperands_S0$D_OUT[130:119], sfd__h17985 } :
		 IF_fpu_div_fOperands_S0_first__6_BITS_65_TO_55_ETC___d385,
	       fpu_div_fOperands_S0$D_OUT[129:119] == 11'd2047 &&
	       fpu_div_fOperands_S0$D_OUT[118:67] != 52'd0 &&
	       !fpu_div_fOperands_S0$D_OUT[118] ||
	       fpu_div_fOperands_S0$D_OUT[65:55] == 11'd2047 &&
	       fpu_div_fOperands_S0$D_OUT[54:3] != 52'd0 &&
	       !fpu_div_fOperands_S0$D_OUT[54] ||
	       (fpu_div_fOperands_S0$D_OUT[129:119] != 11'd2047 ||
		!fpu_div_fOperands_S0$D_OUT[118]) &&
	       (fpu_div_fOperands_S0$D_OUT[65:55] != 11'd2047 ||
		!fpu_div_fOperands_S0$D_OUT[54]) &&
	       fpu_div_fOperands_S0_first__6_BITS_129_TO_119__ETC___d366,
	       (fpu_div_fOperands_S0$D_OUT[129:119] != 11'd2047 ||
		fpu_div_fOperands_S0$D_OUT[118:67] == 52'd0 ||
		fpu_div_fOperands_S0$D_OUT[118]) &&
	       (fpu_div_fOperands_S0$D_OUT[129:119] != 11'd2047 ||
		!fpu_div_fOperands_S0$D_OUT[118]) &&
	       NOT_fpu_div_fOperands_S0_first__6_BITS_129_TO__ETC___d330 &&
	       fpu_div_fOperands_S0$D_OUT[65:55] == 11'd0 &&
	       fpu_div_fOperands_S0$D_OUT[54:3] == 52'd0 &&
	       (fpu_div_fOperands_S0$D_OUT[129:119] != 11'd2047 ||
		fpu_div_fOperands_S0$D_OUT[118:67] != 52'd0),
	       (fpu_div_fOperands_S0$D_OUT[129:119] != 11'd2047 ||
		fpu_div_fOperands_S0$D_OUT[118:67] == 52'd0 ||
		fpu_div_fOperands_S0$D_OUT[118]) &&
	       (fpu_div_fOperands_S0$D_OUT[65:55] != 11'd2047 ||
		fpu_div_fOperands_S0$D_OUT[54:3] == 52'd0 ||
		fpu_div_fOperands_S0$D_OUT[54]) &&
	       (fpu_div_fOperands_S0$D_OUT[129:119] != 11'd2047 ||
		!fpu_div_fOperands_S0$D_OUT[118]) &&
	       (fpu_div_fOperands_S0$D_OUT[65:55] != 11'd2047 ||
		!fpu_div_fOperands_S0$D_OUT[54]) &&
	       (fpu_div_fOperands_S0$D_OUT[65:55] != 11'd0 ||
		fpu_div_fOperands_S0$D_OUT[54:3] != 52'd0) &&
	       (fpu_div_fOperands_S0$D_OUT[129:119] != 11'd2047 ||
		fpu_div_fOperands_S0$D_OUT[118:67] != 52'd0) &&
	       (fpu_div_fOperands_S0$D_OUT[129:119] != 11'd0 ||
		fpu_div_fOperands_S0$D_OUT[118:67] != 52'd0) &&
	       (fpu_div_fOperands_S0$D_OUT[65:55] != 11'd2047 ||
		fpu_div_fOperands_S0$D_OUT[54:3] != 52'd0) &&
	       !IF_fpu_div_fOperands_S0_first__6_BITS_129_TO_1_ETC___d283,
	       (fpu_div_fOperands_S0$D_OUT[129:119] != 11'd2047 ||
		fpu_div_fOperands_S0$D_OUT[118:67] == 52'd0 ||
		fpu_div_fOperands_S0$D_OUT[118]) &&
	       (fpu_div_fOperands_S0$D_OUT[65:55] != 11'd2047 ||
		fpu_div_fOperands_S0$D_OUT[54:3] == 52'd0 ||
		fpu_div_fOperands_S0$D_OUT[54]) &&
	       (fpu_div_fOperands_S0$D_OUT[129:119] != 11'd2047 ||
		!fpu_div_fOperands_S0$D_OUT[118]) &&
	       (fpu_div_fOperands_S0$D_OUT[65:55] != 11'd2047 ||
		!fpu_div_fOperands_S0$D_OUT[54]) &&
	       NOT_fpu_div_fOperands_S0_first__6_BITS_65_TO_5_ETC___d411,
	       (fpu_div_fOperands_S0$D_OUT[129:119] != 11'd2047 ||
		fpu_div_fOperands_S0$D_OUT[118:67] == 52'd0 ||
		fpu_div_fOperands_S0$D_OUT[118]) &&
	       (fpu_div_fOperands_S0$D_OUT[65:55] != 11'd2047 ||
		fpu_div_fOperands_S0$D_OUT[54:3] == 52'd0 ||
		fpu_div_fOperands_S0$D_OUT[54]) &&
	       (fpu_div_fOperands_S0$D_OUT[129:119] != 11'd2047 ||
		!fpu_div_fOperands_S0$D_OUT[118]) &&
	       (fpu_div_fOperands_S0$D_OUT[65:55] != 11'd2047 ||
		!fpu_div_fOperands_S0$D_OUT[54]) &&
	       NOT_fpu_div_fOperands_S0_first__6_BITS_65_TO_5_ETC___d418,
	       fpu_div_fOperands_S0$D_OUT[2:0],
	       !fpu_div_fOperands_S0_first__6_BIT_130_33_EQ_fp_ETC___d335,
	       _theResult___snd_fst_exp__h30412,
	       _theResult___snd_fst_sfd__h30413,
	       x__h30477,
	       x__h30538,
	       x__h30592 } ;
  assign fpu_div_fState_S1$ENQ = CAN_FIRE_RL_fpu_div_s1_stage ;
  assign fpu_div_fState_S1$DEQ = WILL_FIRE_RL_fpu_div_s2_stage ;
  assign fpu_div_fState_S1$CLR = 1'b0 ;
  // submodule fpu_div_fState_S2
  assign fpu_div_fState_S2$D_IN =
	     { fpu_div_fState_S1$D_OUT[318:182],
	       fpu_div_fState_S1$D_OUT[10:0] } ;
  assign fpu_div_fState_S2$ENQ = WILL_FIRE_RL_fpu_div_s2_stage ;
  assign fpu_div_fState_S2$DEQ = CAN_FIRE_RL_fpu_div_s3_stage ;
  assign fpu_div_fState_S2$CLR = 1'b0 ;
  // submodule fpu_div_fState_S3
  assign fpu_div_fState_S3$D_IN =
	     { fpu_div_fState_S2$D_OUT[147:11], x__h32103 } ;
  assign fpu_div_fState_S3$ENQ = CAN_FIRE_RL_fpu_div_s3_stage ;
  assign fpu_div_fState_S3$DEQ = CAN_FIRE_RL_fpu_div_s4_stage ;
  assign fpu_div_fState_S3$CLR = 1'b0 ;
  // submodule fpu_div_fState_S4
  assign fpu_div_fState_S4$D_IN =
	     { (fpu_div_fState_S3$D_OUT[120:110] == 11'd2047) ?
		 fpu_div_fState_S3$D_OUT[57:56] != 2'b0 ||
		 fpu_div_fState_S3$D_OUT[194] :
		 fpu_div_fState_S3$D_OUT[194],
	       (fpu_div_fState_S3$D_OUT[120:110] == 11'd2047) ?
		 ((fpu_div_fState_S3$D_OUT[57:56] == 2'b0) ?
		    fpu_div_fState_S3$D_OUT[193:130] :
		    { CASE_fpu_div_fState_S3D_OUT_BITS_124_TO_122_0_ETC__q174,
		      CASE_fpu_div_fState_S3D_OUT_BITS_124_TO_122_0_ETC__q175 }) :
		 fpu_div_fState_S3$D_OUT[193:130],
	       IF_IF_fpu_div_fState_S3_first__16_BITS_120_TO__ETC___d856,
	       fpu_div_fState_S3$D_OUT[124:122],
	       fpu_div_fState_S3_first__16_BIT_121_37_CONCAT__ETC___d866,
	       x__h41756 } ;
  assign fpu_div_fState_S4$ENQ = CAN_FIRE_RL_fpu_div_s4_stage ;
  assign fpu_div_fState_S4$DEQ = CAN_FIRE_RL_fpu_div_s5_stage ;
  assign fpu_div_fState_S4$CLR = 1'b0 ;
  // submodule fpu_madd_fOperand_S0
  assign fpu_madd_fOperand_S0$D_IN =
	     { iFifo$D_OUT[3:0] != 4'd2,
	       IF_iFifo_first__087_BITS_3_TO_0_088_EQ_0_089_O_ETC___d4623,
	       CASE_iFifoD_OUT_BITS_3_TO_0_0_IF_iFifo_first__ETC__q176,
	       CASE_iFifoD_OUT_BITS_3_TO_0_0_460718241880001_ETC__q177,
	       iFifo$D_OUT[6:4] } ;
  assign fpu_madd_fOperand_S0$ENQ =
	     WILL_FIRE_RL_start_op &&
	     (iFifo$D_OUT[3:0] == 4'd0 || iFifo$D_OUT[3:0] == 4'd1 ||
	      iFifo$D_OUT[3:0] == 4'd2 ||
	      iFifo$D_OUT[3:0] == 4'd5 ||
	      iFifo$D_OUT[3:0] == 4'd6 ||
	      iFifo$D_OUT[3:0] == 4'd7 ||
	      iFifo$D_OUT[3:0] == 4'd8) ;
  assign fpu_madd_fOperand_S0$DEQ = CAN_FIRE_RL_fpu_madd_s1_stage ;
  assign fpu_madd_fOperand_S0$CLR = 1'b0 ;
  // submodule fpu_madd_fProd_S2
  assign fpu_madd_fProd_S2$D_IN =
	     fpu_madd_fState_S1$D_OUT[105:53] *
	     fpu_madd_fState_S1$D_OUT[52:0] ;
  assign fpu_madd_fProd_S2$ENQ = CAN_FIRE_RL_fpu_madd_s2_stage ;
  assign fpu_madd_fProd_S2$DEQ = CAN_FIRE_RL_fpu_madd_s3_stage ;
  assign fpu_madd_fProd_S2$CLR = 1'b0 ;
  // submodule fpu_madd_fProd_S3
  assign fpu_madd_fProd_S3$D_IN = fpu_madd_fProd_S2$D_OUT ;
  assign fpu_madd_fProd_S3$ENQ = CAN_FIRE_RL_fpu_madd_s3_stage ;
  assign fpu_madd_fProd_S3$DEQ = CAN_FIRE_RL_fpu_madd_s4_stage ;
  assign fpu_madd_fProd_S3$CLR = 1'b0 ;
  // submodule fpu_madd_fResult_S9
  assign fpu_madd_fResult_S9$D_IN =
	     fpu_madd_fState_S8$D_OUT[140] ?
	       fpu_madd_fState_S8$D_OUT[139:71] :
	       IF_fpu_madd_fState_S8_first__960_BIT_67_963_AN_ETC___d3081 ;
  assign fpu_madd_fResult_S9$ENQ = CAN_FIRE_RL_fpu_madd_s9_stage ;
  assign fpu_madd_fResult_S9$DEQ = fpu_madd_fResult_S9$EMPTY_N ;
  assign fpu_madd_fResult_S9$CLR = 1'b0 ;
  // submodule fpu_madd_fState_S1
  assign fpu_madd_fState_S1$D_IN =
	     { x__h96539 == 11'd2047 &&
	       _theResult___fst_sfd__h96608 != 52'd0 &&
	       !_theResult___fst_sfd__h96608[51] ||
	       fpu_madd_fOperand_S0$D_OUT[129:119] == 11'd2047 &&
	       fpu_madd_fOperand_S0$D_OUT[118:67] != 52'd0 &&
	       !fpu_madd_fOperand_S0$D_OUT[118] ||
	       fpu_madd_fOperand_S0$D_OUT[65:55] == 11'd2047 &&
	       fpu_madd_fOperand_S0$D_OUT[54:3] != 52'd0 &&
	       !fpu_madd_fOperand_S0$D_OUT[54] ||
	       IF_fpu_madd_fOperand_S0_first__803_BIT_195_804_ETC___d1861,
	       IF_IF_fpu_madd_fOperand_S0_first__803_BIT_195__ETC___d1939,
	       IF_fpu_madd_fOperand_S0_first__803_BIT_195_804_ETC___d1947,
	       4'd0,
	       fpu_madd_fOperand_S0$D_OUT[2:0],
	       fpu_madd_fOperand_S0$D_OUT[195],
	       fpu_madd_fOperand_S0$D_OUT[195] &&
	       fpu_madd_fOperand_S0$D_OUT[194],
	       IF_fpu_madd_fOperand_S0_first__803_BIT_195_804_ETC___d1911,
	       NOT_fpu_madd_fOperand_S0_first__803_BIT_130_85_ETC___d1854,
	       IF_fpu_madd_fOperand_S0_first__803_BITS_129_TO_ETC___d1959 } ;
  assign fpu_madd_fState_S1$ENQ = CAN_FIRE_RL_fpu_madd_s1_stage ;
  assign fpu_madd_fState_S1$DEQ = CAN_FIRE_RL_fpu_madd_s2_stage ;
  assign fpu_madd_fState_S1$CLR = 1'b0 ;
  // submodule fpu_madd_fState_S2
  assign fpu_madd_fState_S2$D_IN = fpu_madd_fState_S1$D_OUT[257:106] ;
  assign fpu_madd_fState_S2$ENQ = CAN_FIRE_RL_fpu_madd_s2_stage ;
  assign fpu_madd_fState_S2$DEQ = CAN_FIRE_RL_fpu_madd_s3_stage ;
  assign fpu_madd_fState_S2$CLR = 1'b0 ;
  // submodule fpu_madd_fState_S3
  assign fpu_madd_fState_S3$D_IN = fpu_madd_fState_S2$D_OUT ;
  assign fpu_madd_fState_S3$ENQ = CAN_FIRE_RL_fpu_madd_s3_stage ;
  assign fpu_madd_fState_S3$DEQ = CAN_FIRE_RL_fpu_madd_s4_stage ;
  assign fpu_madd_fState_S3$CLR = 1'b0 ;
  // submodule fpu_madd_fState_S4
  assign fpu_madd_fState_S4$D_IN =
	     { fpu_madd_fState_S3$D_OUT[151:87],
	       IF_fpu_madd_fState_S3_first__995_BIT_151_996_T_ETC___d2525,
	       fpu_madd_fState_S3$D_OUT[81:14],
	       !fpu_madd_fState_S3$D_OUT[151] && fpu_madd_fState_S3$D_OUT[13],
	       fpu_madd_fState_S3$D_OUT[151] ?
		 63'd0 :
		 IF_fpu_madd_fState_S3_first__995_BITS_12_TO_0__ETC___d2536,
	       x__h131406 } ;
  assign fpu_madd_fState_S4$ENQ = CAN_FIRE_RL_fpu_madd_s4_stage ;
  assign fpu_madd_fState_S4$DEQ = CAN_FIRE_RL_fpu_madd_s5_stage ;
  assign fpu_madd_fState_S4$CLR = 1'b0 ;
  // submodule fpu_madd_fState_S5
  assign fpu_madd_fState_S5$D_IN =
	     { fpu_madd_fState_S4$D_OUT[203:130],
	       fpu_madd_fState_S4$D_OUT[129] != fpu_madd_fState_S4$D_OUT[65],
	       NOT_fpu_madd_fState_S4_first__547_BIT_130_553__ETC___d2584 ?
		 fpu_madd_fState_S4$D_OUT[65] :
		 fpu_madd_fState_S4$D_OUT[129],
	       IF_NOT_fpu_madd_fState_S4_first__547_BIT_130_5_ETC___d2595 } ;
  assign fpu_madd_fState_S5$ENQ = CAN_FIRE_RL_fpu_madd_s5_stage ;
  assign fpu_madd_fState_S5$DEQ = CAN_FIRE_RL_fpu_madd_s6_stage ;
  assign fpu_madd_fState_S5$CLR = 1'b0 ;
  // submodule fpu_madd_fState_S6
  assign fpu_madd_fState_S6$D_IN =
	     { fpu_madd_fState_S5$D_OUT[215:127],
	       fpu_madd_fState_S5$D_OUT[113:57],
	       x__h132359 } ;
  assign fpu_madd_fState_S6$ENQ = CAN_FIRE_RL_fpu_madd_s6_stage ;
  assign fpu_madd_fState_S6$DEQ = CAN_FIRE_RL_fpu_madd_s7_stage ;
  assign fpu_madd_fState_S6$CLR = 1'b0 ;
  // submodule fpu_madd_fState_S7
  assign fpu_madd_fState_S7$D_IN =
	     { fpu_madd_fState_S6$D_OUT[202:114], x__h132871, x__h132880 } ;
  assign fpu_madd_fState_S7$ENQ = CAN_FIRE_RL_fpu_madd_s7_stage ;
  assign fpu_madd_fState_S7$DEQ = CAN_FIRE_RL_fpu_madd_s8_stage ;
  assign fpu_madd_fState_S7$CLR = 1'b0 ;
  // submodule fpu_madd_fState_S8
  assign fpu_madd_fState_S8$D_IN =
	     { fpu_madd_fState_S7$D_OUT[202:138],
	       fpu_madd_fState_S7$D_OUT[202] ?
		 fpu_madd_fState_S7$D_OUT[137:133] :
		 fpu_madd_fState_S7_first__651_BITS_137_TO_133__ETC___d2942,
	       fpu_madd_fState_S7$D_OUT[132:129],
	       !fpu_madd_fState_S7$D_OUT[202] &&
	       fpu_madd_fState_S7$D_OUT[127],
	       fpu_madd_fState_S7$D_OUT[202] ?
		 63'd0 :
		 IF_IF_fpu_madd_fState_S7_first__651_BIT_128_65_ETC___d2952,
	       x__h141760,
	       fpu_madd_fState_S7$D_OUT[128] } ;
  assign fpu_madd_fState_S8$ENQ = CAN_FIRE_RL_fpu_madd_s8_stage ;
  assign fpu_madd_fState_S8$DEQ = CAN_FIRE_RL_fpu_madd_s9_stage ;
  assign fpu_madd_fState_S8$CLR = 1'b0 ;
  // submodule fpu_sqr_fOperand_S0
  assign fpu_sqr_fOperand_S0$D_IN =
	     { IF_iFifo_first__087_BIT_201_115_THEN_IF_iFifo__ETC___d3848,
	       iFifo$D_OUT[6:4] } ;
  assign fpu_sqr_fOperand_S0$ENQ =
	     WILL_FIRE_RL_start_op && iFifo$D_OUT[3:0] == 4'd4 ;
  assign fpu_sqr_fOperand_S0$DEQ = CAN_FIRE_RL_fpu_sqr_s1_stage ;
  assign fpu_sqr_fOperand_S0$CLR = 1'b0 ;
  // submodule fpu_sqr_fResult_S5
  assign fpu_sqr_fResult_S5$D_IN =
	     fpu_sqr_fState_S4$D_OUT[138] ?
	       fpu_sqr_fState_S4$D_OUT[137:69] :
	       { (fpu_sqr_fState_S4$D_OUT[64:54] == 11'd2047) ?
		   fpu_sqr_fState_S4$D_OUT[65:2] :
		   CASE_fpu_sqr_fState_S4D_OUT_BITS_68_TO_66_0_C_ETC__q183,
		 fpu_sqr_fState_S4$D_OUT[73:69] |
		 { 2'd0,
		   _theResult___fst_exp__h95990 == 11'd2047 &&
		   _theResult___fst_sfd__h95991 == 52'd0,
		   1'd0,
		   fpu_sqr_fState_S4$D_OUT[64:54] != 11'd2047 &&
		   fpu_sqr_fState_S4$D_OUT[1:0] != 2'b0 } } ;
  assign fpu_sqr_fResult_S5$ENQ = CAN_FIRE_RL_fpu_sqr_s5_stage ;
  assign fpu_sqr_fResult_S5$DEQ = fpu_sqr_fResult_S5$EMPTY_N ;
  assign fpu_sqr_fResult_S5$CLR = 1'b0 ;
  // submodule fpu_sqr_fState_S1
  assign fpu_sqr_fState_S1$D_IN =
	     (fpu_sqr_fOperand_S0$D_OUT[65:55] == 11'd2047 &&
	      fpu_sqr_fOperand_S0$D_OUT[54:3] != 52'd0 &&
	      !fpu_sqr_fOperand_S0$D_OUT[54]) ?
	       { 1'd1,
		 fpu_sqr_fOperand_S0$D_OUT[66:55],
		 sfd__h45004,
		 130'h20AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA } :
	       IF_fpu_sqr_fOperand_S0_first__059_BITS_65_TO_5_ETC___d1212 ;
  assign fpu_sqr_fState_S1$ENQ = CAN_FIRE_RL_fpu_sqr_s1_stage ;
  assign fpu_sqr_fState_S1$DEQ = WILL_FIRE_RL_fpu_sqr_s2_stage ;
  assign fpu_sqr_fState_S1$CLR = 1'b0 ;
  // submodule fpu_sqr_fState_S2
  assign fpu_sqr_fState_S2$D_IN = fpu_sqr_fState_S1$D_OUT[194:58] ;
  assign fpu_sqr_fState_S2$ENQ = WILL_FIRE_RL_fpu_sqr_s2_stage ;
  assign fpu_sqr_fState_S2$DEQ = CAN_FIRE_RL_fpu_sqr_s3_stage ;
  assign fpu_sqr_fState_S2$CLR = 1'b0 ;
  // submodule fpu_sqr_fState_S3
  assign fpu_sqr_fState_S3$D_IN = { fpu_sqr_fState_S2$D_OUT, x__h86149 } ;
  assign fpu_sqr_fState_S3$ENQ = CAN_FIRE_RL_fpu_sqr_s3_stage ;
  assign fpu_sqr_fState_S3$DEQ = CAN_FIRE_RL_fpu_sqr_s4_stage ;
  assign fpu_sqr_fState_S3$CLR = 1'b0 ;
  // submodule fpu_sqr_fState_S4
  assign fpu_sqr_fState_S4$D_IN =
	     { fpu_sqr_fState_S3$D_OUT[195:131],
	       fpu_sqr_fState_S3$D_OUT[195] && fpu_sqr_fState_S3$D_OUT[130],
	       fpu_sqr_fState_S3$D_OUT[195] && fpu_sqr_fState_S3$D_OUT[129],
	       IF_fpu_sqr_fState_S3_first__375_BIT_195_376_TH_ETC___d1671,
	       fpu_sqr_fState_S3$D_OUT[125:122],
	       fpu_sqr_fState_S3$D_OUT[195] ?
		 fpu_sqr_fState_S3$D_OUT[121:59] :
		 IF_fpu_sqr_fState_S3_first__375_BIT_58_384_AND_ETC___d1678,
	       x__h95138 } ;
  assign fpu_sqr_fState_S4$ENQ = CAN_FIRE_RL_fpu_sqr_s4_stage ;
  assign fpu_sqr_fState_S4$DEQ = CAN_FIRE_RL_fpu_sqr_s5_stage ;
  assign fpu_sqr_fState_S4$CLR = 1'b0 ;
  // submodule iFifo
  assign iFifo$D_IN = server_core_request_put ;
  assign iFifo$ENQ = EN_server_core_request_put ;
  assign iFifo$DEQ = CAN_FIRE_RL_start_op ;
  assign iFifo$CLR = CAN_FIRE_RL_rl_reset ;
  // submodule isDoubleFifo
  assign isDoubleFifo$D_IN = !iFifo$D_OUT[201] ;
  assign isDoubleFifo$ENQ = CAN_FIRE_RL_start_op ;
  assign isDoubleFifo$DEQ = CAN_FIRE_RL_passResult ;
  assign isDoubleFifo$CLR = CAN_FIRE_RL_rl_reset ;
  // submodule isNegateFifo
  assign isNegateFifo$D_IN =
	     iFifo$D_OUT[3:0] == 4'd7 || iFifo$D_OUT[3:0] == 4'd8 ;
  assign isNegateFifo$ENQ = CAN_FIRE_RL_start_op ;
  assign isNegateFifo$DEQ = CAN_FIRE_RL_passResult ;
  assign isNegateFifo$CLR = CAN_FIRE_RL_rl_reset ;
  // submodule oFifo
  assign oFifo$D_IN =
	     { !isDoubleFifo$D_OUT,
	       IF_isDoubleFifo_first__407_THEN_IF_isNegateFif_ETC___d6657,
	       isDoubleFifo$D_OUT ?
		 resWire$wget[4:0] :
		 resWire_wget__410_BITS_4_TO_0_658_OR_NOT_resWi_ETC___d6768 } ;
  assign oFifo$ENQ = CAN_FIRE_RL_passResult ;
  assign oFifo$DEQ = EN_server_core_response_get ;
  assign oFifo$CLR = CAN_FIRE_RL_rl_reset ;
  // submodule resetReqsF
  assign resetReqsF$ENQ = EN_server_reset_request_put ;
  assign resetReqsF$DEQ = CAN_FIRE_RL_rl_reset ;
  assign resetReqsF$CLR = 1'b0 ;
  // submodule resetRspsF
  assign resetRspsF$ENQ = CAN_FIRE_RL_rl_reset ;
  assign resetRspsF$DEQ = EN_server_reset_response_get ;
  assign resetRspsF$CLR = 1'b0 ;
  // submodule rmdFifo
  assign rmdFifo$D_IN = iFifo$D_OUT[6:4] ;
  assign rmdFifo$ENQ = CAN_FIRE_RL_start_op ;
  assign rmdFifo$DEQ = CAN_FIRE_RL_passResult ;
  assign rmdFifo$CLR = CAN_FIRE_RL_rl_reset ;
  // remaining internal signals
  assign IF_0_CONCAT_IF_IF_0b0_CONCAT_NOT_resWire_wget__ETC__q133 =
	     _0_CONCAT_IF_IF_0b0_CONCAT_NOT_resWire_wget__41_ETC___d5769 ?
	       _theResult___snd__h277785 :
	       _theResult____h269613 ;
  assign IF_0_CONCAT_IF_IF_3074_MINUS_SEXT_iFifo_first__ETC__q37 =
	     _0_CONCAT_IF_IF_3074_MINUS_SEXT_iFifo_first__08_ETC___d3574 ?
	       _theResult___snd__h172913 :
	       _theResult____h164612 ;
  assign IF_0_CONCAT_IF_IF_3074_MINUS_SEXT_iFifo_first__ETC__q64 =
	     _0_CONCAT_IF_IF_3074_MINUS_SEXT_iFifo_first__08_ETC___d4282 ?
	       _theResult___snd__h250490 :
	       _theResult____h242189 ;
  assign IF_0_CONCAT_IF_IF_3074_MINUS_SEXT_iFifo_first__ETC__q97 =
	     _0_CONCAT_IF_IF_3074_MINUS_SEXT_iFifo_first__08_ETC___d5057 ?
	       _theResult___snd__h211551 :
	       _theResult____h203250 ;
  assign IF_0_CONCAT_IF_IF_3970_MINUS_SEXT_resWire_wget_ETC__q139 =
	     _0_CONCAT_IF_IF_3970_MINUS_SEXT_resWire_wget__4_ETC___d6280 ?
	       _theResult___snd__h295551 :
	       _theResult____h287250 ;
  assign IF_0_CONCAT_IF_IF_7170_MINUS_fpu_madd_fState_S_ETC__q24 =
	     _0_CONCAT_IF_IF_7170_MINUS_fpu_madd_fState_S3_f_ETC___d2463 ?
	       _theResult___snd__h131023 :
	       _theResult___snd__h131018 ;
  assign IF_0_CONCAT_IF_IF_fpu_div_fState_S3_first__16__ETC__q12 =
	     _0_CONCAT_IF_IF_fpu_div_fState_S3_first__16_BIT_ETC___d813 ?
	       _theResult___snd__h41460 :
	       _theResult___snd__h41455 ;
  assign IF_0_CONCAT_IF_IF_fpu_madd_fState_S7_first__65_ETC__q29 =
	     _0_CONCAT_IF_IF_fpu_madd_fState_S7_first__651_B_ETC___d2904 ?
	       _theResult___snd__h141449 :
	       _theResult___snd__h141444 ;
  assign IF_0_CONCAT_IF_fpu_sqr_fState_S3_first__375_BI_ETC__q19 =
	     _0_CONCAT_IF_fpu_sqr_fState_S3_first__375_BIT_5_ETC___d1633 ?
	       _theResult___snd__h94826 :
	       _theResult___snd__h94821 ;
  assign IF_0_CONCAT_IF_iFifo_first__087_BITS_102_TO_95_ETC__q100 =
	     _0_CONCAT_IF_iFifo_first__087_BITS_102_TO_95_62_ETC___d5107 ?
	       _theResult___snd__h201961 :
	       _theResult___snd__h220273 ;
  assign IF_0_CONCAT_IF_iFifo_first__087_BITS_102_TO_95_ETC__q93 =
	     _0_CONCAT_IF_iFifo_first__087_BITS_102_TO_95_62_ETC___d4759 ?
	       _theResult___snd__h201961 :
	       57'd0 ;
  assign IF_0_CONCAT_IF_iFifo_first__087_BITS_167_TO_16_ETC__q33 =
	     _0_CONCAT_IF_iFifo_first__087_BITS_167_TO_160_1_ETC___d3273 ?
	       _theResult___snd__h163323 :
	       57'd0 ;
  assign IF_0_CONCAT_IF_iFifo_first__087_BITS_167_TO_16_ETC__q40 =
	     _0_CONCAT_IF_iFifo_first__087_BITS_167_TO_160_1_ETC___d3624 ?
	       _theResult___snd__h163323 :
	       _theResult___snd__h181635 ;
  assign IF_0_CONCAT_IF_iFifo_first__087_BITS_37_TO_30__ETC__q60 =
	     _0_CONCAT_IF_iFifo_first__087_BITS_37_TO_30_850_ETC___d3984 ?
	       _theResult___snd__h240900 :
	       57'd0 ;
  assign IF_0_CONCAT_IF_iFifo_first__087_BITS_37_TO_30__ETC__q67 =
	     _0_CONCAT_IF_iFifo_first__087_BITS_37_TO_30_850_ETC___d4332 ?
	       _theResult___snd__h240900 :
	       _theResult___snd__h259212 ;
  assign IF_0_CONCAT_IF_resWire_wget__410_BITS_67_TO_57_ETC__q135 =
	     _0_CONCAT_IF_resWire_wget__410_BITS_67_TO_57_41_ETC___d5984 ?
	       _theResult___snd__h286367 :
	       57'd0 ;
  assign IF_0_CONCAT_IF_resWire_wget__410_BITS_67_TO_57_ETC__q142 =
	     _0_CONCAT_IF_resWire_wget__410_BITS_67_TO_57_41_ETC___d6333 ?
	       _theResult___snd__h286367 :
	       _theResult___snd__h304157 ;
  assign IF_0b0_CONCAT_NOT_fpu_div_fState_S4_first__73__ETC___d910 =
	     sfd__h42033[53] ?
	       ((fpu_div_fState_S4$D_OUT[64:54] == 11'd2046) ?
		  63'h7FF0000000000000 :
		  { din_inc___2_exp__h42617, sfd__h42033[52:1] }) :
	       { IF_fpu_div_fState_S4_first__73_BITS_64_TO_54_7_ETC___d907,
		 sfd__h42033[51:0] } ;
  assign IF_0b0_CONCAT_NOT_fpu_madd_fState_S8_first__96_ETC___d3065 =
	     sfd__h142040[53] ?
	       ((fpu_madd_fState_S8$D_OUT[65:55] == 11'd2046) ?
		  63'h7FF0000000000000 :
		  { din_inc___2_exp__h142626, sfd__h142040[52:1] }) :
	       { IF_fpu_madd_fState_S8_first__960_BITS_65_TO_55_ETC___d2986,
		 sfd__h142040[51:0] } ;
  assign IF_0b0_CONCAT_NOT_fpu_sqr_fState_S4_first__687_ETC___d1724 =
	     sfd__h95416[53] ?
	       ((fpu_sqr_fState_S4$D_OUT[64:54] == 11'd2046) ?
		  63'h7FF0000000000000 :
		  { din_inc___2_exp__h96000, sfd__h95416[52:1] }) :
	       { IF_fpu_sqr_fState_S4_first__687_BITS_64_TO_54__ETC___d1721,
		 sfd__h95416[51:0] } ;
  assign IF_3074_MINUS_0_CONCAT_IF_resWire_wget__410_BI_ETC___d6025 =
	     _3074_MINUS_0_CONCAT_IF_resWire_wget__410_BIT_5_ETC___d5533 ?
	       ((_theResult___fst_exp__h277722 == 8'd255) ?
		  !resWire$wget[68] :
		  IF_rmdFifo_first__778_EQ_0_779_THEN_IF_IF_IF_I_ETC___d5823) :
	       ((_theResult___fst_exp__h286378 == 8'd255) ?
		  !resWire$wget[68] :
		  IF_rmdFifo_first__778_EQ_0_779_THEN_IF_IF_IF_r_ETC___d6023) ;
  assign IF_3074_MINUS_0_CONCAT_IF_resWire_wget__410_BI_ETC___d6399 =
	     _3074_MINUS_0_CONCAT_IF_resWire_wget__410_BIT_5_ETC___d5533 ?
	       ((_theResult___fst_exp__h277722 == 8'd255) ?
		  resWire$wget[68] :
		  IF_rmdFifo_first__778_EQ_0_779_THEN_IF_IF_IF_I_ETC___d6388) :
	       ((_theResult___fst_exp__h286378 == 8'd255) ?
		  resWire$wget[68] :
		  IF_rmdFifo_first__778_EQ_0_779_THEN_IF_IF_IF_r_ETC___d6397) ;
  assign IF_3970_MINUS_0_CONCAT_IF_iFifo_first__087_BIT_ETC___d3317 =
	     _3970_MINUS_0_CONCAT_IF_iFifo_first__087_BIT_15_ETC___d3190 ?
	       (iFifo$D_OUT[6:4] == 3'd0 || iFifo$D_OUT[6:4] == 3'd1 ||
		iFifo$D_OUT[6:4] == 3'd2 ||
		iFifo$D_OUT[6:4] == 3'd3 ||
		iFifo$D_OUT[6:4] == 3'd4) &&
	       iFifo$D_OUT[168] :
	       ((_theResult___fst_exp__h163334 == 11'd2047) ?
		  iFifo$D_OUT[168] :
		  CASE_iFifoD_OUT_BITS_6_TO_4_0_CASE_guard55373_ETC__q55) ;
  assign IF_3970_MINUS_0_CONCAT_IF_iFifo_first__087_BIT_ETC___d4027 =
	     _3970_MINUS_0_CONCAT_IF_iFifo_first__087_BIT_29_ETC___d3910 ?
	       (iFifo$D_OUT[6:4] == 3'd0 || iFifo$D_OUT[6:4] == 3'd1 ||
		iFifo$D_OUT[6:4] == 3'd2 ||
		iFifo$D_OUT[6:4] == 3'd3 ||
		iFifo$D_OUT[6:4] == 3'd4) &&
	       iFifo$D_OUT[38] :
	       ((_theResult___fst_exp__h240911 == 11'd2047) ?
		  iFifo$D_OUT[38] :
		  CASE_iFifoD_OUT_BITS_6_TO_4_0_CASE_guard32950_ETC__q80) ;
  assign IF_3970_MINUS_0_CONCAT_IF_iFifo_first__087_BIT_ETC___d4581 =
	     _3970_MINUS_0_CONCAT_IF_iFifo_first__087_BIT_29_ETC___d3910 ?
	       iFifo$D_OUT[6:4] != 3'd0 && iFifo$D_OUT[6:4] != 3'd1 &&
	       iFifo$D_OUT[6:4] != 3'd2 &&
	       iFifo$D_OUT[6:4] != 3'd3 &&
	       iFifo$D_OUT[6:4] != 3'd4 ||
	       !iFifo$D_OUT[38] :
	       ((_theResult___fst_exp__h240911 == 11'd2047) ?
		  !iFifo$D_OUT[38] :
		  CASE_iFifoD_OUT_BITS_6_TO_4_0_CASE_guard32950_ETC__q88) ;
  assign IF_3970_MINUS_0_CONCAT_IF_iFifo_first__087_BIT_ETC___d4802 =
	     _3970_MINUS_0_CONCAT_IF_iFifo_first__087_BIT_94_ETC___d4685 ?
	       (iFifo$D_OUT[6:4] == 3'd0 || iFifo$D_OUT[6:4] == 3'd1 ||
		iFifo$D_OUT[6:4] == 3'd2 ||
		iFifo$D_OUT[6:4] == 3'd3 ||
		iFifo$D_OUT[6:4] == 3'd4) &&
	       iFifo$D_OUT[103] :
	       ((_theResult___fst_exp__h201972 == 11'd2047) ?
		  iFifo$D_OUT[103] :
		  CASE_iFifoD_OUT_BITS_6_TO_4_0_CASE_guard94011_ETC__q115) ;
  assign IF_3970_MINUS_0_CONCAT_IF_iFifo_first__087_BIT_ETC___d5347 =
	     _3970_MINUS_0_CONCAT_IF_iFifo_first__087_BIT_94_ETC___d4685 ?
	       iFifo$D_OUT[6:4] != 3'd0 && iFifo$D_OUT[6:4] != 3'd1 &&
	       iFifo$D_OUT[6:4] != 3'd2 &&
	       iFifo$D_OUT[6:4] != 3'd3 &&
	       iFifo$D_OUT[6:4] != 3'd4 ||
	       !iFifo$D_OUT[103] :
	       ((_theResult___fst_exp__h201972 == 11'd2047) ?
		  !iFifo$D_OUT[103] :
		  CASE_iFifoD_OUT_BITS_6_TO_4_0_CASE_guard94011_ETC__q121) ;
  assign IF_IF_0b0_CONCAT_NOT_resWire_wget__410_BITS_67_ETC___d5767 =
	     (_theResult____h269613[56] ?
		6'd0 :
		(_theResult____h269613[55] ?
		   6'd1 :
		   (_theResult____h269613[54] ?
		      6'd2 :
		      (_theResult____h269613[53] ?
			 6'd3 :
			 (_theResult____h269613[52] ?
			    6'd4 :
			    (_theResult____h269613[51] ?
			       6'd5 :
			       (_theResult____h269613[50] ?
				  6'd6 :
				  (_theResult____h269613[49] ?
				     6'd7 :
				     (_theResult____h269613[48] ?
					6'd8 :
					(_theResult____h269613[47] ?
					   6'd9 :
					   (_theResult____h269613[46] ?
					      6'd10 :
					      (_theResult____h269613[45] ?
						 6'd11 :
						 (_theResult____h269613[44] ?
						    6'd12 :
						    (_theResult____h269613[43] ?
						       6'd13 :
						       (_theResult____h269613[42] ?
							  6'd14 :
							  (_theResult____h269613[41] ?
							     6'd15 :
							     (_theResult____h269613[40] ?
								6'd16 :
								(_theResult____h269613[39] ?
								   6'd17 :
								   (_theResult____h269613[38] ?
								      6'd18 :
								      (_theResult____h269613[37] ?
									 6'd19 :
									 (_theResult____h269613[36] ?
									    6'd20 :
									    (_theResult____h269613[35] ?
									       6'd21 :
									       (_theResult____h269613[34] ?
										  6'd22 :
										  (_theResult____h269613[33] ?
										     6'd23 :
										     (_theResult____h269613[32] ?
											6'd24 :
											(_theResult____h269613[31] ?
											   6'd25 :
											   (_theResult____h269613[30] ?
											      6'd26 :
											      (_theResult____h269613[29] ?
												 6'd27 :
												 (_theResult____h269613[28] ?
												    6'd28 :
												    (_theResult____h269613[27] ?
												       6'd29 :
												       (_theResult____h269613[26] ?
													  6'd30 :
													  (_theResult____h269613[25] ?
													     6'd31 :
													     (_theResult____h269613[24] ?
														6'd32 :
														(_theResult____h269613[23] ?
														   6'd33 :
														   (_theResult____h269613[22] ?
														      6'd34 :
														      (_theResult____h269613[21] ?
															 6'd35 :
															 (_theResult____h269613[20] ?
															    6'd36 :
															    (_theResult____h269613[19] ?
															       6'd37 :
															       (_theResult____h269613[18] ?
																  6'd38 :
																  (_theResult____h269613[17] ?
																     6'd39 :
																     (_theResult____h269613[16] ?
																	6'd40 :
																	(_theResult____h269613[15] ?
																	   6'd41 :
																	   (_theResult____h269613[14] ?
																	      6'd42 :
																	      (_theResult____h269613[13] ?
																		 6'd43 :
																		 (_theResult____h269613[12] ?
																		    6'd44 :
																		    (_theResult____h269613[11] ?
																		       6'd45 :
																		       (_theResult____h269613[10] ?
																			  6'd46 :
																			  (_theResult____h269613[9] ?
																			     6'd47 :
																			     (_theResult____h269613[8] ?
																				6'd48 :
																				(_theResult____h269613[7] ?
																				   6'd49 :
																				   (_theResult____h269613[6] ?
																				      6'd50 :
																				      (_theResult____h269613[5] ?
																					 6'd51 :
																					 (_theResult____h269613[4] ?
																					    6'd52 :
																					    (_theResult____h269613[3] ?
																					       6'd53 :
																					       (_theResult____h269613[2] ?
																						  6'd54 :
																						  (_theResult____h269613[1] ?
																						     6'd55 :
																						     (_theResult____h269613[0] ?
																							6'd56 :
																							6'd57))))))))))))))))))))))))))))))))))))))))))))))))))))))))) -
	     6'd1 ;
  assign IF_IF_3074_MINUS_SEXT_iFifo_first__087_BITS_10_ETC___d5055 =
	     (_theResult____h203250[56] ?
		6'd0 :
		(_theResult____h203250[55] ?
		   6'd1 :
		   (_theResult____h203250[54] ?
		      6'd2 :
		      (_theResult____h203250[53] ?
			 6'd3 :
			 (_theResult____h203250[52] ?
			    6'd4 :
			    (_theResult____h203250[51] ?
			       6'd5 :
			       (_theResult____h203250[50] ?
				  6'd6 :
				  (_theResult____h203250[49] ?
				     6'd7 :
				     (_theResult____h203250[48] ?
					6'd8 :
					(_theResult____h203250[47] ?
					   6'd9 :
					   (_theResult____h203250[46] ?
					      6'd10 :
					      (_theResult____h203250[45] ?
						 6'd11 :
						 (_theResult____h203250[44] ?
						    6'd12 :
						    (_theResult____h203250[43] ?
						       6'd13 :
						       (_theResult____h203250[42] ?
							  6'd14 :
							  (_theResult____h203250[41] ?
							     6'd15 :
							     (_theResult____h203250[40] ?
								6'd16 :
								(_theResult____h203250[39] ?
								   6'd17 :
								   (_theResult____h203250[38] ?
								      6'd18 :
								      (_theResult____h203250[37] ?
									 6'd19 :
									 (_theResult____h203250[36] ?
									    6'd20 :
									    (_theResult____h203250[35] ?
									       6'd21 :
									       (_theResult____h203250[34] ?
										  6'd22 :
										  (_theResult____h203250[33] ?
										     6'd23 :
										     (_theResult____h203250[32] ?
											6'd24 :
											(_theResult____h203250[31] ?
											   6'd25 :
											   (_theResult____h203250[30] ?
											      6'd26 :
											      (_theResult____h203250[29] ?
												 6'd27 :
												 (_theResult____h203250[28] ?
												    6'd28 :
												    (_theResult____h203250[27] ?
												       6'd29 :
												       (_theResult____h203250[26] ?
													  6'd30 :
													  (_theResult____h203250[25] ?
													     6'd31 :
													     (_theResult____h203250[24] ?
														6'd32 :
														(_theResult____h203250[23] ?
														   6'd33 :
														   (_theResult____h203250[22] ?
														      6'd34 :
														      (_theResult____h203250[21] ?
															 6'd35 :
															 (_theResult____h203250[20] ?
															    6'd36 :
															    (_theResult____h203250[19] ?
															       6'd37 :
															       (_theResult____h203250[18] ?
																  6'd38 :
																  (_theResult____h203250[17] ?
																     6'd39 :
																     (_theResult____h203250[16] ?
																	6'd40 :
																	(_theResult____h203250[15] ?
																	   6'd41 :
																	   (_theResult____h203250[14] ?
																	      6'd42 :
																	      (_theResult____h203250[13] ?
																		 6'd43 :
																		 (_theResult____h203250[12] ?
																		    6'd44 :
																		    (_theResult____h203250[11] ?
																		       6'd45 :
																		       (_theResult____h203250[10] ?
																			  6'd46 :
																			  (_theResult____h203250[9] ?
																			     6'd47 :
																			     (_theResult____h203250[8] ?
																				6'd48 :
																				(_theResult____h203250[7] ?
																				   6'd49 :
																				   (_theResult____h203250[6] ?
																				      6'd50 :
																				      (_theResult____h203250[5] ?
																					 6'd51 :
																					 (_theResult____h203250[4] ?
																					    6'd52 :
																					    (_theResult____h203250[3] ?
																					       6'd53 :
																					       (_theResult____h203250[2] ?
																						  6'd54 :
																						  (_theResult____h203250[1] ?
																						     6'd55 :
																						     (_theResult____h203250[0] ?
																							6'd56 :
																							6'd57))))))))))))))))))))))))))))))))))))))))))))))))))))))))) -
	     6'd1 ;
  assign IF_IF_3074_MINUS_SEXT_iFifo_first__087_BITS_16_ETC___d3572 =
	     (_theResult____h164612[56] ?
		6'd0 :
		(_theResult____h164612[55] ?
		   6'd1 :
		   (_theResult____h164612[54] ?
		      6'd2 :
		      (_theResult____h164612[53] ?
			 6'd3 :
			 (_theResult____h164612[52] ?
			    6'd4 :
			    (_theResult____h164612[51] ?
			       6'd5 :
			       (_theResult____h164612[50] ?
				  6'd6 :
				  (_theResult____h164612[49] ?
				     6'd7 :
				     (_theResult____h164612[48] ?
					6'd8 :
					(_theResult____h164612[47] ?
					   6'd9 :
					   (_theResult____h164612[46] ?
					      6'd10 :
					      (_theResult____h164612[45] ?
						 6'd11 :
						 (_theResult____h164612[44] ?
						    6'd12 :
						    (_theResult____h164612[43] ?
						       6'd13 :
						       (_theResult____h164612[42] ?
							  6'd14 :
							  (_theResult____h164612[41] ?
							     6'd15 :
							     (_theResult____h164612[40] ?
								6'd16 :
								(_theResult____h164612[39] ?
								   6'd17 :
								   (_theResult____h164612[38] ?
								      6'd18 :
								      (_theResult____h164612[37] ?
									 6'd19 :
									 (_theResult____h164612[36] ?
									    6'd20 :
									    (_theResult____h164612[35] ?
									       6'd21 :
									       (_theResult____h164612[34] ?
										  6'd22 :
										  (_theResult____h164612[33] ?
										     6'd23 :
										     (_theResult____h164612[32] ?
											6'd24 :
											(_theResult____h164612[31] ?
											   6'd25 :
											   (_theResult____h164612[30] ?
											      6'd26 :
											      (_theResult____h164612[29] ?
												 6'd27 :
												 (_theResult____h164612[28] ?
												    6'd28 :
												    (_theResult____h164612[27] ?
												       6'd29 :
												       (_theResult____h164612[26] ?
													  6'd30 :
													  (_theResult____h164612[25] ?
													     6'd31 :
													     (_theResult____h164612[24] ?
														6'd32 :
														(_theResult____h164612[23] ?
														   6'd33 :
														   (_theResult____h164612[22] ?
														      6'd34 :
														      (_theResult____h164612[21] ?
															 6'd35 :
															 (_theResult____h164612[20] ?
															    6'd36 :
															    (_theResult____h164612[19] ?
															       6'd37 :
															       (_theResult____h164612[18] ?
																  6'd38 :
																  (_theResult____h164612[17] ?
																     6'd39 :
																     (_theResult____h164612[16] ?
																	6'd40 :
																	(_theResult____h164612[15] ?
																	   6'd41 :
																	   (_theResult____h164612[14] ?
																	      6'd42 :
																	      (_theResult____h164612[13] ?
																		 6'd43 :
																		 (_theResult____h164612[12] ?
																		    6'd44 :
																		    (_theResult____h164612[11] ?
																		       6'd45 :
																		       (_theResult____h164612[10] ?
																			  6'd46 :
																			  (_theResult____h164612[9] ?
																			     6'd47 :
																			     (_theResult____h164612[8] ?
																				6'd48 :
																				(_theResult____h164612[7] ?
																				   6'd49 :
																				   (_theResult____h164612[6] ?
																				      6'd50 :
																				      (_theResult____h164612[5] ?
																					 6'd51 :
																					 (_theResult____h164612[4] ?
																					    6'd52 :
																					    (_theResult____h164612[3] ?
																					       6'd53 :
																					       (_theResult____h164612[2] ?
																						  6'd54 :
																						  (_theResult____h164612[1] ?
																						     6'd55 :
																						     (_theResult____h164612[0] ?
																							6'd56 :
																							6'd57))))))))))))))))))))))))))))))))))))))))))))))))))))))))) -
	     6'd1 ;
  assign IF_IF_3074_MINUS_SEXT_iFifo_first__087_BITS_37_ETC___d4280 =
	     (_theResult____h242189[56] ?
		6'd0 :
		(_theResult____h242189[55] ?
		   6'd1 :
		   (_theResult____h242189[54] ?
		      6'd2 :
		      (_theResult____h242189[53] ?
			 6'd3 :
			 (_theResult____h242189[52] ?
			    6'd4 :
			    (_theResult____h242189[51] ?
			       6'd5 :
			       (_theResult____h242189[50] ?
				  6'd6 :
				  (_theResult____h242189[49] ?
				     6'd7 :
				     (_theResult____h242189[48] ?
					6'd8 :
					(_theResult____h242189[47] ?
					   6'd9 :
					   (_theResult____h242189[46] ?
					      6'd10 :
					      (_theResult____h242189[45] ?
						 6'd11 :
						 (_theResult____h242189[44] ?
						    6'd12 :
						    (_theResult____h242189[43] ?
						       6'd13 :
						       (_theResult____h242189[42] ?
							  6'd14 :
							  (_theResult____h242189[41] ?
							     6'd15 :
							     (_theResult____h242189[40] ?
								6'd16 :
								(_theResult____h242189[39] ?
								   6'd17 :
								   (_theResult____h242189[38] ?
								      6'd18 :
								      (_theResult____h242189[37] ?
									 6'd19 :
									 (_theResult____h242189[36] ?
									    6'd20 :
									    (_theResult____h242189[35] ?
									       6'd21 :
									       (_theResult____h242189[34] ?
										  6'd22 :
										  (_theResult____h242189[33] ?
										     6'd23 :
										     (_theResult____h242189[32] ?
											6'd24 :
											(_theResult____h242189[31] ?
											   6'd25 :
											   (_theResult____h242189[30] ?
											      6'd26 :
											      (_theResult____h242189[29] ?
												 6'd27 :
												 (_theResult____h242189[28] ?
												    6'd28 :
												    (_theResult____h242189[27] ?
												       6'd29 :
												       (_theResult____h242189[26] ?
													  6'd30 :
													  (_theResult____h242189[25] ?
													     6'd31 :
													     (_theResult____h242189[24] ?
														6'd32 :
														(_theResult____h242189[23] ?
														   6'd33 :
														   (_theResult____h242189[22] ?
														      6'd34 :
														      (_theResult____h242189[21] ?
															 6'd35 :
															 (_theResult____h242189[20] ?
															    6'd36 :
															    (_theResult____h242189[19] ?
															       6'd37 :
															       (_theResult____h242189[18] ?
																  6'd38 :
																  (_theResult____h242189[17] ?
																     6'd39 :
																     (_theResult____h242189[16] ?
																	6'd40 :
																	(_theResult____h242189[15] ?
																	   6'd41 :
																	   (_theResult____h242189[14] ?
																	      6'd42 :
																	      (_theResult____h242189[13] ?
																		 6'd43 :
																		 (_theResult____h242189[12] ?
																		    6'd44 :
																		    (_theResult____h242189[11] ?
																		       6'd45 :
																		       (_theResult____h242189[10] ?
																			  6'd46 :
																			  (_theResult____h242189[9] ?
																			     6'd47 :
																			     (_theResult____h242189[8] ?
																				6'd48 :
																				(_theResult____h242189[7] ?
																				   6'd49 :
																				   (_theResult____h242189[6] ?
																				      6'd50 :
																				      (_theResult____h242189[5] ?
																					 6'd51 :
																					 (_theResult____h242189[4] ?
																					    6'd52 :
																					    (_theResult____h242189[3] ?
																					       6'd53 :
																					       (_theResult____h242189[2] ?
																						  6'd54 :
																						  (_theResult____h242189[1] ?
																						     6'd55 :
																						     (_theResult____h242189[0] ?
																							6'd56 :
																							6'd57))))))))))))))))))))))))))))))))))))))))))))))))))))))))) -
	     6'd1 ;
  assign IF_IF_3970_MINUS_SEXT_resWire_wget__410_BITS_6_ETC___d6278 =
	     (_theResult____h287250[56] ?
		6'd0 :
		(_theResult____h287250[55] ?
		   6'd1 :
		   (_theResult____h287250[54] ?
		      6'd2 :
		      (_theResult____h287250[53] ?
			 6'd3 :
			 (_theResult____h287250[52] ?
			    6'd4 :
			    (_theResult____h287250[51] ?
			       6'd5 :
			       (_theResult____h287250[50] ?
				  6'd6 :
				  (_theResult____h287250[49] ?
				     6'd7 :
				     (_theResult____h287250[48] ?
					6'd8 :
					(_theResult____h287250[47] ?
					   6'd9 :
					   (_theResult____h287250[46] ?
					      6'd10 :
					      (_theResult____h287250[45] ?
						 6'd11 :
						 (_theResult____h287250[44] ?
						    6'd12 :
						    (_theResult____h287250[43] ?
						       6'd13 :
						       (_theResult____h287250[42] ?
							  6'd14 :
							  (_theResult____h287250[41] ?
							     6'd15 :
							     (_theResult____h287250[40] ?
								6'd16 :
								(_theResult____h287250[39] ?
								   6'd17 :
								   (_theResult____h287250[38] ?
								      6'd18 :
								      (_theResult____h287250[37] ?
									 6'd19 :
									 (_theResult____h287250[36] ?
									    6'd20 :
									    (_theResult____h287250[35] ?
									       6'd21 :
									       (_theResult____h287250[34] ?
										  6'd22 :
										  (_theResult____h287250[33] ?
										     6'd23 :
										     (_theResult____h287250[32] ?
											6'd24 :
											(_theResult____h287250[31] ?
											   6'd25 :
											   (_theResult____h287250[30] ?
											      6'd26 :
											      (_theResult____h287250[29] ?
												 6'd27 :
												 (_theResult____h287250[28] ?
												    6'd28 :
												    (_theResult____h287250[27] ?
												       6'd29 :
												       (_theResult____h287250[26] ?
													  6'd30 :
													  (_theResult____h287250[25] ?
													     6'd31 :
													     (_theResult____h287250[24] ?
														6'd32 :
														(_theResult____h287250[23] ?
														   6'd33 :
														   (_theResult____h287250[22] ?
														      6'd34 :
														      (_theResult____h287250[21] ?
															 6'd35 :
															 (_theResult____h287250[20] ?
															    6'd36 :
															    (_theResult____h287250[19] ?
															       6'd37 :
															       (_theResult____h287250[18] ?
																  6'd38 :
																  (_theResult____h287250[17] ?
																     6'd39 :
																     (_theResult____h287250[16] ?
																	6'd40 :
																	(_theResult____h287250[15] ?
																	   6'd41 :
																	   (_theResult____h287250[14] ?
																	      6'd42 :
																	      (_theResult____h287250[13] ?
																		 6'd43 :
																		 (_theResult____h287250[12] ?
																		    6'd44 :
																		    (_theResult____h287250[11] ?
																		       6'd45 :
																		       (_theResult____h287250[10] ?
																			  6'd46 :
																			  (_theResult____h287250[9] ?
																			     6'd47 :
																			     (_theResult____h287250[8] ?
																				6'd48 :
																				(_theResult____h287250[7] ?
																				   6'd49 :
																				   (_theResult____h287250[6] ?
																				      6'd50 :
																				      (_theResult____h287250[5] ?
																					 6'd51 :
																					 (_theResult____h287250[4] ?
																					    6'd52 :
																					    (_theResult____h287250[3] ?
																					       6'd53 :
																					       (_theResult____h287250[2] ?
																						  6'd54 :
																						  (_theResult____h287250[1] ?
																						     6'd55 :
																						     (_theResult____h287250[0] ?
																							6'd56 :
																							6'd57))))))))))))))))))))))))))))))))))))))))))))))))))))))))) -
	     6'd1 ;
  assign IF_IF_7170_MINUS_fpu_madd_fState_S3_first__995_ETC___d2031 =
	     (din_exp__h130866 == 11'd0) ?
	       12'd3074 :
	       { din_exp30866_MINUS_1023__q23[10],
		 din_exp30866_MINUS_1023__q23 } ;
  assign IF_IF_7170_MINUS_fpu_madd_fState_S3_first__995_ETC___d2460 =
	     (sfdBC__h115662[105] ?
		7'd0 :
		(sfdBC__h115662[104] ?
		   7'd1 :
		   (sfdBC__h115662[103] ?
		      7'd2 :
		      (sfdBC__h115662[102] ?
			 7'd3 :
			 (sfdBC__h115662[101] ?
			    7'd4 :
			    (sfdBC__h115662[100] ?
			       7'd5 :
			       (sfdBC__h115662[99] ?
				  7'd6 :
				  (sfdBC__h115662[98] ?
				     7'd7 :
				     (sfdBC__h115662[97] ?
					7'd8 :
					(sfdBC__h115662[96] ?
					   7'd9 :
					   (sfdBC__h115662[95] ?
					      7'd10 :
					      (sfdBC__h115662[94] ?
						 7'd11 :
						 (sfdBC__h115662[93] ?
						    7'd12 :
						    (sfdBC__h115662[92] ?
						       7'd13 :
						       (sfdBC__h115662[91] ?
							  7'd14 :
							  (sfdBC__h115662[90] ?
							     7'd15 :
							     (sfdBC__h115662[89] ?
								7'd16 :
								(sfdBC__h115662[88] ?
								   7'd17 :
								   (sfdBC__h115662[87] ?
								      7'd18 :
								      (sfdBC__h115662[86] ?
									 7'd19 :
									 (sfdBC__h115662[85] ?
									    7'd20 :
									    (sfdBC__h115662[84] ?
									       7'd21 :
									       (sfdBC__h115662[83] ?
										  7'd22 :
										  (sfdBC__h115662[82] ?
										     7'd23 :
										     (sfdBC__h115662[81] ?
											7'd24 :
											(sfdBC__h115662[80] ?
											   7'd25 :
											   (sfdBC__h115662[79] ?
											      7'd26 :
											      (sfdBC__h115662[78] ?
												 7'd27 :
												 (sfdBC__h115662[77] ?
												    7'd28 :
												    (sfdBC__h115662[76] ?
												       7'd29 :
												       (sfdBC__h115662[75] ?
													  7'd30 :
													  (sfdBC__h115662[74] ?
													     7'd31 :
													     (sfdBC__h115662[73] ?
														7'd32 :
														(sfdBC__h115662[72] ?
														   7'd33 :
														   (sfdBC__h115662[71] ?
														      7'd34 :
														      (sfdBC__h115662[70] ?
															 7'd35 :
															 (sfdBC__h115662[69] ?
															    7'd36 :
															    (sfdBC__h115662[68] ?
															       7'd37 :
															       (sfdBC__h115662[67] ?
																  7'd38 :
																  (sfdBC__h115662[66] ?
																     7'd39 :
																     (sfdBC__h115662[65] ?
																	7'd40 :
																	(sfdBC__h115662[64] ?
																	   7'd41 :
																	   (sfdBC__h115662[63] ?
																	      7'd42 :
																	      (sfdBC__h115662[62] ?
																		 7'd43 :
																		 (sfdBC__h115662[61] ?
																		    7'd44 :
																		    (sfdBC__h115662[60] ?
																		       7'd45 :
																		       (sfdBC__h115662[59] ?
																			  7'd46 :
																			  (sfdBC__h115662[58] ?
																			     7'd47 :
																			     (sfdBC__h115662[57] ?
																				7'd48 :
																				(sfdBC__h115662[56] ?
																				   7'd49 :
																				   (sfdBC__h115662[55] ?
																				      7'd50 :
																				      (sfdBC__h115662[54] ?
																					 7'd51 :
																					 (sfdBC__h115662[53] ?
																					    7'd52 :
																					    (sfdBC__h115662[52] ?
																					       7'd53 :
																					       (sfdBC__h115662[51] ?
																						  7'd54 :
																						  (sfdBC__h115662[50] ?
																						     7'd55 :
																						     (sfdBC__h115662[49] ?
																							7'd56 :
																							(sfdBC__h115662[48] ?
																							   7'd57 :
																							   (sfdBC__h115662[47] ?
																							      7'd58 :
																							      (sfdBC__h115662[46] ?
																								 7'd59 :
																								 (sfdBC__h115662[45] ?
																								    7'd60 :
																								    (sfdBC__h115662[44] ?
																								       7'd61 :
																								       (sfdBC__h115662[43] ?
																									  7'd62 :
																									  (sfdBC__h115662[42] ?
																									     7'd63 :
																									     (sfdBC__h115662[41] ?
																										7'd64 :
																										(sfdBC__h115662[40] ?
																										   7'd65 :
																										   (sfdBC__h115662[39] ?
																										      7'd66 :
																										      (sfdBC__h115662[38] ?
																											 7'd67 :
																											 (sfdBC__h115662[37] ?
																											    7'd68 :
																											    (sfdBC__h115662[36] ?
																											       7'd69 :
																											       (sfdBC__h115662[35] ?
																												  7'd70 :
																												  (sfdBC__h115662[34] ?
																												     7'd71 :
																												     (sfdBC__h115662[33] ?
																													7'd72 :
																													(sfdBC__h115662[32] ?
																													   7'd73 :
																													   (sfdBC__h115662[31] ?
																													      7'd74 :
																													      (sfdBC__h115662[30] ?
																														 7'd75 :
																														 (sfdBC__h115662[29] ?
																														    7'd76 :
																														    (sfdBC__h115662[28] ?
																														       7'd77 :
																														       (sfdBC__h115662[27] ?
																															  7'd78 :
																															  (sfdBC__h115662[26] ?
																															     7'd79 :
																															     (sfdBC__h115662[25] ?
																																7'd80 :
																																(sfdBC__h115662[24] ?
																																   7'd81 :
																																   (sfdBC__h115662[23] ?
																																      7'd82 :
																																      (sfdBC__h115662[22] ?
																																	 7'd83 :
																																	 (sfdBC__h115662[21] ?
																																	    7'd84 :
																																	    (sfdBC__h115662[20] ?
																																	       7'd85 :
																																	       (sfdBC__h115662[19] ?
																																		  7'd86 :
																																		  (sfdBC__h115662[18] ?
																																		     7'd87 :
																																		     (sfdBC__h115662[17] ?
																																			7'd88 :
																																			(sfdBC__h115662[16] ?
																																			   7'd89 :
																																			   (sfdBC__h115662[15] ?
																																			      7'd90 :
																																			      (sfdBC__h115662[14] ?
																																				 7'd91 :
																																				 (sfdBC__h115662[13] ?
																																				    7'd92 :
																																				    (sfdBC__h115662[12] ?
																																				       7'd93 :
																																				       (sfdBC__h115662[11] ?
																																					  7'd94 :
																																					  (sfdBC__h115662[10] ?
																																					     7'd95 :
																																					     (sfdBC__h115662[9] ?
																																						7'd96 :
																																						(sfdBC__h115662[8] ?
																																						   7'd97 :
																																						   (sfdBC__h115662[7] ?
																																						      7'd98 :
																																						      (sfdBC__h115662[6] ?
																																							 7'd99 :
																																							 (sfdBC__h115662[5] ?
																																							    7'd100 :
																																							    (sfdBC__h115662[4] ?
																																							       7'd101 :
																																							       (sfdBC__h115662[3] ?
																																								  7'd102 :
																																								  (sfdBC__h115662[2] ?
																																								     7'd103 :
																																								     (sfdBC__h115662[1] ?
																																									7'd104 :
																																									(sfdBC__h115662[0] ?
																																									   7'd105 :
																																									   7'd106)))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) -
	     7'd1 ;
  assign IF_IF_7170_MINUS_fpu_madd_fState_S3_first__995_ETC___d2462 =
	     IF_IF_7170_MINUS_fpu_madd_fState_S3_first__995_ETC___d2031 -
	     12'd3074 ;
  assign IF_IF_7170_MINUS_fpu_madd_fState_S3_first__995_ETC___d2534 =
	     (sfdBC__h115662[105] &&
	      IF_IF_7170_MINUS_fpu_madd_fState_S3_first__995_ETC___d2031 ==
	      12'd1023) ?
	       63'h7FEFFFFFFFFFFFFF :
	       { _theResult___fst_exp__h130949, sfdin__h130943[105:54] } ;
  assign IF_IF_IF_IF_0b0_CONCAT_NOT_resWire_wget__410_B_ETC___d6448 =
	     (guard__h269623 == 2'b0 || resWire$wget[68]) ?
	       _theResult___fst_exp__h277722 :
	       _theResult___exp__h278238 ;
  assign IF_IF_IF_IF_0b0_CONCAT_NOT_resWire_wget__410_B_ETC___d6450 =
	     (guard__h269623 == 2'b0) ?
	       _theResult___fst_exp__h277722 :
	       (resWire$wget[68] ?
		  _theResult___exp__h278238 :
		  _theResult___fst_exp__h277722) ;
  assign IF_IF_IF_IF_0b0_CONCAT_NOT_resWire_wget__410_B_ETC___d6576 =
	     (guard__h269623 == 2'b0 || resWire$wget[68]) ?
	       sfdin__h277716[56:34] :
	       _theResult___sfd__h278239 ;
  assign IF_IF_IF_IF_0b0_CONCAT_NOT_resWire_wget__410_B_ETC___d6578 =
	     (guard__h269623 == 2'b0) ?
	       sfdin__h277716[56:34] :
	       (resWire$wget[68] ?
		  _theResult___sfd__h278239 :
		  sfdin__h277716[56:34]) ;
  assign IF_IF_IF_IF_3074_MINUS_SEXT_iFifo_first__087_B_ETC___d3729 =
	     (guard__h164622 == 2'b0 || iFifo$D_OUT[168]) ?
	       _theResult___fst_exp__h172850 :
	       _theResult___exp__h173569 ;
  assign IF_IF_IF_IF_3074_MINUS_SEXT_iFifo_first__087_B_ETC___d3731 =
	     (guard__h164622 == 2'b0) ?
	       _theResult___fst_exp__h172850 :
	       (iFifo$D_OUT[168] ?
		  _theResult___exp__h173569 :
		  _theResult___fst_exp__h172850) ;
  assign IF_IF_IF_IF_3074_MINUS_SEXT_iFifo_first__087_B_ETC___d3813 =
	     (guard__h164622 == 2'b0 || iFifo$D_OUT[168]) ?
	       sfdin__h172844[56:5] :
	       _theResult___sfd__h173570 ;
  assign IF_IF_IF_IF_3074_MINUS_SEXT_iFifo_first__087_B_ETC___d3815 =
	     (guard__h164622 == 2'b0) ?
	       sfdin__h172844[56:5] :
	       (iFifo$D_OUT[168] ?
		  _theResult___sfd__h173570 :
		  sfdin__h172844[56:5]) ;
  assign IF_IF_IF_IF_3074_MINUS_SEXT_iFifo_first__087_B_ETC___d4436 =
	     (guard__h242199 == 2'b0 || iFifo$D_OUT[38]) ?
	       _theResult___fst_exp__h250427 :
	       _theResult___exp__h251146 ;
  assign IF_IF_IF_IF_3074_MINUS_SEXT_iFifo_first__087_B_ETC___d4438 =
	     (guard__h242199 == 2'b0) ?
	       _theResult___fst_exp__h250427 :
	       (iFifo$D_OUT[38] ?
		  _theResult___exp__h251146 :
		  _theResult___fst_exp__h250427) ;
  assign IF_IF_IF_IF_3074_MINUS_SEXT_iFifo_first__087_B_ETC___d4519 =
	     (guard__h242199 == 2'b0 || iFifo$D_OUT[38]) ?
	       sfdin__h250421[56:5] :
	       _theResult___sfd__h251147 ;
  assign IF_IF_IF_IF_3074_MINUS_SEXT_iFifo_first__087_B_ETC___d4521 =
	     (guard__h242199 == 2'b0) ?
	       sfdin__h250421[56:5] :
	       (iFifo$D_OUT[38] ?
		  _theResult___sfd__h251147 :
		  sfdin__h250421[56:5]) ;
  assign IF_IF_IF_IF_3074_MINUS_SEXT_iFifo_first__087_B_ETC___d5211 =
	     (guard__h203260 == 2'b0 || iFifo$D_OUT[103]) ?
	       _theResult___fst_exp__h211488 :
	       _theResult___exp__h212207 ;
  assign IF_IF_IF_IF_3074_MINUS_SEXT_iFifo_first__087_B_ETC___d5213 =
	     (guard__h203260 == 2'b0) ?
	       _theResult___fst_exp__h211488 :
	       (iFifo$D_OUT[103] ?
		  _theResult___exp__h212207 :
		  _theResult___fst_exp__h211488) ;
  assign IF_IF_IF_IF_3074_MINUS_SEXT_iFifo_first__087_B_ETC___d5294 =
	     (guard__h203260 == 2'b0 || iFifo$D_OUT[103]) ?
	       sfdin__h211482[56:5] :
	       _theResult___sfd__h212208 ;
  assign IF_IF_IF_IF_3074_MINUS_SEXT_iFifo_first__087_B_ETC___d5296 =
	     (guard__h203260 == 2'b0) ?
	       sfdin__h211482[56:5] :
	       (iFifo$D_OUT[103] ?
		  _theResult___sfd__h212208 :
		  sfdin__h211482[56:5]) ;
  assign IF_IF_IF_IF_3970_MINUS_SEXT_resWire_wget__410__ETC___d6518 =
	     (guard__h287260 == 2'b0 || resWire$wget[68]) ?
	       _theResult___fst_exp__h295488 :
	       _theResult___exp__h296004 ;
  assign IF_IF_IF_IF_3970_MINUS_SEXT_resWire_wget__410__ETC___d6520 =
	     (guard__h287260 == 2'b0) ?
	       _theResult___fst_exp__h295488 :
	       (resWire$wget[68] ?
		  _theResult___exp__h296004 :
		  _theResult___fst_exp__h295488) ;
  assign IF_IF_IF_IF_3970_MINUS_SEXT_resWire_wget__410__ETC___d6622 =
	     (guard__h287260 == 2'b0 || resWire$wget[68]) ?
	       sfdin__h295482[56:34] :
	       _theResult___sfd__h296005 ;
  assign IF_IF_IF_IF_3970_MINUS_SEXT_resWire_wget__410__ETC___d6624 =
	     (guard__h287260 == 2'b0) ?
	       sfdin__h295482[56:34] :
	       (resWire$wget[68] ?
		  _theResult___sfd__h296005 :
		  sfdin__h295482[56:34]) ;
  assign IF_IF_IF_iFifo_first__087_BITS_102_TO_95_625_E_ETC___d5173 =
	     (guard__h194011 == 2'b0 || iFifo$D_OUT[103]) ?
	       _theResult___fst_exp__h201972 :
	       _theResult___exp__h202617 ;
  assign IF_IF_IF_iFifo_first__087_BITS_102_TO_95_625_E_ETC___d5175 =
	     (guard__h194011 == 2'b0) ?
	       _theResult___fst_exp__h201972 :
	       (iFifo$D_OUT[103] ?
		  _theResult___exp__h202617 :
		  _theResult___fst_exp__h201972) ;
  assign IF_IF_IF_iFifo_first__087_BITS_102_TO_95_625_E_ETC___d5242 =
	     (guard__h212299 == 2'b0 || iFifo$D_OUT[103]) ?
	       _theResult___fst_exp__h220289 :
	       _theResult___exp__h220959 ;
  assign IF_IF_IF_iFifo_first__087_BITS_102_TO_95_625_E_ETC___d5244 =
	     (guard__h212299 == 2'b0) ?
	       _theResult___fst_exp__h220289 :
	       (iFifo$D_OUT[103] ?
		  _theResult___exp__h220959 :
		  _theResult___fst_exp__h220289) ;
  assign IF_IF_IF_iFifo_first__087_BITS_102_TO_95_625_E_ETC___d5268 =
	     (guard__h194011 == 2'b0 || iFifo$D_OUT[103]) ?
	       _theResult___snd__h201923[56:5] :
	       _theResult___sfd__h202618 ;
  assign IF_IF_IF_iFifo_first__087_BITS_102_TO_95_625_E_ETC___d5270 =
	     (guard__h194011 == 2'b0) ?
	       _theResult___snd__h201923[56:5] :
	       (iFifo$D_OUT[103] ?
		  _theResult___sfd__h202618 :
		  _theResult___snd__h201923[56:5]) ;
  assign IF_IF_IF_iFifo_first__087_BITS_102_TO_95_625_E_ETC___d5313 =
	     (guard__h212299 == 2'b0 || iFifo$D_OUT[103]) ?
	       _theResult___snd__h220235[56:5] :
	       _theResult___sfd__h220960 ;
  assign IF_IF_IF_iFifo_first__087_BITS_102_TO_95_625_E_ETC___d5315 =
	     (guard__h212299 == 2'b0) ?
	       _theResult___snd__h220235[56:5] :
	       (iFifo$D_OUT[103] ?
		  _theResult___sfd__h220960 :
		  _theResult___snd__h220235[56:5]) ;
  assign IF_IF_IF_iFifo_first__087_BITS_167_TO_160_130__ETC___d3690 =
	     (guard__h155373 == 2'b0 || iFifo$D_OUT[168]) ?
	       _theResult___fst_exp__h163334 :
	       _theResult___exp__h163979 ;
  assign IF_IF_IF_iFifo_first__087_BITS_167_TO_160_130__ETC___d3692 =
	     (guard__h155373 == 2'b0) ?
	       _theResult___fst_exp__h163334 :
	       (iFifo$D_OUT[168] ?
		  _theResult___exp__h163979 :
		  _theResult___fst_exp__h163334) ;
  assign IF_IF_IF_iFifo_first__087_BITS_167_TO_160_130__ETC___d3760 =
	     (guard__h173661 == 2'b0 || iFifo$D_OUT[168]) ?
	       _theResult___fst_exp__h181651 :
	       _theResult___exp__h182321 ;
  assign IF_IF_IF_iFifo_first__087_BITS_167_TO_160_130__ETC___d3762 =
	     (guard__h173661 == 2'b0) ?
	       _theResult___fst_exp__h181651 :
	       (iFifo$D_OUT[168] ?
		  _theResult___exp__h182321 :
		  _theResult___fst_exp__h181651) ;
  assign IF_IF_IF_iFifo_first__087_BITS_167_TO_160_130__ETC___d3786 =
	     (guard__h155373 == 2'b0 || iFifo$D_OUT[168]) ?
	       _theResult___snd__h163285[56:5] :
	       _theResult___sfd__h163980 ;
  assign IF_IF_IF_iFifo_first__087_BITS_167_TO_160_130__ETC___d3788 =
	     (guard__h155373 == 2'b0) ?
	       _theResult___snd__h163285[56:5] :
	       (iFifo$D_OUT[168] ?
		  _theResult___sfd__h163980 :
		  _theResult___snd__h163285[56:5]) ;
  assign IF_IF_IF_iFifo_first__087_BITS_167_TO_160_130__ETC___d3832 =
	     (guard__h173661 == 2'b0 || iFifo$D_OUT[168]) ?
	       _theResult___snd__h181597[56:5] :
	       _theResult___sfd__h182322 ;
  assign IF_IF_IF_iFifo_first__087_BITS_167_TO_160_130__ETC___d3834 =
	     (guard__h173661 == 2'b0) ?
	       _theResult___snd__h181597[56:5] :
	       (iFifo$D_OUT[168] ?
		  _theResult___sfd__h182322 :
		  _theResult___snd__h181597[56:5]) ;
  assign IF_IF_IF_iFifo_first__087_BITS_37_TO_30_850_EQ_ETC___d4398 =
	     (guard__h232950 == 2'b0 || iFifo$D_OUT[38]) ?
	       _theResult___fst_exp__h240911 :
	       _theResult___exp__h241556 ;
  assign IF_IF_IF_iFifo_first__087_BITS_37_TO_30_850_EQ_ETC___d4400 =
	     (guard__h232950 == 2'b0) ?
	       _theResult___fst_exp__h240911 :
	       (iFifo$D_OUT[38] ?
		  _theResult___exp__h241556 :
		  _theResult___fst_exp__h240911) ;
  assign IF_IF_IF_iFifo_first__087_BITS_37_TO_30_850_EQ_ETC___d4467 =
	     (guard__h251238 == 2'b0 || iFifo$D_OUT[38]) ?
	       _theResult___fst_exp__h259228 :
	       _theResult___exp__h259898 ;
  assign IF_IF_IF_iFifo_first__087_BITS_37_TO_30_850_EQ_ETC___d4469 =
	     (guard__h251238 == 2'b0) ?
	       _theResult___fst_exp__h259228 :
	       (iFifo$D_OUT[38] ?
		  _theResult___exp__h259898 :
		  _theResult___fst_exp__h259228) ;
  assign IF_IF_IF_iFifo_first__087_BITS_37_TO_30_850_EQ_ETC___d4493 =
	     (guard__h232950 == 2'b0 || iFifo$D_OUT[38]) ?
	       _theResult___snd__h240862[56:5] :
	       _theResult___sfd__h241557 ;
  assign IF_IF_IF_iFifo_first__087_BITS_37_TO_30_850_EQ_ETC___d4495 =
	     (guard__h232950 == 2'b0) ?
	       _theResult___snd__h240862[56:5] :
	       (iFifo$D_OUT[38] ?
		  _theResult___sfd__h241557 :
		  _theResult___snd__h240862[56:5]) ;
  assign IF_IF_IF_iFifo_first__087_BITS_37_TO_30_850_EQ_ETC___d4538 =
	     (guard__h251238 == 2'b0 || iFifo$D_OUT[38]) ?
	       _theResult___snd__h259174[56:5] :
	       _theResult___sfd__h259899 ;
  assign IF_IF_IF_iFifo_first__087_BITS_37_TO_30_850_EQ_ETC___d4540 =
	     (guard__h251238 == 2'b0) ?
	       _theResult___snd__h259174[56:5] :
	       (iFifo$D_OUT[38] ?
		  _theResult___sfd__h259899 :
		  _theResult___snd__h259174[56:5]) ;
  assign IF_IF_IF_resWire_wget__410_BITS_67_TO_57_416_E_ETC___d6479 =
	     (guard__h278330 == 2'b0 || resWire$wget[68]) ?
	       _theResult___fst_exp__h286378 :
	       _theResult___exp__h286820 ;
  assign IF_IF_IF_resWire_wget__410_BITS_67_TO_57_416_E_ETC___d6481 =
	     (guard__h278330 == 2'b0) ?
	       _theResult___fst_exp__h286378 :
	       (resWire$wget[68] ?
		  _theResult___exp__h286820 :
		  _theResult___fst_exp__h286378) ;
  assign IF_IF_IF_resWire_wget__410_BITS_67_TO_57_416_E_ETC___d6549 =
	     (guard__h296096 == 2'b0 || resWire$wget[68]) ?
	       _theResult___fst_exp__h304173 :
	       _theResult___exp__h304640 ;
  assign IF_IF_IF_resWire_wget__410_BITS_67_TO_57_416_E_ETC___d6551 =
	     (guard__h296096 == 2'b0) ?
	       _theResult___fst_exp__h304173 :
	       (resWire$wget[68] ?
		  _theResult___exp__h304640 :
		  _theResult___fst_exp__h304173) ;
  assign IF_IF_IF_resWire_wget__410_BITS_67_TO_57_416_E_ETC___d6595 =
	     (guard__h278330 == 2'b0 || resWire$wget[68]) ?
	       _theResult___snd__h286329[56:34] :
	       _theResult___sfd__h286821 ;
  assign IF_IF_IF_resWire_wget__410_BITS_67_TO_57_416_E_ETC___d6597 =
	     (guard__h278330 == 2'b0) ?
	       _theResult___snd__h286329[56:34] :
	       (resWire$wget[68] ?
		  _theResult___sfd__h286821 :
		  _theResult___snd__h286329[56:34]) ;
  assign IF_IF_IF_resWire_wget__410_BITS_67_TO_57_416_E_ETC___d6641 =
	     (guard__h296096 == 2'b0 || resWire$wget[68]) ?
	       _theResult___snd__h304119[56:34] :
	       _theResult___sfd__h304641 ;
  assign IF_IF_IF_resWire_wget__410_BITS_67_TO_57_416_E_ETC___d6643 =
	     (guard__h296096 == 2'b0) ?
	       _theResult___snd__h304119[56:34] :
	       (resWire$wget[68] ?
		  _theResult___sfd__h304641 :
		  _theResult___snd__h304119[56:34]) ;
  assign IF_IF_fpu_div_fState_S3_first__16_BITS_120_TO__ETC___d573 =
	     (_theResult___fst_exp__h41341 == 11'd0) ?
	       12'd3074 :
	       { theResult___fst_exp1341_MINUS_1023__q11[10],
		 theResult___fst_exp1341_MINUS_1023__q11 } ;
  assign IF_IF_fpu_div_fState_S3_first__16_BITS_120_TO__ETC___d810 =
	     (sfdin__h33169[57] ?
		6'd0 :
		(sfdin__h33169[56] ?
		   6'd1 :
		   (sfdin__h33169[55] ?
		      6'd2 :
		      (sfdin__h33169[54] ?
			 6'd3 :
			 (sfdin__h33169[53] ?
			    6'd4 :
			    (sfdin__h33169[52] ?
			       6'd5 :
			       (sfdin__h33169[51] ?
				  6'd6 :
				  (sfdin__h33169[50] ?
				     6'd7 :
				     (sfdin__h33169[49] ?
					6'd8 :
					(sfdin__h33169[48] ?
					   6'd9 :
					   (sfdin__h33169[47] ?
					      6'd10 :
					      (sfdin__h33169[46] ?
						 6'd11 :
						 (sfdin__h33169[45] ?
						    6'd12 :
						    (sfdin__h33169[44] ?
						       6'd13 :
						       (sfdin__h33169[43] ?
							  6'd14 :
							  (sfdin__h33169[42] ?
							     6'd15 :
							     (sfdin__h33169[41] ?
								6'd16 :
								(sfdin__h33169[40] ?
								   6'd17 :
								   (sfdin__h33169[39] ?
								      6'd18 :
								      (sfdin__h33169[38] ?
									 6'd19 :
									 (sfdin__h33169[37] ?
									    6'd20 :
									    (sfdin__h33169[36] ?
									       6'd21 :
									       (sfdin__h33169[35] ?
										  6'd22 :
										  (sfdin__h33169[34] ?
										     6'd23 :
										     (sfdin__h33169[33] ?
											6'd24 :
											(sfdin__h33169[32] ?
											   6'd25 :
											   (sfdin__h33169[31] ?
											      6'd26 :
											      (sfdin__h33169[30] ?
												 6'd27 :
												 (sfdin__h33169[29] ?
												    6'd28 :
												    (sfdin__h33169[28] ?
												       6'd29 :
												       (sfdin__h33169[27] ?
													  6'd30 :
													  (sfdin__h33169[26] ?
													     6'd31 :
													     (sfdin__h33169[25] ?
														6'd32 :
														(sfdin__h33169[24] ?
														   6'd33 :
														   (sfdin__h33169[23] ?
														      6'd34 :
														      (sfdin__h33169[22] ?
															 6'd35 :
															 (sfdin__h33169[21] ?
															    6'd36 :
															    (sfdin__h33169[20] ?
															       6'd37 :
															       (sfdin__h33169[19] ?
																  6'd38 :
																  (sfdin__h33169[18] ?
																     6'd39 :
																     (sfdin__h33169[17] ?
																	6'd40 :
																	(sfdin__h33169[16] ?
																	   6'd41 :
																	   (sfdin__h33169[15] ?
																	      6'd42 :
																	      (sfdin__h33169[14] ?
																		 6'd43 :
																		 (sfdin__h33169[13] ?
																		    6'd44 :
																		    (sfdin__h33169[12] ?
																		       6'd45 :
																		       (sfdin__h33169[11] ?
																			  6'd46 :
																			  (sfdin__h33169[10] ?
																			     6'd47 :
																			     (sfdin__h33169[9] ?
																				6'd48 :
																				(sfdin__h33169[8] ?
																				   6'd49 :
																				   (sfdin__h33169[7] ?
																				      6'd50 :
																				      (sfdin__h33169[6] ?
																					 6'd51 :
																					 (sfdin__h33169[5] ?
																					    6'd52 :
																					    (sfdin__h33169[4] ?
																					       6'd53 :
																					       (sfdin__h33169[3] ?
																						  6'd54 :
																						  (sfdin__h33169[2] ?
																						     6'd55 :
																						     (sfdin__h33169[1] ?
																							6'd56 :
																							(sfdin__h33169[0] ?
																							   6'd57 :
																							   6'd58)))))))))))))))))))))))))))))))))))))))))))))))))))))))))) -
	     6'd1 ;
  assign IF_IF_fpu_div_fState_S3_first__16_BITS_120_TO__ETC___d812 =
	     IF_IF_fpu_div_fState_S3_first__16_BITS_120_TO__ETC___d573 -
	     12'd3074 ;
  assign IF_IF_fpu_div_fState_S3_first__16_BITS_120_TO__ETC___d856 =
	     IF_fpu_div_fState_S3_first__16_BITS_120_TO_110_ETC___d527 ?
	       IF_fpu_div_fState_S3_first__16_BITS_120_TO_110_ETC___d851 :
	       { fpu_div_fState_S3$D_OUT[129:128],
		 (fpu_div_fState_S3$D_OUT[120:110] == 11'd2047) ?
		   fpu_div_fState_S3$D_OUT[57:56] != 2'b0 ||
		   fpu_div_fState_S3$D_OUT[127] :
		   fpu_div_fState_S3$D_OUT[127],
		 fpu_div_fState_S3$D_OUT[126],
		 (fpu_div_fState_S3$D_OUT[120:110] == 11'd2047) ?
		   fpu_div_fState_S3$D_OUT[57:56] != 2'b0 ||
		   fpu_div_fState_S3$D_OUT[125] :
		   fpu_div_fState_S3$D_OUT[125] } ;
  assign IF_IF_fpu_div_fState_S3_first__16_BITS_120_TO__ETC___d859 =
	     (sfdin__h33169[57] &&
	      IF_IF_fpu_div_fState_S3_first__16_BITS_120_TO__ETC___d573 ==
	      12'd1023) ?
	       63'h7FEFFFFFFFFFFFFF :
	       { _theResult___fst_exp__h41384, sfdin__h41378[57:6] } ;
  assign IF_IF_fpu_madd_fOperand_S0_first__803_BIT_195__ETC___d1922 =
	     (x__h96539 == 11'd2047 &&
	      _theResult___fst_sfd__h96608 == 52'd0) ?
	       fpu_madd_fOperand_S0$D_OUT[195] &&
	       fpu_madd_fOperand_S0$D_OUT[194] :
	       ((fpu_madd_fOperand_S0$D_OUT[129:119] == 11'd2047 &&
		 fpu_madd_fOperand_S0$D_OUT[118:67] == 52'd0 ||
		 fpu_madd_fOperand_S0$D_OUT[65:55] == 11'd2047 &&
		 fpu_madd_fOperand_S0$D_OUT[54:3] == 52'd0) ?
		  NOT_fpu_madd_fOperand_S0_first__803_BIT_130_85_ETC___d1854 :
		  fpu_madd_fOperand_S0$D_OUT[195] &&
		  fpu_madd_fOperand_S0$D_OUT[194]) ;
  assign IF_IF_fpu_madd_fOperand_S0_first__803_BIT_195__ETC___d1931 =
	     (x__h96539 == 11'd2047 &&
	      _theResult___fst_sfd__h96608 == 52'd0) ?
	       IF_fpu_madd_fOperand_S0_first__803_BIT_195_804_ETC___d1911 :
	       ((fpu_madd_fOperand_S0$D_OUT[129:119] == 11'd2047 &&
		 fpu_madd_fOperand_S0$D_OUT[118:67] == 52'd0 ||
		 fpu_madd_fOperand_S0$D_OUT[65:55] == 11'd2047 &&
		 fpu_madd_fOperand_S0$D_OUT[54:3] == 52'd0) ?
		  63'h7FF0000000000000 :
		  IF_fpu_madd_fOperand_S0_first__803_BIT_195_804_ETC___d1911) ;
  assign IF_IF_fpu_madd_fOperand_S0_first__803_BIT_195__ETC___d1936 =
	     (x__h96539 == 11'd2047 && _theResult___fst_sfd__h96608[51]) ?
	       { fpu_madd_fOperand_S0$D_OUT[195] &&
		 fpu_madd_fOperand_S0$D_OUT[194],
		 IF_fpu_madd_fOperand_S0_first__803_BIT_195_804_ETC___d1911 } :
	       ((fpu_madd_fOperand_S0$D_OUT[129:119] == 11'd2047 &&
		 fpu_madd_fOperand_S0$D_OUT[118]) ?
		  fpu_madd_fOperand_S0$D_OUT[130:67] :
		  ((fpu_madd_fOperand_S0$D_OUT[65:55] == 11'd2047 &&
		    fpu_madd_fOperand_S0$D_OUT[54]) ?
		     fpu_madd_fOperand_S0$D_OUT[66:3] :
		     { NOT_fpu_madd_fOperand_S0_first__803_BITS_129_T_ETC___d1923,
		       IF_fpu_madd_fOperand_S0_first__803_BITS_129_TO_ETC___d1932 })) ;
  assign IF_IF_fpu_madd_fOperand_S0_first__803_BIT_195__ETC___d1939 =
	     (x__h96539 == 11'd2047 &&
	      _theResult___fst_sfd__h96608 != 52'd0 &&
	      !_theResult___fst_sfd__h96608[51]) ?
	       { fpu_madd_fOperand_S0$D_OUT[195] &&
		 fpu_madd_fOperand_S0$D_OUT[194],
		 x__h96539,
		 sfd__h99402 } :
	       IF_fpu_madd_fOperand_S0_first__803_BITS_129_TO_ETC___d1938 ;
  assign IF_IF_fpu_madd_fState_S7_first__651_BIT_128_65_ETC___d2901 =
	     (sfd__h133119[56] ?
		6'd0 :
		(sfd__h133119[55] ?
		   6'd1 :
		   (sfd__h133119[54] ?
		      6'd2 :
		      (sfd__h133119[53] ?
			 6'd3 :
			 (sfd__h133119[52] ?
			    6'd4 :
			    (sfd__h133119[51] ?
			       6'd5 :
			       (sfd__h133119[50] ?
				  6'd6 :
				  (sfd__h133119[49] ?
				     6'd7 :
				     (sfd__h133119[48] ?
					6'd8 :
					(sfd__h133119[47] ?
					   6'd9 :
					   (sfd__h133119[46] ?
					      6'd10 :
					      (sfd__h133119[45] ?
						 6'd11 :
						 (sfd__h133119[44] ?
						    6'd12 :
						    (sfd__h133119[43] ?
						       6'd13 :
						       (sfd__h133119[42] ?
							  6'd14 :
							  (sfd__h133119[41] ?
							     6'd15 :
							     (sfd__h133119[40] ?
								6'd16 :
								(sfd__h133119[39] ?
								   6'd17 :
								   (sfd__h133119[38] ?
								      6'd18 :
								      (sfd__h133119[37] ?
									 6'd19 :
									 (sfd__h133119[36] ?
									    6'd20 :
									    (sfd__h133119[35] ?
									       6'd21 :
									       (sfd__h133119[34] ?
										  6'd22 :
										  (sfd__h133119[33] ?
										     6'd23 :
										     (sfd__h133119[32] ?
											6'd24 :
											(sfd__h133119[31] ?
											   6'd25 :
											   (sfd__h133119[30] ?
											      6'd26 :
											      (sfd__h133119[29] ?
												 6'd27 :
												 (sfd__h133119[28] ?
												    6'd28 :
												    (sfd__h133119[27] ?
												       6'd29 :
												       (sfd__h133119[26] ?
													  6'd30 :
													  (sfd__h133119[25] ?
													     6'd31 :
													     (sfd__h133119[24] ?
														6'd32 :
														(sfd__h133119[23] ?
														   6'd33 :
														   (sfd__h133119[22] ?
														      6'd34 :
														      (sfd__h133119[21] ?
															 6'd35 :
															 (sfd__h133119[20] ?
															    6'd36 :
															    (sfd__h133119[19] ?
															       6'd37 :
															       (sfd__h133119[18] ?
																  6'd38 :
																  (sfd__h133119[17] ?
																     6'd39 :
																     (sfd__h133119[16] ?
																	6'd40 :
																	(sfd__h133119[15] ?
																	   6'd41 :
																	   (sfd__h133119[14] ?
																	      6'd42 :
																	      (sfd__h133119[13] ?
																		 6'd43 :
																		 (sfd__h133119[12] ?
																		    6'd44 :
																		    (sfd__h133119[11] ?
																		       6'd45 :
																		       (sfd__h133119[10] ?
																			  6'd46 :
																			  (sfd__h133119[9] ?
																			     6'd47 :
																			     (sfd__h133119[8] ?
																				6'd48 :
																				(sfd__h133119[7] ?
																				   6'd49 :
																				   (sfd__h133119[6] ?
																				      6'd50 :
																				      (sfd__h133119[5] ?
																					 6'd51 :
																					 (sfd__h133119[4] ?
																					    6'd52 :
																					    (sfd__h133119[3] ?
																					       6'd53 :
																					       (sfd__h133119[2] ?
																						  6'd54 :
																						  (sfd__h133119[1] ?
																						     6'd55 :
																						     (sfd__h133119[0] ?
																							6'd56 :
																							6'd57))))))))))))))))))))))))))))))))))))))))))))))))))))))))) -
	     6'd1 ;
  assign IF_IF_fpu_madd_fState_S7_first__651_BIT_128_65_ETC___d2952 =
	     (sfd__h133119[56] &&
	      IF_fpu_madd_fState_S7_first__651_BITS_126_TO_1_ETC___d2668 ==
	      12'd1023) ?
	       63'h7FEFFFFFFFFFFFFF :
	       { _theResult___fst_exp__h141375, sfdin__h141369[56:5] } ;
  assign IF_IF_rg_index_1_87_ULE_58_91_THEN_NOT_rg_b_92_ETC___d1028 =
	     IF_rg_index_1_87_ULE_58_91_THEN_NOT_rg_b_92_EQ_ETC___d1009 ?
	       ((IF_rg_index_1_87_ULE_58_91_THEN_IF_rg_res_94_B_ETC___d1002 ==
		 116'd0) ?
		  IF_rg_index_1_87_ULE_58_91_THEN_IF_rg_res_94_B_ETC___d1022 :
		  IF_rg_index_1_87_ULE_58_91_THEN_IF_rg_res_94_B_ETC___d1026) :
	       IF_rg_index_1_87_ULE_58_91_THEN_IF_rg_res_94_B_ETC___d1026 ;
  assign IF_NOT_fpu_madd_fState_S3_first__995_BITS_12_T_ETC___d2503 =
	     (!fpu_madd_fState_S3_first__995_BITS_12_TO_0_001_ETC___d2002 ||
	      fpu_madd_fState_S3_first__995_BITS_12_TO_0_001_ETC___d2004) ?
	       fpu_madd_fState_S3$D_OUT[86] :
	       fpu_madd_fState_S3_first__995_BITS_86_TO_82_00_ETC___d2501[4] ;
  assign IF_NOT_fpu_madd_fState_S3_first__995_BITS_12_T_ETC___d2506 =
	     (!fpu_madd_fState_S3_first__995_BITS_12_TO_0_001_ETC___d2002 ||
	      fpu_madd_fState_S3_first__995_BITS_12_TO_0_001_ETC___d2004) ?
	       fpu_madd_fState_S3$D_OUT[85] :
	       fpu_madd_fState_S3_first__995_BITS_86_TO_82_00_ETC___d2501[3] ;
  assign IF_NOT_fpu_madd_fState_S4_first__547_BIT_130_5_ETC___d2595 =
	     { NOT_fpu_madd_fState_S4_first__547_BIT_130_553__ETC___d2584 ?
		 IF_fpu_madd_fState_S4_first__547_BITS_64_TO_54_ETC___d2563 :
		 IF_fpu_madd_fState_S4_first__547_BITS_128_TO_1_ETC___d2568,
	       NOT_fpu_madd_fState_S4_first__547_BIT_130_553__ETC___d2584 ?
		 IF_fpu_madd_fState_S4_first__547_BITS_64_TO_54_ETC___d2563 -
		 IF_fpu_madd_fState_S4_first__547_BITS_128_TO_1_ETC___d2568 :
		 IF_fpu_madd_fState_S4_first__547_BITS_128_TO_1_ETC___d2568 -
		 IF_fpu_madd_fState_S4_first__547_BITS_64_TO_54_ETC___d2563,
	       x__h131940,
	       x__h131944 } ;
  assign IF_SEXT_iFifo_first__087_BITS_102_TO_95_625_MI_ETC___d5106 =
	     ((SEXT_iFifo_first__087_BITS_102_TO_95_625_MINUS_ETC__q96[10:0] ==
	       11'd0) ?
		12'd3074 :
		{ SEXT_iFifo_first__087_BITS_102_TO_95_625_MINUS_ETC__q99[10],
		  SEXT_iFifo_first__087_BITS_102_TO_95_625_MINUS_ETC__q99 }) -
	     12'd3074 ;
  assign IF_SEXT_iFifo_first__087_BITS_102_TO_95_625_MI_ETC___d5146 =
	     SEXT_iFifo_first__087_BITS_102_TO_95_625_MINUS_ETC___d4808 ?
	       ((_theResult___fst_exp__h211488 == 11'd2047) ?
		  iFifo$D_OUT[103] :
		  CASE_iFifoD_OUT_BITS_6_TO_4_0_CASE_guard03260_ETC__q117) :
	       ((_theResult___fst_exp__h220289 == 11'd2047) ?
		  iFifo$D_OUT[103] :
		  CASE_iFifoD_OUT_BITS_6_TO_4_0_CASE_guard12299_ETC__q119) ;
  assign IF_SEXT_iFifo_first__087_BITS_102_TO_95_625_MI_ETC___d5374 =
	     SEXT_iFifo_first__087_BITS_102_TO_95_625_MINUS_ETC___d4808 ?
	       ((_theResult___fst_exp__h211488 == 11'd2047) ?
		  !iFifo$D_OUT[103] :
		  CASE_iFifoD_OUT_BITS_6_TO_4_0_CASE_guard03260_ETC__q123) :
	       ((_theResult___fst_exp__h220289 == 11'd2047) ?
		  !iFifo$D_OUT[103] :
		  CASE_iFifoD_OUT_BITS_6_TO_4_0_CASE_guard12299_ETC__q125) ;
  assign IF_SEXT_iFifo_first__087_BITS_167_TO_160_130_M_ETC___d3623 =
	     ((SEXT_iFifo_first__087_BITS_167_TO_160_130_MINU_ETC__q36[10:0] ==
	       11'd0) ?
		12'd3074 :
		{ SEXT_iFifo_first__087_BITS_167_TO_160_130_MINU_ETC__q39[10],
		  SEXT_iFifo_first__087_BITS_167_TO_160_130_MINU_ETC__q39 }) -
	     12'd3074 ;
  assign IF_SEXT_iFifo_first__087_BITS_167_TO_160_130_M_ETC___d3663 =
	     SEXT_iFifo_first__087_BITS_167_TO_160_130_MINU_ETC___d3325 ?
	       ((_theResult___fst_exp__h172850 == 11'd2047) ?
		  iFifo$D_OUT[168] :
		  CASE_iFifoD_OUT_BITS_6_TO_4_0_CASE_guard64622_ETC__q57) :
	       ((_theResult___fst_exp__h181651 == 11'd2047) ?
		  iFifo$D_OUT[168] :
		  CASE_iFifoD_OUT_BITS_6_TO_4_0_CASE_guard73661_ETC__q59) ;
  assign IF_SEXT_iFifo_first__087_BITS_37_TO_30_850_MIN_ETC___d4331 =
	     ((SEXT_iFifo_first__087_BITS_37_TO_30_850_MINUS__ETC__q63[10:0] ==
	       11'd0) ?
		12'd3074 :
		{ SEXT_iFifo_first__087_BITS_37_TO_30_850_MINUS__ETC__q66[10],
		  SEXT_iFifo_first__087_BITS_37_TO_30_850_MINUS__ETC__q66 }) -
	     12'd3074 ;
  assign IF_SEXT_iFifo_first__087_BITS_37_TO_30_850_MIN_ETC___d4371 =
	     SEXT_iFifo_first__087_BITS_37_TO_30_850_MINUS__ETC___d4033 ?
	       ((_theResult___fst_exp__h250427 == 11'd2047) ?
		  iFifo$D_OUT[38] :
		  CASE_iFifoD_OUT_BITS_6_TO_4_0_CASE_guard42199_ETC__q84) :
	       ((_theResult___fst_exp__h259228 == 11'd2047) ?
		  iFifo$D_OUT[38] :
		  CASE_iFifoD_OUT_BITS_6_TO_4_0_CASE_guard51238_ETC__q86) ;
  assign IF_SEXT_iFifo_first__087_BITS_37_TO_30_850_MIN_ETC___d4608 =
	     SEXT_iFifo_first__087_BITS_37_TO_30_850_MINUS__ETC___d4033 ?
	       ((_theResult___fst_exp__h250427 == 11'd2047) ?
		  !iFifo$D_OUT[38] :
		  CASE_iFifoD_OUT_BITS_6_TO_4_0_CASE_guard42199_ETC__q90) :
	       ((_theResult___fst_exp__h259228 == 11'd2047) ?
		  !iFifo$D_OUT[38] :
		  CASE_iFifoD_OUT_BITS_6_TO_4_0_CASE_guard51238_ETC__q92) ;
  assign IF_SEXT_resWire_wget__410_BITS_67_TO_57_416_MI_ETC___d6332 =
	     ((SEXT_resWire_wget__410_BITS_67_TO_57_416_MINUS_ETC__q138[7:0] ==
	       8'd0) ?
		9'd386 :
		{ SEXT_resWire_wget__410_BITS_67_TO_57_416_MINUS_ETC__q141[7],
		  SEXT_resWire_wget__410_BITS_67_TO_57_416_MINUS_ETC__q141 }) -
	     9'd386 ;
  assign IF_SEXT_resWire_wget__410_BITS_67_TO_57_416_MI_ETC___d6375 =
	     SEXT_resWire_wget__410_BITS_67_TO_57_416_MINUS_ETC___d6033 ?
	       ((_theResult___fst_exp__h295488 == 8'd255) ?
		  !resWire$wget[68] :
		  IF_rmdFifo_first__778_EQ_0_779_THEN_IF_IF_IF_I_ETC___d6324) :
	       ((_theResult___fst_exp__h304173 == 8'd255) ?
		  !resWire$wget[68] :
		  IF_rmdFifo_first__778_EQ_0_779_THEN_IF_IF_IF_r_ETC___d6373) ;
  assign IF_SEXT_resWire_wget__410_BITS_67_TO_57_416_MI_ETC___d6420 =
	     SEXT_resWire_wget__410_BITS_67_TO_57_416_MINUS_ETC___d6033 ?
	       ((_theResult___fst_exp__h295488 == 8'd255) ?
		  resWire$wget[68] :
		  IF_rmdFifo_first__778_EQ_0_779_THEN_IF_IF_IF_I_ETC___d6409) :
	       ((_theResult___fst_exp__h304173 == 8'd255) ?
		  resWire$wget[68] :
		  IF_rmdFifo_first__778_EQ_0_779_THEN_IF_IF_IF_r_ETC___d6418) ;
  assign IF_SEXT_resWire_wget__410_BITS_67_TO_57_416_MI_ETC___d6734 =
	     SEXT_resWire_wget__410_BITS_67_TO_57_416_MINUS_ETC___d6033 ?
	       _0_CONCAT_IF_IF_3970_MINUS_SEXT_resWire_wget__4_ETC___d6705[2] :
	       _theResult___fst_exp__h304721 == 8'd255 &&
	       _theResult___fst_sfd__h304722 == 23'd0 ;
  assign IF_SEXT_resWire_wget__410_BITS_67_TO_57_416_MI_ETC___d6747 =
	     SEXT_resWire_wget__410_BITS_67_TO_57_416_MINUS_ETC___d6033 ?
	       _0_CONCAT_IF_IF_3970_MINUS_SEXT_resWire_wget__4_ETC___d6705[1] :
	       _theResult___fst_exp__h304173 == 8'd0 &&
	       guard__h296096 != 2'b0 ;
  assign IF_SEXT_resWire_wget__410_BITS_67_TO_57_416_MI_ETC___d6760 =
	     SEXT_resWire_wget__410_BITS_67_TO_57_416_MINUS_ETC___d6033 ?
	       _0_CONCAT_IF_IF_3970_MINUS_SEXT_resWire_wget__4_ETC___d6705[0] :
	       _theResult___fst_exp__h304173 != 8'd255 &&
	       guard__h296096 != 2'b0 ;
  assign IF_fpu_div_fOperands_S0_first__6_BITS_129_TO_1_ETC___d282 =
	     (((fpu_div_fOperands_S0$D_OUT[129:119] == 11'd0) ?
		 13'd7170 :
		 { {2{fpu_div_fOperands_S0D_OUT_BITS_129_TO_119_MIN_ETC__q7[10]}},
		   fpu_div_fOperands_S0D_OUT_BITS_129_TO_119_MIN_ETC__q7 }) -
	      { 7'd0, b__h3090 }) -
	     (((fpu_div_fOperands_S0$D_OUT[65:55] == 11'd0) ?
		 13'd7170 :
		 { {2{fpu_div_fOperands_S0D_OUT_BITS_65_TO_55_MINUS_ETC__q8[10]}},
		   fpu_div_fOperands_S0D_OUT_BITS_65_TO_55_MINUS_ETC__q8 }) -
	      { 7'd0, b__h10508 }) ;
  assign IF_fpu_div_fOperands_S0_first__6_BITS_129_TO_1_ETC___d283 =
	     (IF_fpu_div_fOperands_S0_first__6_BITS_129_TO_1_ETC___d282 ^
	      13'h1000) <=
	     13'd5120 ;
  assign IF_fpu_div_fOperands_S0_first__6_BITS_129_TO_1_ETC___d285 =
	     (IF_fpu_div_fOperands_S0_first__6_BITS_129_TO_1_ETC___d282 ^
	      13'h1000) <
	     13'd3020 ;
  assign IF_fpu_div_fOperands_S0_first__6_BITS_129_TO_1_ETC___d429 =
	     (IF_fpu_div_fOperands_S0_first__6_BITS_129_TO_1_ETC___d282 ^
	      13'h1000) <
	     13'd3074 ;
  assign IF_fpu_div_fOperands_S0_first__6_BITS_65_TO_55_ETC___d352 =
	     (fpu_div_fOperands_S0$D_OUT[65:55] == 11'd0 &&
	      fpu_div_fOperands_S0$D_OUT[54:3] == 52'd0 ||
	      fpu_div_fOperands_S0_first__6_BITS_129_TO_119__ETC___d331) ?
	       !fpu_div_fOperands_S0_first__6_BIT_130_33_EQ_fp_ETC___d335 :
	       CASE_fpu_div_fOperands_S0D_OUT_BITS_2_TO_0_0__ETC__q9 ;
  assign IF_fpu_div_fOperands_S0_first__6_BITS_65_TO_55_ETC___d363 =
	     (fpu_div_fOperands_S0$D_OUT[65:55] == 11'd0 &&
	      fpu_div_fOperands_S0$D_OUT[54:3] == 52'd0 ||
	      fpu_div_fOperands_S0$D_OUT[129:119] == 11'd2047 &&
	      fpu_div_fOperands_S0$D_OUT[118:67] == 52'd0) ?
	       11'd2047 :
	       ((fpu_div_fOperands_S0$D_OUT[129:119] == 11'd0 &&
		 fpu_div_fOperands_S0$D_OUT[118:67] == 52'd0 ||
		 fpu_div_fOperands_S0$D_OUT[65:55] == 11'd2047 &&
		 fpu_div_fOperands_S0$D_OUT[54:3] == 52'd0 ||
		 IF_fpu_div_fOperands_S0_first__6_BITS_129_TO_1_ETC___d283) ?
		  11'd0 :
		  _theResult___fst_exp__h18518) ;
  assign IF_fpu_div_fOperands_S0_first__6_BITS_65_TO_55_ETC___d380 =
	     (fpu_div_fOperands_S0$D_OUT[65:55] == 11'd0 &&
	      fpu_div_fOperands_S0$D_OUT[54:3] == 52'd0 ||
	      fpu_div_fOperands_S0_first__6_BITS_129_TO_119__ETC___d331) ?
	       52'd0 :
	       (IF_fpu_div_fOperands_S0_first__6_BITS_129_TO_1_ETC___d283 ?
		  _theResult___fst_sfd__h19008 :
		  _theResult___fst_sfd__h18519) ;
  assign IF_fpu_div_fOperands_S0_first__6_BITS_65_TO_55_ETC___d385 =
	     (fpu_div_fOperands_S0$D_OUT[65:55] == 11'd2047 &&
	      fpu_div_fOperands_S0$D_OUT[54:3] != 52'd0 &&
	      !fpu_div_fOperands_S0$D_OUT[54]) ?
	       { fpu_div_fOperands_S0$D_OUT[66:55], sfd__h17988 } :
	       ((fpu_div_fOperands_S0$D_OUT[129:119] == 11'd2047 &&
		 fpu_div_fOperands_S0$D_OUT[118]) ?
		  fpu_div_fOperands_S0$D_OUT[130:67] :
		  ((fpu_div_fOperands_S0$D_OUT[65:55] == 11'd2047 &&
		    fpu_div_fOperands_S0$D_OUT[54]) ?
		     fpu_div_fOperands_S0$D_OUT[66:3] :
		     NOT_fpu_div_fOperands_S0_first__6_BITS_129_TO__ETC___d382)) ;
  assign IF_fpu_div_fState_S3_first__16_BITS_120_TO_110_ETC___d527 =
	     (fpu_div_fState_S3$D_OUT[120:110] == 11'd2047) ?
	       fpu_div_fState_S3$D_OUT[57:56] == 2'b0 &&
	       !fpu_div_fState_S3$D_OUT[194] :
	       !fpu_div_fState_S3$D_OUT[194] ;
  assign IF_fpu_div_fState_S3_first__16_BITS_120_TO_110_ETC___d851 =
	     ((fpu_div_fState_S3$D_OUT[120:110] == 11'd2047) ?
		{ fpu_div_fState_S3$D_OUT[129:128],
		  fpu_div_fState_S3$D_OUT[57:56] != 2'b0 ||
		  fpu_div_fState_S3$D_OUT[127],
		  fpu_div_fState_S3$D_OUT[126],
		  fpu_div_fState_S3$D_OUT[57:56] != 2'b0 ||
		  fpu_div_fState_S3$D_OUT[125] } :
		fpu_div_fState_S3$D_OUT[129:125]) |
	     { 2'd0,
	       sfdin__h33169[57] &&
	       IF_IF_fpu_div_fState_S3_first__16_BITS_120_TO__ETC___d573 ==
	       12'd1023,
	       _theResult___fst_exp__h41387 == 11'd0 && guard__h32997 != 2'd0,
	       sfdin__h33169[57] &&
	       IF_IF_fpu_div_fState_S3_first__16_BITS_120_TO__ETC___d573 ==
	       12'd1023 } ;
  assign IF_fpu_div_fState_S4_first__73_BITS_64_TO_54_7_ETC___d907 =
	     (fpu_div_fState_S4$D_OUT[64:54] == 11'd0 &&
	      sfd__h42033[53:52] == 2'b01) ?
	       11'd1 :
	       fpu_div_fState_S4$D_OUT[64:54] ;
  assign IF_fpu_madd_fOperand_S0_first__803_BITS_129_TO_ETC___d1932 =
	     (fpu_madd_fOperand_S0_first__803_BITS_129_TO_11_ETC___d1926 ||
	      IF_fpu_madd_fOperand_S0_first__803_BIT_195_804_ETC___d1927 &&
	      !fpu_madd_fOperand_S0_first__803_BIT_195_804_AN_ETC___d1855) ?
	       63'h7FF8000000000000 :
	       IF_IF_fpu_madd_fOperand_S0_first__803_BIT_195__ETC___d1931 ;
  assign IF_fpu_madd_fOperand_S0_first__803_BITS_129_TO_ETC___d1938 =
	     (fpu_madd_fOperand_S0$D_OUT[129:119] == 11'd2047 &&
	      fpu_madd_fOperand_S0$D_OUT[118:67] != 52'd0 &&
	      !fpu_madd_fOperand_S0$D_OUT[118]) ?
	       { fpu_madd_fOperand_S0$D_OUT[130:119], sfd__h99405 } :
	       ((fpu_madd_fOperand_S0$D_OUT[65:55] == 11'd2047 &&
		 fpu_madd_fOperand_S0$D_OUT[54:3] != 52'd0 &&
		 !fpu_madd_fOperand_S0$D_OUT[54]) ?
		  { fpu_madd_fOperand_S0$D_OUT[66:55], sfd__h99408 } :
		  IF_IF_fpu_madd_fOperand_S0_first__803_BIT_195__ETC___d1936) ;
  assign IF_fpu_madd_fOperand_S0_first__803_BITS_129_TO_ETC___d1959 =
	     { ((fpu_madd_fOperand_S0$D_OUT[129:119] == 11'd0) ?
		  13'd7170 :
		  { {2{fpu_madd_fOperand_S0D_OUT_BITS_129_TO_119_MIN_ETC__q128[10]}},
		    fpu_madd_fOperand_S0D_OUT_BITS_129_TO_119_MIN_ETC__q128 }) +
	       ((fpu_madd_fOperand_S0$D_OUT[65:55] == 11'd0) ?
		  13'd7170 :
		  { {2{fpu_madd_fOperand_S0D_OUT_BITS_65_TO_55_MINUS_ETC__q129[10]}},
		    fpu_madd_fOperand_S0D_OUT_BITS_65_TO_55_MINUS_ETC__q129 }),
	       x__h114243,
	       x__h114255 } ;
  assign IF_fpu_madd_fOperand_S0_first__803_BIT_195_804_ETC___d1861 =
	     x__h96539 == 11'd2047 && _theResult___fst_sfd__h96608[51] ||
	     fpu_madd_fOperand_S0$D_OUT[129:119] == 11'd2047 &&
	     fpu_madd_fOperand_S0$D_OUT[118] ||
	     fpu_madd_fOperand_S0$D_OUT[65:55] == 11'd2047 &&
	     fpu_madd_fOperand_S0$D_OUT[54] ||
	     x__h96539 == 11'd2047 && _theResult___fst_sfd__h96608 == 52'd0 ||
	     fpu_madd_fOperand_S0_first__803_BITS_129_TO_11_ETC___d1857 ;
  assign IF_fpu_madd_fOperand_S0_first__803_BIT_195_804_ETC___d1911 =
	     fpu_madd_fOperand_S0$D_OUT[195] ?
	       fpu_madd_fOperand_S0$D_OUT[193:131] :
	       63'd0 ;
  assign IF_fpu_madd_fOperand_S0_first__803_BIT_195_804_ETC___d1927 =
	     x__h96539 == 11'd2047 && _theResult___fst_sfd__h96608 == 52'd0 &&
	     (fpu_madd_fOperand_S0$D_OUT[129:119] == 11'd2047 &&
	      fpu_madd_fOperand_S0$D_OUT[118:67] == 52'd0 ||
	      fpu_madd_fOperand_S0$D_OUT[65:55] == 11'd2047 &&
	      fpu_madd_fOperand_S0$D_OUT[54:3] == 52'd0) ;
  assign IF_fpu_madd_fOperand_S0_first__803_BIT_195_804_ETC___d1947 =
	     x__h96539 == 11'd2047 && _theResult___fst_sfd__h96608 != 52'd0 &&
	     !_theResult___fst_sfd__h96608[51] ||
	     fpu_madd_fOperand_S0$D_OUT[129:119] == 11'd2047 &&
	     fpu_madd_fOperand_S0$D_OUT[118:67] != 52'd0 &&
	     !fpu_madd_fOperand_S0$D_OUT[118] ||
	     fpu_madd_fOperand_S0$D_OUT[65:55] == 11'd2047 &&
	     fpu_madd_fOperand_S0$D_OUT[54:3] != 52'd0 &&
	     !fpu_madd_fOperand_S0$D_OUT[54] ||
	     NOT_IF_fpu_madd_fOperand_S0_first__803_BIT_195_ETC___d1946 ;
  assign IF_fpu_madd_fState_S3_first__995_BITS_12_TO_0__ETC___d2516 =
	     fpu_madd_fState_S3_first__995_BITS_12_TO_0_001_ETC___d2004 ?
	       fpu_madd_fProd_S3$D_OUT != 106'd0 ||
	       fpu_madd_fState_S3$D_OUT[83] :
	       fpu_madd_fState_S3_first__995_BITS_86_TO_82_00_ETC___d2501[1] ;
  assign IF_fpu_madd_fState_S3_first__995_BITS_12_TO_0__ETC___d2521 =
	     fpu_madd_fState_S3_first__995_BITS_12_TO_0_001_ETC___d2004 ?
	       fpu_madd_fProd_S3$D_OUT != 106'd0 ||
	       fpu_madd_fState_S3$D_OUT[82] :
	       fpu_madd_fState_S3_first__995_BITS_86_TO_82_00_ETC___d2501[0] ;
  assign IF_fpu_madd_fState_S3_first__995_BITS_12_TO_0__ETC___d2536 =
	     fpu_madd_fState_S3_first__995_BITS_12_TO_0_001_ETC___d2002 ?
	       (fpu_madd_fState_S3_first__995_BITS_12_TO_0_001_ETC___d2004 ?
		  63'd0 :
		  IF_IF_7170_MINUS_fpu_madd_fState_S3_first__995_ETC___d2534) :
	       63'h7FEFFFFFFFFFFFFF ;
  assign IF_fpu_madd_fState_S3_first__995_BIT_151_996_T_ETC___d2525 =
	     fpu_madd_fState_S3$D_OUT[151] ?
	       fpu_madd_fState_S3$D_OUT[86:82] :
	       { IF_NOT_fpu_madd_fState_S3_first__995_BITS_12_T_ETC___d2503,
		 IF_NOT_fpu_madd_fState_S3_first__995_BITS_12_T_ETC___d2506,
		 NOT_fpu_madd_fState_S3_first__995_BITS_12_TO_0_ETC___d2523 } ;
  assign IF_fpu_madd_fState_S4_first__547_BITS_128_TO_1_ETC___d2568 =
	     (fpu_madd_fState_S4$D_OUT[128:118] == 11'd0) ?
	       13'd7170 :
	       { {2{fpu_madd_fState_S4D_OUT_BITS_128_TO_118_MINUS_ETC__q26[10]}},
		 fpu_madd_fState_S4D_OUT_BITS_128_TO_118_MINUS_ETC__q26 } ;
  assign IF_fpu_madd_fState_S4_first__547_BITS_64_TO_54_ETC___d2563 =
	     (fpu_madd_fState_S4$D_OUT[64:54] == 11'd0) ?
	       13'd7170 :
	       { {2{fpu_madd_fState_S4D_OUT_BITS_64_TO_54_MINUS_1023__q27[10]}},
		 fpu_madd_fState_S4D_OUT_BITS_64_TO_54_MINUS_1023__q27 } ;
  assign IF_fpu_madd_fState_S7_first__651_BITS_126_TO_1_ETC___d2668 =
	     (value__h141307[10:0] == 11'd0) ?
	       12'd3074 :
	       { value41307_BITS_10_TO_0_MINUS_1023__q28[10],
		 value41307_BITS_10_TO_0_MINUS_1023__q28 } ;
  assign IF_fpu_madd_fState_S7_first__651_BITS_126_TO_1_ETC___d2903 =
	     IF_fpu_madd_fState_S7_first__651_BITS_126_TO_1_ETC___d2668 -
	     12'd3074 ;
  assign IF_fpu_madd_fState_S8_first__960_BITS_65_TO_55_ETC___d2986 =
	     (fpu_madd_fState_S8$D_OUT[65:55] == 11'd0 &&
	      sfd__h142040[53:52] == 2'b01) ?
	       11'd1 :
	       fpu_madd_fState_S8$D_OUT[65:55] ;
  assign IF_fpu_madd_fState_S8_first__960_BITS_65_TO_55_ETC___d3011 =
	     (fpu_madd_fState_S8$D_OUT[65:55] == 11'd2047) ?
	       fpu_madd_fState_S8$D_OUT[65:55] :
	       _theResult___fst_exp__h142619 ;
  assign IF_fpu_madd_fState_S8_first__960_BIT_67_963_AN_ETC___d3060 =
	     (fpu_madd_fState_S8$D_OUT[67] &&
	      IF_fpu_madd_fState_S8_first__960_BITS_65_TO_55_ETC___d3011 ==
	      11'd0 &&
	      ((fpu_madd_fState_S8$D_OUT[65:55] == 11'd2047) ?
		 fpu_madd_fState_S8$D_OUT[54:3] :
		 _theResult___fst_sfd__h142620) ==
	      52'd0 &&
	      !fpu_madd_fState_S8_first__960_BITS_75_TO_71_03_ETC___d3043[0] &&
	      fpu_madd_fState_S8$D_OUT[0]) ?
	       fpu_madd_fState_S8$D_OUT[70:68] == 3'd3 :
	       ((fpu_madd_fState_S8$D_OUT[65:55] == 11'd2047) ?
		  fpu_madd_fState_S8$D_OUT[66] :
		  CASE_fpu_madd_fState_S8D_OUT_BITS_70_TO_68_0__ETC__q127) ;
  assign IF_fpu_madd_fState_S8_first__960_BIT_67_963_AN_ETC___d3081 =
	     { IF_fpu_madd_fState_S8_first__960_BIT_67_963_AN_ETC___d3060,
	       (fpu_madd_fState_S8$D_OUT[65:55] == 11'd2047) ?
		 fpu_madd_fState_S8$D_OUT[65:3] :
		 CASE_fpu_madd_fState_S8D_OUT_BITS_70_TO_68_0__ETC__q132,
	       fpu_madd_fState_S8_first__960_BITS_75_TO_71_03_ETC___d3043 } ;
  assign IF_fpu_sqr_fOperand_S0_first__059_BITS_65_TO_5_ETC___d1193 =
	     (fpu_sqr_fOperand_S0$D_OUT[65:55] == 11'd0) ?
	       (fpu_sqr_fOperand_S0$D_OUT[54] ?
		  6'd2 :
		  (fpu_sqr_fOperand_S0$D_OUT[53] ?
		     6'd3 :
		     (fpu_sqr_fOperand_S0$D_OUT[52] ?
			6'd4 :
			(fpu_sqr_fOperand_S0$D_OUT[51] ?
			   6'd5 :
			   (fpu_sqr_fOperand_S0$D_OUT[50] ?
			      6'd6 :
			      (fpu_sqr_fOperand_S0$D_OUT[49] ?
				 6'd7 :
				 (fpu_sqr_fOperand_S0$D_OUT[48] ?
				    6'd8 :
				    (fpu_sqr_fOperand_S0$D_OUT[47] ?
				       6'd9 :
				       (fpu_sqr_fOperand_S0$D_OUT[46] ?
					  6'd10 :
					  (fpu_sqr_fOperand_S0$D_OUT[45] ?
					     6'd11 :
					     (fpu_sqr_fOperand_S0$D_OUT[44] ?
						6'd12 :
						(fpu_sqr_fOperand_S0$D_OUT[43] ?
						   6'd13 :
						   (fpu_sqr_fOperand_S0$D_OUT[42] ?
						      6'd14 :
						      (fpu_sqr_fOperand_S0$D_OUT[41] ?
							 6'd15 :
							 (fpu_sqr_fOperand_S0$D_OUT[40] ?
							    6'd16 :
							    (fpu_sqr_fOperand_S0$D_OUT[39] ?
							       6'd17 :
							       (fpu_sqr_fOperand_S0$D_OUT[38] ?
								  6'd18 :
								  (fpu_sqr_fOperand_S0$D_OUT[37] ?
								     6'd19 :
								     (fpu_sqr_fOperand_S0$D_OUT[36] ?
									6'd20 :
									(fpu_sqr_fOperand_S0$D_OUT[35] ?
									   6'd21 :
									   (fpu_sqr_fOperand_S0$D_OUT[34] ?
									      6'd22 :
									      (fpu_sqr_fOperand_S0$D_OUT[33] ?
										 6'd23 :
										 (fpu_sqr_fOperand_S0$D_OUT[32] ?
										    6'd24 :
										    (fpu_sqr_fOperand_S0$D_OUT[31] ?
										       6'd25 :
										       (fpu_sqr_fOperand_S0$D_OUT[30] ?
											  6'd26 :
											  (fpu_sqr_fOperand_S0$D_OUT[29] ?
											     6'd27 :
											     (fpu_sqr_fOperand_S0$D_OUT[28] ?
												6'd28 :
												(fpu_sqr_fOperand_S0$D_OUT[27] ?
												   6'd29 :
												   (fpu_sqr_fOperand_S0$D_OUT[26] ?
												      6'd30 :
												      (fpu_sqr_fOperand_S0$D_OUT[25] ?
													 6'd31 :
													 (fpu_sqr_fOperand_S0$D_OUT[24] ?
													    6'd32 :
													    (fpu_sqr_fOperand_S0$D_OUT[23] ?
													       6'd33 :
													       (fpu_sqr_fOperand_S0$D_OUT[22] ?
														  6'd34 :
														  (fpu_sqr_fOperand_S0$D_OUT[21] ?
														     6'd35 :
														     (fpu_sqr_fOperand_S0$D_OUT[20] ?
															6'd36 :
															(fpu_sqr_fOperand_S0$D_OUT[19] ?
															   6'd37 :
															   (fpu_sqr_fOperand_S0$D_OUT[18] ?
															      6'd38 :
															      (fpu_sqr_fOperand_S0$D_OUT[17] ?
																 6'd39 :
																 (fpu_sqr_fOperand_S0$D_OUT[16] ?
																    6'd40 :
																    (fpu_sqr_fOperand_S0$D_OUT[15] ?
																       6'd41 :
																       (fpu_sqr_fOperand_S0$D_OUT[14] ?
																	  6'd42 :
																	  (fpu_sqr_fOperand_S0$D_OUT[13] ?
																	     6'd43 :
																	     (fpu_sqr_fOperand_S0$D_OUT[12] ?
																		6'd44 :
																		(fpu_sqr_fOperand_S0$D_OUT[11] ?
																		   6'd45 :
																		   (fpu_sqr_fOperand_S0$D_OUT[10] ?
																		      6'd46 :
																		      (fpu_sqr_fOperand_S0$D_OUT[9] ?
																			 6'd47 :
																			 (fpu_sqr_fOperand_S0$D_OUT[8] ?
																			    6'd48 :
																			    (fpu_sqr_fOperand_S0$D_OUT[7] ?
																			       6'd49 :
																			       (fpu_sqr_fOperand_S0$D_OUT[6] ?
																				  6'd50 :
																				  (fpu_sqr_fOperand_S0$D_OUT[5] ?
																				     6'd51 :
																				     (fpu_sqr_fOperand_S0$D_OUT[4] ?
																					6'd52 :
																					(fpu_sqr_fOperand_S0$D_OUT[3] ?
																					   6'd53 :
																					   6'd58)))))))))))))))))))))))))))))))))))))))))))))))))))) :
	       6'd1 ;
  assign IF_fpu_sqr_fOperand_S0_first__059_BITS_65_TO_5_ETC___d1195 =
	     ((fpu_sqr_fOperand_S0$D_OUT[65:55] == 11'd0) ?
		13'd7170 :
		{ {2{fpu_sqr_fOperand_S0D_OUT_BITS_65_TO_55_MINUS__ETC__q16[10]}},
		  fpu_sqr_fOperand_S0D_OUT_BITS_65_TO_55_MINUS__ETC__q16 }) -
	     { 7'd0,
	       IF_fpu_sqr_fOperand_S0_first__059_BITS_65_TO_5_ETC___d1193 } ;
  assign IF_fpu_sqr_fOperand_S0_first__059_BITS_65_TO_5_ETC___d1212 =
	     (fpu_sqr_fOperand_S0$D_OUT[65:55] == 11'd2047 &&
	      fpu_sqr_fOperand_S0$D_OUT[54] ||
	      fpu_sqr_fOperand_S0$D_OUT[65:55] == 11'd0 &&
	      fpu_sqr_fOperand_S0$D_OUT[54:3] == 52'd0 ||
	      fpu_sqr_fOperand_S0$D_OUT[65:55] == 11'd2047 &&
	      fpu_sqr_fOperand_S0$D_OUT[54:3] == 52'd0 &&
	      !fpu_sqr_fOperand_S0$D_OUT[66]) ?
	       { 1'd1,
		 fpu_sqr_fOperand_S0$D_OUT[66:3],
		 130'h00AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA } :
	       (fpu_sqr_fOperand_S0$D_OUT[66] ?
		  195'h5FFE00000000000020AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA :
		  { 70'h155555555555555540,
		    fpu_sqr_fOperand_S0$D_OUT[2:0],
		    fpu_sqr_fOperand_S0$D_OUT[66],
		    x__h52551[10:0],
		    fpu_sqr_fOperand_S0$D_OUT[54:3],
		    x__h60693 }) ;
  assign IF_fpu_sqr_fOperand_S0_first__059_BITS_65_TO_5_ETC__q17 =
	     IF_fpu_sqr_fOperand_S0_first__059_BITS_65_TO_5_ETC___d1195[12:1] ;
  assign IF_fpu_sqr_fState_S1_first__216_BIT_57_226_THE_ETC___d1342 =
	     (fpu_sqr_fState_S1$D_OUT[57] ?
		7'd0 :
		(fpu_sqr_fState_S1$D_OUT[56] ?
		   7'd1 :
		   (fpu_sqr_fState_S1$D_OUT[55] ?
		      7'd2 :
		      (fpu_sqr_fState_S1$D_OUT[54] ?
			 7'd3 :
			 (fpu_sqr_fState_S1$D_OUT[53] ?
			    7'd4 :
			    (fpu_sqr_fState_S1$D_OUT[52] ?
			       7'd5 :
			       (fpu_sqr_fState_S1$D_OUT[51] ?
				  7'd6 :
				  (fpu_sqr_fState_S1$D_OUT[50] ?
				     7'd7 :
				     (fpu_sqr_fState_S1$D_OUT[49] ?
					7'd8 :
					(fpu_sqr_fState_S1$D_OUT[48] ?
					   7'd9 :
					   (fpu_sqr_fState_S1$D_OUT[47] ?
					      7'd10 :
					      (fpu_sqr_fState_S1$D_OUT[46] ?
						 7'd11 :
						 (fpu_sqr_fState_S1$D_OUT[45] ?
						    7'd12 :
						    (fpu_sqr_fState_S1$D_OUT[44] ?
						       7'd13 :
						       (fpu_sqr_fState_S1$D_OUT[43] ?
							  7'd14 :
							  (fpu_sqr_fState_S1$D_OUT[42] ?
							     7'd15 :
							     (fpu_sqr_fState_S1$D_OUT[41] ?
								7'd16 :
								(fpu_sqr_fState_S1$D_OUT[40] ?
								   7'd17 :
								   (fpu_sqr_fState_S1$D_OUT[39] ?
								      7'd18 :
								      (fpu_sqr_fState_S1$D_OUT[38] ?
									 7'd19 :
									 (fpu_sqr_fState_S1$D_OUT[37] ?
									    7'd20 :
									    (fpu_sqr_fState_S1$D_OUT[36] ?
									       7'd21 :
									       (fpu_sqr_fState_S1$D_OUT[35] ?
										  7'd22 :
										  (fpu_sqr_fState_S1$D_OUT[34] ?
										     7'd23 :
										     (fpu_sqr_fState_S1$D_OUT[33] ?
											7'd24 :
											(fpu_sqr_fState_S1$D_OUT[32] ?
											   7'd25 :
											   (fpu_sqr_fState_S1$D_OUT[31] ?
											      7'd26 :
											      (fpu_sqr_fState_S1$D_OUT[30] ?
												 7'd27 :
												 (fpu_sqr_fState_S1$D_OUT[29] ?
												    7'd28 :
												    (fpu_sqr_fState_S1$D_OUT[28] ?
												       7'd29 :
												       (fpu_sqr_fState_S1$D_OUT[27] ?
													  7'd30 :
													  (fpu_sqr_fState_S1$D_OUT[26] ?
													     7'd31 :
													     (fpu_sqr_fState_S1$D_OUT[25] ?
														7'd32 :
														(fpu_sqr_fState_S1$D_OUT[24] ?
														   7'd33 :
														   (fpu_sqr_fState_S1$D_OUT[23] ?
														      7'd34 :
														      (fpu_sqr_fState_S1$D_OUT[22] ?
															 7'd35 :
															 (fpu_sqr_fState_S1$D_OUT[21] ?
															    7'd36 :
															    (fpu_sqr_fState_S1$D_OUT[20] ?
															       7'd37 :
															       (fpu_sqr_fState_S1$D_OUT[19] ?
																  7'd38 :
																  (fpu_sqr_fState_S1$D_OUT[18] ?
																     7'd39 :
																     (fpu_sqr_fState_S1$D_OUT[17] ?
																	7'd40 :
																	(fpu_sqr_fState_S1$D_OUT[16] ?
																	   7'd41 :
																	   (fpu_sqr_fState_S1$D_OUT[15] ?
																	      7'd42 :
																	      (fpu_sqr_fState_S1$D_OUT[14] ?
																		 7'd43 :
																		 (fpu_sqr_fState_S1$D_OUT[13] ?
																		    7'd44 :
																		    (fpu_sqr_fState_S1$D_OUT[12] ?
																		       7'd45 :
																		       (fpu_sqr_fState_S1$D_OUT[11] ?
																			  7'd46 :
																			  (fpu_sqr_fState_S1$D_OUT[10] ?
																			     7'd47 :
																			     (fpu_sqr_fState_S1$D_OUT[9] ?
																				7'd48 :
																				(fpu_sqr_fState_S1$D_OUT[8] ?
																				   7'd49 :
																				   (fpu_sqr_fState_S1$D_OUT[7] ?
																				      7'd50 :
																				      (fpu_sqr_fState_S1$D_OUT[6] ?
																					 7'd51 :
																					 (fpu_sqr_fState_S1$D_OUT[5] ?
																					    7'd52 :
																					    (fpu_sqr_fState_S1$D_OUT[4] ?
																					       7'd53 :
																					       (fpu_sqr_fState_S1$D_OUT[3] ?
																						  7'd54 :
																						  (fpu_sqr_fState_S1$D_OUT[2] ?
																						     7'd55 :
																						     (fpu_sqr_fState_S1$D_OUT[1] ?
																							7'd56 :
																							(fpu_sqr_fState_S1$D_OUT[0] ?
																							   7'd57 :
																							   7'd116)))))))))))))))))))))))))))))))))))))))))))))))))))))))))) -
	     7'd1 ;
  assign IF_fpu_sqr_fState_S3_first__375_BITS_121_TO_11_ETC___d1389 =
	     (fpu_sqr_fState_S3$D_OUT[121:111] == 11'd0) ?
	       12'd3074 :
	       { fpu_sqr_fState_S3D_OUT_BITS_121_TO_111_MINUS__ETC__q18[10],
		 fpu_sqr_fState_S3D_OUT_BITS_121_TO_111_MINUS__ETC__q18 } ;
  assign IF_fpu_sqr_fState_S3_first__375_BITS_121_TO_11_ETC___d1632 =
	     IF_fpu_sqr_fState_S3_first__375_BITS_121_TO_11_ETC___d1389 -
	     12'd3074 ;
  assign IF_fpu_sqr_fState_S3_first__375_BIT_195_376_TH_ETC___d1671 =
	     fpu_sqr_fState_S3$D_OUT[195] ?
	       fpu_sqr_fState_S3$D_OUT[128:126] :
	       { fpu_sqr_fState_S3$D_OUT[58] &&
		 IF_fpu_sqr_fState_S3_first__375_BITS_121_TO_11_ETC___d1389 ==
		 12'd1023,
		 _theResult___fst_exp__h94753 == 11'd0 &&
		 guard__h86435 != 2'd0,
		 fpu_sqr_fState_S3$D_OUT[58] &&
		 IF_fpu_sqr_fState_S3_first__375_BITS_121_TO_11_ETC___d1389 ==
		 12'd1023 } ;
  assign IF_fpu_sqr_fState_S3_first__375_BIT_58_384_AND_ETC___d1678 =
	     (fpu_sqr_fState_S3$D_OUT[58] &&
	      IF_fpu_sqr_fState_S3_first__375_BITS_121_TO_11_ETC___d1389 ==
	      12'd1023) ?
	       63'h7FEFFFFFFFFFFFFF :
	       { _theResult___fst_exp__h94750, sfdin__h94744[58:7] } ;
  assign IF_fpu_sqr_fState_S3_first__375_BIT_58_384_THE_ETC___d1630 =
	     (fpu_sqr_fState_S3$D_OUT[58] ?
		6'd0 :
		(fpu_sqr_fState_S3$D_OUT[57] ?
		   6'd1 :
		   (fpu_sqr_fState_S3$D_OUT[56] ?
		      6'd2 :
		      (fpu_sqr_fState_S3$D_OUT[55] ?
			 6'd3 :
			 (fpu_sqr_fState_S3$D_OUT[54] ?
			    6'd4 :
			    (fpu_sqr_fState_S3$D_OUT[53] ?
			       6'd5 :
			       (fpu_sqr_fState_S3$D_OUT[52] ?
				  6'd6 :
				  (fpu_sqr_fState_S3$D_OUT[51] ?
				     6'd7 :
				     (fpu_sqr_fState_S3$D_OUT[50] ?
					6'd8 :
					(fpu_sqr_fState_S3$D_OUT[49] ?
					   6'd9 :
					   (fpu_sqr_fState_S3$D_OUT[48] ?
					      6'd10 :
					      (fpu_sqr_fState_S3$D_OUT[47] ?
						 6'd11 :
						 (fpu_sqr_fState_S3$D_OUT[46] ?
						    6'd12 :
						    (fpu_sqr_fState_S3$D_OUT[45] ?
						       6'd13 :
						       (fpu_sqr_fState_S3$D_OUT[44] ?
							  6'd14 :
							  (fpu_sqr_fState_S3$D_OUT[43] ?
							     6'd15 :
							     (fpu_sqr_fState_S3$D_OUT[42] ?
								6'd16 :
								(fpu_sqr_fState_S3$D_OUT[41] ?
								   6'd17 :
								   (fpu_sqr_fState_S3$D_OUT[40] ?
								      6'd18 :
								      (fpu_sqr_fState_S3$D_OUT[39] ?
									 6'd19 :
									 (fpu_sqr_fState_S3$D_OUT[38] ?
									    6'd20 :
									    (fpu_sqr_fState_S3$D_OUT[37] ?
									       6'd21 :
									       (fpu_sqr_fState_S3$D_OUT[36] ?
										  6'd22 :
										  (fpu_sqr_fState_S3$D_OUT[35] ?
										     6'd23 :
										     (fpu_sqr_fState_S3$D_OUT[34] ?
											6'd24 :
											(fpu_sqr_fState_S3$D_OUT[33] ?
											   6'd25 :
											   (fpu_sqr_fState_S3$D_OUT[32] ?
											      6'd26 :
											      (fpu_sqr_fState_S3$D_OUT[31] ?
												 6'd27 :
												 (fpu_sqr_fState_S3$D_OUT[30] ?
												    6'd28 :
												    (fpu_sqr_fState_S3$D_OUT[29] ?
												       6'd29 :
												       (fpu_sqr_fState_S3$D_OUT[28] ?
													  6'd30 :
													  (fpu_sqr_fState_S3$D_OUT[27] ?
													     6'd31 :
													     (fpu_sqr_fState_S3$D_OUT[26] ?
														6'd32 :
														(fpu_sqr_fState_S3$D_OUT[25] ?
														   6'd33 :
														   (fpu_sqr_fState_S3$D_OUT[24] ?
														      6'd34 :
														      (fpu_sqr_fState_S3$D_OUT[23] ?
															 6'd35 :
															 (fpu_sqr_fState_S3$D_OUT[22] ?
															    6'd36 :
															    (fpu_sqr_fState_S3$D_OUT[21] ?
															       6'd37 :
															       (fpu_sqr_fState_S3$D_OUT[20] ?
																  6'd38 :
																  (fpu_sqr_fState_S3$D_OUT[19] ?
																     6'd39 :
																     (fpu_sqr_fState_S3$D_OUT[18] ?
																	6'd40 :
																	(fpu_sqr_fState_S3$D_OUT[17] ?
																	   6'd41 :
																	   (fpu_sqr_fState_S3$D_OUT[16] ?
																	      6'd42 :
																	      (fpu_sqr_fState_S3$D_OUT[15] ?
																		 6'd43 :
																		 (fpu_sqr_fState_S3$D_OUT[14] ?
																		    6'd44 :
																		    (fpu_sqr_fState_S3$D_OUT[13] ?
																		       6'd45 :
																		       (fpu_sqr_fState_S3$D_OUT[12] ?
																			  6'd46 :
																			  (fpu_sqr_fState_S3$D_OUT[11] ?
																			     6'd47 :
																			     (fpu_sqr_fState_S3$D_OUT[10] ?
																				6'd48 :
																				(fpu_sqr_fState_S3$D_OUT[9] ?
																				   6'd49 :
																				   (fpu_sqr_fState_S3$D_OUT[8] ?
																				      6'd50 :
																				      (fpu_sqr_fState_S3$D_OUT[7] ?
																					 6'd51 :
																					 (fpu_sqr_fState_S3$D_OUT[6] ?
																					    6'd52 :
																					    (fpu_sqr_fState_S3$D_OUT[5] ?
																					       6'd53 :
																					       (fpu_sqr_fState_S3$D_OUT[4] ?
																						  6'd54 :
																						  (fpu_sqr_fState_S3$D_OUT[3] ?
																						     6'd55 :
																						     (fpu_sqr_fState_S3$D_OUT[2] ?
																							6'd56 :
																							(fpu_sqr_fState_S3$D_OUT[1] ?
																							   6'd57 :
																							   (fpu_sqr_fState_S3$D_OUT[0] ?
																							      6'd58 :
																							      6'd59))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) -
	     6'd1 ;
  assign IF_fpu_sqr_fState_S4_first__687_BITS_64_TO_54__ETC___d1721 =
	     (fpu_sqr_fState_S4$D_OUT[64:54] == 11'd0 &&
	      sfd__h95416[53:52] == 2'b01) ?
	       11'd1 :
	       fpu_sqr_fState_S4$D_OUT[64:54] ;
  assign IF_iFifo_first__087_BITS_102_TO_95_625_EQ_0_63_ETC___d4757 =
	     ((iFifo$D_OUT[102:95] == 8'd0) ?
		(iFifo$D_OUT[94] ?
		   6'd2 :
		   (iFifo$D_OUT[93] ?
		      6'd3 :
		      (iFifo$D_OUT[92] ?
			 6'd4 :
			 (iFifo$D_OUT[91] ?
			    6'd5 :
			    (iFifo$D_OUT[90] ?
			       6'd6 :
			       (iFifo$D_OUT[89] ?
				  6'd7 :
				  (iFifo$D_OUT[88] ?
				     6'd8 :
				     (iFifo$D_OUT[87] ?
					6'd9 :
					(iFifo$D_OUT[86] ?
					   6'd10 :
					   (iFifo$D_OUT[85] ?
					      6'd11 :
					      (iFifo$D_OUT[84] ?
						 6'd12 :
						 (iFifo$D_OUT[83] ?
						    6'd13 :
						    (iFifo$D_OUT[82] ?
						       6'd14 :
						       (iFifo$D_OUT[81] ?
							  6'd15 :
							  (iFifo$D_OUT[80] ?
							     6'd16 :
							     (iFifo$D_OUT[79] ?
								6'd17 :
								(iFifo$D_OUT[78] ?
								   6'd18 :
								   (iFifo$D_OUT[77] ?
								      6'd19 :
								      (iFifo$D_OUT[76] ?
									 6'd20 :
									 (iFifo$D_OUT[75] ?
									    6'd21 :
									    (iFifo$D_OUT[74] ?
									       6'd22 :
									       (iFifo$D_OUT[73] ?
										  6'd23 :
										  (iFifo$D_OUT[72] ?
										     6'd24 :
										     6'd57))))))))))))))))))))))) :
		6'd1) -
	     6'd1 ;
  assign IF_iFifo_first__087_BITS_102_TO_95_625_EQ_0_63_ETC___d5148 =
	     (iFifo$D_OUT[102:95] == 8'd0) ?
	       (_3970_MINUS_0_CONCAT_IF_iFifo_first__087_BIT_94_ETC___d4684 ?
		  IF_3970_MINUS_0_CONCAT_IF_iFifo_first__087_BIT_ETC___d4802 :
		  IF_iFifo_first__087_BITS_6_TO_4_118_EQ_0_191_O_ETC___d4803) :
	       (SEXT_iFifo_first__087_BITS_102_TO_95_625_MINUS_ETC___d4807 ?
		  IF_SEXT_iFifo_first__087_BITS_102_TO_95_625_MI_ETC___d5146 :
		  IF_iFifo_first__087_BITS_6_TO_4_118_EQ_0_191_O_ETC___d4803) ;
  assign IF_iFifo_first__087_BITS_102_TO_95_625_EQ_0_63_ETC___d5376 =
	     (iFifo$D_OUT[102:95] == 8'd0) ?
	       (_3970_MINUS_0_CONCAT_IF_iFifo_first__087_BIT_94_ETC___d4684 ?
		  IF_3970_MINUS_0_CONCAT_IF_iFifo_first__087_BIT_ETC___d5347 :
		  IF_iFifo_first__087_BITS_6_TO_4_118_EQ_0_191_O_ETC___d5348) :
	       (SEXT_iFifo_first__087_BITS_102_TO_95_625_MINUS_ETC___d4807 ?
		  IF_SEXT_iFifo_first__087_BITS_102_TO_95_625_MI_ETC___d5374 :
		  IF_iFifo_first__087_BITS_6_TO_4_118_EQ_0_191_O_ETC___d5348) ;
  assign IF_iFifo_first__087_BITS_102_TO_95_625_EQ_255__ETC___d5327 =
	     { (iFifo$D_OUT[102:95] == 8'd255) ?
		 11'd2047 :
		 _theResult___fst_exp__h221052,
	       (iFifo$D_OUT[102:95] == 8'd255 &&
		iFifo$D_OUT[94:72] != 23'd0) ?
		 _theResult___snd_fst_sfd__h183124 :
		 _theResult___fst_sfd__h221056 } ;
  assign IF_iFifo_first__087_BITS_102_TO_95_625_EQ_255__ETC___d5328 =
	     { (iFifo$D_OUT[102:95] == 8'd255 &&
		iFifo$D_OUT[94:72] != 23'd0 ||
		(iFifo$D_OUT[102:95] == 8'd255 ||
		 iFifo$D_OUT[102:95] == 8'd0) &&
		iFifo$D_OUT[94:72] == 23'd0) ?
		 iFifo$D_OUT[103] :
		 IF_iFifo_first__087_BITS_102_TO_95_625_EQ_0_63_ETC___d5148,
	       IF_iFifo_first__087_BITS_102_TO_95_625_EQ_255__ETC___d5327 } ;
  assign IF_iFifo_first__087_BITS_102_TO_95_625_EQ_255__ETC___d5378 =
	     { (iFifo$D_OUT[102:95] == 8'd255 &&
		iFifo$D_OUT[94:72] != 23'd0 ||
		(iFifo$D_OUT[102:95] == 8'd255 ||
		 iFifo$D_OUT[102:95] == 8'd0) &&
		iFifo$D_OUT[94:72] == 23'd0) ?
		 !iFifo$D_OUT[103] :
		 IF_iFifo_first__087_BITS_102_TO_95_625_EQ_0_63_ETC___d5376,
	       IF_iFifo_first__087_BITS_102_TO_95_625_EQ_255__ETC___d5327 } ;
  assign IF_iFifo_first__087_BITS_167_TO_160_130_EQ_0_1_ETC___d3271 =
	     ((iFifo$D_OUT[167:160] == 8'd0) ?
		(iFifo$D_OUT[159] ?
		   6'd2 :
		   (iFifo$D_OUT[158] ?
		      6'd3 :
		      (iFifo$D_OUT[157] ?
			 6'd4 :
			 (iFifo$D_OUT[156] ?
			    6'd5 :
			    (iFifo$D_OUT[155] ?
			       6'd6 :
			       (iFifo$D_OUT[154] ?
				  6'd7 :
				  (iFifo$D_OUT[153] ?
				     6'd8 :
				     (iFifo$D_OUT[152] ?
					6'd9 :
					(iFifo$D_OUT[151] ?
					   6'd10 :
					   (iFifo$D_OUT[150] ?
					      6'd11 :
					      (iFifo$D_OUT[149] ?
						 6'd12 :
						 (iFifo$D_OUT[148] ?
						    6'd13 :
						    (iFifo$D_OUT[147] ?
						       6'd14 :
						       (iFifo$D_OUT[146] ?
							  6'd15 :
							  (iFifo$D_OUT[145] ?
							     6'd16 :
							     (iFifo$D_OUT[144] ?
								6'd17 :
								(iFifo$D_OUT[143] ?
								   6'd18 :
								   (iFifo$D_OUT[142] ?
								      6'd19 :
								      (iFifo$D_OUT[141] ?
									 6'd20 :
									 (iFifo$D_OUT[140] ?
									    6'd21 :
									    (iFifo$D_OUT[139] ?
									       6'd22 :
									       (iFifo$D_OUT[138] ?
										  6'd23 :
										  (iFifo$D_OUT[137] ?
										     6'd24 :
										     6'd57))))))))))))))))))))))) :
		6'd1) -
	     6'd1 ;
  assign IF_iFifo_first__087_BITS_167_TO_160_130_EQ_0_1_ETC___d3665 =
	     (iFifo$D_OUT[167:160] == 8'd0) ?
	       (_3970_MINUS_0_CONCAT_IF_iFifo_first__087_BIT_15_ETC___d3189 ?
		  IF_3970_MINUS_0_CONCAT_IF_iFifo_first__087_BIT_ETC___d3317 :
		  IF_iFifo_first__087_BITS_6_TO_4_118_EQ_0_191_O_ETC___d3320) :
	       (SEXT_iFifo_first__087_BITS_167_TO_160_130_MINU_ETC___d3324 ?
		  IF_SEXT_iFifo_first__087_BITS_167_TO_160_130_M_ETC___d3663 :
		  IF_iFifo_first__087_BITS_6_TO_4_118_EQ_0_191_O_ETC___d3320) ;
  assign IF_iFifo_first__087_BITS_167_TO_160_130_EQ_255_ETC___d3846 =
	     { (iFifo$D_OUT[167:160] == 8'd255 &&
		iFifo$D_OUT[159:137] != 23'd0 ||
		(iFifo$D_OUT[167:160] == 8'd255 ||
		 iFifo$D_OUT[167:160] == 8'd0) &&
		iFifo$D_OUT[159:137] == 23'd0) ?
		 iFifo$D_OUT[168] :
		 IF_iFifo_first__087_BITS_167_TO_160_130_EQ_0_1_ETC___d3665,
	       (iFifo$D_OUT[167:160] == 8'd255) ?
		 11'd2047 :
		 _theResult___fst_exp__h182414,
	       (iFifo$D_OUT[167:160] == 8'd255 &&
		iFifo$D_OUT[159:137] != 23'd0) ?
		 _theResult___snd_fst_sfd__h144484 :
		 _theResult___fst_sfd__h182418 } ;
  assign IF_iFifo_first__087_BITS_37_TO_30_850_EQ_0_856_ETC___d3982 =
	     ((iFifo$D_OUT[37:30] == 8'd0) ?
		(iFifo$D_OUT[29] ?
		   6'd2 :
		   (iFifo$D_OUT[28] ?
		      6'd3 :
		      (iFifo$D_OUT[27] ?
			 6'd4 :
			 (iFifo$D_OUT[26] ?
			    6'd5 :
			    (iFifo$D_OUT[25] ?
			       6'd6 :
			       (iFifo$D_OUT[24] ?
				  6'd7 :
				  (iFifo$D_OUT[23] ?
				     6'd8 :
				     (iFifo$D_OUT[22] ?
					6'd9 :
					(iFifo$D_OUT[21] ?
					   6'd10 :
					   (iFifo$D_OUT[20] ?
					      6'd11 :
					      (iFifo$D_OUT[19] ?
						 6'd12 :
						 (iFifo$D_OUT[18] ?
						    6'd13 :
						    (iFifo$D_OUT[17] ?
						       6'd14 :
						       (iFifo$D_OUT[16] ?
							  6'd15 :
							  (iFifo$D_OUT[15] ?
							     6'd16 :
							     (iFifo$D_OUT[14] ?
								6'd17 :
								(iFifo$D_OUT[13] ?
								   6'd18 :
								   (iFifo$D_OUT[12] ?
								      6'd19 :
								      (iFifo$D_OUT[11] ?
									 6'd20 :
									 (iFifo$D_OUT[10] ?
									    6'd21 :
									    (iFifo$D_OUT[9] ?
									       6'd22 :
									       (iFifo$D_OUT[8] ?
										  6'd23 :
										  (iFifo$D_OUT[7] ?
										     6'd24 :
										     6'd57))))))))))))))))))))))) :
		6'd1) -
	     6'd1 ;
  assign IF_iFifo_first__087_BITS_37_TO_30_850_EQ_0_856_ETC___d4373 =
	     (iFifo$D_OUT[37:30] == 8'd0) ?
	       (_3970_MINUS_0_CONCAT_IF_iFifo_first__087_BIT_29_ETC___d3909 ?
		  IF_3970_MINUS_0_CONCAT_IF_iFifo_first__087_BIT_ETC___d4027 :
		  IF_iFifo_first__087_BITS_6_TO_4_118_EQ_0_191_O_ETC___d4028) :
	       (SEXT_iFifo_first__087_BITS_37_TO_30_850_MINUS__ETC___d4032 ?
		  IF_SEXT_iFifo_first__087_BITS_37_TO_30_850_MIN_ETC___d4371 :
		  IF_iFifo_first__087_BITS_6_TO_4_118_EQ_0_191_O_ETC___d4028) ;
  assign IF_iFifo_first__087_BITS_37_TO_30_850_EQ_0_856_ETC___d4610 =
	     (iFifo$D_OUT[37:30] == 8'd0) ?
	       (_3970_MINUS_0_CONCAT_IF_iFifo_first__087_BIT_29_ETC___d3909 ?
		  IF_3970_MINUS_0_CONCAT_IF_iFifo_first__087_BIT_ETC___d4581 :
		  IF_iFifo_first__087_BITS_6_TO_4_118_EQ_0_191_O_ETC___d4582) :
	       (SEXT_iFifo_first__087_BITS_37_TO_30_850_MINUS__ETC___d4032 ?
		  IF_SEXT_iFifo_first__087_BITS_37_TO_30_850_MIN_ETC___d4608 :
		  IF_iFifo_first__087_BITS_6_TO_4_118_EQ_0_191_O_ETC___d4582) ;
  assign IF_iFifo_first__087_BITS_37_TO_30_850_EQ_255_8_ETC___d4552 =
	     { (iFifo$D_OUT[37:30] == 8'd255) ?
		 11'd2047 :
		 _theResult___fst_exp__h259991,
	       (iFifo$D_OUT[37:30] == 8'd255 && iFifo$D_OUT[29:7] != 23'd0) ?
		 _theResult___snd_fst_sfd__h222063 :
		 _theResult___fst_sfd__h259995 } ;
  assign IF_iFifo_first__087_BITS_37_TO_30_850_EQ_255_8_ETC___d4553 =
	     { (iFifo$D_OUT[37:30] == 8'd255 && iFifo$D_OUT[29:7] != 23'd0 ||
		(iFifo$D_OUT[37:30] == 8'd255 ||
		 iFifo$D_OUT[37:30] == 8'd0) &&
		iFifo$D_OUT[29:7] == 23'd0) ?
		 iFifo$D_OUT[38] :
		 IF_iFifo_first__087_BITS_37_TO_30_850_EQ_0_856_ETC___d4373,
	       IF_iFifo_first__087_BITS_37_TO_30_850_EQ_255_8_ETC___d4552 } ;
  assign IF_iFifo_first__087_BITS_37_TO_30_850_EQ_255_8_ETC___d4612 =
	     { (iFifo$D_OUT[37:30] == 8'd255 && iFifo$D_OUT[29:7] != 23'd0 ||
		(iFifo$D_OUT[37:30] == 8'd255 ||
		 iFifo$D_OUT[37:30] == 8'd0) &&
		iFifo$D_OUT[29:7] == 23'd0) ?
		 !iFifo$D_OUT[38] :
		 IF_iFifo_first__087_BITS_37_TO_30_850_EQ_0_856_ETC___d4610,
	       IF_iFifo_first__087_BITS_37_TO_30_850_EQ_255_8_ETC___d4552 } ;
  assign IF_iFifo_first__087_BIT_136_624_THEN_IF_iFifo__ETC___d5330 =
	     iFifo$D_OUT[136] ?
	       IF_iFifo_first__087_BITS_102_TO_95_625_EQ_255__ETC___d5328 :
	       iFifo$D_OUT[135:72] ;
  assign IF_iFifo_first__087_BIT_201_115_THEN_IF_iFifo__ETC___d3848 =
	     iFifo$D_OUT[201] ?
	       IF_iFifo_first__087_BITS_167_TO_160_130_EQ_255_ETC___d3846 :
	       iFifo$D_OUT[200:137] ;
  assign IF_iFifo_first__087_BIT_71_849_THEN_IF_iFifo_f_ETC___d4555 =
	     iFifo$D_OUT[71] ?
	       IF_iFifo_first__087_BITS_37_TO_30_850_EQ_255_8_ETC___d4553 :
	       iFifo$D_OUT[70:7] ;
  assign IF_iFifo_first__087_BIT_71_849_THEN_IF_iFifo_f_ETC___d4618 =
	     iFifo$D_OUT[71] ?
	       IF_iFifo_first__087_BITS_37_TO_30_850_EQ_255_8_ETC___d4612 :
	       { iFifo$D_OUT[71] || !iFifo$D_OUT[70], iFifo$D_OUT[69:7] } ;
  assign IF_isDoubleFifo_first__407_THEN_IF_isNegateFif_ETC___d6657 =
	     isDoubleFifo$D_OUT ?
	       { isNegateFifo$D_OUT ^ resWire$wget[68], resWire$wget[67:5] } :
	       { 32'hAAAAAAAA,
		 IF_isNegateFifo_first__409_THEN_IF_resWire_wge_ETC___d6424,
		 exp__h304742,
		 sfd__h304743 } ;
  assign IF_isNegateFifo_first__409_THEN_IF_resWire_wge_ETC___d6424 =
	     isNegateFifo$D_OUT ?
	       ((resWire$wget[67:57] == 11'd2047 &&
		 resWire$wget[56:5] != 52'd0 ||
		 (resWire$wget[67:57] == 11'd2047 ||
		  resWire$wget[67:57] == 11'd0) &&
		 resWire$wget[56:5] == 52'd0) ?
		  !resWire$wget[68] :
		  IF_resWire_wget__410_BITS_67_TO_57_416_EQ_0_42_ETC___d6377) :
	       ((resWire$wget[67:57] == 11'd2047 &&
		 resWire$wget[56:5] != 52'd0 ||
		 (resWire$wget[67:57] == 11'd2047 ||
		  resWire$wget[67:57] == 11'd0) &&
		 resWire$wget[56:5] == 52'd0) ?
		  resWire$wget[68] :
		  IF_resWire_wget__410_BITS_67_TO_57_416_EQ_0_42_ETC___d6422) ;
  assign IF_resWire_wget__410_BITS_67_TO_57_416_EQ_0_42_ETC___d5982 =
	     ((resWire$wget[67:57] == 11'd0) ?
		(resWire$wget[56] ?
		   6'd2 :
		   (resWire$wget[55] ?
		      6'd3 :
		      (resWire$wget[54] ?
			 6'd4 :
			 (resWire$wget[53] ?
			    6'd5 :
			    (resWire$wget[52] ?
			       6'd6 :
			       (resWire$wget[51] ?
				  6'd7 :
				  (resWire$wget[50] ?
				     6'd8 :
				     (resWire$wget[49] ?
					6'd9 :
					(resWire$wget[48] ?
					   6'd10 :
					   (resWire$wget[47] ?
					      6'd11 :
					      (resWire$wget[46] ?
						 6'd12 :
						 (resWire$wget[45] ?
						    6'd13 :
						    (resWire$wget[44] ?
						       6'd14 :
						       (resWire$wget[43] ?
							  6'd15 :
							  (resWire$wget[42] ?
							     6'd16 :
							     (resWire$wget[41] ?
								6'd17 :
								(resWire$wget[40] ?
								   6'd18 :
								   (resWire$wget[39] ?
								      6'd19 :
								      (resWire$wget[38] ?
									 6'd20 :
									 (resWire$wget[37] ?
									    6'd21 :
									    (resWire$wget[36] ?
									       6'd22 :
									       (resWire$wget[35] ?
										  6'd23 :
										  (resWire$wget[34] ?
										     6'd24 :
										     (resWire$wget[33] ?
											6'd25 :
											(resWire$wget[32] ?
											   6'd26 :
											   (resWire$wget[31] ?
											      6'd27 :
											      (resWire$wget[30] ?
												 6'd28 :
												 (resWire$wget[29] ?
												    6'd29 :
												    (resWire$wget[28] ?
												       6'd30 :
												       (resWire$wget[27] ?
													  6'd31 :
													  (resWire$wget[26] ?
													     6'd32 :
													     (resWire$wget[25] ?
														6'd33 :
														(resWire$wget[24] ?
														   6'd34 :
														   (resWire$wget[23] ?
														      6'd35 :
														      (resWire$wget[22] ?
															 6'd36 :
															 (resWire$wget[21] ?
															    6'd37 :
															    (resWire$wget[20] ?
															       6'd38 :
															       (resWire$wget[19] ?
																  6'd39 :
																  (resWire$wget[18] ?
																     6'd40 :
																     (resWire$wget[17] ?
																	6'd41 :
																	(resWire$wget[16] ?
																	   6'd42 :
																	   (resWire$wget[15] ?
																	      6'd43 :
																	      (resWire$wget[14] ?
																		 6'd44 :
																		 (resWire$wget[13] ?
																		    6'd45 :
																		    (resWire$wget[12] ?
																		       6'd46 :
																		       (resWire$wget[11] ?
																			  6'd47 :
																			  (resWire$wget[10] ?
																			     6'd48 :
																			     (resWire$wget[9] ?
																				6'd49 :
																				(resWire$wget[8] ?
																				   6'd50 :
																				   (resWire$wget[7] ?
																				      6'd51 :
																				      (resWire$wget[6] ?
																					 6'd52 :
																					 (resWire$wget[5] ?
																					    6'd53 :
																					    6'd57)))))))))))))))))))))))))))))))))))))))))))))))))))) :
		6'd1) -
	     6'd1 ;
  assign IF_resWire_wget__410_BITS_67_TO_57_416_EQ_0_42_ETC___d6377 =
	     (resWire$wget[67:57] == 11'd0) ?
	       (_3074_MINUS_0_CONCAT_IF_resWire_wget__410_BIT_5_ETC___d5532 ?
		  IF_3074_MINUS_0_CONCAT_IF_resWire_wget__410_BI_ETC___d6025 :
		  IF_rmdFifo_first__778_EQ_0_779_OR_rmdFifo_firs_ETC___d6028) :
	       (SEXT_resWire_wget__410_BITS_67_TO_57_416_MINUS_ETC___d6032 ?
		  IF_SEXT_resWire_wget__410_BITS_67_TO_57_416_MI_ETC___d6375 :
		  IF_rmdFifo_first__778_EQ_0_779_OR_rmdFifo_firs_ETC___d6028) ;
  assign IF_resWire_wget__410_BITS_67_TO_57_416_EQ_0_42_ETC___d6422 =
	     (resWire$wget[67:57] == 11'd0) ?
	       (_3074_MINUS_0_CONCAT_IF_resWire_wget__410_BIT_5_ETC___d5532 ?
		  IF_3074_MINUS_0_CONCAT_IF_resWire_wget__410_BI_ETC___d6399 :
		  IF_rmdFifo_first__778_EQ_0_779_OR_rmdFifo_firs_ETC___d6400) :
	       (SEXT_resWire_wget__410_BITS_67_TO_57_416_MINUS_ETC___d6032 ?
		  IF_SEXT_resWire_wget__410_BITS_67_TO_57_416_MI_ETC___d6420 :
		  IF_rmdFifo_first__778_EQ_0_779_OR_rmdFifo_firs_ETC___d6400) ;
  assign IF_resWire_wget__410_BITS_67_TO_57_416_EQ_0_42_ETC___d6709 =
	     (resWire$wget[67:57] == 11'd0) ?
	       _3074_MINUS_0_CONCAT_IF_resWire_wget__410_BIT_5_ETC___d6691 :
	       SEXT_resWire_wget__410_BITS_67_TO_57_416_MINUS_ETC___d6032 &&
	       SEXT_resWire_wget__410_BITS_67_TO_57_416_MINUS_ETC___d6033 &&
	       _0_CONCAT_IF_IF_3970_MINUS_SEXT_resWire_wget__4_ETC___d6705[4] ;
  assign IF_resWire_wget__410_BITS_67_TO_57_416_EQ_0_42_ETC___d6720 =
	     (resWire$wget[67:57] == 11'd0) ?
	       _3074_MINUS_0_CONCAT_IF_resWire_wget__410_BIT_5_ETC___d6716 :
	       SEXT_resWire_wget__410_BITS_67_TO_57_416_MINUS_ETC___d6032 &&
	       SEXT_resWire_wget__410_BITS_67_TO_57_416_MINUS_ETC___d6033 &&
	       _0_CONCAT_IF_IF_3970_MINUS_SEXT_resWire_wget__4_ETC___d6705[3] ;
  assign IF_resWire_wget__410_BITS_67_TO_57_416_EQ_0_42_ETC___d6736 =
	     (resWire$wget[67:57] == 11'd0) ?
	       NOT_3074_MINUS_0_CONCAT_IF_resWire_wget__410_B_ETC___d6728 :
	       !SEXT_resWire_wget__410_BITS_67_TO_57_416_MINUS_ETC___d6032 ||
	       IF_SEXT_resWire_wget__410_BITS_67_TO_57_416_MI_ETC___d6734 ;
  assign IF_resWire_wget__410_BITS_67_TO_57_416_EQ_0_42_ETC___d6749 =
	     (resWire$wget[67:57] == 11'd0) ?
	       _3074_MINUS_0_CONCAT_IF_resWire_wget__410_BIT_5_ETC___d6743 :
	       SEXT_resWire_wget__410_BITS_67_TO_57_416_MINUS_ETC___d6032 &&
	       IF_SEXT_resWire_wget__410_BITS_67_TO_57_416_MI_ETC___d6747 ;
  assign IF_resWire_wget__410_BITS_67_TO_57_416_EQ_0_42_ETC___d6762 =
	     (resWire$wget[67:57] == 11'd0) ?
	       NOT_3074_MINUS_0_CONCAT_IF_resWire_wget__410_B_ETC___d6756 :
	       !SEXT_resWire_wget__410_BITS_67_TO_57_416_MINUS_ETC___d6032 ||
	       IF_SEXT_resWire_wget__410_BITS_67_TO_57_416_MI_ETC___d6760 ;
  assign IF_rg_index_1_87_ULE_58_91_THEN_IF_rg_res_94_B_ETC___d1002 =
	     rg_index_1_87_ULE_58___d991 ? _theResult___fst__h43537 : rg_b ;
  assign IF_rg_index_1_87_ULE_58_91_THEN_IF_rg_res_94_B_ETC___d1022 =
	     rg_index_1_87_ULE_58___d991 ?
	       _theResult___snd_snd_snd__h43542 :
	       rg_r_1 ;
  assign IF_rg_index_1_87_ULE_58_91_THEN_IF_rg_res_94_B_ETC___d1026 =
	     rg_index_1_87_ULE_58___d991 ?
	       IF_rg_res_94_BIT_116_95_THEN_rg_res_94_BITS_11_ETC___d1025 :
	       rg_res[115:0] ;
  assign IF_rg_index_1_87_ULE_58_91_THEN_IF_rg_res_94_B_ETC___d1036 =
	     rg_index_1_87_ULE_58___d991 ?
	       _theResult___snd_fst__h43539 :
	       rg_s ;
  assign IF_rg_index_1_87_ULE_58_91_THEN_IF_rg_res_94_B_ETC___d1038 =
	     IF_rg_index_1_87_ULE_58_91_THEN_IF_rg_res_94_B_ETC___d1036 <
	     sum__h43732 ;
  assign IF_rg_index_1_87_ULE_58_91_THEN_NOT_rg_b_92_EQ_ETC___d1009 =
	     rg_index_1_87_ULE_58___d991 ?
	       rg_b != 116'd0 && !rg_res[116] :
	       !rg_res[116] ;
  assign IF_rg_index_1_87_ULE_58_91_THEN_rg_b_92_EQ_0_9_ETC___d997 =
	     rg_index_1_87_ULE_58___d991 ?
	       rg_b == 116'd0 || rg_res[116] :
	       rg_res[116] ;
  assign IF_rg_index_ULE_57_THEN_IF_rg_r_0_BIT_115_1_TH_ETC___d22 =
	     rg_index_ULE_57___d7 ?
	       (rg_r[115] ?
		  { rg_r[114:0], 1'd0 } + b__h31634 :
		  { rg_r[114:0], 1'd0 } - b__h31634) :
	       rg_r ;
  assign IF_rg_index_ULE_57_THEN_rg_q_BITS_56_TO_0_CONC_ETC___d14 =
	     rg_index_ULE_57___d7 ? { rg_q[56:0], !rg_r[115] } : rg_q ;
  assign IF_rg_r_BIT_115_THEN_rg_q_PLUS_NEG_INV_rg_q_89_ETC__q10 =
	     rg_r[115] ?
	       rg_q_PLUS_NEG_INV_rg_q_89_90___d491 - 58'd1 :
	       rg_q_PLUS_NEG_INV_rg_q_89_90___d491 ;
  assign IF_rg_res_94_BIT_116_95_THEN_rg_res_94_BITS_11_ETC___d1025 =
	     rg_res[116] ?
	       rg_res[115:0] :
	       ((rg_b == 116'd0) ? rg_r_1 : rg_res[115:0]) ;
  assign IF_sfdin11482_BIT_4_THEN_2_ELSE_0__q98 =
	     sfdin__h211482[4] ? 2'd2 : 2'd0 ;
  assign IF_sfdin1378_BIT_5_THEN_2_ELSE_0__q13 =
	     sfdin__h41378[5] ? 2'd2 : 2'd0 ;
  assign IF_sfdin30943_BIT_53_THEN_2_ELSE_0__q25 =
	     sfdin__h130943[53] ? 2'd2 : 2'd0 ;
  assign IF_sfdin41369_BIT_4_THEN_2_ELSE_0__q30 =
	     sfdin__h141369[4] ? 2'd2 : 2'd0 ;
  assign IF_sfdin4744_BIT_6_THEN_2_ELSE_0__q20 =
	     sfdin__h94744[6] ? 2'd2 : 2'd0 ;
  assign IF_sfdin50421_BIT_4_THEN_2_ELSE_0__q65 =
	     sfdin__h250421[4] ? 2'd2 : 2'd0 ;
  assign IF_sfdin72844_BIT_4_THEN_2_ELSE_0__q38 =
	     sfdin__h172844[4] ? 2'd2 : 2'd0 ;
  assign IF_sfdin77716_BIT_33_THEN_2_ELSE_0__q134 =
	     sfdin__h277716[33] ? 2'd2 : 2'd0 ;
  assign IF_sfdin95482_BIT_33_THEN_2_ELSE_0__q140 =
	     sfdin__h295482[33] ? 2'd2 : 2'd0 ;
  assign IF_theResult___snd01923_BIT_4_THEN_2_ELSE_0__q94 =
	     _theResult___snd__h201923[4] ? 2'd2 : 2'd0 ;
  assign IF_theResult___snd04119_BIT_33_THEN_2_ELSE_0__q143 =
	     _theResult___snd__h304119[33] ? 2'd2 : 2'd0 ;
  assign IF_theResult___snd20235_BIT_4_THEN_2_ELSE_0__q101 =
	     _theResult___snd__h220235[4] ? 2'd2 : 2'd0 ;
  assign IF_theResult___snd40862_BIT_4_THEN_2_ELSE_0__q61 =
	     _theResult___snd__h240862[4] ? 2'd2 : 2'd0 ;
  assign IF_theResult___snd59174_BIT_4_THEN_2_ELSE_0__q68 =
	     _theResult___snd__h259174[4] ? 2'd2 : 2'd0 ;
  assign IF_theResult___snd63285_BIT_4_THEN_2_ELSE_0__q34 =
	     _theResult___snd__h163285[4] ? 2'd2 : 2'd0 ;
  assign IF_theResult___snd81597_BIT_4_THEN_2_ELSE_0__q41 =
	     _theResult___snd__h181597[4] ? 2'd2 : 2'd0 ;
  assign IF_theResult___snd86329_BIT_33_THEN_2_ELSE_0__q136 =
	     _theResult___snd__h286329[33] ? 2'd2 : 2'd0 ;
  assign NOT_3074_MINUS_0_CONCAT_IF_resWire_wget__410_B_ETC___d6728 =
	     !_3074_MINUS_0_CONCAT_IF_resWire_wget__410_BIT_5_ETC___d5532 ||
	     (_3074_MINUS_0_CONCAT_IF_resWire_wget__410_BIT_5_ETC___d5533 ?
		_0_CONCAT_IF_IF_0b0_CONCAT_NOT_resWire_wget__41_ETC___d6676[2] :
		_0_CONCAT_IF_resWire_wget__410_BITS_67_TO_57_41_ETC___d6688[2]) ;
  assign NOT_3074_MINUS_0_CONCAT_IF_resWire_wget__410_B_ETC___d6756 =
	     !_3074_MINUS_0_CONCAT_IF_resWire_wget__410_BIT_5_ETC___d5532 ||
	     (_3074_MINUS_0_CONCAT_IF_resWire_wget__410_BIT_5_ETC___d5533 ?
		_0_CONCAT_IF_IF_0b0_CONCAT_NOT_resWire_wget__41_ETC___d6676[0] :
		_0_CONCAT_IF_resWire_wget__410_BITS_67_TO_57_41_ETC___d6688[0]) ;
  assign NOT_IF_fpu_madd_fOperand_S0_first__803_BIT_195_ETC___d1946 =
	     (x__h96539 != 11'd2047 || !_theResult___fst_sfd__h96608[51]) &&
	     (fpu_madd_fOperand_S0$D_OUT[129:119] != 11'd2047 ||
	      !fpu_madd_fOperand_S0$D_OUT[118]) &&
	     (fpu_madd_fOperand_S0$D_OUT[65:55] != 11'd2047 ||
	      !fpu_madd_fOperand_S0$D_OUT[54]) &&
	     (fpu_madd_fOperand_S0_first__803_BITS_129_TO_11_ETC___d1926 ||
	      IF_fpu_madd_fOperand_S0_first__803_BIT_195_804_ETC___d1927 &&
	      !fpu_madd_fOperand_S0_first__803_BIT_195_804_AN_ETC___d1855) ;
  assign NOT_fpu_div_fOperands_S0_first__6_BITS_129_TO__ETC___d330 =
	     (fpu_div_fOperands_S0$D_OUT[129:119] != 11'd2047 ||
	      fpu_div_fOperands_S0$D_OUT[118:67] != 52'd0 ||
	      fpu_div_fOperands_S0$D_OUT[65:55] != 11'd2047 ||
	      fpu_div_fOperands_S0$D_OUT[54:3] != 52'd0) &&
	     (fpu_div_fOperands_S0$D_OUT[129:119] != 11'd0 ||
	      fpu_div_fOperands_S0$D_OUT[118:67] != 52'd0 ||
	      fpu_div_fOperands_S0$D_OUT[65:55] != 11'd0 ||
	      fpu_div_fOperands_S0$D_OUT[54:3] != 52'd0) ;
  assign NOT_fpu_div_fOperands_S0_first__6_BITS_129_TO__ETC___d382 =
	     { NOT_fpu_div_fOperands_S0_first__6_BITS_129_TO__ETC___d330 &&
	       IF_fpu_div_fOperands_S0_first__6_BITS_65_TO_55_ETC___d352,
	       IF_fpu_div_fOperands_S0_first__6_BITS_65_TO_55_ETC___d363,
	       fpu_div_fOperands_S0_first__6_BITS_129_TO_119__ETC___d366 ?
		 52'h8000000000000 :
		 IF_fpu_div_fOperands_S0_first__6_BITS_65_TO_55_ETC___d380 } ;
  assign NOT_fpu_div_fOperands_S0_first__6_BITS_65_TO_5_ETC___d411 =
	     (fpu_div_fOperands_S0$D_OUT[65:55] != 11'd0 ||
	      fpu_div_fOperands_S0$D_OUT[54:3] != 52'd0) &&
	     (fpu_div_fOperands_S0$D_OUT[129:119] != 11'd2047 ||
	      fpu_div_fOperands_S0$D_OUT[118:67] != 52'd0) &&
	     (fpu_div_fOperands_S0$D_OUT[129:119] != 11'd0 ||
	      fpu_div_fOperands_S0$D_OUT[118:67] != 52'd0) &&
	     (fpu_div_fOperands_S0$D_OUT[65:55] != 11'd2047 ||
	      fpu_div_fOperands_S0$D_OUT[54:3] != 52'd0) &&
	     IF_fpu_div_fOperands_S0_first__6_BITS_129_TO_1_ETC___d283 &&
	     IF_fpu_div_fOperands_S0_first__6_BITS_129_TO_1_ETC___d285 ;
  assign NOT_fpu_div_fOperands_S0_first__6_BITS_65_TO_5_ETC___d418 =
	     (fpu_div_fOperands_S0$D_OUT[65:55] != 11'd0 ||
	      fpu_div_fOperands_S0$D_OUT[54:3] != 52'd0) &&
	     (fpu_div_fOperands_S0$D_OUT[129:119] != 11'd2047 ||
	      fpu_div_fOperands_S0$D_OUT[118:67] != 52'd0) &&
	     (fpu_div_fOperands_S0$D_OUT[129:119] != 11'd0 ||
	      fpu_div_fOperands_S0$D_OUT[118:67] != 52'd0) &&
	     (fpu_div_fOperands_S0$D_OUT[65:55] != 11'd2047 ||
	      fpu_div_fOperands_S0$D_OUT[54:3] != 52'd0) &&
	     (!IF_fpu_div_fOperands_S0_first__6_BITS_129_TO_1_ETC___d283 ||
	      IF_fpu_div_fOperands_S0_first__6_BITS_129_TO_1_ETC___d285) ;
  assign NOT_fpu_madd_fOperand_S0_first__803_BITS_129_T_ETC___d1923 =
	     (fpu_madd_fOperand_S0$D_OUT[129:119] != 11'd2047 ||
	      fpu_madd_fOperand_S0$D_OUT[118:67] != 52'd0 ||
	      fpu_madd_fOperand_S0$D_OUT[65:55] != 11'd0 ||
	      fpu_madd_fOperand_S0$D_OUT[54:3] != 52'd0) &&
	     (fpu_madd_fOperand_S0$D_OUT[129:119] != 11'd0 ||
	      fpu_madd_fOperand_S0$D_OUT[118:67] != 52'd0 ||
	      fpu_madd_fOperand_S0$D_OUT[65:55] != 11'd2047 ||
	      fpu_madd_fOperand_S0$D_OUT[54:3] != 52'd0) &&
	     (x__h96539 != 11'd2047 ||
	      _theResult___fst_sfd__h96608 != 52'd0 ||
	      (fpu_madd_fOperand_S0$D_OUT[129:119] != 11'd2047 ||
	       fpu_madd_fOperand_S0$D_OUT[118:67] != 52'd0) &&
	      (fpu_madd_fOperand_S0$D_OUT[65:55] != 11'd2047 ||
	       fpu_madd_fOperand_S0$D_OUT[54:3] != 52'd0) ||
	      fpu_madd_fOperand_S0_first__803_BIT_195_804_AN_ETC___d1855) &&
	     IF_IF_fpu_madd_fOperand_S0_first__803_BIT_195__ETC___d1922 ;
  assign NOT_fpu_madd_fOperand_S0_first__803_BIT_130_85_ETC___d1854 =
	     fpu_madd_fOperand_S0$D_OUT[130] !=
	     fpu_madd_fOperand_S0$D_OUT[66] ;
  assign NOT_fpu_madd_fState_S3_first__995_BITS_12_TO_0_ETC___d2510 =
	     !fpu_madd_fState_S3_first__995_BITS_12_TO_0_001_ETC___d2002 ||
	     (fpu_madd_fState_S3_first__995_BITS_12_TO_0_001_ETC___d2004 ?
		fpu_madd_fState_S3$D_OUT[84] :
		fpu_madd_fState_S3_first__995_BITS_86_TO_82_00_ETC___d2501[2]) ;
  assign NOT_fpu_madd_fState_S3_first__995_BITS_12_TO_0_ETC___d2523 =
	     { NOT_fpu_madd_fState_S3_first__995_BITS_12_TO_0_ETC___d2510,
	       fpu_madd_fState_S3_first__995_BITS_12_TO_0_001_ETC___d2002 ?
		 IF_fpu_madd_fState_S3_first__995_BITS_12_TO_0__ETC___d2516 :
		 fpu_madd_fState_S3$D_OUT[83],
	       !fpu_madd_fState_S3_first__995_BITS_12_TO_0_001_ETC___d2002 ||
	       IF_fpu_madd_fState_S3_first__995_BITS_12_TO_0__ETC___d2521 } ;
  assign NOT_fpu_madd_fState_S4_first__547_BIT_130_553__ETC___d2584 =
	     !fpu_madd_fState_S4$D_OUT[130] ||
	     (IF_fpu_madd_fState_S4_first__547_BITS_64_TO_54_ETC___d2563 ^
	      13'h1000) >
	     (IF_fpu_madd_fState_S4_first__547_BITS_128_TO_1_ETC___d2568 ^
	      13'h1000) ||
	     IF_fpu_madd_fState_S4_first__547_BITS_64_TO_54_ETC___d2563 ==
	     IF_fpu_madd_fState_S4_first__547_BITS_128_TO_1_ETC___d2568 &&
	     sfdBC__h131578 > sfdA__h131577 ;
  assign NOT_iFifo_first__087_BIT_158_142_202_AND_NOT_i_ETC___d3244 =
	     !iFifo$D_OUT[158] && !iFifo$D_OUT[157] && !iFifo$D_OUT[156] &&
	     !iFifo$D_OUT[155] &&
	     !iFifo$D_OUT[154] &&
	     !iFifo$D_OUT[153] &&
	     !iFifo$D_OUT[152] &&
	     !iFifo$D_OUT[151] &&
	     !iFifo$D_OUT[150] &&
	     !iFifo$D_OUT[149] &&
	     !iFifo$D_OUT[148] &&
	     !iFifo$D_OUT[147] &&
	     !iFifo$D_OUT[146] &&
	     !iFifo$D_OUT[145] &&
	     !iFifo$D_OUT[144] &&
	     !iFifo$D_OUT[143] &&
	     !iFifo$D_OUT[142] &&
	     !iFifo$D_OUT[141] &&
	     !iFifo$D_OUT[140] &&
	     !iFifo$D_OUT[139] &&
	     !iFifo$D_OUT[138] &&
	     !iFifo$D_OUT[137] ;
  assign NOT_iFifo_first__087_BIT_28_862_913_AND_NOT_iF_ETC___d3955 =
	     !iFifo$D_OUT[28] && !iFifo$D_OUT[27] && !iFifo$D_OUT[26] &&
	     !iFifo$D_OUT[25] &&
	     !iFifo$D_OUT[24] &&
	     !iFifo$D_OUT[23] &&
	     !iFifo$D_OUT[22] &&
	     !iFifo$D_OUT[21] &&
	     !iFifo$D_OUT[20] &&
	     !iFifo$D_OUT[19] &&
	     !iFifo$D_OUT[18] &&
	     !iFifo$D_OUT[17] &&
	     !iFifo$D_OUT[16] &&
	     !iFifo$D_OUT[15] &&
	     !iFifo$D_OUT[14] &&
	     !iFifo$D_OUT[13] &&
	     !iFifo$D_OUT[12] &&
	     !iFifo$D_OUT[11] &&
	     !iFifo$D_OUT[10] &&
	     !iFifo$D_OUT[9] &&
	     !iFifo$D_OUT[8] &&
	     !iFifo$D_OUT[7] ;
  assign NOT_iFifo_first__087_BIT_93_637_688_AND_NOT_iF_ETC___d4730 =
	     !iFifo$D_OUT[93] && !iFifo$D_OUT[92] && !iFifo$D_OUT[91] &&
	     !iFifo$D_OUT[90] &&
	     !iFifo$D_OUT[89] &&
	     !iFifo$D_OUT[88] &&
	     !iFifo$D_OUT[87] &&
	     !iFifo$D_OUT[86] &&
	     !iFifo$D_OUT[85] &&
	     !iFifo$D_OUT[84] &&
	     !iFifo$D_OUT[83] &&
	     !iFifo$D_OUT[82] &&
	     !iFifo$D_OUT[81] &&
	     !iFifo$D_OUT[80] &&
	     !iFifo$D_OUT[79] &&
	     !iFifo$D_OUT[78] &&
	     !iFifo$D_OUT[77] &&
	     !iFifo$D_OUT[76] &&
	     !iFifo$D_OUT[75] &&
	     !iFifo$D_OUT[74] &&
	     !iFifo$D_OUT[73] &&
	     !iFifo$D_OUT[72] ;
  assign NOT_resWire_wget__410_BIT_56_426_825_AND_NOT_r_ETC___d5927 =
	     !resWire$wget[56] && !resWire$wget[55] && !resWire$wget[54] &&
	     !resWire$wget[53] &&
	     !resWire$wget[52] &&
	     !resWire$wget[51] &&
	     !resWire$wget[50] &&
	     !resWire$wget[49] &&
	     !resWire$wget[48] &&
	     !resWire$wget[47] &&
	     !resWire$wget[46] &&
	     !resWire$wget[45] &&
	     !resWire$wget[44] &&
	     !resWire$wget[43] &&
	     !resWire$wget[42] &&
	     !resWire$wget[41] &&
	     !resWire$wget[40] &&
	     !resWire$wget[39] &&
	     !resWire$wget[38] &&
	     !resWire$wget[37] &&
	     !resWire$wget[36] &&
	     !resWire$wget[35] &&
	     !resWire$wget[34] &&
	     !resWire$wget[33] &&
	     !resWire$wget[32] &&
	     !resWire$wget[31] &&
	     !resWire$wget[30] &&
	     !resWire$wget[29] &&
	     !resWire$wget[28] &&
	     !resWire$wget[27] &&
	     !resWire$wget[26] &&
	     !resWire$wget[25] &&
	     !resWire$wget[24] &&
	     !resWire$wget[23] &&
	     !resWire$wget[22] &&
	     !resWire$wget[21] &&
	     !resWire$wget[20] &&
	     !resWire$wget[19] &&
	     !resWire$wget[18] &&
	     !resWire$wget[17] &&
	     !resWire$wget[16] &&
	     !resWire$wget[15] &&
	     !resWire$wget[14] &&
	     !resWire$wget[13] &&
	     !resWire$wget[12] &&
	     !resWire$wget[11] &&
	     !resWire$wget[10] &&
	     !resWire$wget[9] &&
	     !resWire$wget[8] &&
	     !resWire$wget[7] &&
	     !resWire$wget[6] &&
	     !resWire$wget[5] ;
  assign SEXT_iFifo_first__087_BITS_102_TO_95_625_MINUS_ETC___d4806 =
	     { {4{iFifoD_OUT_BITS_102_TO_95_MINUS_127__q95[7]}},
	       iFifoD_OUT_BITS_102_TO_95_MINUS_127__q95 } ;
  assign SEXT_iFifo_first__087_BITS_102_TO_95_625_MINUS_ETC___d4807 =
	     (SEXT_iFifo_first__087_BITS_102_TO_95_625_MINUS_ETC___d4806 ^
	      12'h800) <=
	     12'd3071 ;
  assign SEXT_iFifo_first__087_BITS_102_TO_95_625_MINUS_ETC___d4808 =
	     (SEXT_iFifo_first__087_BITS_102_TO_95_625_MINUS_ETC___d4806 ^
	      12'h800) <
	     12'd1026 ;
  assign SEXT_iFifo_first__087_BITS_102_TO_95_625_MINUS_ETC__q96 =
	     SEXT_iFifo_first__087_BITS_102_TO_95_625_MINUS_ETC___d4806 +
	     12'd1023 ;
  assign SEXT_iFifo_first__087_BITS_102_TO_95_625_MINUS_ETC__q99 =
	     SEXT_iFifo_first__087_BITS_102_TO_95_625_MINUS_ETC__q96[10:0] -
	     11'd1023 ;
  assign SEXT_iFifo_first__087_BITS_167_TO_160_130_MINU_ETC___d3323 =
	     { {4{iFifoD_OUT_BITS_167_TO_160_MINUS_127__q35[7]}},
	       iFifoD_OUT_BITS_167_TO_160_MINUS_127__q35 } ;
  assign SEXT_iFifo_first__087_BITS_167_TO_160_130_MINU_ETC___d3324 =
	     (SEXT_iFifo_first__087_BITS_167_TO_160_130_MINU_ETC___d3323 ^
	      12'h800) <=
	     12'd3071 ;
  assign SEXT_iFifo_first__087_BITS_167_TO_160_130_MINU_ETC___d3325 =
	     (SEXT_iFifo_first__087_BITS_167_TO_160_130_MINU_ETC___d3323 ^
	      12'h800) <
	     12'd1026 ;
  assign SEXT_iFifo_first__087_BITS_167_TO_160_130_MINU_ETC__q36 =
	     SEXT_iFifo_first__087_BITS_167_TO_160_130_MINU_ETC___d3323 +
	     12'd1023 ;
  assign SEXT_iFifo_first__087_BITS_167_TO_160_130_MINU_ETC__q39 =
	     SEXT_iFifo_first__087_BITS_167_TO_160_130_MINU_ETC__q36[10:0] -
	     11'd1023 ;
  assign SEXT_iFifo_first__087_BITS_37_TO_30_850_MINUS__ETC___d4031 =
	     { {4{iFifoD_OUT_BITS_37_TO_30_MINUS_127__q62[7]}},
	       iFifoD_OUT_BITS_37_TO_30_MINUS_127__q62 } ;
  assign SEXT_iFifo_first__087_BITS_37_TO_30_850_MINUS__ETC___d4032 =
	     (SEXT_iFifo_first__087_BITS_37_TO_30_850_MINUS__ETC___d4031 ^
	      12'h800) <=
	     12'd3071 ;
  assign SEXT_iFifo_first__087_BITS_37_TO_30_850_MINUS__ETC___d4033 =
	     (SEXT_iFifo_first__087_BITS_37_TO_30_850_MINUS__ETC___d4031 ^
	      12'h800) <
	     12'd1026 ;
  assign SEXT_iFifo_first__087_BITS_37_TO_30_850_MINUS__ETC__q63 =
	     SEXT_iFifo_first__087_BITS_37_TO_30_850_MINUS__ETC___d4031 +
	     12'd1023 ;
  assign SEXT_iFifo_first__087_BITS_37_TO_30_850_MINUS__ETC__q66 =
	     SEXT_iFifo_first__087_BITS_37_TO_30_850_MINUS__ETC__q63[10:0] -
	     11'd1023 ;
  assign SEXT_resWire_wget__410_BITS_67_TO_57_416_MINUS_ETC___d6031 =
	     { resWirewget_BITS_67_TO_57_MINUS_1023__q137[10],
	       resWirewget_BITS_67_TO_57_MINUS_1023__q137 } ;
  assign SEXT_resWire_wget__410_BITS_67_TO_57_416_MINUS_ETC___d6032 =
	     (SEXT_resWire_wget__410_BITS_67_TO_57_416_MINUS_ETC___d6031 ^
	      12'h800) <=
	     12'd2175 ;
  assign SEXT_resWire_wget__410_BITS_67_TO_57_416_MINUS_ETC___d6033 =
	     (SEXT_resWire_wget__410_BITS_67_TO_57_416_MINUS_ETC___d6031 ^
	      12'h800) <
	     12'd1922 ;
  assign SEXT_resWire_wget__410_BITS_67_TO_57_416_MINUS_ETC__q138 =
	     SEXT_resWire_wget__410_BITS_67_TO_57_416_MINUS_ETC___d6031 +
	     12'd127 ;
  assign SEXT_resWire_wget__410_BITS_67_TO_57_416_MINUS_ETC__q141 =
	     SEXT_resWire_wget__410_BITS_67_TO_57_416_MINUS_ETC__q138[7:0] -
	     8'd127 ;
  assign _0_CONCAT_IF_IF_0b0_CONCAT_NOT_resWire_wget__41_ETC___d5769 =
	     ({ 3'd0,
		IF_IF_0b0_CONCAT_NOT_resWire_wget__410_BITS_67_ETC___d5767 } ^
	      9'h100) <=
	     9'd256 ;
  assign _0_CONCAT_IF_IF_0b0_CONCAT_NOT_resWire_wget__41_ETC___d6676 =
	     { 3'd0,
	       _theResult___fst_exp__h277722 == 8'd0 &&
	       (sfdin__h277716[56:34] == 23'd0 || guard__h269623 != 2'b0),
	       1'd0 } |
	     { 2'd0,
	       _theResult___fst_exp__h278319 == 8'd255 &&
	       _theResult___fst_sfd__h278320 == 23'd0,
	       1'd0,
	       _theResult___fst_exp__h277722 != 8'd255 &&
	       guard__h269623 != 2'b0 } ;
  assign _0_CONCAT_IF_IF_3074_MINUS_SEXT_iFifo_first__08_ETC___d3574 =
	     ({ 6'd0,
		IF_IF_3074_MINUS_SEXT_iFifo_first__087_BITS_16_ETC___d3572 } ^
	      12'h800) <=
	     12'd2048 ;
  assign _0_CONCAT_IF_IF_3074_MINUS_SEXT_iFifo_first__08_ETC___d4282 =
	     ({ 6'd0,
		IF_IF_3074_MINUS_SEXT_iFifo_first__087_BITS_37_ETC___d4280 } ^
	      12'h800) <=
	     12'd2048 ;
  assign _0_CONCAT_IF_IF_3074_MINUS_SEXT_iFifo_first__08_ETC___d5057 =
	     ({ 6'd0,
		IF_IF_3074_MINUS_SEXT_iFifo_first__087_BITS_10_ETC___d5055 } ^
	      12'h800) <=
	     12'd2048 ;
  assign _0_CONCAT_IF_IF_3970_MINUS_SEXT_resWire_wget__4_ETC___d6280 =
	     ({ 3'd0,
		IF_IF_3970_MINUS_SEXT_resWire_wget__410_BITS_6_ETC___d6278 } ^
	      9'h100) <=
	     9'd256 ;
  assign _0_CONCAT_IF_IF_3970_MINUS_SEXT_resWire_wget__4_ETC___d6705 =
	     { 3'd0,
	       _theResult___fst_exp__h295488 == 8'd0 &&
	       (sfdin__h295482[56:34] == 23'd0 || guard__h287260 != 2'b0),
	       1'd0 } |
	     { 2'd0,
	       _theResult___fst_exp__h296085 == 8'd255 &&
	       _theResult___fst_sfd__h296086 == 23'd0,
	       1'd0,
	       _theResult___fst_exp__h295488 != 8'd255 &&
	       guard__h287260 != 2'b0 } ;
  assign _0_CONCAT_IF_IF_7170_MINUS_fpu_madd_fState_S3_f_ETC___d2463 =
	     ({ 5'd0,
		IF_IF_7170_MINUS_fpu_madd_fState_S3_first__995_ETC___d2460 } ^
	      12'h800) <=
	     (IF_IF_7170_MINUS_fpu_madd_fState_S3_first__995_ETC___d2462 ^
	      12'h800) ;
  assign _0_CONCAT_IF_IF_fpu_div_fState_S3_first__16_BIT_ETC___d813 =
	     ({ 6'd0,
		IF_IF_fpu_div_fState_S3_first__16_BITS_120_TO__ETC___d810 } ^
	      12'h800) <=
	     (IF_IF_fpu_div_fState_S3_first__16_BITS_120_TO__ETC___d812 ^
	      12'h800) ;
  assign _0_CONCAT_IF_IF_fpu_madd_fState_S7_first__651_B_ETC___d2904 =
	     ({ 6'd0,
		IF_IF_fpu_madd_fState_S7_first__651_BIT_128_65_ETC___d2901 } ^
	      12'h800) <=
	     (IF_fpu_madd_fState_S7_first__651_BITS_126_TO_1_ETC___d2903 ^
	      12'h800) ;
  assign _0_CONCAT_IF_fpu_sqr_fState_S3_first__375_BIT_5_ETC___d1633 =
	     ({ 6'd0,
		IF_fpu_sqr_fState_S3_first__375_BIT_58_384_THE_ETC___d1630 } ^
	      12'h800) <=
	     (IF_fpu_sqr_fState_S3_first__375_BITS_121_TO_11_ETC___d1632 ^
	      12'h800) ;
  assign _0_CONCAT_IF_iFifo_first__087_BITS_102_TO_95_62_ETC___d4759 =
	     ({ 6'd0,
		IF_iFifo_first__087_BITS_102_TO_95_625_EQ_0_63_ETC___d4757 } ^
	      12'h800) <=
	     12'd2944 ;
  assign _0_CONCAT_IF_iFifo_first__087_BITS_102_TO_95_62_ETC___d5107 =
	     ({ 6'd0,
		IF_iFifo_first__087_BITS_102_TO_95_625_EQ_0_63_ETC___d4757 } ^
	      12'h800) <=
	     (IF_SEXT_iFifo_first__087_BITS_102_TO_95_625_MI_ETC___d5106 ^
	      12'h800) ;
  assign _0_CONCAT_IF_iFifo_first__087_BITS_167_TO_160_1_ETC___d3273 =
	     ({ 6'd0,
		IF_iFifo_first__087_BITS_167_TO_160_130_EQ_0_1_ETC___d3271 } ^
	      12'h800) <=
	     12'd2944 ;
  assign _0_CONCAT_IF_iFifo_first__087_BITS_167_TO_160_1_ETC___d3624 =
	     ({ 6'd0,
		IF_iFifo_first__087_BITS_167_TO_160_130_EQ_0_1_ETC___d3271 } ^
	      12'h800) <=
	     (IF_SEXT_iFifo_first__087_BITS_167_TO_160_130_M_ETC___d3623 ^
	      12'h800) ;
  assign _0_CONCAT_IF_iFifo_first__087_BITS_37_TO_30_850_ETC___d3984 =
	     ({ 6'd0,
		IF_iFifo_first__087_BITS_37_TO_30_850_EQ_0_856_ETC___d3982 } ^
	      12'h800) <=
	     12'd2944 ;
  assign _0_CONCAT_IF_iFifo_first__087_BITS_37_TO_30_850_ETC___d4332 =
	     ({ 6'd0,
		IF_iFifo_first__087_BITS_37_TO_30_850_EQ_0_856_ETC___d3982 } ^
	      12'h800) <=
	     (IF_SEXT_iFifo_first__087_BITS_37_TO_30_850_MIN_ETC___d4331 ^
	      12'h800) ;
  assign _0_CONCAT_IF_resWire_wget__410_BITS_67_TO_57_41_ETC___d5984 =
	     ({ 3'd0,
		IF_resWire_wget__410_BITS_67_TO_57_416_EQ_0_42_ETC___d5982 } ^
	      9'h100) <=
	     9'd384 ;
  assign _0_CONCAT_IF_resWire_wget__410_BITS_67_TO_57_41_ETC___d6333 =
	     ({ 3'd0,
		IF_resWire_wget__410_BITS_67_TO_57_416_EQ_0_42_ETC___d5982 } ^
	      9'h100) <=
	     (IF_SEXT_resWire_wget__410_BITS_67_TO_57_416_MI_ETC___d6332 ^
	      9'h100) ;
  assign _0_CONCAT_IF_resWire_wget__410_BITS_67_TO_57_41_ETC___d6688 =
	     { 3'd0,
	       _theResult___fst_exp__h286378 == 8'd0 &&
	       guard__h278330 != 2'b0,
	       1'd0 } |
	     { 2'd0,
	       _theResult___fst_exp__h286901 == 8'd255 &&
	       _theResult___fst_sfd__h286902 == 23'd0,
	       1'd0,
	       _theResult___fst_exp__h286378 != 8'd255 &&
	       guard__h278330 != 2'b0 } ;
  assign _0b0_CONCAT_NOT_iFifo_first__087_BITS_102_TO_95_ETC___d4813 =
	     sfd__h183174 >>
	     _3074_MINUS_SEXT_iFifo_first__087_BITS_102_TO_9_ETC___d4809 ;
  assign _0b0_CONCAT_NOT_iFifo_first__087_BITS_167_TO_16_ETC___d3330 =
	     sfd__h144534 >>
	     _3074_MINUS_SEXT_iFifo_first__087_BITS_167_TO_1_ETC___d3326 ;
  assign _0b0_CONCAT_NOT_iFifo_first__087_BITS_37_TO_30__ETC___d4038 =
	     sfd__h222113 >>
	     _3074_MINUS_SEXT_iFifo_first__087_BITS_37_TO_30_ETC___d4034 ;
  assign _0b0_CONCAT_NOT_resWire_wget__410_BITS_67_TO_57_ETC___d6038 =
	     sfd__h262011 >>
	     _3970_MINUS_SEXT_resWire_wget__410_BITS_67_TO_5_ETC___d6034 ;
  assign _3074_MINUS_0_CONCAT_IF_resWire_wget__410_BIT_5_ETC___d5531 =
	     12'd3074 -
	     { 6'd0,
	       resWire$wget[56] ?
		 6'd0 :
		 (resWire$wget[55] ?
		    6'd1 :
		    (resWire$wget[54] ?
		       6'd2 :
		       (resWire$wget[53] ?
			  6'd3 :
			  (resWire$wget[52] ?
			     6'd4 :
			     (resWire$wget[51] ?
				6'd5 :
				(resWire$wget[50] ?
				   6'd6 :
				   (resWire$wget[49] ?
				      6'd7 :
				      (resWire$wget[48] ?
					 6'd8 :
					 (resWire$wget[47] ?
					    6'd9 :
					    (resWire$wget[46] ?
					       6'd10 :
					       (resWire$wget[45] ?
						  6'd11 :
						  (resWire$wget[44] ?
						     6'd12 :
						     (resWire$wget[43] ?
							6'd13 :
							(resWire$wget[42] ?
							   6'd14 :
							   (resWire$wget[41] ?
							      6'd15 :
							      (resWire$wget[40] ?
								 6'd16 :
								 (resWire$wget[39] ?
								    6'd17 :
								    (resWire$wget[38] ?
								       6'd18 :
								       (resWire$wget[37] ?
									  6'd19 :
									  (resWire$wget[36] ?
									     6'd20 :
									     (resWire$wget[35] ?
										6'd21 :
										(resWire$wget[34] ?
										   6'd22 :
										   (resWire$wget[33] ?
										      6'd23 :
										      (resWire$wget[32] ?
											 6'd24 :
											 (resWire$wget[31] ?
											    6'd25 :
											    (resWire$wget[30] ?
											       6'd26 :
											       (resWire$wget[29] ?
												  6'd27 :
												  (resWire$wget[28] ?
												     6'd28 :
												     (resWire$wget[27] ?
													6'd29 :
													(resWire$wget[26] ?
													   6'd30 :
													   (resWire$wget[25] ?
													      6'd31 :
													      (resWire$wget[24] ?
														 6'd32 :
														 (resWire$wget[23] ?
														    6'd33 :
														    (resWire$wget[22] ?
														       6'd34 :
														       (resWire$wget[21] ?
															  6'd35 :
															  (resWire$wget[20] ?
															     6'd36 :
															     (resWire$wget[19] ?
																6'd37 :
																(resWire$wget[18] ?
																   6'd38 :
																   (resWire$wget[17] ?
																      6'd39 :
																      (resWire$wget[16] ?
																	 6'd40 :
																	 (resWire$wget[15] ?
																	    6'd41 :
																	    (resWire$wget[14] ?
																	       6'd42 :
																	       (resWire$wget[13] ?
																		  6'd43 :
																		  (resWire$wget[12] ?
																		     6'd44 :
																		     (resWire$wget[11] ?
																			6'd45 :
																			(resWire$wget[10] ?
																			   6'd46 :
																			   (resWire$wget[9] ?
																			      6'd47 :
																			      (resWire$wget[8] ?
																				 6'd48 :
																				 (resWire$wget[7] ?
																				    6'd49 :
																				    (resWire$wget[6] ?
																				       6'd50 :
																				       (resWire$wget[5] ?
																					  6'd51 :
																					  6'd52))))))))))))))))))))))))))))))))))))))))))))))))))) } ;
  assign _3074_MINUS_0_CONCAT_IF_resWire_wget__410_BIT_5_ETC___d5532 =
	     (_3074_MINUS_0_CONCAT_IF_resWire_wget__410_BIT_5_ETC___d5531 ^
	      12'h800) <=
	     12'd2175 ;
  assign _3074_MINUS_0_CONCAT_IF_resWire_wget__410_BIT_5_ETC___d5533 =
	     (_3074_MINUS_0_CONCAT_IF_resWire_wget__410_BIT_5_ETC___d5531 ^
	      12'h800) <
	     12'd1922 ;
  assign _3074_MINUS_0_CONCAT_IF_resWire_wget__410_BIT_5_ETC___d6691 =
	     _3074_MINUS_0_CONCAT_IF_resWire_wget__410_BIT_5_ETC___d5532 &&
	     (_3074_MINUS_0_CONCAT_IF_resWire_wget__410_BIT_5_ETC___d5533 ?
		_0_CONCAT_IF_IF_0b0_CONCAT_NOT_resWire_wget__41_ETC___d6676[4] :
		_0_CONCAT_IF_resWire_wget__410_BITS_67_TO_57_41_ETC___d6688[4]) ;
  assign _3074_MINUS_0_CONCAT_IF_resWire_wget__410_BIT_5_ETC___d6716 =
	     _3074_MINUS_0_CONCAT_IF_resWire_wget__410_BIT_5_ETC___d5532 &&
	     (_3074_MINUS_0_CONCAT_IF_resWire_wget__410_BIT_5_ETC___d5533 ?
		_0_CONCAT_IF_IF_0b0_CONCAT_NOT_resWire_wget__41_ETC___d6676[3] :
		_0_CONCAT_IF_resWire_wget__410_BITS_67_TO_57_41_ETC___d6688[3]) ;
  assign _3074_MINUS_0_CONCAT_IF_resWire_wget__410_BIT_5_ETC___d6743 =
	     _3074_MINUS_0_CONCAT_IF_resWire_wget__410_BIT_5_ETC___d5532 &&
	     (_3074_MINUS_0_CONCAT_IF_resWire_wget__410_BIT_5_ETC___d5533 ?
		_0_CONCAT_IF_IF_0b0_CONCAT_NOT_resWire_wget__41_ETC___d6676[1] :
		_0_CONCAT_IF_resWire_wget__410_BITS_67_TO_57_41_ETC___d6688[1]) ;
  assign _3074_MINUS_SEXT_iFifo_first__087_BITS_102_TO_9_ETC___d4809 =
	     12'd3074 -
	     SEXT_iFifo_first__087_BITS_102_TO_95_625_MINUS_ETC___d4806 ;
  assign _3074_MINUS_SEXT_iFifo_first__087_BITS_167_TO_1_ETC___d3326 =
	     12'd3074 -
	     SEXT_iFifo_first__087_BITS_167_TO_160_130_MINU_ETC___d3323 ;
  assign _3074_MINUS_SEXT_iFifo_first__087_BITS_37_TO_30_ETC___d4034 =
	     12'd3074 -
	     SEXT_iFifo_first__087_BITS_37_TO_30_850_MINUS__ETC___d4031 ;
  assign _3970_MINUS_0_CONCAT_IF_iFifo_first__087_BIT_15_ETC___d3188 =
	     12'd3970 -
	     { 7'd0,
	       iFifo$D_OUT[159] ?
		 5'd0 :
		 (iFifo$D_OUT[158] ?
		    5'd1 :
		    (iFifo$D_OUT[157] ?
		       5'd2 :
		       (iFifo$D_OUT[156] ?
			  5'd3 :
			  (iFifo$D_OUT[155] ?
			     5'd4 :
			     (iFifo$D_OUT[154] ?
				5'd5 :
				(iFifo$D_OUT[153] ?
				   5'd6 :
				   (iFifo$D_OUT[152] ?
				      5'd7 :
				      (iFifo$D_OUT[151] ?
					 5'd8 :
					 (iFifo$D_OUT[150] ?
					    5'd9 :
					    (iFifo$D_OUT[149] ?
					       5'd10 :
					       (iFifo$D_OUT[148] ?
						  5'd11 :
						  (iFifo$D_OUT[147] ?
						     5'd12 :
						     (iFifo$D_OUT[146] ?
							5'd13 :
							(iFifo$D_OUT[145] ?
							   5'd14 :
							   (iFifo$D_OUT[144] ?
							      5'd15 :
							      (iFifo$D_OUT[143] ?
								 5'd16 :
								 (iFifo$D_OUT[142] ?
								    5'd17 :
								    (iFifo$D_OUT[141] ?
								       5'd18 :
								       (iFifo$D_OUT[140] ?
									  5'd19 :
									  (iFifo$D_OUT[139] ?
									     5'd20 :
									     (iFifo$D_OUT[138] ?
										5'd21 :
										(iFifo$D_OUT[137] ?
										   5'd22 :
										   5'd23)))))))))))))))))))))) } ;
  assign _3970_MINUS_0_CONCAT_IF_iFifo_first__087_BIT_15_ETC___d3189 =
	     (_3970_MINUS_0_CONCAT_IF_iFifo_first__087_BIT_15_ETC___d3188 ^
	      12'h800) <=
	     12'd3071 ;
  assign _3970_MINUS_0_CONCAT_IF_iFifo_first__087_BIT_15_ETC___d3190 =
	     (_3970_MINUS_0_CONCAT_IF_iFifo_first__087_BIT_15_ETC___d3188 ^
	      12'h800) <
	     12'd1026 ;
  assign _3970_MINUS_0_CONCAT_IF_iFifo_first__087_BIT_29_ETC___d3908 =
	     12'd3970 -
	     { 7'd0,
	       iFifo$D_OUT[29] ?
		 5'd0 :
		 (iFifo$D_OUT[28] ?
		    5'd1 :
		    (iFifo$D_OUT[27] ?
		       5'd2 :
		       (iFifo$D_OUT[26] ?
			  5'd3 :
			  (iFifo$D_OUT[25] ?
			     5'd4 :
			     (iFifo$D_OUT[24] ?
				5'd5 :
				(iFifo$D_OUT[23] ?
				   5'd6 :
				   (iFifo$D_OUT[22] ?
				      5'd7 :
				      (iFifo$D_OUT[21] ?
					 5'd8 :
					 (iFifo$D_OUT[20] ?
					    5'd9 :
					    (iFifo$D_OUT[19] ?
					       5'd10 :
					       (iFifo$D_OUT[18] ?
						  5'd11 :
						  (iFifo$D_OUT[17] ?
						     5'd12 :
						     (iFifo$D_OUT[16] ?
							5'd13 :
							(iFifo$D_OUT[15] ?
							   5'd14 :
							   (iFifo$D_OUT[14] ?
							      5'd15 :
							      (iFifo$D_OUT[13] ?
								 5'd16 :
								 (iFifo$D_OUT[12] ?
								    5'd17 :
								    (iFifo$D_OUT[11] ?
								       5'd18 :
								       (iFifo$D_OUT[10] ?
									  5'd19 :
									  (iFifo$D_OUT[9] ?
									     5'd20 :
									     (iFifo$D_OUT[8] ?
										5'd21 :
										(iFifo$D_OUT[7] ?
										   5'd22 :
										   5'd23)))))))))))))))))))))) } ;
  assign _3970_MINUS_0_CONCAT_IF_iFifo_first__087_BIT_29_ETC___d3909 =
	     (_3970_MINUS_0_CONCAT_IF_iFifo_first__087_BIT_29_ETC___d3908 ^
	      12'h800) <=
	     12'd3071 ;
  assign _3970_MINUS_0_CONCAT_IF_iFifo_first__087_BIT_29_ETC___d3910 =
	     (_3970_MINUS_0_CONCAT_IF_iFifo_first__087_BIT_29_ETC___d3908 ^
	      12'h800) <
	     12'd1026 ;
  assign _3970_MINUS_0_CONCAT_IF_iFifo_first__087_BIT_94_ETC___d4683 =
	     12'd3970 -
	     { 7'd0,
	       iFifo$D_OUT[94] ?
		 5'd0 :
		 (iFifo$D_OUT[93] ?
		    5'd1 :
		    (iFifo$D_OUT[92] ?
		       5'd2 :
		       (iFifo$D_OUT[91] ?
			  5'd3 :
			  (iFifo$D_OUT[90] ?
			     5'd4 :
			     (iFifo$D_OUT[89] ?
				5'd5 :
				(iFifo$D_OUT[88] ?
				   5'd6 :
				   (iFifo$D_OUT[87] ?
				      5'd7 :
				      (iFifo$D_OUT[86] ?
					 5'd8 :
					 (iFifo$D_OUT[85] ?
					    5'd9 :
					    (iFifo$D_OUT[84] ?
					       5'd10 :
					       (iFifo$D_OUT[83] ?
						  5'd11 :
						  (iFifo$D_OUT[82] ?
						     5'd12 :
						     (iFifo$D_OUT[81] ?
							5'd13 :
							(iFifo$D_OUT[80] ?
							   5'd14 :
							   (iFifo$D_OUT[79] ?
							      5'd15 :
							      (iFifo$D_OUT[78] ?
								 5'd16 :
								 (iFifo$D_OUT[77] ?
								    5'd17 :
								    (iFifo$D_OUT[76] ?
								       5'd18 :
								       (iFifo$D_OUT[75] ?
									  5'd19 :
									  (iFifo$D_OUT[74] ?
									     5'd20 :
									     (iFifo$D_OUT[73] ?
										5'd21 :
										(iFifo$D_OUT[72] ?
										   5'd22 :
										   5'd23)))))))))))))))))))))) } ;
  assign _3970_MINUS_0_CONCAT_IF_iFifo_first__087_BIT_94_ETC___d4684 =
	     (_3970_MINUS_0_CONCAT_IF_iFifo_first__087_BIT_94_ETC___d4683 ^
	      12'h800) <=
	     12'd3071 ;
  assign _3970_MINUS_0_CONCAT_IF_iFifo_first__087_BIT_94_ETC___d4685 =
	     (_3970_MINUS_0_CONCAT_IF_iFifo_first__087_BIT_94_ETC___d4683 ^
	      12'h800) <
	     12'd1026 ;
  assign _3970_MINUS_SEXT_resWire_wget__410_BITS_67_TO_5_ETC___d6034 =
	     12'd3970 -
	     SEXT_resWire_wget__410_BITS_67_TO_57_416_MINUS_ETC___d6031 ;
  assign _7170_MINUS_fpu_madd_fState_S3_first__995_BITS__ETC___d2007 =
	     13'd7170 - fpu_madd_fState_S3$D_OUT[12:0] ;
  assign _7170_MINUS_fpu_madd_fState_S3_first__995_BITS__ETC___d2008 =
	     (_7170_MINUS_fpu_madd_fState_S3_first__995_BITS__ETC___d2007 ^
	      13'h1000) <=
	     13'd4096 ;
  assign _theResult____h164612 =
	     ((_3074_MINUS_SEXT_iFifo_first__087_BITS_167_TO_1_ETC___d3326 ^
	       12'h800) <
	      12'd2105) ?
	       result__h165225 :
	       ((value__h148921 == 25'd0) ? sfd__h144534 : 57'd1) ;
  assign _theResult____h203250 =
	     ((_3074_MINUS_SEXT_iFifo_first__087_BITS_102_TO_9_ETC___d4809 ^
	       12'h800) <
	      12'd2105) ?
	       result__h203863 :
	       ((value__h187559 == 25'd0) ? sfd__h183174 : 57'd1) ;
  assign _theResult____h242189 =
	     ((_3074_MINUS_SEXT_iFifo_first__087_BITS_37_TO_30_ETC___d4034 ^
	       12'h800) <
	      12'd2105) ?
	       result__h242802 :
	       ((value__h226498 == 25'd0) ? sfd__h222113 : 57'd1) ;
  assign _theResult____h269613 =
	     (value__h270233 == 54'd0) ? sfd__h262011 : 57'd1 ;
  assign _theResult____h287250 =
	     ((_3970_MINUS_SEXT_resWire_wget__410_BITS_67_TO_5_ETC___d6034 ^
	       12'h800) <
	      12'd2105) ?
	       result__h287863 :
	       _theResult____h269613 ;
  assign _theResult____h31574 =
	     (fpu_div_fState_S2$D_OUT[10:0] < 11'd58) ?
	       result__h31699 :
	       result__h31874 ;
  assign _theResult___exp__h142541 =
	     sfd__h142040[53] ?
	       ((fpu_madd_fState_S8$D_OUT[65:55] == 11'd2046) ?
		  11'd2047 :
		  din_inc___2_exp__h142626) :
	       IF_fpu_madd_fState_S8_first__960_BITS_65_TO_55_ETC___d2986 ;
  assign _theResult___exp__h163979 =
	     sfd__h163352[53] ?
	       ((_theResult___fst_exp__h163334 == 11'd2046) ?
		  11'd2047 :
		  din_inc___2_exp__h182467) :
	       ((_theResult___fst_exp__h163334 == 11'd0 &&
		 sfd__h163352[53:52] == 2'b01) ?
		  11'd1 :
		  _theResult___fst_exp__h163334) ;
  assign _theResult___exp__h173569 =
	     sfd__h172942[53] ?
	       ((_theResult___fst_exp__h172850 == 11'd2046) ?
		  11'd2047 :
		  din_inc___2_exp__h182502) :
	       ((_theResult___fst_exp__h172850 == 11'd0 &&
		 sfd__h172942[53:52] == 2'b01) ?
		  11'd1 :
		  _theResult___fst_exp__h172850) ;
  assign _theResult___exp__h182321 =
	     sfd__h181670[53] ?
	       ((_theResult___fst_exp__h181651 == 11'd2046) ?
		  11'd2047 :
		  din_inc___2_exp__h182528) :
	       ((_theResult___fst_exp__h181651 == 11'd0 &&
		 sfd__h181670[53:52] == 2'b01) ?
		  11'd1 :
		  _theResult___fst_exp__h181651) ;
  assign _theResult___exp__h202617 =
	     sfd__h201990[53] ?
	       ((_theResult___fst_exp__h201972 == 11'd2046) ?
		  11'd2047 :
		  din_inc___2_exp__h221105) :
	       ((_theResult___fst_exp__h201972 == 11'd0 &&
		 sfd__h201990[53:52] == 2'b01) ?
		  11'd1 :
		  _theResult___fst_exp__h201972) ;
  assign _theResult___exp__h212207 =
	     sfd__h211580[53] ?
	       ((_theResult___fst_exp__h211488 == 11'd2046) ?
		  11'd2047 :
		  din_inc___2_exp__h221140) :
	       ((_theResult___fst_exp__h211488 == 11'd0 &&
		 sfd__h211580[53:52] == 2'b01) ?
		  11'd1 :
		  _theResult___fst_exp__h211488) ;
  assign _theResult___exp__h220959 =
	     sfd__h220308[53] ?
	       ((_theResult___fst_exp__h220289 == 11'd2046) ?
		  11'd2047 :
		  din_inc___2_exp__h221166) :
	       ((_theResult___fst_exp__h220289 == 11'd0 &&
		 sfd__h220308[53:52] == 2'b01) ?
		  11'd1 :
		  _theResult___fst_exp__h220289) ;
  assign _theResult___exp__h241556 =
	     sfd__h240929[53] ?
	       ((_theResult___fst_exp__h240911 == 11'd2046) ?
		  11'd2047 :
		  din_inc___2_exp__h260044) :
	       ((_theResult___fst_exp__h240911 == 11'd0 &&
		 sfd__h240929[53:52] == 2'b01) ?
		  11'd1 :
		  _theResult___fst_exp__h240911) ;
  assign _theResult___exp__h251146 =
	     sfd__h250519[53] ?
	       ((_theResult___fst_exp__h250427 == 11'd2046) ?
		  11'd2047 :
		  din_inc___2_exp__h260079) :
	       ((_theResult___fst_exp__h250427 == 11'd0 &&
		 sfd__h250519[53:52] == 2'b01) ?
		  11'd1 :
		  _theResult___fst_exp__h250427) ;
  assign _theResult___exp__h259898 =
	     sfd__h259247[53] ?
	       ((_theResult___fst_exp__h259228 == 11'd2046) ?
		  11'd2047 :
		  din_inc___2_exp__h260105) :
	       ((_theResult___fst_exp__h259228 == 11'd0 &&
		 sfd__h259247[53:52] == 2'b01) ?
		  11'd1 :
		  _theResult___fst_exp__h259228) ;
  assign _theResult___exp__h278238 =
	     sfd__h277814[24] ?
	       ((_theResult___fst_exp__h277722 == 8'd254) ?
		  8'd255 :
		  din_inc___2_exp__h304759) :
	       ((_theResult___fst_exp__h277722 == 8'd0 &&
		 sfd__h277814[24:23] == 2'b01) ?
		  8'd1 :
		  _theResult___fst_exp__h277722) ;
  assign _theResult___exp__h286820 =
	     sfd__h286396[24] ?
	       ((_theResult___fst_exp__h286378 == 8'd254) ?
		  8'd255 :
		  din_inc___2_exp__h304785) :
	       ((_theResult___fst_exp__h286378 == 8'd0 &&
		 sfd__h286396[24:23] == 2'b01) ?
		  8'd1 :
		  _theResult___fst_exp__h286378) ;
  assign _theResult___exp__h296004 =
	     sfd__h295580[24] ?
	       ((_theResult___fst_exp__h295488 == 8'd254) ?
		  8'd255 :
		  din_inc___2_exp__h304820) :
	       ((_theResult___fst_exp__h295488 == 8'd0 &&
		 sfd__h295580[24:23] == 2'b01) ?
		  8'd1 :
		  _theResult___fst_exp__h295488) ;
  assign _theResult___exp__h304640 =
	     sfd__h304192[24] ?
	       ((_theResult___fst_exp__h304173 == 8'd254) ?
		  8'd255 :
		  din_inc___2_exp__h304846) :
	       ((_theResult___fst_exp__h304173 == 8'd0 &&
		 sfd__h304192[24:23] == 2'b01) ?
		  8'd1 :
		  _theResult___fst_exp__h304173) ;
  assign _theResult___exp__h42526 =
	     sfd__h42033[53] ?
	       ((fpu_div_fState_S4$D_OUT[64:54] == 11'd2046) ?
		  11'd2047 :
		  din_inc___2_exp__h42617) :
	       IF_fpu_div_fState_S4_first__73_BITS_64_TO_54_7_ETC___d907 ;
  assign _theResult___exp__h95909 =
	     sfd__h95416[53] ?
	       ((fpu_sqr_fState_S4$D_OUT[64:54] == 11'd2046) ?
		  11'd2047 :
		  din_inc___2_exp__h96000) :
	       IF_fpu_sqr_fState_S4_first__687_BITS_64_TO_54__ETC___d1721 ;
  assign _theResult___fst__h116827 =
	     { fpu_madd_fProd_S3_first__009_SRL_IF_7170_MINUS_ETC___d2012[105:1],
	       fpu_madd_fProd_S3_first__009_SRL_IF_7170_MINUS_ETC___d2012[0] |
	       sfdlsb__h116825 } ;
  assign _theResult___fst__h30373 =
	     IF_fpu_div_fOperands_S0_first__6_BITS_129_TO_1_ETC___d429 ?
	       value__h30601[10:0] :
	       11'd0 ;
  assign _theResult___fst__h43498 =
	     IF_rg_index_1_87_ULE_58_91_THEN_NOT_rg_b_92_EQ_ETC___d1009 ?
	       _theResult___fst__h43622 :
	       IF_rg_index_1_87_ULE_58_91_THEN_IF_rg_res_94_B_ETC___d1002 ;
  assign _theResult___fst__h43537 =
	     (rg_res[116] || rg_b == 116'd0) ? rg_b : b__h43630 ;
  assign _theResult___fst__h43622 =
	     (IF_rg_index_1_87_ULE_58_91_THEN_IF_rg_res_94_B_ETC___d1002 ==
	      116'd0) ?
	       IF_rg_index_1_87_ULE_58_91_THEN_IF_rg_res_94_B_ETC___d1002 :
	       b__h43734 ;
  assign _theResult___fst_exp__h130949 =
	     sfdBC__h115662[105] ?
	       _theResult___fst_exp__h130971 :
	       _theResult___fst_exp__h131034 ;
  assign _theResult___fst_exp__h130952 =
	     (sfdBC__h115662[105] &&
	      IF_IF_7170_MINUS_fpu_madd_fState_S3_first__995_ETC___d2031 ==
	      12'd1023) ?
	       11'd2046 :
	       _theResult___fst_exp__h130949 ;
  assign _theResult___fst_exp__h130971 =
	     (din_exp__h130866 == 11'd0) ? 11'd2 : din_exp__h130866 + 11'd1 ;
  assign _theResult___fst_exp__h130986 =
	     (din_exp__h130866 == 11'd0) ? 11'd1 : din_exp__h130866 ;
  assign _theResult___fst_exp__h131025 =
	     din_exp__h130866 -
	     { 4'd0,
	       IF_IF_7170_MINUS_fpu_madd_fState_S3_first__995_ETC___d2460 } ;
  assign _theResult___fst_exp__h131031 =
	     (!sfdBC__h115662[105] && !sfdBC__h115662[104] &&
	      !sfdBC__h115662[103] &&
	      !sfdBC__h115662[102] &&
	      !sfdBC__h115662[101] &&
	      !sfdBC__h115662[100] &&
	      !sfdBC__h115662[99] &&
	      !sfdBC__h115662[98] &&
	      !sfdBC__h115662[97] &&
	      !sfdBC__h115662[96] &&
	      !sfdBC__h115662[95] &&
	      !sfdBC__h115662[94] &&
	      !sfdBC__h115662[93] &&
	      !sfdBC__h115662[92] &&
	      !sfdBC__h115662[91] &&
	      !sfdBC__h115662[90] &&
	      !sfdBC__h115662[89] &&
	      !sfdBC__h115662[88] &&
	      !sfdBC__h115662[87] &&
	      !sfdBC__h115662[86] &&
	      !sfdBC__h115662[85] &&
	      !sfdBC__h115662[84] &&
	      !sfdBC__h115662[83] &&
	      !sfdBC__h115662[82] &&
	      !sfdBC__h115662[81] &&
	      !sfdBC__h115662[80] &&
	      !sfdBC__h115662[79] &&
	      !sfdBC__h115662[78] &&
	      !sfdBC__h115662[77] &&
	      !sfdBC__h115662[76] &&
	      !sfdBC__h115662[75] &&
	      !sfdBC__h115662[74] &&
	      !sfdBC__h115662[73] &&
	      !sfdBC__h115662[72] &&
	      !sfdBC__h115662[71] &&
	      !sfdBC__h115662[70] &&
	      !sfdBC__h115662[69] &&
	      !sfdBC__h115662[68] &&
	      !sfdBC__h115662[67] &&
	      !sfdBC__h115662[66] &&
	      !sfdBC__h115662[65] &&
	      !sfdBC__h115662[64] &&
	      !sfdBC__h115662[63] &&
	      !sfdBC__h115662[62] &&
	      !sfdBC__h115662[61] &&
	      !sfdBC__h115662[60] &&
	      !sfdBC__h115662[59] &&
	      !sfdBC__h115662[58] &&
	      !sfdBC__h115662[57] &&
	      !sfdBC__h115662[56] &&
	      !sfdBC__h115662[55] &&
	      !sfdBC__h115662[54] &&
	      !sfdBC__h115662[53] &&
	      !sfdBC__h115662[52] &&
	      !sfdBC__h115662[51] &&
	      !sfdBC__h115662[50] &&
	      !sfdBC__h115662[49] &&
	      !sfdBC__h115662[48] &&
	      !sfdBC__h115662[47] &&
	      !sfdBC__h115662[46] &&
	      !sfdBC__h115662[45] &&
	      !sfdBC__h115662[44] &&
	      !sfdBC__h115662[43] &&
	      !sfdBC__h115662[42] &&
	      !sfdBC__h115662[41] &&
	      !sfdBC__h115662[40] &&
	      !sfdBC__h115662[39] &&
	      !sfdBC__h115662[38] &&
	      !sfdBC__h115662[37] &&
	      !sfdBC__h115662[36] &&
	      !sfdBC__h115662[35] &&
	      !sfdBC__h115662[34] &&
	      !sfdBC__h115662[33] &&
	      !sfdBC__h115662[32] &&
	      !sfdBC__h115662[31] &&
	      !sfdBC__h115662[30] &&
	      !sfdBC__h115662[29] &&
	      !sfdBC__h115662[28] &&
	      !sfdBC__h115662[27] &&
	      !sfdBC__h115662[26] &&
	      !sfdBC__h115662[25] &&
	      !sfdBC__h115662[24] &&
	      !sfdBC__h115662[23] &&
	      !sfdBC__h115662[22] &&
	      !sfdBC__h115662[21] &&
	      !sfdBC__h115662[20] &&
	      !sfdBC__h115662[19] &&
	      !sfdBC__h115662[18] &&
	      !sfdBC__h115662[17] &&
	      !sfdBC__h115662[16] &&
	      !sfdBC__h115662[15] &&
	      !sfdBC__h115662[14] &&
	      !sfdBC__h115662[13] &&
	      !sfdBC__h115662[12] &&
	      !sfdBC__h115662[11] &&
	      !sfdBC__h115662[10] &&
	      !sfdBC__h115662[9] &&
	      !sfdBC__h115662[8] &&
	      !sfdBC__h115662[7] &&
	      !sfdBC__h115662[6] &&
	      !sfdBC__h115662[5] &&
	      !sfdBC__h115662[4] &&
	      !sfdBC__h115662[3] &&
	      !sfdBC__h115662[2] &&
	      !sfdBC__h115662[1] &&
	      !sfdBC__h115662[0] ||
	      !_0_CONCAT_IF_IF_7170_MINUS_fpu_madd_fState_S3_f_ETC___d2463) ?
	       11'd0 :
	       _theResult___fst_exp__h131025 ;
  assign _theResult___fst_exp__h131034 =
	     (!sfdBC__h115662[105] && sfdBC__h115662[104]) ?
	       _theResult___fst_exp__h130986 :
	       _theResult___fst_exp__h131031 ;
  assign _theResult___fst_exp__h141375 =
	     sfd__h133119[56] ?
	       _theResult___fst_exp__h141397 :
	       _theResult___fst_exp__h141460 ;
  assign _theResult___fst_exp__h141378 =
	     (sfd__h133119[56] &&
	      IF_fpu_madd_fState_S7_first__651_BITS_126_TO_1_ETC___d2668 ==
	      12'd1023) ?
	       11'd2046 :
	       _theResult___fst_exp__h141375 ;
  assign _theResult___fst_exp__h141397 =
	     (value__h141307[10:0] == 11'd0) ?
	       11'd2 :
	       value__h141307[10:0] + 11'd1 ;
  assign _theResult___fst_exp__h141412 =
	     (value__h141307[10:0] == 11'd0) ? 11'd1 : value__h141307[10:0] ;
  assign _theResult___fst_exp__h141451 =
	     value__h141307[10:0] -
	     { 5'd0,
	       IF_IF_fpu_madd_fState_S7_first__651_BIT_128_65_ETC___d2901 } ;
  assign _theResult___fst_exp__h141457 =
	     (!sfd__h133119[56] && !sfd__h133119[55] && !sfd__h133119[54] &&
	      !sfd__h133119[53] &&
	      !sfd__h133119[52] &&
	      !sfd__h133119[51] &&
	      !sfd__h133119[50] &&
	      !sfd__h133119[49] &&
	      !sfd__h133119[48] &&
	      !sfd__h133119[47] &&
	      !sfd__h133119[46] &&
	      !sfd__h133119[45] &&
	      !sfd__h133119[44] &&
	      !sfd__h133119[43] &&
	      !sfd__h133119[42] &&
	      !sfd__h133119[41] &&
	      !sfd__h133119[40] &&
	      !sfd__h133119[39] &&
	      !sfd__h133119[38] &&
	      !sfd__h133119[37] &&
	      !sfd__h133119[36] &&
	      !sfd__h133119[35] &&
	      !sfd__h133119[34] &&
	      !sfd__h133119[33] &&
	      !sfd__h133119[32] &&
	      !sfd__h133119[31] &&
	      !sfd__h133119[30] &&
	      !sfd__h133119[29] &&
	      !sfd__h133119[28] &&
	      !sfd__h133119[27] &&
	      !sfd__h133119[26] &&
	      !sfd__h133119[25] &&
	      !sfd__h133119[24] &&
	      !sfd__h133119[23] &&
	      !sfd__h133119[22] &&
	      !sfd__h133119[21] &&
	      !sfd__h133119[20] &&
	      !sfd__h133119[19] &&
	      !sfd__h133119[18] &&
	      !sfd__h133119[17] &&
	      !sfd__h133119[16] &&
	      !sfd__h133119[15] &&
	      !sfd__h133119[14] &&
	      !sfd__h133119[13] &&
	      !sfd__h133119[12] &&
	      !sfd__h133119[11] &&
	      !sfd__h133119[10] &&
	      !sfd__h133119[9] &&
	      !sfd__h133119[8] &&
	      !sfd__h133119[7] &&
	      !sfd__h133119[6] &&
	      !sfd__h133119[5] &&
	      !sfd__h133119[4] &&
	      !sfd__h133119[3] &&
	      !sfd__h133119[2] &&
	      !sfd__h133119[1] &&
	      !sfd__h133119[0] ||
	      !_0_CONCAT_IF_IF_fpu_madd_fState_S7_first__651_B_ETC___d2904) ?
	       11'd0 :
	       _theResult___fst_exp__h141451 ;
  assign _theResult___fst_exp__h141460 =
	     (!sfd__h133119[56] && sfd__h133119[55]) ?
	       _theResult___fst_exp__h141412 :
	       _theResult___fst_exp__h141457 ;
  assign _theResult___fst_exp__h163325 =
	     11'd897 -
	     { 5'd0,
	       IF_iFifo_first__087_BITS_167_TO_160_130_EQ_0_1_ETC___d3271 } ;
  assign _theResult___fst_exp__h163331 =
	     (iFifo$D_OUT[167:160] == 8'd0 && !iFifo$D_OUT[159] &&
	      NOT_iFifo_first__087_BIT_158_142_202_AND_NOT_i_ETC___d3244 ||
	      !_0_CONCAT_IF_iFifo_first__087_BITS_167_TO_160_1_ETC___d3273) ?
	       11'd0 :
	       _theResult___fst_exp__h163325 ;
  assign _theResult___fst_exp__h163334 =
	     (iFifo$D_OUT[167:160] == 8'd0) ?
	       _theResult___fst_exp__h163331 :
	       11'd897 ;
  assign _theResult___fst_exp__h164060 =
	     (_theResult___fst_exp__h163334 == 11'd2047) ?
	       _theResult___fst_exp__h163334 :
	       _theResult___fst_exp__h164057 ;
  assign _theResult___fst_exp__h172850 =
	     _theResult____h164612[56] ?
	       11'd2 :
	       _theResult___fst_exp__h172924 ;
  assign _theResult___fst_exp__h172915 =
	     11'd0 -
	     { 5'd0,
	       IF_IF_3074_MINUS_SEXT_iFifo_first__087_BITS_16_ETC___d3572 } ;
  assign _theResult___fst_exp__h172921 =
	     (!_theResult____h164612[56] && !_theResult____h164612[55] &&
	      !_theResult____h164612[54] &&
	      !_theResult____h164612[53] &&
	      !_theResult____h164612[52] &&
	      !_theResult____h164612[51] &&
	      !_theResult____h164612[50] &&
	      !_theResult____h164612[49] &&
	      !_theResult____h164612[48] &&
	      !_theResult____h164612[47] &&
	      !_theResult____h164612[46] &&
	      !_theResult____h164612[45] &&
	      !_theResult____h164612[44] &&
	      !_theResult____h164612[43] &&
	      !_theResult____h164612[42] &&
	      !_theResult____h164612[41] &&
	      !_theResult____h164612[40] &&
	      !_theResult____h164612[39] &&
	      !_theResult____h164612[38] &&
	      !_theResult____h164612[37] &&
	      !_theResult____h164612[36] &&
	      !_theResult____h164612[35] &&
	      !_theResult____h164612[34] &&
	      !_theResult____h164612[33] &&
	      !_theResult____h164612[32] &&
	      !_theResult____h164612[31] &&
	      !_theResult____h164612[30] &&
	      !_theResult____h164612[29] &&
	      !_theResult____h164612[28] &&
	      !_theResult____h164612[27] &&
	      !_theResult____h164612[26] &&
	      !_theResult____h164612[25] &&
	      !_theResult____h164612[24] &&
	      !_theResult____h164612[23] &&
	      !_theResult____h164612[22] &&
	      !_theResult____h164612[21] &&
	      !_theResult____h164612[20] &&
	      !_theResult____h164612[19] &&
	      !_theResult____h164612[18] &&
	      !_theResult____h164612[17] &&
	      !_theResult____h164612[16] &&
	      !_theResult____h164612[15] &&
	      !_theResult____h164612[14] &&
	      !_theResult____h164612[13] &&
	      !_theResult____h164612[12] &&
	      !_theResult____h164612[11] &&
	      !_theResult____h164612[10] &&
	      !_theResult____h164612[9] &&
	      !_theResult____h164612[8] &&
	      !_theResult____h164612[7] &&
	      !_theResult____h164612[6] &&
	      !_theResult____h164612[5] &&
	      !_theResult____h164612[4] &&
	      !_theResult____h164612[3] &&
	      !_theResult____h164612[2] &&
	      !_theResult____h164612[1] &&
	      !_theResult____h164612[0] ||
	      !_0_CONCAT_IF_IF_3074_MINUS_SEXT_iFifo_first__08_ETC___d3574) ?
	       11'd0 :
	       _theResult___fst_exp__h172915 ;
  assign _theResult___fst_exp__h172924 =
	     (!_theResult____h164612[56] && _theResult____h164612[55]) ?
	       11'd1 :
	       _theResult___fst_exp__h172921 ;
  assign _theResult___fst_exp__h173650 =
	     (_theResult___fst_exp__h172850 == 11'd2047) ?
	       _theResult___fst_exp__h172850 :
	       _theResult___fst_exp__h173647 ;
  assign _theResult___fst_exp__h181603 =
	     (SEXT_iFifo_first__087_BITS_167_TO_160_130_MINU_ETC__q36[10:0] ==
	      11'd0) ?
	       11'd1 :
	       SEXT_iFifo_first__087_BITS_167_TO_160_130_MINU_ETC__q36[10:0] ;
  assign _theResult___fst_exp__h181642 =
	     SEXT_iFifo_first__087_BITS_167_TO_160_130_MINU_ETC__q36[10:0] -
	     { 5'd0,
	       IF_iFifo_first__087_BITS_167_TO_160_130_EQ_0_1_ETC___d3271 } ;
  assign _theResult___fst_exp__h181648 =
	     (iFifo$D_OUT[167:160] == 8'd0 && !iFifo$D_OUT[159] &&
	      NOT_iFifo_first__087_BIT_158_142_202_AND_NOT_i_ETC___d3244 ||
	      !_0_CONCAT_IF_iFifo_first__087_BITS_167_TO_160_1_ETC___d3624) ?
	       11'd0 :
	       _theResult___fst_exp__h181642 ;
  assign _theResult___fst_exp__h181651 =
	     (iFifo$D_OUT[167:160] == 8'd0) ?
	       _theResult___fst_exp__h181648 :
	       _theResult___fst_exp__h181603 ;
  assign _theResult___fst_exp__h182402 =
	     (_theResult___fst_exp__h181651 == 11'd2047) ?
	       _theResult___fst_exp__h181651 :
	       _theResult___fst_exp__h182399 ;
  assign _theResult___fst_exp__h182411 =
	     (iFifo$D_OUT[167:160] == 8'd0) ?
	       (_3970_MINUS_0_CONCAT_IF_iFifo_first__087_BIT_15_ETC___d3189 ?
		  _theResult___snd_fst_exp__h164063 :
		  _theResult___fst_exp__h148289) :
	       (SEXT_iFifo_first__087_BITS_167_TO_160_130_MINU_ETC___d3324 ?
		  _theResult___snd_fst_exp__h182405 :
		  _theResult___fst_exp__h148289) ;
  assign _theResult___fst_exp__h182414 =
	     (iFifo$D_OUT[167:160] == 8'd0 && iFifo$D_OUT[159:137] == 23'd0) ?
	       11'd0 :
	       _theResult___fst_exp__h182411 ;
  assign _theResult___fst_exp__h201963 =
	     11'd897 -
	     { 5'd0,
	       IF_iFifo_first__087_BITS_102_TO_95_625_EQ_0_63_ETC___d4757 } ;
  assign _theResult___fst_exp__h201969 =
	     (iFifo$D_OUT[102:95] == 8'd0 && !iFifo$D_OUT[94] &&
	      NOT_iFifo_first__087_BIT_93_637_688_AND_NOT_iF_ETC___d4730 ||
	      !_0_CONCAT_IF_iFifo_first__087_BITS_102_TO_95_62_ETC___d4759) ?
	       11'd0 :
	       _theResult___fst_exp__h201963 ;
  assign _theResult___fst_exp__h201972 =
	     (iFifo$D_OUT[102:95] == 8'd0) ?
	       _theResult___fst_exp__h201969 :
	       11'd897 ;
  assign _theResult___fst_exp__h202698 =
	     (_theResult___fst_exp__h201972 == 11'd2047) ?
	       _theResult___fst_exp__h201972 :
	       _theResult___fst_exp__h202695 ;
  assign _theResult___fst_exp__h211488 =
	     _theResult____h203250[56] ?
	       11'd2 :
	       _theResult___fst_exp__h211562 ;
  assign _theResult___fst_exp__h211553 =
	     11'd0 -
	     { 5'd0,
	       IF_IF_3074_MINUS_SEXT_iFifo_first__087_BITS_10_ETC___d5055 } ;
  assign _theResult___fst_exp__h211559 =
	     (!_theResult____h203250[56] && !_theResult____h203250[55] &&
	      !_theResult____h203250[54] &&
	      !_theResult____h203250[53] &&
	      !_theResult____h203250[52] &&
	      !_theResult____h203250[51] &&
	      !_theResult____h203250[50] &&
	      !_theResult____h203250[49] &&
	      !_theResult____h203250[48] &&
	      !_theResult____h203250[47] &&
	      !_theResult____h203250[46] &&
	      !_theResult____h203250[45] &&
	      !_theResult____h203250[44] &&
	      !_theResult____h203250[43] &&
	      !_theResult____h203250[42] &&
	      !_theResult____h203250[41] &&
	      !_theResult____h203250[40] &&
	      !_theResult____h203250[39] &&
	      !_theResult____h203250[38] &&
	      !_theResult____h203250[37] &&
	      !_theResult____h203250[36] &&
	      !_theResult____h203250[35] &&
	      !_theResult____h203250[34] &&
	      !_theResult____h203250[33] &&
	      !_theResult____h203250[32] &&
	      !_theResult____h203250[31] &&
	      !_theResult____h203250[30] &&
	      !_theResult____h203250[29] &&
	      !_theResult____h203250[28] &&
	      !_theResult____h203250[27] &&
	      !_theResult____h203250[26] &&
	      !_theResult____h203250[25] &&
	      !_theResult____h203250[24] &&
	      !_theResult____h203250[23] &&
	      !_theResult____h203250[22] &&
	      !_theResult____h203250[21] &&
	      !_theResult____h203250[20] &&
	      !_theResult____h203250[19] &&
	      !_theResult____h203250[18] &&
	      !_theResult____h203250[17] &&
	      !_theResult____h203250[16] &&
	      !_theResult____h203250[15] &&
	      !_theResult____h203250[14] &&
	      !_theResult____h203250[13] &&
	      !_theResult____h203250[12] &&
	      !_theResult____h203250[11] &&
	      !_theResult____h203250[10] &&
	      !_theResult____h203250[9] &&
	      !_theResult____h203250[8] &&
	      !_theResult____h203250[7] &&
	      !_theResult____h203250[6] &&
	      !_theResult____h203250[5] &&
	      !_theResult____h203250[4] &&
	      !_theResult____h203250[3] &&
	      !_theResult____h203250[2] &&
	      !_theResult____h203250[1] &&
	      !_theResult____h203250[0] ||
	      !_0_CONCAT_IF_IF_3074_MINUS_SEXT_iFifo_first__08_ETC___d5057) ?
	       11'd0 :
	       _theResult___fst_exp__h211553 ;
  assign _theResult___fst_exp__h211562 =
	     (!_theResult____h203250[56] && _theResult____h203250[55]) ?
	       11'd1 :
	       _theResult___fst_exp__h211559 ;
  assign _theResult___fst_exp__h212288 =
	     (_theResult___fst_exp__h211488 == 11'd2047) ?
	       _theResult___fst_exp__h211488 :
	       _theResult___fst_exp__h212285 ;
  assign _theResult___fst_exp__h220241 =
	     (SEXT_iFifo_first__087_BITS_102_TO_95_625_MINUS_ETC__q96[10:0] ==
	      11'd0) ?
	       11'd1 :
	       SEXT_iFifo_first__087_BITS_102_TO_95_625_MINUS_ETC__q96[10:0] ;
  assign _theResult___fst_exp__h220280 =
	     SEXT_iFifo_first__087_BITS_102_TO_95_625_MINUS_ETC__q96[10:0] -
	     { 5'd0,
	       IF_iFifo_first__087_BITS_102_TO_95_625_EQ_0_63_ETC___d4757 } ;
  assign _theResult___fst_exp__h220286 =
	     (iFifo$D_OUT[102:95] == 8'd0 && !iFifo$D_OUT[94] &&
	      NOT_iFifo_first__087_BIT_93_637_688_AND_NOT_iF_ETC___d4730 ||
	      !_0_CONCAT_IF_iFifo_first__087_BITS_102_TO_95_62_ETC___d5107) ?
	       11'd0 :
	       _theResult___fst_exp__h220280 ;
  assign _theResult___fst_exp__h220289 =
	     (iFifo$D_OUT[102:95] == 8'd0) ?
	       _theResult___fst_exp__h220286 :
	       _theResult___fst_exp__h220241 ;
  assign _theResult___fst_exp__h221040 =
	     (_theResult___fst_exp__h220289 == 11'd2047) ?
	       _theResult___fst_exp__h220289 :
	       _theResult___fst_exp__h221037 ;
  assign _theResult___fst_exp__h221049 =
	     (iFifo$D_OUT[102:95] == 8'd0) ?
	       (_3970_MINUS_0_CONCAT_IF_iFifo_first__087_BIT_94_ETC___d4684 ?
		  _theResult___snd_fst_exp__h202701 :
		  _theResult___fst_exp__h186929) :
	       (SEXT_iFifo_first__087_BITS_102_TO_95_625_MINUS_ETC___d4807 ?
		  _theResult___snd_fst_exp__h221043 :
		  _theResult___fst_exp__h186929) ;
  assign _theResult___fst_exp__h221052 =
	     (iFifo$D_OUT[102:95] == 8'd0 && iFifo$D_OUT[94:72] == 23'd0) ?
	       11'd0 :
	       _theResult___fst_exp__h221049 ;
  assign _theResult___fst_exp__h240902 =
	     11'd897 -
	     { 5'd0,
	       IF_iFifo_first__087_BITS_37_TO_30_850_EQ_0_856_ETC___d3982 } ;
  assign _theResult___fst_exp__h240908 =
	     (iFifo$D_OUT[37:30] == 8'd0 && !iFifo$D_OUT[29] &&
	      NOT_iFifo_first__087_BIT_28_862_913_AND_NOT_iF_ETC___d3955 ||
	      !_0_CONCAT_IF_iFifo_first__087_BITS_37_TO_30_850_ETC___d3984) ?
	       11'd0 :
	       _theResult___fst_exp__h240902 ;
  assign _theResult___fst_exp__h240911 =
	     (iFifo$D_OUT[37:30] == 8'd0) ?
	       _theResult___fst_exp__h240908 :
	       11'd897 ;
  assign _theResult___fst_exp__h241637 =
	     (_theResult___fst_exp__h240911 == 11'd2047) ?
	       _theResult___fst_exp__h240911 :
	       _theResult___fst_exp__h241634 ;
  assign _theResult___fst_exp__h250427 =
	     _theResult____h242189[56] ?
	       11'd2 :
	       _theResult___fst_exp__h250501 ;
  assign _theResult___fst_exp__h250492 =
	     11'd0 -
	     { 5'd0,
	       IF_IF_3074_MINUS_SEXT_iFifo_first__087_BITS_37_ETC___d4280 } ;
  assign _theResult___fst_exp__h250498 =
	     (!_theResult____h242189[56] && !_theResult____h242189[55] &&
	      !_theResult____h242189[54] &&
	      !_theResult____h242189[53] &&
	      !_theResult____h242189[52] &&
	      !_theResult____h242189[51] &&
	      !_theResult____h242189[50] &&
	      !_theResult____h242189[49] &&
	      !_theResult____h242189[48] &&
	      !_theResult____h242189[47] &&
	      !_theResult____h242189[46] &&
	      !_theResult____h242189[45] &&
	      !_theResult____h242189[44] &&
	      !_theResult____h242189[43] &&
	      !_theResult____h242189[42] &&
	      !_theResult____h242189[41] &&
	      !_theResult____h242189[40] &&
	      !_theResult____h242189[39] &&
	      !_theResult____h242189[38] &&
	      !_theResult____h242189[37] &&
	      !_theResult____h242189[36] &&
	      !_theResult____h242189[35] &&
	      !_theResult____h242189[34] &&
	      !_theResult____h242189[33] &&
	      !_theResult____h242189[32] &&
	      !_theResult____h242189[31] &&
	      !_theResult____h242189[30] &&
	      !_theResult____h242189[29] &&
	      !_theResult____h242189[28] &&
	      !_theResult____h242189[27] &&
	      !_theResult____h242189[26] &&
	      !_theResult____h242189[25] &&
	      !_theResult____h242189[24] &&
	      !_theResult____h242189[23] &&
	      !_theResult____h242189[22] &&
	      !_theResult____h242189[21] &&
	      !_theResult____h242189[20] &&
	      !_theResult____h242189[19] &&
	      !_theResult____h242189[18] &&
	      !_theResult____h242189[17] &&
	      !_theResult____h242189[16] &&
	      !_theResult____h242189[15] &&
	      !_theResult____h242189[14] &&
	      !_theResult____h242189[13] &&
	      !_theResult____h242189[12] &&
	      !_theResult____h242189[11] &&
	      !_theResult____h242189[10] &&
	      !_theResult____h242189[9] &&
	      !_theResult____h242189[8] &&
	      !_theResult____h242189[7] &&
	      !_theResult____h242189[6] &&
	      !_theResult____h242189[5] &&
	      !_theResult____h242189[4] &&
	      !_theResult____h242189[3] &&
	      !_theResult____h242189[2] &&
	      !_theResult____h242189[1] &&
	      !_theResult____h242189[0] ||
	      !_0_CONCAT_IF_IF_3074_MINUS_SEXT_iFifo_first__08_ETC___d4282) ?
	       11'd0 :
	       _theResult___fst_exp__h250492 ;
  assign _theResult___fst_exp__h250501 =
	     (!_theResult____h242189[56] && _theResult____h242189[55]) ?
	       11'd1 :
	       _theResult___fst_exp__h250498 ;
  assign _theResult___fst_exp__h251227 =
	     (_theResult___fst_exp__h250427 == 11'd2047) ?
	       _theResult___fst_exp__h250427 :
	       _theResult___fst_exp__h251224 ;
  assign _theResult___fst_exp__h259180 =
	     (SEXT_iFifo_first__087_BITS_37_TO_30_850_MINUS__ETC__q63[10:0] ==
	      11'd0) ?
	       11'd1 :
	       SEXT_iFifo_first__087_BITS_37_TO_30_850_MINUS__ETC__q63[10:0] ;
  assign _theResult___fst_exp__h259219 =
	     SEXT_iFifo_first__087_BITS_37_TO_30_850_MINUS__ETC__q63[10:0] -
	     { 5'd0,
	       IF_iFifo_first__087_BITS_37_TO_30_850_EQ_0_856_ETC___d3982 } ;
  assign _theResult___fst_exp__h259225 =
	     (iFifo$D_OUT[37:30] == 8'd0 && !iFifo$D_OUT[29] &&
	      NOT_iFifo_first__087_BIT_28_862_913_AND_NOT_iF_ETC___d3955 ||
	      !_0_CONCAT_IF_iFifo_first__087_BITS_37_TO_30_850_ETC___d4332) ?
	       11'd0 :
	       _theResult___fst_exp__h259219 ;
  assign _theResult___fst_exp__h259228 =
	     (iFifo$D_OUT[37:30] == 8'd0) ?
	       _theResult___fst_exp__h259225 :
	       _theResult___fst_exp__h259180 ;
  assign _theResult___fst_exp__h259979 =
	     (_theResult___fst_exp__h259228 == 11'd2047) ?
	       _theResult___fst_exp__h259228 :
	       _theResult___fst_exp__h259976 ;
  assign _theResult___fst_exp__h259988 =
	     (iFifo$D_OUT[37:30] == 8'd0) ?
	       (_3970_MINUS_0_CONCAT_IF_iFifo_first__087_BIT_29_ETC___d3909 ?
		  _theResult___snd_fst_exp__h241640 :
		  _theResult___fst_exp__h225868) :
	       (SEXT_iFifo_first__087_BITS_37_TO_30_850_MINUS__ETC___d4032 ?
		  _theResult___snd_fst_exp__h259982 :
		  _theResult___fst_exp__h225868) ;
  assign _theResult___fst_exp__h259991 =
	     (iFifo$D_OUT[37:30] == 8'd0 && iFifo$D_OUT[29:7] == 23'd0) ?
	       11'd0 :
	       _theResult___fst_exp__h259988 ;
  assign _theResult___fst_exp__h277722 =
	     _theResult____h269613[56] ?
	       8'd2 :
	       _theResult___fst_exp__h277796 ;
  assign _theResult___fst_exp__h277787 =
	     8'd0 -
	     { 2'd0,
	       IF_IF_0b0_CONCAT_NOT_resWire_wget__410_BITS_67_ETC___d5767 } ;
  assign _theResult___fst_exp__h277793 =
	     (!_theResult____h269613[56] && !_theResult____h269613[55] &&
	      !_theResult____h269613[54] &&
	      !_theResult____h269613[53] &&
	      !_theResult____h269613[52] &&
	      !_theResult____h269613[51] &&
	      !_theResult____h269613[50] &&
	      !_theResult____h269613[49] &&
	      !_theResult____h269613[48] &&
	      !_theResult____h269613[47] &&
	      !_theResult____h269613[46] &&
	      !_theResult____h269613[45] &&
	      !_theResult____h269613[44] &&
	      !_theResult____h269613[43] &&
	      !_theResult____h269613[42] &&
	      !_theResult____h269613[41] &&
	      !_theResult____h269613[40] &&
	      !_theResult____h269613[39] &&
	      !_theResult____h269613[38] &&
	      !_theResult____h269613[37] &&
	      !_theResult____h269613[36] &&
	      !_theResult____h269613[35] &&
	      !_theResult____h269613[34] &&
	      !_theResult____h269613[33] &&
	      !_theResult____h269613[32] &&
	      !_theResult____h269613[31] &&
	      !_theResult____h269613[30] &&
	      !_theResult____h269613[29] &&
	      !_theResult____h269613[28] &&
	      !_theResult____h269613[27] &&
	      !_theResult____h269613[26] &&
	      !_theResult____h269613[25] &&
	      !_theResult____h269613[24] &&
	      !_theResult____h269613[23] &&
	      !_theResult____h269613[22] &&
	      !_theResult____h269613[21] &&
	      !_theResult____h269613[20] &&
	      !_theResult____h269613[19] &&
	      !_theResult____h269613[18] &&
	      !_theResult____h269613[17] &&
	      !_theResult____h269613[16] &&
	      !_theResult____h269613[15] &&
	      !_theResult____h269613[14] &&
	      !_theResult____h269613[13] &&
	      !_theResult____h269613[12] &&
	      !_theResult____h269613[11] &&
	      !_theResult____h269613[10] &&
	      !_theResult____h269613[9] &&
	      !_theResult____h269613[8] &&
	      !_theResult____h269613[7] &&
	      !_theResult____h269613[6] &&
	      !_theResult____h269613[5] &&
	      !_theResult____h269613[4] &&
	      !_theResult____h269613[3] &&
	      !_theResult____h269613[2] &&
	      !_theResult____h269613[1] &&
	      !_theResult____h269613[0] ||
	      !_0_CONCAT_IF_IF_0b0_CONCAT_NOT_resWire_wget__41_ETC___d5769) ?
	       8'd0 :
	       _theResult___fst_exp__h277787 ;
  assign _theResult___fst_exp__h277796 =
	     (!_theResult____h269613[56] && _theResult____h269613[55]) ?
	       8'd1 :
	       _theResult___fst_exp__h277793 ;
  assign _theResult___fst_exp__h278319 =
	     (_theResult___fst_exp__h277722 == 8'd255) ?
	       _theResult___fst_exp__h277722 :
	       _theResult___fst_exp__h278316 ;
  assign _theResult___fst_exp__h286369 =
	     8'd129 -
	     { 2'd0,
	       IF_resWire_wget__410_BITS_67_TO_57_416_EQ_0_42_ETC___d5982 } ;
  assign _theResult___fst_exp__h286375 =
	     (resWire$wget[67:57] == 11'd0 &&
	      NOT_resWire_wget__410_BIT_56_426_825_AND_NOT_r_ETC___d5927 ||
	      !_0_CONCAT_IF_resWire_wget__410_BITS_67_TO_57_41_ETC___d5984) ?
	       8'd0 :
	       _theResult___fst_exp__h286369 ;
  assign _theResult___fst_exp__h286378 =
	     (resWire$wget[67:57] == 11'd0) ?
	       _theResult___fst_exp__h286375 :
	       8'd129 ;
  assign _theResult___fst_exp__h286901 =
	     (_theResult___fst_exp__h286378 == 8'd255) ?
	       _theResult___fst_exp__h286378 :
	       _theResult___fst_exp__h286898 ;
  assign _theResult___fst_exp__h295488 =
	     _theResult____h287250[56] ?
	       8'd2 :
	       _theResult___fst_exp__h295562 ;
  assign _theResult___fst_exp__h295553 =
	     8'd0 -
	     { 2'd0,
	       IF_IF_3970_MINUS_SEXT_resWire_wget__410_BITS_6_ETC___d6278 } ;
  assign _theResult___fst_exp__h295559 =
	     (!_theResult____h287250[56] && !_theResult____h287250[55] &&
	      !_theResult____h287250[54] &&
	      !_theResult____h287250[53] &&
	      !_theResult____h287250[52] &&
	      !_theResult____h287250[51] &&
	      !_theResult____h287250[50] &&
	      !_theResult____h287250[49] &&
	      !_theResult____h287250[48] &&
	      !_theResult____h287250[47] &&
	      !_theResult____h287250[46] &&
	      !_theResult____h287250[45] &&
	      !_theResult____h287250[44] &&
	      !_theResult____h287250[43] &&
	      !_theResult____h287250[42] &&
	      !_theResult____h287250[41] &&
	      !_theResult____h287250[40] &&
	      !_theResult____h287250[39] &&
	      !_theResult____h287250[38] &&
	      !_theResult____h287250[37] &&
	      !_theResult____h287250[36] &&
	      !_theResult____h287250[35] &&
	      !_theResult____h287250[34] &&
	      !_theResult____h287250[33] &&
	      !_theResult____h287250[32] &&
	      !_theResult____h287250[31] &&
	      !_theResult____h287250[30] &&
	      !_theResult____h287250[29] &&
	      !_theResult____h287250[28] &&
	      !_theResult____h287250[27] &&
	      !_theResult____h287250[26] &&
	      !_theResult____h287250[25] &&
	      !_theResult____h287250[24] &&
	      !_theResult____h287250[23] &&
	      !_theResult____h287250[22] &&
	      !_theResult____h287250[21] &&
	      !_theResult____h287250[20] &&
	      !_theResult____h287250[19] &&
	      !_theResult____h287250[18] &&
	      !_theResult____h287250[17] &&
	      !_theResult____h287250[16] &&
	      !_theResult____h287250[15] &&
	      !_theResult____h287250[14] &&
	      !_theResult____h287250[13] &&
	      !_theResult____h287250[12] &&
	      !_theResult____h287250[11] &&
	      !_theResult____h287250[10] &&
	      !_theResult____h287250[9] &&
	      !_theResult____h287250[8] &&
	      !_theResult____h287250[7] &&
	      !_theResult____h287250[6] &&
	      !_theResult____h287250[5] &&
	      !_theResult____h287250[4] &&
	      !_theResult____h287250[3] &&
	      !_theResult____h287250[2] &&
	      !_theResult____h287250[1] &&
	      !_theResult____h287250[0] ||
	      !_0_CONCAT_IF_IF_3970_MINUS_SEXT_resWire_wget__4_ETC___d6280) ?
	       8'd0 :
	       _theResult___fst_exp__h295553 ;
  assign _theResult___fst_exp__h295562 =
	     (!_theResult____h287250[56] && _theResult____h287250[55]) ?
	       8'd1 :
	       _theResult___fst_exp__h295559 ;
  assign _theResult___fst_exp__h296085 =
	     (_theResult___fst_exp__h295488 == 8'd255) ?
	       _theResult___fst_exp__h295488 :
	       _theResult___fst_exp__h296082 ;
  assign _theResult___fst_exp__h304125 =
	     (SEXT_resWire_wget__410_BITS_67_TO_57_416_MINUS_ETC__q138[7:0] ==
	      8'd0) ?
	       8'd1 :
	       SEXT_resWire_wget__410_BITS_67_TO_57_416_MINUS_ETC__q138[7:0] ;
  assign _theResult___fst_exp__h304164 =
	     SEXT_resWire_wget__410_BITS_67_TO_57_416_MINUS_ETC__q138[7:0] -
	     { 2'd0,
	       IF_resWire_wget__410_BITS_67_TO_57_416_EQ_0_42_ETC___d5982 } ;
  assign _theResult___fst_exp__h304170 =
	     (resWire$wget[67:57] == 11'd0 &&
	      NOT_resWire_wget__410_BIT_56_426_825_AND_NOT_r_ETC___d5927 ||
	      !_0_CONCAT_IF_resWire_wget__410_BITS_67_TO_57_41_ETC___d6333) ?
	       8'd0 :
	       _theResult___fst_exp__h304164 ;
  assign _theResult___fst_exp__h304173 =
	     (resWire$wget[67:57] == 11'd0) ?
	       _theResult___fst_exp__h304170 :
	       _theResult___fst_exp__h304125 ;
  assign _theResult___fst_exp__h304721 =
	     (_theResult___fst_exp__h304173 == 8'd255) ?
	       _theResult___fst_exp__h304173 :
	       _theResult___fst_exp__h304718 ;
  assign _theResult___fst_exp__h304730 =
	     (resWire$wget[67:57] == 11'd0) ?
	       (_3074_MINUS_0_CONCAT_IF_resWire_wget__410_BIT_5_ETC___d5532 ?
		  _theResult___snd_fst_exp__h286904 :
		  _theResult___fst_exp__h269595) :
	       (SEXT_resWire_wget__410_BITS_67_TO_57_416_MINUS_ETC___d6032 ?
		  _theResult___snd_fst_exp__h304724 :
		  _theResult___fst_exp__h269595) ;
  assign _theResult___fst_exp__h304733 =
	     (resWire$wget[67:57] == 11'd0 && resWire$wget[56:5] == 52'd0) ?
	       8'd0 :
	       _theResult___fst_exp__h304730 ;
  assign _theResult___fst_exp__h41335 =
	     fpu_div_fState_S3$D_OUT[120:110] - 11'd1 ;
  assign _theResult___fst_exp__h41338 =
	     (fpu_div_fState_S3$D_OUT[57:56] == 2'b0) ?
	       _theResult___fst_exp__h41335 :
	       11'd2046 ;
  assign _theResult___fst_exp__h41341 =
	     (fpu_div_fState_S3$D_OUT[120:110] == 11'd2047) ?
	       _theResult___fst_exp__h41338 :
	       fpu_div_fState_S3$D_OUT[120:110] ;
  assign _theResult___fst_exp__h41384 =
	     sfdin__h33169[57] ?
	       _theResult___fst_exp__h41407 :
	       _theResult___fst_exp__h41471 ;
  assign _theResult___fst_exp__h41387 =
	     (sfdin__h33169[57] &&
	      IF_IF_fpu_div_fState_S3_first__16_BITS_120_TO__ETC___d573 ==
	      12'd1023) ?
	       11'd2046 :
	       _theResult___fst_exp__h41384 ;
  assign _theResult___fst_exp__h41407 =
	     (_theResult___fst_exp__h41341 == 11'd0) ?
	       11'd2 :
	       _theResult___fst_exp__h41341 + 11'd1 ;
  assign _theResult___fst_exp__h41423 =
	     (_theResult___fst_exp__h41341 == 11'd0) ?
	       11'd1 :
	       _theResult___fst_exp__h41341 ;
  assign _theResult___fst_exp__h41462 =
	     _theResult___fst_exp__h41341 -
	     { 5'd0,
	       IF_IF_fpu_div_fState_S3_first__16_BITS_120_TO__ETC___d810 } ;
  assign _theResult___fst_exp__h41468 =
	     (!sfdin__h33169[57] && !sfdin__h33169[56] &&
	      !sfdin__h33169[55] &&
	      !sfdin__h33169[54] &&
	      !sfdin__h33169[53] &&
	      !sfdin__h33169[52] &&
	      !sfdin__h33169[51] &&
	      !sfdin__h33169[50] &&
	      !sfdin__h33169[49] &&
	      !sfdin__h33169[48] &&
	      !sfdin__h33169[47] &&
	      !sfdin__h33169[46] &&
	      !sfdin__h33169[45] &&
	      !sfdin__h33169[44] &&
	      !sfdin__h33169[43] &&
	      !sfdin__h33169[42] &&
	      !sfdin__h33169[41] &&
	      !sfdin__h33169[40] &&
	      !sfdin__h33169[39] &&
	      !sfdin__h33169[38] &&
	      !sfdin__h33169[37] &&
	      !sfdin__h33169[36] &&
	      !sfdin__h33169[35] &&
	      !sfdin__h33169[34] &&
	      !sfdin__h33169[33] &&
	      !sfdin__h33169[32] &&
	      !sfdin__h33169[31] &&
	      !sfdin__h33169[30] &&
	      !sfdin__h33169[29] &&
	      !sfdin__h33169[28] &&
	      !sfdin__h33169[27] &&
	      !sfdin__h33169[26] &&
	      !sfdin__h33169[25] &&
	      !sfdin__h33169[24] &&
	      !sfdin__h33169[23] &&
	      !sfdin__h33169[22] &&
	      !sfdin__h33169[21] &&
	      !sfdin__h33169[20] &&
	      !sfdin__h33169[19] &&
	      !sfdin__h33169[18] &&
	      !sfdin__h33169[17] &&
	      !sfdin__h33169[16] &&
	      !sfdin__h33169[15] &&
	      !sfdin__h33169[14] &&
	      !sfdin__h33169[13] &&
	      !sfdin__h33169[12] &&
	      !sfdin__h33169[11] &&
	      !sfdin__h33169[10] &&
	      !sfdin__h33169[9] &&
	      !sfdin__h33169[8] &&
	      !sfdin__h33169[7] &&
	      !sfdin__h33169[6] &&
	      !sfdin__h33169[5] &&
	      !sfdin__h33169[4] &&
	      !sfdin__h33169[3] &&
	      !sfdin__h33169[2] &&
	      !sfdin__h33169[1] &&
	      !sfdin__h33169[0] ||
	      !_0_CONCAT_IF_IF_fpu_div_fState_S3_first__16_BIT_ETC___d813) ?
	       11'd0 :
	       _theResult___fst_exp__h41462 ;
  assign _theResult___fst_exp__h41471 =
	     (!sfdin__h33169[57] && sfdin__h33169[56]) ?
	       _theResult___fst_exp__h41423 :
	       _theResult___fst_exp__h41468 ;
  assign _theResult___fst_exp__h42607 =
	     (fpu_div_fState_S4$D_OUT[64:54] == 11'd2047) ?
	       fpu_div_fState_S4$D_OUT[64:54] :
	       _theResult___fst_exp__h42604 ;
  assign _theResult___fst_exp__h94750 =
	     fpu_sqr_fState_S3$D_OUT[58] ?
	       _theResult___fst_exp__h94773 :
	       _theResult___fst_exp__h94837 ;
  assign _theResult___fst_exp__h94753 =
	     (fpu_sqr_fState_S3$D_OUT[58] &&
	      IF_fpu_sqr_fState_S3_first__375_BITS_121_TO_11_ETC___d1389 ==
	      12'd1023) ?
	       11'd2046 :
	       _theResult___fst_exp__h94750 ;
  assign _theResult___fst_exp__h94773 =
	     (fpu_sqr_fState_S3$D_OUT[121:111] == 11'd0) ?
	       11'd2 :
	       fpu_sqr_fState_S3$D_OUT[121:111] + 11'd1 ;
  assign _theResult___fst_exp__h94789 =
	     (fpu_sqr_fState_S3$D_OUT[121:111] == 11'd0) ?
	       11'd1 :
	       fpu_sqr_fState_S3$D_OUT[121:111] ;
  assign _theResult___fst_exp__h94828 =
	     fpu_sqr_fState_S3$D_OUT[121:111] -
	     { 5'd0,
	       IF_fpu_sqr_fState_S3_first__375_BIT_58_384_THE_ETC___d1630 } ;
  assign _theResult___fst_exp__h94834 =
	     (!fpu_sqr_fState_S3$D_OUT[58] && !fpu_sqr_fState_S3$D_OUT[57] &&
	      !fpu_sqr_fState_S3$D_OUT[56] &&
	      !fpu_sqr_fState_S3$D_OUT[55] &&
	      !fpu_sqr_fState_S3$D_OUT[54] &&
	      !fpu_sqr_fState_S3$D_OUT[53] &&
	      !fpu_sqr_fState_S3$D_OUT[52] &&
	      !fpu_sqr_fState_S3$D_OUT[51] &&
	      !fpu_sqr_fState_S3$D_OUT[50] &&
	      !fpu_sqr_fState_S3$D_OUT[49] &&
	      !fpu_sqr_fState_S3$D_OUT[48] &&
	      !fpu_sqr_fState_S3$D_OUT[47] &&
	      !fpu_sqr_fState_S3$D_OUT[46] &&
	      !fpu_sqr_fState_S3$D_OUT[45] &&
	      !fpu_sqr_fState_S3$D_OUT[44] &&
	      !fpu_sqr_fState_S3$D_OUT[43] &&
	      !fpu_sqr_fState_S3$D_OUT[42] &&
	      !fpu_sqr_fState_S3$D_OUT[41] &&
	      !fpu_sqr_fState_S3$D_OUT[40] &&
	      !fpu_sqr_fState_S3$D_OUT[39] &&
	      !fpu_sqr_fState_S3$D_OUT[38] &&
	      !fpu_sqr_fState_S3$D_OUT[37] &&
	      !fpu_sqr_fState_S3$D_OUT[36] &&
	      !fpu_sqr_fState_S3$D_OUT[35] &&
	      !fpu_sqr_fState_S3$D_OUT[34] &&
	      !fpu_sqr_fState_S3$D_OUT[33] &&
	      !fpu_sqr_fState_S3$D_OUT[32] &&
	      !fpu_sqr_fState_S3$D_OUT[31] &&
	      !fpu_sqr_fState_S3$D_OUT[30] &&
	      !fpu_sqr_fState_S3$D_OUT[29] &&
	      !fpu_sqr_fState_S3$D_OUT[28] &&
	      !fpu_sqr_fState_S3$D_OUT[27] &&
	      !fpu_sqr_fState_S3$D_OUT[26] &&
	      !fpu_sqr_fState_S3$D_OUT[25] &&
	      !fpu_sqr_fState_S3$D_OUT[24] &&
	      !fpu_sqr_fState_S3$D_OUT[23] &&
	      !fpu_sqr_fState_S3$D_OUT[22] &&
	      !fpu_sqr_fState_S3$D_OUT[21] &&
	      !fpu_sqr_fState_S3$D_OUT[20] &&
	      !fpu_sqr_fState_S3$D_OUT[19] &&
	      !fpu_sqr_fState_S3$D_OUT[18] &&
	      !fpu_sqr_fState_S3$D_OUT[17] &&
	      !fpu_sqr_fState_S3$D_OUT[16] &&
	      !fpu_sqr_fState_S3$D_OUT[15] &&
	      !fpu_sqr_fState_S3$D_OUT[14] &&
	      !fpu_sqr_fState_S3$D_OUT[13] &&
	      !fpu_sqr_fState_S3$D_OUT[12] &&
	      !fpu_sqr_fState_S3$D_OUT[11] &&
	      !fpu_sqr_fState_S3$D_OUT[10] &&
	      !fpu_sqr_fState_S3$D_OUT[9] &&
	      !fpu_sqr_fState_S3$D_OUT[8] &&
	      !fpu_sqr_fState_S3$D_OUT[7] &&
	      !fpu_sqr_fState_S3$D_OUT[6] &&
	      !fpu_sqr_fState_S3$D_OUT[5] &&
	      !fpu_sqr_fState_S3$D_OUT[4] &&
	      !fpu_sqr_fState_S3$D_OUT[3] &&
	      !fpu_sqr_fState_S3$D_OUT[2] &&
	      !fpu_sqr_fState_S3$D_OUT[1] &&
	      !fpu_sqr_fState_S3$D_OUT[0] ||
	      !_0_CONCAT_IF_fpu_sqr_fState_S3_first__375_BIT_5_ETC___d1633) ?
	       11'd0 :
	       _theResult___fst_exp__h94828 ;
  assign _theResult___fst_exp__h94837 =
	     (!fpu_sqr_fState_S3$D_OUT[58] && fpu_sqr_fState_S3$D_OUT[57]) ?
	       _theResult___fst_exp__h94789 :
	       _theResult___fst_exp__h94834 ;
  assign _theResult___fst_exp__h95990 =
	     (fpu_sqr_fState_S4$D_OUT[64:54] == 11'd2047) ?
	       fpu_sqr_fState_S4$D_OUT[64:54] :
	       _theResult___fst_exp__h95987 ;
  assign _theResult___fst_sfd__h164061 =
	     (_theResult___fst_exp__h163334 == 11'd2047) ?
	       _theResult___snd__h163285[56:5] :
	       _theResult___fst_sfd__h164058 ;
  assign _theResult___fst_sfd__h173651 =
	     (_theResult___fst_exp__h172850 == 11'd2047) ?
	       sfdin__h172844[56:5] :
	       _theResult___fst_sfd__h173648 ;
  assign _theResult___fst_sfd__h182403 =
	     (_theResult___fst_exp__h181651 == 11'd2047) ?
	       _theResult___snd__h181597[56:5] :
	       _theResult___fst_sfd__h182400 ;
  assign _theResult___fst_sfd__h182412 =
	     (iFifo$D_OUT[167:160] == 8'd0) ?
	       (_3970_MINUS_0_CONCAT_IF_iFifo_first__087_BIT_15_ETC___d3189 ?
		  _theResult___snd_fst_sfd__h164064 :
		  _theResult___fst_sfd__h148290) :
	       (SEXT_iFifo_first__087_BITS_167_TO_160_130_MINU_ETC___d3324 ?
		  _theResult___snd_fst_sfd__h182406 :
		  _theResult___fst_sfd__h148290) ;
  assign _theResult___fst_sfd__h182418 =
	     ((iFifo$D_OUT[167:160] == 8'd255 ||
	       iFifo$D_OUT[167:160] == 8'd0) &&
	      iFifo$D_OUT[159:137] == 23'd0) ?
	       52'd0 :
	       _theResult___fst_sfd__h182412 ;
  assign _theResult___fst_sfd__h202699 =
	     (_theResult___fst_exp__h201972 == 11'd2047) ?
	       _theResult___snd__h201923[56:5] :
	       _theResult___fst_sfd__h202696 ;
  assign _theResult___fst_sfd__h212289 =
	     (_theResult___fst_exp__h211488 == 11'd2047) ?
	       sfdin__h211482[56:5] :
	       _theResult___fst_sfd__h212286 ;
  assign _theResult___fst_sfd__h221041 =
	     (_theResult___fst_exp__h220289 == 11'd2047) ?
	       _theResult___snd__h220235[56:5] :
	       _theResult___fst_sfd__h221038 ;
  assign _theResult___fst_sfd__h221050 =
	     (iFifo$D_OUT[102:95] == 8'd0) ?
	       (_3970_MINUS_0_CONCAT_IF_iFifo_first__087_BIT_94_ETC___d4684 ?
		  _theResult___snd_fst_sfd__h202702 :
		  _theResult___fst_sfd__h186930) :
	       (SEXT_iFifo_first__087_BITS_102_TO_95_625_MINUS_ETC___d4807 ?
		  _theResult___snd_fst_sfd__h221044 :
		  _theResult___fst_sfd__h186930) ;
  assign _theResult___fst_sfd__h221056 =
	     ((iFifo$D_OUT[102:95] == 8'd255 ||
	       iFifo$D_OUT[102:95] == 8'd0) &&
	      iFifo$D_OUT[94:72] == 23'd0) ?
	       52'd0 :
	       _theResult___fst_sfd__h221050 ;
  assign _theResult___fst_sfd__h241638 =
	     (_theResult___fst_exp__h240911 == 11'd2047) ?
	       _theResult___snd__h240862[56:5] :
	       _theResult___fst_sfd__h241635 ;
  assign _theResult___fst_sfd__h251228 =
	     (_theResult___fst_exp__h250427 == 11'd2047) ?
	       sfdin__h250421[56:5] :
	       _theResult___fst_sfd__h251225 ;
  assign _theResult___fst_sfd__h259980 =
	     (_theResult___fst_exp__h259228 == 11'd2047) ?
	       _theResult___snd__h259174[56:5] :
	       _theResult___fst_sfd__h259977 ;
  assign _theResult___fst_sfd__h259989 =
	     (iFifo$D_OUT[37:30] == 8'd0) ?
	       (_3970_MINUS_0_CONCAT_IF_iFifo_first__087_BIT_29_ETC___d3909 ?
		  _theResult___snd_fst_sfd__h241641 :
		  _theResult___fst_sfd__h225869) :
	       (SEXT_iFifo_first__087_BITS_37_TO_30_850_MINUS__ETC___d4032 ?
		  _theResult___snd_fst_sfd__h259983 :
		  _theResult___fst_sfd__h225869) ;
  assign _theResult___fst_sfd__h259995 =
	     ((iFifo$D_OUT[37:30] == 8'd255 || iFifo$D_OUT[37:30] == 8'd0) &&
	      iFifo$D_OUT[29:7] == 23'd0) ?
	       52'd0 :
	       _theResult___fst_sfd__h259989 ;
  assign _theResult___fst_sfd__h278320 =
	     (_theResult___fst_exp__h277722 == 8'd255) ?
	       sfdin__h277716[56:34] :
	       _theResult___fst_sfd__h278317 ;
  assign _theResult___fst_sfd__h286902 =
	     (_theResult___fst_exp__h286378 == 8'd255) ?
	       _theResult___snd__h286329[56:34] :
	       _theResult___fst_sfd__h286899 ;
  assign _theResult___fst_sfd__h296086 =
	     (_theResult___fst_exp__h295488 == 8'd255) ?
	       sfdin__h295482[56:34] :
	       _theResult___fst_sfd__h296083 ;
  assign _theResult___fst_sfd__h304722 =
	     (_theResult___fst_exp__h304173 == 8'd255) ?
	       _theResult___snd__h304119[56:34] :
	       _theResult___fst_sfd__h304719 ;
  assign _theResult___fst_sfd__h304731 =
	     (resWire$wget[67:57] == 11'd0) ?
	       (_3074_MINUS_0_CONCAT_IF_resWire_wget__410_BIT_5_ETC___d5532 ?
		  _theResult___snd_fst_sfd__h286905 :
		  _theResult___fst_sfd__h269596) :
	       (SEXT_resWire_wget__410_BITS_67_TO_57_416_MINUS_ETC___d6032 ?
		  _theResult___snd_fst_sfd__h304725 :
		  _theResult___fst_sfd__h269596) ;
  assign _theResult___fst_sfd__h304737 =
	     ((resWire$wget[67:57] == 11'd2047 ||
	       resWire$wget[67:57] == 11'd0) &&
	      resWire$wget[56:5] == 52'd0) ?
	       23'd0 :
	       _theResult___fst_sfd__h304731 ;
  assign _theResult___fst_sfd__h42608 =
	     (fpu_div_fState_S4$D_OUT[64:54] == 11'd2047) ?
	       fpu_div_fState_S4$D_OUT[53:2] :
	       _theResult___fst_sfd__h42605 ;
  assign _theResult___fst_sfd__h95991 =
	     (fpu_sqr_fState_S4$D_OUT[64:54] == 11'd2047) ?
	       fpu_sqr_fState_S4$D_OUT[53:2] :
	       _theResult___fst_sfd__h95988 ;
  assign _theResult___fst_sfd__h96608 =
	     fpu_madd_fOperand_S0$D_OUT[195] ?
	       fpu_madd_fOperand_S0$D_OUT[182:131] :
	       52'd0 ;
  assign _theResult___sfd__h142542 =
	     sfd__h142040[53] ?
	       ((fpu_madd_fState_S8$D_OUT[65:55] == 11'd2046) ?
		  52'd0 :
		  sfd__h142040[52:1]) :
	       sfd__h142040[51:0] ;
  assign _theResult___sfd__h163980 =
	     sfd__h163352[53] ?
	       ((_theResult___fst_exp__h163334 == 11'd2046) ?
		  52'd0 :
		  sfd__h163352[52:1]) :
	       sfd__h163352[51:0] ;
  assign _theResult___sfd__h173570 =
	     sfd__h172942[53] ?
	       ((_theResult___fst_exp__h172850 == 11'd2046) ?
		  52'd0 :
		  sfd__h172942[52:1]) :
	       sfd__h172942[51:0] ;
  assign _theResult___sfd__h182322 =
	     sfd__h181670[53] ?
	       ((_theResult___fst_exp__h181651 == 11'd2046) ?
		  52'd0 :
		  sfd__h181670[52:1]) :
	       sfd__h181670[51:0] ;
  assign _theResult___sfd__h202618 =
	     sfd__h201990[53] ?
	       ((_theResult___fst_exp__h201972 == 11'd2046) ?
		  52'd0 :
		  sfd__h201990[52:1]) :
	       sfd__h201990[51:0] ;
  assign _theResult___sfd__h212208 =
	     sfd__h211580[53] ?
	       ((_theResult___fst_exp__h211488 == 11'd2046) ?
		  52'd0 :
		  sfd__h211580[52:1]) :
	       sfd__h211580[51:0] ;
  assign _theResult___sfd__h220960 =
	     sfd__h220308[53] ?
	       ((_theResult___fst_exp__h220289 == 11'd2046) ?
		  52'd0 :
		  sfd__h220308[52:1]) :
	       sfd__h220308[51:0] ;
  assign _theResult___sfd__h241557 =
	     sfd__h240929[53] ?
	       ((_theResult___fst_exp__h240911 == 11'd2046) ?
		  52'd0 :
		  sfd__h240929[52:1]) :
	       sfd__h240929[51:0] ;
  assign _theResult___sfd__h251147 =
	     sfd__h250519[53] ?
	       ((_theResult___fst_exp__h250427 == 11'd2046) ?
		  52'd0 :
		  sfd__h250519[52:1]) :
	       sfd__h250519[51:0] ;
  assign _theResult___sfd__h259899 =
	     sfd__h259247[53] ?
	       ((_theResult___fst_exp__h259228 == 11'd2046) ?
		  52'd0 :
		  sfd__h259247[52:1]) :
	       sfd__h259247[51:0] ;
  assign _theResult___sfd__h278239 =
	     sfd__h277814[24] ?
	       ((_theResult___fst_exp__h277722 == 8'd254) ?
		  23'd0 :
		  sfd__h277814[23:1]) :
	       sfd__h277814[22:0] ;
  assign _theResult___sfd__h286821 =
	     sfd__h286396[24] ?
	       ((_theResult___fst_exp__h286378 == 8'd254) ?
		  23'd0 :
		  sfd__h286396[23:1]) :
	       sfd__h286396[22:0] ;
  assign _theResult___sfd__h296005 =
	     sfd__h295580[24] ?
	       ((_theResult___fst_exp__h295488 == 8'd254) ?
		  23'd0 :
		  sfd__h295580[23:1]) :
	       sfd__h295580[22:0] ;
  assign _theResult___sfd__h304641 =
	     sfd__h304192[24] ?
	       ((_theResult___fst_exp__h304173 == 8'd254) ?
		  23'd0 :
		  sfd__h304192[23:1]) :
	       sfd__h304192[22:0] ;
  assign _theResult___sfd__h42527 =
	     sfd__h42033[53] ?
	       ((fpu_div_fState_S4$D_OUT[64:54] == 11'd2046) ?
		  52'd0 :
		  sfd__h42033[52:1]) :
	       sfd__h42033[51:0] ;
  assign _theResult___sfd__h95910 =
	     sfd__h95416[53] ?
	       ((fpu_sqr_fState_S4$D_OUT[64:54] == 11'd2046) ?
		  52'd0 :
		  sfd__h95416[52:1]) :
	       sfd__h95416[51:0] ;
  assign _theResult___snd__h130966 = { sfdBC__h115662[104:0], 1'd0 } ;
  assign _theResult___snd__h130980 =
	     (!sfdBC__h115662[105] && sfdBC__h115662[104]) ?
	       _theResult___snd__h130982 :
	       _theResult___snd__h130994 ;
  assign _theResult___snd__h130982 = { sfdBC__h115662[103:0], 2'd0 } ;
  assign _theResult___snd__h130994 =
	     (!sfdBC__h115662[105] && !sfdBC__h115662[104] &&
	      !sfdBC__h115662[103] &&
	      !sfdBC__h115662[102] &&
	      !sfdBC__h115662[101] &&
	      !sfdBC__h115662[100] &&
	      !sfdBC__h115662[99] &&
	      !sfdBC__h115662[98] &&
	      !sfdBC__h115662[97] &&
	      !sfdBC__h115662[96] &&
	      !sfdBC__h115662[95] &&
	      !sfdBC__h115662[94] &&
	      !sfdBC__h115662[93] &&
	      !sfdBC__h115662[92] &&
	      !sfdBC__h115662[91] &&
	      !sfdBC__h115662[90] &&
	      !sfdBC__h115662[89] &&
	      !sfdBC__h115662[88] &&
	      !sfdBC__h115662[87] &&
	      !sfdBC__h115662[86] &&
	      !sfdBC__h115662[85] &&
	      !sfdBC__h115662[84] &&
	      !sfdBC__h115662[83] &&
	      !sfdBC__h115662[82] &&
	      !sfdBC__h115662[81] &&
	      !sfdBC__h115662[80] &&
	      !sfdBC__h115662[79] &&
	      !sfdBC__h115662[78] &&
	      !sfdBC__h115662[77] &&
	      !sfdBC__h115662[76] &&
	      !sfdBC__h115662[75] &&
	      !sfdBC__h115662[74] &&
	      !sfdBC__h115662[73] &&
	      !sfdBC__h115662[72] &&
	      !sfdBC__h115662[71] &&
	      !sfdBC__h115662[70] &&
	      !sfdBC__h115662[69] &&
	      !sfdBC__h115662[68] &&
	      !sfdBC__h115662[67] &&
	      !sfdBC__h115662[66] &&
	      !sfdBC__h115662[65] &&
	      !sfdBC__h115662[64] &&
	      !sfdBC__h115662[63] &&
	      !sfdBC__h115662[62] &&
	      !sfdBC__h115662[61] &&
	      !sfdBC__h115662[60] &&
	      !sfdBC__h115662[59] &&
	      !sfdBC__h115662[58] &&
	      !sfdBC__h115662[57] &&
	      !sfdBC__h115662[56] &&
	      !sfdBC__h115662[55] &&
	      !sfdBC__h115662[54] &&
	      !sfdBC__h115662[53] &&
	      !sfdBC__h115662[52] &&
	      !sfdBC__h115662[51] &&
	      !sfdBC__h115662[50] &&
	      !sfdBC__h115662[49] &&
	      !sfdBC__h115662[48] &&
	      !sfdBC__h115662[47] &&
	      !sfdBC__h115662[46] &&
	      !sfdBC__h115662[45] &&
	      !sfdBC__h115662[44] &&
	      !sfdBC__h115662[43] &&
	      !sfdBC__h115662[42] &&
	      !sfdBC__h115662[41] &&
	      !sfdBC__h115662[40] &&
	      !sfdBC__h115662[39] &&
	      !sfdBC__h115662[38] &&
	      !sfdBC__h115662[37] &&
	      !sfdBC__h115662[36] &&
	      !sfdBC__h115662[35] &&
	      !sfdBC__h115662[34] &&
	      !sfdBC__h115662[33] &&
	      !sfdBC__h115662[32] &&
	      !sfdBC__h115662[31] &&
	      !sfdBC__h115662[30] &&
	      !sfdBC__h115662[29] &&
	      !sfdBC__h115662[28] &&
	      !sfdBC__h115662[27] &&
	      !sfdBC__h115662[26] &&
	      !sfdBC__h115662[25] &&
	      !sfdBC__h115662[24] &&
	      !sfdBC__h115662[23] &&
	      !sfdBC__h115662[22] &&
	      !sfdBC__h115662[21] &&
	      !sfdBC__h115662[20] &&
	      !sfdBC__h115662[19] &&
	      !sfdBC__h115662[18] &&
	      !sfdBC__h115662[17] &&
	      !sfdBC__h115662[16] &&
	      !sfdBC__h115662[15] &&
	      !sfdBC__h115662[14] &&
	      !sfdBC__h115662[13] &&
	      !sfdBC__h115662[12] &&
	      !sfdBC__h115662[11] &&
	      !sfdBC__h115662[10] &&
	      !sfdBC__h115662[9] &&
	      !sfdBC__h115662[8] &&
	      !sfdBC__h115662[7] &&
	      !sfdBC__h115662[6] &&
	      !sfdBC__h115662[5] &&
	      !sfdBC__h115662[4] &&
	      !sfdBC__h115662[3] &&
	      !sfdBC__h115662[2] &&
	      !sfdBC__h115662[1] &&
	      !sfdBC__h115662[0]) ?
	       sfdBC__h115662 :
	       _theResult___snd__h131000 ;
  assign _theResult___snd__h131000 =
	     { IF_0_CONCAT_IF_IF_7170_MINUS_fpu_madd_fState_S_ETC__q24[103:0],
	       2'd0 } ;
  assign _theResult___snd__h131018 =
	     sfdBC__h115662 <<
	     IF_IF_7170_MINUS_fpu_madd_fState_S3_first__995_ETC___d2462 ;
  assign _theResult___snd__h131023 =
	     sfdBC__h115662 <<
	     IF_IF_7170_MINUS_fpu_madd_fState_S3_first__995_ETC___d2460 ;
  assign _theResult___snd__h141392 = { sfd__h133119[55:0], 1'd0 } ;
  assign _theResult___snd__h141406 =
	     (!sfd__h133119[56] && sfd__h133119[55]) ?
	       _theResult___snd__h141408 :
	       _theResult___snd__h141420 ;
  assign _theResult___snd__h141408 = { sfd__h133119[54:0], 2'd0 } ;
  assign _theResult___snd__h141420 =
	     (!sfd__h133119[56] && !sfd__h133119[55] && !sfd__h133119[54] &&
	      !sfd__h133119[53] &&
	      !sfd__h133119[52] &&
	      !sfd__h133119[51] &&
	      !sfd__h133119[50] &&
	      !sfd__h133119[49] &&
	      !sfd__h133119[48] &&
	      !sfd__h133119[47] &&
	      !sfd__h133119[46] &&
	      !sfd__h133119[45] &&
	      !sfd__h133119[44] &&
	      !sfd__h133119[43] &&
	      !sfd__h133119[42] &&
	      !sfd__h133119[41] &&
	      !sfd__h133119[40] &&
	      !sfd__h133119[39] &&
	      !sfd__h133119[38] &&
	      !sfd__h133119[37] &&
	      !sfd__h133119[36] &&
	      !sfd__h133119[35] &&
	      !sfd__h133119[34] &&
	      !sfd__h133119[33] &&
	      !sfd__h133119[32] &&
	      !sfd__h133119[31] &&
	      !sfd__h133119[30] &&
	      !sfd__h133119[29] &&
	      !sfd__h133119[28] &&
	      !sfd__h133119[27] &&
	      !sfd__h133119[26] &&
	      !sfd__h133119[25] &&
	      !sfd__h133119[24] &&
	      !sfd__h133119[23] &&
	      !sfd__h133119[22] &&
	      !sfd__h133119[21] &&
	      !sfd__h133119[20] &&
	      !sfd__h133119[19] &&
	      !sfd__h133119[18] &&
	      !sfd__h133119[17] &&
	      !sfd__h133119[16] &&
	      !sfd__h133119[15] &&
	      !sfd__h133119[14] &&
	      !sfd__h133119[13] &&
	      !sfd__h133119[12] &&
	      !sfd__h133119[11] &&
	      !sfd__h133119[10] &&
	      !sfd__h133119[9] &&
	      !sfd__h133119[8] &&
	      !sfd__h133119[7] &&
	      !sfd__h133119[6] &&
	      !sfd__h133119[5] &&
	      !sfd__h133119[4] &&
	      !sfd__h133119[3] &&
	      !sfd__h133119[2] &&
	      !sfd__h133119[1] &&
	      !sfd__h133119[0]) ?
	       sfd__h133119 :
	       _theResult___snd__h141426 ;
  assign _theResult___snd__h141426 =
	     { IF_0_CONCAT_IF_IF_fpu_madd_fState_S7_first__65_ETC__q29[54:0],
	       2'd0 } ;
  assign _theResult___snd__h141444 =
	     sfd__h133119 <<
	     IF_fpu_madd_fState_S7_first__651_BITS_126_TO_1_ETC___d2903 ;
  assign _theResult___snd__h141449 =
	     sfd__h133119 <<
	     IF_IF_fpu_madd_fState_S7_first__651_BIT_128_65_ETC___d2901 ;
  assign _theResult___snd__h163285 =
	     (iFifo$D_OUT[167:160] == 8'd0) ?
	       _theResult___snd__h163294 :
	       _theResult___snd__h163287 ;
  assign _theResult___snd__h163287 = { iFifo$D_OUT[159:137], 34'd0 } ;
  assign _theResult___snd__h163294 =
	     (iFifo$D_OUT[167:160] == 8'd0 && !iFifo$D_OUT[159] &&
	      NOT_iFifo_first__087_BIT_158_142_202_AND_NOT_i_ETC___d3244) ?
	       sfd__h144534 :
	       _theResult___snd__h163300 ;
  assign _theResult___snd__h163300 =
	     { IF_0_CONCAT_IF_iFifo_first__087_BITS_167_TO_16_ETC__q33[54:0],
	       2'd0 } ;
  assign _theResult___snd__h163323 =
	     sfd__h144534 <<
	     IF_iFifo_first__087_BITS_167_TO_160_130_EQ_0_1_ETC___d3271 ;
  assign _theResult___snd__h172861 = { _theResult____h164612[55:0], 1'd0 } ;
  assign _theResult___snd__h172872 =
	     (!_theResult____h164612[56] && _theResult____h164612[55]) ?
	       _theResult___snd__h172874 :
	       _theResult___snd__h172884 ;
  assign _theResult___snd__h172874 = { _theResult____h164612[54:0], 2'd0 } ;
  assign _theResult___snd__h172884 =
	     (!_theResult____h164612[56] && !_theResult____h164612[55] &&
	      !_theResult____h164612[54] &&
	      !_theResult____h164612[53] &&
	      !_theResult____h164612[52] &&
	      !_theResult____h164612[51] &&
	      !_theResult____h164612[50] &&
	      !_theResult____h164612[49] &&
	      !_theResult____h164612[48] &&
	      !_theResult____h164612[47] &&
	      !_theResult____h164612[46] &&
	      !_theResult____h164612[45] &&
	      !_theResult____h164612[44] &&
	      !_theResult____h164612[43] &&
	      !_theResult____h164612[42] &&
	      !_theResult____h164612[41] &&
	      !_theResult____h164612[40] &&
	      !_theResult____h164612[39] &&
	      !_theResult____h164612[38] &&
	      !_theResult____h164612[37] &&
	      !_theResult____h164612[36] &&
	      !_theResult____h164612[35] &&
	      !_theResult____h164612[34] &&
	      !_theResult____h164612[33] &&
	      !_theResult____h164612[32] &&
	      !_theResult____h164612[31] &&
	      !_theResult____h164612[30] &&
	      !_theResult____h164612[29] &&
	      !_theResult____h164612[28] &&
	      !_theResult____h164612[27] &&
	      !_theResult____h164612[26] &&
	      !_theResult____h164612[25] &&
	      !_theResult____h164612[24] &&
	      !_theResult____h164612[23] &&
	      !_theResult____h164612[22] &&
	      !_theResult____h164612[21] &&
	      !_theResult____h164612[20] &&
	      !_theResult____h164612[19] &&
	      !_theResult____h164612[18] &&
	      !_theResult____h164612[17] &&
	      !_theResult____h164612[16] &&
	      !_theResult____h164612[15] &&
	      !_theResult____h164612[14] &&
	      !_theResult____h164612[13] &&
	      !_theResult____h164612[12] &&
	      !_theResult____h164612[11] &&
	      !_theResult____h164612[10] &&
	      !_theResult____h164612[9] &&
	      !_theResult____h164612[8] &&
	      !_theResult____h164612[7] &&
	      !_theResult____h164612[6] &&
	      !_theResult____h164612[5] &&
	      !_theResult____h164612[4] &&
	      !_theResult____h164612[3] &&
	      !_theResult____h164612[2] &&
	      !_theResult____h164612[1] &&
	      !_theResult____h164612[0]) ?
	       _theResult____h164612 :
	       _theResult___snd__h172890 ;
  assign _theResult___snd__h172890 =
	     { IF_0_CONCAT_IF_IF_3074_MINUS_SEXT_iFifo_first__ETC__q37[54:0],
	       2'd0 } ;
  assign _theResult___snd__h172913 =
	     _theResult____h164612 <<
	     IF_IF_3074_MINUS_SEXT_iFifo_first__087_BITS_16_ETC___d3572 ;
  assign _theResult___snd__h181597 =
	     (iFifo$D_OUT[167:160] == 8'd0) ?
	       _theResult___snd__h181611 :
	       _theResult___snd__h163287 ;
  assign _theResult___snd__h181611 =
	     (iFifo$D_OUT[167:160] == 8'd0 && !iFifo$D_OUT[159] &&
	      NOT_iFifo_first__087_BIT_158_142_202_AND_NOT_i_ETC___d3244) ?
	       sfd__h144534 :
	       _theResult___snd__h181617 ;
  assign _theResult___snd__h181617 =
	     { IF_0_CONCAT_IF_iFifo_first__087_BITS_167_TO_16_ETC__q40[54:0],
	       2'd0 } ;
  assign _theResult___snd__h181635 =
	     sfd__h144534 <<
	     IF_SEXT_iFifo_first__087_BITS_167_TO_160_130_M_ETC___d3623 ;
  assign _theResult___snd__h201923 =
	     (iFifo$D_OUT[102:95] == 8'd0) ?
	       _theResult___snd__h201932 :
	       _theResult___snd__h201925 ;
  assign _theResult___snd__h201925 = { iFifo$D_OUT[94:72], 34'd0 } ;
  assign _theResult___snd__h201932 =
	     (iFifo$D_OUT[102:95] == 8'd0 && !iFifo$D_OUT[94] &&
	      NOT_iFifo_first__087_BIT_93_637_688_AND_NOT_iF_ETC___d4730) ?
	       sfd__h183174 :
	       _theResult___snd__h201938 ;
  assign _theResult___snd__h201938 =
	     { IF_0_CONCAT_IF_iFifo_first__087_BITS_102_TO_95_ETC__q93[54:0],
	       2'd0 } ;
  assign _theResult___snd__h201961 =
	     sfd__h183174 <<
	     IF_iFifo_first__087_BITS_102_TO_95_625_EQ_0_63_ETC___d4757 ;
  assign _theResult___snd__h211499 = { _theResult____h203250[55:0], 1'd0 } ;
  assign _theResult___snd__h211510 =
	     (!_theResult____h203250[56] && _theResult____h203250[55]) ?
	       _theResult___snd__h211512 :
	       _theResult___snd__h211522 ;
  assign _theResult___snd__h211512 = { _theResult____h203250[54:0], 2'd0 } ;
  assign _theResult___snd__h211522 =
	     (!_theResult____h203250[56] && !_theResult____h203250[55] &&
	      !_theResult____h203250[54] &&
	      !_theResult____h203250[53] &&
	      !_theResult____h203250[52] &&
	      !_theResult____h203250[51] &&
	      !_theResult____h203250[50] &&
	      !_theResult____h203250[49] &&
	      !_theResult____h203250[48] &&
	      !_theResult____h203250[47] &&
	      !_theResult____h203250[46] &&
	      !_theResult____h203250[45] &&
	      !_theResult____h203250[44] &&
	      !_theResult____h203250[43] &&
	      !_theResult____h203250[42] &&
	      !_theResult____h203250[41] &&
	      !_theResult____h203250[40] &&
	      !_theResult____h203250[39] &&
	      !_theResult____h203250[38] &&
	      !_theResult____h203250[37] &&
	      !_theResult____h203250[36] &&
	      !_theResult____h203250[35] &&
	      !_theResult____h203250[34] &&
	      !_theResult____h203250[33] &&
	      !_theResult____h203250[32] &&
	      !_theResult____h203250[31] &&
	      !_theResult____h203250[30] &&
	      !_theResult____h203250[29] &&
	      !_theResult____h203250[28] &&
	      !_theResult____h203250[27] &&
	      !_theResult____h203250[26] &&
	      !_theResult____h203250[25] &&
	      !_theResult____h203250[24] &&
	      !_theResult____h203250[23] &&
	      !_theResult____h203250[22] &&
	      !_theResult____h203250[21] &&
	      !_theResult____h203250[20] &&
	      !_theResult____h203250[19] &&
	      !_theResult____h203250[18] &&
	      !_theResult____h203250[17] &&
	      !_theResult____h203250[16] &&
	      !_theResult____h203250[15] &&
	      !_theResult____h203250[14] &&
	      !_theResult____h203250[13] &&
	      !_theResult____h203250[12] &&
	      !_theResult____h203250[11] &&
	      !_theResult____h203250[10] &&
	      !_theResult____h203250[9] &&
	      !_theResult____h203250[8] &&
	      !_theResult____h203250[7] &&
	      !_theResult____h203250[6] &&
	      !_theResult____h203250[5] &&
	      !_theResult____h203250[4] &&
	      !_theResult____h203250[3] &&
	      !_theResult____h203250[2] &&
	      !_theResult____h203250[1] &&
	      !_theResult____h203250[0]) ?
	       _theResult____h203250 :
	       _theResult___snd__h211528 ;
  assign _theResult___snd__h211528 =
	     { IF_0_CONCAT_IF_IF_3074_MINUS_SEXT_iFifo_first__ETC__q97[54:0],
	       2'd0 } ;
  assign _theResult___snd__h211551 =
	     _theResult____h203250 <<
	     IF_IF_3074_MINUS_SEXT_iFifo_first__087_BITS_10_ETC___d5055 ;
  assign _theResult___snd__h220235 =
	     (iFifo$D_OUT[102:95] == 8'd0) ?
	       _theResult___snd__h220249 :
	       _theResult___snd__h201925 ;
  assign _theResult___snd__h220249 =
	     (iFifo$D_OUT[102:95] == 8'd0 && !iFifo$D_OUT[94] &&
	      NOT_iFifo_first__087_BIT_93_637_688_AND_NOT_iF_ETC___d4730) ?
	       sfd__h183174 :
	       _theResult___snd__h220255 ;
  assign _theResult___snd__h220255 =
	     { IF_0_CONCAT_IF_iFifo_first__087_BITS_102_TO_95_ETC__q100[54:0],
	       2'd0 } ;
  assign _theResult___snd__h220273 =
	     sfd__h183174 <<
	     IF_SEXT_iFifo_first__087_BITS_102_TO_95_625_MI_ETC___d5106 ;
  assign _theResult___snd__h240862 =
	     (iFifo$D_OUT[37:30] == 8'd0) ?
	       _theResult___snd__h240871 :
	       _theResult___snd__h240864 ;
  assign _theResult___snd__h240864 = { iFifo$D_OUT[29:7], 34'd0 } ;
  assign _theResult___snd__h240871 =
	     (iFifo$D_OUT[37:30] == 8'd0 && !iFifo$D_OUT[29] &&
	      NOT_iFifo_first__087_BIT_28_862_913_AND_NOT_iF_ETC___d3955) ?
	       sfd__h222113 :
	       _theResult___snd__h240877 ;
  assign _theResult___snd__h240877 =
	     { IF_0_CONCAT_IF_iFifo_first__087_BITS_37_TO_30__ETC__q60[54:0],
	       2'd0 } ;
  assign _theResult___snd__h240900 =
	     sfd__h222113 <<
	     IF_iFifo_first__087_BITS_37_TO_30_850_EQ_0_856_ETC___d3982 ;
  assign _theResult___snd__h250438 = { _theResult____h242189[55:0], 1'd0 } ;
  assign _theResult___snd__h250449 =
	     (!_theResult____h242189[56] && _theResult____h242189[55]) ?
	       _theResult___snd__h250451 :
	       _theResult___snd__h250461 ;
  assign _theResult___snd__h250451 = { _theResult____h242189[54:0], 2'd0 } ;
  assign _theResult___snd__h250461 =
	     (!_theResult____h242189[56] && !_theResult____h242189[55] &&
	      !_theResult____h242189[54] &&
	      !_theResult____h242189[53] &&
	      !_theResult____h242189[52] &&
	      !_theResult____h242189[51] &&
	      !_theResult____h242189[50] &&
	      !_theResult____h242189[49] &&
	      !_theResult____h242189[48] &&
	      !_theResult____h242189[47] &&
	      !_theResult____h242189[46] &&
	      !_theResult____h242189[45] &&
	      !_theResult____h242189[44] &&
	      !_theResult____h242189[43] &&
	      !_theResult____h242189[42] &&
	      !_theResult____h242189[41] &&
	      !_theResult____h242189[40] &&
	      !_theResult____h242189[39] &&
	      !_theResult____h242189[38] &&
	      !_theResult____h242189[37] &&
	      !_theResult____h242189[36] &&
	      !_theResult____h242189[35] &&
	      !_theResult____h242189[34] &&
	      !_theResult____h242189[33] &&
	      !_theResult____h242189[32] &&
	      !_theResult____h242189[31] &&
	      !_theResult____h242189[30] &&
	      !_theResult____h242189[29] &&
	      !_theResult____h242189[28] &&
	      !_theResult____h242189[27] &&
	      !_theResult____h242189[26] &&
	      !_theResult____h242189[25] &&
	      !_theResult____h242189[24] &&
	      !_theResult____h242189[23] &&
	      !_theResult____h242189[22] &&
	      !_theResult____h242189[21] &&
	      !_theResult____h242189[20] &&
	      !_theResult____h242189[19] &&
	      !_theResult____h242189[18] &&
	      !_theResult____h242189[17] &&
	      !_theResult____h242189[16] &&
	      !_theResult____h242189[15] &&
	      !_theResult____h242189[14] &&
	      !_theResult____h242189[13] &&
	      !_theResult____h242189[12] &&
	      !_theResult____h242189[11] &&
	      !_theResult____h242189[10] &&
	      !_theResult____h242189[9] &&
	      !_theResult____h242189[8] &&
	      !_theResult____h242189[7] &&
	      !_theResult____h242189[6] &&
	      !_theResult____h242189[5] &&
	      !_theResult____h242189[4] &&
	      !_theResult____h242189[3] &&
	      !_theResult____h242189[2] &&
	      !_theResult____h242189[1] &&
	      !_theResult____h242189[0]) ?
	       _theResult____h242189 :
	       _theResult___snd__h250467 ;
  assign _theResult___snd__h250467 =
	     { IF_0_CONCAT_IF_IF_3074_MINUS_SEXT_iFifo_first__ETC__q64[54:0],
	       2'd0 } ;
  assign _theResult___snd__h250490 =
	     _theResult____h242189 <<
	     IF_IF_3074_MINUS_SEXT_iFifo_first__087_BITS_37_ETC___d4280 ;
  assign _theResult___snd__h259174 =
	     (iFifo$D_OUT[37:30] == 8'd0) ?
	       _theResult___snd__h259188 :
	       _theResult___snd__h240864 ;
  assign _theResult___snd__h259188 =
	     (iFifo$D_OUT[37:30] == 8'd0 && !iFifo$D_OUT[29] &&
	      NOT_iFifo_first__087_BIT_28_862_913_AND_NOT_iF_ETC___d3955) ?
	       sfd__h222113 :
	       _theResult___snd__h259194 ;
  assign _theResult___snd__h259194 =
	     { IF_0_CONCAT_IF_iFifo_first__087_BITS_37_TO_30__ETC__q67[54:0],
	       2'd0 } ;
  assign _theResult___snd__h259212 =
	     sfd__h222113 <<
	     IF_SEXT_iFifo_first__087_BITS_37_TO_30_850_MIN_ETC___d4331 ;
  assign _theResult___snd__h277733 = { _theResult____h269613[55:0], 1'd0 } ;
  assign _theResult___snd__h277744 =
	     (!_theResult____h269613[56] && _theResult____h269613[55]) ?
	       _theResult___snd__h277746 :
	       _theResult___snd__h277756 ;
  assign _theResult___snd__h277746 = { _theResult____h269613[54:0], 2'd0 } ;
  assign _theResult___snd__h277756 =
	     (!_theResult____h269613[56] && !_theResult____h269613[55] &&
	      !_theResult____h269613[54] &&
	      !_theResult____h269613[53] &&
	      !_theResult____h269613[52] &&
	      !_theResult____h269613[51] &&
	      !_theResult____h269613[50] &&
	      !_theResult____h269613[49] &&
	      !_theResult____h269613[48] &&
	      !_theResult____h269613[47] &&
	      !_theResult____h269613[46] &&
	      !_theResult____h269613[45] &&
	      !_theResult____h269613[44] &&
	      !_theResult____h269613[43] &&
	      !_theResult____h269613[42] &&
	      !_theResult____h269613[41] &&
	      !_theResult____h269613[40] &&
	      !_theResult____h269613[39] &&
	      !_theResult____h269613[38] &&
	      !_theResult____h269613[37] &&
	      !_theResult____h269613[36] &&
	      !_theResult____h269613[35] &&
	      !_theResult____h269613[34] &&
	      !_theResult____h269613[33] &&
	      !_theResult____h269613[32] &&
	      !_theResult____h269613[31] &&
	      !_theResult____h269613[30] &&
	      !_theResult____h269613[29] &&
	      !_theResult____h269613[28] &&
	      !_theResult____h269613[27] &&
	      !_theResult____h269613[26] &&
	      !_theResult____h269613[25] &&
	      !_theResult____h269613[24] &&
	      !_theResult____h269613[23] &&
	      !_theResult____h269613[22] &&
	      !_theResult____h269613[21] &&
	      !_theResult____h269613[20] &&
	      !_theResult____h269613[19] &&
	      !_theResult____h269613[18] &&
	      !_theResult____h269613[17] &&
	      !_theResult____h269613[16] &&
	      !_theResult____h269613[15] &&
	      !_theResult____h269613[14] &&
	      !_theResult____h269613[13] &&
	      !_theResult____h269613[12] &&
	      !_theResult____h269613[11] &&
	      !_theResult____h269613[10] &&
	      !_theResult____h269613[9] &&
	      !_theResult____h269613[8] &&
	      !_theResult____h269613[7] &&
	      !_theResult____h269613[6] &&
	      !_theResult____h269613[5] &&
	      !_theResult____h269613[4] &&
	      !_theResult____h269613[3] &&
	      !_theResult____h269613[2] &&
	      !_theResult____h269613[1] &&
	      !_theResult____h269613[0]) ?
	       _theResult____h269613 :
	       _theResult___snd__h277762 ;
  assign _theResult___snd__h277762 =
	     { IF_0_CONCAT_IF_IF_0b0_CONCAT_NOT_resWire_wget__ETC__q133[54:0],
	       2'd0 } ;
  assign _theResult___snd__h277785 =
	     _theResult____h269613 <<
	     IF_IF_0b0_CONCAT_NOT_resWire_wget__410_BITS_67_ETC___d5767 ;
  assign _theResult___snd__h286329 =
	     (resWire$wget[67:57] == 11'd0) ?
	       _theResult___snd__h286338 :
	       _theResult___snd__h286331 ;
  assign _theResult___snd__h286331 = { resWire$wget[56:5], 5'd0 } ;
  assign _theResult___snd__h286338 =
	     (resWire$wget[67:57] == 11'd0 &&
	      NOT_resWire_wget__410_BIT_56_426_825_AND_NOT_r_ETC___d5927) ?
	       sfd__h262011 :
	       _theResult___snd__h286344 ;
  assign _theResult___snd__h286344 =
	     { IF_0_CONCAT_IF_resWire_wget__410_BITS_67_TO_57_ETC__q135[54:0],
	       2'd0 } ;
  assign _theResult___snd__h286367 =
	     sfd__h262011 <<
	     IF_resWire_wget__410_BITS_67_TO_57_416_EQ_0_42_ETC___d5982 ;
  assign _theResult___snd__h295499 = { _theResult____h287250[55:0], 1'd0 } ;
  assign _theResult___snd__h295510 =
	     (!_theResult____h287250[56] && _theResult____h287250[55]) ?
	       _theResult___snd__h295512 :
	       _theResult___snd__h295522 ;
  assign _theResult___snd__h295512 = { _theResult____h287250[54:0], 2'd0 } ;
  assign _theResult___snd__h295522 =
	     (!_theResult____h287250[56] && !_theResult____h287250[55] &&
	      !_theResult____h287250[54] &&
	      !_theResult____h287250[53] &&
	      !_theResult____h287250[52] &&
	      !_theResult____h287250[51] &&
	      !_theResult____h287250[50] &&
	      !_theResult____h287250[49] &&
	      !_theResult____h287250[48] &&
	      !_theResult____h287250[47] &&
	      !_theResult____h287250[46] &&
	      !_theResult____h287250[45] &&
	      !_theResult____h287250[44] &&
	      !_theResult____h287250[43] &&
	      !_theResult____h287250[42] &&
	      !_theResult____h287250[41] &&
	      !_theResult____h287250[40] &&
	      !_theResult____h287250[39] &&
	      !_theResult____h287250[38] &&
	      !_theResult____h287250[37] &&
	      !_theResult____h287250[36] &&
	      !_theResult____h287250[35] &&
	      !_theResult____h287250[34] &&
	      !_theResult____h287250[33] &&
	      !_theResult____h287250[32] &&
	      !_theResult____h287250[31] &&
	      !_theResult____h287250[30] &&
	      !_theResult____h287250[29] &&
	      !_theResult____h287250[28] &&
	      !_theResult____h287250[27] &&
	      !_theResult____h287250[26] &&
	      !_theResult____h287250[25] &&
	      !_theResult____h287250[24] &&
	      !_theResult____h287250[23] &&
	      !_theResult____h287250[22] &&
	      !_theResult____h287250[21] &&
	      !_theResult____h287250[20] &&
	      !_theResult____h287250[19] &&
	      !_theResult____h287250[18] &&
	      !_theResult____h287250[17] &&
	      !_theResult____h287250[16] &&
	      !_theResult____h287250[15] &&
	      !_theResult____h287250[14] &&
	      !_theResult____h287250[13] &&
	      !_theResult____h287250[12] &&
	      !_theResult____h287250[11] &&
	      !_theResult____h287250[10] &&
	      !_theResult____h287250[9] &&
	      !_theResult____h287250[8] &&
	      !_theResult____h287250[7] &&
	      !_theResult____h287250[6] &&
	      !_theResult____h287250[5] &&
	      !_theResult____h287250[4] &&
	      !_theResult____h287250[3] &&
	      !_theResult____h287250[2] &&
	      !_theResult____h287250[1] &&
	      !_theResult____h287250[0]) ?
	       _theResult____h287250 :
	       _theResult___snd__h295528 ;
  assign _theResult___snd__h295528 =
	     { IF_0_CONCAT_IF_IF_3970_MINUS_SEXT_resWire_wget_ETC__q139[54:0],
	       2'd0 } ;
  assign _theResult___snd__h295551 =
	     _theResult____h287250 <<
	     IF_IF_3970_MINUS_SEXT_resWire_wget__410_BITS_6_ETC___d6278 ;
  assign _theResult___snd__h304119 =
	     (resWire$wget[67:57] == 11'd0) ?
	       _theResult___snd__h304133 :
	       _theResult___snd__h286331 ;
  assign _theResult___snd__h304133 =
	     (resWire$wget[67:57] == 11'd0 &&
	      NOT_resWire_wget__410_BIT_56_426_825_AND_NOT_r_ETC___d5927) ?
	       sfd__h262011 :
	       _theResult___snd__h304139 ;
  assign _theResult___snd__h304139 =
	     { IF_0_CONCAT_IF_resWire_wget__410_BITS_67_TO_57_ETC__q142[54:0],
	       2'd0 } ;
  assign _theResult___snd__h304157 =
	     sfd__h262011 <<
	     IF_SEXT_resWire_wget__410_BITS_67_TO_57_416_MI_ETC___d6332 ;
  assign _theResult___snd__h33766 = { fpu_div_fState_S3$D_OUT[56:0], 1'd0 } ;
  assign _theResult___snd__h41401 = { sfdin__h33169[56:0], 1'd0 } ;
  assign _theResult___snd__h41416 =
	     (!sfdin__h33169[57] && sfdin__h33169[56]) ?
	       _theResult___snd__h41418 :
	       _theResult___snd__h41431 ;
  assign _theResult___snd__h41418 = { sfdin__h33169[55:0], 2'd0 } ;
  assign _theResult___snd__h41431 =
	     (!sfdin__h33169[57] && !sfdin__h33169[56] &&
	      !sfdin__h33169[55] &&
	      !sfdin__h33169[54] &&
	      !sfdin__h33169[53] &&
	      !sfdin__h33169[52] &&
	      !sfdin__h33169[51] &&
	      !sfdin__h33169[50] &&
	      !sfdin__h33169[49] &&
	      !sfdin__h33169[48] &&
	      !sfdin__h33169[47] &&
	      !sfdin__h33169[46] &&
	      !sfdin__h33169[45] &&
	      !sfdin__h33169[44] &&
	      !sfdin__h33169[43] &&
	      !sfdin__h33169[42] &&
	      !sfdin__h33169[41] &&
	      !sfdin__h33169[40] &&
	      !sfdin__h33169[39] &&
	      !sfdin__h33169[38] &&
	      !sfdin__h33169[37] &&
	      !sfdin__h33169[36] &&
	      !sfdin__h33169[35] &&
	      !sfdin__h33169[34] &&
	      !sfdin__h33169[33] &&
	      !sfdin__h33169[32] &&
	      !sfdin__h33169[31] &&
	      !sfdin__h33169[30] &&
	      !sfdin__h33169[29] &&
	      !sfdin__h33169[28] &&
	      !sfdin__h33169[27] &&
	      !sfdin__h33169[26] &&
	      !sfdin__h33169[25] &&
	      !sfdin__h33169[24] &&
	      !sfdin__h33169[23] &&
	      !sfdin__h33169[22] &&
	      !sfdin__h33169[21] &&
	      !sfdin__h33169[20] &&
	      !sfdin__h33169[19] &&
	      !sfdin__h33169[18] &&
	      !sfdin__h33169[17] &&
	      !sfdin__h33169[16] &&
	      !sfdin__h33169[15] &&
	      !sfdin__h33169[14] &&
	      !sfdin__h33169[13] &&
	      !sfdin__h33169[12] &&
	      !sfdin__h33169[11] &&
	      !sfdin__h33169[10] &&
	      !sfdin__h33169[9] &&
	      !sfdin__h33169[8] &&
	      !sfdin__h33169[7] &&
	      !sfdin__h33169[6] &&
	      !sfdin__h33169[5] &&
	      !sfdin__h33169[4] &&
	      !sfdin__h33169[3] &&
	      !sfdin__h33169[2] &&
	      !sfdin__h33169[1] &&
	      !sfdin__h33169[0]) ?
	       sfdin__h33169 :
	       _theResult___snd__h41437 ;
  assign _theResult___snd__h41437 =
	     { IF_0_CONCAT_IF_IF_fpu_div_fState_S3_first__16__ETC__q12[55:0],
	       2'd0 } ;
  assign _theResult___snd__h41455 =
	     sfdin__h33169 <<
	     IF_IF_fpu_div_fState_S3_first__16_BITS_120_TO__ETC___d812 ;
  assign _theResult___snd__h41460 =
	     sfdin__h33169 <<
	     IF_IF_fpu_div_fState_S3_first__16_BITS_120_TO__ETC___d810 ;
  assign _theResult___snd__h94767 = { fpu_sqr_fState_S3$D_OUT[57:0], 1'd0 } ;
  assign _theResult___snd__h94782 =
	     (!fpu_sqr_fState_S3$D_OUT[58] && fpu_sqr_fState_S3$D_OUT[57]) ?
	       _theResult___snd__h94784 :
	       _theResult___snd__h94797 ;
  assign _theResult___snd__h94784 = { fpu_sqr_fState_S3$D_OUT[56:0], 2'd0 } ;
  assign _theResult___snd__h94797 =
	     (!fpu_sqr_fState_S3$D_OUT[58] && !fpu_sqr_fState_S3$D_OUT[57] &&
	      !fpu_sqr_fState_S3$D_OUT[56] &&
	      !fpu_sqr_fState_S3$D_OUT[55] &&
	      !fpu_sqr_fState_S3$D_OUT[54] &&
	      !fpu_sqr_fState_S3$D_OUT[53] &&
	      !fpu_sqr_fState_S3$D_OUT[52] &&
	      !fpu_sqr_fState_S3$D_OUT[51] &&
	      !fpu_sqr_fState_S3$D_OUT[50] &&
	      !fpu_sqr_fState_S3$D_OUT[49] &&
	      !fpu_sqr_fState_S3$D_OUT[48] &&
	      !fpu_sqr_fState_S3$D_OUT[47] &&
	      !fpu_sqr_fState_S3$D_OUT[46] &&
	      !fpu_sqr_fState_S3$D_OUT[45] &&
	      !fpu_sqr_fState_S3$D_OUT[44] &&
	      !fpu_sqr_fState_S3$D_OUT[43] &&
	      !fpu_sqr_fState_S3$D_OUT[42] &&
	      !fpu_sqr_fState_S3$D_OUT[41] &&
	      !fpu_sqr_fState_S3$D_OUT[40] &&
	      !fpu_sqr_fState_S3$D_OUT[39] &&
	      !fpu_sqr_fState_S3$D_OUT[38] &&
	      !fpu_sqr_fState_S3$D_OUT[37] &&
	      !fpu_sqr_fState_S3$D_OUT[36] &&
	      !fpu_sqr_fState_S3$D_OUT[35] &&
	      !fpu_sqr_fState_S3$D_OUT[34] &&
	      !fpu_sqr_fState_S3$D_OUT[33] &&
	      !fpu_sqr_fState_S3$D_OUT[32] &&
	      !fpu_sqr_fState_S3$D_OUT[31] &&
	      !fpu_sqr_fState_S3$D_OUT[30] &&
	      !fpu_sqr_fState_S3$D_OUT[29] &&
	      !fpu_sqr_fState_S3$D_OUT[28] &&
	      !fpu_sqr_fState_S3$D_OUT[27] &&
	      !fpu_sqr_fState_S3$D_OUT[26] &&
	      !fpu_sqr_fState_S3$D_OUT[25] &&
	      !fpu_sqr_fState_S3$D_OUT[24] &&
	      !fpu_sqr_fState_S3$D_OUT[23] &&
	      !fpu_sqr_fState_S3$D_OUT[22] &&
	      !fpu_sqr_fState_S3$D_OUT[21] &&
	      !fpu_sqr_fState_S3$D_OUT[20] &&
	      !fpu_sqr_fState_S3$D_OUT[19] &&
	      !fpu_sqr_fState_S3$D_OUT[18] &&
	      !fpu_sqr_fState_S3$D_OUT[17] &&
	      !fpu_sqr_fState_S3$D_OUT[16] &&
	      !fpu_sqr_fState_S3$D_OUT[15] &&
	      !fpu_sqr_fState_S3$D_OUT[14] &&
	      !fpu_sqr_fState_S3$D_OUT[13] &&
	      !fpu_sqr_fState_S3$D_OUT[12] &&
	      !fpu_sqr_fState_S3$D_OUT[11] &&
	      !fpu_sqr_fState_S3$D_OUT[10] &&
	      !fpu_sqr_fState_S3$D_OUT[9] &&
	      !fpu_sqr_fState_S3$D_OUT[8] &&
	      !fpu_sqr_fState_S3$D_OUT[7] &&
	      !fpu_sqr_fState_S3$D_OUT[6] &&
	      !fpu_sqr_fState_S3$D_OUT[5] &&
	      !fpu_sqr_fState_S3$D_OUT[4] &&
	      !fpu_sqr_fState_S3$D_OUT[3] &&
	      !fpu_sqr_fState_S3$D_OUT[2] &&
	      !fpu_sqr_fState_S3$D_OUT[1] &&
	      !fpu_sqr_fState_S3$D_OUT[0]) ?
	       fpu_sqr_fState_S3$D_OUT[58:0] :
	       _theResult___snd__h94803 ;
  assign _theResult___snd__h94803 =
	     { IF_0_CONCAT_IF_fpu_sqr_fState_S3_first__375_BI_ETC__q19[56:0],
	       2'd0 } ;
  assign _theResult___snd__h94821 =
	     fpu_sqr_fState_S3$D_OUT[58:0] <<
	     IF_fpu_sqr_fState_S3_first__375_BITS_121_TO_11_ETC___d1632 ;
  assign _theResult___snd__h94826 =
	     fpu_sqr_fState_S3$D_OUT[58:0] <<
	     IF_fpu_sqr_fState_S3_first__375_BIT_58_384_THE_ETC___d1630 ;
  assign _theResult___snd_fst__h131051 =
	     { IF_sfdin30943_BIT_53_THEN_2_ELSE_0__q25[1],
	       { sfdin__h130943[52:0], 52'd0 } != 105'd0 } ;
  assign _theResult___snd_fst__h141477 =
	     { IF_sfdin41369_BIT_4_THEN_2_ELSE_0__q30[1],
	       { sfdin__h141369[3:0], 52'd0 } != 56'd0 } ;
  assign _theResult___snd_fst__h41490 =
	     { IF_sfdin1378_BIT_5_THEN_2_ELSE_0__q13[1],
	       { sfdin__h41378[4:0], 52'd0 } != 57'd0 } ;
  assign _theResult___snd_fst__h43500 =
	     IF_rg_index_1_87_ULE_58_91_THEN_NOT_rg_b_92_EQ_ETC___d1009 ?
	       _theResult___snd_fst__h43624 :
	       IF_rg_index_1_87_ULE_58_91_THEN_IF_rg_res_94_B_ETC___d1036 ;
  assign _theResult___snd_fst__h43539 =
	     (rg_res[116] || rg_b == 116'd0 ||
	      rg_s_014_ULT_rg_r_1_013_PLUS_rg_b_92_015___d1016) ?
	       rg_s :
	       s__h43680 ;
  assign _theResult___snd_fst__h43624 =
	     (IF_rg_index_1_87_ULE_58_91_THEN_IF_rg_res_94_B_ETC___d1002 ==
	      116'd0 ||
	      IF_rg_index_1_87_ULE_58_91_THEN_IF_rg_res_94_B_ETC___d1038) ?
	       IF_rg_index_1_87_ULE_58_91_THEN_IF_rg_res_94_B_ETC___d1036 :
	       s__h43745 ;
  assign _theResult___snd_fst__h94856 =
	     { IF_sfdin4744_BIT_6_THEN_2_ELSE_0__q20[1],
	       { sfdin__h94744[5:0], 52'd0 } != 58'd0 } ;
  assign _theResult___snd_fst_exp__h164063 =
	     _3970_MINUS_0_CONCAT_IF_iFifo_first__087_BIT_15_ETC___d3190 ?
	       11'd0 :
	       _theResult___fst_exp__h164060 ;
  assign _theResult___snd_fst_exp__h182405 =
	     SEXT_iFifo_first__087_BITS_167_TO_160_130_MINU_ETC___d3325 ?
	       _theResult___fst_exp__h173650 :
	       _theResult___fst_exp__h182402 ;
  assign _theResult___snd_fst_exp__h202701 =
	     _3970_MINUS_0_CONCAT_IF_iFifo_first__087_BIT_94_ETC___d4685 ?
	       11'd0 :
	       _theResult___fst_exp__h202698 ;
  assign _theResult___snd_fst_exp__h221043 =
	     SEXT_iFifo_first__087_BITS_102_TO_95_625_MINUS_ETC___d4808 ?
	       _theResult___fst_exp__h212288 :
	       _theResult___fst_exp__h221040 ;
  assign _theResult___snd_fst_exp__h241640 =
	     _3970_MINUS_0_CONCAT_IF_iFifo_first__087_BIT_29_ETC___d3910 ?
	       11'd0 :
	       _theResult___fst_exp__h241637 ;
  assign _theResult___snd_fst_exp__h259982 =
	     SEXT_iFifo_first__087_BITS_37_TO_30_850_MINUS__ETC___d4033 ?
	       _theResult___fst_exp__h251227 :
	       _theResult___fst_exp__h259979 ;
  assign _theResult___snd_fst_exp__h286904 =
	     _3074_MINUS_0_CONCAT_IF_resWire_wget__410_BIT_5_ETC___d5533 ?
	       _theResult___fst_exp__h278319 :
	       _theResult___fst_exp__h286901 ;
  assign _theResult___snd_fst_exp__h30385 =
	     (IF_fpu_div_fOperands_S0_first__6_BITS_129_TO_1_ETC___d285 ||
	      IF_fpu_div_fOperands_S0_first__6_BITS_129_TO_1_ETC___d429) ?
	       11'd0 :
	       value__h30425[10:0] ;
  assign _theResult___snd_fst_exp__h30388 =
	     IF_fpu_div_fOperands_S0_first__6_BITS_129_TO_1_ETC___d283 ?
	       _theResult___snd_fst_exp__h30385 :
	       11'd2046 ;
  assign _theResult___snd_fst_exp__h30412 =
	     fpu_div_fOperands_S0_first__6_BITS_129_TO_119__ETC___d428 ?
	       11'd0 :
	       _theResult___snd_fst_exp__h30388 ;
  assign _theResult___snd_fst_exp__h304724 =
	     SEXT_resWire_wget__410_BITS_67_TO_57_416_MINUS_ETC___d6033 ?
	       _theResult___fst_exp__h296085 :
	       _theResult___fst_exp__h304721 ;
  assign _theResult___snd_fst_sfd__h144484 =
	     (iFifo$D_OUT[159:137] == 23'd0) ?
	       52'h4000000000000 :
	       out___1_sfd__h144233 ;
  assign _theResult___snd_fst_sfd__h164064 =
	     _3970_MINUS_0_CONCAT_IF_iFifo_first__087_BIT_15_ETC___d3190 ?
	       52'd0 :
	       _theResult___fst_sfd__h164061 ;
  assign _theResult___snd_fst_sfd__h182406 =
	     SEXT_iFifo_first__087_BITS_167_TO_160_130_MINU_ETC___d3325 ?
	       _theResult___fst_sfd__h173651 :
	       _theResult___fst_sfd__h182403 ;
  assign _theResult___snd_fst_sfd__h183124 =
	     (iFifo$D_OUT[94:72] == 23'd0) ?
	       52'h4000000000000 :
	       out___1_sfd__h182873 ;
  assign _theResult___snd_fst_sfd__h202702 =
	     _3970_MINUS_0_CONCAT_IF_iFifo_first__087_BIT_94_ETC___d4685 ?
	       52'd0 :
	       _theResult___fst_sfd__h202699 ;
  assign _theResult___snd_fst_sfd__h221044 =
	     SEXT_iFifo_first__087_BITS_102_TO_95_625_MINUS_ETC___d4808 ?
	       _theResult___fst_sfd__h212289 :
	       _theResult___fst_sfd__h221041 ;
  assign _theResult___snd_fst_sfd__h222063 =
	     (iFifo$D_OUT[29:7] == 23'd0) ?
	       52'h4000000000000 :
	       out___1_sfd__h221812 ;
  assign _theResult___snd_fst_sfd__h241641 =
	     _3970_MINUS_0_CONCAT_IF_iFifo_first__087_BIT_29_ETC___d3910 ?
	       52'd0 :
	       _theResult___fst_sfd__h241638 ;
  assign _theResult___snd_fst_sfd__h259983 =
	     SEXT_iFifo_first__087_BITS_37_TO_30_850_MINUS__ETC___d4033 ?
	       _theResult___fst_sfd__h251228 :
	       _theResult___fst_sfd__h259980 ;
  assign _theResult___snd_fst_sfd__h261961 =
	     (resWire$wget[56:34] == 23'd0) ?
	       23'd2097152 :
	       resWire$wget[56:34] ;
  assign _theResult___snd_fst_sfd__h286905 =
	     _3074_MINUS_0_CONCAT_IF_resWire_wget__410_BIT_5_ETC___d5533 ?
	       _theResult___fst_sfd__h278320 :
	       _theResult___fst_sfd__h286902 ;
  assign _theResult___snd_fst_sfd__h30413 =
	     (fpu_div_fOperands_S0_first__6_BITS_129_TO_119__ETC___d428 ||
	      IF_fpu_div_fOperands_S0_first__6_BITS_129_TO_1_ETC___d283) ?
	       52'd0 :
	       52'hFFFFFFFFFFFFF ;
  assign _theResult___snd_fst_sfd__h304725 =
	     SEXT_resWire_wget__410_BITS_67_TO_57_416_MINUS_ETC___d6033 ?
	       _theResult___fst_sfd__h296086 :
	       _theResult___fst_sfd__h304722 ;
  assign _theResult___snd_snd__h131371 =
	     (fpu_madd_fProd_S3$D_OUT == 106'd0) ? 2'd0 : 2'd1 ;
  assign _theResult___snd_snd__h43671 =
	     rg_s_014_ULT_rg_r_1_013_PLUS_rg_b_92_015___d1016 ?
	       r__h43685 :
	       r__h43681 ;
  assign _theResult___snd_snd__h43737 =
	     IF_rg_index_1_87_ULE_58_91_THEN_IF_rg_res_94_B_ETC___d1038 ?
	       r__h43775 :
	       r__h43746 ;
  assign _theResult___snd_snd_snd__h131369 =
	     fpu_madd_fState_S3_first__995_BITS_12_TO_0_001_ETC___d2004 ?
	       _theResult___snd_snd__h131371 :
	       guardBC__h115666 ;
  assign _theResult___snd_snd_snd__h33014 =
	     (fpu_div_fState_S3$D_OUT[57:56] == 2'b0) ?
	       _theResult___snd__h33766 :
	       fpu_div_fState_S3$D_OUT[57:0] ;
  assign _theResult___snd_snd_snd__h43503 =
	     IF_rg_index_1_87_ULE_58_91_THEN_NOT_rg_b_92_EQ_ETC___d1009 ?
	       _theResult___snd_snd_snd__h43627 :
	       IF_rg_index_1_87_ULE_58_91_THEN_IF_rg_res_94_B_ETC___d1022 ;
  assign _theResult___snd_snd_snd__h43542 =
	     (rg_res[116] || rg_b == 116'd0) ?
	       rg_r_1 :
	       _theResult___snd_snd__h43671 ;
  assign _theResult___snd_snd_snd__h43627 =
	     (IF_rg_index_1_87_ULE_58_91_THEN_IF_rg_res_94_B_ETC___d1002 ==
	      116'd0) ?
	       IF_rg_index_1_87_ULE_58_91_THEN_IF_rg_res_94_B_ETC___d1022 :
	       _theResult___snd_snd__h43737 ;
  assign b___1__h77160 = 116'h40000000000000000000000000000 >> x__h85465 ;
  assign b__h10508 =
	     (fpu_div_fOperands_S0$D_OUT[65:55] == 11'd0) ?
	       (fpu_div_fOperands_S0$D_OUT[54] ?
		  6'd1 :
		  (fpu_div_fOperands_S0$D_OUT[53] ?
		     6'd2 :
		     (fpu_div_fOperands_S0$D_OUT[52] ?
			6'd3 :
			(fpu_div_fOperands_S0$D_OUT[51] ?
			   6'd4 :
			   (fpu_div_fOperands_S0$D_OUT[50] ?
			      6'd5 :
			      (fpu_div_fOperands_S0$D_OUT[49] ?
				 6'd6 :
				 (fpu_div_fOperands_S0$D_OUT[48] ?
				    6'd7 :
				    (fpu_div_fOperands_S0$D_OUT[47] ?
				       6'd8 :
				       (fpu_div_fOperands_S0$D_OUT[46] ?
					  6'd9 :
					  (fpu_div_fOperands_S0$D_OUT[45] ?
					     6'd10 :
					     (fpu_div_fOperands_S0$D_OUT[44] ?
						6'd11 :
						(fpu_div_fOperands_S0$D_OUT[43] ?
						   6'd12 :
						   (fpu_div_fOperands_S0$D_OUT[42] ?
						      6'd13 :
						      (fpu_div_fOperands_S0$D_OUT[41] ?
							 6'd14 :
							 (fpu_div_fOperands_S0$D_OUT[40] ?
							    6'd15 :
							    (fpu_div_fOperands_S0$D_OUT[39] ?
							       6'd16 :
							       (fpu_div_fOperands_S0$D_OUT[38] ?
								  6'd17 :
								  (fpu_div_fOperands_S0$D_OUT[37] ?
								     6'd18 :
								     (fpu_div_fOperands_S0$D_OUT[36] ?
									6'd19 :
									(fpu_div_fOperands_S0$D_OUT[35] ?
									   6'd20 :
									   (fpu_div_fOperands_S0$D_OUT[34] ?
									      6'd21 :
									      (fpu_div_fOperands_S0$D_OUT[33] ?
										 6'd22 :
										 (fpu_div_fOperands_S0$D_OUT[32] ?
										    6'd23 :
										    (fpu_div_fOperands_S0$D_OUT[31] ?
										       6'd24 :
										       (fpu_div_fOperands_S0$D_OUT[30] ?
											  6'd25 :
											  (fpu_div_fOperands_S0$D_OUT[29] ?
											     6'd26 :
											     (fpu_div_fOperands_S0$D_OUT[28] ?
												6'd27 :
												(fpu_div_fOperands_S0$D_OUT[27] ?
												   6'd28 :
												   (fpu_div_fOperands_S0$D_OUT[26] ?
												      6'd29 :
												      (fpu_div_fOperands_S0$D_OUT[25] ?
													 6'd30 :
													 (fpu_div_fOperands_S0$D_OUT[24] ?
													    6'd31 :
													    (fpu_div_fOperands_S0$D_OUT[23] ?
													       6'd32 :
													       (fpu_div_fOperands_S0$D_OUT[22] ?
														  6'd33 :
														  (fpu_div_fOperands_S0$D_OUT[21] ?
														     6'd34 :
														     (fpu_div_fOperands_S0$D_OUT[20] ?
															6'd35 :
															(fpu_div_fOperands_S0$D_OUT[19] ?
															   6'd36 :
															   (fpu_div_fOperands_S0$D_OUT[18] ?
															      6'd37 :
															      (fpu_div_fOperands_S0$D_OUT[17] ?
																 6'd38 :
																 (fpu_div_fOperands_S0$D_OUT[16] ?
																    6'd39 :
																    (fpu_div_fOperands_S0$D_OUT[15] ?
																       6'd40 :
																       (fpu_div_fOperands_S0$D_OUT[14] ?
																	  6'd41 :
																	  (fpu_div_fOperands_S0$D_OUT[13] ?
																	     6'd42 :
																	     (fpu_div_fOperands_S0$D_OUT[12] ?
																		6'd43 :
																		(fpu_div_fOperands_S0$D_OUT[11] ?
																		   6'd44 :
																		   (fpu_div_fOperands_S0$D_OUT[10] ?
																		      6'd45 :
																		      (fpu_div_fOperands_S0$D_OUT[9] ?
																			 6'd46 :
																			 (fpu_div_fOperands_S0$D_OUT[8] ?
																			    6'd47 :
																			    (fpu_div_fOperands_S0$D_OUT[7] ?
																			       6'd48 :
																			       (fpu_div_fOperands_S0$D_OUT[6] ?
																				  6'd49 :
																				  (fpu_div_fOperands_S0$D_OUT[5] ?
																				     6'd50 :
																				     (fpu_div_fOperands_S0$D_OUT[4] ?
																					6'd51 :
																					(fpu_div_fOperands_S0$D_OUT[3] ?
																					   6'd52 :
																					   6'd53)))))))))))))))))))))))))))))))))))))))))))))))))))) :
	       6'd0 ;
  assign b__h3090 =
	     (fpu_div_fOperands_S0$D_OUT[129:119] == 11'd0) ?
	       (fpu_div_fOperands_S0$D_OUT[118] ?
		  6'd1 :
		  (fpu_div_fOperands_S0$D_OUT[117] ?
		     6'd2 :
		     (fpu_div_fOperands_S0$D_OUT[116] ?
			6'd3 :
			(fpu_div_fOperands_S0$D_OUT[115] ?
			   6'd4 :
			   (fpu_div_fOperands_S0$D_OUT[114] ?
			      6'd5 :
			      (fpu_div_fOperands_S0$D_OUT[113] ?
				 6'd6 :
				 (fpu_div_fOperands_S0$D_OUT[112] ?
				    6'd7 :
				    (fpu_div_fOperands_S0$D_OUT[111] ?
				       6'd8 :
				       (fpu_div_fOperands_S0$D_OUT[110] ?
					  6'd9 :
					  (fpu_div_fOperands_S0$D_OUT[109] ?
					     6'd10 :
					     (fpu_div_fOperands_S0$D_OUT[108] ?
						6'd11 :
						(fpu_div_fOperands_S0$D_OUT[107] ?
						   6'd12 :
						   (fpu_div_fOperands_S0$D_OUT[106] ?
						      6'd13 :
						      (fpu_div_fOperands_S0$D_OUT[105] ?
							 6'd14 :
							 (fpu_div_fOperands_S0$D_OUT[104] ?
							    6'd15 :
							    (fpu_div_fOperands_S0$D_OUT[103] ?
							       6'd16 :
							       (fpu_div_fOperands_S0$D_OUT[102] ?
								  6'd17 :
								  (fpu_div_fOperands_S0$D_OUT[101] ?
								     6'd18 :
								     (fpu_div_fOperands_S0$D_OUT[100] ?
									6'd19 :
									(fpu_div_fOperands_S0$D_OUT[99] ?
									   6'd20 :
									   (fpu_div_fOperands_S0$D_OUT[98] ?
									      6'd21 :
									      (fpu_div_fOperands_S0$D_OUT[97] ?
										 6'd22 :
										 (fpu_div_fOperands_S0$D_OUT[96] ?
										    6'd23 :
										    (fpu_div_fOperands_S0$D_OUT[95] ?
										       6'd24 :
										       (fpu_div_fOperands_S0$D_OUT[94] ?
											  6'd25 :
											  (fpu_div_fOperands_S0$D_OUT[93] ?
											     6'd26 :
											     (fpu_div_fOperands_S0$D_OUT[92] ?
												6'd27 :
												(fpu_div_fOperands_S0$D_OUT[91] ?
												   6'd28 :
												   (fpu_div_fOperands_S0$D_OUT[90] ?
												      6'd29 :
												      (fpu_div_fOperands_S0$D_OUT[89] ?
													 6'd30 :
													 (fpu_div_fOperands_S0$D_OUT[88] ?
													    6'd31 :
													    (fpu_div_fOperands_S0$D_OUT[87] ?
													       6'd32 :
													       (fpu_div_fOperands_S0$D_OUT[86] ?
														  6'd33 :
														  (fpu_div_fOperands_S0$D_OUT[85] ?
														     6'd34 :
														     (fpu_div_fOperands_S0$D_OUT[84] ?
															6'd35 :
															(fpu_div_fOperands_S0$D_OUT[83] ?
															   6'd36 :
															   (fpu_div_fOperands_S0$D_OUT[82] ?
															      6'd37 :
															      (fpu_div_fOperands_S0$D_OUT[81] ?
																 6'd38 :
																 (fpu_div_fOperands_S0$D_OUT[80] ?
																    6'd39 :
																    (fpu_div_fOperands_S0$D_OUT[79] ?
																       6'd40 :
																       (fpu_div_fOperands_S0$D_OUT[78] ?
																	  6'd41 :
																	  (fpu_div_fOperands_S0$D_OUT[77] ?
																	     6'd42 :
																	     (fpu_div_fOperands_S0$D_OUT[76] ?
																		6'd43 :
																		(fpu_div_fOperands_S0$D_OUT[75] ?
																		   6'd44 :
																		   (fpu_div_fOperands_S0$D_OUT[74] ?
																		      6'd45 :
																		      (fpu_div_fOperands_S0$D_OUT[73] ?
																			 6'd46 :
																			 (fpu_div_fOperands_S0$D_OUT[72] ?
																			    6'd47 :
																			    (fpu_div_fOperands_S0$D_OUT[71] ?
																			       6'd48 :
																			       (fpu_div_fOperands_S0$D_OUT[70] ?
																				  6'd49 :
																				  (fpu_div_fOperands_S0$D_OUT[69] ?
																				     6'd50 :
																				     (fpu_div_fOperands_S0$D_OUT[68] ?
																					6'd51 :
																					(fpu_div_fOperands_S0$D_OUT[67] ?
																					   6'd52 :
																					   6'd53)))))))))))))))))))))))))))))))))))))))))))))))))))) :
	       6'd0 ;
  assign b__h31634 = { rg_d, 58'd0 } ;
  assign b__h43630 = { 2'd0, rg_b[115:2] } ;
  assign b__h43734 =
	     { 2'd0,
	       IF_rg_index_1_87_ULE_58_91_THEN_IF_rg_res_94_B_ETC___d1002[115:2] } ;
  assign din_exp30866_MINUS_1023__q23 = din_exp__h130866 - 11'd1023 ;
  assign din_exp__h130866 =
	     _7170_MINUS_fpu_madd_fState_S3_first__995_BITS__ETC___d2008 ?
	       value__h130883[10:0] :
	       11'd0 ;
  assign din_inc___2_exp__h142626 = fpu_madd_fState_S8$D_OUT[65:55] + 11'd1 ;
  assign din_inc___2_exp__h182467 = _theResult___fst_exp__h163334 + 11'd1 ;
  assign din_inc___2_exp__h182502 = _theResult___fst_exp__h172850 + 11'd1 ;
  assign din_inc___2_exp__h182528 = _theResult___fst_exp__h181651 + 11'd1 ;
  assign din_inc___2_exp__h221105 = _theResult___fst_exp__h201972 + 11'd1 ;
  assign din_inc___2_exp__h221140 = _theResult___fst_exp__h211488 + 11'd1 ;
  assign din_inc___2_exp__h221166 = _theResult___fst_exp__h220289 + 11'd1 ;
  assign din_inc___2_exp__h260044 = _theResult___fst_exp__h240911 + 11'd1 ;
  assign din_inc___2_exp__h260079 = _theResult___fst_exp__h250427 + 11'd1 ;
  assign din_inc___2_exp__h260105 = _theResult___fst_exp__h259228 + 11'd1 ;
  assign din_inc___2_exp__h304759 = _theResult___fst_exp__h277722 + 8'd1 ;
  assign din_inc___2_exp__h304785 = _theResult___fst_exp__h286378 + 8'd1 ;
  assign din_inc___2_exp__h304820 = _theResult___fst_exp__h295488 + 8'd1 ;
  assign din_inc___2_exp__h304846 = _theResult___fst_exp__h304173 + 8'd1 ;
  assign din_inc___2_exp__h42617 = fpu_div_fState_S4$D_OUT[64:54] + 11'd1 ;
  assign din_inc___2_exp__h96000 = fpu_sqr_fState_S4$D_OUT[64:54] + 11'd1 ;
  assign exp__h304742 =
	     (resWire$wget[67:57] == 11'd2047) ?
	       8'd255 :
	       _theResult___fst_exp__h304733 ;
  assign fpu_div_fOperands_S0D_OUT_BITS_129_TO_119_MIN_ETC__q7 =
	     fpu_div_fOperands_S0$D_OUT[129:119] - 11'd1023 ;
  assign fpu_div_fOperands_S0D_OUT_BITS_65_TO_55_MINUS_ETC__q8 =
	     fpu_div_fOperands_S0$D_OUT[65:55] - 11'd1023 ;
  assign fpu_div_fOperands_S0_first__6_BITS_129_TO_119__ETC___d293 =
	     fpu_div_fOperands_S0$D_OUT[129:119] == 11'd2047 &&
	     fpu_div_fOperands_S0$D_OUT[118:67] != 52'd0 &&
	     !fpu_div_fOperands_S0$D_OUT[118] ||
	     fpu_div_fOperands_S0$D_OUT[65:55] == 11'd2047 &&
	     fpu_div_fOperands_S0$D_OUT[54:3] != 52'd0 &&
	     !fpu_div_fOperands_S0$D_OUT[54] ||
	     fpu_div_fOperands_S0$D_OUT[129:119] == 11'd2047 &&
	     fpu_div_fOperands_S0$D_OUT[118] ||
	     fpu_div_fOperands_S0$D_OUT[65:55] == 11'd2047 &&
	     fpu_div_fOperands_S0$D_OUT[54] ||
	     fpu_div_fOperands_S0_first__6_BITS_65_TO_55_6__ETC___d289 ;
  assign fpu_div_fOperands_S0_first__6_BITS_129_TO_119__ETC___d331 =
	     fpu_div_fOperands_S0$D_OUT[129:119] == 11'd2047 &&
	     fpu_div_fOperands_S0$D_OUT[118:67] == 52'd0 ||
	     fpu_div_fOperands_S0$D_OUT[129:119] == 11'd0 &&
	     fpu_div_fOperands_S0$D_OUT[118:67] == 52'd0 ||
	     fpu_div_fOperands_S0$D_OUT[65:55] == 11'd2047 &&
	     fpu_div_fOperands_S0$D_OUT[54:3] == 52'd0 ;
  assign fpu_div_fOperands_S0_first__6_BITS_129_TO_119__ETC___d366 =
	     fpu_div_fOperands_S0$D_OUT[129:119] == 11'd2047 &&
	     fpu_div_fOperands_S0$D_OUT[118:67] == 52'd0 &&
	     fpu_div_fOperands_S0$D_OUT[65:55] == 11'd2047 &&
	     fpu_div_fOperands_S0$D_OUT[54:3] == 52'd0 ||
	     fpu_div_fOperands_S0$D_OUT[129:119] == 11'd0 &&
	     fpu_div_fOperands_S0$D_OUT[118:67] == 52'd0 &&
	     fpu_div_fOperands_S0$D_OUT[65:55] == 11'd0 &&
	     fpu_div_fOperands_S0$D_OUT[54:3] == 52'd0 ;
  assign fpu_div_fOperands_S0_first__6_BITS_129_TO_119__ETC___d428 =
	     fpu_div_fOperands_S0$D_OUT[129:119] == 11'd2047 &&
	     fpu_div_fOperands_S0$D_OUT[118:67] != 52'd0 &&
	     !fpu_div_fOperands_S0$D_OUT[118] ||
	     fpu_div_fOperands_S0$D_OUT[65:55] == 11'd2047 &&
	     fpu_div_fOperands_S0$D_OUT[54:3] != 52'd0 &&
	     !fpu_div_fOperands_S0$D_OUT[54] ||
	     fpu_div_fOperands_S0$D_OUT[129:119] == 11'd2047 &&
	     fpu_div_fOperands_S0$D_OUT[118] ||
	     fpu_div_fOperands_S0$D_OUT[65:55] == 11'd2047 &&
	     fpu_div_fOperands_S0$D_OUT[54] ||
	     fpu_div_fOperands_S0$D_OUT[65:55] == 11'd0 &&
	     fpu_div_fOperands_S0$D_OUT[54:3] == 52'd0 ||
	     fpu_div_fOperands_S0_first__6_BITS_129_TO_119__ETC___d331 ;
  assign fpu_div_fOperands_S0_first__6_BITS_65_TO_55_6__ETC___d289 =
	     fpu_div_fOperands_S0$D_OUT[65:55] == 11'd0 &&
	     fpu_div_fOperands_S0$D_OUT[54:3] == 52'd0 ||
	     fpu_div_fOperands_S0$D_OUT[129:119] == 11'd2047 &&
	     fpu_div_fOperands_S0$D_OUT[118:67] == 52'd0 ||
	     fpu_div_fOperands_S0$D_OUT[129:119] == 11'd0 &&
	     fpu_div_fOperands_S0$D_OUT[118:67] == 52'd0 ||
	     fpu_div_fOperands_S0$D_OUT[65:55] == 11'd2047 &&
	     fpu_div_fOperands_S0$D_OUT[54:3] == 52'd0 ||
	     !IF_fpu_div_fOperands_S0_first__6_BITS_129_TO_1_ETC___d283 ||
	     IF_fpu_div_fOperands_S0_first__6_BITS_129_TO_1_ETC___d285 ;
  assign fpu_div_fOperands_S0_first__6_BIT_130_33_EQ_fp_ETC___d335 =
	     fpu_div_fOperands_S0$D_OUT[130] ==
	     fpu_div_fOperands_S0$D_OUT[66] ;
  assign fpu_div_fState_S3_first__16_BIT_121_37_CONCAT__ETC___d866 =
	     { fpu_div_fState_S3$D_OUT[121],
	       IF_fpu_div_fState_S3_first__16_BITS_120_TO_110_ETC___d527 ?
		 IF_IF_fpu_div_fState_S3_first__16_BITS_120_TO__ETC___d859 :
		 ((fpu_div_fState_S3$D_OUT[120:110] == 11'd2047) ?
		    ((fpu_div_fState_S3$D_OUT[57:56] == 2'b0) ?
		       { _theResult___fst_exp__h41335,
			 fpu_div_fState_S3$D_OUT[109:58] } :
		       63'h7FEFFFFFFFFFFFFF) :
		    fpu_div_fState_S3$D_OUT[120:58]) } ;
  assign fpu_madd_fOperand_S0D_OUT_BITS_129_TO_119_MIN_ETC__q128 =
	     fpu_madd_fOperand_S0$D_OUT[129:119] - 11'd1023 ;
  assign fpu_madd_fOperand_S0D_OUT_BITS_65_TO_55_MINUS_ETC__q129 =
	     fpu_madd_fOperand_S0$D_OUT[65:55] - 11'd1023 ;
  assign fpu_madd_fOperand_S0_first__803_BITS_129_TO_11_ETC___d1857 =
	     fpu_madd_fOperand_S0$D_OUT[129:119] == 11'd2047 &&
	     fpu_madd_fOperand_S0$D_OUT[118:67] == 52'd0 ||
	     fpu_madd_fOperand_S0$D_OUT[65:55] == 11'd2047 &&
	     fpu_madd_fOperand_S0$D_OUT[54:3] == 52'd0 ||
	     x__h96539 == 11'd0 && _theResult___fst_sfd__h96608 == 52'd0 &&
	     (fpu_madd_fOperand_S0$D_OUT[129:119] == 11'd0 &&
	      fpu_madd_fOperand_S0$D_OUT[118:67] == 52'd0 ||
	      fpu_madd_fOperand_S0$D_OUT[65:55] == 11'd0 &&
	      fpu_madd_fOperand_S0$D_OUT[54:3] == 52'd0) &&
	     fpu_madd_fOperand_S0_first__803_BIT_195_804_AN_ETC___d1855 ;
  assign fpu_madd_fOperand_S0_first__803_BITS_129_TO_11_ETC___d1926 =
	     fpu_madd_fOperand_S0$D_OUT[129:119] == 11'd2047 &&
	     fpu_madd_fOperand_S0$D_OUT[118:67] == 52'd0 &&
	     fpu_madd_fOperand_S0$D_OUT[65:55] == 11'd0 &&
	     fpu_madd_fOperand_S0$D_OUT[54:3] == 52'd0 ||
	     fpu_madd_fOperand_S0$D_OUT[129:119] == 11'd0 &&
	     fpu_madd_fOperand_S0$D_OUT[118:67] == 52'd0 &&
	     fpu_madd_fOperand_S0$D_OUT[65:55] == 11'd2047 &&
	     fpu_madd_fOperand_S0$D_OUT[54:3] == 52'd0 ;
  assign fpu_madd_fOperand_S0_first__803_BIT_195_804_AN_ETC___d1855 =
	     (fpu_madd_fOperand_S0$D_OUT[195] &&
	      fpu_madd_fOperand_S0$D_OUT[194]) ==
	     NOT_fpu_madd_fOperand_S0_first__803_BIT_130_85_ETC___d1854 ;
  assign fpu_madd_fProd_S3_first__009_SRL_IF_7170_MINUS_ETC___d2012 =
	     fpu_madd_fProd_S3$D_OUT >>
	     _7170_MINUS_fpu_madd_fState_S3_first__995_BITS__ETC___d2007 ;
  assign fpu_madd_fState_S3_first__995_BITS_12_TO_0_001_ETC___d2002 =
	     (fpu_madd_fState_S3$D_OUT[12:0] ^ 13'h1000) <= 13'd5119 ;
  assign fpu_madd_fState_S3_first__995_BITS_12_TO_0_001_ETC___d2004 =
	     (fpu_madd_fState_S3$D_OUT[12:0] ^ 13'h1000) < 13'd3020 ;
  assign fpu_madd_fState_S3_first__995_BITS_86_TO_82_00_ETC___d2501 =
	     fpu_madd_fState_S3$D_OUT[86:82] |
	     { 2'd0,
	       sfdBC__h115662[105] &&
	       IF_IF_7170_MINUS_fpu_madd_fState_S3_first__995_ETC___d2031 ==
	       12'd1023,
	       _theResult___fst_exp__h130952 == 11'd0 &&
	       guardBC__h115666 != 2'd0,
	       sfdBC__h115662[105] &&
	       IF_IF_7170_MINUS_fpu_madd_fState_S3_first__995_ETC___d2031 ==
	       12'd1023 } ;
  assign fpu_madd_fState_S4D_OUT_BITS_128_TO_118_MINUS_ETC__q26 =
	     fpu_madd_fState_S4$D_OUT[128:118] - 11'd1023 ;
  assign fpu_madd_fState_S4D_OUT_BITS_64_TO_54_MINUS_1023__q27 =
	     fpu_madd_fState_S4$D_OUT[64:54] - 11'd1023 ;
  assign fpu_madd_fState_S5_first__601_BITS_56_TO_0_610_ETC___d2615 =
	     fpu_madd_fState_S5$D_OUT[56:0] >>
	     fpu_madd_fState_S5$D_OUT[126:114] ;
  assign fpu_madd_fState_S7_first__651_BITS_137_TO_133__ETC___d2942 =
	     fpu_madd_fState_S7$D_OUT[137:133] |
	     { 2'd0,
	       sfd__h133119[56] &&
	       IF_fpu_madd_fState_S7_first__651_BITS_126_TO_1_ETC___d2668 ==
	       12'd1023,
	       _theResult___fst_exp__h141378 == 11'd0 &&
	       guard__h133123 != 2'd0,
	       sfd__h133119[56] &&
	       IF_fpu_madd_fState_S7_first__651_BITS_126_TO_1_ETC___d2668 ==
	       12'd1023 } ;
  assign fpu_madd_fState_S8_first__960_BITS_75_TO_71_03_ETC___d3043 =
	     fpu_madd_fState_S8$D_OUT[75:71] |
	     { 2'd0,
	       IF_fpu_madd_fState_S8_first__960_BITS_65_TO_55_ETC___d3011 ==
	       11'd2047 &&
	       ((fpu_madd_fState_S8$D_OUT[65:55] == 11'd2047) ?
		  fpu_madd_fState_S8$D_OUT[54:3] :
		  _theResult___fst_sfd__h142620) ==
	       52'd0,
	       1'd0,
	       fpu_madd_fState_S8$D_OUT[65:55] != 11'd2047 &&
	       fpu_madd_fState_S8$D_OUT[2:1] != 2'b0 } ;
  assign fpu_sqr_fOperand_S0D_OUT_BITS_65_TO_55_MINUS__ETC__q16 =
	     fpu_sqr_fOperand_S0$D_OUT[65:55] - 11'd1023 ;
  assign fpu_sqr_fState_S3D_OUT_BITS_121_TO_111_MINUS__ETC__q18 =
	     fpu_sqr_fState_S3$D_OUT[121:111] - 11'd1023 ;
  assign guardBC__h115666 =
	     (sfdBC__h115662[105] &&
	      IF_IF_7170_MINUS_fpu_madd_fState_S3_first__995_ETC___d2031 ==
	      12'd1023) ?
	       2'd3 :
	       _theResult___snd_fst__h131051 ;
  assign guard__h132367 = fpu_madd_fState_S5$D_OUT[56:0] << x__h132471 ;
  assign guard__h133123 =
	     (sfd__h133119[56] &&
	      IF_fpu_madd_fState_S7_first__651_BITS_126_TO_1_ETC___d2668 ==
	      12'd1023) ?
	       2'd3 :
	       _theResult___snd_fst__h141477 ;
  assign guard__h155373 =
	     { IF_theResult___snd63285_BIT_4_THEN_2_ELSE_0__q34[1],
	       { _theResult___snd__h163285[3:0], 52'd0 } != 56'd0 } ;
  assign guard__h164622 =
	     { IF_sfdin72844_BIT_4_THEN_2_ELSE_0__q38[1],
	       { sfdin__h172844[3:0], 52'd0 } != 56'd0 } ;
  assign guard__h165220 = x__h165322 != 57'd0 ;
  assign guard__h173661 =
	     { IF_theResult___snd81597_BIT_4_THEN_2_ELSE_0__q41[1],
	       { _theResult___snd__h181597[3:0], 52'd0 } != 56'd0 } ;
  assign guard__h194011 =
	     { IF_theResult___snd01923_BIT_4_THEN_2_ELSE_0__q94[1],
	       { _theResult___snd__h201923[3:0], 52'd0 } != 56'd0 } ;
  assign guard__h203260 =
	     { IF_sfdin11482_BIT_4_THEN_2_ELSE_0__q98[1],
	       { sfdin__h211482[3:0], 52'd0 } != 56'd0 } ;
  assign guard__h203858 = x__h203960 != 57'd0 ;
  assign guard__h212299 =
	     { IF_theResult___snd20235_BIT_4_THEN_2_ELSE_0__q101[1],
	       { _theResult___snd__h220235[3:0], 52'd0 } != 56'd0 } ;
  assign guard__h232950 =
	     { IF_theResult___snd40862_BIT_4_THEN_2_ELSE_0__q61[1],
	       { _theResult___snd__h240862[3:0], 52'd0 } != 56'd0 } ;
  assign guard__h242199 =
	     { IF_sfdin50421_BIT_4_THEN_2_ELSE_0__q65[1],
	       { sfdin__h250421[3:0], 52'd0 } != 56'd0 } ;
  assign guard__h242797 = x__h242899 != 57'd0 ;
  assign guard__h251238 =
	     { IF_theResult___snd59174_BIT_4_THEN_2_ELSE_0__q68[1],
	       { _theResult___snd__h259174[3:0], 52'd0 } != 56'd0 } ;
  assign guard__h269623 =
	     { IF_sfdin77716_BIT_33_THEN_2_ELSE_0__q134[1],
	       { sfdin__h277716[32:0], 23'd0 } != 56'd0 } ;
  assign guard__h278330 =
	     { IF_theResult___snd86329_BIT_33_THEN_2_ELSE_0__q136[1],
	       { _theResult___snd__h286329[32:0], 23'd0 } != 56'd0 } ;
  assign guard__h287260 =
	     { IF_sfdin95482_BIT_33_THEN_2_ELSE_0__q140[1],
	       { sfdin__h295482[32:0], 23'd0 } != 56'd0 } ;
  assign guard__h287858 = x__h287960 != 57'd0 ;
  assign guard__h296096 =
	     { IF_theResult___snd04119_BIT_33_THEN_2_ELSE_0__q143[1],
	       { _theResult___snd__h304119[32:0], 23'd0 } != 56'd0 } ;
  assign guard__h32997 = x__h41756 ;
  assign guard__h86435 = x__h95138 ;
  assign iFifoD_OUT_BITS_102_TO_95_MINUS_127__q95 =
	     iFifo$D_OUT[102:95] - 8'd127 ;
  assign iFifoD_OUT_BITS_167_TO_160_MINUS_127__q35 =
	     iFifo$D_OUT[167:160] - 8'd127 ;
  assign iFifoD_OUT_BITS_37_TO_30_MINUS_127__q62 =
	     iFifo$D_OUT[37:30] - 8'd127 ;
  assign out___1_sfd__h144233 = { iFifo$D_OUT[159:137], 29'd0 } ;
  assign out___1_sfd__h182873 = { iFifo$D_OUT[94:72], 29'd0 } ;
  assign out___1_sfd__h221812 = { iFifo$D_OUT[29:7], 29'd0 } ;
  assign out_exp__h142544 =
	     fpu_madd_fState_S8$D_OUT[3] ?
	       _theResult___exp__h142541 :
	       fpu_madd_fState_S8$D_OUT[65:55] ;
  assign out_exp__h163982 =
	     _theResult___snd__h163285[5] ?
	       _theResult___exp__h163979 :
	       _theResult___fst_exp__h163334 ;
  assign out_exp__h173572 =
	     sfdin__h172844[5] ?
	       _theResult___exp__h173569 :
	       _theResult___fst_exp__h172850 ;
  assign out_exp__h182324 =
	     _theResult___snd__h181597[5] ?
	       _theResult___exp__h182321 :
	       _theResult___fst_exp__h181651 ;
  assign out_exp__h202620 =
	     _theResult___snd__h201923[5] ?
	       _theResult___exp__h202617 :
	       _theResult___fst_exp__h201972 ;
  assign out_exp__h212210 =
	     sfdin__h211482[5] ?
	       _theResult___exp__h212207 :
	       _theResult___fst_exp__h211488 ;
  assign out_exp__h220962 =
	     _theResult___snd__h220235[5] ?
	       _theResult___exp__h220959 :
	       _theResult___fst_exp__h220289 ;
  assign out_exp__h241559 =
	     _theResult___snd__h240862[5] ?
	       _theResult___exp__h241556 :
	       _theResult___fst_exp__h240911 ;
  assign out_exp__h251149 =
	     sfdin__h250421[5] ?
	       _theResult___exp__h251146 :
	       _theResult___fst_exp__h250427 ;
  assign out_exp__h259901 =
	     _theResult___snd__h259174[5] ?
	       _theResult___exp__h259898 :
	       _theResult___fst_exp__h259228 ;
  assign out_exp__h278241 =
	     sfdin__h277716[34] ?
	       _theResult___exp__h278238 :
	       _theResult___fst_exp__h277722 ;
  assign out_exp__h286823 =
	     _theResult___snd__h286329[34] ?
	       _theResult___exp__h286820 :
	       _theResult___fst_exp__h286378 ;
  assign out_exp__h296007 =
	     sfdin__h295482[34] ?
	       _theResult___exp__h296004 :
	       _theResult___fst_exp__h295488 ;
  assign out_exp__h304643 =
	     _theResult___snd__h304119[34] ?
	       _theResult___exp__h304640 :
	       _theResult___fst_exp__h304173 ;
  assign out_exp__h42529 =
	     fpu_div_fState_S4$D_OUT[2] ?
	       _theResult___exp__h42526 :
	       fpu_div_fState_S4$D_OUT[64:54] ;
  assign out_exp__h95912 =
	     fpu_sqr_fState_S4$D_OUT[2] ?
	       _theResult___exp__h95909 :
	       fpu_sqr_fState_S4$D_OUT[64:54] ;
  assign out_sfd__h142545 =
	     fpu_madd_fState_S8$D_OUT[3] ?
	       _theResult___sfd__h142542 :
	       fpu_madd_fState_S8$D_OUT[54:3] ;
  assign out_sfd__h163983 =
	     _theResult___snd__h163285[5] ?
	       _theResult___sfd__h163980 :
	       _theResult___snd__h163285[56:5] ;
  assign out_sfd__h173573 =
	     sfdin__h172844[5] ?
	       _theResult___sfd__h173570 :
	       sfdin__h172844[56:5] ;
  assign out_sfd__h182325 =
	     _theResult___snd__h181597[5] ?
	       _theResult___sfd__h182322 :
	       _theResult___snd__h181597[56:5] ;
  assign out_sfd__h202621 =
	     _theResult___snd__h201923[5] ?
	       _theResult___sfd__h202618 :
	       _theResult___snd__h201923[56:5] ;
  assign out_sfd__h212211 =
	     sfdin__h211482[5] ?
	       _theResult___sfd__h212208 :
	       sfdin__h211482[56:5] ;
  assign out_sfd__h220963 =
	     _theResult___snd__h220235[5] ?
	       _theResult___sfd__h220960 :
	       _theResult___snd__h220235[56:5] ;
  assign out_sfd__h241560 =
	     _theResult___snd__h240862[5] ?
	       _theResult___sfd__h241557 :
	       _theResult___snd__h240862[56:5] ;
  assign out_sfd__h251150 =
	     sfdin__h250421[5] ?
	       _theResult___sfd__h251147 :
	       sfdin__h250421[56:5] ;
  assign out_sfd__h259902 =
	     _theResult___snd__h259174[5] ?
	       _theResult___sfd__h259899 :
	       _theResult___snd__h259174[56:5] ;
  assign out_sfd__h278242 =
	     sfdin__h277716[34] ?
	       _theResult___sfd__h278239 :
	       sfdin__h277716[56:34] ;
  assign out_sfd__h286824 =
	     _theResult___snd__h286329[34] ?
	       _theResult___sfd__h286821 :
	       _theResult___snd__h286329[56:34] ;
  assign out_sfd__h296008 =
	     sfdin__h295482[34] ?
	       _theResult___sfd__h296005 :
	       sfdin__h295482[56:34] ;
  assign out_sfd__h304644 =
	     _theResult___snd__h304119[34] ?
	       _theResult___sfd__h304641 :
	       _theResult___snd__h304119[56:34] ;
  assign out_sfd__h42530 =
	     fpu_div_fState_S4$D_OUT[2] ?
	       _theResult___sfd__h42527 :
	       fpu_div_fState_S4$D_OUT[53:2] ;
  assign out_sfd__h95913 =
	     fpu_sqr_fState_S4$D_OUT[2] ?
	       _theResult___sfd__h95910 :
	       fpu_sqr_fState_S4$D_OUT[53:2] ;
  assign r__h43681 = r__h43685 + rg_b ;
  assign r__h43685 = { 1'd0, rg_r_1[115:1] } ;
  assign r__h43746 =
	     r__h43775 +
	     IF_rg_index_1_87_ULE_58_91_THEN_IF_rg_res_94_B_ETC___d1002 ;
  assign r__h43775 =
	     { 1'd0,
	       IF_rg_index_1_87_ULE_58_91_THEN_IF_rg_res_94_B_ETC___d1022[115:1] } ;
  assign resWire_wget__410_BITS_4_TO_0_658_OR_NOT_resWi_ETC___d6768 =
	     resWire$wget[4:0] |
	     { (resWire$wget[67:57] != 11'd2047 ||
		resWire$wget[56:5] == 52'd0) &&
	       (resWire$wget[67:57] != 11'd2047 ||
		resWire$wget[56:5] != 52'd0) &&
	       (resWire$wget[67:57] != 11'd0 ||
		resWire$wget[56:5] != 52'd0) &&
	       IF_resWire_wget__410_BITS_67_TO_57_416_EQ_0_42_ETC___d6709,
	       (resWire$wget[67:57] != 11'd2047 ||
		resWire$wget[56:5] == 52'd0) &&
	       (resWire$wget[67:57] != 11'd2047 ||
		resWire$wget[56:5] != 52'd0) &&
	       (resWire$wget[67:57] != 11'd0 ||
		resWire$wget[56:5] != 52'd0) &&
	       IF_resWire_wget__410_BITS_67_TO_57_416_EQ_0_42_ETC___d6720,
	       (resWire$wget[67:57] != 11'd2047 ||
		resWire$wget[56:5] == 52'd0) &&
	       (resWire$wget[67:57] != 11'd2047 ||
		resWire$wget[56:5] != 52'd0) &&
	       (resWire$wget[67:57] != 11'd0 ||
		resWire$wget[56:5] != 52'd0) &&
	       IF_resWire_wget__410_BITS_67_TO_57_416_EQ_0_42_ETC___d6736,
	       (resWire$wget[67:57] != 11'd2047 ||
		resWire$wget[56:5] == 52'd0) &&
	       (resWire$wget[67:57] != 11'd2047 ||
		resWire$wget[56:5] != 52'd0) &&
	       (resWire$wget[67:57] != 11'd0 ||
		resWire$wget[56:5] != 52'd0) &&
	       IF_resWire_wget__410_BITS_67_TO_57_416_EQ_0_42_ETC___d6749,
	       (resWire$wget[67:57] != 11'd2047 ||
		resWire$wget[56:5] == 52'd0) &&
	       (resWire$wget[67:57] != 11'd2047 ||
		resWire$wget[56:5] != 52'd0) &&
	       (resWire$wget[67:57] != 11'd0 ||
		resWire$wget[56:5] != 52'd0) &&
	       IF_resWire_wget__410_BITS_67_TO_57_416_EQ_0_42_ETC___d6762 } ;
  assign resWirewget_BITS_67_TO_57_MINUS_1023__q137 =
	     resWire$wget[67:57] - 11'd1023 ;
  assign result__h132372 =
	     { fpu_madd_fState_S5_first__601_BITS_56_TO_0_610_ETC___d2615[56:1],
	       fpu_madd_fState_S5_first__601_BITS_56_TO_0_610_ETC___d2615[0] |
	       guard__h132367 != 57'd0 } ;
  assign result__h165225 =
	     { _0b0_CONCAT_NOT_iFifo_first__087_BITS_167_TO_16_ETC___d3330[56:1],
	       _0b0_CONCAT_NOT_iFifo_first__087_BITS_167_TO_16_ETC___d3330[0] |
	       guard__h165220 } ;
  assign result__h203863 =
	     { _0b0_CONCAT_NOT_iFifo_first__087_BITS_102_TO_95_ETC___d4813[56:1],
	       _0b0_CONCAT_NOT_iFifo_first__087_BITS_102_TO_95_ETC___d4813[0] |
	       guard__h203858 } ;
  assign result__h242802 =
	     { _0b0_CONCAT_NOT_iFifo_first__087_BITS_37_TO_30__ETC___d4038[56:1],
	       _0b0_CONCAT_NOT_iFifo_first__087_BITS_37_TO_30__ETC___d4038[0] |
	       guard__h242797 } ;
  assign result__h287863 =
	     { _0b0_CONCAT_NOT_resWire_wget__410_BITS_67_TO_57_ETC___d6038[56:1],
	       _0b0_CONCAT_NOT_resWire_wget__410_BITS_67_TO_57_ETC___d6038[0] |
	       guard__h287858 } ;
  assign result__h31668 = { _theResult____h31574[57:1], 1'd1 } ;
  assign result__h31699 =
	     { 1'd0,
	       value__h31712[56:1],
	       value__h31712[0] | sfdlsb__h31694 } ;
  assign result__h31874 =
	     (IF_rg_r_BIT_115_THEN_rg_q_PLUS_NEG_INV_rg_q_89_ETC__q10[56:0] ==
	      57'd0) ?
	       58'd0 :
	       58'd1 ;
  assign result__h85925 = { x__h85931[58:1], 1'd1 } ;
  assign rg_index_1_87_PLUS_1_89_ULE_58___d990 = rg_index_1 + 6'd1 <= 6'd58 ;
  assign rg_index_1_87_ULE_58___d991 = rg_index_1 <= 6'd58 ;
  assign rg_index_PLUS_1_ULE_57___d6 = rg_index + 6'd1 <= 6'd57 ;
  assign rg_index_ULE_57___d7 = rg_index <= 6'd57 ;
  assign rg_q_PLUS_NEG_INV_rg_q_89_90___d491 = rg_q + -(~rg_q) ;
  assign rg_s_014_ULT_rg_r_1_013_PLUS_rg_b_92_015___d1016 =
	     rg_s < sum__h43628 ;
  assign s__h43680 = rg_s - sum__h43628 ;
  assign s__h43745 =
	     IF_rg_index_1_87_ULE_58_91_THEN_IF_rg_res_94_B_ETC___d1036 -
	     sum__h43732 ;
  assign sfdA__h1086 =
	     { fpu_div_fOperands_S0$D_OUT[129:119] != 11'd0,
	       fpu_div_fOperands_S0$D_OUT[118:67] } ;
  assign sfdA__h1090 = sfdA__h1086 << b__h3090 ;
  assign sfdA__h131577 =
	     { 1'b0,
	       fpu_madd_fState_S4$D_OUT[128:118] != 11'd0,
	       fpu_madd_fState_S4$D_OUT[117:66],
	       3'b0 } ;
  assign sfdBC__h115662 =
	     _7170_MINUS_fpu_madd_fState_S3_first__995_BITS__ETC___d2008 ?
	       fpu_madd_fProd_S3$D_OUT :
	       _theResult___fst__h116827 ;
  assign sfdBC__h131578 =
	     { 1'b0,
	       fpu_madd_fState_S4$D_OUT[64:54] != 11'd0,
	       fpu_madd_fState_S4$D_OUT[53:0],
	       1'b0 } ;
  assign sfdB__h1087 =
	     { fpu_div_fOperands_S0$D_OUT[65:55] != 11'd0,
	       fpu_div_fOperands_S0$D_OUT[54:3] } ;
  assign sfdB__h1092 = sfdB__h1087 << b__h10508 ;
  assign sfd___1__h60702 = { 1'd0, sfd__h44953[57:1] } ;
  assign sfd__h133119 =
	     fpu_madd_fState_S7$D_OUT[128] ?
	       fpu_madd_fState_S7$D_OUT[56:0] :
	       fpu_madd_fState_S7$D_OUT[113:57] ;
  assign sfd__h142040 =
	     { 1'b0,
	       fpu_madd_fState_S8$D_OUT[65:55] != 11'd0,
	       fpu_madd_fState_S8$D_OUT[54:3] } +
	     54'd1 ;
  assign sfd__h144534 = { value__h148921, 32'd0 } ;
  assign sfd__h163352 =
	     { 1'b0,
	       _theResult___fst_exp__h163334 != 11'd0,
	       _theResult___snd__h163285[56:5] } +
	     54'd1 ;
  assign sfd__h172942 =
	     { 1'b0,
	       _theResult___fst_exp__h172850 != 11'd0,
	       sfdin__h172844[56:5] } +
	     54'd1 ;
  assign sfd__h17985 = { 1'd1, fpu_div_fOperands_S0$D_OUT[117:67] } ;
  assign sfd__h17988 = { 1'd1, fpu_div_fOperands_S0$D_OUT[53:3] } ;
  assign sfd__h181670 =
	     { 1'b0,
	       _theResult___fst_exp__h181651 != 11'd0,
	       _theResult___snd__h181597[56:5] } +
	     54'd1 ;
  assign sfd__h183174 = { value__h187559, 32'd0 } ;
  assign sfd__h201990 =
	     { 1'b0,
	       _theResult___fst_exp__h201972 != 11'd0,
	       _theResult___snd__h201923[56:5] } +
	     54'd1 ;
  assign sfd__h211580 =
	     { 1'b0,
	       _theResult___fst_exp__h211488 != 11'd0,
	       sfdin__h211482[56:5] } +
	     54'd1 ;
  assign sfd__h220308 =
	     { 1'b0,
	       _theResult___fst_exp__h220289 != 11'd0,
	       _theResult___snd__h220235[56:5] } +
	     54'd1 ;
  assign sfd__h222113 = { value__h226498, 32'd0 } ;
  assign sfd__h240929 =
	     { 1'b0,
	       _theResult___fst_exp__h240911 != 11'd0,
	       _theResult___snd__h240862[56:5] } +
	     54'd1 ;
  assign sfd__h250519 =
	     { 1'b0,
	       _theResult___fst_exp__h250427 != 11'd0,
	       sfdin__h250421[56:5] } +
	     54'd1 ;
  assign sfd__h259247 =
	     { 1'b0,
	       _theResult___fst_exp__h259228 != 11'd0,
	       _theResult___snd__h259174[56:5] } +
	     54'd1 ;
  assign sfd__h262011 = { value__h270233, 3'd0 } ;
  assign sfd__h277814 =
	     { 1'b0,
	       _theResult___fst_exp__h277722 != 8'd0,
	       sfdin__h277716[56:34] } +
	     25'd1 ;
  assign sfd__h286396 =
	     { 1'b0,
	       _theResult___fst_exp__h286378 != 8'd0,
	       _theResult___snd__h286329[56:34] } +
	     25'd1 ;
  assign sfd__h295580 =
	     { 1'b0,
	       _theResult___fst_exp__h295488 != 8'd0,
	       sfdin__h295482[56:34] } +
	     25'd1 ;
  assign sfd__h304192 =
	     { 1'b0,
	       _theResult___fst_exp__h304173 != 8'd0,
	       _theResult___snd__h304119[56:34] } +
	     25'd1 ;
  assign sfd__h304743 =
	     (resWire$wget[67:57] == 11'd2047 &&
	      resWire$wget[56:5] != 52'd0) ?
	       _theResult___snd_fst_sfd__h261961 :
	       _theResult___fst_sfd__h304737 ;
  assign sfd__h42033 =
	     { 1'b0,
	       fpu_div_fState_S4$D_OUT[64:54] != 11'd0,
	       fpu_div_fState_S4$D_OUT[53:2] } +
	     54'd1 ;
  assign sfd__h44951 = { value__h53174, 4'd0 } ;
  assign sfd__h44953 = sfd__h44951 << x__h60732 ;
  assign sfd__h45004 = { 1'd1, fpu_sqr_fOperand_S0$D_OUT[53:3] } ;
  assign sfd__h95416 =
	     { 1'b0,
	       fpu_sqr_fState_S4$D_OUT[64:54] != 11'd0,
	       fpu_sqr_fState_S4$D_OUT[53:2] } +
	     54'd1 ;
  assign sfd__h99402 = { 1'd1, _theResult___fst_sfd__h96608[50:0] } ;
  assign sfd__h99405 = { 1'd1, fpu_madd_fOperand_S0$D_OUT[117:67] } ;
  assign sfd__h99408 = { 1'd1, fpu_madd_fOperand_S0$D_OUT[53:3] } ;
  assign sfdin__h130943 =
	     sfdBC__h115662[105] ?
	       _theResult___snd__h130966 :
	       _theResult___snd__h130980 ;
  assign sfdin__h141369 =
	     sfd__h133119[56] ?
	       _theResult___snd__h141392 :
	       _theResult___snd__h141406 ;
  assign sfdin__h172844 =
	     _theResult____h164612[56] ?
	       _theResult___snd__h172861 :
	       _theResult___snd__h172872 ;
  assign sfdin__h211482 =
	     _theResult____h203250[56] ?
	       _theResult___snd__h211499 :
	       _theResult___snd__h211510 ;
  assign sfdin__h250421 =
	     _theResult____h242189[56] ?
	       _theResult___snd__h250438 :
	       _theResult___snd__h250449 ;
  assign sfdin__h277716 =
	     _theResult____h269613[56] ?
	       _theResult___snd__h277733 :
	       _theResult___snd__h277744 ;
  assign sfdin__h295482 =
	     _theResult____h287250[56] ?
	       _theResult___snd__h295499 :
	       _theResult___snd__h295510 ;
  assign sfdin__h33169 =
	     (fpu_div_fState_S3$D_OUT[120:110] == 11'd2047) ?
	       _theResult___snd_snd_snd__h33014 :
	       fpu_div_fState_S3$D_OUT[57:0] ;
  assign sfdin__h41378 =
	     sfdin__h33169[57] ?
	       _theResult___snd__h41401 :
	       _theResult___snd__h41416 ;
  assign sfdin__h94744 =
	     fpu_sqr_fState_S3$D_OUT[58] ?
	       _theResult___snd__h94767 :
	       _theResult___snd__h94782 ;
  assign sfdlsb__h116825 = x__h116896 != 106'd0 ;
  assign sfdlsb__h31694 = x__h31813 != 58'd0 ;
  assign sum__h43628 = rg_r_1 + rg_b ;
  assign sum__h43732 =
	     IF_rg_index_1_87_ULE_58_91_THEN_IF_rg_res_94_B_ETC___d1022 +
	     IF_rg_index_1_87_ULE_58_91_THEN_IF_rg_res_94_B_ETC___d1002 ;
  assign theResult___fst_exp1341_MINUS_1023__q11 =
	     _theResult___fst_exp__h41341 - 11'd1023 ;
  assign value41307_BITS_10_TO_0_MINUS_1023__q28 =
	     value__h141307[10:0] - 11'd1023 ;
  assign value_BIT_52___h53270 = fpu_sqr_fOperand_S0$D_OUT[65:55] != 11'd0 ;
  assign value__h130883 = fpu_madd_fState_S3$D_OUT[12:0] + 13'd1023 ;
  assign value__h141307 = fpu_madd_fState_S7$D_OUT[126:114] + 13'd1023 ;
  assign value__h148921 =
	     { 1'b0, iFifo$D_OUT[167:160] != 8'd0, iFifo$D_OUT[159:137] } ;
  assign value__h187559 =
	     { 1'b0, iFifo$D_OUT[102:95] != 8'd0, iFifo$D_OUT[94:72] } ;
  assign value__h226498 =
	     { 1'b0, iFifo$D_OUT[37:30] != 8'd0, iFifo$D_OUT[29:7] } ;
  assign value__h270233 =
	     { 1'b0, resWire$wget[67:57] != 11'd0, resWire$wget[56:5] } ;
  assign value__h30425 =
	     IF_fpu_div_fOperands_S0_first__6_BITS_129_TO_1_ETC___d282 +
	     13'd1023 ;
  assign value__h30480 = { 1'b0, sfdA__h1090 } ;
  assign value__h30601 =
	     13'd7170 -
	     IF_fpu_div_fOperands_S0_first__6_BITS_129_TO_1_ETC___d282 ;
  assign value__h31592 = rg_r[115] ? rg_r + b__h31634 : rg_r ;
  assign value__h31712 =
	     IF_rg_r_BIT_115_THEN_rg_q_PLUS_NEG_INV_rg_q_89_ETC__q10[56:0] >>
	     fpu_div_fState_S2$D_OUT[10:0] ;
  assign value__h53174 =
	     { 1'b0,
	       value_BIT_52___h53270,
	       fpu_sqr_fOperand_S0$D_OUT[54:3] } ;
  assign x__h114243 =
	     { fpu_madd_fOperand_S0$D_OUT[129:119] != 11'd0,
	       fpu_madd_fOperand_S0$D_OUT[118:67] } ;
  assign x__h114255 =
	     { fpu_madd_fOperand_S0$D_OUT[65:55] != 11'd0,
	       fpu_madd_fOperand_S0$D_OUT[54:3] } ;
  assign x__h116896 = fpu_madd_fProd_S3$D_OUT << x__h116929 ;
  assign x__h116929 =
	     13'd106 -
	     _7170_MINUS_fpu_madd_fState_S3_first__995_BITS__ETC___d2007 ;
  assign x__h131406 =
	     fpu_madd_fState_S3_first__995_BITS_12_TO_0_001_ETC___d2002 ?
	       _theResult___snd_snd_snd__h131369 :
	       2'd3 ;
  assign x__h131940 =
	     { 1'b0,
	       NOT_fpu_madd_fState_S4_first__547_BIT_130_553__ETC___d2584 ?
		 { fpu_madd_fState_S4$D_OUT[64:54] != 11'd0,
		   fpu_madd_fState_S4$D_OUT[53:0],
		   1'b0 } :
		 { fpu_madd_fState_S4$D_OUT[128:118] != 11'd0,
		   fpu_madd_fState_S4$D_OUT[117:66],
		   3'b0 } } ;
  assign x__h131944 =
	     { 1'b0,
	       NOT_fpu_madd_fState_S4_first__547_BIT_130_553__ETC___d2584 ?
		 { fpu_madd_fState_S4$D_OUT[128:118] != 11'd0,
		   fpu_madd_fState_S4$D_OUT[117:66],
		   3'b0 } :
		 { fpu_madd_fState_S4$D_OUT[64:54] != 11'd0,
		   fpu_madd_fState_S4$D_OUT[53:0],
		   1'b0 } } ;
  assign x__h132359 =
	     fpu_madd_fState_S5$D_OUT[215] ?
	       fpu_madd_fState_S5$D_OUT[56:0] :
	       (((fpu_madd_fState_S5$D_OUT[126:114] ^ 13'h1000) < 13'd4153) ?
		  result__h132372 :
		  ((fpu_madd_fState_S5$D_OUT[56:0] == 57'd0) ?
		     fpu_madd_fState_S5$D_OUT[56:0] :
		     57'd1)) ;
  assign x__h132471 = 13'd57 - fpu_madd_fState_S5$D_OUT[126:114] ;
  assign x__h132871 =
	     fpu_madd_fState_S6$D_OUT[113:57] +
	     fpu_madd_fState_S6$D_OUT[56:0] ;
  assign x__h132880 =
	     fpu_madd_fState_S6$D_OUT[113:57] -
	     fpu_madd_fState_S6$D_OUT[56:0] ;
  assign x__h141760 = fpu_madd_fState_S7$D_OUT[202] ? 2'd0 : guard__h133123 ;
  assign x__h165322 = sfd__h144534 << x__h165355 ;
  assign x__h165355 =
	     12'd57 -
	     _3074_MINUS_SEXT_iFifo_first__087_BITS_167_TO_1_ETC___d3326 ;
  assign x__h203960 = sfd__h183174 << x__h203993 ;
  assign x__h203993 =
	     12'd57 -
	     _3074_MINUS_SEXT_iFifo_first__087_BITS_102_TO_9_ETC___d4809 ;
  assign x__h242899 = sfd__h222113 << x__h242932 ;
  assign x__h242932 =
	     12'd57 -
	     _3074_MINUS_SEXT_iFifo_first__087_BITS_37_TO_30_ETC___d4034 ;
  assign x__h287960 = sfd__h262011 << x__h287993 ;
  assign x__h287993 =
	     12'd57 -
	     _3970_MINUS_SEXT_resWire_wget__410_BITS_67_TO_5_ETC___d6034 ;
  assign x__h30477 = { value__h30480, 60'd0 } ;
  assign x__h30538 = { sfdB__h1092, 4'b0 } ;
  assign x__h30592 =
	     fpu_div_fOperands_S0_first__6_BITS_129_TO_119__ETC___d293 ?
	       11'd0 :
	       _theResult___fst__h30373 ;
  assign x__h31813 =
	     { 1'd0,
	       IF_rg_r_BIT_115_THEN_rg_q_PLUS_NEG_INV_rg_q_89_ETC__q10[56:0] } <<
	     x__h31820 ;
  assign x__h31820 = 11'd58 - fpu_div_fState_S2$D_OUT[10:0] ;
  assign x__h32103 =
	     (value__h31592[114:58] == 57'd0) ?
	       _theResult____h31574 :
	       result__h31668 ;
  assign x__h41756 =
	     (sfdin__h33169[57] &&
	      IF_IF_fpu_div_fState_S3_first__16_BITS_120_TO__ETC___d573 ==
	      12'd1023) ?
	       2'd3 :
	       _theResult___snd_fst__h41490 ;
  assign x__h52551 = x__h52569 + 13'd1024 ;
  assign x__h52569 =
	     { IF_fpu_sqr_fOperand_S0_first__059_BITS_65_TO_5_ETC__q17[11],
	       IF_fpu_sqr_fOperand_S0_first__059_BITS_65_TO_5_ETC__q17 } ;
  assign x__h60693 =
	     IF_fpu_sqr_fOperand_S0_first__059_BITS_65_TO_5_ETC___d1195[0] ?
	       sfd__h44953 :
	       sfd___1__h60702 ;
  assign x__h60732 =
	     IF_fpu_sqr_fOperand_S0_first__059_BITS_65_TO_5_ETC___d1193 -
	     6'd1 ;
  assign x__h85465 =
	     IF_fpu_sqr_fState_S1_first__216_BIT_57_226_THE_ETC___d1342[0] ?
	       IF_fpu_sqr_fState_S1_first__216_BIT_57_226_THE_ETC___d1342 +
	       7'd1 :
	       IF_fpu_sqr_fState_S1_first__216_BIT_57_226_THE_ETC___d1342 ;
  assign x__h85931 = rg_res[116] ? rg_res[115:0] : 116'd0 ;
  assign x__h86149 = (rg_s == 116'd0) ? x__h85931[58:0] : result__h85925 ;
  assign x__h95138 =
	     (fpu_sqr_fState_S3$D_OUT[58] &&
	      IF_fpu_sqr_fState_S3_first__375_BITS_121_TO_11_ETC___d1389 ==
	      12'd1023) ?
	       2'd3 :
	       _theResult___snd_fst__h94856 ;
  assign x__h96539 =
	     fpu_madd_fOperand_S0$D_OUT[195] ?
	       fpu_madd_fOperand_S0$D_OUT[193:183] :
	       11'd0 ;
  always@(fpu_div_fState_S4$D_OUT or
	  out_sfd__h42530 or _theResult___sfd__h42527)
  begin
    case (fpu_div_fState_S4$D_OUT[1:0])
      2'b0, 2'b01:
	  CASE_fpu_div_fState_S4D_OUT_BITS_1_TO_0_0b0_f_ETC__q1 =
	      fpu_div_fState_S4$D_OUT[53:2];
      2'b10:
	  CASE_fpu_div_fState_S4D_OUT_BITS_1_TO_0_0b0_f_ETC__q1 =
	      out_sfd__h42530;
      2'b11:
	  CASE_fpu_div_fState_S4D_OUT_BITS_1_TO_0_0b0_f_ETC__q1 =
	      _theResult___sfd__h42527;
    endcase
  end
  always@(fpu_div_fState_S4$D_OUT or _theResult___sfd__h42527)
  begin
    case (fpu_div_fState_S4$D_OUT[1:0])
      2'b0:
	  CASE_fpu_div_fState_S4D_OUT_BITS_1_TO_0_0b0_f_ETC__q2 =
	      fpu_div_fState_S4$D_OUT[53:2];
      2'b01, 2'b10, 2'b11:
	  CASE_fpu_div_fState_S4D_OUT_BITS_1_TO_0_0b0_f_ETC__q2 =
	      _theResult___sfd__h42527;
    endcase
  end
  always@(fpu_div_fState_S4$D_OUT or
	  CASE_fpu_div_fState_S4D_OUT_BITS_1_TO_0_0b0_f_ETC__q1 or
	  CASE_fpu_div_fState_S4D_OUT_BITS_1_TO_0_0b0_f_ETC__q2 or
	  _theResult___sfd__h42527)
  begin
    case (fpu_div_fState_S4$D_OUT[68:66])
      3'd0:
	  _theResult___fst_sfd__h42605 =
	      CASE_fpu_div_fState_S4D_OUT_BITS_1_TO_0_0b0_f_ETC__q1;
      3'd1:
	  _theResult___fst_sfd__h42605 =
	      CASE_fpu_div_fState_S4D_OUT_BITS_1_TO_0_0b0_f_ETC__q2;
      3'd2:
	  _theResult___fst_sfd__h42605 =
	      (fpu_div_fState_S4$D_OUT[1:0] == 2'b0 ||
	       fpu_div_fState_S4$D_OUT[65]) ?
		fpu_div_fState_S4$D_OUT[53:2] :
		_theResult___sfd__h42527;
      3'd3:
	  _theResult___fst_sfd__h42605 =
	      (fpu_div_fState_S4$D_OUT[1:0] == 2'b0) ?
		fpu_div_fState_S4$D_OUT[53:2] :
		(fpu_div_fState_S4$D_OUT[65] ?
		   _theResult___sfd__h42527 :
		   fpu_div_fState_S4$D_OUT[53:2]);
      3'd4: _theResult___fst_sfd__h42605 = fpu_div_fState_S4$D_OUT[53:2];
      default: _theResult___fst_sfd__h42605 = 52'd0;
    endcase
  end
  always@(fpu_sqr_fState_S4$D_OUT or
	  out_sfd__h95913 or _theResult___sfd__h95910)
  begin
    case (fpu_sqr_fState_S4$D_OUT[1:0])
      2'b0, 2'b01:
	  CASE_fpu_sqr_fState_S4D_OUT_BITS_1_TO_0_0b0_f_ETC__q3 =
	      fpu_sqr_fState_S4$D_OUT[53:2];
      2'b10:
	  CASE_fpu_sqr_fState_S4D_OUT_BITS_1_TO_0_0b0_f_ETC__q3 =
	      out_sfd__h95913;
      2'b11:
	  CASE_fpu_sqr_fState_S4D_OUT_BITS_1_TO_0_0b0_f_ETC__q3 =
	      _theResult___sfd__h95910;
    endcase
  end
  always@(fpu_sqr_fState_S4$D_OUT or _theResult___sfd__h95910)
  begin
    case (fpu_sqr_fState_S4$D_OUT[1:0])
      2'b0:
	  CASE_fpu_sqr_fState_S4D_OUT_BITS_1_TO_0_0b0_f_ETC__q4 =
	      fpu_sqr_fState_S4$D_OUT[53:2];
      2'b01, 2'b10, 2'b11:
	  CASE_fpu_sqr_fState_S4D_OUT_BITS_1_TO_0_0b0_f_ETC__q4 =
	      _theResult___sfd__h95910;
    endcase
  end
  always@(fpu_sqr_fState_S4$D_OUT or
	  CASE_fpu_sqr_fState_S4D_OUT_BITS_1_TO_0_0b0_f_ETC__q3 or
	  CASE_fpu_sqr_fState_S4D_OUT_BITS_1_TO_0_0b0_f_ETC__q4 or
	  _theResult___sfd__h95910)
  begin
    case (fpu_sqr_fState_S4$D_OUT[68:66])
      3'd0:
	  _theResult___fst_sfd__h95988 =
	      CASE_fpu_sqr_fState_S4D_OUT_BITS_1_TO_0_0b0_f_ETC__q3;
      3'd1:
	  _theResult___fst_sfd__h95988 =
	      CASE_fpu_sqr_fState_S4D_OUT_BITS_1_TO_0_0b0_f_ETC__q4;
      3'd2:
	  _theResult___fst_sfd__h95988 =
	      (fpu_sqr_fState_S4$D_OUT[1:0] == 2'b0 ||
	       fpu_sqr_fState_S4$D_OUT[65]) ?
		fpu_sqr_fState_S4$D_OUT[53:2] :
		_theResult___sfd__h95910;
      3'd3:
	  _theResult___fst_sfd__h95988 =
	      (fpu_sqr_fState_S4$D_OUT[1:0] == 2'b0) ?
		fpu_sqr_fState_S4$D_OUT[53:2] :
		(fpu_sqr_fState_S4$D_OUT[65] ?
		   _theResult___sfd__h95910 :
		   fpu_sqr_fState_S4$D_OUT[53:2]);
      3'd4: _theResult___fst_sfd__h95988 = fpu_sqr_fState_S4$D_OUT[53:2];
      default: _theResult___fst_sfd__h95988 = 52'd0;
    endcase
  end
  always@(fpu_madd_fState_S8$D_OUT or
	  out_sfd__h142545 or _theResult___sfd__h142542)
  begin
    case (fpu_madd_fState_S8$D_OUT[2:1])
      2'b0, 2'b01:
	  CASE_fpu_madd_fState_S8D_OUT_BITS_2_TO_1_0b0__ETC__q5 =
	      fpu_madd_fState_S8$D_OUT[54:3];
      2'b10:
	  CASE_fpu_madd_fState_S8D_OUT_BITS_2_TO_1_0b0__ETC__q5 =
	      out_sfd__h142545;
      2'b11:
	  CASE_fpu_madd_fState_S8D_OUT_BITS_2_TO_1_0b0__ETC__q5 =
	      _theResult___sfd__h142542;
    endcase
  end
  always@(fpu_madd_fState_S8$D_OUT or _theResult___sfd__h142542)
  begin
    case (fpu_madd_fState_S8$D_OUT[2:1])
      2'b0:
	  CASE_fpu_madd_fState_S8D_OUT_BITS_2_TO_1_0b0__ETC__q6 =
	      fpu_madd_fState_S8$D_OUT[54:3];
      2'b01, 2'b10, 2'b11:
	  CASE_fpu_madd_fState_S8D_OUT_BITS_2_TO_1_0b0__ETC__q6 =
	      _theResult___sfd__h142542;
    endcase
  end
  always@(fpu_madd_fState_S8$D_OUT or
	  CASE_fpu_madd_fState_S8D_OUT_BITS_2_TO_1_0b0__ETC__q5 or
	  CASE_fpu_madd_fState_S8D_OUT_BITS_2_TO_1_0b0__ETC__q6 or
	  _theResult___sfd__h142542)
  begin
    case (fpu_madd_fState_S8$D_OUT[70:68])
      3'd0:
	  _theResult___fst_sfd__h142620 =
	      CASE_fpu_madd_fState_S8D_OUT_BITS_2_TO_1_0b0__ETC__q5;
      3'd1:
	  _theResult___fst_sfd__h142620 =
	      CASE_fpu_madd_fState_S8D_OUT_BITS_2_TO_1_0b0__ETC__q6;
      3'd2:
	  _theResult___fst_sfd__h142620 =
	      (fpu_madd_fState_S8$D_OUT[2:1] == 2'b0 ||
	       fpu_madd_fState_S8$D_OUT[66]) ?
		fpu_madd_fState_S8$D_OUT[54:3] :
		_theResult___sfd__h142542;
      3'd3:
	  _theResult___fst_sfd__h142620 =
	      (fpu_madd_fState_S8$D_OUT[2:1] == 2'b0) ?
		fpu_madd_fState_S8$D_OUT[54:3] :
		(fpu_madd_fState_S8$D_OUT[66] ?
		   _theResult___sfd__h142542 :
		   fpu_madd_fState_S8$D_OUT[54:3]);
      3'd4: _theResult___fst_sfd__h142620 = fpu_madd_fState_S8$D_OUT[54:3];
      default: _theResult___fst_sfd__h142620 = 52'd0;
    endcase
  end
  always@(iFifo$D_OUT)
  begin
    case (iFifo$D_OUT[6:4])
      3'd0, 3'd1: _theResult___fst_exp__h148289 = 11'd2047;
      3'd2:
	  _theResult___fst_exp__h148289 =
	      iFifo$D_OUT[168] ? 11'd2046 : 11'd2047;
      3'd3:
	  _theResult___fst_exp__h148289 =
	      iFifo$D_OUT[168] ? 11'd2047 : 11'd2046;
      3'd4: _theResult___fst_exp__h148289 = 11'd2046;
      default: _theResult___fst_exp__h148289 = 11'd0;
    endcase
  end
  always@(iFifo$D_OUT)
  begin
    case (iFifo$D_OUT[6:4])
      3'd0, 3'd1: _theResult___fst_sfd__h148290 = 52'd0;
      3'd2:
	  _theResult___fst_sfd__h148290 =
	      iFifo$D_OUT[168] ? 52'hFFFFFFFFFFFFF : 52'd0;
      3'd3:
	  _theResult___fst_sfd__h148290 =
	      iFifo$D_OUT[168] ? 52'd0 : 52'hFFFFFFFFFFFFF;
      3'd4: _theResult___fst_sfd__h148290 = 52'hFFFFFFFFFFFFF;
      default: _theResult___fst_sfd__h148290 = 52'd0;
    endcase
  end
  always@(iFifo$D_OUT)
  begin
    case (iFifo$D_OUT[6:4])
      3'd0, 3'd1: _theResult___fst_exp__h186929 = 11'd2047;
      3'd2:
	  _theResult___fst_exp__h186929 =
	      iFifo$D_OUT[103] ? 11'd2046 : 11'd2047;
      3'd3:
	  _theResult___fst_exp__h186929 =
	      iFifo$D_OUT[103] ? 11'd2047 : 11'd2046;
      3'd4: _theResult___fst_exp__h186929 = 11'd2046;
      default: _theResult___fst_exp__h186929 = 11'd0;
    endcase
  end
  always@(iFifo$D_OUT)
  begin
    case (iFifo$D_OUT[6:4])
      3'd0, 3'd1: _theResult___fst_exp__h225868 = 11'd2047;
      3'd2:
	  _theResult___fst_exp__h225868 =
	      iFifo$D_OUT[38] ? 11'd2046 : 11'd2047;
      3'd3:
	  _theResult___fst_exp__h225868 =
	      iFifo$D_OUT[38] ? 11'd2047 : 11'd2046;
      3'd4: _theResult___fst_exp__h225868 = 11'd2046;
      default: _theResult___fst_exp__h225868 = 11'd0;
    endcase
  end
  always@(iFifo$D_OUT)
  begin
    case (iFifo$D_OUT[6:4])
      3'd0, 3'd1: _theResult___fst_sfd__h186930 = 52'd0;
      3'd2:
	  _theResult___fst_sfd__h186930 =
	      iFifo$D_OUT[103] ? 52'hFFFFFFFFFFFFF : 52'd0;
      3'd3:
	  _theResult___fst_sfd__h186930 =
	      iFifo$D_OUT[103] ? 52'd0 : 52'hFFFFFFFFFFFFF;
      3'd4: _theResult___fst_sfd__h186930 = 52'hFFFFFFFFFFFFF;
      default: _theResult___fst_sfd__h186930 = 52'd0;
    endcase
  end
  always@(iFifo$D_OUT)
  begin
    case (iFifo$D_OUT[6:4])
      3'd0, 3'd1: _theResult___fst_sfd__h225869 = 52'd0;
      3'd2:
	  _theResult___fst_sfd__h225869 =
	      iFifo$D_OUT[38] ? 52'hFFFFFFFFFFFFF : 52'd0;
      3'd3:
	  _theResult___fst_sfd__h225869 =
	      iFifo$D_OUT[38] ? 52'd0 : 52'hFFFFFFFFFFFFF;
      3'd4: _theResult___fst_sfd__h225869 = 52'hFFFFFFFFFFFFF;
      default: _theResult___fst_sfd__h225869 = 52'd0;
    endcase
  end
  always@(fpu_div_fOperands_S0$D_OUT or
	  fpu_div_fOperands_S0_first__6_BIT_130_33_EQ_fp_ETC___d335)
  begin
    case (fpu_div_fOperands_S0$D_OUT[2:0])
      3'd0, 3'd1: _theResult___fst_exp__h18518 = 11'd2047;
      3'd2:
	  _theResult___fst_exp__h18518 =
	      fpu_div_fOperands_S0_first__6_BIT_130_33_EQ_fp_ETC___d335 ?
		11'd2047 :
		11'd2046;
      3'd3:
	  _theResult___fst_exp__h18518 =
	      fpu_div_fOperands_S0_first__6_BIT_130_33_EQ_fp_ETC___d335 ?
		11'd2046 :
		11'd2047;
      3'd4: _theResult___fst_exp__h18518 = 11'd2046;
      default: _theResult___fst_exp__h18518 = 11'd0;
    endcase
  end
  always@(fpu_div_fOperands_S0$D_OUT or
	  fpu_div_fOperands_S0_first__6_BIT_130_33_EQ_fp_ETC___d335)
  begin
    case (fpu_div_fOperands_S0$D_OUT[2:0])
      3'd0, 3'd1: _theResult___fst_sfd__h18519 = 52'd0;
      3'd2:
	  _theResult___fst_sfd__h18519 =
	      fpu_div_fOperands_S0_first__6_BIT_130_33_EQ_fp_ETC___d335 ?
		52'd0 :
		52'hFFFFFFFFFFFFF;
      3'd3:
	  _theResult___fst_sfd__h18519 =
	      fpu_div_fOperands_S0_first__6_BIT_130_33_EQ_fp_ETC___d335 ?
		52'hFFFFFFFFFFFFF :
		52'd0;
      3'd4: _theResult___fst_sfd__h18519 = 52'hFFFFFFFFFFFFF;
      default: _theResult___fst_sfd__h18519 = 52'd0;
    endcase
  end
  always@(fpu_div_fOperands_S0$D_OUT or
	  fpu_div_fOperands_S0_first__6_BIT_130_33_EQ_fp_ETC___d335)
  begin
    case (fpu_div_fOperands_S0$D_OUT[2:0])
      3'd0: _theResult___fst_sfd__h19008 = 52'd0;
      3'd1: _theResult___fst_sfd__h19008 = 52'd1;
      3'd2:
	  _theResult___fst_sfd__h19008 =
	      fpu_div_fOperands_S0_first__6_BIT_130_33_EQ_fp_ETC___d335 ?
		52'd1 :
		52'd0;
      3'd3:
	  _theResult___fst_sfd__h19008 =
	      fpu_div_fOperands_S0_first__6_BIT_130_33_EQ_fp_ETC___d335 ?
		52'd0 :
		52'd1;
      default: _theResult___fst_sfd__h19008 = 52'd0;
    endcase
  end
  always@(fpu_div_fOperands_S0$D_OUT or
	  fpu_div_fOperands_S0_first__6_BIT_130_33_EQ_fp_ETC___d335)
  begin
    case (fpu_div_fOperands_S0$D_OUT[2:0])
      3'd0, 3'd1, 3'd2, 3'd3:
	  CASE_fpu_div_fOperands_S0D_OUT_BITS_2_TO_0_0__ETC__q9 =
	      !fpu_div_fOperands_S0_first__6_BIT_130_33_EQ_fp_ETC___d335;
      default: CASE_fpu_div_fOperands_S0D_OUT_BITS_2_TO_0_0__ETC__q9 =
		   fpu_div_fOperands_S0$D_OUT[2:0] == 3'd4 &&
		   !fpu_div_fOperands_S0_first__6_BIT_130_33_EQ_fp_ETC___d335;
    endcase
  end
  always@(fpu_div_fState_S4$D_OUT or
	  out_exp__h42529 or _theResult___exp__h42526)
  begin
    case (fpu_div_fState_S4$D_OUT[1:0])
      2'b0, 2'b01:
	  CASE_fpu_div_fState_S4D_OUT_BITS_1_TO_0_0b0_f_ETC__q14 =
	      fpu_div_fState_S4$D_OUT[64:54];
      2'b10:
	  CASE_fpu_div_fState_S4D_OUT_BITS_1_TO_0_0b0_f_ETC__q14 =
	      out_exp__h42529;
      2'b11:
	  CASE_fpu_div_fState_S4D_OUT_BITS_1_TO_0_0b0_f_ETC__q14 =
	      _theResult___exp__h42526;
    endcase
  end
  always@(fpu_div_fState_S4$D_OUT or _theResult___exp__h42526)
  begin
    case (fpu_div_fState_S4$D_OUT[1:0])
      2'b0:
	  CASE_fpu_div_fState_S4D_OUT_BITS_1_TO_0_0b0_f_ETC__q15 =
	      fpu_div_fState_S4$D_OUT[64:54];
      2'b01, 2'b10, 2'b11:
	  CASE_fpu_div_fState_S4D_OUT_BITS_1_TO_0_0b0_f_ETC__q15 =
	      _theResult___exp__h42526;
    endcase
  end
  always@(fpu_div_fState_S4$D_OUT or
	  CASE_fpu_div_fState_S4D_OUT_BITS_1_TO_0_0b0_f_ETC__q14 or
	  CASE_fpu_div_fState_S4D_OUT_BITS_1_TO_0_0b0_f_ETC__q15 or
	  _theResult___exp__h42526)
  begin
    case (fpu_div_fState_S4$D_OUT[68:66])
      3'd0:
	  _theResult___fst_exp__h42604 =
	      CASE_fpu_div_fState_S4D_OUT_BITS_1_TO_0_0b0_f_ETC__q14;
      3'd1:
	  _theResult___fst_exp__h42604 =
	      CASE_fpu_div_fState_S4D_OUT_BITS_1_TO_0_0b0_f_ETC__q15;
      3'd2:
	  _theResult___fst_exp__h42604 =
	      (fpu_div_fState_S4$D_OUT[1:0] == 2'b0 ||
	       fpu_div_fState_S4$D_OUT[65]) ?
		fpu_div_fState_S4$D_OUT[64:54] :
		_theResult___exp__h42526;
      3'd3:
	  _theResult___fst_exp__h42604 =
	      (fpu_div_fState_S4$D_OUT[1:0] == 2'b0) ?
		fpu_div_fState_S4$D_OUT[64:54] :
		(fpu_div_fState_S4$D_OUT[65] ?
		   _theResult___exp__h42526 :
		   fpu_div_fState_S4$D_OUT[64:54]);
      3'd4: _theResult___fst_exp__h42604 = fpu_div_fState_S4$D_OUT[64:54];
      default: _theResult___fst_exp__h42604 = 11'd0;
    endcase
  end
  always@(fpu_sqr_fState_S4$D_OUT or
	  out_exp__h95912 or _theResult___exp__h95909)
  begin
    case (fpu_sqr_fState_S4$D_OUT[1:0])
      2'b0, 2'b01:
	  CASE_fpu_sqr_fState_S4D_OUT_BITS_1_TO_0_0b0_f_ETC__q21 =
	      fpu_sqr_fState_S4$D_OUT[64:54];
      2'b10:
	  CASE_fpu_sqr_fState_S4D_OUT_BITS_1_TO_0_0b0_f_ETC__q21 =
	      out_exp__h95912;
      2'b11:
	  CASE_fpu_sqr_fState_S4D_OUT_BITS_1_TO_0_0b0_f_ETC__q21 =
	      _theResult___exp__h95909;
    endcase
  end
  always@(fpu_sqr_fState_S4$D_OUT or _theResult___exp__h95909)
  begin
    case (fpu_sqr_fState_S4$D_OUT[1:0])
      2'b0:
	  CASE_fpu_sqr_fState_S4D_OUT_BITS_1_TO_0_0b0_f_ETC__q22 =
	      fpu_sqr_fState_S4$D_OUT[64:54];
      2'b01, 2'b10, 2'b11:
	  CASE_fpu_sqr_fState_S4D_OUT_BITS_1_TO_0_0b0_f_ETC__q22 =
	      _theResult___exp__h95909;
    endcase
  end
  always@(fpu_sqr_fState_S4$D_OUT or
	  CASE_fpu_sqr_fState_S4D_OUT_BITS_1_TO_0_0b0_f_ETC__q21 or
	  CASE_fpu_sqr_fState_S4D_OUT_BITS_1_TO_0_0b0_f_ETC__q22 or
	  _theResult___exp__h95909)
  begin
    case (fpu_sqr_fState_S4$D_OUT[68:66])
      3'd0:
	  _theResult___fst_exp__h95987 =
	      CASE_fpu_sqr_fState_S4D_OUT_BITS_1_TO_0_0b0_f_ETC__q21;
      3'd1:
	  _theResult___fst_exp__h95987 =
	      CASE_fpu_sqr_fState_S4D_OUT_BITS_1_TO_0_0b0_f_ETC__q22;
      3'd2:
	  _theResult___fst_exp__h95987 =
	      (fpu_sqr_fState_S4$D_OUT[1:0] == 2'b0 ||
	       fpu_sqr_fState_S4$D_OUT[65]) ?
		fpu_sqr_fState_S4$D_OUT[64:54] :
		_theResult___exp__h95909;
      3'd3:
	  _theResult___fst_exp__h95987 =
	      (fpu_sqr_fState_S4$D_OUT[1:0] == 2'b0) ?
		fpu_sqr_fState_S4$D_OUT[64:54] :
		(fpu_sqr_fState_S4$D_OUT[65] ?
		   _theResult___exp__h95909 :
		   fpu_sqr_fState_S4$D_OUT[64:54]);
      3'd4: _theResult___fst_exp__h95987 = fpu_sqr_fState_S4$D_OUT[64:54];
      default: _theResult___fst_exp__h95987 = 11'd0;
    endcase
  end
  always@(fpu_madd_fState_S8$D_OUT or
	  out_exp__h142544 or _theResult___exp__h142541)
  begin
    case (fpu_madd_fState_S8$D_OUT[2:1])
      2'b0, 2'b01:
	  CASE_fpu_madd_fState_S8D_OUT_BITS_2_TO_1_0b0__ETC__q31 =
	      fpu_madd_fState_S8$D_OUT[65:55];
      2'b10:
	  CASE_fpu_madd_fState_S8D_OUT_BITS_2_TO_1_0b0__ETC__q31 =
	      out_exp__h142544;
      2'b11:
	  CASE_fpu_madd_fState_S8D_OUT_BITS_2_TO_1_0b0__ETC__q31 =
	      _theResult___exp__h142541;
    endcase
  end
  always@(fpu_madd_fState_S8$D_OUT or _theResult___exp__h142541)
  begin
    case (fpu_madd_fState_S8$D_OUT[2:1])
      2'b0:
	  CASE_fpu_madd_fState_S8D_OUT_BITS_2_TO_1_0b0__ETC__q32 =
	      fpu_madd_fState_S8$D_OUT[65:55];
      2'b01, 2'b10, 2'b11:
	  CASE_fpu_madd_fState_S8D_OUT_BITS_2_TO_1_0b0__ETC__q32 =
	      _theResult___exp__h142541;
    endcase
  end
  always@(fpu_madd_fState_S8$D_OUT or
	  CASE_fpu_madd_fState_S8D_OUT_BITS_2_TO_1_0b0__ETC__q31 or
	  CASE_fpu_madd_fState_S8D_OUT_BITS_2_TO_1_0b0__ETC__q32 or
	  _theResult___exp__h142541)
  begin
    case (fpu_madd_fState_S8$D_OUT[70:68])
      3'd0:
	  _theResult___fst_exp__h142619 =
	      CASE_fpu_madd_fState_S8D_OUT_BITS_2_TO_1_0b0__ETC__q31;
      3'd1:
	  _theResult___fst_exp__h142619 =
	      CASE_fpu_madd_fState_S8D_OUT_BITS_2_TO_1_0b0__ETC__q32;
      3'd2:
	  _theResult___fst_exp__h142619 =
	      (fpu_madd_fState_S8$D_OUT[2:1] == 2'b0 ||
	       fpu_madd_fState_S8$D_OUT[66]) ?
		fpu_madd_fState_S8$D_OUT[65:55] :
		_theResult___exp__h142541;
      3'd3:
	  _theResult___fst_exp__h142619 =
	      (fpu_madd_fState_S8$D_OUT[2:1] == 2'b0) ?
		fpu_madd_fState_S8$D_OUT[65:55] :
		(fpu_madd_fState_S8$D_OUT[66] ?
		   _theResult___exp__h142541 :
		   fpu_madd_fState_S8$D_OUT[65:55]);
      3'd4: _theResult___fst_exp__h142619 = fpu_madd_fState_S8$D_OUT[65:55];
      default: _theResult___fst_exp__h142619 = 11'd0;
    endcase
  end
  always@(guard__h155373 or
	  _theResult___fst_exp__h163334 or
	  out_exp__h163982 or _theResult___exp__h163979)
  begin
    case (guard__h155373)
      2'b0, 2'b01:
	  CASE_guard55373_0b0_theResult___fst_exp63334_0_ETC__q42 =
	      _theResult___fst_exp__h163334;
      2'b10:
	  CASE_guard55373_0b0_theResult___fst_exp63334_0_ETC__q42 =
	      out_exp__h163982;
      2'b11:
	  CASE_guard55373_0b0_theResult___fst_exp63334_0_ETC__q42 =
	      _theResult___exp__h163979;
    endcase
  end
  always@(guard__h155373 or
	  _theResult___fst_exp__h163334 or _theResult___exp__h163979)
  begin
    case (guard__h155373)
      2'b0:
	  CASE_guard55373_0b0_theResult___fst_exp63334_0_ETC__q43 =
	      _theResult___fst_exp__h163334;
      2'b01, 2'b10, 2'b11:
	  CASE_guard55373_0b0_theResult___fst_exp63334_0_ETC__q43 =
	      _theResult___exp__h163979;
    endcase
  end
  always@(iFifo$D_OUT or
	  CASE_guard55373_0b0_theResult___fst_exp63334_0_ETC__q42 or
	  CASE_guard55373_0b0_theResult___fst_exp63334_0_ETC__q43 or
	  IF_IF_IF_iFifo_first__087_BITS_167_TO_160_130__ETC___d3690 or
	  IF_IF_IF_iFifo_first__087_BITS_167_TO_160_130__ETC___d3692 or
	  _theResult___fst_exp__h163334)
  begin
    case (iFifo$D_OUT[6:4])
      3'd0:
	  _theResult___fst_exp__h164057 =
	      CASE_guard55373_0b0_theResult___fst_exp63334_0_ETC__q42;
      3'd1:
	  _theResult___fst_exp__h164057 =
	      CASE_guard55373_0b0_theResult___fst_exp63334_0_ETC__q43;
      3'd2:
	  _theResult___fst_exp__h164057 =
	      IF_IF_IF_iFifo_first__087_BITS_167_TO_160_130__ETC___d3690;
      3'd3:
	  _theResult___fst_exp__h164057 =
	      IF_IF_IF_iFifo_first__087_BITS_167_TO_160_130__ETC___d3692;
      3'd4: _theResult___fst_exp__h164057 = _theResult___fst_exp__h163334;
      default: _theResult___fst_exp__h164057 = 11'd0;
    endcase
  end
  always@(guard__h164622 or
	  _theResult___fst_exp__h172850 or
	  out_exp__h173572 or _theResult___exp__h173569)
  begin
    case (guard__h164622)
      2'b0, 2'b01:
	  CASE_guard64622_0b0_theResult___fst_exp72850_0_ETC__q44 =
	      _theResult___fst_exp__h172850;
      2'b10:
	  CASE_guard64622_0b0_theResult___fst_exp72850_0_ETC__q44 =
	      out_exp__h173572;
      2'b11:
	  CASE_guard64622_0b0_theResult___fst_exp72850_0_ETC__q44 =
	      _theResult___exp__h173569;
    endcase
  end
  always@(guard__h164622 or
	  _theResult___fst_exp__h172850 or _theResult___exp__h173569)
  begin
    case (guard__h164622)
      2'b0:
	  CASE_guard64622_0b0_theResult___fst_exp72850_0_ETC__q45 =
	      _theResult___fst_exp__h172850;
      2'b01, 2'b10, 2'b11:
	  CASE_guard64622_0b0_theResult___fst_exp72850_0_ETC__q45 =
	      _theResult___exp__h173569;
    endcase
  end
  always@(iFifo$D_OUT or
	  CASE_guard64622_0b0_theResult___fst_exp72850_0_ETC__q44 or
	  CASE_guard64622_0b0_theResult___fst_exp72850_0_ETC__q45 or
	  IF_IF_IF_IF_3074_MINUS_SEXT_iFifo_first__087_B_ETC___d3729 or
	  IF_IF_IF_IF_3074_MINUS_SEXT_iFifo_first__087_B_ETC___d3731 or
	  _theResult___fst_exp__h172850)
  begin
    case (iFifo$D_OUT[6:4])
      3'd0:
	  _theResult___fst_exp__h173647 =
	      CASE_guard64622_0b0_theResult___fst_exp72850_0_ETC__q44;
      3'd1:
	  _theResult___fst_exp__h173647 =
	      CASE_guard64622_0b0_theResult___fst_exp72850_0_ETC__q45;
      3'd2:
	  _theResult___fst_exp__h173647 =
	      IF_IF_IF_IF_3074_MINUS_SEXT_iFifo_first__087_B_ETC___d3729;
      3'd3:
	  _theResult___fst_exp__h173647 =
	      IF_IF_IF_IF_3074_MINUS_SEXT_iFifo_first__087_B_ETC___d3731;
      3'd4: _theResult___fst_exp__h173647 = _theResult___fst_exp__h172850;
      default: _theResult___fst_exp__h173647 = 11'd0;
    endcase
  end
  always@(guard__h173661 or
	  _theResult___fst_exp__h181651 or
	  out_exp__h182324 or _theResult___exp__h182321)
  begin
    case (guard__h173661)
      2'b0, 2'b01:
	  CASE_guard73661_0b0_theResult___fst_exp81651_0_ETC__q46 =
	      _theResult___fst_exp__h181651;
      2'b10:
	  CASE_guard73661_0b0_theResult___fst_exp81651_0_ETC__q46 =
	      out_exp__h182324;
      2'b11:
	  CASE_guard73661_0b0_theResult___fst_exp81651_0_ETC__q46 =
	      _theResult___exp__h182321;
    endcase
  end
  always@(guard__h173661 or
	  _theResult___fst_exp__h181651 or _theResult___exp__h182321)
  begin
    case (guard__h173661)
      2'b0:
	  CASE_guard73661_0b0_theResult___fst_exp81651_0_ETC__q47 =
	      _theResult___fst_exp__h181651;
      2'b01, 2'b10, 2'b11:
	  CASE_guard73661_0b0_theResult___fst_exp81651_0_ETC__q47 =
	      _theResult___exp__h182321;
    endcase
  end
  always@(iFifo$D_OUT or
	  CASE_guard73661_0b0_theResult___fst_exp81651_0_ETC__q46 or
	  CASE_guard73661_0b0_theResult___fst_exp81651_0_ETC__q47 or
	  IF_IF_IF_iFifo_first__087_BITS_167_TO_160_130__ETC___d3760 or
	  IF_IF_IF_iFifo_first__087_BITS_167_TO_160_130__ETC___d3762 or
	  _theResult___fst_exp__h181651)
  begin
    case (iFifo$D_OUT[6:4])
      3'd0:
	  _theResult___fst_exp__h182399 =
	      CASE_guard73661_0b0_theResult___fst_exp81651_0_ETC__q46;
      3'd1:
	  _theResult___fst_exp__h182399 =
	      CASE_guard73661_0b0_theResult___fst_exp81651_0_ETC__q47;
      3'd2:
	  _theResult___fst_exp__h182399 =
	      IF_IF_IF_iFifo_first__087_BITS_167_TO_160_130__ETC___d3760;
      3'd3:
	  _theResult___fst_exp__h182399 =
	      IF_IF_IF_iFifo_first__087_BITS_167_TO_160_130__ETC___d3762;
      3'd4: _theResult___fst_exp__h182399 = _theResult___fst_exp__h181651;
      default: _theResult___fst_exp__h182399 = 11'd0;
    endcase
  end
  always@(guard__h155373 or
	  _theResult___snd__h163285 or
	  out_sfd__h163983 or _theResult___sfd__h163980)
  begin
    case (guard__h155373)
      2'b0, 2'b01:
	  CASE_guard55373_0b0_theResult___snd63285_BITS__ETC__q48 =
	      _theResult___snd__h163285[56:5];
      2'b10:
	  CASE_guard55373_0b0_theResult___snd63285_BITS__ETC__q48 =
	      out_sfd__h163983;
      2'b11:
	  CASE_guard55373_0b0_theResult___snd63285_BITS__ETC__q48 =
	      _theResult___sfd__h163980;
    endcase
  end
  always@(guard__h155373 or
	  _theResult___snd__h163285 or _theResult___sfd__h163980)
  begin
    case (guard__h155373)
      2'b0:
	  CASE_guard55373_0b0_theResult___snd63285_BITS__ETC__q49 =
	      _theResult___snd__h163285[56:5];
      2'b01, 2'b10, 2'b11:
	  CASE_guard55373_0b0_theResult___snd63285_BITS__ETC__q49 =
	      _theResult___sfd__h163980;
    endcase
  end
  always@(iFifo$D_OUT or
	  CASE_guard55373_0b0_theResult___snd63285_BITS__ETC__q48 or
	  CASE_guard55373_0b0_theResult___snd63285_BITS__ETC__q49 or
	  IF_IF_IF_iFifo_first__087_BITS_167_TO_160_130__ETC___d3786 or
	  IF_IF_IF_iFifo_first__087_BITS_167_TO_160_130__ETC___d3788 or
	  _theResult___snd__h163285)
  begin
    case (iFifo$D_OUT[6:4])
      3'd0:
	  _theResult___fst_sfd__h164058 =
	      CASE_guard55373_0b0_theResult___snd63285_BITS__ETC__q48;
      3'd1:
	  _theResult___fst_sfd__h164058 =
	      CASE_guard55373_0b0_theResult___snd63285_BITS__ETC__q49;
      3'd2:
	  _theResult___fst_sfd__h164058 =
	      IF_IF_IF_iFifo_first__087_BITS_167_TO_160_130__ETC___d3786;
      3'd3:
	  _theResult___fst_sfd__h164058 =
	      IF_IF_IF_iFifo_first__087_BITS_167_TO_160_130__ETC___d3788;
      3'd4: _theResult___fst_sfd__h164058 = _theResult___snd__h163285[56:5];
      default: _theResult___fst_sfd__h164058 = 52'd0;
    endcase
  end
  always@(guard__h164622 or
	  sfdin__h172844 or out_sfd__h173573 or _theResult___sfd__h173570)
  begin
    case (guard__h164622)
      2'b0, 2'b01:
	  CASE_guard64622_0b0_sfdin72844_BITS_56_TO_5_0b_ETC__q50 =
	      sfdin__h172844[56:5];
      2'b10:
	  CASE_guard64622_0b0_sfdin72844_BITS_56_TO_5_0b_ETC__q50 =
	      out_sfd__h173573;
      2'b11:
	  CASE_guard64622_0b0_sfdin72844_BITS_56_TO_5_0b_ETC__q50 =
	      _theResult___sfd__h173570;
    endcase
  end
  always@(guard__h164622 or sfdin__h172844 or _theResult___sfd__h173570)
  begin
    case (guard__h164622)
      2'b0:
	  CASE_guard64622_0b0_sfdin72844_BITS_56_TO_5_0b_ETC__q51 =
	      sfdin__h172844[56:5];
      2'b01, 2'b10, 2'b11:
	  CASE_guard64622_0b0_sfdin72844_BITS_56_TO_5_0b_ETC__q51 =
	      _theResult___sfd__h173570;
    endcase
  end
  always@(iFifo$D_OUT or
	  CASE_guard64622_0b0_sfdin72844_BITS_56_TO_5_0b_ETC__q50 or
	  CASE_guard64622_0b0_sfdin72844_BITS_56_TO_5_0b_ETC__q51 or
	  IF_IF_IF_IF_3074_MINUS_SEXT_iFifo_first__087_B_ETC___d3813 or
	  IF_IF_IF_IF_3074_MINUS_SEXT_iFifo_first__087_B_ETC___d3815 or
	  sfdin__h172844)
  begin
    case (iFifo$D_OUT[6:4])
      3'd0:
	  _theResult___fst_sfd__h173648 =
	      CASE_guard64622_0b0_sfdin72844_BITS_56_TO_5_0b_ETC__q50;
      3'd1:
	  _theResult___fst_sfd__h173648 =
	      CASE_guard64622_0b0_sfdin72844_BITS_56_TO_5_0b_ETC__q51;
      3'd2:
	  _theResult___fst_sfd__h173648 =
	      IF_IF_IF_IF_3074_MINUS_SEXT_iFifo_first__087_B_ETC___d3813;
      3'd3:
	  _theResult___fst_sfd__h173648 =
	      IF_IF_IF_IF_3074_MINUS_SEXT_iFifo_first__087_B_ETC___d3815;
      3'd4: _theResult___fst_sfd__h173648 = sfdin__h172844[56:5];
      default: _theResult___fst_sfd__h173648 = 52'd0;
    endcase
  end
  always@(guard__h173661 or
	  _theResult___snd__h181597 or
	  out_sfd__h182325 or _theResult___sfd__h182322)
  begin
    case (guard__h173661)
      2'b0, 2'b01:
	  CASE_guard73661_0b0_theResult___snd81597_BITS__ETC__q52 =
	      _theResult___snd__h181597[56:5];
      2'b10:
	  CASE_guard73661_0b0_theResult___snd81597_BITS__ETC__q52 =
	      out_sfd__h182325;
      2'b11:
	  CASE_guard73661_0b0_theResult___snd81597_BITS__ETC__q52 =
	      _theResult___sfd__h182322;
    endcase
  end
  always@(guard__h173661 or
	  _theResult___snd__h181597 or _theResult___sfd__h182322)
  begin
    case (guard__h173661)
      2'b0:
	  CASE_guard73661_0b0_theResult___snd81597_BITS__ETC__q53 =
	      _theResult___snd__h181597[56:5];
      2'b01, 2'b10, 2'b11:
	  CASE_guard73661_0b0_theResult___snd81597_BITS__ETC__q53 =
	      _theResult___sfd__h182322;
    endcase
  end
  always@(iFifo$D_OUT or
	  CASE_guard73661_0b0_theResult___snd81597_BITS__ETC__q52 or
	  CASE_guard73661_0b0_theResult___snd81597_BITS__ETC__q53 or
	  IF_IF_IF_iFifo_first__087_BITS_167_TO_160_130__ETC___d3832 or
	  IF_IF_IF_iFifo_first__087_BITS_167_TO_160_130__ETC___d3834 or
	  _theResult___snd__h181597)
  begin
    case (iFifo$D_OUT[6:4])
      3'd0:
	  _theResult___fst_sfd__h182400 =
	      CASE_guard73661_0b0_theResult___snd81597_BITS__ETC__q52;
      3'd1:
	  _theResult___fst_sfd__h182400 =
	      CASE_guard73661_0b0_theResult___snd81597_BITS__ETC__q53;
      3'd2:
	  _theResult___fst_sfd__h182400 =
	      IF_IF_IF_iFifo_first__087_BITS_167_TO_160_130__ETC___d3832;
      3'd3:
	  _theResult___fst_sfd__h182400 =
	      IF_IF_IF_iFifo_first__087_BITS_167_TO_160_130__ETC___d3834;
      3'd4: _theResult___fst_sfd__h182400 = _theResult___snd__h181597[56:5];
      default: _theResult___fst_sfd__h182400 = 52'd0;
    endcase
  end
  always@(guard__h155373 or iFifo$D_OUT)
  begin
    case (guard__h155373)
      2'b0, 2'b01, 2'b10:
	  CASE_guard55373_0b0_iFifoD_OUT_BIT_168_0b1_iF_ETC__q54 =
	      iFifo$D_OUT[168];
      2'd3:
	  CASE_guard55373_0b0_iFifoD_OUT_BIT_168_0b1_iF_ETC__q54 =
	      guard__h155373 == 2'b11 && iFifo$D_OUT[168];
    endcase
  end
  always@(iFifo$D_OUT or
	  CASE_guard55373_0b0_iFifoD_OUT_BIT_168_0b1_iF_ETC__q54 or
	  guard__h155373)
  begin
    case (iFifo$D_OUT[6:4])
      3'd0:
	  CASE_iFifoD_OUT_BITS_6_TO_4_0_CASE_guard55373_ETC__q55 =
	      CASE_guard55373_0b0_iFifoD_OUT_BIT_168_0b1_iF_ETC__q54;
      3'd1:
	  CASE_iFifoD_OUT_BITS_6_TO_4_0_CASE_guard55373_ETC__q55 =
	      (guard__h155373 == 2'b0) ?
		iFifo$D_OUT[168] :
		(guard__h155373 == 2'b01 || guard__h155373 == 2'b10 ||
		 guard__h155373 == 2'b11) &&
		iFifo$D_OUT[168];
      3'd2, 3'd3:
	  CASE_iFifoD_OUT_BITS_6_TO_4_0_CASE_guard55373_ETC__q55 =
	      iFifo$D_OUT[168];
      default: CASE_iFifoD_OUT_BITS_6_TO_4_0_CASE_guard55373_ETC__q55 =
		   iFifo$D_OUT[6:4] == 3'd4 && iFifo$D_OUT[168];
    endcase
  end
  always@(iFifo$D_OUT)
  begin
    case (iFifo$D_OUT[6:4])
      3'd0, 3'd1, 3'd2, 3'd3:
	  IF_iFifo_first__087_BITS_6_TO_4_118_EQ_0_191_O_ETC___d3320 =
	      iFifo$D_OUT[168];
      default: IF_iFifo_first__087_BITS_6_TO_4_118_EQ_0_191_O_ETC___d3320 =
		   iFifo$D_OUT[6:4] == 3'd4 && iFifo$D_OUT[168];
    endcase
  end
  always@(guard__h164622 or iFifo$D_OUT)
  begin
    case (guard__h164622)
      2'b0, 2'b01, 2'b10:
	  CASE_guard64622_0b0_iFifoD_OUT_BIT_168_0b1_iF_ETC__q56 =
	      iFifo$D_OUT[168];
      2'd3:
	  CASE_guard64622_0b0_iFifoD_OUT_BIT_168_0b1_iF_ETC__q56 =
	      guard__h164622 == 2'b11 && iFifo$D_OUT[168];
    endcase
  end
  always@(iFifo$D_OUT or
	  CASE_guard64622_0b0_iFifoD_OUT_BIT_168_0b1_iF_ETC__q56 or
	  guard__h164622)
  begin
    case (iFifo$D_OUT[6:4])
      3'd0:
	  CASE_iFifoD_OUT_BITS_6_TO_4_0_CASE_guard64622_ETC__q57 =
	      CASE_guard64622_0b0_iFifoD_OUT_BIT_168_0b1_iF_ETC__q56;
      3'd1:
	  CASE_iFifoD_OUT_BITS_6_TO_4_0_CASE_guard64622_ETC__q57 =
	      (guard__h164622 == 2'b0) ?
		iFifo$D_OUT[168] :
		(guard__h164622 == 2'b01 || guard__h164622 == 2'b10 ||
		 guard__h164622 == 2'b11) &&
		iFifo$D_OUT[168];
      3'd2, 3'd3:
	  CASE_iFifoD_OUT_BITS_6_TO_4_0_CASE_guard64622_ETC__q57 =
	      iFifo$D_OUT[168];
      default: CASE_iFifoD_OUT_BITS_6_TO_4_0_CASE_guard64622_ETC__q57 =
		   iFifo$D_OUT[6:4] == 3'd4 && iFifo$D_OUT[168];
    endcase
  end
  always@(guard__h173661 or iFifo$D_OUT)
  begin
    case (guard__h173661)
      2'b0, 2'b01, 2'b10:
	  CASE_guard73661_0b0_iFifoD_OUT_BIT_168_0b1_iF_ETC__q58 =
	      iFifo$D_OUT[168];
      2'd3:
	  CASE_guard73661_0b0_iFifoD_OUT_BIT_168_0b1_iF_ETC__q58 =
	      guard__h173661 == 2'b11 && iFifo$D_OUT[168];
    endcase
  end
  always@(iFifo$D_OUT or
	  CASE_guard73661_0b0_iFifoD_OUT_BIT_168_0b1_iF_ETC__q58 or
	  guard__h173661)
  begin
    case (iFifo$D_OUT[6:4])
      3'd0:
	  CASE_iFifoD_OUT_BITS_6_TO_4_0_CASE_guard73661_ETC__q59 =
	      CASE_guard73661_0b0_iFifoD_OUT_BIT_168_0b1_iF_ETC__q58;
      3'd1:
	  CASE_iFifoD_OUT_BITS_6_TO_4_0_CASE_guard73661_ETC__q59 =
	      (guard__h173661 == 2'b0) ?
		iFifo$D_OUT[168] :
		(guard__h173661 == 2'b01 || guard__h173661 == 2'b10 ||
		 guard__h173661 == 2'b11) &&
		iFifo$D_OUT[168];
      3'd2, 3'd3:
	  CASE_iFifoD_OUT_BITS_6_TO_4_0_CASE_guard73661_ETC__q59 =
	      iFifo$D_OUT[168];
      default: CASE_iFifoD_OUT_BITS_6_TO_4_0_CASE_guard73661_ETC__q59 =
		   iFifo$D_OUT[6:4] == 3'd4 && iFifo$D_OUT[168];
    endcase
  end
  always@(guard__h232950 or
	  _theResult___fst_exp__h240911 or
	  out_exp__h241559 or _theResult___exp__h241556)
  begin
    case (guard__h232950)
      2'b0, 2'b01:
	  CASE_guard32950_0b0_theResult___fst_exp40911_0_ETC__q69 =
	      _theResult___fst_exp__h240911;
      2'b10:
	  CASE_guard32950_0b0_theResult___fst_exp40911_0_ETC__q69 =
	      out_exp__h241559;
      2'b11:
	  CASE_guard32950_0b0_theResult___fst_exp40911_0_ETC__q69 =
	      _theResult___exp__h241556;
    endcase
  end
  always@(guard__h232950 or
	  _theResult___fst_exp__h240911 or _theResult___exp__h241556)
  begin
    case (guard__h232950)
      2'b0:
	  CASE_guard32950_0b0_theResult___fst_exp40911_0_ETC__q70 =
	      _theResult___fst_exp__h240911;
      2'b01, 2'b10, 2'b11:
	  CASE_guard32950_0b0_theResult___fst_exp40911_0_ETC__q70 =
	      _theResult___exp__h241556;
    endcase
  end
  always@(iFifo$D_OUT or
	  CASE_guard32950_0b0_theResult___fst_exp40911_0_ETC__q69 or
	  CASE_guard32950_0b0_theResult___fst_exp40911_0_ETC__q70 or
	  IF_IF_IF_iFifo_first__087_BITS_37_TO_30_850_EQ_ETC___d4398 or
	  IF_IF_IF_iFifo_first__087_BITS_37_TO_30_850_EQ_ETC___d4400 or
	  _theResult___fst_exp__h240911)
  begin
    case (iFifo$D_OUT[6:4])
      3'd0:
	  _theResult___fst_exp__h241634 =
	      CASE_guard32950_0b0_theResult___fst_exp40911_0_ETC__q69;
      3'd1:
	  _theResult___fst_exp__h241634 =
	      CASE_guard32950_0b0_theResult___fst_exp40911_0_ETC__q70;
      3'd2:
	  _theResult___fst_exp__h241634 =
	      IF_IF_IF_iFifo_first__087_BITS_37_TO_30_850_EQ_ETC___d4398;
      3'd3:
	  _theResult___fst_exp__h241634 =
	      IF_IF_IF_iFifo_first__087_BITS_37_TO_30_850_EQ_ETC___d4400;
      3'd4: _theResult___fst_exp__h241634 = _theResult___fst_exp__h240911;
      default: _theResult___fst_exp__h241634 = 11'd0;
    endcase
  end
  always@(guard__h242199 or
	  _theResult___fst_exp__h250427 or
	  out_exp__h251149 or _theResult___exp__h251146)
  begin
    case (guard__h242199)
      2'b0, 2'b01:
	  CASE_guard42199_0b0_theResult___fst_exp50427_0_ETC__q71 =
	      _theResult___fst_exp__h250427;
      2'b10:
	  CASE_guard42199_0b0_theResult___fst_exp50427_0_ETC__q71 =
	      out_exp__h251149;
      2'b11:
	  CASE_guard42199_0b0_theResult___fst_exp50427_0_ETC__q71 =
	      _theResult___exp__h251146;
    endcase
  end
  always@(guard__h242199 or
	  _theResult___fst_exp__h250427 or _theResult___exp__h251146)
  begin
    case (guard__h242199)
      2'b0:
	  CASE_guard42199_0b0_theResult___fst_exp50427_0_ETC__q72 =
	      _theResult___fst_exp__h250427;
      2'b01, 2'b10, 2'b11:
	  CASE_guard42199_0b0_theResult___fst_exp50427_0_ETC__q72 =
	      _theResult___exp__h251146;
    endcase
  end
  always@(iFifo$D_OUT or
	  CASE_guard42199_0b0_theResult___fst_exp50427_0_ETC__q71 or
	  CASE_guard42199_0b0_theResult___fst_exp50427_0_ETC__q72 or
	  IF_IF_IF_IF_3074_MINUS_SEXT_iFifo_first__087_B_ETC___d4436 or
	  IF_IF_IF_IF_3074_MINUS_SEXT_iFifo_first__087_B_ETC___d4438 or
	  _theResult___fst_exp__h250427)
  begin
    case (iFifo$D_OUT[6:4])
      3'd0:
	  _theResult___fst_exp__h251224 =
	      CASE_guard42199_0b0_theResult___fst_exp50427_0_ETC__q71;
      3'd1:
	  _theResult___fst_exp__h251224 =
	      CASE_guard42199_0b0_theResult___fst_exp50427_0_ETC__q72;
      3'd2:
	  _theResult___fst_exp__h251224 =
	      IF_IF_IF_IF_3074_MINUS_SEXT_iFifo_first__087_B_ETC___d4436;
      3'd3:
	  _theResult___fst_exp__h251224 =
	      IF_IF_IF_IF_3074_MINUS_SEXT_iFifo_first__087_B_ETC___d4438;
      3'd4: _theResult___fst_exp__h251224 = _theResult___fst_exp__h250427;
      default: _theResult___fst_exp__h251224 = 11'd0;
    endcase
  end
  always@(guard__h251238 or
	  _theResult___fst_exp__h259228 or
	  out_exp__h259901 or _theResult___exp__h259898)
  begin
    case (guard__h251238)
      2'b0, 2'b01:
	  CASE_guard51238_0b0_theResult___fst_exp59228_0_ETC__q73 =
	      _theResult___fst_exp__h259228;
      2'b10:
	  CASE_guard51238_0b0_theResult___fst_exp59228_0_ETC__q73 =
	      out_exp__h259901;
      2'b11:
	  CASE_guard51238_0b0_theResult___fst_exp59228_0_ETC__q73 =
	      _theResult___exp__h259898;
    endcase
  end
  always@(guard__h251238 or
	  _theResult___fst_exp__h259228 or _theResult___exp__h259898)
  begin
    case (guard__h251238)
      2'b0:
	  CASE_guard51238_0b0_theResult___fst_exp59228_0_ETC__q74 =
	      _theResult___fst_exp__h259228;
      2'b01, 2'b10, 2'b11:
	  CASE_guard51238_0b0_theResult___fst_exp59228_0_ETC__q74 =
	      _theResult___exp__h259898;
    endcase
  end
  always@(iFifo$D_OUT or
	  CASE_guard51238_0b0_theResult___fst_exp59228_0_ETC__q73 or
	  CASE_guard51238_0b0_theResult___fst_exp59228_0_ETC__q74 or
	  IF_IF_IF_iFifo_first__087_BITS_37_TO_30_850_EQ_ETC___d4467 or
	  IF_IF_IF_iFifo_first__087_BITS_37_TO_30_850_EQ_ETC___d4469 or
	  _theResult___fst_exp__h259228)
  begin
    case (iFifo$D_OUT[6:4])
      3'd0:
	  _theResult___fst_exp__h259976 =
	      CASE_guard51238_0b0_theResult___fst_exp59228_0_ETC__q73;
      3'd1:
	  _theResult___fst_exp__h259976 =
	      CASE_guard51238_0b0_theResult___fst_exp59228_0_ETC__q74;
      3'd2:
	  _theResult___fst_exp__h259976 =
	      IF_IF_IF_iFifo_first__087_BITS_37_TO_30_850_EQ_ETC___d4467;
      3'd3:
	  _theResult___fst_exp__h259976 =
	      IF_IF_IF_iFifo_first__087_BITS_37_TO_30_850_EQ_ETC___d4469;
      3'd4: _theResult___fst_exp__h259976 = _theResult___fst_exp__h259228;
      default: _theResult___fst_exp__h259976 = 11'd0;
    endcase
  end
  always@(guard__h232950 or
	  _theResult___snd__h240862 or
	  out_sfd__h241560 or _theResult___sfd__h241557)
  begin
    case (guard__h232950)
      2'b0, 2'b01:
	  CASE_guard32950_0b0_theResult___snd40862_BITS__ETC__q75 =
	      _theResult___snd__h240862[56:5];
      2'b10:
	  CASE_guard32950_0b0_theResult___snd40862_BITS__ETC__q75 =
	      out_sfd__h241560;
      2'b11:
	  CASE_guard32950_0b0_theResult___snd40862_BITS__ETC__q75 =
	      _theResult___sfd__h241557;
    endcase
  end
  always@(guard__h232950 or
	  _theResult___snd__h240862 or _theResult___sfd__h241557)
  begin
    case (guard__h232950)
      2'b0:
	  CASE_guard32950_0b0_theResult___snd40862_BITS__ETC__q76 =
	      _theResult___snd__h240862[56:5];
      2'b01, 2'b10, 2'b11:
	  CASE_guard32950_0b0_theResult___snd40862_BITS__ETC__q76 =
	      _theResult___sfd__h241557;
    endcase
  end
  always@(iFifo$D_OUT or
	  CASE_guard32950_0b0_theResult___snd40862_BITS__ETC__q75 or
	  CASE_guard32950_0b0_theResult___snd40862_BITS__ETC__q76 or
	  IF_IF_IF_iFifo_first__087_BITS_37_TO_30_850_EQ_ETC___d4493 or
	  IF_IF_IF_iFifo_first__087_BITS_37_TO_30_850_EQ_ETC___d4495 or
	  _theResult___snd__h240862)
  begin
    case (iFifo$D_OUT[6:4])
      3'd0:
	  _theResult___fst_sfd__h241635 =
	      CASE_guard32950_0b0_theResult___snd40862_BITS__ETC__q75;
      3'd1:
	  _theResult___fst_sfd__h241635 =
	      CASE_guard32950_0b0_theResult___snd40862_BITS__ETC__q76;
      3'd2:
	  _theResult___fst_sfd__h241635 =
	      IF_IF_IF_iFifo_first__087_BITS_37_TO_30_850_EQ_ETC___d4493;
      3'd3:
	  _theResult___fst_sfd__h241635 =
	      IF_IF_IF_iFifo_first__087_BITS_37_TO_30_850_EQ_ETC___d4495;
      3'd4: _theResult___fst_sfd__h241635 = _theResult___snd__h240862[56:5];
      default: _theResult___fst_sfd__h241635 = 52'd0;
    endcase
  end
  always@(guard__h242199 or
	  sfdin__h250421 or out_sfd__h251150 or _theResult___sfd__h251147)
  begin
    case (guard__h242199)
      2'b0, 2'b01:
	  CASE_guard42199_0b0_sfdin50421_BITS_56_TO_5_0b_ETC__q77 =
	      sfdin__h250421[56:5];
      2'b10:
	  CASE_guard42199_0b0_sfdin50421_BITS_56_TO_5_0b_ETC__q77 =
	      out_sfd__h251150;
      2'b11:
	  CASE_guard42199_0b0_sfdin50421_BITS_56_TO_5_0b_ETC__q77 =
	      _theResult___sfd__h251147;
    endcase
  end
  always@(guard__h242199 or sfdin__h250421 or _theResult___sfd__h251147)
  begin
    case (guard__h242199)
      2'b0:
	  CASE_guard42199_0b0_sfdin50421_BITS_56_TO_5_0b_ETC__q78 =
	      sfdin__h250421[56:5];
      2'b01, 2'b10, 2'b11:
	  CASE_guard42199_0b0_sfdin50421_BITS_56_TO_5_0b_ETC__q78 =
	      _theResult___sfd__h251147;
    endcase
  end
  always@(iFifo$D_OUT or
	  CASE_guard42199_0b0_sfdin50421_BITS_56_TO_5_0b_ETC__q77 or
	  CASE_guard42199_0b0_sfdin50421_BITS_56_TO_5_0b_ETC__q78 or
	  IF_IF_IF_IF_3074_MINUS_SEXT_iFifo_first__087_B_ETC___d4519 or
	  IF_IF_IF_IF_3074_MINUS_SEXT_iFifo_first__087_B_ETC___d4521 or
	  sfdin__h250421)
  begin
    case (iFifo$D_OUT[6:4])
      3'd0:
	  _theResult___fst_sfd__h251225 =
	      CASE_guard42199_0b0_sfdin50421_BITS_56_TO_5_0b_ETC__q77;
      3'd1:
	  _theResult___fst_sfd__h251225 =
	      CASE_guard42199_0b0_sfdin50421_BITS_56_TO_5_0b_ETC__q78;
      3'd2:
	  _theResult___fst_sfd__h251225 =
	      IF_IF_IF_IF_3074_MINUS_SEXT_iFifo_first__087_B_ETC___d4519;
      3'd3:
	  _theResult___fst_sfd__h251225 =
	      IF_IF_IF_IF_3074_MINUS_SEXT_iFifo_first__087_B_ETC___d4521;
      3'd4: _theResult___fst_sfd__h251225 = sfdin__h250421[56:5];
      default: _theResult___fst_sfd__h251225 = 52'd0;
    endcase
  end
  always@(guard__h232950 or iFifo$D_OUT)
  begin
    case (guard__h232950)
      2'b0, 2'b01, 2'b10:
	  CASE_guard32950_0b0_iFifoD_OUT_BIT_38_0b1_iFi_ETC__q79 =
	      iFifo$D_OUT[38];
      2'd3:
	  CASE_guard32950_0b0_iFifoD_OUT_BIT_38_0b1_iFi_ETC__q79 =
	      guard__h232950 == 2'b11 && iFifo$D_OUT[38];
    endcase
  end
  always@(iFifo$D_OUT or
	  CASE_guard32950_0b0_iFifoD_OUT_BIT_38_0b1_iFi_ETC__q79 or
	  guard__h232950)
  begin
    case (iFifo$D_OUT[6:4])
      3'd0:
	  CASE_iFifoD_OUT_BITS_6_TO_4_0_CASE_guard32950_ETC__q80 =
	      CASE_guard32950_0b0_iFifoD_OUT_BIT_38_0b1_iFi_ETC__q79;
      3'd1:
	  CASE_iFifoD_OUT_BITS_6_TO_4_0_CASE_guard32950_ETC__q80 =
	      (guard__h232950 == 2'b0) ?
		iFifo$D_OUT[38] :
		(guard__h232950 == 2'b01 || guard__h232950 == 2'b10 ||
		 guard__h232950 == 2'b11) &&
		iFifo$D_OUT[38];
      3'd2, 3'd3:
	  CASE_iFifoD_OUT_BITS_6_TO_4_0_CASE_guard32950_ETC__q80 =
	      iFifo$D_OUT[38];
      default: CASE_iFifoD_OUT_BITS_6_TO_4_0_CASE_guard32950_ETC__q80 =
		   iFifo$D_OUT[6:4] == 3'd4 && iFifo$D_OUT[38];
    endcase
  end
  always@(guard__h251238 or
	  _theResult___snd__h259174 or
	  out_sfd__h259902 or _theResult___sfd__h259899)
  begin
    case (guard__h251238)
      2'b0, 2'b01:
	  CASE_guard51238_0b0_theResult___snd59174_BITS__ETC__q81 =
	      _theResult___snd__h259174[56:5];
      2'b10:
	  CASE_guard51238_0b0_theResult___snd59174_BITS__ETC__q81 =
	      out_sfd__h259902;
      2'b11:
	  CASE_guard51238_0b0_theResult___snd59174_BITS__ETC__q81 =
	      _theResult___sfd__h259899;
    endcase
  end
  always@(guard__h251238 or
	  _theResult___snd__h259174 or _theResult___sfd__h259899)
  begin
    case (guard__h251238)
      2'b0:
	  CASE_guard51238_0b0_theResult___snd59174_BITS__ETC__q82 =
	      _theResult___snd__h259174[56:5];
      2'b01, 2'b10, 2'b11:
	  CASE_guard51238_0b0_theResult___snd59174_BITS__ETC__q82 =
	      _theResult___sfd__h259899;
    endcase
  end
  always@(iFifo$D_OUT or
	  CASE_guard51238_0b0_theResult___snd59174_BITS__ETC__q81 or
	  CASE_guard51238_0b0_theResult___snd59174_BITS__ETC__q82 or
	  IF_IF_IF_iFifo_first__087_BITS_37_TO_30_850_EQ_ETC___d4538 or
	  IF_IF_IF_iFifo_first__087_BITS_37_TO_30_850_EQ_ETC___d4540 or
	  _theResult___snd__h259174)
  begin
    case (iFifo$D_OUT[6:4])
      3'd0:
	  _theResult___fst_sfd__h259977 =
	      CASE_guard51238_0b0_theResult___snd59174_BITS__ETC__q81;
      3'd1:
	  _theResult___fst_sfd__h259977 =
	      CASE_guard51238_0b0_theResult___snd59174_BITS__ETC__q82;
      3'd2:
	  _theResult___fst_sfd__h259977 =
	      IF_IF_IF_iFifo_first__087_BITS_37_TO_30_850_EQ_ETC___d4538;
      3'd3:
	  _theResult___fst_sfd__h259977 =
	      IF_IF_IF_iFifo_first__087_BITS_37_TO_30_850_EQ_ETC___d4540;
      3'd4: _theResult___fst_sfd__h259977 = _theResult___snd__h259174[56:5];
      default: _theResult___fst_sfd__h259977 = 52'd0;
    endcase
  end
  always@(iFifo$D_OUT)
  begin
    case (iFifo$D_OUT[6:4])
      3'd0, 3'd1, 3'd2, 3'd3:
	  IF_iFifo_first__087_BITS_6_TO_4_118_EQ_0_191_O_ETC___d4028 =
	      iFifo$D_OUT[38];
      default: IF_iFifo_first__087_BITS_6_TO_4_118_EQ_0_191_O_ETC___d4028 =
		   iFifo$D_OUT[6:4] == 3'd4 && iFifo$D_OUT[38];
    endcase
  end
  always@(guard__h242199 or iFifo$D_OUT)
  begin
    case (guard__h242199)
      2'b0, 2'b01, 2'b10:
	  CASE_guard42199_0b0_iFifoD_OUT_BIT_38_0b1_iFi_ETC__q83 =
	      iFifo$D_OUT[38];
      2'd3:
	  CASE_guard42199_0b0_iFifoD_OUT_BIT_38_0b1_iFi_ETC__q83 =
	      guard__h242199 == 2'b11 && iFifo$D_OUT[38];
    endcase
  end
  always@(iFifo$D_OUT or
	  CASE_guard42199_0b0_iFifoD_OUT_BIT_38_0b1_iFi_ETC__q83 or
	  guard__h242199)
  begin
    case (iFifo$D_OUT[6:4])
      3'd0:
	  CASE_iFifoD_OUT_BITS_6_TO_4_0_CASE_guard42199_ETC__q84 =
	      CASE_guard42199_0b0_iFifoD_OUT_BIT_38_0b1_iFi_ETC__q83;
      3'd1:
	  CASE_iFifoD_OUT_BITS_6_TO_4_0_CASE_guard42199_ETC__q84 =
	      (guard__h242199 == 2'b0) ?
		iFifo$D_OUT[38] :
		(guard__h242199 == 2'b01 || guard__h242199 == 2'b10 ||
		 guard__h242199 == 2'b11) &&
		iFifo$D_OUT[38];
      3'd2, 3'd3:
	  CASE_iFifoD_OUT_BITS_6_TO_4_0_CASE_guard42199_ETC__q84 =
	      iFifo$D_OUT[38];
      default: CASE_iFifoD_OUT_BITS_6_TO_4_0_CASE_guard42199_ETC__q84 =
		   iFifo$D_OUT[6:4] == 3'd4 && iFifo$D_OUT[38];
    endcase
  end
  always@(guard__h251238 or iFifo$D_OUT)
  begin
    case (guard__h251238)
      2'b0, 2'b01, 2'b10:
	  CASE_guard51238_0b0_iFifoD_OUT_BIT_38_0b1_iFi_ETC__q85 =
	      iFifo$D_OUT[38];
      2'd3:
	  CASE_guard51238_0b0_iFifoD_OUT_BIT_38_0b1_iFi_ETC__q85 =
	      guard__h251238 == 2'b11 && iFifo$D_OUT[38];
    endcase
  end
  always@(iFifo$D_OUT or
	  CASE_guard51238_0b0_iFifoD_OUT_BIT_38_0b1_iFi_ETC__q85 or
	  guard__h251238)
  begin
    case (iFifo$D_OUT[6:4])
      3'd0:
	  CASE_iFifoD_OUT_BITS_6_TO_4_0_CASE_guard51238_ETC__q86 =
	      CASE_guard51238_0b0_iFifoD_OUT_BIT_38_0b1_iFi_ETC__q85;
      3'd1:
	  CASE_iFifoD_OUT_BITS_6_TO_4_0_CASE_guard51238_ETC__q86 =
	      (guard__h251238 == 2'b0) ?
		iFifo$D_OUT[38] :
		(guard__h251238 == 2'b01 || guard__h251238 == 2'b10 ||
		 guard__h251238 == 2'b11) &&
		iFifo$D_OUT[38];
      3'd2, 3'd3:
	  CASE_iFifoD_OUT_BITS_6_TO_4_0_CASE_guard51238_ETC__q86 =
	      iFifo$D_OUT[38];
      default: CASE_iFifoD_OUT_BITS_6_TO_4_0_CASE_guard51238_ETC__q86 =
		   iFifo$D_OUT[6:4] == 3'd4 && iFifo$D_OUT[38];
    endcase
  end
  always@(guard__h232950 or iFifo$D_OUT)
  begin
    case (guard__h232950)
      2'b0, 2'b01, 2'b10:
	  CASE_guard32950_0b0_NOT_iFifoD_OUT_BIT_38_0b1_ETC__q87 =
	      !iFifo$D_OUT[38];
      2'd3:
	  CASE_guard32950_0b0_NOT_iFifoD_OUT_BIT_38_0b1_ETC__q87 =
	      guard__h232950 != 2'b11 || !iFifo$D_OUT[38];
    endcase
  end
  always@(iFifo$D_OUT or
	  CASE_guard32950_0b0_NOT_iFifoD_OUT_BIT_38_0b1_ETC__q87 or
	  guard__h232950)
  begin
    case (iFifo$D_OUT[6:4])
      3'd0:
	  CASE_iFifoD_OUT_BITS_6_TO_4_0_CASE_guard32950_ETC__q88 =
	      CASE_guard32950_0b0_NOT_iFifoD_OUT_BIT_38_0b1_ETC__q87;
      3'd1:
	  CASE_iFifoD_OUT_BITS_6_TO_4_0_CASE_guard32950_ETC__q88 =
	      (guard__h232950 == 2'b0) ?
		!iFifo$D_OUT[38] :
		guard__h232950 != 2'b01 && guard__h232950 != 2'b10 &&
		guard__h232950 != 2'b11 ||
		!iFifo$D_OUT[38];
      3'd2, 3'd3:
	  CASE_iFifoD_OUT_BITS_6_TO_4_0_CASE_guard32950_ETC__q88 =
	      !iFifo$D_OUT[38];
      default: CASE_iFifoD_OUT_BITS_6_TO_4_0_CASE_guard32950_ETC__q88 =
		   iFifo$D_OUT[6:4] != 3'd4 || !iFifo$D_OUT[38];
    endcase
  end
  always@(guard__h242199 or iFifo$D_OUT)
  begin
    case (guard__h242199)
      2'b0, 2'b01, 2'b10:
	  CASE_guard42199_0b0_NOT_iFifoD_OUT_BIT_38_0b1_ETC__q89 =
	      !iFifo$D_OUT[38];
      2'd3:
	  CASE_guard42199_0b0_NOT_iFifoD_OUT_BIT_38_0b1_ETC__q89 =
	      guard__h242199 != 2'b11 || !iFifo$D_OUT[38];
    endcase
  end
  always@(iFifo$D_OUT or
	  CASE_guard42199_0b0_NOT_iFifoD_OUT_BIT_38_0b1_ETC__q89 or
	  guard__h242199)
  begin
    case (iFifo$D_OUT[6:4])
      3'd0:
	  CASE_iFifoD_OUT_BITS_6_TO_4_0_CASE_guard42199_ETC__q90 =
	      CASE_guard42199_0b0_NOT_iFifoD_OUT_BIT_38_0b1_ETC__q89;
      3'd1:
	  CASE_iFifoD_OUT_BITS_6_TO_4_0_CASE_guard42199_ETC__q90 =
	      (guard__h242199 == 2'b0) ?
		!iFifo$D_OUT[38] :
		guard__h242199 != 2'b01 && guard__h242199 != 2'b10 &&
		guard__h242199 != 2'b11 ||
		!iFifo$D_OUT[38];
      3'd2, 3'd3:
	  CASE_iFifoD_OUT_BITS_6_TO_4_0_CASE_guard42199_ETC__q90 =
	      !iFifo$D_OUT[38];
      default: CASE_iFifoD_OUT_BITS_6_TO_4_0_CASE_guard42199_ETC__q90 =
		   iFifo$D_OUT[6:4] != 3'd4 || !iFifo$D_OUT[38];
    endcase
  end
  always@(guard__h251238 or iFifo$D_OUT)
  begin
    case (guard__h251238)
      2'b0, 2'b01, 2'b10:
	  CASE_guard51238_0b0_NOT_iFifoD_OUT_BIT_38_0b1_ETC__q91 =
	      !iFifo$D_OUT[38];
      2'd3:
	  CASE_guard51238_0b0_NOT_iFifoD_OUT_BIT_38_0b1_ETC__q91 =
	      guard__h251238 != 2'b11 || !iFifo$D_OUT[38];
    endcase
  end
  always@(iFifo$D_OUT or
	  CASE_guard51238_0b0_NOT_iFifoD_OUT_BIT_38_0b1_ETC__q91 or
	  guard__h251238)
  begin
    case (iFifo$D_OUT[6:4])
      3'd0:
	  CASE_iFifoD_OUT_BITS_6_TO_4_0_CASE_guard51238_ETC__q92 =
	      CASE_guard51238_0b0_NOT_iFifoD_OUT_BIT_38_0b1_ETC__q91;
      3'd1:
	  CASE_iFifoD_OUT_BITS_6_TO_4_0_CASE_guard51238_ETC__q92 =
	      (guard__h251238 == 2'b0) ?
		!iFifo$D_OUT[38] :
		guard__h251238 != 2'b01 && guard__h251238 != 2'b10 &&
		guard__h251238 != 2'b11 ||
		!iFifo$D_OUT[38];
      3'd2, 3'd3:
	  CASE_iFifoD_OUT_BITS_6_TO_4_0_CASE_guard51238_ETC__q92 =
	      !iFifo$D_OUT[38];
      default: CASE_iFifoD_OUT_BITS_6_TO_4_0_CASE_guard51238_ETC__q92 =
		   iFifo$D_OUT[6:4] != 3'd4 || !iFifo$D_OUT[38];
    endcase
  end
  always@(iFifo$D_OUT)
  begin
    case (iFifo$D_OUT[6:4])
      3'd0, 3'd1, 3'd2, 3'd3:
	  IF_iFifo_first__087_BITS_6_TO_4_118_EQ_0_191_O_ETC___d4582 =
	      !iFifo$D_OUT[38];
      default: IF_iFifo_first__087_BITS_6_TO_4_118_EQ_0_191_O_ETC___d4582 =
		   iFifo$D_OUT[6:4] != 3'd4 || !iFifo$D_OUT[38];
    endcase
  end
  always@(guard__h194011 or
	  _theResult___fst_exp__h201972 or
	  out_exp__h202620 or _theResult___exp__h202617)
  begin
    case (guard__h194011)
      2'b0, 2'b01:
	  CASE_guard94011_0b0_theResult___fst_exp01972_0_ETC__q102 =
	      _theResult___fst_exp__h201972;
      2'b10:
	  CASE_guard94011_0b0_theResult___fst_exp01972_0_ETC__q102 =
	      out_exp__h202620;
      2'b11:
	  CASE_guard94011_0b0_theResult___fst_exp01972_0_ETC__q102 =
	      _theResult___exp__h202617;
    endcase
  end
  always@(guard__h194011 or
	  _theResult___fst_exp__h201972 or _theResult___exp__h202617)
  begin
    case (guard__h194011)
      2'b0:
	  CASE_guard94011_0b0_theResult___fst_exp01972_0_ETC__q103 =
	      _theResult___fst_exp__h201972;
      2'b01, 2'b10, 2'b11:
	  CASE_guard94011_0b0_theResult___fst_exp01972_0_ETC__q103 =
	      _theResult___exp__h202617;
    endcase
  end
  always@(iFifo$D_OUT or
	  CASE_guard94011_0b0_theResult___fst_exp01972_0_ETC__q102 or
	  CASE_guard94011_0b0_theResult___fst_exp01972_0_ETC__q103 or
	  IF_IF_IF_iFifo_first__087_BITS_102_TO_95_625_E_ETC___d5173 or
	  IF_IF_IF_iFifo_first__087_BITS_102_TO_95_625_E_ETC___d5175 or
	  _theResult___fst_exp__h201972)
  begin
    case (iFifo$D_OUT[6:4])
      3'd0:
	  _theResult___fst_exp__h202695 =
	      CASE_guard94011_0b0_theResult___fst_exp01972_0_ETC__q102;
      3'd1:
	  _theResult___fst_exp__h202695 =
	      CASE_guard94011_0b0_theResult___fst_exp01972_0_ETC__q103;
      3'd2:
	  _theResult___fst_exp__h202695 =
	      IF_IF_IF_iFifo_first__087_BITS_102_TO_95_625_E_ETC___d5173;
      3'd3:
	  _theResult___fst_exp__h202695 =
	      IF_IF_IF_iFifo_first__087_BITS_102_TO_95_625_E_ETC___d5175;
      3'd4: _theResult___fst_exp__h202695 = _theResult___fst_exp__h201972;
      default: _theResult___fst_exp__h202695 = 11'd0;
    endcase
  end
  always@(guard__h203260 or
	  _theResult___fst_exp__h211488 or
	  out_exp__h212210 or _theResult___exp__h212207)
  begin
    case (guard__h203260)
      2'b0, 2'b01:
	  CASE_guard03260_0b0_theResult___fst_exp11488_0_ETC__q104 =
	      _theResult___fst_exp__h211488;
      2'b10:
	  CASE_guard03260_0b0_theResult___fst_exp11488_0_ETC__q104 =
	      out_exp__h212210;
      2'b11:
	  CASE_guard03260_0b0_theResult___fst_exp11488_0_ETC__q104 =
	      _theResult___exp__h212207;
    endcase
  end
  always@(guard__h203260 or
	  _theResult___fst_exp__h211488 or _theResult___exp__h212207)
  begin
    case (guard__h203260)
      2'b0:
	  CASE_guard03260_0b0_theResult___fst_exp11488_0_ETC__q105 =
	      _theResult___fst_exp__h211488;
      2'b01, 2'b10, 2'b11:
	  CASE_guard03260_0b0_theResult___fst_exp11488_0_ETC__q105 =
	      _theResult___exp__h212207;
    endcase
  end
  always@(iFifo$D_OUT or
	  CASE_guard03260_0b0_theResult___fst_exp11488_0_ETC__q104 or
	  CASE_guard03260_0b0_theResult___fst_exp11488_0_ETC__q105 or
	  IF_IF_IF_IF_3074_MINUS_SEXT_iFifo_first__087_B_ETC___d5211 or
	  IF_IF_IF_IF_3074_MINUS_SEXT_iFifo_first__087_B_ETC___d5213 or
	  _theResult___fst_exp__h211488)
  begin
    case (iFifo$D_OUT[6:4])
      3'd0:
	  _theResult___fst_exp__h212285 =
	      CASE_guard03260_0b0_theResult___fst_exp11488_0_ETC__q104;
      3'd1:
	  _theResult___fst_exp__h212285 =
	      CASE_guard03260_0b0_theResult___fst_exp11488_0_ETC__q105;
      3'd2:
	  _theResult___fst_exp__h212285 =
	      IF_IF_IF_IF_3074_MINUS_SEXT_iFifo_first__087_B_ETC___d5211;
      3'd3:
	  _theResult___fst_exp__h212285 =
	      IF_IF_IF_IF_3074_MINUS_SEXT_iFifo_first__087_B_ETC___d5213;
      3'd4: _theResult___fst_exp__h212285 = _theResult___fst_exp__h211488;
      default: _theResult___fst_exp__h212285 = 11'd0;
    endcase
  end
  always@(guard__h212299 or
	  _theResult___fst_exp__h220289 or
	  out_exp__h220962 or _theResult___exp__h220959)
  begin
    case (guard__h212299)
      2'b0, 2'b01:
	  CASE_guard12299_0b0_theResult___fst_exp20289_0_ETC__q106 =
	      _theResult___fst_exp__h220289;
      2'b10:
	  CASE_guard12299_0b0_theResult___fst_exp20289_0_ETC__q106 =
	      out_exp__h220962;
      2'b11:
	  CASE_guard12299_0b0_theResult___fst_exp20289_0_ETC__q106 =
	      _theResult___exp__h220959;
    endcase
  end
  always@(guard__h212299 or
	  _theResult___fst_exp__h220289 or _theResult___exp__h220959)
  begin
    case (guard__h212299)
      2'b0:
	  CASE_guard12299_0b0_theResult___fst_exp20289_0_ETC__q107 =
	      _theResult___fst_exp__h220289;
      2'b01, 2'b10, 2'b11:
	  CASE_guard12299_0b0_theResult___fst_exp20289_0_ETC__q107 =
	      _theResult___exp__h220959;
    endcase
  end
  always@(iFifo$D_OUT or
	  CASE_guard12299_0b0_theResult___fst_exp20289_0_ETC__q106 or
	  CASE_guard12299_0b0_theResult___fst_exp20289_0_ETC__q107 or
	  IF_IF_IF_iFifo_first__087_BITS_102_TO_95_625_E_ETC___d5242 or
	  IF_IF_IF_iFifo_first__087_BITS_102_TO_95_625_E_ETC___d5244 or
	  _theResult___fst_exp__h220289)
  begin
    case (iFifo$D_OUT[6:4])
      3'd0:
	  _theResult___fst_exp__h221037 =
	      CASE_guard12299_0b0_theResult___fst_exp20289_0_ETC__q106;
      3'd1:
	  _theResult___fst_exp__h221037 =
	      CASE_guard12299_0b0_theResult___fst_exp20289_0_ETC__q107;
      3'd2:
	  _theResult___fst_exp__h221037 =
	      IF_IF_IF_iFifo_first__087_BITS_102_TO_95_625_E_ETC___d5242;
      3'd3:
	  _theResult___fst_exp__h221037 =
	      IF_IF_IF_iFifo_first__087_BITS_102_TO_95_625_E_ETC___d5244;
      3'd4: _theResult___fst_exp__h221037 = _theResult___fst_exp__h220289;
      default: _theResult___fst_exp__h221037 = 11'd0;
    endcase
  end
  always@(guard__h194011 or
	  _theResult___snd__h201923 or
	  out_sfd__h202621 or _theResult___sfd__h202618)
  begin
    case (guard__h194011)
      2'b0, 2'b01:
	  CASE_guard94011_0b0_theResult___snd01923_BITS__ETC__q108 =
	      _theResult___snd__h201923[56:5];
      2'b10:
	  CASE_guard94011_0b0_theResult___snd01923_BITS__ETC__q108 =
	      out_sfd__h202621;
      2'b11:
	  CASE_guard94011_0b0_theResult___snd01923_BITS__ETC__q108 =
	      _theResult___sfd__h202618;
    endcase
  end
  always@(guard__h194011 or
	  _theResult___snd__h201923 or _theResult___sfd__h202618)
  begin
    case (guard__h194011)
      2'b0:
	  CASE_guard94011_0b0_theResult___snd01923_BITS__ETC__q109 =
	      _theResult___snd__h201923[56:5];
      2'b01, 2'b10, 2'b11:
	  CASE_guard94011_0b0_theResult___snd01923_BITS__ETC__q109 =
	      _theResult___sfd__h202618;
    endcase
  end
  always@(iFifo$D_OUT or
	  CASE_guard94011_0b0_theResult___snd01923_BITS__ETC__q108 or
	  CASE_guard94011_0b0_theResult___snd01923_BITS__ETC__q109 or
	  IF_IF_IF_iFifo_first__087_BITS_102_TO_95_625_E_ETC___d5268 or
	  IF_IF_IF_iFifo_first__087_BITS_102_TO_95_625_E_ETC___d5270 or
	  _theResult___snd__h201923)
  begin
    case (iFifo$D_OUT[6:4])
      3'd0:
	  _theResult___fst_sfd__h202696 =
	      CASE_guard94011_0b0_theResult___snd01923_BITS__ETC__q108;
      3'd1:
	  _theResult___fst_sfd__h202696 =
	      CASE_guard94011_0b0_theResult___snd01923_BITS__ETC__q109;
      3'd2:
	  _theResult___fst_sfd__h202696 =
	      IF_IF_IF_iFifo_first__087_BITS_102_TO_95_625_E_ETC___d5268;
      3'd3:
	  _theResult___fst_sfd__h202696 =
	      IF_IF_IF_iFifo_first__087_BITS_102_TO_95_625_E_ETC___d5270;
      3'd4: _theResult___fst_sfd__h202696 = _theResult___snd__h201923[56:5];
      default: _theResult___fst_sfd__h202696 = 52'd0;
    endcase
  end
  always@(guard__h203260 or
	  sfdin__h211482 or out_sfd__h212211 or _theResult___sfd__h212208)
  begin
    case (guard__h203260)
      2'b0, 2'b01:
	  CASE_guard03260_0b0_sfdin11482_BITS_56_TO_5_0b_ETC__q110 =
	      sfdin__h211482[56:5];
      2'b10:
	  CASE_guard03260_0b0_sfdin11482_BITS_56_TO_5_0b_ETC__q110 =
	      out_sfd__h212211;
      2'b11:
	  CASE_guard03260_0b0_sfdin11482_BITS_56_TO_5_0b_ETC__q110 =
	      _theResult___sfd__h212208;
    endcase
  end
  always@(guard__h203260 or sfdin__h211482 or _theResult___sfd__h212208)
  begin
    case (guard__h203260)
      2'b0:
	  CASE_guard03260_0b0_sfdin11482_BITS_56_TO_5_0b_ETC__q111 =
	      sfdin__h211482[56:5];
      2'b01, 2'b10, 2'b11:
	  CASE_guard03260_0b0_sfdin11482_BITS_56_TO_5_0b_ETC__q111 =
	      _theResult___sfd__h212208;
    endcase
  end
  always@(iFifo$D_OUT or
	  CASE_guard03260_0b0_sfdin11482_BITS_56_TO_5_0b_ETC__q110 or
	  CASE_guard03260_0b0_sfdin11482_BITS_56_TO_5_0b_ETC__q111 or
	  IF_IF_IF_IF_3074_MINUS_SEXT_iFifo_first__087_B_ETC___d5294 or
	  IF_IF_IF_IF_3074_MINUS_SEXT_iFifo_first__087_B_ETC___d5296 or
	  sfdin__h211482)
  begin
    case (iFifo$D_OUT[6:4])
      3'd0:
	  _theResult___fst_sfd__h212286 =
	      CASE_guard03260_0b0_sfdin11482_BITS_56_TO_5_0b_ETC__q110;
      3'd1:
	  _theResult___fst_sfd__h212286 =
	      CASE_guard03260_0b0_sfdin11482_BITS_56_TO_5_0b_ETC__q111;
      3'd2:
	  _theResult___fst_sfd__h212286 =
	      IF_IF_IF_IF_3074_MINUS_SEXT_iFifo_first__087_B_ETC___d5294;
      3'd3:
	  _theResult___fst_sfd__h212286 =
	      IF_IF_IF_IF_3074_MINUS_SEXT_iFifo_first__087_B_ETC___d5296;
      3'd4: _theResult___fst_sfd__h212286 = sfdin__h211482[56:5];
      default: _theResult___fst_sfd__h212286 = 52'd0;
    endcase
  end
  always@(guard__h212299 or
	  _theResult___snd__h220235 or
	  out_sfd__h220963 or _theResult___sfd__h220960)
  begin
    case (guard__h212299)
      2'b0, 2'b01:
	  CASE_guard12299_0b0_theResult___snd20235_BITS__ETC__q112 =
	      _theResult___snd__h220235[56:5];
      2'b10:
	  CASE_guard12299_0b0_theResult___snd20235_BITS__ETC__q112 =
	      out_sfd__h220963;
      2'b11:
	  CASE_guard12299_0b0_theResult___snd20235_BITS__ETC__q112 =
	      _theResult___sfd__h220960;
    endcase
  end
  always@(guard__h212299 or
	  _theResult___snd__h220235 or _theResult___sfd__h220960)
  begin
    case (guard__h212299)
      2'b0:
	  CASE_guard12299_0b0_theResult___snd20235_BITS__ETC__q113 =
	      _theResult___snd__h220235[56:5];
      2'b01, 2'b10, 2'b11:
	  CASE_guard12299_0b0_theResult___snd20235_BITS__ETC__q113 =
	      _theResult___sfd__h220960;
    endcase
  end
  always@(iFifo$D_OUT or
	  CASE_guard12299_0b0_theResult___snd20235_BITS__ETC__q112 or
	  CASE_guard12299_0b0_theResult___snd20235_BITS__ETC__q113 or
	  IF_IF_IF_iFifo_first__087_BITS_102_TO_95_625_E_ETC___d5313 or
	  IF_IF_IF_iFifo_first__087_BITS_102_TO_95_625_E_ETC___d5315 or
	  _theResult___snd__h220235)
  begin
    case (iFifo$D_OUT[6:4])
      3'd0:
	  _theResult___fst_sfd__h221038 =
	      CASE_guard12299_0b0_theResult___snd20235_BITS__ETC__q112;
      3'd1:
	  _theResult___fst_sfd__h221038 =
	      CASE_guard12299_0b0_theResult___snd20235_BITS__ETC__q113;
      3'd2:
	  _theResult___fst_sfd__h221038 =
	      IF_IF_IF_iFifo_first__087_BITS_102_TO_95_625_E_ETC___d5313;
      3'd3:
	  _theResult___fst_sfd__h221038 =
	      IF_IF_IF_iFifo_first__087_BITS_102_TO_95_625_E_ETC___d5315;
      3'd4: _theResult___fst_sfd__h221038 = _theResult___snd__h220235[56:5];
      default: _theResult___fst_sfd__h221038 = 52'd0;
    endcase
  end
  always@(guard__h194011 or iFifo$D_OUT)
  begin
    case (guard__h194011)
      2'b0, 2'b01, 2'b10:
	  CASE_guard94011_0b0_iFifoD_OUT_BIT_103_0b1_iF_ETC__q114 =
	      iFifo$D_OUT[103];
      2'd3:
	  CASE_guard94011_0b0_iFifoD_OUT_BIT_103_0b1_iF_ETC__q114 =
	      guard__h194011 == 2'b11 && iFifo$D_OUT[103];
    endcase
  end
  always@(iFifo$D_OUT or
	  CASE_guard94011_0b0_iFifoD_OUT_BIT_103_0b1_iF_ETC__q114 or
	  guard__h194011)
  begin
    case (iFifo$D_OUT[6:4])
      3'd0:
	  CASE_iFifoD_OUT_BITS_6_TO_4_0_CASE_guard94011_ETC__q115 =
	      CASE_guard94011_0b0_iFifoD_OUT_BIT_103_0b1_iF_ETC__q114;
      3'd1:
	  CASE_iFifoD_OUT_BITS_6_TO_4_0_CASE_guard94011_ETC__q115 =
	      (guard__h194011 == 2'b0) ?
		iFifo$D_OUT[103] :
		(guard__h194011 == 2'b01 || guard__h194011 == 2'b10 ||
		 guard__h194011 == 2'b11) &&
		iFifo$D_OUT[103];
      3'd2, 3'd3:
	  CASE_iFifoD_OUT_BITS_6_TO_4_0_CASE_guard94011_ETC__q115 =
	      iFifo$D_OUT[103];
      default: CASE_iFifoD_OUT_BITS_6_TO_4_0_CASE_guard94011_ETC__q115 =
		   iFifo$D_OUT[6:4] == 3'd4 && iFifo$D_OUT[103];
    endcase
  end
  always@(iFifo$D_OUT)
  begin
    case (iFifo$D_OUT[6:4])
      3'd0, 3'd1, 3'd2, 3'd3:
	  IF_iFifo_first__087_BITS_6_TO_4_118_EQ_0_191_O_ETC___d4803 =
	      iFifo$D_OUT[103];
      default: IF_iFifo_first__087_BITS_6_TO_4_118_EQ_0_191_O_ETC___d4803 =
		   iFifo$D_OUT[6:4] == 3'd4 && iFifo$D_OUT[103];
    endcase
  end
  always@(guard__h203260 or iFifo$D_OUT)
  begin
    case (guard__h203260)
      2'b0, 2'b01, 2'b10:
	  CASE_guard03260_0b0_iFifoD_OUT_BIT_103_0b1_iF_ETC__q116 =
	      iFifo$D_OUT[103];
      2'd3:
	  CASE_guard03260_0b0_iFifoD_OUT_BIT_103_0b1_iF_ETC__q116 =
	      guard__h203260 == 2'b11 && iFifo$D_OUT[103];
    endcase
  end
  always@(iFifo$D_OUT or
	  CASE_guard03260_0b0_iFifoD_OUT_BIT_103_0b1_iF_ETC__q116 or
	  guard__h203260)
  begin
    case (iFifo$D_OUT[6:4])
      3'd0:
	  CASE_iFifoD_OUT_BITS_6_TO_4_0_CASE_guard03260_ETC__q117 =
	      CASE_guard03260_0b0_iFifoD_OUT_BIT_103_0b1_iF_ETC__q116;
      3'd1:
	  CASE_iFifoD_OUT_BITS_6_TO_4_0_CASE_guard03260_ETC__q117 =
	      (guard__h203260 == 2'b0) ?
		iFifo$D_OUT[103] :
		(guard__h203260 == 2'b01 || guard__h203260 == 2'b10 ||
		 guard__h203260 == 2'b11) &&
		iFifo$D_OUT[103];
      3'd2, 3'd3:
	  CASE_iFifoD_OUT_BITS_6_TO_4_0_CASE_guard03260_ETC__q117 =
	      iFifo$D_OUT[103];
      default: CASE_iFifoD_OUT_BITS_6_TO_4_0_CASE_guard03260_ETC__q117 =
		   iFifo$D_OUT[6:4] == 3'd4 && iFifo$D_OUT[103];
    endcase
  end
  always@(guard__h212299 or iFifo$D_OUT)
  begin
    case (guard__h212299)
      2'b0, 2'b01, 2'b10:
	  CASE_guard12299_0b0_iFifoD_OUT_BIT_103_0b1_iF_ETC__q118 =
	      iFifo$D_OUT[103];
      2'd3:
	  CASE_guard12299_0b0_iFifoD_OUT_BIT_103_0b1_iF_ETC__q118 =
	      guard__h212299 == 2'b11 && iFifo$D_OUT[103];
    endcase
  end
  always@(iFifo$D_OUT or
	  CASE_guard12299_0b0_iFifoD_OUT_BIT_103_0b1_iF_ETC__q118 or
	  guard__h212299)
  begin
    case (iFifo$D_OUT[6:4])
      3'd0:
	  CASE_iFifoD_OUT_BITS_6_TO_4_0_CASE_guard12299_ETC__q119 =
	      CASE_guard12299_0b0_iFifoD_OUT_BIT_103_0b1_iF_ETC__q118;
      3'd1:
	  CASE_iFifoD_OUT_BITS_6_TO_4_0_CASE_guard12299_ETC__q119 =
	      (guard__h212299 == 2'b0) ?
		iFifo$D_OUT[103] :
		(guard__h212299 == 2'b01 || guard__h212299 == 2'b10 ||
		 guard__h212299 == 2'b11) &&
		iFifo$D_OUT[103];
      3'd2, 3'd3:
	  CASE_iFifoD_OUT_BITS_6_TO_4_0_CASE_guard12299_ETC__q119 =
	      iFifo$D_OUT[103];
      default: CASE_iFifoD_OUT_BITS_6_TO_4_0_CASE_guard12299_ETC__q119 =
		   iFifo$D_OUT[6:4] == 3'd4 && iFifo$D_OUT[103];
    endcase
  end
  always@(guard__h194011 or iFifo$D_OUT)
  begin
    case (guard__h194011)
      2'b0, 2'b01, 2'b10:
	  CASE_guard94011_0b0_NOT_iFifoD_OUT_BIT_103_0b_ETC__q120 =
	      !iFifo$D_OUT[103];
      2'd3:
	  CASE_guard94011_0b0_NOT_iFifoD_OUT_BIT_103_0b_ETC__q120 =
	      guard__h194011 != 2'b11 || !iFifo$D_OUT[103];
    endcase
  end
  always@(iFifo$D_OUT or
	  CASE_guard94011_0b0_NOT_iFifoD_OUT_BIT_103_0b_ETC__q120 or
	  guard__h194011)
  begin
    case (iFifo$D_OUT[6:4])
      3'd0:
	  CASE_iFifoD_OUT_BITS_6_TO_4_0_CASE_guard94011_ETC__q121 =
	      CASE_guard94011_0b0_NOT_iFifoD_OUT_BIT_103_0b_ETC__q120;
      3'd1:
	  CASE_iFifoD_OUT_BITS_6_TO_4_0_CASE_guard94011_ETC__q121 =
	      (guard__h194011 == 2'b0) ?
		!iFifo$D_OUT[103] :
		guard__h194011 != 2'b01 && guard__h194011 != 2'b10 &&
		guard__h194011 != 2'b11 ||
		!iFifo$D_OUT[103];
      3'd2, 3'd3:
	  CASE_iFifoD_OUT_BITS_6_TO_4_0_CASE_guard94011_ETC__q121 =
	      !iFifo$D_OUT[103];
      default: CASE_iFifoD_OUT_BITS_6_TO_4_0_CASE_guard94011_ETC__q121 =
		   iFifo$D_OUT[6:4] != 3'd4 || !iFifo$D_OUT[103];
    endcase
  end
  always@(guard__h203260 or iFifo$D_OUT)
  begin
    case (guard__h203260)
      2'b0, 2'b01, 2'b10:
	  CASE_guard03260_0b0_NOT_iFifoD_OUT_BIT_103_0b_ETC__q122 =
	      !iFifo$D_OUT[103];
      2'd3:
	  CASE_guard03260_0b0_NOT_iFifoD_OUT_BIT_103_0b_ETC__q122 =
	      guard__h203260 != 2'b11 || !iFifo$D_OUT[103];
    endcase
  end
  always@(iFifo$D_OUT or
	  CASE_guard03260_0b0_NOT_iFifoD_OUT_BIT_103_0b_ETC__q122 or
	  guard__h203260)
  begin
    case (iFifo$D_OUT[6:4])
      3'd0:
	  CASE_iFifoD_OUT_BITS_6_TO_4_0_CASE_guard03260_ETC__q123 =
	      CASE_guard03260_0b0_NOT_iFifoD_OUT_BIT_103_0b_ETC__q122;
      3'd1:
	  CASE_iFifoD_OUT_BITS_6_TO_4_0_CASE_guard03260_ETC__q123 =
	      (guard__h203260 == 2'b0) ?
		!iFifo$D_OUT[103] :
		guard__h203260 != 2'b01 && guard__h203260 != 2'b10 &&
		guard__h203260 != 2'b11 ||
		!iFifo$D_OUT[103];
      3'd2, 3'd3:
	  CASE_iFifoD_OUT_BITS_6_TO_4_0_CASE_guard03260_ETC__q123 =
	      !iFifo$D_OUT[103];
      default: CASE_iFifoD_OUT_BITS_6_TO_4_0_CASE_guard03260_ETC__q123 =
		   iFifo$D_OUT[6:4] != 3'd4 || !iFifo$D_OUT[103];
    endcase
  end
  always@(guard__h212299 or iFifo$D_OUT)
  begin
    case (guard__h212299)
      2'b0, 2'b01, 2'b10:
	  CASE_guard12299_0b0_NOT_iFifoD_OUT_BIT_103_0b_ETC__q124 =
	      !iFifo$D_OUT[103];
      2'd3:
	  CASE_guard12299_0b0_NOT_iFifoD_OUT_BIT_103_0b_ETC__q124 =
	      guard__h212299 != 2'b11 || !iFifo$D_OUT[103];
    endcase
  end
  always@(iFifo$D_OUT or
	  CASE_guard12299_0b0_NOT_iFifoD_OUT_BIT_103_0b_ETC__q124 or
	  guard__h212299)
  begin
    case (iFifo$D_OUT[6:4])
      3'd0:
	  CASE_iFifoD_OUT_BITS_6_TO_4_0_CASE_guard12299_ETC__q125 =
	      CASE_guard12299_0b0_NOT_iFifoD_OUT_BIT_103_0b_ETC__q124;
      3'd1:
	  CASE_iFifoD_OUT_BITS_6_TO_4_0_CASE_guard12299_ETC__q125 =
	      (guard__h212299 == 2'b0) ?
		!iFifo$D_OUT[103] :
		guard__h212299 != 2'b01 && guard__h212299 != 2'b10 &&
		guard__h212299 != 2'b11 ||
		!iFifo$D_OUT[103];
      3'd2, 3'd3:
	  CASE_iFifoD_OUT_BITS_6_TO_4_0_CASE_guard12299_ETC__q125 =
	      !iFifo$D_OUT[103];
      default: CASE_iFifoD_OUT_BITS_6_TO_4_0_CASE_guard12299_ETC__q125 =
		   iFifo$D_OUT[6:4] != 3'd4 || !iFifo$D_OUT[103];
    endcase
  end
  always@(iFifo$D_OUT)
  begin
    case (iFifo$D_OUT[6:4])
      3'd0, 3'd1, 3'd2, 3'd3:
	  IF_iFifo_first__087_BITS_6_TO_4_118_EQ_0_191_O_ETC___d5348 =
	      !iFifo$D_OUT[103];
      default: IF_iFifo_first__087_BITS_6_TO_4_118_EQ_0_191_O_ETC___d5348 =
		   iFifo$D_OUT[6:4] != 3'd4 || !iFifo$D_OUT[103];
    endcase
  end
  always@(fpu_madd_fState_S8$D_OUT)
  begin
    case (fpu_madd_fState_S8$D_OUT[2:1])
      2'b0, 2'b01, 2'b10:
	  CASE_fpu_madd_fState_S8D_OUT_BITS_2_TO_1_0b0__ETC__q126 =
	      fpu_madd_fState_S8$D_OUT[66];
      2'd3:
	  CASE_fpu_madd_fState_S8D_OUT_BITS_2_TO_1_0b0__ETC__q126 =
	      fpu_madd_fState_S8$D_OUT[2:1] == 2'b11 &&
	      fpu_madd_fState_S8$D_OUT[66];
    endcase
  end
  always@(fpu_madd_fState_S8$D_OUT or
	  CASE_fpu_madd_fState_S8D_OUT_BITS_2_TO_1_0b0__ETC__q126)
  begin
    case (fpu_madd_fState_S8$D_OUT[70:68])
      3'd0:
	  CASE_fpu_madd_fState_S8D_OUT_BITS_70_TO_68_0__ETC__q127 =
	      CASE_fpu_madd_fState_S8D_OUT_BITS_2_TO_1_0b0__ETC__q126;
      3'd1:
	  CASE_fpu_madd_fState_S8D_OUT_BITS_70_TO_68_0__ETC__q127 =
	      (fpu_madd_fState_S8$D_OUT[2:1] == 2'b0) ?
		fpu_madd_fState_S8$D_OUT[66] :
		(fpu_madd_fState_S8$D_OUT[2:1] == 2'b01 ||
		 fpu_madd_fState_S8$D_OUT[2:1] == 2'b10 ||
		 fpu_madd_fState_S8$D_OUT[2:1] == 2'b11) &&
		fpu_madd_fState_S8$D_OUT[66];
      3'd2, 3'd3:
	  CASE_fpu_madd_fState_S8D_OUT_BITS_70_TO_68_0__ETC__q127 =
	      fpu_madd_fState_S8$D_OUT[66];
      default: CASE_fpu_madd_fState_S8D_OUT_BITS_70_TO_68_0__ETC__q127 =
		   fpu_madd_fState_S8$D_OUT[70:68] == 3'd4 &&
		   fpu_madd_fState_S8$D_OUT[66];
    endcase
  end
  always@(iFifo$D_OUT or
	  IF_iFifo_first__087_BIT_71_849_THEN_IF_iFifo_f_ETC___d4618 or
	  IF_iFifo_first__087_BIT_201_115_THEN_IF_iFifo__ETC___d3848 or
	  IF_iFifo_first__087_BIT_71_849_THEN_IF_iFifo_f_ETC___d4555)
  begin
    case (iFifo$D_OUT[3:0])
      4'd0, 4'd1:
	  IF_iFifo_first__087_BITS_3_TO_0_088_EQ_0_089_O_ETC___d4623 =
	      IF_iFifo_first__087_BIT_201_115_THEN_IF_iFifo__ETC___d3848;
      4'd5, 4'd7:
	  IF_iFifo_first__087_BITS_3_TO_0_088_EQ_0_089_O_ETC___d4623 =
	      IF_iFifo_first__087_BIT_71_849_THEN_IF_iFifo_f_ETC___d4555;
      4'd6:
	  IF_iFifo_first__087_BITS_3_TO_0_088_EQ_0_089_O_ETC___d4623 =
	      IF_iFifo_first__087_BIT_71_849_THEN_IF_iFifo_f_ETC___d4618;
      default: IF_iFifo_first__087_BITS_3_TO_0_088_EQ_0_089_O_ETC___d4623 =
		   IF_iFifo_first__087_BIT_71_849_THEN_IF_iFifo_f_ETC___d4618;
    endcase
  end
  always@(iFifo$D_OUT or
	  fpu_madd_fOperand_S0$FULL_N or
	  fpu_div_fOperands_S0$FULL_N or fpu_sqr_fOperand_S0$FULL_N)
  begin
    case (iFifo$D_OUT[3:0])
      4'd0, 4'd1, 4'd2, 4'd5, 4'd6, 4'd7:
	  IF_iFifo_first__087_BITS_3_TO_0_088_EQ_0_089_O_ETC___d3110 =
	      fpu_madd_fOperand_S0$FULL_N;
      4'd3:
	  IF_iFifo_first__087_BITS_3_TO_0_088_EQ_0_089_O_ETC___d3110 =
	      fpu_div_fOperands_S0$FULL_N;
      4'd4:
	  IF_iFifo_first__087_BITS_3_TO_0_088_EQ_0_089_O_ETC___d3110 =
	      fpu_sqr_fOperand_S0$FULL_N;
      default: IF_iFifo_first__087_BITS_3_TO_0_088_EQ_0_089_O_ETC___d3110 =
		   iFifo$D_OUT[3:0] != 4'd8 || fpu_madd_fOperand_S0$FULL_N;
    endcase
  end
  always@(fpu_madd_fState_S8$D_OUT or
	  IF_0b0_CONCAT_NOT_fpu_madd_fState_S8_first__96_ETC___d3065)
  begin
    case (fpu_madd_fState_S8$D_OUT[2:1])
      2'b0, 2'b01:
	  CASE_fpu_madd_fState_S8D_OUT_BITS_2_TO_1_0b0__ETC__q130 =
	      fpu_madd_fState_S8$D_OUT[65:3];
      2'b10:
	  CASE_fpu_madd_fState_S8D_OUT_BITS_2_TO_1_0b0__ETC__q130 =
	      fpu_madd_fState_S8$D_OUT[3] ?
		IF_0b0_CONCAT_NOT_fpu_madd_fState_S8_first__96_ETC___d3065 :
		fpu_madd_fState_S8$D_OUT[65:3];
      2'b11:
	  CASE_fpu_madd_fState_S8D_OUT_BITS_2_TO_1_0b0__ETC__q130 =
	      IF_0b0_CONCAT_NOT_fpu_madd_fState_S8_first__96_ETC___d3065;
    endcase
  end
  always@(fpu_madd_fState_S8$D_OUT or
	  IF_0b0_CONCAT_NOT_fpu_madd_fState_S8_first__96_ETC___d3065)
  begin
    case (fpu_madd_fState_S8$D_OUT[2:1])
      2'b0:
	  CASE_fpu_madd_fState_S8D_OUT_BITS_2_TO_1_0b0__ETC__q131 =
	      fpu_madd_fState_S8$D_OUT[65:3];
      2'b01, 2'b10, 2'b11:
	  CASE_fpu_madd_fState_S8D_OUT_BITS_2_TO_1_0b0__ETC__q131 =
	      IF_0b0_CONCAT_NOT_fpu_madd_fState_S8_first__96_ETC___d3065;
    endcase
  end
  always@(fpu_madd_fState_S8$D_OUT or
	  CASE_fpu_madd_fState_S8D_OUT_BITS_2_TO_1_0b0__ETC__q130 or
	  CASE_fpu_madd_fState_S8D_OUT_BITS_2_TO_1_0b0__ETC__q131 or
	  IF_0b0_CONCAT_NOT_fpu_madd_fState_S8_first__96_ETC___d3065)
  begin
    case (fpu_madd_fState_S8$D_OUT[70:68])
      3'd0:
	  CASE_fpu_madd_fState_S8D_OUT_BITS_70_TO_68_0__ETC__q132 =
	      CASE_fpu_madd_fState_S8D_OUT_BITS_2_TO_1_0b0__ETC__q130;
      3'd1:
	  CASE_fpu_madd_fState_S8D_OUT_BITS_70_TO_68_0__ETC__q132 =
	      CASE_fpu_madd_fState_S8D_OUT_BITS_2_TO_1_0b0__ETC__q131;
      3'd2:
	  CASE_fpu_madd_fState_S8D_OUT_BITS_70_TO_68_0__ETC__q132 =
	      (fpu_madd_fState_S8$D_OUT[2:1] == 2'b0 ||
	       fpu_madd_fState_S8$D_OUT[66]) ?
		fpu_madd_fState_S8$D_OUT[65:3] :
		IF_0b0_CONCAT_NOT_fpu_madd_fState_S8_first__96_ETC___d3065;
      3'd3:
	  CASE_fpu_madd_fState_S8D_OUT_BITS_70_TO_68_0__ETC__q132 =
	      (fpu_madd_fState_S8$D_OUT[2:1] == 2'b0) ?
		fpu_madd_fState_S8$D_OUT[65:3] :
		(fpu_madd_fState_S8$D_OUT[66] ?
		   IF_0b0_CONCAT_NOT_fpu_madd_fState_S8_first__96_ETC___d3065 :
		   fpu_madd_fState_S8$D_OUT[65:3]);
      3'd4:
	  CASE_fpu_madd_fState_S8D_OUT_BITS_70_TO_68_0__ETC__q132 =
	      fpu_madd_fState_S8$D_OUT[65:3];
      default: CASE_fpu_madd_fState_S8D_OUT_BITS_70_TO_68_0__ETC__q132 =
		   63'd0;
    endcase
  end
  always@(rmdFifo$D_OUT or resWire$wget)
  begin
    case (rmdFifo$D_OUT)
      3'd0, 3'd1: _theResult___fst_exp__h269595 = 8'd255;
      3'd2:
	  _theResult___fst_exp__h269595 = resWire$wget[68] ? 8'd254 : 8'd255;
      3'd3:
	  _theResult___fst_exp__h269595 = resWire$wget[68] ? 8'd255 : 8'd254;
      3'd4: _theResult___fst_exp__h269595 = 8'd254;
      default: _theResult___fst_exp__h269595 = 8'd0;
    endcase
  end
  always@(rmdFifo$D_OUT or resWire$wget)
  begin
    case (rmdFifo$D_OUT)
      3'd0, 3'd1: _theResult___fst_sfd__h269596 = 23'd0;
      3'd2:
	  _theResult___fst_sfd__h269596 =
	      resWire$wget[68] ? 23'd8388607 : 23'd0;
      3'd3:
	  _theResult___fst_sfd__h269596 =
	      resWire$wget[68] ? 23'd0 : 23'd8388607;
      3'd4: _theResult___fst_sfd__h269596 = 23'd8388607;
      default: _theResult___fst_sfd__h269596 = 23'd0;
    endcase
  end
  always@(guard__h269623 or resWire$wget)
  begin
    case (guard__h269623)
      2'b0, 2'b01, 2'b10:
	  CASE_guard69623_0b0_resWirewget_BIT_68_0b1_re_ETC__q144 =
	      resWire$wget[68];
      2'd3:
	  CASE_guard69623_0b0_resWirewget_BIT_68_0b1_re_ETC__q144 =
	      guard__h269623 == 2'b11 && resWire$wget[68];
    endcase
  end
  always@(rmdFifo$D_OUT or
	  resWire$wget or
	  CASE_guard69623_0b0_resWirewget_BIT_68_0b1_re_ETC__q144 or
	  guard__h269623)
  begin
    case (rmdFifo$D_OUT)
      3'd0:
	  IF_rmdFifo_first__778_EQ_0_779_THEN_IF_IF_IF_I_ETC___d6388 =
	      CASE_guard69623_0b0_resWirewget_BIT_68_0b1_re_ETC__q144;
      3'd1:
	  IF_rmdFifo_first__778_EQ_0_779_THEN_IF_IF_IF_I_ETC___d6388 =
	      (guard__h269623 == 2'b0) ?
		resWire$wget[68] :
		(guard__h269623 == 2'b01 || guard__h269623 == 2'b10 ||
		 guard__h269623 == 2'b11) &&
		resWire$wget[68];
      3'd2, 3'd3:
	  IF_rmdFifo_first__778_EQ_0_779_THEN_IF_IF_IF_I_ETC___d6388 =
	      resWire$wget[68];
      default: IF_rmdFifo_first__778_EQ_0_779_THEN_IF_IF_IF_I_ETC___d6388 =
		   rmdFifo$D_OUT == 3'd4 && resWire$wget[68];
    endcase
  end
  always@(guard__h269623 or resWire$wget)
  begin
    case (guard__h269623)
      2'b0, 2'b01, 2'b10:
	  CASE_guard69623_0b0_NOT_resWirewget_BIT_68_0b_ETC__q145 =
	      !resWire$wget[68];
      2'd3:
	  CASE_guard69623_0b0_NOT_resWirewget_BIT_68_0b_ETC__q145 =
	      guard__h269623 != 2'b11 || !resWire$wget[68];
    endcase
  end
  always@(rmdFifo$D_OUT or
	  resWire$wget or
	  CASE_guard69623_0b0_NOT_resWirewget_BIT_68_0b_ETC__q145 or
	  guard__h269623)
  begin
    case (rmdFifo$D_OUT)
      3'd0:
	  IF_rmdFifo_first__778_EQ_0_779_THEN_IF_IF_IF_I_ETC___d5823 =
	      CASE_guard69623_0b0_NOT_resWirewget_BIT_68_0b_ETC__q145;
      3'd1:
	  IF_rmdFifo_first__778_EQ_0_779_THEN_IF_IF_IF_I_ETC___d5823 =
	      (guard__h269623 == 2'b0) ?
		!resWire$wget[68] :
		guard__h269623 != 2'b01 && guard__h269623 != 2'b10 &&
		guard__h269623 != 2'b11 ||
		!resWire$wget[68];
      3'd2, 3'd3:
	  IF_rmdFifo_first__778_EQ_0_779_THEN_IF_IF_IF_I_ETC___d5823 =
	      !resWire$wget[68];
      default: IF_rmdFifo_first__778_EQ_0_779_THEN_IF_IF_IF_I_ETC___d5823 =
		   rmdFifo$D_OUT != 3'd4 || !resWire$wget[68];
    endcase
  end
  always@(guard__h278330 or resWire$wget)
  begin
    case (guard__h278330)
      2'b0, 2'b01, 2'b10:
	  CASE_guard78330_0b0_resWirewget_BIT_68_0b1_re_ETC__q146 =
	      resWire$wget[68];
      2'd3:
	  CASE_guard78330_0b0_resWirewget_BIT_68_0b1_re_ETC__q146 =
	      guard__h278330 == 2'b11 && resWire$wget[68];
    endcase
  end
  always@(rmdFifo$D_OUT or
	  resWire$wget or
	  CASE_guard78330_0b0_resWirewget_BIT_68_0b1_re_ETC__q146 or
	  guard__h278330)
  begin
    case (rmdFifo$D_OUT)
      3'd0:
	  IF_rmdFifo_first__778_EQ_0_779_THEN_IF_IF_IF_r_ETC___d6397 =
	      CASE_guard78330_0b0_resWirewget_BIT_68_0b1_re_ETC__q146;
      3'd1:
	  IF_rmdFifo_first__778_EQ_0_779_THEN_IF_IF_IF_r_ETC___d6397 =
	      (guard__h278330 == 2'b0) ?
		resWire$wget[68] :
		(guard__h278330 == 2'b01 || guard__h278330 == 2'b10 ||
		 guard__h278330 == 2'b11) &&
		resWire$wget[68];
      3'd2, 3'd3:
	  IF_rmdFifo_first__778_EQ_0_779_THEN_IF_IF_IF_r_ETC___d6397 =
	      resWire$wget[68];
      default: IF_rmdFifo_first__778_EQ_0_779_THEN_IF_IF_IF_r_ETC___d6397 =
		   rmdFifo$D_OUT == 3'd4 && resWire$wget[68];
    endcase
  end
  always@(guard__h278330 or resWire$wget)
  begin
    case (guard__h278330)
      2'b0, 2'b01, 2'b10:
	  CASE_guard78330_0b0_NOT_resWirewget_BIT_68_0b_ETC__q147 =
	      !resWire$wget[68];
      2'd3:
	  CASE_guard78330_0b0_NOT_resWirewget_BIT_68_0b_ETC__q147 =
	      guard__h278330 != 2'b11 || !resWire$wget[68];
    endcase
  end
  always@(rmdFifo$D_OUT or
	  resWire$wget or
	  CASE_guard78330_0b0_NOT_resWirewget_BIT_68_0b_ETC__q147 or
	  guard__h278330)
  begin
    case (rmdFifo$D_OUT)
      3'd0:
	  IF_rmdFifo_first__778_EQ_0_779_THEN_IF_IF_IF_r_ETC___d6023 =
	      CASE_guard78330_0b0_NOT_resWirewget_BIT_68_0b_ETC__q147;
      3'd1:
	  IF_rmdFifo_first__778_EQ_0_779_THEN_IF_IF_IF_r_ETC___d6023 =
	      (guard__h278330 == 2'b0) ?
		!resWire$wget[68] :
		guard__h278330 != 2'b01 && guard__h278330 != 2'b10 &&
		guard__h278330 != 2'b11 ||
		!resWire$wget[68];
      3'd2, 3'd3:
	  IF_rmdFifo_first__778_EQ_0_779_THEN_IF_IF_IF_r_ETC___d6023 =
	      !resWire$wget[68];
      default: IF_rmdFifo_first__778_EQ_0_779_THEN_IF_IF_IF_r_ETC___d6023 =
		   rmdFifo$D_OUT != 3'd4 || !resWire$wget[68];
    endcase
  end
  always@(guard__h287260 or resWire$wget)
  begin
    case (guard__h287260)
      2'b0, 2'b01, 2'b10:
	  CASE_guard87260_0b0_resWirewget_BIT_68_0b1_re_ETC__q148 =
	      resWire$wget[68];
      2'd3:
	  CASE_guard87260_0b0_resWirewget_BIT_68_0b1_re_ETC__q148 =
	      guard__h287260 == 2'b11 && resWire$wget[68];
    endcase
  end
  always@(rmdFifo$D_OUT or
	  resWire$wget or
	  CASE_guard87260_0b0_resWirewget_BIT_68_0b1_re_ETC__q148 or
	  guard__h287260)
  begin
    case (rmdFifo$D_OUT)
      3'd0:
	  IF_rmdFifo_first__778_EQ_0_779_THEN_IF_IF_IF_I_ETC___d6409 =
	      CASE_guard87260_0b0_resWirewget_BIT_68_0b1_re_ETC__q148;
      3'd1:
	  IF_rmdFifo_first__778_EQ_0_779_THEN_IF_IF_IF_I_ETC___d6409 =
	      (guard__h287260 == 2'b0) ?
		resWire$wget[68] :
		(guard__h287260 == 2'b01 || guard__h287260 == 2'b10 ||
		 guard__h287260 == 2'b11) &&
		resWire$wget[68];
      3'd2, 3'd3:
	  IF_rmdFifo_first__778_EQ_0_779_THEN_IF_IF_IF_I_ETC___d6409 =
	      resWire$wget[68];
      default: IF_rmdFifo_first__778_EQ_0_779_THEN_IF_IF_IF_I_ETC___d6409 =
		   rmdFifo$D_OUT == 3'd4 && resWire$wget[68];
    endcase
  end
  always@(guard__h287260 or resWire$wget)
  begin
    case (guard__h287260)
      2'b0, 2'b01, 2'b10:
	  CASE_guard87260_0b0_NOT_resWirewget_BIT_68_0b_ETC__q149 =
	      !resWire$wget[68];
      2'd3:
	  CASE_guard87260_0b0_NOT_resWirewget_BIT_68_0b_ETC__q149 =
	      guard__h287260 != 2'b11 || !resWire$wget[68];
    endcase
  end
  always@(rmdFifo$D_OUT or
	  resWire$wget or
	  CASE_guard87260_0b0_NOT_resWirewget_BIT_68_0b_ETC__q149 or
	  guard__h287260)
  begin
    case (rmdFifo$D_OUT)
      3'd0:
	  IF_rmdFifo_first__778_EQ_0_779_THEN_IF_IF_IF_I_ETC___d6324 =
	      CASE_guard87260_0b0_NOT_resWirewget_BIT_68_0b_ETC__q149;
      3'd1:
	  IF_rmdFifo_first__778_EQ_0_779_THEN_IF_IF_IF_I_ETC___d6324 =
	      (guard__h287260 == 2'b0) ?
		!resWire$wget[68] :
		guard__h287260 != 2'b01 && guard__h287260 != 2'b10 &&
		guard__h287260 != 2'b11 ||
		!resWire$wget[68];
      3'd2, 3'd3:
	  IF_rmdFifo_first__778_EQ_0_779_THEN_IF_IF_IF_I_ETC___d6324 =
	      !resWire$wget[68];
      default: IF_rmdFifo_first__778_EQ_0_779_THEN_IF_IF_IF_I_ETC___d6324 =
		   rmdFifo$D_OUT != 3'd4 || !resWire$wget[68];
    endcase
  end
  always@(guard__h296096 or resWire$wget)
  begin
    case (guard__h296096)
      2'b0, 2'b01, 2'b10:
	  CASE_guard96096_0b0_resWirewget_BIT_68_0b1_re_ETC__q150 =
	      resWire$wget[68];
      2'd3:
	  CASE_guard96096_0b0_resWirewget_BIT_68_0b1_re_ETC__q150 =
	      guard__h296096 == 2'b11 && resWire$wget[68];
    endcase
  end
  always@(rmdFifo$D_OUT or
	  resWire$wget or
	  CASE_guard96096_0b0_resWirewget_BIT_68_0b1_re_ETC__q150 or
	  guard__h296096)
  begin
    case (rmdFifo$D_OUT)
      3'd0:
	  IF_rmdFifo_first__778_EQ_0_779_THEN_IF_IF_IF_r_ETC___d6418 =
	      CASE_guard96096_0b0_resWirewget_BIT_68_0b1_re_ETC__q150;
      3'd1:
	  IF_rmdFifo_first__778_EQ_0_779_THEN_IF_IF_IF_r_ETC___d6418 =
	      (guard__h296096 == 2'b0) ?
		resWire$wget[68] :
		(guard__h296096 == 2'b01 || guard__h296096 == 2'b10 ||
		 guard__h296096 == 2'b11) &&
		resWire$wget[68];
      3'd2, 3'd3:
	  IF_rmdFifo_first__778_EQ_0_779_THEN_IF_IF_IF_r_ETC___d6418 =
	      resWire$wget[68];
      default: IF_rmdFifo_first__778_EQ_0_779_THEN_IF_IF_IF_r_ETC___d6418 =
		   rmdFifo$D_OUT == 3'd4 && resWire$wget[68];
    endcase
  end
  always@(guard__h296096 or resWire$wget)
  begin
    case (guard__h296096)
      2'b0, 2'b01, 2'b10:
	  CASE_guard96096_0b0_NOT_resWirewget_BIT_68_0b_ETC__q151 =
	      !resWire$wget[68];
      2'd3:
	  CASE_guard96096_0b0_NOT_resWirewget_BIT_68_0b_ETC__q151 =
	      guard__h296096 != 2'b11 || !resWire$wget[68];
    endcase
  end
  always@(rmdFifo$D_OUT or
	  resWire$wget or
	  CASE_guard96096_0b0_NOT_resWirewget_BIT_68_0b_ETC__q151 or
	  guard__h296096)
  begin
    case (rmdFifo$D_OUT)
      3'd0:
	  IF_rmdFifo_first__778_EQ_0_779_THEN_IF_IF_IF_r_ETC___d6373 =
	      CASE_guard96096_0b0_NOT_resWirewget_BIT_68_0b_ETC__q151;
      3'd1:
	  IF_rmdFifo_first__778_EQ_0_779_THEN_IF_IF_IF_r_ETC___d6373 =
	      (guard__h296096 == 2'b0) ?
		!resWire$wget[68] :
		guard__h296096 != 2'b01 && guard__h296096 != 2'b10 &&
		guard__h296096 != 2'b11 ||
		!resWire$wget[68];
      3'd2, 3'd3:
	  IF_rmdFifo_first__778_EQ_0_779_THEN_IF_IF_IF_r_ETC___d6373 =
	      !resWire$wget[68];
      default: IF_rmdFifo_first__778_EQ_0_779_THEN_IF_IF_IF_r_ETC___d6373 =
		   rmdFifo$D_OUT != 3'd4 || !resWire$wget[68];
    endcase
  end
  always@(rmdFifo$D_OUT or resWire$wget)
  begin
    case (rmdFifo$D_OUT)
      3'd0, 3'd1, 3'd2, 3'd3:
	  IF_rmdFifo_first__778_EQ_0_779_OR_rmdFifo_firs_ETC___d6400 =
	      resWire$wget[68];
      default: IF_rmdFifo_first__778_EQ_0_779_OR_rmdFifo_firs_ETC___d6400 =
		   rmdFifo$D_OUT == 3'd4 && resWire$wget[68];
    endcase
  end
  always@(rmdFifo$D_OUT or resWire$wget)
  begin
    case (rmdFifo$D_OUT)
      3'd0, 3'd1, 3'd2, 3'd3:
	  IF_rmdFifo_first__778_EQ_0_779_OR_rmdFifo_firs_ETC___d6028 =
	      !resWire$wget[68];
      default: IF_rmdFifo_first__778_EQ_0_779_OR_rmdFifo_firs_ETC___d6028 =
		   rmdFifo$D_OUT != 3'd4 || !resWire$wget[68];
    endcase
  end
  always@(guard__h278330 or
	  _theResult___fst_exp__h286378 or
	  out_exp__h286823 or _theResult___exp__h286820)
  begin
    case (guard__h278330)
      2'b0, 2'b01:
	  CASE_guard78330_0b0_theResult___fst_exp86378_0_ETC__q152 =
	      _theResult___fst_exp__h286378;
      2'b10:
	  CASE_guard78330_0b0_theResult___fst_exp86378_0_ETC__q152 =
	      out_exp__h286823;
      2'b11:
	  CASE_guard78330_0b0_theResult___fst_exp86378_0_ETC__q152 =
	      _theResult___exp__h286820;
    endcase
  end
  always@(guard__h278330 or
	  _theResult___fst_exp__h286378 or _theResult___exp__h286820)
  begin
    case (guard__h278330)
      2'b0:
	  CASE_guard78330_0b0_theResult___fst_exp86378_0_ETC__q153 =
	      _theResult___fst_exp__h286378;
      2'b01, 2'b10, 2'b11:
	  CASE_guard78330_0b0_theResult___fst_exp86378_0_ETC__q153 =
	      _theResult___exp__h286820;
    endcase
  end
  always@(rmdFifo$D_OUT or
	  CASE_guard78330_0b0_theResult___fst_exp86378_0_ETC__q152 or
	  CASE_guard78330_0b0_theResult___fst_exp86378_0_ETC__q153 or
	  IF_IF_IF_resWire_wget__410_BITS_67_TO_57_416_E_ETC___d6479 or
	  IF_IF_IF_resWire_wget__410_BITS_67_TO_57_416_E_ETC___d6481 or
	  _theResult___fst_exp__h286378)
  begin
    case (rmdFifo$D_OUT)
      3'd0:
	  _theResult___fst_exp__h286898 =
	      CASE_guard78330_0b0_theResult___fst_exp86378_0_ETC__q152;
      3'd1:
	  _theResult___fst_exp__h286898 =
	      CASE_guard78330_0b0_theResult___fst_exp86378_0_ETC__q153;
      3'd2:
	  _theResult___fst_exp__h286898 =
	      IF_IF_IF_resWire_wget__410_BITS_67_TO_57_416_E_ETC___d6479;
      3'd3:
	  _theResult___fst_exp__h286898 =
	      IF_IF_IF_resWire_wget__410_BITS_67_TO_57_416_E_ETC___d6481;
      3'd4: _theResult___fst_exp__h286898 = _theResult___fst_exp__h286378;
      default: _theResult___fst_exp__h286898 = 8'd0;
    endcase
  end
  always@(guard__h269623 or
	  _theResult___fst_exp__h277722 or
	  out_exp__h278241 or _theResult___exp__h278238)
  begin
    case (guard__h269623)
      2'b0, 2'b01:
	  CASE_guard69623_0b0_theResult___fst_exp77722_0_ETC__q154 =
	      _theResult___fst_exp__h277722;
      2'b10:
	  CASE_guard69623_0b0_theResult___fst_exp77722_0_ETC__q154 =
	      out_exp__h278241;
      2'b11:
	  CASE_guard69623_0b0_theResult___fst_exp77722_0_ETC__q154 =
	      _theResult___exp__h278238;
    endcase
  end
  always@(guard__h269623 or
	  _theResult___fst_exp__h277722 or _theResult___exp__h278238)
  begin
    case (guard__h269623)
      2'b0:
	  CASE_guard69623_0b0_theResult___fst_exp77722_0_ETC__q155 =
	      _theResult___fst_exp__h277722;
      2'b01, 2'b10, 2'b11:
	  CASE_guard69623_0b0_theResult___fst_exp77722_0_ETC__q155 =
	      _theResult___exp__h278238;
    endcase
  end
  always@(rmdFifo$D_OUT or
	  CASE_guard69623_0b0_theResult___fst_exp77722_0_ETC__q154 or
	  CASE_guard69623_0b0_theResult___fst_exp77722_0_ETC__q155 or
	  IF_IF_IF_IF_0b0_CONCAT_NOT_resWire_wget__410_B_ETC___d6448 or
	  IF_IF_IF_IF_0b0_CONCAT_NOT_resWire_wget__410_B_ETC___d6450 or
	  _theResult___fst_exp__h277722)
  begin
    case (rmdFifo$D_OUT)
      3'd0:
	  _theResult___fst_exp__h278316 =
	      CASE_guard69623_0b0_theResult___fst_exp77722_0_ETC__q154;
      3'd1:
	  _theResult___fst_exp__h278316 =
	      CASE_guard69623_0b0_theResult___fst_exp77722_0_ETC__q155;
      3'd2:
	  _theResult___fst_exp__h278316 =
	      IF_IF_IF_IF_0b0_CONCAT_NOT_resWire_wget__410_B_ETC___d6448;
      3'd3:
	  _theResult___fst_exp__h278316 =
	      IF_IF_IF_IF_0b0_CONCAT_NOT_resWire_wget__410_B_ETC___d6450;
      3'd4: _theResult___fst_exp__h278316 = _theResult___fst_exp__h277722;
      default: _theResult___fst_exp__h278316 = 8'd0;
    endcase
  end
  always@(guard__h287260 or
	  _theResult___fst_exp__h295488 or
	  out_exp__h296007 or _theResult___exp__h296004)
  begin
    case (guard__h287260)
      2'b0, 2'b01:
	  CASE_guard87260_0b0_theResult___fst_exp95488_0_ETC__q156 =
	      _theResult___fst_exp__h295488;
      2'b10:
	  CASE_guard87260_0b0_theResult___fst_exp95488_0_ETC__q156 =
	      out_exp__h296007;
      2'b11:
	  CASE_guard87260_0b0_theResult___fst_exp95488_0_ETC__q156 =
	      _theResult___exp__h296004;
    endcase
  end
  always@(guard__h287260 or
	  _theResult___fst_exp__h295488 or _theResult___exp__h296004)
  begin
    case (guard__h287260)
      2'b0:
	  CASE_guard87260_0b0_theResult___fst_exp95488_0_ETC__q157 =
	      _theResult___fst_exp__h295488;
      2'b01, 2'b10, 2'b11:
	  CASE_guard87260_0b0_theResult___fst_exp95488_0_ETC__q157 =
	      _theResult___exp__h296004;
    endcase
  end
  always@(rmdFifo$D_OUT or
	  CASE_guard87260_0b0_theResult___fst_exp95488_0_ETC__q156 or
	  CASE_guard87260_0b0_theResult___fst_exp95488_0_ETC__q157 or
	  IF_IF_IF_IF_3970_MINUS_SEXT_resWire_wget__410__ETC___d6518 or
	  IF_IF_IF_IF_3970_MINUS_SEXT_resWire_wget__410__ETC___d6520 or
	  _theResult___fst_exp__h295488)
  begin
    case (rmdFifo$D_OUT)
      3'd0:
	  _theResult___fst_exp__h296082 =
	      CASE_guard87260_0b0_theResult___fst_exp95488_0_ETC__q156;
      3'd1:
	  _theResult___fst_exp__h296082 =
	      CASE_guard87260_0b0_theResult___fst_exp95488_0_ETC__q157;
      3'd2:
	  _theResult___fst_exp__h296082 =
	      IF_IF_IF_IF_3970_MINUS_SEXT_resWire_wget__410__ETC___d6518;
      3'd3:
	  _theResult___fst_exp__h296082 =
	      IF_IF_IF_IF_3970_MINUS_SEXT_resWire_wget__410__ETC___d6520;
      3'd4: _theResult___fst_exp__h296082 = _theResult___fst_exp__h295488;
      default: _theResult___fst_exp__h296082 = 8'd0;
    endcase
  end
  always@(guard__h296096 or
	  _theResult___fst_exp__h304173 or
	  out_exp__h304643 or _theResult___exp__h304640)
  begin
    case (guard__h296096)
      2'b0, 2'b01:
	  CASE_guard96096_0b0_theResult___fst_exp04173_0_ETC__q158 =
	      _theResult___fst_exp__h304173;
      2'b10:
	  CASE_guard96096_0b0_theResult___fst_exp04173_0_ETC__q158 =
	      out_exp__h304643;
      2'b11:
	  CASE_guard96096_0b0_theResult___fst_exp04173_0_ETC__q158 =
	      _theResult___exp__h304640;
    endcase
  end
  always@(guard__h296096 or
	  _theResult___fst_exp__h304173 or _theResult___exp__h304640)
  begin
    case (guard__h296096)
      2'b0:
	  CASE_guard96096_0b0_theResult___fst_exp04173_0_ETC__q159 =
	      _theResult___fst_exp__h304173;
      2'b01, 2'b10, 2'b11:
	  CASE_guard96096_0b0_theResult___fst_exp04173_0_ETC__q159 =
	      _theResult___exp__h304640;
    endcase
  end
  always@(rmdFifo$D_OUT or
	  CASE_guard96096_0b0_theResult___fst_exp04173_0_ETC__q158 or
	  CASE_guard96096_0b0_theResult___fst_exp04173_0_ETC__q159 or
	  IF_IF_IF_resWire_wget__410_BITS_67_TO_57_416_E_ETC___d6549 or
	  IF_IF_IF_resWire_wget__410_BITS_67_TO_57_416_E_ETC___d6551 or
	  _theResult___fst_exp__h304173)
  begin
    case (rmdFifo$D_OUT)
      3'd0:
	  _theResult___fst_exp__h304718 =
	      CASE_guard96096_0b0_theResult___fst_exp04173_0_ETC__q158;
      3'd1:
	  _theResult___fst_exp__h304718 =
	      CASE_guard96096_0b0_theResult___fst_exp04173_0_ETC__q159;
      3'd2:
	  _theResult___fst_exp__h304718 =
	      IF_IF_IF_resWire_wget__410_BITS_67_TO_57_416_E_ETC___d6549;
      3'd3:
	  _theResult___fst_exp__h304718 =
	      IF_IF_IF_resWire_wget__410_BITS_67_TO_57_416_E_ETC___d6551;
      3'd4: _theResult___fst_exp__h304718 = _theResult___fst_exp__h304173;
      default: _theResult___fst_exp__h304718 = 8'd0;
    endcase
  end
  always@(guard__h278330 or
	  _theResult___snd__h286329 or
	  out_sfd__h286824 or _theResult___sfd__h286821)
  begin
    case (guard__h278330)
      2'b0, 2'b01:
	  CASE_guard78330_0b0_theResult___snd86329_BITS__ETC__q160 =
	      _theResult___snd__h286329[56:34];
      2'b10:
	  CASE_guard78330_0b0_theResult___snd86329_BITS__ETC__q160 =
	      out_sfd__h286824;
      2'b11:
	  CASE_guard78330_0b0_theResult___snd86329_BITS__ETC__q160 =
	      _theResult___sfd__h286821;
    endcase
  end
  always@(guard__h278330 or
	  _theResult___snd__h286329 or _theResult___sfd__h286821)
  begin
    case (guard__h278330)
      2'b0:
	  CASE_guard78330_0b0_theResult___snd86329_BITS__ETC__q161 =
	      _theResult___snd__h286329[56:34];
      2'b01, 2'b10, 2'b11:
	  CASE_guard78330_0b0_theResult___snd86329_BITS__ETC__q161 =
	      _theResult___sfd__h286821;
    endcase
  end
  always@(rmdFifo$D_OUT or
	  CASE_guard78330_0b0_theResult___snd86329_BITS__ETC__q160 or
	  CASE_guard78330_0b0_theResult___snd86329_BITS__ETC__q161 or
	  IF_IF_IF_resWire_wget__410_BITS_67_TO_57_416_E_ETC___d6595 or
	  IF_IF_IF_resWire_wget__410_BITS_67_TO_57_416_E_ETC___d6597 or
	  _theResult___snd__h286329)
  begin
    case (rmdFifo$D_OUT)
      3'd0:
	  _theResult___fst_sfd__h286899 =
	      CASE_guard78330_0b0_theResult___snd86329_BITS__ETC__q160;
      3'd1:
	  _theResult___fst_sfd__h286899 =
	      CASE_guard78330_0b0_theResult___snd86329_BITS__ETC__q161;
      3'd2:
	  _theResult___fst_sfd__h286899 =
	      IF_IF_IF_resWire_wget__410_BITS_67_TO_57_416_E_ETC___d6595;
      3'd3:
	  _theResult___fst_sfd__h286899 =
	      IF_IF_IF_resWire_wget__410_BITS_67_TO_57_416_E_ETC___d6597;
      3'd4: _theResult___fst_sfd__h286899 = _theResult___snd__h286329[56:34];
      default: _theResult___fst_sfd__h286899 = 23'd0;
    endcase
  end
  always@(guard__h269623 or
	  sfdin__h277716 or out_sfd__h278242 or _theResult___sfd__h278239)
  begin
    case (guard__h269623)
      2'b0, 2'b01:
	  CASE_guard69623_0b0_sfdin77716_BITS_56_TO_34_0_ETC__q162 =
	      sfdin__h277716[56:34];
      2'b10:
	  CASE_guard69623_0b0_sfdin77716_BITS_56_TO_34_0_ETC__q162 =
	      out_sfd__h278242;
      2'b11:
	  CASE_guard69623_0b0_sfdin77716_BITS_56_TO_34_0_ETC__q162 =
	      _theResult___sfd__h278239;
    endcase
  end
  always@(guard__h269623 or sfdin__h277716 or _theResult___sfd__h278239)
  begin
    case (guard__h269623)
      2'b0:
	  CASE_guard69623_0b0_sfdin77716_BITS_56_TO_34_0_ETC__q163 =
	      sfdin__h277716[56:34];
      2'b01, 2'b10, 2'b11:
	  CASE_guard69623_0b0_sfdin77716_BITS_56_TO_34_0_ETC__q163 =
	      _theResult___sfd__h278239;
    endcase
  end
  always@(rmdFifo$D_OUT or
	  CASE_guard69623_0b0_sfdin77716_BITS_56_TO_34_0_ETC__q162 or
	  CASE_guard69623_0b0_sfdin77716_BITS_56_TO_34_0_ETC__q163 or
	  IF_IF_IF_IF_0b0_CONCAT_NOT_resWire_wget__410_B_ETC___d6576 or
	  IF_IF_IF_IF_0b0_CONCAT_NOT_resWire_wget__410_B_ETC___d6578 or
	  sfdin__h277716)
  begin
    case (rmdFifo$D_OUT)
      3'd0:
	  _theResult___fst_sfd__h278317 =
	      CASE_guard69623_0b0_sfdin77716_BITS_56_TO_34_0_ETC__q162;
      3'd1:
	  _theResult___fst_sfd__h278317 =
	      CASE_guard69623_0b0_sfdin77716_BITS_56_TO_34_0_ETC__q163;
      3'd2:
	  _theResult___fst_sfd__h278317 =
	      IF_IF_IF_IF_0b0_CONCAT_NOT_resWire_wget__410_B_ETC___d6576;
      3'd3:
	  _theResult___fst_sfd__h278317 =
	      IF_IF_IF_IF_0b0_CONCAT_NOT_resWire_wget__410_B_ETC___d6578;
      3'd4: _theResult___fst_sfd__h278317 = sfdin__h277716[56:34];
      default: _theResult___fst_sfd__h278317 = 23'd0;
    endcase
  end
  always@(guard__h287260 or
	  sfdin__h295482 or out_sfd__h296008 or _theResult___sfd__h296005)
  begin
    case (guard__h287260)
      2'b0, 2'b01:
	  CASE_guard87260_0b0_sfdin95482_BITS_56_TO_34_0_ETC__q164 =
	      sfdin__h295482[56:34];
      2'b10:
	  CASE_guard87260_0b0_sfdin95482_BITS_56_TO_34_0_ETC__q164 =
	      out_sfd__h296008;
      2'b11:
	  CASE_guard87260_0b0_sfdin95482_BITS_56_TO_34_0_ETC__q164 =
	      _theResult___sfd__h296005;
    endcase
  end
  always@(guard__h287260 or sfdin__h295482 or _theResult___sfd__h296005)
  begin
    case (guard__h287260)
      2'b0:
	  CASE_guard87260_0b0_sfdin95482_BITS_56_TO_34_0_ETC__q165 =
	      sfdin__h295482[56:34];
      2'b01, 2'b10, 2'b11:
	  CASE_guard87260_0b0_sfdin95482_BITS_56_TO_34_0_ETC__q165 =
	      _theResult___sfd__h296005;
    endcase
  end
  always@(rmdFifo$D_OUT or
	  CASE_guard87260_0b0_sfdin95482_BITS_56_TO_34_0_ETC__q164 or
	  CASE_guard87260_0b0_sfdin95482_BITS_56_TO_34_0_ETC__q165 or
	  IF_IF_IF_IF_3970_MINUS_SEXT_resWire_wget__410__ETC___d6622 or
	  IF_IF_IF_IF_3970_MINUS_SEXT_resWire_wget__410__ETC___d6624 or
	  sfdin__h295482)
  begin
    case (rmdFifo$D_OUT)
      3'd0:
	  _theResult___fst_sfd__h296083 =
	      CASE_guard87260_0b0_sfdin95482_BITS_56_TO_34_0_ETC__q164;
      3'd1:
	  _theResult___fst_sfd__h296083 =
	      CASE_guard87260_0b0_sfdin95482_BITS_56_TO_34_0_ETC__q165;
      3'd2:
	  _theResult___fst_sfd__h296083 =
	      IF_IF_IF_IF_3970_MINUS_SEXT_resWire_wget__410__ETC___d6622;
      3'd3:
	  _theResult___fst_sfd__h296083 =
	      IF_IF_IF_IF_3970_MINUS_SEXT_resWire_wget__410__ETC___d6624;
      3'd4: _theResult___fst_sfd__h296083 = sfdin__h295482[56:34];
      default: _theResult___fst_sfd__h296083 = 23'd0;
    endcase
  end
  always@(guard__h296096 or
	  _theResult___snd__h304119 or
	  out_sfd__h304644 or _theResult___sfd__h304641)
  begin
    case (guard__h296096)
      2'b0, 2'b01:
	  CASE_guard96096_0b0_theResult___snd04119_BITS__ETC__q166 =
	      _theResult___snd__h304119[56:34];
      2'b10:
	  CASE_guard96096_0b0_theResult___snd04119_BITS__ETC__q166 =
	      out_sfd__h304644;
      2'b11:
	  CASE_guard96096_0b0_theResult___snd04119_BITS__ETC__q166 =
	      _theResult___sfd__h304641;
    endcase
  end
  always@(guard__h296096 or
	  _theResult___snd__h304119 or _theResult___sfd__h304641)
  begin
    case (guard__h296096)
      2'b0:
	  CASE_guard96096_0b0_theResult___snd04119_BITS__ETC__q167 =
	      _theResult___snd__h304119[56:34];
      2'b01, 2'b10, 2'b11:
	  CASE_guard96096_0b0_theResult___snd04119_BITS__ETC__q167 =
	      _theResult___sfd__h304641;
    endcase
  end
  always@(rmdFifo$D_OUT or
	  CASE_guard96096_0b0_theResult___snd04119_BITS__ETC__q166 or
	  CASE_guard96096_0b0_theResult___snd04119_BITS__ETC__q167 or
	  IF_IF_IF_resWire_wget__410_BITS_67_TO_57_416_E_ETC___d6641 or
	  IF_IF_IF_resWire_wget__410_BITS_67_TO_57_416_E_ETC___d6643 or
	  _theResult___snd__h304119)
  begin
    case (rmdFifo$D_OUT)
      3'd0:
	  _theResult___fst_sfd__h304719 =
	      CASE_guard96096_0b0_theResult___snd04119_BITS__ETC__q166;
      3'd1:
	  _theResult___fst_sfd__h304719 =
	      CASE_guard96096_0b0_theResult___snd04119_BITS__ETC__q167;
      3'd2:
	  _theResult___fst_sfd__h304719 =
	      IF_IF_IF_resWire_wget__410_BITS_67_TO_57_416_E_ETC___d6641;
      3'd3:
	  _theResult___fst_sfd__h304719 =
	      IF_IF_IF_resWire_wget__410_BITS_67_TO_57_416_E_ETC___d6643;
      3'd4: _theResult___fst_sfd__h304719 = _theResult___snd__h304119[56:34];
      default: _theResult___fst_sfd__h304719 = 23'd0;
    endcase
  end
  always@(fpu_div_fState_S4$D_OUT)
  begin
    case (fpu_div_fState_S4$D_OUT[68:66])
      3'd2, 3'd3:
	  CASE_fpu_div_fState_S4D_OUT_BITS_68_TO_66_2_f_ETC__q168 =
	      fpu_div_fState_S4$D_OUT[65];
      default: CASE_fpu_div_fState_S4D_OUT_BITS_68_TO_66_2_f_ETC__q168 =
		   fpu_div_fState_S4$D_OUT[68:66] == 3'd4 &&
		   fpu_div_fState_S4$D_OUT[65];
    endcase
  end
  always@(fpu_div_fState_S4$D_OUT or
	  IF_0b0_CONCAT_NOT_fpu_div_fState_S4_first__73__ETC___d910)
  begin
    case (fpu_div_fState_S4$D_OUT[68:66])
      3'd2:
	  CASE_fpu_div_fState_S4D_OUT_BITS_68_TO_66_2_I_ETC__q169 =
	      (fpu_div_fState_S4$D_OUT[1:0] == 2'b0 ||
	       fpu_div_fState_S4$D_OUT[65]) ?
		fpu_div_fState_S4$D_OUT[64:2] :
		IF_0b0_CONCAT_NOT_fpu_div_fState_S4_first__73__ETC___d910;
      3'd3:
	  CASE_fpu_div_fState_S4D_OUT_BITS_68_TO_66_2_I_ETC__q169 =
	      (fpu_div_fState_S4$D_OUT[1:0] == 2'b0) ?
		fpu_div_fState_S4$D_OUT[64:2] :
		(fpu_div_fState_S4$D_OUT[65] ?
		   IF_0b0_CONCAT_NOT_fpu_div_fState_S4_first__73__ETC___d910 :
		   fpu_div_fState_S4$D_OUT[64:2]);
      3'd4:
	  CASE_fpu_div_fState_S4D_OUT_BITS_68_TO_66_2_I_ETC__q169 =
	      fpu_div_fState_S4$D_OUT[64:2];
      default: CASE_fpu_div_fState_S4D_OUT_BITS_68_TO_66_2_I_ETC__q169 =
		   63'd0;
    endcase
  end
  always@(fpu_div_fState_S4$D_OUT)
  begin
    case (fpu_div_fState_S4$D_OUT[1:0])
      2'b0, 2'b01, 2'b10:
	  CASE_fpu_div_fState_S4D_OUT_BITS_1_TO_0_0b0_f_ETC__q170 =
	      fpu_div_fState_S4$D_OUT[65];
      2'd3:
	  CASE_fpu_div_fState_S4D_OUT_BITS_1_TO_0_0b0_f_ETC__q170 =
	      fpu_div_fState_S4$D_OUT[1:0] == 2'b11 &&
	      fpu_div_fState_S4$D_OUT[65];
    endcase
  end
  always@(fpu_div_fState_S4$D_OUT or
	  IF_0b0_CONCAT_NOT_fpu_div_fState_S4_first__73__ETC___d910)
  begin
    case (fpu_div_fState_S4$D_OUT[1:0])
      2'b0, 2'b01:
	  CASE_fpu_div_fState_S4D_OUT_BITS_1_TO_0_0b0_f_ETC__q171 =
	      fpu_div_fState_S4$D_OUT[64:2];
      2'b10:
	  CASE_fpu_div_fState_S4D_OUT_BITS_1_TO_0_0b0_f_ETC__q171 =
	      fpu_div_fState_S4$D_OUT[2] ?
		IF_0b0_CONCAT_NOT_fpu_div_fState_S4_first__73__ETC___d910 :
		fpu_div_fState_S4$D_OUT[64:2];
      2'b11:
	  CASE_fpu_div_fState_S4D_OUT_BITS_1_TO_0_0b0_f_ETC__q171 =
	      IF_0b0_CONCAT_NOT_fpu_div_fState_S4_first__73__ETC___d910;
    endcase
  end
  always@(fpu_div_fState_S4$D_OUT or
	  IF_0b0_CONCAT_NOT_fpu_div_fState_S4_first__73__ETC___d910)
  begin
    case (fpu_div_fState_S4$D_OUT[1:0])
      2'd0: CASE_fpu_div_fState_S4D_OUT_BITS_1_TO_0_0_0_0_ETC__q172 = 63'd0;
      2'b01, 2'b10, 2'b11:
	  CASE_fpu_div_fState_S4D_OUT_BITS_1_TO_0_0_0_0_ETC__q172 =
	      IF_0b0_CONCAT_NOT_fpu_div_fState_S4_first__73__ETC___d910;
    endcase
  end
  always@(fpu_div_fState_S4$D_OUT or
	  CASE_fpu_div_fState_S4D_OUT_BITS_68_TO_66_2_f_ETC__q168 or
	  CASE_fpu_div_fState_S4D_OUT_BITS_68_TO_66_2_I_ETC__q169 or
	  CASE_fpu_div_fState_S4D_OUT_BITS_1_TO_0_0b0_f_ETC__q170 or
	  CASE_fpu_div_fState_S4D_OUT_BITS_1_TO_0_0b0_f_ETC__q171 or
	  CASE_fpu_div_fState_S4D_OUT_BITS_1_TO_0_0_0_0_ETC__q172)
  begin
    case (fpu_div_fState_S4$D_OUT[68:66])
      3'd0:
	  CASE_fpu_div_fState_S4D_OUT_BITS_68_TO_66_0_C_ETC__q173 =
	      { CASE_fpu_div_fState_S4D_OUT_BITS_1_TO_0_0b0_f_ETC__q170,
		CASE_fpu_div_fState_S4D_OUT_BITS_1_TO_0_0b0_f_ETC__q171 };
      3'd1:
	  CASE_fpu_div_fState_S4D_OUT_BITS_68_TO_66_0_C_ETC__q173 =
	      (fpu_div_fState_S4$D_OUT[1:0] == 2'b0) ?
		fpu_div_fState_S4$D_OUT[65:2] :
		{ (fpu_div_fState_S4$D_OUT[1:0] == 2'b01 ||
		   fpu_div_fState_S4$D_OUT[1:0] == 2'b10 ||
		   fpu_div_fState_S4$D_OUT[1:0] == 2'b11) &&
		  fpu_div_fState_S4$D_OUT[65],
		  CASE_fpu_div_fState_S4D_OUT_BITS_1_TO_0_0_0_0_ETC__q172 };
      default: CASE_fpu_div_fState_S4D_OUT_BITS_68_TO_66_0_C_ETC__q173 =
		   { CASE_fpu_div_fState_S4D_OUT_BITS_68_TO_66_2_f_ETC__q168,
		     CASE_fpu_div_fState_S4D_OUT_BITS_68_TO_66_2_I_ETC__q169 };
    endcase
  end
  always@(fpu_div_fState_S3$D_OUT)
  begin
    case (fpu_div_fState_S3$D_OUT[124:122])
      3'd0, 3'd1, 3'd2, 3'd3:
	  CASE_fpu_div_fState_S3D_OUT_BITS_124_TO_122_0_ETC__q174 =
	      fpu_div_fState_S3$D_OUT[121];
      default: CASE_fpu_div_fState_S3D_OUT_BITS_124_TO_122_0_ETC__q174 =
		   fpu_div_fState_S3$D_OUT[124:122] == 3'd4 &&
		   fpu_div_fState_S3$D_OUT[121];
    endcase
  end
  always@(fpu_div_fState_S3$D_OUT)
  begin
    case (fpu_div_fState_S3$D_OUT[124:122])
      3'd0, 3'd1:
	  CASE_fpu_div_fState_S3D_OUT_BITS_124_TO_122_0_ETC__q175 =
	      63'h7FF0000000000000;
      3'd2:
	  CASE_fpu_div_fState_S3D_OUT_BITS_124_TO_122_0_ETC__q175 =
	      fpu_div_fState_S3$D_OUT[121] ?
		63'h7FEFFFFFFFFFFFFF :
		63'h7FF0000000000000;
      3'd3:
	  CASE_fpu_div_fState_S3D_OUT_BITS_124_TO_122_0_ETC__q175 =
	      fpu_div_fState_S3$D_OUT[121] ?
		63'h7FF0000000000000 :
		63'h7FEFFFFFFFFFFFFF;
      3'd4:
	  CASE_fpu_div_fState_S3D_OUT_BITS_124_TO_122_0_ETC__q175 =
	      63'h7FEFFFFFFFFFFFFF;
      default: CASE_fpu_div_fState_S3D_OUT_BITS_124_TO_122_0_ETC__q175 =
		   63'd0;
    endcase
  end
  always@(iFifo$D_OUT or
	  IF_iFifo_first__087_BIT_201_115_THEN_IF_iFifo__ETC___d3848 or
	  IF_iFifo_first__087_BIT_136_624_THEN_IF_iFifo__ETC___d5330 or
	  IF_iFifo_first__087_BITS_102_TO_95_625_EQ_255__ETC___d5378)
  begin
    case (iFifo$D_OUT[3:0])
      4'd0:
	  CASE_iFifoD_OUT_BITS_3_TO_0_0_IF_iFifo_first__ETC__q176 =
	      IF_iFifo_first__087_BIT_136_624_THEN_IF_iFifo__ETC___d5330;
      4'd1:
	  CASE_iFifoD_OUT_BITS_3_TO_0_0_IF_iFifo_first__ETC__q176 =
	      iFifo$D_OUT[136] ?
		IF_iFifo_first__087_BITS_102_TO_95_625_EQ_255__ETC___d5378 :
		{ iFifo$D_OUT[136] || !iFifo$D_OUT[135],
		  iFifo$D_OUT[134:72] };
      default: CASE_iFifoD_OUT_BITS_3_TO_0_0_IF_iFifo_first__ETC__q176 =
		   IF_iFifo_first__087_BIT_201_115_THEN_IF_iFifo__ETC___d3848;
    endcase
  end
  always@(iFifo$D_OUT or
	  IF_iFifo_first__087_BIT_136_624_THEN_IF_iFifo__ETC___d5330)
  begin
    case (iFifo$D_OUT[3:0])
      4'd0, 4'd1:
	  CASE_iFifoD_OUT_BITS_3_TO_0_0_460718241880001_ETC__q177 =
	      64'h3FF0000000000000;
      default: CASE_iFifoD_OUT_BITS_3_TO_0_0_460718241880001_ETC__q177 =
		   IF_iFifo_first__087_BIT_136_624_THEN_IF_iFifo__ETC___d5330;
    endcase
  end
  always@(fpu_sqr_fState_S4$D_OUT)
  begin
    case (fpu_sqr_fState_S4$D_OUT[68:66])
      3'd2, 3'd3:
	  CASE_fpu_sqr_fState_S4D_OUT_BITS_68_TO_66_2_f_ETC__q178 =
	      fpu_sqr_fState_S4$D_OUT[65];
      default: CASE_fpu_sqr_fState_S4D_OUT_BITS_68_TO_66_2_f_ETC__q178 =
		   fpu_sqr_fState_S4$D_OUT[68:66] == 3'd4 &&
		   fpu_sqr_fState_S4$D_OUT[65];
    endcase
  end
  always@(fpu_sqr_fState_S4$D_OUT or
	  IF_0b0_CONCAT_NOT_fpu_sqr_fState_S4_first__687_ETC___d1724)
  begin
    case (fpu_sqr_fState_S4$D_OUT[68:66])
      3'd2:
	  CASE_fpu_sqr_fState_S4D_OUT_BITS_68_TO_66_2_I_ETC__q179 =
	      (fpu_sqr_fState_S4$D_OUT[1:0] == 2'b0 ||
	       fpu_sqr_fState_S4$D_OUT[65]) ?
		fpu_sqr_fState_S4$D_OUT[64:2] :
		IF_0b0_CONCAT_NOT_fpu_sqr_fState_S4_first__687_ETC___d1724;
      3'd3:
	  CASE_fpu_sqr_fState_S4D_OUT_BITS_68_TO_66_2_I_ETC__q179 =
	      (fpu_sqr_fState_S4$D_OUT[1:0] == 2'b0) ?
		fpu_sqr_fState_S4$D_OUT[64:2] :
		(fpu_sqr_fState_S4$D_OUT[65] ?
		   IF_0b0_CONCAT_NOT_fpu_sqr_fState_S4_first__687_ETC___d1724 :
		   fpu_sqr_fState_S4$D_OUT[64:2]);
      3'd4:
	  CASE_fpu_sqr_fState_S4D_OUT_BITS_68_TO_66_2_I_ETC__q179 =
	      fpu_sqr_fState_S4$D_OUT[64:2];
      default: CASE_fpu_sqr_fState_S4D_OUT_BITS_68_TO_66_2_I_ETC__q179 =
		   63'd0;
    endcase
  end
  always@(fpu_sqr_fState_S4$D_OUT)
  begin
    case (fpu_sqr_fState_S4$D_OUT[1:0])
      2'b0, 2'b01, 2'b10:
	  CASE_fpu_sqr_fState_S4D_OUT_BITS_1_TO_0_0b0_f_ETC__q180 =
	      fpu_sqr_fState_S4$D_OUT[65];
      2'd3:
	  CASE_fpu_sqr_fState_S4D_OUT_BITS_1_TO_0_0b0_f_ETC__q180 =
	      fpu_sqr_fState_S4$D_OUT[1:0] == 2'b11 &&
	      fpu_sqr_fState_S4$D_OUT[65];
    endcase
  end
  always@(fpu_sqr_fState_S4$D_OUT or
	  IF_0b0_CONCAT_NOT_fpu_sqr_fState_S4_first__687_ETC___d1724)
  begin
    case (fpu_sqr_fState_S4$D_OUT[1:0])
      2'b0, 2'b01:
	  CASE_fpu_sqr_fState_S4D_OUT_BITS_1_TO_0_0b0_f_ETC__q181 =
	      fpu_sqr_fState_S4$D_OUT[64:2];
      2'b10:
	  CASE_fpu_sqr_fState_S4D_OUT_BITS_1_TO_0_0b0_f_ETC__q181 =
	      fpu_sqr_fState_S4$D_OUT[2] ?
		IF_0b0_CONCAT_NOT_fpu_sqr_fState_S4_first__687_ETC___d1724 :
		fpu_sqr_fState_S4$D_OUT[64:2];
      2'b11:
	  CASE_fpu_sqr_fState_S4D_OUT_BITS_1_TO_0_0b0_f_ETC__q181 =
	      IF_0b0_CONCAT_NOT_fpu_sqr_fState_S4_first__687_ETC___d1724;
    endcase
  end
  always@(fpu_sqr_fState_S4$D_OUT or
	  IF_0b0_CONCAT_NOT_fpu_sqr_fState_S4_first__687_ETC___d1724)
  begin
    case (fpu_sqr_fState_S4$D_OUT[1:0])
      2'd0: CASE_fpu_sqr_fState_S4D_OUT_BITS_1_TO_0_0_0_0_ETC__q182 = 63'd0;
      2'b01, 2'b10, 2'b11:
	  CASE_fpu_sqr_fState_S4D_OUT_BITS_1_TO_0_0_0_0_ETC__q182 =
	      IF_0b0_CONCAT_NOT_fpu_sqr_fState_S4_first__687_ETC___d1724;
    endcase
  end
  always@(fpu_sqr_fState_S4$D_OUT or
	  CASE_fpu_sqr_fState_S4D_OUT_BITS_68_TO_66_2_f_ETC__q178 or
	  CASE_fpu_sqr_fState_S4D_OUT_BITS_68_TO_66_2_I_ETC__q179 or
	  CASE_fpu_sqr_fState_S4D_OUT_BITS_1_TO_0_0b0_f_ETC__q180 or
	  CASE_fpu_sqr_fState_S4D_OUT_BITS_1_TO_0_0b0_f_ETC__q181 or
	  CASE_fpu_sqr_fState_S4D_OUT_BITS_1_TO_0_0_0_0_ETC__q182)
  begin
    case (fpu_sqr_fState_S4$D_OUT[68:66])
      3'd0:
	  CASE_fpu_sqr_fState_S4D_OUT_BITS_68_TO_66_0_C_ETC__q183 =
	      { CASE_fpu_sqr_fState_S4D_OUT_BITS_1_TO_0_0b0_f_ETC__q180,
		CASE_fpu_sqr_fState_S4D_OUT_BITS_1_TO_0_0b0_f_ETC__q181 };
      3'd1:
	  CASE_fpu_sqr_fState_S4D_OUT_BITS_68_TO_66_0_C_ETC__q183 =
	      (fpu_sqr_fState_S4$D_OUT[1:0] == 2'b0) ?
		fpu_sqr_fState_S4$D_OUT[65:2] :
		{ (fpu_sqr_fState_S4$D_OUT[1:0] == 2'b01 ||
		   fpu_sqr_fState_S4$D_OUT[1:0] == 2'b10 ||
		   fpu_sqr_fState_S4$D_OUT[1:0] == 2'b11) &&
		  fpu_sqr_fState_S4$D_OUT[65],
		  CASE_fpu_sqr_fState_S4D_OUT_BITS_1_TO_0_0_0_0_ETC__q182 };
      default: CASE_fpu_sqr_fState_S4D_OUT_BITS_68_TO_66_0_C_ETC__q183 =
		   { CASE_fpu_sqr_fState_S4D_OUT_BITS_68_TO_66_2_f_ETC__q178,
		     CASE_fpu_sqr_fState_S4D_OUT_BITS_68_TO_66_2_I_ETC__q179 };
    endcase
  end
  // handling of inlined registers
  always@(posedge CLK)
  begin
    if (RST_N == `BSV_RESET_VALUE)
      begin
        crg_done <= `BSV_ASSIGNMENT_DELAY 1'd0;
	crg_done_1 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	rg_busy <= `BSV_ASSIGNMENT_DELAY 1'd0;
	rg_busy_1 <= `BSV_ASSIGNMENT_DELAY 1'd0;
      end
    else
      begin
        if (crg_done$EN) crg_done <= `BSV_ASSIGNMENT_DELAY crg_done$D_IN;
	if (crg_done_1$EN)
	  crg_done_1 <= `BSV_ASSIGNMENT_DELAY crg_done_1$D_IN;
	if (rg_busy$EN) rg_busy <= `BSV_ASSIGNMENT_DELAY rg_busy$D_IN;
	if (rg_busy_1$EN) rg_busy_1 <= `BSV_ASSIGNMENT_DELAY rg_busy_1$D_IN;
      end
    if (rg_b$EN) rg_b <= `BSV_ASSIGNMENT_DELAY rg_b$D_IN;
    if (rg_d$EN) rg_d <= `BSV_ASSIGNMENT_DELAY rg_d$D_IN;
    if (rg_index$EN) rg_index <= `BSV_ASSIGNMENT_DELAY rg_index$D_IN;
    if (rg_index_1$EN) rg_index_1 <= `BSV_ASSIGNMENT_DELAY rg_index_1$D_IN;
    if (rg_q$EN) rg_q <= `BSV_ASSIGNMENT_DELAY rg_q$D_IN;
    if (rg_r$EN) rg_r <= `BSV_ASSIGNMENT_DELAY rg_r$D_IN;
    if (rg_r_1$EN) rg_r_1 <= `BSV_ASSIGNMENT_DELAY rg_r_1$D_IN;
    if (rg_res$EN) rg_res <= `BSV_ASSIGNMENT_DELAY rg_res$D_IN;
    if (rg_s$EN) rg_s <= `BSV_ASSIGNMENT_DELAY rg_s$D_IN;
  end
  // synopsys translate_off
  `ifdef BSV_NO_INITIAL_BLOCKS
  `else // not BSV_NO_INITIAL_BLOCKS
  initial
  begin
    crg_done = 1'h0;
    crg_done_1 = 1'h0;
    rg_b = 116'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
    rg_busy = 1'h0;
    rg_busy_1 = 1'h0;
    rg_d = 58'h2AAAAAAAAAAAAAA;
    rg_index = 6'h2A;
    rg_index_1 = 6'h2A;
    rg_q = 58'h2AAAAAAAAAAAAAA;
    rg_r = 116'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
    rg_r_1 = 116'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
    rg_res = 117'h0AAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
    rg_s = 116'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
  end
  `endif // BSV_NO_INITIAL_BLOCKS
  // synopsys translate_on
  // handling of system tasks
  // synopsys translate_off
  always@(negedge CLK)
  begin
    #0;
    if (RST_N != `BSV_RESET_VALUE)
      if (fpu_madd_fResult_S9$EMPTY_N && fpu_div_fResult_S5$EMPTY_N)
	$display("Error: \"../../src_Core/CPU/FPU.bsv\", line 152, column 15: (R0001)\n  Mutually exclusive rules (from the ME sets [RL_getResFromPipe] and\n  [RL_getResFromPipe_1] ) fired in the same clock cycle.\n");
    if (RST_N != `BSV_RESET_VALUE)
      if ((fpu_madd_fResult_S9$EMPTY_N || fpu_div_fResult_S5$EMPTY_N) &&
	  fpu_sqr_fResult_S5$EMPTY_N)
	$display("Error: \"../../src_Core/CPU/FPU.bsv\", line 152, column 15: (R0001)\n  Mutually exclusive rules (from the ME sets [RL_getResFromPipe,\n  RL_getResFromPipe_1] and [RL_getResFromPipe_2] ) fired in the same clock\n  cycle.\n");
  end
  // synopsys translate_on
endmodule