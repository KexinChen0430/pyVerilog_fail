module ecrc(
   sys_clk ,
   rst_n ,
   data_in ,
   enable_crc ,
   half_data ,
   rst_crc ,
   crc_out64 ,
   crc_out32
   ) ;
input                  sys_clk ;
input                  rst_n ;
input  [15:0]          data_in ;
input                  enable_crc ;
input                  half_data ;
input                  rst_crc ;
output [31:0]          crc_out64 ;
output [31:0]          crc_out32 ;
reg  [31:0]            ohb435d ;
reg  [31:0]            ira1aec ;
reg  [31:0]            epd764 ;
reg  [31:0]            nr6bb24 ;
reg  [31:0]            zk5d927 ;
reg  [63:0]            hbec93a ;
reg  [63:0]            bl649d6 ;
reg  [31:0]            ym24eb6 ;
reg  [31:0]            db275b0 ;
reg  [31:0]            pu3ad86 ;
reg  [31:0]            uvd6c32 ;
reg                    qib6195 ;
wire [7:0]             dbb0ca9 ;
wire [7:0]             ba8654f ;
wire [7:0]             ph32a7b ;
wire [7:0]             qv953de ;
wire [7:0]             ksa9ef5 ;
wire [7:0]             zx4f7a8 ;
wire [7:0]             dz7bd47 ;
wire [7:0]             aydea3e ;
wire [31:0]            crc_out64 ;
wire [31:0]            crc_out32 ;
reg [15 : 0] uvf7ec2;
reg mg8d12e;
reg xwf1091;
reg aa8848a;
reg [31 : 0] fa42450;
reg [31 : 0] ux12283;
reg [31 : 0] ph9141c;
reg [31 : 0] ep8a0e7;
reg [31 : 0] rt5073d;
reg [63 : 0] tw839ef;
reg [63 : 0] zz1cf7a;
reg [31 : 0] gbe7bd6;
reg [31 : 0] tj3deb5;
reg [31 : 0] cmef5af;
reg [31 : 0] mr7ad78;
reg wjd6bc4;
reg [7 : 0] jrb5e25;
reg [7 : 0] zzaf12f;
reg [7 : 0] me7897e;
reg [7 : 0] ykc4bf1;
reg [7 : 0] pu25f89;
reg [7 : 0] hq2fc4a;
reg [7 : 0] fn7e253;
reg [7 : 0] vif129f;
reg [2047:0] necf6c2;
wire [23:0] ld7b613;
localparam qgdb09f = 24,nrd84f8 = 32'hfdffd14b;
localparam [31:0] thc27c7 = nrd84f8;
localparam mt9f1ff = nrd84f8 & 4'hf;
localparam [11:0] fnc7fe5 = 'h7ff;
wire  [(1 << mt9f1ff)  -1:0] suff972;
reg    [qgdb09f-1:0] cme5c87;
reg [mt9f1ff-1:0] qg721c0 [0:1];
reg [mt9f1ff-1:0] ym8700c;
reg rv38061;
integer jcc030e;
integer vk1872;
always @(uvf7ec2 or fa42450) begin   hbec93a = uvf7ec2;   bl649d6 = {          tw839ef[56], tw839ef[57], tw839ef[58], tw839ef[59], tw839ef[60], tw839ef[61], tw839ef[62], tw839ef[63],          tw839ef[48], tw839ef[49], tw839ef[50], tw839ef[51], tw839ef[52], tw839ef[53], tw839ef[54], tw839ef[55],          tw839ef[40], tw839ef[41], tw839ef[42], tw839ef[43], tw839ef[44], tw839ef[45], tw839ef[46], tw839ef[47],          tw839ef[32], tw839ef[33], tw839ef[34], tw839ef[35], tw839ef[36], tw839ef[37], tw839ef[38], tw839ef[39],          tw839ef[24], tw839ef[25], tw839ef[26], tw839ef[27], tw839ef[28], tw839ef[29], tw839ef[30], tw839ef[31],          tw839ef[16], tw839ef[17], tw839ef[18], tw839ef[19], tw839ef[20], tw839ef[21], tw839ef[22], tw839ef[23],          tw839ef[8], tw839ef[9], tw839ef[10], tw839ef[11], tw839ef[12], tw839ef[13], tw839ef[14], tw839ef[15],          tw839ef[0], tw839ef[1], tw839ef[2], tw839ef[3], tw839ef[4], tw839ef[5], tw839ef[6], tw839ef[7]         } ;   ym24eb6 = fa42450;   epd764[0] = zz1cf7a[63] ^ zz1cf7a[61] ^ zz1cf7a[60] ^ zz1cf7a[58] ^ zz1cf7a[55] ^ zz1cf7a[54] ^ zz1cf7a[53] ^                  zz1cf7a[50] ^ zz1cf7a[48] ^ zz1cf7a[47] ^ zz1cf7a[45] ^ zz1cf7a[44] ^ zz1cf7a[37] ^ zz1cf7a[34] ^                  zz1cf7a[32] ^ zz1cf7a[31] ^ zz1cf7a[30] ^ zz1cf7a[29] ^ zz1cf7a[28] ^ zz1cf7a[26] ^ zz1cf7a[25] ^                  zz1cf7a[24] ^ zz1cf7a[16] ^ zz1cf7a[12] ^ zz1cf7a[10] ^ zz1cf7a[9] ^ zz1cf7a[6] ^ zz1cf7a[0] ^                  gbe7bd6[0] ^ gbe7bd6[2] ^ gbe7bd6[5] ^ gbe7bd6[12] ^ gbe7bd6[13] ^ gbe7bd6[15] ^ gbe7bd6[16] ^                  gbe7bd6[18] ^ gbe7bd6[21] ^ gbe7bd6[22] ^ gbe7bd6[23] ^ gbe7bd6[26] ^ gbe7bd6[28] ^ gbe7bd6[29] ^                  gbe7bd6[31];   epd764[1] = zz1cf7a[63] ^ zz1cf7a[62] ^ zz1cf7a[60] ^ zz1cf7a[59] ^ zz1cf7a[58] ^ zz1cf7a[56] ^ zz1cf7a[53] ^                  zz1cf7a[51] ^ zz1cf7a[50] ^ zz1cf7a[49] ^ zz1cf7a[47] ^ zz1cf7a[46] ^ zz1cf7a[44] ^ zz1cf7a[38] ^                  zz1cf7a[37] ^ zz1cf7a[35] ^ zz1cf7a[34] ^ zz1cf7a[33] ^ zz1cf7a[28] ^ zz1cf7a[27] ^ zz1cf7a[24] ^                  zz1cf7a[17] ^ zz1cf7a[16] ^ zz1cf7a[13] ^ zz1cf7a[12] ^ zz1cf7a[11] ^ zz1cf7a[9] ^ zz1cf7a[7] ^                  zz1cf7a[6] ^ zz1cf7a[1] ^ zz1cf7a[0] ^ gbe7bd6[1] ^ gbe7bd6[2] ^ gbe7bd6[3] ^ gbe7bd6[5] ^ gbe7bd6[6] ^                  gbe7bd6[12] ^ gbe7bd6[14] ^ gbe7bd6[15] ^ gbe7bd6[17] ^ gbe7bd6[18] ^ gbe7bd6[19] ^ gbe7bd6[21] ^                  gbe7bd6[24] ^ gbe7bd6[26] ^ gbe7bd6[27] ^ gbe7bd6[28] ^ gbe7bd6[30] ^ gbe7bd6[31];   epd764[2] = zz1cf7a[59] ^ zz1cf7a[58] ^ zz1cf7a[57] ^ zz1cf7a[55] ^ zz1cf7a[53] ^ zz1cf7a[52] ^ zz1cf7a[51] ^                  zz1cf7a[44] ^ zz1cf7a[39] ^ zz1cf7a[38] ^ zz1cf7a[37] ^ zz1cf7a[36] ^ zz1cf7a[35] ^ zz1cf7a[32] ^                  zz1cf7a[31] ^ zz1cf7a[30] ^ zz1cf7a[26] ^ zz1cf7a[24] ^ zz1cf7a[18] ^ zz1cf7a[17] ^ zz1cf7a[16] ^                  zz1cf7a[14] ^ zz1cf7a[13] ^ zz1cf7a[9] ^ zz1cf7a[8] ^ zz1cf7a[7] ^ zz1cf7a[6] ^ zz1cf7a[2] ^                  zz1cf7a[1] ^ zz1cf7a[0] ^ gbe7bd6[0] ^ gbe7bd6[3] ^ gbe7bd6[4] ^ gbe7bd6[5] ^ gbe7bd6[6] ^ gbe7bd6[7] ^                  gbe7bd6[12] ^ gbe7bd6[19] ^ gbe7bd6[20] ^ gbe7bd6[21] ^ gbe7bd6[23] ^ gbe7bd6[25] ^ gbe7bd6[26] ^                  gbe7bd6[27];   epd764[3] = zz1cf7a[60] ^ zz1cf7a[59] ^ zz1cf7a[58] ^ zz1cf7a[56] ^ zz1cf7a[54] ^ zz1cf7a[53] ^ zz1cf7a[52] ^                  zz1cf7a[45] ^ zz1cf7a[40] ^ zz1cf7a[39] ^ zz1cf7a[38] ^ zz1cf7a[37] ^ zz1cf7a[36] ^ zz1cf7a[33] ^                  zz1cf7a[32] ^ zz1cf7a[31] ^ zz1cf7a[27] ^ zz1cf7a[25] ^ zz1cf7a[19] ^ zz1cf7a[18] ^ zz1cf7a[17] ^                  zz1cf7a[15] ^ zz1cf7a[14] ^ zz1cf7a[10] ^ zz1cf7a[9] ^ zz1cf7a[8] ^ zz1cf7a[7] ^ zz1cf7a[3] ^                  zz1cf7a[2] ^ zz1cf7a[1] ^ gbe7bd6[0] ^ gbe7bd6[1] ^ gbe7bd6[4] ^ gbe7bd6[5] ^ gbe7bd6[6] ^ gbe7bd6[7] ^                  gbe7bd6[8] ^ gbe7bd6[13] ^ gbe7bd6[20] ^ gbe7bd6[21] ^ gbe7bd6[22] ^ gbe7bd6[24] ^ gbe7bd6[26] ^                  gbe7bd6[27] ^ gbe7bd6[28];   epd764[4] = zz1cf7a[63] ^ zz1cf7a[59] ^ zz1cf7a[58] ^ zz1cf7a[57] ^ zz1cf7a[50] ^ zz1cf7a[48] ^ zz1cf7a[47] ^                  zz1cf7a[46] ^ zz1cf7a[45] ^ zz1cf7a[44] ^ zz1cf7a[41] ^ zz1cf7a[40] ^ zz1cf7a[39] ^ zz1cf7a[38] ^                  zz1cf7a[33] ^ zz1cf7a[31] ^ zz1cf7a[30] ^ zz1cf7a[29] ^ zz1cf7a[25] ^ zz1cf7a[24] ^ zz1cf7a[20] ^                  zz1cf7a[19] ^ zz1cf7a[18] ^ zz1cf7a[15] ^ zz1cf7a[12] ^ zz1cf7a[11] ^ zz1cf7a[8] ^ zz1cf7a[6] ^                  zz1cf7a[4] ^ zz1cf7a[3] ^ zz1cf7a[2] ^ zz1cf7a[0] ^ gbe7bd6[1] ^ gbe7bd6[6] ^ gbe7bd6[7] ^ gbe7bd6[8] ^                  gbe7bd6[9] ^ gbe7bd6[12] ^ gbe7bd6[13] ^ gbe7bd6[14] ^ gbe7bd6[15] ^ gbe7bd6[16] ^ gbe7bd6[18] ^                  gbe7bd6[25] ^ gbe7bd6[26] ^ gbe7bd6[27] ^ gbe7bd6[31];   epd764[5] = zz1cf7a[63] ^ zz1cf7a[61] ^ zz1cf7a[59] ^ zz1cf7a[55] ^ zz1cf7a[54] ^ zz1cf7a[53] ^ zz1cf7a[51] ^                  zz1cf7a[50] ^ zz1cf7a[49] ^ zz1cf7a[46] ^ zz1cf7a[44] ^ zz1cf7a[42] ^ zz1cf7a[41] ^ zz1cf7a[40] ^                  zz1cf7a[39] ^ zz1cf7a[37] ^ zz1cf7a[29] ^ zz1cf7a[28] ^ zz1cf7a[24] ^ zz1cf7a[21] ^ zz1cf7a[20] ^                  zz1cf7a[19] ^ zz1cf7a[13] ^ zz1cf7a[10] ^ zz1cf7a[7] ^ zz1cf7a[6] ^ zz1cf7a[5] ^ zz1cf7a[4] ^                  zz1cf7a[3] ^ zz1cf7a[1] ^ zz1cf7a[0] ^ gbe7bd6[5] ^ gbe7bd6[7] ^ gbe7bd6[8] ^ gbe7bd6[9] ^ gbe7bd6[10] ^                  gbe7bd6[12] ^ gbe7bd6[14] ^ gbe7bd6[17] ^ gbe7bd6[18] ^ gbe7bd6[19] ^ gbe7bd6[21] ^ gbe7bd6[22] ^                  gbe7bd6[23] ^ gbe7bd6[27] ^ gbe7bd6[29] ^ gbe7bd6[31];   epd764[6] = zz1cf7a[62] ^ zz1cf7a[60] ^ zz1cf7a[56] ^ zz1cf7a[55] ^ zz1cf7a[54] ^ zz1cf7a[52] ^ zz1cf7a[51] ^                  zz1cf7a[50] ^ zz1cf7a[47] ^ zz1cf7a[45] ^ zz1cf7a[43] ^ zz1cf7a[42] ^ zz1cf7a[41] ^ zz1cf7a[40] ^                  zz1cf7a[38] ^ zz1cf7a[30] ^ zz1cf7a[29] ^ zz1cf7a[25] ^ zz1cf7a[22] ^ zz1cf7a[21] ^ zz1cf7a[20] ^                  zz1cf7a[14] ^ zz1cf7a[11] ^ zz1cf7a[8] ^ zz1cf7a[7] ^ zz1cf7a[6] ^ zz1cf7a[5] ^ zz1cf7a[4] ^                  zz1cf7a[2] ^ zz1cf7a[1] ^ gbe7bd6[6] ^ gbe7bd6[8] ^ gbe7bd6[9] ^ gbe7bd6[10] ^ gbe7bd6[11] ^                  gbe7bd6[13] ^ gbe7bd6[15] ^ gbe7bd6[18] ^ gbe7bd6[19] ^ gbe7bd6[20] ^ gbe7bd6[22] ^ gbe7bd6[23] ^                  gbe7bd6[24] ^ gbe7bd6[28] ^ gbe7bd6[30];   epd764[7] = zz1cf7a[60] ^ zz1cf7a[58] ^ zz1cf7a[57] ^ zz1cf7a[56] ^ zz1cf7a[54] ^ zz1cf7a[52] ^ zz1cf7a[51] ^                  zz1cf7a[50] ^ zz1cf7a[47] ^ zz1cf7a[46] ^ zz1cf7a[45] ^ zz1cf7a[43] ^ zz1cf7a[42] ^ zz1cf7a[41] ^                  zz1cf7a[39] ^ zz1cf7a[37] ^ zz1cf7a[34] ^ zz1cf7a[32] ^ zz1cf7a[29] ^ zz1cf7a[28] ^ zz1cf7a[25] ^                  zz1cf7a[24] ^ zz1cf7a[23] ^ zz1cf7a[22] ^ zz1cf7a[21] ^ zz1cf7a[16] ^ zz1cf7a[15] ^ zz1cf7a[10] ^                  zz1cf7a[8] ^ zz1cf7a[7] ^ zz1cf7a[5] ^ zz1cf7a[3] ^ zz1cf7a[2] ^ zz1cf7a[0] ^ gbe7bd6[0] ^ gbe7bd6[2] ^                  gbe7bd6[5] ^ gbe7bd6[7] ^ gbe7bd6[9] ^ gbe7bd6[10] ^ gbe7bd6[11] ^ gbe7bd6[13] ^ gbe7bd6[14] ^                  gbe7bd6[15] ^ gbe7bd6[18] ^ gbe7bd6[19] ^ gbe7bd6[20] ^ gbe7bd6[22] ^ gbe7bd6[24] ^ gbe7bd6[25] ^                  gbe7bd6[26] ^ gbe7bd6[28];   epd764[8] = zz1cf7a[63] ^ zz1cf7a[60] ^ zz1cf7a[59] ^ zz1cf7a[57] ^ zz1cf7a[54] ^ zz1cf7a[52] ^ zz1cf7a[51] ^                  zz1cf7a[50] ^ zz1cf7a[46] ^ zz1cf7a[45] ^ zz1cf7a[43] ^ zz1cf7a[42] ^ zz1cf7a[40] ^ zz1cf7a[38] ^                  zz1cf7a[37] ^ zz1cf7a[35] ^ zz1cf7a[34] ^ zz1cf7a[33] ^ zz1cf7a[32] ^ zz1cf7a[31] ^ zz1cf7a[28] ^                  zz1cf7a[23] ^ zz1cf7a[22] ^ zz1cf7a[17] ^ zz1cf7a[12] ^ zz1cf7a[11] ^ zz1cf7a[10] ^ zz1cf7a[8] ^                  zz1cf7a[4] ^ zz1cf7a[3] ^ zz1cf7a[1] ^ zz1cf7a[0] ^ gbe7bd6[0] ^ gbe7bd6[1] ^ gbe7bd6[2] ^ gbe7bd6[3] ^                  gbe7bd6[5] ^ gbe7bd6[6] ^ gbe7bd6[8] ^ gbe7bd6[10] ^ gbe7bd6[11] ^ gbe7bd6[13] ^ gbe7bd6[14] ^                  gbe7bd6[18] ^ gbe7bd6[19] ^ gbe7bd6[20] ^ gbe7bd6[22] ^ gbe7bd6[25] ^ gbe7bd6[27] ^ gbe7bd6[28] ^                  gbe7bd6[31];   epd764[9] = zz1cf7a[61] ^ zz1cf7a[60] ^ zz1cf7a[58] ^ zz1cf7a[55] ^ zz1cf7a[53] ^ zz1cf7a[52] ^ zz1cf7a[51] ^                  zz1cf7a[47] ^ zz1cf7a[46] ^ zz1cf7a[44] ^ zz1cf7a[43] ^ zz1cf7a[41] ^ zz1cf7a[39] ^ zz1cf7a[38] ^                  zz1cf7a[36] ^ zz1cf7a[35] ^ zz1cf7a[34] ^ zz1cf7a[33] ^
zz1cf7a[32] ^ zz1cf7a[29] ^ zz1cf7a[24] ^                  zz1cf7a[23] ^ zz1cf7a[18] ^ zz1cf7a[13] ^ zz1cf7a[12] ^ zz1cf7a[11] ^ zz1cf7a[9] ^ zz1cf7a[5] ^                  zz1cf7a[4] ^ zz1cf7a[2] ^ zz1cf7a[1] ^ gbe7bd6[0] ^ gbe7bd6[1] ^ gbe7bd6[2] ^ gbe7bd6[3] ^ gbe7bd6[4] ^                  gbe7bd6[6] ^ gbe7bd6[7] ^ gbe7bd6[9] ^ gbe7bd6[11] ^ gbe7bd6[12] ^ gbe7bd6[14] ^ gbe7bd6[15] ^                  gbe7bd6[19] ^ gbe7bd6[20] ^ gbe7bd6[21] ^ gbe7bd6[23] ^ gbe7bd6[26] ^ gbe7bd6[28] ^ gbe7bd6[29];   epd764[10] = zz1cf7a[63] ^ zz1cf7a[62] ^ zz1cf7a[60] ^ zz1cf7a[59] ^ zz1cf7a[58] ^ zz1cf7a[56] ^ zz1cf7a[55] ^                   zz1cf7a[52] ^ zz1cf7a[50] ^ zz1cf7a[42] ^ zz1cf7a[40] ^ zz1cf7a[39] ^ zz1cf7a[36] ^ zz1cf7a[35] ^                   zz1cf7a[33] ^ zz1cf7a[32] ^ zz1cf7a[31] ^ zz1cf7a[29] ^ zz1cf7a[28] ^ zz1cf7a[26] ^ zz1cf7a[19] ^                   zz1cf7a[16] ^ zz1cf7a[14] ^ zz1cf7a[13] ^ zz1cf7a[9] ^ zz1cf7a[5] ^ zz1cf7a[3] ^ zz1cf7a[2] ^                   zz1cf7a[0] ^ gbe7bd6[0] ^ gbe7bd6[1] ^ gbe7bd6[3] ^ gbe7bd6[4] ^ gbe7bd6[7] ^ gbe7bd6[8] ^ gbe7bd6[10] ^                   gbe7bd6[18] ^ gbe7bd6[20] ^ gbe7bd6[23] ^ gbe7bd6[24] ^ gbe7bd6[26] ^ gbe7bd6[27] ^ gbe7bd6[28] ^                   gbe7bd6[30] ^ gbe7bd6[31];   epd764[11] = zz1cf7a[59] ^ zz1cf7a[58] ^ zz1cf7a[57] ^ zz1cf7a[56] ^ zz1cf7a[55] ^ zz1cf7a[54] ^ zz1cf7a[51] ^                   zz1cf7a[50] ^ zz1cf7a[48] ^ zz1cf7a[47] ^ zz1cf7a[45] ^ zz1cf7a[44] ^ zz1cf7a[43] ^ zz1cf7a[41] ^                   zz1cf7a[40] ^ zz1cf7a[36] ^ zz1cf7a[33] ^ zz1cf7a[31] ^ zz1cf7a[28] ^ zz1cf7a[27] ^ zz1cf7a[26] ^                   zz1cf7a[25] ^ zz1cf7a[24] ^ zz1cf7a[20] ^ zz1cf7a[17] ^ zz1cf7a[16] ^ zz1cf7a[15] ^ zz1cf7a[14] ^                   zz1cf7a[12] ^ zz1cf7a[9] ^ zz1cf7a[4] ^ zz1cf7a[3] ^ zz1cf7a[1] ^ zz1cf7a[0] ^ gbe7bd6[1] ^ gbe7bd6[4] ^                   gbe7bd6[8] ^ gbe7bd6[9] ^ gbe7bd6[11] ^ gbe7bd6[12] ^ gbe7bd6[13] ^ gbe7bd6[15] ^ gbe7bd6[16] ^                   gbe7bd6[18] ^ gbe7bd6[19] ^ gbe7bd6[22] ^ gbe7bd6[23] ^ gbe7bd6[24] ^ gbe7bd6[25] ^ gbe7bd6[26] ^                   gbe7bd6[27];   epd764[12] = zz1cf7a[63] ^ zz1cf7a[61] ^ zz1cf7a[59] ^ zz1cf7a[57] ^ zz1cf7a[56] ^ zz1cf7a[54] ^ zz1cf7a[53] ^                   zz1cf7a[52] ^ zz1cf7a[51] ^ zz1cf7a[50] ^ zz1cf7a[49] ^ zz1cf7a[47] ^ zz1cf7a[46] ^ zz1cf7a[42] ^                   zz1cf7a[41] ^ zz1cf7a[31] ^ zz1cf7a[30] ^ zz1cf7a[27] ^ zz1cf7a[24] ^ zz1cf7a[21] ^ zz1cf7a[18] ^                   zz1cf7a[17] ^ zz1cf7a[15] ^ zz1cf7a[13] ^ zz1cf7a[12] ^ zz1cf7a[9] ^ zz1cf7a[6] ^ zz1cf7a[5] ^                   zz1cf7a[4] ^ zz1cf7a[2] ^ zz1cf7a[1] ^ zz1cf7a[0] ^ gbe7bd6[9] ^ gbe7bd6[10] ^ gbe7bd6[14] ^                   gbe7bd6[15] ^ gbe7bd6[17] ^ gbe7bd6[18] ^ gbe7bd6[19] ^ gbe7bd6[20] ^ gbe7bd6[21] ^ gbe7bd6[22] ^                   gbe7bd6[24] ^ gbe7bd6[25] ^ gbe7bd6[27] ^ gbe7bd6[29] ^ gbe7bd6[31];   epd764[13] = zz1cf7a[62] ^ zz1cf7a[60] ^ zz1cf7a[58] ^ zz1cf7a[57] ^ zz1cf7a[55] ^ zz1cf7a[54] ^ zz1cf7a[53] ^                   zz1cf7a[52] ^ zz1cf7a[51] ^ zz1cf7a[50] ^ zz1cf7a[48] ^ zz1cf7a[47] ^ zz1cf7a[43] ^ zz1cf7a[42] ^                   zz1cf7a[32] ^ zz1cf7a[31] ^ zz1cf7a[28] ^ zz1cf7a[25] ^ zz1cf7a[22] ^ zz1cf7a[19] ^ zz1cf7a[18] ^                   zz1cf7a[16] ^ zz1cf7a[14] ^ zz1cf7a[13] ^ zz1cf7a[10] ^ zz1cf7a[7] ^ zz1cf7a[6] ^ zz1cf7a[5] ^                   zz1cf7a[3] ^ zz1cf7a[2] ^ zz1cf7a[1] ^ gbe7bd6[0] ^ gbe7bd6[10] ^ gbe7bd6[11] ^ gbe7bd6[15] ^                   gbe7bd6[16] ^ gbe7bd6[18] ^ gbe7bd6[19] ^ gbe7bd6[20] ^ gbe7bd6[21] ^ gbe7bd6[22] ^ gbe7bd6[23] ^                   gbe7bd6[25] ^ gbe7bd6[26] ^ gbe7bd6[28] ^ gbe7bd6[30];   epd764[14] = zz1cf7a[63] ^ zz1cf7a[61] ^ zz1cf7a[59] ^ zz1cf7a[58] ^ zz1cf7a[56] ^ zz1cf7a[55] ^ zz1cf7a[54] ^                   zz1cf7a[53] ^ zz1cf7a[52] ^ zz1cf7a[51] ^ zz1cf7a[49] ^ zz1cf7a[48] ^ zz1cf7a[44] ^ zz1cf7a[43] ^                   zz1cf7a[33] ^ zz1cf7a[32] ^ zz1cf7a[29] ^ zz1cf7a[26] ^ zz1cf7a[23] ^ zz1cf7a[20] ^ zz1cf7a[19] ^                   zz1cf7a[17] ^ zz1cf7a[15] ^ zz1cf7a[14] ^ zz1cf7a[11] ^ zz1cf7a[8] ^ zz1cf7a[7] ^ zz1cf7a[6] ^                   zz1cf7a[4] ^ zz1cf7a[3] ^ zz1cf7a[2] ^ gbe7bd6[0] ^ gbe7bd6[1] ^ gbe7bd6[11] ^ gbe7bd6[12] ^                   gbe7bd6[16] ^ gbe7bd6[17] ^ gbe7bd6[19] ^ gbe7bd6[20] ^ gbe7bd6[21] ^ gbe7bd6[22] ^ gbe7bd6[23] ^                   gbe7bd6[24] ^ gbe7bd6[26] ^ gbe7bd6[27] ^ gbe7bd6[29] ^ gbe7bd6[31];   epd764[15] = zz1cf7a[62] ^ zz1cf7a[60] ^ zz1cf7a[59] ^ zz1cf7a[57] ^ zz1cf7a[56] ^ zz1cf7a[55] ^ zz1cf7a[54] ^                   zz1cf7a[53] ^ zz1cf7a[52] ^ zz1cf7a[50] ^ zz1cf7a[49] ^ zz1cf7a[45] ^ zz1cf7a[44] ^ zz1cf7a[34] ^                   zz1cf7a[33] ^ zz1cf7a[30] ^ zz1cf7a[27] ^ zz1cf7a[24] ^ zz1cf7a[21] ^ zz1cf7a[20] ^ zz1cf7a[18] ^                   zz1cf7a[16] ^ zz1cf7a[15] ^ zz1cf7a[12] ^ zz1cf7a[9] ^ zz1cf7a[8] ^ zz1cf7a[7] ^ zz1cf7a[5] ^                   zz1cf7a[4] ^ zz1cf7a[3] ^ gbe7bd6[1] ^ gbe7bd6[2] ^ gbe7bd6[12] ^ gbe7bd6[13] ^ gbe7bd6[17] ^                   gbe7bd6[18] ^ gbe7bd6[20] ^ gbe7bd6[21] ^ gbe7bd6[22] ^ gbe7bd6[23] ^ gbe7bd6[24] ^ gbe7bd6[25] ^                   gbe7bd6[27] ^ gbe7bd6[28] ^ gbe7bd6[30];   epd764[16] = zz1cf7a[57] ^ zz1cf7a[56] ^ zz1cf7a[51] ^ zz1cf7a[48] ^ zz1cf7a[47] ^ zz1cf7a[46] ^ zz1cf7a[44] ^                   zz1cf7a[37] ^ zz1cf7a[35] ^ zz1cf7a[32] ^ zz1cf7a[30] ^ zz1cf7a[29] ^ zz1cf7a[26] ^ zz1cf7a[24] ^                   zz1cf7a[22] ^ zz1cf7a[21] ^ zz1cf7a[19] ^ zz1cf7a[17] ^ zz1cf7a[13] ^ zz1cf7a[12] ^ zz1cf7a[8] ^                   zz1cf7a[5] ^ zz1cf7a[4] ^ zz1cf7a[0] ^ gbe7bd6[0] ^ gbe7bd6[3] ^ gbe7bd6[5] ^ gbe7bd6[12] ^ gbe7bd6[14] ^                   gbe7bd6[15] ^ gbe7bd6[16] ^ gbe7bd6[19] ^ gbe7bd6[24] ^ gbe7bd6[25];   epd764[17] = zz1cf7a[58] ^ zz1cf7a[57] ^ zz1cf7a[52] ^ zz1cf7a[49] ^ zz1cf7a[48] ^ zz1cf7a[47] ^ zz1cf7a[45] ^                   zz1cf7a[38] ^ zz1cf7a[36] ^ zz1cf7a[33] ^ zz1cf7a[31] ^ zz1cf7a[30] ^ zz1cf7a[27] ^ zz1cf7a[25] ^                   zz1cf7a[23] ^ zz1cf7a[22] ^ zz1cf7a[20] ^ zz1cf7a[18] ^ zz1cf7a[14] ^ zz1cf7a[13] ^ zz1cf7a[9] ^                   zz1cf7a[6] ^ zz1cf7a[5] ^ zz1cf7a[1] ^ gbe7bd6[1] ^ gbe7bd6[4] ^ gbe7bd6[6] ^ gbe7bd6[13] ^ gbe7bd6[15] ^                   gbe7bd6[16] ^ gbe7bd6[17] ^ gbe7bd6[20] ^ gbe7bd6[25] ^ gbe7bd6[26];   epd764[18] = zz1cf7a[59] ^ zz1cf7a[58] ^ zz1cf7a[53] ^ zz1cf7a[50] ^ zz1cf7a[49] ^ zz1cf7a[48] ^ zz1cf7a[46] ^                   zz1cf7a[39] ^ zz1cf7a[37] ^ zz1cf7a[34] ^ zz1cf7a[32] ^ zz1cf7a[31] ^ zz1cf7a[28] ^ zz1cf7a[26] ^                   zz1cf7a[24] ^ zz1cf7a[23] ^ zz1cf7a[21] ^ zz1cf7a[19] ^ zz1cf7a[15] ^ zz1cf7a[14] ^ zz1cf7a[10] ^                   zz1cf7a[7] ^ zz1cf7a[6] ^ zz1cf7a[2] ^ gbe7bd6[0] ^ gbe7bd6[2] ^ gbe7bd6[5] ^ gbe7bd6[7] ^ gbe7bd6[14] ^                   gbe7bd6[16] ^ gbe7bd6[17] ^ gbe7bd6[18] ^ gbe7bd6[21] ^ gbe7bd6[26] ^ gbe7bd6[27];   epd764[19] = zz1cf7a[60] ^ zz1cf7a[59] ^ zz1cf7a[54] ^ zz1cf7a[51] ^ zz1cf7a[50] ^ zz1cf7a[49] ^ zz1cf7a[47] ^                   zz1cf7a[40] ^ zz1cf7a[38] ^ zz1cf7a[35] ^ zz1cf7a[33] ^ zz1cf7a[32] ^ zz1cf7a[29] ^ zz1cf7a[27] ^                   zz1cf7a[25] ^ zz1cf7a[24] ^ zz1cf7a[22] ^ zz1cf7a[20] ^ zz1cf7a[16] ^ zz1cf7a[15] ^ zz1cf7a[11] ^                   zz1cf7a[8] ^ zz1cf7a[7] ^ zz1cf7a[3] ^ gbe7bd6[0] ^ gbe7bd6[1] ^ gbe7bd6[3] ^ gbe7bd6[6] ^ gbe7bd6[8] ^                   gbe7bd6[15] ^ gbe7bd6[17] ^ gbe7bd6[18] ^ gbe7bd6[19] ^ gbe7bd6[22] ^ gbe7bd6[27] ^ gbe7bd6[28];   epd764[20] = zz1cf7a[61] ^ zz1cf7a[60] ^ zz1cf7a[55] ^ zz1cf7a[52] ^ zz1cf7a[51] ^ zz1cf7a[50] ^ zz1cf7a[48] ^                   zz1cf7a[41] ^ zz1cf7a[39] ^ zz1cf7a[36] ^ zz1cf7a[34] ^ zz1cf7a[33] ^ zz1cf7a[30] ^ zz1cf7a[28] ^                   zz1cf7a[26] ^ zz1cf7a[25] ^ zz1cf7a[23] ^ zz1cf7a[21] ^ zz1cf7a[17] ^ zz1cf7a[16] ^ zz1cf7a[12] ^                   zz1cf7a[9] ^ zz1cf7a[8] ^ zz1cf7a[4] ^ gbe7bd6[1] ^ gbe7bd6[2] ^ gbe7bd6[4] ^ gbe7bd6[7] ^ gbe7bd6[9] ^                   gbe7bd6[16] ^ gbe7bd6[18] ^ gbe7bd6[19] ^ gbe7bd6[20] ^ gbe7bd6[23] ^ gbe7bd6[28] ^ gbe7bd6[29];   epd764[21] = zz1cf7a[62] ^ zz1cf7a[61] ^ zz1cf7a[56] ^ zz1cf7a[53] ^ zz1cf7a[52] ^ zz1cf7a[51] ^ zz1cf7a[49] ^                   zz1cf7a[42] ^ zz1cf7a[40] ^ zz1cf7a[37] ^ zz1cf7a[35] ^ zz1cf7a[34] ^ zz1cf7a[31] ^
 zz1cf7a[29] ^                   zz1cf7a[27] ^ zz1cf7a[26] ^ zz1cf7a[24] ^ zz1cf7a[22] ^ zz1cf7a[18] ^ zz1cf7a[17] ^ zz1cf7a[13] ^                   zz1cf7a[10] ^ zz1cf7a[9] ^ zz1cf7a[5] ^ gbe7bd6[2] ^ gbe7bd6[3] ^ gbe7bd6[5] ^ gbe7bd6[8] ^ gbe7bd6[10] ^                   gbe7bd6[17] ^ gbe7bd6[19] ^ gbe7bd6[20] ^ gbe7bd6[21] ^ gbe7bd6[24] ^ gbe7bd6[29] ^ gbe7bd6[30];   epd764[22] = zz1cf7a[62] ^ zz1cf7a[61] ^ zz1cf7a[60] ^ zz1cf7a[58] ^ zz1cf7a[57] ^ zz1cf7a[55] ^ zz1cf7a[52] ^                   zz1cf7a[48] ^ zz1cf7a[47] ^ zz1cf7a[45] ^ zz1cf7a[44] ^ zz1cf7a[43] ^ zz1cf7a[41] ^ zz1cf7a[38] ^                   zz1cf7a[37] ^ zz1cf7a[36] ^ zz1cf7a[35] ^ zz1cf7a[34] ^ zz1cf7a[31] ^ zz1cf7a[29] ^ zz1cf7a[27] ^                   zz1cf7a[26] ^ zz1cf7a[24] ^ zz1cf7a[23] ^ zz1cf7a[19] ^ zz1cf7a[18] ^ zz1cf7a[16] ^ zz1cf7a[14] ^                   zz1cf7a[12] ^ zz1cf7a[11] ^ zz1cf7a[9] ^ zz1cf7a[0] ^ gbe7bd6[2] ^ gbe7bd6[3] ^ gbe7bd6[4] ^                   gbe7bd6[5] ^ gbe7bd6[6] ^ gbe7bd6[9] ^ gbe7bd6[11] ^ gbe7bd6[12] ^ gbe7bd6[13] ^ gbe7bd6[15] ^                   gbe7bd6[16] ^ gbe7bd6[20] ^ gbe7bd6[23] ^ gbe7bd6[25] ^ gbe7bd6[26] ^ gbe7bd6[28] ^ gbe7bd6[29] ^                   gbe7bd6[30];   epd764[23] = zz1cf7a[62] ^ zz1cf7a[60] ^ zz1cf7a[59] ^ zz1cf7a[56] ^ zz1cf7a[55] ^ zz1cf7a[54] ^ zz1cf7a[50] ^                   zz1cf7a[49] ^ zz1cf7a[47] ^ zz1cf7a[46] ^ zz1cf7a[42] ^ zz1cf7a[39] ^ zz1cf7a[38] ^ zz1cf7a[36] ^                   zz1cf7a[35] ^ zz1cf7a[34] ^ zz1cf7a[31] ^ zz1cf7a[29] ^ zz1cf7a[27] ^ zz1cf7a[26] ^ zz1cf7a[20] ^                   zz1cf7a[19] ^ zz1cf7a[17] ^ zz1cf7a[16] ^ zz1cf7a[15] ^ zz1cf7a[13] ^ zz1cf7a[9] ^ zz1cf7a[6] ^                   zz1cf7a[1] ^ zz1cf7a[0] ^ gbe7bd6[2] ^ gbe7bd6[3] ^ gbe7bd6[4] ^ gbe7bd6[6] ^ gbe7bd6[7] ^ gbe7bd6[10] ^                   gbe7bd6[14] ^ gbe7bd6[15] ^ gbe7bd6[17] ^ gbe7bd6[18] ^ gbe7bd6[22] ^ gbe7bd6[23] ^ gbe7bd6[24] ^                   gbe7bd6[27] ^ gbe7bd6[28] ^ gbe7bd6[30];   epd764[24] = zz1cf7a[63] ^ zz1cf7a[61] ^ zz1cf7a[60] ^ zz1cf7a[57] ^ zz1cf7a[56] ^ zz1cf7a[55] ^ zz1cf7a[51] ^                   zz1cf7a[50] ^ zz1cf7a[48] ^ zz1cf7a[47] ^ zz1cf7a[43] ^ zz1cf7a[40] ^ zz1cf7a[39] ^ zz1cf7a[37] ^                   zz1cf7a[36] ^ zz1cf7a[35] ^ zz1cf7a[32] ^ zz1cf7a[30] ^ zz1cf7a[28] ^ zz1cf7a[27] ^ zz1cf7a[21] ^                   zz1cf7a[20] ^ zz1cf7a[18] ^ zz1cf7a[17] ^ zz1cf7a[16] ^ zz1cf7a[14] ^ zz1cf7a[10] ^ zz1cf7a[7] ^                   zz1cf7a[2] ^ zz1cf7a[1] ^ gbe7bd6[0] ^ gbe7bd6[3] ^ gbe7bd6[4] ^ gbe7bd6[5] ^ gbe7bd6[7] ^ gbe7bd6[8] ^                   gbe7bd6[11] ^ gbe7bd6[15] ^ gbe7bd6[16] ^ gbe7bd6[18] ^ gbe7bd6[19] ^ gbe7bd6[23] ^ gbe7bd6[24] ^                   gbe7bd6[25] ^ gbe7bd6[28] ^ gbe7bd6[29] ^ gbe7bd6[31];   epd764[25] = zz1cf7a[62] ^ zz1cf7a[61] ^ zz1cf7a[58] ^ zz1cf7a[57] ^ zz1cf7a[56] ^ zz1cf7a[52] ^ zz1cf7a[51] ^                   zz1cf7a[49] ^ zz1cf7a[48] ^ zz1cf7a[44] ^ zz1cf7a[41] ^ zz1cf7a[40] ^ zz1cf7a[38] ^ zz1cf7a[37] ^                   zz1cf7a[36] ^ zz1cf7a[33] ^ zz1cf7a[31] ^ zz1cf7a[29] ^ zz1cf7a[28] ^ zz1cf7a[22] ^ zz1cf7a[21] ^                   zz1cf7a[19] ^ zz1cf7a[18] ^ zz1cf7a[17] ^ zz1cf7a[15] ^ zz1cf7a[11] ^ zz1cf7a[8] ^ zz1cf7a[3] ^                   zz1cf7a[2] ^ gbe7bd6[1] ^ gbe7bd6[4] ^ gbe7bd6[5] ^ gbe7bd6[6] ^ gbe7bd6[8] ^ gbe7bd6[9] ^ gbe7bd6[12] ^                   gbe7bd6[16] ^ gbe7bd6[17] ^ gbe7bd6[19] ^ gbe7bd6[20] ^ gbe7bd6[24] ^ gbe7bd6[25] ^ gbe7bd6[26] ^                   gbe7bd6[29] ^ gbe7bd6[30];   epd764[26] = zz1cf7a[62] ^ zz1cf7a[61] ^ zz1cf7a[60] ^ zz1cf7a[59] ^ zz1cf7a[57] ^ zz1cf7a[55] ^ zz1cf7a[54] ^                   zz1cf7a[52] ^ zz1cf7a[49] ^ zz1cf7a[48] ^ zz1cf7a[47] ^ zz1cf7a[44] ^ zz1cf7a[42] ^ zz1cf7a[41] ^                   zz1cf7a[39] ^ zz1cf7a[38] ^ zz1cf7a[31] ^ zz1cf7a[28] ^ zz1cf7a[26] ^ zz1cf7a[25] ^ zz1cf7a[24] ^                   zz1cf7a[23] ^ zz1cf7a[22] ^ zz1cf7a[20] ^ zz1cf7a[19] ^ zz1cf7a[18] ^ zz1cf7a[10] ^ zz1cf7a[6] ^                   zz1cf7a[4] ^ zz1cf7a[3] ^ zz1cf7a[0] ^ gbe7bd6[6] ^ gbe7bd6[7] ^ gbe7bd6[9] ^ gbe7bd6[10] ^ gbe7bd6[12] ^                   gbe7bd6[15] ^ gbe7bd6[16] ^ gbe7bd6[17] ^ gbe7bd6[20] ^ gbe7bd6[22] ^ gbe7bd6[23] ^ gbe7bd6[25] ^                   gbe7bd6[27] ^ gbe7bd6[28] ^ gbe7bd6[29] ^ gbe7bd6[30];   epd764[27] = zz1cf7a[63] ^ zz1cf7a[62] ^ zz1cf7a[61] ^ zz1cf7a[60] ^ zz1cf7a[58] ^ zz1cf7a[56] ^ zz1cf7a[55] ^                   zz1cf7a[53] ^ zz1cf7a[50] ^ zz1cf7a[49] ^ zz1cf7a[48] ^ zz1cf7a[45] ^ zz1cf7a[43] ^ zz1cf7a[42] ^                   zz1cf7a[40] ^ zz1cf7a[39] ^ zz1cf7a[32] ^ zz1cf7a[29] ^ zz1cf7a[27] ^ zz1cf7a[26] ^ zz1cf7a[25] ^                   zz1cf7a[24] ^ zz1cf7a[23] ^ zz1cf7a[21] ^ zz1cf7a[20] ^ zz1cf7a[19] ^ zz1cf7a[11] ^ zz1cf7a[7] ^                   zz1cf7a[5] ^ zz1cf7a[4] ^ zz1cf7a[1] ^ gbe7bd6[0] ^ gbe7bd6[7] ^ gbe7bd6[8] ^ gbe7bd6[10] ^ gbe7bd6[11] ^                   gbe7bd6[13] ^ gbe7bd6[16] ^ gbe7bd6[17] ^ gbe7bd6[18] ^ gbe7bd6[21] ^ gbe7bd6[23] ^ gbe7bd6[24] ^                   gbe7bd6[26] ^ gbe7bd6[28] ^ gbe7bd6[29] ^ gbe7bd6[30] ^ gbe7bd6[31];   epd764[28] = zz1cf7a[63] ^ zz1cf7a[62] ^ zz1cf7a[61] ^ zz1cf7a[59] ^ zz1cf7a[57] ^ zz1cf7a[56] ^ zz1cf7a[54] ^                   zz1cf7a[51] ^ zz1cf7a[50] ^ zz1cf7a[49] ^ zz1cf7a[46] ^ zz1cf7a[44] ^ zz1cf7a[43] ^ zz1cf7a[41] ^                   zz1cf7a[40] ^ zz1cf7a[33] ^ zz1cf7a[30] ^ zz1cf7a[28] ^ zz1cf7a[27] ^ zz1cf7a[26] ^ zz1cf7a[25] ^                   zz1cf7a[24] ^ zz1cf7a[22] ^ zz1cf7a[21] ^ zz1cf7a[20] ^ zz1cf7a[12] ^ zz1cf7a[8] ^ zz1cf7a[6] ^                   zz1cf7a[5] ^ zz1cf7a[2] ^ gbe7bd6[1] ^ gbe7bd6[8] ^ gbe7bd6[9] ^ gbe7bd6[11] ^ gbe7bd6[12] ^                   gbe7bd6[14] ^ gbe7bd6[17] ^ gbe7bd6[18] ^ gbe7bd6[19] ^ gbe7bd6[22] ^ gbe7bd6[24] ^ gbe7bd6[25] ^                   gbe7bd6[27] ^ gbe7bd6[29] ^ gbe7bd6[30] ^ gbe7bd6[31];   epd764[29] = zz1cf7a[63] ^ zz1cf7a[62] ^ zz1cf7a[60] ^ zz1cf7a[58] ^ zz1cf7a[57] ^ zz1cf7a[55] ^ zz1cf7a[52] ^                   zz1cf7a[51] ^ zz1cf7a[50] ^ zz1cf7a[47] ^ zz1cf7a[45] ^ zz1cf7a[44] ^ zz1cf7a[42] ^ zz1cf7a[41] ^                   zz1cf7a[34] ^ zz1cf7a[31] ^ zz1cf7a[29] ^ zz1cf7a[28] ^ zz1cf7a[27] ^ zz1cf7a[26] ^ zz1cf7a[25] ^                   zz1cf7a[23] ^ zz1cf7a[22] ^ zz1cf7a[21] ^ zz1cf7a[13] ^ zz1cf7a[9] ^ zz1cf7a[7] ^ zz1cf7a[6] ^                   zz1cf7a[3] ^ gbe7bd6[2] ^ gbe7bd6[9] ^ gbe7bd6[10] ^ gbe7bd6[12] ^ gbe7bd6[13] ^ gbe7bd6[15] ^                   gbe7bd6[18] ^ gbe7bd6[19] ^ gbe7bd6[20] ^ gbe7bd6[23] ^ gbe7bd6[25] ^ gbe7bd6[26] ^ gbe7bd6[28] ^                   gbe7bd6[30] ^ gbe7bd6[31];   epd764[30] = zz1cf7a[63] ^ zz1cf7a[61] ^ zz1cf7a[59] ^ zz1cf7a[58] ^ zz1cf7a[56] ^ zz1cf7a[53] ^ zz1cf7a[52] ^                   zz1cf7a[51] ^ zz1cf7a[48] ^ zz1cf7a[46] ^ zz1cf7a[45] ^ zz1cf7a[43] ^ zz1cf7a[42] ^ zz1cf7a[35] ^                   zz1cf7a[32] ^ zz1cf7a[30] ^ zz1cf7a[29] ^ zz1cf7a[28] ^ zz1cf7a[27] ^ zz1cf7a[26] ^ zz1cf7a[24] ^                   zz1cf7a[23] ^ zz1cf7a[22] ^ zz1cf7a[14] ^ zz1cf7a[10] ^ zz1cf7a[8] ^ zz1cf7a[7] ^ zz1cf7a[4] ^                   gbe7bd6[0] ^ gbe7bd6[3] ^ gbe7bd6[10] ^ gbe7bd6[11] ^ gbe7bd6[13] ^ gbe7bd6[14] ^ gbe7bd6[16] ^                   gbe7bd6[19] ^ gbe7bd6[20] ^ gbe7bd6[21] ^ gbe7bd6[24] ^ gbe7bd6[26] ^ gbe7bd6[27] ^ gbe7bd6[29] ^                   gbe7bd6[31];   epd764[31] = zz1cf7a[62] ^ zz1cf7a[60] ^ zz1cf7a[59] ^ zz1cf7a[57] ^ zz1cf7a[54] ^ zz1cf7a[53] ^ zz1cf7a[52] ^                   zz1cf7a[49] ^ zz1cf7a[47] ^ zz1cf7a[46] ^ zz1cf7a[44] ^ zz1cf7a[43] ^ zz1cf7a[36] ^ zz1cf7a[33] ^                   zz1cf7a[31] ^ zz1cf7a[30] ^ zz1cf7a[29] ^ zz1cf7a[28] ^ zz1cf7a[27] ^ zz1cf7a[25] ^ zz1cf7a[24] ^                   zz1cf7a[23] ^ zz1cf7a[15] ^ zz1cf7a[11] ^ zz1cf7a[9] ^ zz1cf7a[8] ^ zz1cf7a[5] ^ gbe7bd6[1] ^                   gbe7bd6[4] ^ gbe7bd6[11] ^ gbe7bd6[12] ^ gbe7bd6[14] ^ gbe7bd6[15] ^ gbe7bd6[17] ^ gbe7bd6[20] ^                   gbe7bd6[21] ^ gbe7bd6[22] ^ gbe7bd6[25] ^ gbe7bd6[27] ^ gbe7bd6[28] ^ gbe7bd6[30];
end
always @(rt5073d or ux12283) begin   db275b0 = rt5073d;   pu3ad86 = {          tj3deb5[24], tj3deb5[25], tj3deb5[26], tj3deb5[27], tj3deb5[28], tj3deb5[29], tj3deb5[30], tj3deb5[31],          tj3deb5[16], tj3deb5[17], tj3deb5[18], tj3deb5[19], tj3deb5[20], tj3deb5[21], tj3deb5[22], tj3deb5[23],          tj3deb5[8], tj3deb5[9], tj3deb5[10], tj3deb5[11], tj3deb5[12], tj3deb5[13], tj3deb5[14], tj3deb5[15],          tj3deb5[0], tj3deb5[1], tj3deb5[2], tj3deb5[3], tj3deb5[4], tj3deb5[5], tj3deb5[6], tj3deb5[7]         } ;   uvd6c32 = ux12283;   nr6bb24[0] = cmef5af[31] ^ cmef5af[30] ^ cmef5af[29] ^ cmef5af[28] ^ cmef5af[26] ^ cmef5af[25] ^ cmef5af[24] ^                  cmef5af[16] ^ cmef5af[12] ^ cmef5af[10] ^ cmef5af[9] ^ cmef5af[6] ^ cmef5af[0] ^ mr7ad78[0] ^                  mr7ad78[6] ^ mr7ad78[9] ^ mr7ad78[10] ^ mr7ad78[12] ^ mr7ad78[16] ^ mr7ad78[24] ^ mr7ad78[25] ^                  mr7ad78[26] ^ mr7ad78[28] ^ mr7ad78[29] ^ mr7ad78[30] ^ mr7ad78[31];   nr6bb24[1] = cmef5af[28] ^ cmef5af[27] ^ cmef5af[24] ^ cmef5af[17] ^ cmef5af[16] ^ cmef5af[13] ^ cmef5af[12] ^                  cmef5af[11] ^ cmef5af[9] ^ cmef5af[7] ^ cmef5af[6] ^ cmef5af[1] ^ cmef5af[0] ^ mr7ad78[0] ^ mr7ad78[1] ^                  mr7ad78[6] ^ mr7ad78[7] ^ mr7ad78[9] ^ mr7ad78[11] ^ mr7ad78[12] ^ mr7ad78[13] ^ mr7ad78[16] ^                  mr7ad78[17] ^ mr7ad78[24] ^ mr7ad78[27] ^ mr7ad78[28];   nr6bb24[2] = cmef5af[31] ^ cmef5af[30] ^ cmef5af[26] ^ cmef5af[24] ^ cmef5af[18] ^ cmef5af[17] ^ cmef5af[16] ^                  cmef5af[14] ^ cmef5af[13] ^ cmef5af[9] ^ cmef5af[8] ^ cmef5af[7] ^ cmef5af[6] ^ cmef5af[2] ^                  cmef5af[1] ^ cmef5af[0] ^ mr7ad78[0] ^ mr7ad78[1] ^ mr7ad78[2] ^ mr7ad78[6] ^ mr7ad78[7] ^ mr7ad78[8] ^                  mr7ad78[9] ^ mr7ad78[13] ^ mr7ad78[14] ^ mr7ad78[16] ^ mr7ad78[17] ^ mr7ad78[18] ^ mr7ad78[24] ^                  mr7ad78[26] ^ mr7ad78[30] ^ mr7ad78[31];   nr6bb24[3] = cmef5af[31] ^ cmef5af[27] ^ cmef5af[25] ^ cmef5af[19] ^ cmef5af[18] ^ cmef5af[17] ^ cmef5af[15] ^                  cmef5af[14] ^ cmef5af[10] ^ cmef5af[9] ^ cmef5af[8] ^ cmef5af[7] ^ cmef5af[3] ^ cmef5af[2] ^                  cmef5af[1] ^ mr7ad78[1] ^ mr7ad78[2] ^ mr7ad78[3] ^ mr7ad78[7] ^ mr7ad78[8] ^ mr7ad78[9] ^ mr7ad78[10] ^                  mr7ad78[14] ^ mr7ad78[15] ^ mr7ad78[17] ^ mr7ad78[18] ^ mr7ad78[19] ^ mr7ad78[25] ^ mr7ad78[27] ^                  mr7ad78[31];   nr6bb24[4] = cmef5af[31] ^ cmef5af[30] ^ cmef5af[29] ^ cmef5af[25] ^ cmef5af[24] ^ cmef5af[20] ^ cmef5af[19] ^                  cmef5af[18] ^ cmef5af[15] ^ cmef5af[12] ^ cmef5af[11] ^ cmef5af[8] ^ cmef5af[6] ^ cmef5af[4] ^                  cmef5af[3] ^ cmef5af[2] ^ cmef5af[0] ^ mr7ad78[0] ^ mr7ad78[2] ^ mr7ad78[3] ^ mr7ad78[4] ^ mr7ad78[6] ^                  mr7ad78[8] ^ mr7ad78[11] ^ mr7ad78[12] ^ mr7ad78[15] ^ mr7ad78[18] ^ mr7ad78[19] ^ mr7ad78[20] ^                  mr7ad78[24] ^ mr7ad78[25] ^ mr7ad78[29] ^ mr7ad78[30] ^ mr7ad78[31];   nr6bb24[5] = cmef5af[29] ^ cmef5af[28] ^ cmef5af[24] ^ cmef5af[21] ^ cmef5af[20] ^ cmef5af[19] ^ cmef5af[13] ^                  cmef5af[10] ^ cmef5af[7] ^ cmef5af[6] ^ cmef5af[5] ^ cmef5af[4] ^ cmef5af[3] ^ cmef5af[1] ^ cmef5af[0] ^                  mr7ad78[0] ^ mr7ad78[1] ^ mr7ad78[3] ^ mr7ad78[4] ^ mr7ad78[5] ^ mr7ad78[6] ^ mr7ad78[7] ^ mr7ad78[10] ^                  mr7ad78[13] ^ mr7ad78[19] ^ mr7ad78[20] ^ mr7ad78[21] ^ mr7ad78[24] ^ mr7ad78[28] ^ mr7ad78[29];   nr6bb24[6] = cmef5af[30] ^ cmef5af[29] ^ cmef5af[25] ^ cmef5af[22] ^ cmef5af[21] ^ cmef5af[20] ^ cmef5af[14] ^                  cmef5af[11] ^ cmef5af[8] ^ cmef5af[7] ^ cmef5af[6] ^ cmef5af[5] ^ cmef5af[4] ^ cmef5af[2] ^ cmef5af[1] ^                  mr7ad78[1] ^ mr7ad78[2] ^ mr7ad78[4] ^ mr7ad78[5] ^ mr7ad78[6] ^ mr7ad78[7] ^ mr7ad78[8] ^ mr7ad78[11] ^                  mr7ad78[14] ^ mr7ad78[20] ^ mr7ad78[21] ^ mr7ad78[22] ^ mr7ad78[25] ^ mr7ad78[29] ^ mr7ad78[30];   nr6bb24[7] = cmef5af[29] ^ cmef5af[28] ^ cmef5af[25] ^ cmef5af[24] ^ cmef5af[23] ^ cmef5af[22] ^ cmef5af[21] ^                  cmef5af[16] ^ cmef5af[15] ^ cmef5af[10] ^ cmef5af[8] ^ cmef5af[7] ^ cmef5af[5] ^ cmef5af[3] ^                  cmef5af[2] ^ cmef5af[0] ^ mr7ad78[0] ^ mr7ad78[2] ^ mr7ad78[3] ^ mr7ad78[5] ^ mr7ad78[7] ^ mr7ad78[8] ^                  mr7ad78[10] ^ mr7ad78[15] ^ mr7ad78[16] ^ mr7ad78[21] ^ mr7ad78[22] ^ mr7ad78[23] ^ mr7ad78[24] ^                  mr7ad78[25] ^ mr7ad78[28] ^ mr7ad78[29];   nr6bb24[8] = cmef5af[31] ^ cmef5af[28] ^ cmef5af[23] ^ cmef5af[22] ^ cmef5af[17] ^ cmef5af[12] ^ cmef5af[11] ^                  cmef5af[10] ^ cmef5af[8] ^ cmef5af[4] ^ cmef5af[3] ^ cmef5af[1] ^ cmef5af[0] ^ mr7ad78[0] ^ mr7ad78[1] ^                  mr7ad78[3] ^ mr7ad78[4] ^ mr7ad78[8] ^ mr7ad78[10] ^ mr7ad78[11] ^ mr7ad78[12] ^ mr7ad78[17] ^                  mr7ad78[22] ^ mr7ad78[23] ^ mr7ad78[28] ^ mr7ad78[31];   nr6bb24[9] = cmef5af[29] ^ cmef5af[24] ^ cmef5af[23] ^ cmef5af[18] ^ cmef5af[13] ^ cmef5af[12] ^ cmef5af[11] ^                  cmef5af[9] ^ cmef5af[5] ^ cmef5af[4] ^ cmef5af[2] ^ cmef5af[1] ^ mr7ad78[1] ^ mr7ad78[2] ^ mr7ad78[4] ^                  mr7ad78[5] ^ mr7ad78[9] ^ mr7ad78[11] ^ mr7ad78[12] ^ mr7ad78[13] ^ mr7ad78[18] ^ mr7ad78[23] ^                  mr7ad78[24] ^ mr7ad78[29];   nr6bb24[10] = cmef5af[31] ^ cmef5af[29] ^ cmef5af[28] ^ cmef5af[26] ^ cmef5af[19] ^ cmef5af[16] ^ cmef5af[14] ^                   cmef5af[13] ^ cmef5af[9] ^ cmef5af[5] ^ cmef5af[3] ^ cmef5af[2] ^ cmef5af[0] ^ mr7ad78[0] ^ mr7ad78[2] ^                   mr7ad78[3] ^ mr7ad78[5] ^ mr7ad78[9] ^ mr7ad78[13] ^ mr7ad78[14] ^ mr7ad78[16] ^ mr7ad78[19] ^                   mr7ad78[26] ^ mr7ad78[28] ^ mr7ad78[29] ^ mr7ad78[31];   nr6bb24[11] = cmef5af[31] ^ cmef5af[28] ^ cmef5af[27] ^ cmef5af[26] ^ cmef5af[25] ^ cmef5af[24] ^ cmef5af[20] ^                   cmef5af[17] ^ cmef5af[16] ^ cmef5af[15] ^ cmef5af[14] ^ cmef5af[12] ^ cmef5af[9] ^ cmef5af[4] ^                   cmef5af[3] ^ cmef5af[1] ^ cmef5af[0] ^ mr7ad78[0] ^ mr7ad78[1] ^ mr7ad78[3] ^ mr7ad78[4] ^ mr7ad78[9] ^                   mr7ad78[12] ^ mr7ad78[14] ^ mr7ad78[15] ^ mr7ad78[16] ^ mr7ad78[17] ^ mr7ad78[20] ^ mr7ad78[24] ^                   mr7ad78[25] ^ mr7ad78[26] ^ mr7ad78[27] ^ mr7ad78[28] ^ mr7ad78[31];   nr6bb24[12] = cmef5af[31] ^ cmef5af[30] ^ cmef5af[27] ^ cmef5af[24] ^ cmef5af[21] ^ cmef5af[18] ^ cmef5af[17] ^                   cmef5af[15] ^ cmef5af[13] ^ cmef5af[12] ^ cmef5af[9] ^ cmef5af[6] ^ cmef5af[5] ^ cmef5af[4] ^                   cmef5af[2] ^ cmef5af[1] ^ cmef5af[0] ^ mr7ad78[0] ^ mr7ad78[1] ^ mr7ad78[2] ^ mr7ad78[4] ^ mr7ad78[5] ^                   mr7ad78[6] ^ mr7ad78[9] ^ mr7ad78[12] ^ mr7ad78[13] ^ mr7ad78[15] ^ mr7ad78[17] ^ mr7ad78[18] ^                   mr7ad78[21] ^ mr7ad78[24] ^ mr7ad78[27] ^ mr7ad78[30] ^ mr7ad78[31];   nr6bb24[13] = cmef5af[31] ^ cmef5af[28] ^ cmef5af[25] ^ cmef5af[22] ^ cmef5af[19] ^ cmef5af[18] ^ cmef5af[16] ^                   cmef5af[14] ^ cmef5af[13] ^ cmef5af[10] ^ cmef5af[7] ^ cmef5af[6] ^ cmef5af[5] ^ cmef5af[3] ^                   cmef5af[2] ^ cmef5af[1] ^ mr7ad78[1] ^ mr7ad78[2] ^ mr7ad78[3] ^ mr7ad78[5] ^ mr7ad78[6] ^ mr7ad78[7] ^                   mr7ad78[10] ^ mr7ad78[13] ^ mr7ad78[14] ^ mr7ad78[16] ^ mr7ad78[18] ^ mr7ad78[19] ^ mr7ad78[22] ^                   mr7ad78[25] ^ mr7ad78[28] ^ mr7ad78[31];   nr6bb24[14] = cmef5af[29] ^ cmef5af[26] ^ cmef5af[23] ^ cmef5af[20] ^ cmef5af[19] ^ cmef5af[17] ^ cmef5af[15] ^                   cmef5af[14] ^ cmef5af[11] ^ cmef5af[8] ^ cmef5af[7] ^ cmef5af[6] ^ cmef5af[4] ^ cmef5af[3] ^                   cmef5af[2] ^ mr7ad78[2] ^ mr7ad78[3] ^ mr7ad78[4] ^ mr7ad78[6] ^ mr7ad78[7] ^ mr7ad78[8] ^ mr7ad78[11] ^                   mr7ad78[14] ^ mr7ad78[15] ^ mr7ad78[17] ^ mr7ad78[19] ^ mr7ad78[20] ^ mr7ad78[23] ^ mr7ad78[26] ^                   mr7ad78[29];   nr6bb24[15] = cmef5af[30] ^ cmef5af[27] ^ cmef5af[24] ^ cmef5af[21] ^ cmef5af[20] ^ cmef5af[18] ^ cmef5af[16] ^                   cmef5af[15] ^ cmef5af[12] ^ cmef5af[9] ^ cmef5af[8] ^ cmef5af[7] ^ cmef5af[5] ^ cmef5af[4] ^                   cmef5af[3] ^ mr7ad78[3] ^ mr7ad78[4] ^ mr7ad78[5] ^ mr7ad78[7] ^ mr7ad78[8] ^ mr7ad78[9] ^ mr7ad78[12] ^                   mr7ad78[15] ^ mr7ad78[16] ^ mr7ad78[18] ^ mr7ad78[20] ^ mr7ad78[21] ^
mr7ad78[24] ^ mr7ad78[27] ^                   mr7ad78[30];   nr6bb24[16] = cmef5af[30] ^ cmef5af[29] ^ cmef5af[26] ^ cmef5af[24] ^ cmef5af[22] ^ cmef5af[21] ^ cmef5af[19] ^                   cmef5af[17] ^ cmef5af[13] ^ cmef5af[12] ^ cmef5af[8] ^ cmef5af[5] ^ cmef5af[4] ^ cmef5af[0] ^                   mr7ad78[0] ^ mr7ad78[4] ^ mr7ad78[5] ^ mr7ad78[8] ^ mr7ad78[12] ^ mr7ad78[13] ^ mr7ad78[17] ^                   mr7ad78[19] ^ mr7ad78[21] ^ mr7ad78[22] ^ mr7ad78[24] ^ mr7ad78[26] ^ mr7ad78[29] ^ mr7ad78[30];   nr6bb24[17] = cmef5af[31] ^ cmef5af[30] ^ cmef5af[27] ^ cmef5af[25] ^ cmef5af[23] ^ cmef5af[22] ^ cmef5af[20] ^                   cmef5af[18] ^ cmef5af[14] ^ cmef5af[13] ^ cmef5af[9] ^ cmef5af[6] ^ cmef5af[5] ^ cmef5af[1] ^                   mr7ad78[1] ^ mr7ad78[5] ^ mr7ad78[6] ^ mr7ad78[9] ^ mr7ad78[13] ^ mr7ad78[14] ^ mr7ad78[18] ^                   mr7ad78[20] ^ mr7ad78[22] ^ mr7ad78[23] ^ mr7ad78[25] ^ mr7ad78[27] ^ mr7ad78[30] ^ mr7ad78[31];   nr6bb24[18] = cmef5af[31] ^ cmef5af[28] ^ cmef5af[26] ^ cmef5af[24] ^ cmef5af[23] ^ cmef5af[21] ^ cmef5af[19] ^                   cmef5af[15] ^ cmef5af[14] ^ cmef5af[10] ^ cmef5af[7] ^ cmef5af[6] ^ cmef5af[2] ^ mr7ad78[2] ^                   mr7ad78[6] ^ mr7ad78[7] ^ mr7ad78[10] ^ mr7ad78[14] ^ mr7ad78[15] ^ mr7ad78[19] ^ mr7ad78[21] ^                   mr7ad78[23] ^ mr7ad78[24] ^ mr7ad78[26] ^ mr7ad78[28] ^ mr7ad78[31];   nr6bb24[19] = cmef5af[29] ^ cmef5af[27] ^ cmef5af[25] ^ cmef5af[24] ^ cmef5af[22] ^ cmef5af[20] ^ cmef5af[16] ^                   cmef5af[15] ^ cmef5af[11] ^ cmef5af[8] ^ cmef5af[7] ^ cmef5af[3] ^ mr7ad78[3] ^ mr7ad78[7] ^                   mr7ad78[8] ^ mr7ad78[11] ^ mr7ad78[15] ^ mr7ad78[16] ^ mr7ad78[20] ^ mr7ad78[22] ^ mr7ad78[24] ^                   mr7ad78[25] ^ mr7ad78[27] ^ mr7ad78[29];   nr6bb24[20] = cmef5af[30] ^ cmef5af[28] ^ cmef5af[26] ^ cmef5af[25] ^ cmef5af[23] ^ cmef5af[21] ^ cmef5af[17] ^                   cmef5af[16] ^ cmef5af[12] ^ cmef5af[9] ^ cmef5af[8] ^ cmef5af[4] ^ mr7ad78[4] ^ mr7ad78[8] ^                   mr7ad78[9] ^ mr7ad78[12] ^ mr7ad78[16] ^ mr7ad78[17] ^ mr7ad78[21] ^ mr7ad78[23] ^ mr7ad78[25] ^                   mr7ad78[26] ^ mr7ad78[28] ^ mr7ad78[30];   nr6bb24[21] = cmef5af[31] ^ cmef5af[29] ^ cmef5af[27] ^ cmef5af[26] ^ cmef5af[24] ^ cmef5af[22] ^ cmef5af[18] ^                   cmef5af[17] ^ cmef5af[13] ^ cmef5af[10] ^ cmef5af[9] ^ cmef5af[5] ^ mr7ad78[5] ^ mr7ad78[9] ^                   mr7ad78[10] ^ mr7ad78[13] ^ mr7ad78[17] ^ mr7ad78[18] ^ mr7ad78[22] ^ mr7ad78[24] ^ mr7ad78[26] ^                   mr7ad78[27] ^ mr7ad78[29] ^ mr7ad78[31];   nr6bb24[22] = cmef5af[31] ^ cmef5af[29] ^ cmef5af[27] ^ cmef5af[26] ^ cmef5af[24] ^ cmef5af[23] ^ cmef5af[19] ^                   cmef5af[18] ^ cmef5af[16] ^ cmef5af[14] ^ cmef5af[12] ^ cmef5af[11] ^ cmef5af[9] ^ cmef5af[0] ^                   mr7ad78[0] ^ mr7ad78[9] ^ mr7ad78[11] ^ mr7ad78[12] ^ mr7ad78[14] ^ mr7ad78[16] ^ mr7ad78[18] ^                   mr7ad78[19] ^ mr7ad78[23] ^ mr7ad78[24] ^ mr7ad78[26] ^ mr7ad78[27] ^ mr7ad78[29] ^ mr7ad78[31];   nr6bb24[23] = cmef5af[31] ^ cmef5af[29] ^ cmef5af[27] ^ cmef5af[26] ^ cmef5af[20] ^ cmef5af[19] ^ cmef5af[17] ^                   cmef5af[16] ^ cmef5af[15] ^ cmef5af[13] ^ cmef5af[9] ^ cmef5af[6] ^ cmef5af[1] ^ cmef5af[0] ^                   mr7ad78[0] ^ mr7ad78[1] ^ mr7ad78[6] ^ mr7ad78[9] ^ mr7ad78[13] ^ mr7ad78[15] ^ mr7ad78[16] ^                   mr7ad78[17] ^ mr7ad78[19] ^ mr7ad78[20] ^ mr7ad78[26] ^ mr7ad78[27] ^ mr7ad78[29] ^ mr7ad78[31];   nr6bb24[24] = cmef5af[30] ^ cmef5af[28] ^ cmef5af[27] ^ cmef5af[21] ^ cmef5af[20] ^ cmef5af[18] ^ cmef5af[17] ^                   cmef5af[16] ^ cmef5af[14] ^ cmef5af[10] ^ cmef5af[7] ^ cmef5af[2] ^ cmef5af[1] ^ mr7ad78[1] ^                   mr7ad78[2] ^ mr7ad78[7] ^ mr7ad78[10] ^ mr7ad78[14] ^ mr7ad78[16] ^ mr7ad78[17] ^ mr7ad78[18] ^                   mr7ad78[20] ^ mr7ad78[21] ^ mr7ad78[27] ^ mr7ad78[28] ^ mr7ad78[30];   nr6bb24[25] = cmef5af[31] ^ cmef5af[29] ^ cmef5af[28] ^ cmef5af[22] ^ cmef5af[21] ^ cmef5af[19] ^ cmef5af[18] ^                   cmef5af[17] ^ cmef5af[15] ^ cmef5af[11] ^ cmef5af[8] ^ cmef5af[3] ^ cmef5af[2] ^ mr7ad78[2] ^                   mr7ad78[3] ^ mr7ad78[8] ^ mr7ad78[11] ^ mr7ad78[15] ^ mr7ad78[17] ^ mr7ad78[18] ^ mr7ad78[19] ^                   mr7ad78[21] ^ mr7ad78[22] ^ mr7ad78[28] ^ mr7ad78[29] ^ mr7ad78[31];   nr6bb24[26] = cmef5af[31] ^ cmef5af[28] ^ cmef5af[26] ^ cmef5af[25] ^ cmef5af[24] ^ cmef5af[23] ^ cmef5af[22] ^                   cmef5af[20] ^ cmef5af[19] ^ cmef5af[18] ^ cmef5af[10] ^ cmef5af[6] ^ cmef5af[4] ^ cmef5af[3] ^                   cmef5af[0] ^ mr7ad78[0] ^ mr7ad78[3] ^ mr7ad78[4] ^ mr7ad78[6] ^ mr7ad78[10] ^ mr7ad78[18] ^                   mr7ad78[19] ^ mr7ad78[20] ^ mr7ad78[22] ^ mr7ad78[23] ^ mr7ad78[24] ^ mr7ad78[25] ^ mr7ad78[26] ^                   mr7ad78[28] ^ mr7ad78[31];   nr6bb24[27] = cmef5af[29] ^ cmef5af[27] ^ cmef5af[26] ^ cmef5af[25] ^ cmef5af[24] ^ cmef5af[23] ^ cmef5af[21] ^                   cmef5af[20] ^ cmef5af[19] ^ cmef5af[11] ^ cmef5af[7] ^ cmef5af[5] ^ cmef5af[4] ^ cmef5af[1] ^                   mr7ad78[1] ^ mr7ad78[4] ^ mr7ad78[5] ^ mr7ad78[7] ^ mr7ad78[11] ^ mr7ad78[19] ^ mr7ad78[20] ^                   mr7ad78[21] ^ mr7ad78[23] ^ mr7ad78[24] ^ mr7ad78[25] ^ mr7ad78[26] ^ mr7ad78[27] ^ mr7ad78[29];   nr6bb24[28] = cmef5af[30] ^ cmef5af[28] ^ cmef5af[27] ^ cmef5af[26] ^ cmef5af[25] ^ cmef5af[24] ^ cmef5af[22] ^                   cmef5af[21] ^ cmef5af[20] ^ cmef5af[12] ^ cmef5af[8] ^ cmef5af[6] ^ cmef5af[5] ^ cmef5af[2] ^                   mr7ad78[2] ^ mr7ad78[5] ^ mr7ad78[6] ^ mr7ad78[8] ^ mr7ad78[12] ^ mr7ad78[20] ^ mr7ad78[21] ^                   mr7ad78[22] ^ mr7ad78[24] ^ mr7ad78[25] ^ mr7ad78[26] ^ mr7ad78[27] ^ mr7ad78[28] ^ mr7ad78[30];   nr6bb24[29] = cmef5af[31] ^ cmef5af[29] ^ cmef5af[28] ^ cmef5af[27] ^ cmef5af[26] ^ cmef5af[25] ^ cmef5af[23] ^                   cmef5af[22] ^ cmef5af[21] ^ cmef5af[13] ^ cmef5af[9] ^ cmef5af[7] ^ cmef5af[6] ^ cmef5af[3] ^                   mr7ad78[3] ^ mr7ad78[6] ^ mr7ad78[7] ^ mr7ad78[9] ^ mr7ad78[13] ^ mr7ad78[21] ^ mr7ad78[22] ^                   mr7ad78[23] ^ mr7ad78[25] ^ mr7ad78[26] ^ mr7ad78[27] ^ mr7ad78[28] ^ mr7ad78[29] ^ mr7ad78[31];   nr6bb24[30] = cmef5af[30] ^ cmef5af[29] ^ cmef5af[28] ^ cmef5af[27] ^ cmef5af[26] ^ cmef5af[24] ^ cmef5af[23] ^                   cmef5af[22] ^ cmef5af[14] ^ cmef5af[10] ^ cmef5af[8] ^ cmef5af[7] ^ cmef5af[4] ^ mr7ad78[4] ^                   mr7ad78[7] ^ mr7ad78[8] ^ mr7ad78[10] ^ mr7ad78[14] ^ mr7ad78[22] ^ mr7ad78[23] ^ mr7ad78[24] ^                   mr7ad78[26] ^ mr7ad78[27] ^ mr7ad78[28] ^ mr7ad78[29] ^ mr7ad78[30];   nr6bb24[31] = cmef5af[31] ^ cmef5af[30] ^ cmef5af[29] ^ cmef5af[28] ^ cmef5af[27] ^ cmef5af[25] ^ cmef5af[24] ^                   cmef5af[23] ^ cmef5af[15] ^ cmef5af[11] ^ cmef5af[9] ^ cmef5af[8] ^ cmef5af[5] ^ mr7ad78[5] ^                   mr7ad78[8] ^ mr7ad78[9] ^ mr7ad78[11] ^ mr7ad78[15] ^ mr7ad78[23] ^ mr7ad78[24] ^ mr7ad78[25] ^                   mr7ad78[27] ^ mr7ad78[28] ^ mr7ad78[29] ^ mr7ad78[30] ^ mr7ad78[31];
end
always @( posedge sys_clk or negedge rst_n ) begin   if (!rst_n)      ohb435d <= 32'hFFFF_FFFF ;   else if (aa8848a)      ohb435d <= 32'hFFFF_FFFF ;   else if (mg8d12e)      ohb435d <= ph9141c ;   else      ohb435d <= fa42450 ;
end
always @( posedge sys_clk or negedge rst_n ) begin   if (!rst_n)      ira1aec <= 32'h0000_0000 ;   else if (xwf1091)      ira1aec <= fa42450 ;   else if (wjd6bc4)      ira1aec <= ep8a0e7 ;   else            ira1aec <= ux12283 ;
end
always @( posedge sys_clk or negedge rst_n ) begin   if (!rst_n)      zk5d927 <= 32'h0000_0000 ;   else if (xwf1091)      zk5d927 <= uvf7ec2[63:32] ;   else      zk5d927 <= 32'h0000_0000 ;
end
always @( posedge sys_clk or negedge rst_n ) begin   if (!rst_n)      qib6195  <= 1'b0 ;   else      qib6195  <= xwf1091 ;
end
assign dbb0ca9 = { ~fa42450[24], ~fa42450[25], ~fa42450[26], ~fa42450[27],                        ~fa42450[28], ~fa42450[29], ~fa42450[30], ~fa42450[31] } ;
assign ba8654f = { ~fa42450[16], ~fa42450[17], ~fa42450[18], ~fa42450[19],                        ~fa42450[20], ~fa42450[21], ~fa42450[22], ~fa42450[23] } ;
assign ph32a7b = { ~fa42450[8], ~fa42450[9], ~fa42450[10], ~fa42450[11],                        ~fa42450[12], ~fa42450[13], ~fa42450[14], ~fa42450[15] } ;
assign qv953de = { ~fa42450[0], ~fa42450[1], ~fa42450[2], ~fa42450[3],                        ~fa42450[4], ~fa42450[5], ~fa42450[6], ~fa42450[7] } ;
assign ksa9ef5 = { ~ux12283[24], ~ux12283[25], ~ux12283[26], ~ux12283[27],                        ~ux12283[28], ~ux12283[29], ~ux12283[30], ~ux12283[31] } ;
assign zx4f7a8 = { ~ux12283[16], ~ux12283[17], ~ux12283[18], ~ux12283[19],                        ~ux12283[20], ~ux12283[21], ~ux12283[22], ~ux12283[23] } ;
assign dz7bd47 = { ~ux12283[8], ~ux12283[9], ~ux12283[10], ~ux12283[11],                        ~ux12283[12], ~ux12283[13], ~ux12283[14], ~ux12283[15] } ;
assign aydea3e = { ~ux12283[0], ~ux12283[1], ~ux12283[2], ~ux12283[3],                        ~ux12283[4], ~ux12283[5], ~ux12283[6], ~ux12283[7] } ;
assign crc_out64 = {jrb5e25, zzaf12f, me7897e, ykc4bf1} ;
assign crc_out32 = {pu25f89, hq2fc4a, fn7e253, vif129f} ;
always@* begin uvf7ec2<={data_in>>1,ld7b613[0]};mg8d12e<=ld7b613[1];xwf1091<=ld7b613[2];aa8848a<=ld7b613[3];fa42450<={ohb435d>>1,ld7b613[4]};ux12283<={ira1aec>>1,ld7b613[5]};ph9141c<={epd764>>1,ld7b613[6]};ep8a0e7<={nr6bb24>>1,ld7b613[7]};rt5073d<={zk5d927>>1,ld7b613[8]};tw839ef<={hbec93a>>1,ld7b613[9]};zz1cf7a<={bl649d6>>1,ld7b613[10]};gbe7bd6<={ym24eb6>>1,ld7b613[11]};tj3deb5<={db275b0>>1,ld7b613[12]};cmef5af<={pu3ad86>>1,ld7b613[13]};mr7ad78<={uvd6c32>>1,ld7b613[14]};wjd6bc4<=ld7b613[15];jrb5e25<={dbb0ca9>>1,ld7b613[16]};zzaf12f<={ba8654f>>1,ld7b613[17]};me7897e<={ph32a7b>>1,ld7b613[18]};ykc4bf1<={qv953de>>1,ld7b613[19]};pu25f89<={ksa9ef5>>1,ld7b613[20]};hq2fc4a<={zx4f7a8>>1,ld7b613[21]};fn7e253<={dz7bd47>>1,ld7b613[22]};vif129f<={aydea3e>>1,ld7b613[23]};end
always@* begin necf6c2[2047]<=enable_crc;necf6c2[2046]<=half_data;necf6c2[2044]<=rst_crc;necf6c2[2040]<=ohb435d[0];necf6c2[2033]<=ira1aec[0];necf6c2[2019]<=epd764[0];necf6c2[1990]<=nr6bb24[0];necf6c2[1939]<=ph32a7b[0];necf6c2[1933]<=zk5d927[0];necf6c2[1831]<=qv953de[0];necf6c2[1819]<=hbec93a[0];necf6c2[1778]<=qib6195;necf6c2[1615]<=ksa9ef5[0];necf6c2[1591]<=bl649d6[0];necf6c2[1508]<=dbb0ca9[0];necf6c2[1182]<=zx4f7a8[0];necf6c2[1135]<=ym24eb6[0];necf6c2[1023]<=data_in[0];necf6c2[969]<=ba8654f[0];necf6c2[889]<=uvd6c32[0];necf6c2[635]<=aydea3e[0];necf6c2[444]<=pu3ad86[0];necf6c2[317]<=dz7bd47[0];necf6c2[222]<=db275b0[0];end         assign suff972 = necf6c2,ld7b613 = cme5c87;   initial begin   jcc030e = $fopen(".fred");   $fdisplay( jcc030e, "%3h\n%3h", (thc27c7 >> 4) & fnc7fe5, (thc27c7 >> (mt9f1ff+4)) & fnc7fe5 );   $fclose(jcc030e);   $readmemh(".fred", qg721c0);   end   always @ (suff972) begin   ym8700c = qg721c0[1];       for (vk1872=0; vk1872<qgdb09f; vk1872=vk1872+1) begin           cme5c87[vk1872] = suff972[ym8700c];       rv38061  = ^(ym8700c & qg721c0[0]);       ym8700c =  {ym8700c, rv38061};       end   end
endmodule