module header
	// Internal signals
	// Generated Signal List
	// End of Generated Signal List
	// %COMPILER_OPTS%
	// Generated Signal Assignments
	// Generated Instances and Port Mappings
		// Generated Instance Port Map for inst_ea
		inst_ea_e inst_ea (
		);
		// End of Generated Instance Port Map for inst_ea
endmodule