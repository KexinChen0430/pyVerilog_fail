module not_a_bug315;
   typedef int supply_net_t;
   input int i;
   input imp_test_pkg::byte_t i;
   input supply_net_t bug316;
endmodule