module cla_adder(
	input [31:0] A,
	input [31:0] B,
	input Cin,
	output [31:0] Sum,
	output Cout
 );
	wire [31:0] a_plus_b_cin_0;
	wire [31:0] a_plus_b_cin_1;
	full_adder fa_00_cin_0
	full_adder fa_01_cin_0
	full_adder fa_02_cin_0
	full_adder fa_03_cin_0
	full_adder fa_00_cin_0
	full_adder fa_00_cin_0
	full_adder fa_00_cin_0
	full_adder fa_00_cin_0
	full_adder fa_00_cin_0
	full_adder fa_00_cin_0
	full_adder fa_00_cin_0
	full_adder fa_00_cin_0
	full_adder fa_00_cin_0
	full_adder fa_0_cin_0
	full_adder fa_0_cin_0
	full_adder fa_0_cin_0
	full_adder fa_0_cin_0
	full_adder fa_0_cin_0
	full_adder fa_0_cin_0
	full_adder fa_0_cin_0
	full_adder fa_0_cin_0
	full_adder fa_0_cin_0
	full_adder fa_0_cin_0
	full_adder fa_0_cin_0
	full_adder fa_0_cin_0
	full_adder fa_0_cin_0
	full_adder fa_0_cin_0
	full_adder fa_0_cin_0
	full_adder fa_0_cin_0
	full_adder fa_0_cin_0
	full_adder fa_0_cin_0
	full_adder fa_0_cin_0
	full_adder fa_0_cin_0
	full_adder fa_0_cin_0
	full_adder fa_0_cin_0
	full_adder fa_0_cin_0
	full_adder fa_0_cin_0
endmodule