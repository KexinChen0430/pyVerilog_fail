module's unterminated outputs)
   wire o_A_internal = 1'h0;
   wire o_A_outsideo = 1'h0;
   // End of automatics
endmodule