module VCU #(
`ifdef XIL_TIMING
  parameter LOC = "UNPLACED",
`endif
  parameter integer CORECLKREQ = 667,
  parameter integer DECHORRESOLUTION = 3840,
  parameter DECODERCHROMAFORMAT = "4_2_2",
  parameter DECODERCODING = "H.265",
  parameter integer DECODERCOLORDEPTH = 10,
  parameter integer DECODERNUMCORES = 2,
  parameter integer DECVERTRESOLUTION = 2160,
  parameter ENABLEDECODER = "TRUE",
  parameter ENABLEENCODER = "TRUE",
  parameter integer ENCHORRESOLUTION = 3840,
  parameter ENCODERCHROMAFORMAT = "4_2_2",
  parameter ENCODERCODING = "H.265",
  parameter integer ENCODERCOLORDEPTH = 10,
  parameter integer ENCODERNUMCORES = 4,
  parameter integer ENCVERTRESOLUTION = 2160
)(
  output VCUPLARREADYAXILITEAPB,
  output VCUPLAWREADYAXILITEAPB,
  output [1:0] VCUPLBRESPAXILITEAPB,
  output VCUPLBVALIDAXILITEAPB,
  output VCUPLCORESTATUSCLKPLL,
  output [43:0] VCUPLDECARADDR0,
  output [43:0] VCUPLDECARADDR1,
  output [1:0] VCUPLDECARBURST0,
  output [1:0] VCUPLDECARBURST1,
  output [3:0] VCUPLDECARCACHE0,
  output [3:0] VCUPLDECARCACHE1,
  output [3:0] VCUPLDECARID0,
  output [3:0] VCUPLDECARID1,
  output [7:0] VCUPLDECARLEN0,
  output [7:0] VCUPLDECARLEN1,
  output VCUPLDECARPROT0,
  output VCUPLDECARPROT1,
  output [3:0] VCUPLDECARQOS0,
  output [3:0] VCUPLDECARQOS1,
  output [2:0] VCUPLDECARSIZE0,
  output [2:0] VCUPLDECARSIZE1,
  output VCUPLDECARVALID0,
  output VCUPLDECARVALID1,
  output [43:0] VCUPLDECAWADDR0,
  output [43:0] VCUPLDECAWADDR1,
  output [1:0] VCUPLDECAWBURST0,
  output [1:0] VCUPLDECAWBURST1,
  output [3:0] VCUPLDECAWCACHE0,
  output [3:0] VCUPLDECAWCACHE1,
  output [3:0] VCUPLDECAWID0,
  output [3:0] VCUPLDECAWID1,
  output [7:0] VCUPLDECAWLEN0,
  output [7:0] VCUPLDECAWLEN1,
  output VCUPLDECAWPROT0,
  output VCUPLDECAWPROT1,
  output [3:0] VCUPLDECAWQOS0,
  output [3:0] VCUPLDECAWQOS1,
  output [2:0] VCUPLDECAWSIZE0,
  output [2:0] VCUPLDECAWSIZE1,
  output VCUPLDECAWVALID0,
  output VCUPLDECAWVALID1,
  output VCUPLDECBREADY0,
  output VCUPLDECBREADY1,
  output VCUPLDECRREADY0,
  output VCUPLDECRREADY1,
  output [127:0] VCUPLDECWDATA0,
  output [127:0] VCUPLDECWDATA1,
  output VCUPLDECWLAST0,
  output VCUPLDECWLAST1,
  output VCUPLDECWVALID0,
  output VCUPLDECWVALID1,
  output [16:0] VCUPLENCALL2CADDR,
  output VCUPLENCALL2CRVALID,
  output [319:0] VCUPLENCALL2CWDATA,
  output VCUPLENCALL2CWVALID,
  output [43:0] VCUPLENCARADDR0,
  output [43:0] VCUPLENCARADDR1,
  output [1:0] VCUPLENCARBURST0,
  output [1:0] VCUPLENCARBURST1,
  output [3:0] VCUPLENCARCACHE0,
  output [3:0] VCUPLENCARCACHE1,
  output [3:0] VCUPLENCARID0,
  output [3:0] VCUPLENCARID1,
  output [7:0] VCUPLENCARLEN0,
  output [7:0] VCUPLENCARLEN1,
  output VCUPLENCARPROT0,
  output VCUPLENCARPROT1,
  output [3:0] VCUPLENCARQOS0,
  output [3:0] VCUPLENCARQOS1,
  output [2:0] VCUPLENCARSIZE0,
  output [2:0] VCUPLENCARSIZE1,
  output VCUPLENCARVALID0,
  output VCUPLENCARVALID1,
  output [43:0] VCUPLENCAWADDR0,
  output [43:0] VCUPLENCAWADDR1,
  output [1:0] VCUPLENCAWBURST0,
  output [1:0] VCUPLENCAWBURST1,
  output [3:0] VCUPLENCAWCACHE0,
  output [3:0] VCUPLENCAWCACHE1,
  output [3:0] VCUPLENCAWID0,
  output [3:0] VCUPLENCAWID1,
  output [7:0] VCUPLENCAWLEN0,
  output [7:0] VCUPLENCAWLEN1,
  output VCUPLENCAWPROT0,
  output VCUPLENCAWPROT1,
  output [3:0] VCUPLENCAWQOS0,
  output [3:0] VCUPLENCAWQOS1,
  output [2:0] VCUPLENCAWSIZE0,
  output [2:0] VCUPLENCAWSIZE1,
  output VCUPLENCAWVALID0,
  output VCUPLENCAWVALID1,
  output VCUPLENCBREADY0,
  output VCUPLENCBREADY1,
  output VCUPLENCRREADY0,
  output VCUPLENCRREADY1,
  output [127:0] VCUPLENCWDATA0,
  output [127:0] VCUPLENCWDATA1,
  output VCUPLENCWLAST0,
  output VCUPLENCWLAST1,
  output VCUPLENCWVALID0,
  output VCUPLENCWVALID1,
  output [43:0] VCUPLMCUMAXIICDCARADDR,
  output [1:0] VCUPLMCUMAXIICDCARBURST,
  output [3:0] VCUPLMCUMAXIICDCARCACHE,
  output [2:0] VCUPLMCUMAXIICDCARID,
  output [7:0] VCUPLMCUMAXIICDCARLEN,
  output VCUPLMCUMAXIICDCARLOCK,
  output [2:0] VCUPLMCUMAXIICDCARPROT,
  output [3:0] VCUPLMCUMAXIICDCARQOS,
  output [2:0] VCUPLMCUMAXIICDCARSIZE,
  output VCUPLMCUMAXIICDCARVALID,
  output [43:0] VCUPLMCUMAXIICDCAWADDR,
  output [1:0] VCUPLMCUMAXIICDCAWBURST,
  output [3:0] VCUPLMCUMAXIICDCAWCACHE,
  output [2:0] VCUPLMCUMAXIICDCAWID,
  output [7:0] VCUPLMCUMAXIICDCAWLEN,
  output VCUPLMCUMAXIICDCAWLOCK,
  output [2:0] VCUPLMCUMAXIICDCAWPROT,
  output [3:0] VCUPLMCUMAXIICDCAWQOS,
  output [2:0] VCUPLMCUMAXIICDCAWSIZE,
  output VCUPLMCUMAXIICDCAWVALID,
  output VCUPLMCUMAXIICDCBREADY,
  output VCUPLMCUMAXIICDCRREADY,
  output [31:0] VCUPLMCUMAXIICDCWDATA,
  output VCUPLMCUMAXIICDCWLAST,
  output [3:0] VCUPLMCUMAXIICDCWSTRB,
  output VCUPLMCUMAXIICDCWVALID,
  output VCUPLMCUSTATUSCLKPLL,
  output VCUPLPINTREQ,
  output VCUPLPLLSTATUSPLLLOCK,
  output VCUPLPWRSUPPLYSTATUSVCCAUX,
  output VCUPLPWRSUPPLYSTATUSVCUINT,
  output [31:0] VCUPLRDATAAXILITEAPB,
  output [1:0] VCUPLRRESPAXILITEAPB,
  output VCUPLRVALIDAXILITEAPB,
  output VCUPLWREADYAXILITEAPB,
  input INITPLVCUGASKETCLAMPCONTROLLVLSHVCCINTD,
  input [19:0] PLVCUARADDRAXILITEAPB,
  input [2:0] PLVCUARPROTAXILITEAPB,
  input PLVCUARVALIDAXILITEAPB,
  input [19:0] PLVCUAWADDRAXILITEAPB,
  input [2:0] PLVCUAWPROTAXILITEAPB,
  input PLVCUAWVALIDAXILITEAPB,
  input PLVCUAXIDECCLK,
  input PLVCUAXIENCCLK,
  input PLVCUAXILITECLK,
  input PLVCUAXIMCUCLK,
  input PLVCUBREADYAXILITEAPB,
  input PLVCUCORECLK,
  input PLVCUDECARREADY0,
  input PLVCUDECARREADY1,
  input PLVCUDECAWREADY0,
  input PLVCUDECAWREADY1,
  input [3:0] PLVCUDECBID0,
  input [3:0] PLVCUDECBID1,
  input [1:0] PLVCUDECBRESP0,
  input [1:0] PLVCUDECBRESP1,
  input PLVCUDECBVALID0,
  input PLVCUDECBVALID1,
  input [127:0] PLVCUDECRDATA0,
  input [127:0] PLVCUDECRDATA1,
  input [3:0] PLVCUDECRID0,
  input [3:0] PLVCUDECRID1,
  input PLVCUDECRLAST0,
  input PLVCUDECRLAST1,
  input [1:0] PLVCUDECRRESP0,
  input [1:0] PLVCUDECRRESP1,
  input PLVCUDECRVALID0,
  input PLVCUDECRVALID1,
  input PLVCUDECWREADY0,
  input PLVCUDECWREADY1,
  input [319:0] PLVCUENCALL2CRDATA,
  input PLVCUENCALL2CRREADY,
  input PLVCUENCARREADY0,
  input PLVCUENCARREADY1,
  input PLVCUENCAWREADY0,
  input PLVCUENCAWREADY1,
  input [3:0] PLVCUENCBID0,
  input [3:0] PLVCUENCBID1,
  input [1:0] PLVCUENCBRESP0,
  input [1:0] PLVCUENCBRESP1,
  input PLVCUENCBVALID0,
  input PLVCUENCBVALID1,
  input PLVCUENCL2CCLK,
  input [127:0] PLVCUENCRDATA0,
  input [127:0] PLVCUENCRDATA1,
  input [3:0] PLVCUENCRID0,
  input [3:0] PLVCUENCRID1,
  input PLVCUENCRLAST0,
  input PLVCUENCRLAST1,
  input [1:0] PLVCUENCRRESP0,
  input [1:0] PLVCUENCRRESP1,
  input PLVCUENCRVALID0,
  input PLVCUENCRVALID1,
  input PLVCUENCWREADY0,
  input PLVCUENCWREADY1,
  input PLVCUMCUCLK,
  input PLVCUMCUMAXIICDCARREADY,
  input PLVCUMCUMAXIICDCAWREADY,
  input [2:0] PLVCUMCUMAXIICDCBID,
  input [1:0] PLVCUMCUMAXIICDCBRESP,
  input PLVCUMCUMAXIICDCBVALID,
  input [31:0] PLVCUMCUMAXIICDCRDATA,
  input [2:0] PLVCUMCUMAXIICDCRID,
  input PLVCUMCUMAXIICDCRLAST,
  input [1:0] PLVCUMCUMAXIICDCRRESP,
  input PLVCUMCUMAXIICDCRVALID,
  input PLVCUMCUMAXIICDCWREADY,
  input PLVCUPLLREFCLKPL,
  input PLVCURAWRSTN,
  input PLVCURREADYAXILITEAPB,
  input [31:0] PLVCUWDATAAXILITEAPB,
  input [3:0] PLVCUWSTRBAXILITEAPB,
  input PLVCUWVALIDAXILITEAPB
);
// define constants
  localparam MODULE_NAME = "VCU";
// Parameter encodings and registers
  localparam DECODERCHROMAFORMAT_4_2_0 = 1;
  localparam DECODERCHROMAFORMAT_4_2_2 = 0;
  localparam DECODERCODING_H_264 = 1;
  localparam DECODERCODING_H_265 = 0;
  localparam ENABLEDECODER_FALSE = 1;
  localparam ENABLEDECODER_TRUE = 0;
  localparam ENABLEENCODER_FALSE = 1;
  localparam ENABLEENCODER_TRUE = 0;
  localparam ENCODERCHROMAFORMAT_4_2_0 = 1;
  localparam ENCODERCHROMAFORMAT_4_2_2 = 0;
  localparam ENCODERCODING_H_264 = 1;
  localparam ENCODERCODING_H_265 = 0;
  reg trig_attr = 1'b0;
// include dynamic registers - XILINX test only
`ifdef XIL_DR
  `include "VCU_dr.v"
`else
  reg [31:0] CORECLKREQ_REG = CORECLKREQ;
  reg [31:0] DECHORRESOLUTION_REG = DECHORRESOLUTION;
  reg [40:1] DECODERCHROMAFORMAT_REG = DECODERCHROMAFORMAT;
  reg [40:1] DECODERCODING_REG = DECODERCODING;
  reg [31:0] DECODERCOLORDEPTH_REG = DECODERCOLORDEPTH;
  reg [31:0] DECODERNUMCORES_REG = DECODERNUMCORES;
  reg [31:0] DECVERTRESOLUTION_REG = DECVERTRESOLUTION;
  reg [40:1] ENABLEDECODER_REG = ENABLEDECODER;
  reg [40:1] ENABLEENCODER_REG = ENABLEENCODER;
  reg [31:0] ENCHORRESOLUTION_REG = ENCHORRESOLUTION;
  reg [40:1] ENCODERCHROMAFORMAT_REG = ENCODERCHROMAFORMAT;
  reg [40:1] ENCODERCODING_REG = ENCODERCODING;
  reg [31:0] ENCODERCOLORDEPTH_REG = ENCODERCOLORDEPTH;
  reg [31:0] ENCODERNUMCORES_REG = ENCODERNUMCORES;
  reg [31:0] ENCVERTRESOLUTION_REG = ENCVERTRESOLUTION;
`endif
`ifdef XIL_XECLIB
  wire [9:0] CORECLKREQ_BIN;
  wire [13:0] DECHORRESOLUTION_BIN;
  wire DECODERCHROMAFORMAT_BIN;
  wire DECODERCODING_BIN;
  wire [3:0] DECODERCOLORDEPTH_BIN;
  wire [1:0] DECODERNUMCORES_BIN;
  wire [12:0] DECVERTRESOLUTION_BIN;
  wire ENABLEDECODER_BIN;
  wire ENABLEENCODER_BIN;
  wire [13:0] ENCHORRESOLUTION_BIN;
  wire ENCODERCHROMAFORMAT_BIN;
  wire ENCODERCODING_BIN;
  wire [3:0] ENCODERCOLORDEPTH_BIN;
  wire [2:0] ENCODERNUMCORES_BIN;
  wire [12:0] ENCVERTRESOLUTION_BIN;
`else
  reg [9:0] CORECLKREQ_BIN;
  reg [13:0] DECHORRESOLUTION_BIN;
  reg DECODERCHROMAFORMAT_BIN;
  reg DECODERCODING_BIN;
  reg [3:0] DECODERCOLORDEPTH_BIN;
  reg [1:0] DECODERNUMCORES_BIN;
  reg [12:0] DECVERTRESOLUTION_BIN;
  reg ENABLEDECODER_BIN;
  reg ENABLEENCODER_BIN;
  reg [13:0] ENCHORRESOLUTION_BIN;
  reg ENCODERCHROMAFORMAT_BIN;
  reg ENCODERCODING_BIN;
  reg [3:0] ENCODERCOLORDEPTH_BIN;
  reg [2:0] ENCODERNUMCORES_BIN;
  reg [12:0] ENCVERTRESOLUTION_BIN;
`endif
`ifdef XIL_ATTR_TEST
  reg attr_test = 1'b1;
`else
  reg attr_test = 1'b0;
`endif
  reg attr_err = 1'b0;
  tri0 glblGSR = glbl.GSR;
//  reg VCUPLCORESTATUSCLKPLL_out;
//  reg VCUPLMCUSTATUSCLKPLL_out;
  reg VCUPLARREADYAXILITEAPB_out;
  reg VCUPLAWREADYAXILITEAPB_out;
  reg [1:0] VCUPLBRESPAXILITEAPB_out;
  reg VCUPLBVALIDAXILITEAPB_out;
  reg VCUPLCORESTATUSCLKPLL_out;
  reg [43:0] VCUPLDECARADDR0_out;
  reg [43:0] VCUPLDECARADDR1_out;
  reg [1:0] VCUPLDECARBURST0_out;
  reg [1:0] VCUPLDECARBURST1_out;
  reg [3:0] VCUPLDECARCACHE0_out;
  reg [3:0] VCUPLDECARCACHE1_out;
  reg [3:0] VCUPLDECARID0_out;
  reg [3:0] VCUPLDECARID1_out;
  reg [7:0] VCUPLDECARLEN0_out;
  reg [7:0] VCUPLDECARLEN1_out;
  reg VCUPLDECARPROT0_out;
  reg VCUPLDECARPROT1_out;
  reg [3:0] VCUPLDECARQOS0_out;
  reg [3:0] VCUPLDECARQOS1_out;
  reg [2:0] VCUPLDECARSIZE0_out;
  reg [2:0] VCUPLDECARSIZE1_out;
  reg VCUPLDECARVALID0_out;
  reg VCUPLDECARVALID1_out;
  reg [43:0] VCUPLDECAWADDR0_out;
  reg [43:0] VCUPLDECAWADDR1_out;
  reg [1:0] VCUPLDECAWBURST0_out;
  reg [1:0] VCUPLDECAWBURST1_out;
  reg [3:0] VCUPLDECAWCACHE0_out;
  reg [3:0] VCUPLDECAWCACHE1_out;
  reg [3:0] VCUPLDECAWID0_out;
  reg [3:0] VCUPLDECAWID1_out;
  reg [7:0] VCUPLDECAWLEN0_out;
  reg [7:0] VCUPLDECAWLEN1_out;
  reg VCUPLDECAWPROT0_out;
  reg VCUPLDECAWPROT1_out;
  reg [3:0] VCUPLDECAWQOS0_out;
  reg [3:0] VCUPLDECAWQOS1_out;
  reg [2:0] VCUPLDECAWSIZE0_out;
  reg [2:0] VCUPLDECAWSIZE1_out;
  reg VCUPLDECAWVALID0_out;
  reg VCUPLDECAWVALID1_out;
  reg VCUPLDECBREADY0_out;
  reg VCUPLDECBREADY1_out;
  reg VCUPLDECRREADY0_out;
  reg VCUPLDECRREADY1_out;
  reg [127:0] VCUPLDECWDATA0_out;
  reg [127:0] VCUPLDECWDATA1_out;
  reg VCUPLDECWLAST0_out;
  reg VCUPLDECWLAST1_out;
  reg VCUPLDECWVALID0_out;
  reg VCUPLDECWVALID1_out;
  reg [16:0] VCUPLENCALL2CADDR_out;
  reg VCUPLENCALL2CRVALID_out;
  reg [319:0] VCUPLENCALL2CWDATA_out;
  reg VCUPLENCALL2CWVALID_out;
  reg [43:0] VCUPLENCARADDR0_out;
  reg [43:0] VCUPLENCARADDR1_out;
  reg [1:0] VCUPLENCARBURST0_out;
  reg [1:0] VCUPLENCARBURST1_out;
  reg [3:0] VCUPLENCARCACHE0_out;
  reg [3:0] VCUPLENCARCACHE1_out;
  reg [3:0] VCUPLENCARID0_out;
  reg [3:0] VCUPLENCARID1_out;
  reg [7:0] VCUPLENCARLEN0_out;
  reg [7:0] VCUPLENCARLEN1_out;
  reg VCUPLENCARPROT0_out;
  reg VCUPLENCARPROT1_out;
  reg [3:0] VCUPLENCARQOS0_out;
  reg [3:0] VCUPLENCARQOS1_out;
  reg [2:0] VCUPLENCARSIZE0_out;
  reg [2:0] VCUPLENCARSIZE1_out;
  reg VCUPLENCARVALID0_out;
  reg VCUPLENCARVALID1_out;
  reg [43:0] VCUPLENCAWADDR0_out;
  reg [43:0] VCUPLENCAWADDR1_out;
  reg [1:0] VCUPLENCAWBURST0_out;
  reg [1:0] VCUPLENCAWBURST1_out;
  reg [3:0] VCUPLENCAWCACHE0_out;
  reg [3:0] VCUPLENCAWCACHE1_out;
  reg [3:0] VCUPLENCAWID0_out;
  reg [3:0] VCUPLENCAWID1_out;
  reg [7:0] VCUPLENCAWLEN0_out;
  reg [7:0] VCUPLENCAWLEN1_out;
  reg VCUPLENCAWPROT0_out;
  reg VCUPLENCAWPROT1_out;
  reg [3:0] VCUPLENCAWQOS0_out;
  reg [3:0] VCUPLENCAWQOS1_out;
  reg [2:0] VCUPLENCAWSIZE0_out;
  reg [2:0] VCUPLENCAWSIZE1_out;
  reg VCUPLENCAWVALID0_out;
  reg VCUPLENCAWVALID1_out;
  reg VCUPLENCBREADY0_out;
  reg VCUPLENCBREADY1_out;
  reg VCUPLENCRREADY0_out;
  reg VCUPLENCRREADY1_out;
  reg [127:0] VCUPLENCWDATA0_out;
  reg [127:0] VCUPLENCWDATA1_out;
  reg VCUPLENCWLAST0_out;
  reg VCUPLENCWLAST1_out;
  reg VCUPLENCWVALID0_out;
  reg VCUPLENCWVALID1_out;
  reg [43:0] VCUPLMCUMAXIICDCARADDR_out;
  reg [1:0] VCUPLMCUMAXIICDCARBURST_out;
  reg [3:0] VCUPLMCUMAXIICDCARCACHE_out;
  reg [2:0] VCUPLMCUMAXIICDCARID_out;
  reg [7:0] VCUPLMCUMAXIICDCARLEN_out;
  reg VCUPLMCUMAXIICDCARLOCK_out;
  reg [2:0] VCUPLMCUMAXIICDCARPROT_out;
  reg [3:0] VCUPLMCUMAXIICDCARQOS_out;
  reg [2:0] VCUPLMCUMAXIICDCARSIZE_out;
  reg VCUPLMCUMAXIICDCARVALID_out;
  reg [43:0] VCUPLMCUMAXIICDCAWADDR_out;
  reg [1:0] VCUPLMCUMAXIICDCAWBURST_out;
  reg [3:0] VCUPLMCUMAXIICDCAWCACHE_out;
  reg [2:0] VCUPLMCUMAXIICDCAWID_out;
  reg [7:0] VCUPLMCUMAXIICDCAWLEN_out;
  reg VCUPLMCUMAXIICDCAWLOCK_out;
  reg [2:0] VCUPLMCUMAXIICDCAWPROT_out;
  reg [3:0] VCUPLMCUMAXIICDCAWQOS_out;
  reg [2:0] VCUPLMCUMAXIICDCAWSIZE_out;
  reg VCUPLMCUMAXIICDCAWVALID_out;
  reg VCUPLMCUMAXIICDCBREADY_out;
  reg VCUPLMCUMAXIICDCRREADY_out;
  reg [31:0] VCUPLMCUMAXIICDCWDATA_out;
  reg VCUPLMCUMAXIICDCWLAST_out;
  reg [3:0] VCUPLMCUMAXIICDCWSTRB_out;
  reg VCUPLMCUMAXIICDCWVALID_out;
  reg VCUPLMCUSTATUSCLKPLL_out;
  reg VCUPLPINTREQ_out;
  reg VCUPLPLLSTATUSPLLLOCK_out;
  reg VCUPLPWRSUPPLYSTATUSVCCAUX_out;
  reg VCUPLPWRSUPPLYSTATUSVCUINT_out;
  reg [31:0] VCUPLRDATAAXILITEAPB_out;
  reg [1:0] VCUPLRRESPAXILITEAPB_out;
  reg VCUPLRVALIDAXILITEAPB_out;
  reg VCUPLWREADYAXILITEAPB_out;
  wire INITPLVCUGASKETCLAMPCONTROLLVLSHVCCINTD_in;
  wire PLVCUARVALIDAXILITEAPB_in;
  wire PLVCUAWVALIDAXILITEAPB_in;
  wire PLVCUAXIDECCLK_in;
  wire PLVCUAXIENCCLK_in;
  wire PLVCUAXILITECLK_in;
  wire PLVCUAXIMCUCLK_in;
  wire PLVCUBREADYAXILITEAPB_in;
  wire PLVCUCORECLK_in;
  wire PLVCUDECARREADY0_in;
  wire PLVCUDECARREADY1_in;
  wire PLVCUDECAWREADY0_in;
  wire PLVCUDECAWREADY1_in;
  wire PLVCUDECBVALID0_in;
  wire PLVCUDECBVALID1_in;
  wire PLVCUDECRLAST0_in;
  wire PLVCUDECRLAST1_in;
  wire PLVCUDECRVALID0_in;
  wire PLVCUDECRVALID1_in;
  wire PLVCUDECWREADY0_in;
  wire PLVCUDECWREADY1_in;
  wire PLVCUENCALL2CRREADY_in;
  wire PLVCUENCARREADY0_in;
  wire PLVCUENCARREADY1_in;
  wire PLVCUENCAWREADY0_in;
  wire PLVCUENCAWREADY1_in;
  wire PLVCUENCBVALID0_in;
  wire PLVCUENCBVALID1_in;
  wire PLVCUENCL2CCLK_in;
  wire PLVCUENCRLAST0_in;
  wire PLVCUENCRLAST1_in;
  wire PLVCUENCRVALID0_in;
  wire PLVCUENCRVALID1_in;
  wire PLVCUENCWREADY0_in;
  wire PLVCUENCWREADY1_in;
  wire PLVCUMCUCLK_in;
  wire PLVCUMCUMAXIICDCARREADY_in;
  wire PLVCUMCUMAXIICDCAWREADY_in;
  wire PLVCUMCUMAXIICDCBVALID_in;
  wire PLVCUMCUMAXIICDCRLAST_in;
  wire PLVCUMCUMAXIICDCRVALID_in;
  wire PLVCUMCUMAXIICDCWREADY_in;
  wire PLVCUPLLREFCLKPL_in;
  wire PLVCURAWRSTN_in;
  wire PLVCURREADYAXILITEAPB_in;
  wire PLVCUWVALIDAXILITEAPB_in;
  wire [127:0] PLVCUDECRDATA0_in;
  wire [127:0] PLVCUDECRDATA1_in;
  wire [127:0] PLVCUENCRDATA0_in;
  wire [127:0] PLVCUENCRDATA1_in;
  wire [19:0] PLVCUARADDRAXILITEAPB_in;
  wire [19:0] PLVCUAWADDRAXILITEAPB_in;
  wire [1:0] PLVCUDECBRESP0_in;
  wire [1:0] PLVCUDECBRESP1_in;
  wire [1:0] PLVCUDECRRESP0_in;
  wire [1:0] PLVCUDECRRESP1_in;
  wire [1:0] PLVCUENCBRESP0_in;
  wire [1:0] PLVCUENCBRESP1_in;
  wire [1:0] PLVCUENCRRESP0_in;
  wire [1:0] PLVCUENCRRESP1_in;
  wire [1:0] PLVCUMCUMAXIICDCBRESP_in;
  wire [1:0] PLVCUMCUMAXIICDCRRESP_in;
  wire [2:0] PLVCUARPROTAXILITEAPB_in;
  wire [2:0] PLVCUAWPROTAXILITEAPB_in;
  wire [2:0] PLVCUMCUMAXIICDCBID_in;
  wire [2:0] PLVCUMCUMAXIICDCRID_in;
  wire [319:0] PLVCUENCALL2CRDATA_in;
  wire [31:0] PLVCUMCUMAXIICDCRDATA_in;
  wire [31:0] PLVCUWDATAAXILITEAPB_in;
  wire [3:0] PLVCUDECBID0_in;
  wire [3:0] PLVCUDECBID1_in;
  wire [3:0] PLVCUDECRID0_in;
  wire [3:0] PLVCUDECRID1_in;
  wire [3:0] PLVCUENCBID0_in;
  wire [3:0] PLVCUENCBID1_in;
  wire [3:0] PLVCUENCRID0_in;
  wire [3:0] PLVCUENCRID1_in;
  wire [3:0] PLVCUWSTRBAXILITEAPB_in;
`ifdef XIL_TIMING
  wire PLVCUARVALIDAXILITEAPB_delay;
  wire PLVCUAWVALIDAXILITEAPB_delay;
  wire PLVCUAXIDECCLK_delay;
  wire PLVCUAXIENCCLK_delay;
  wire PLVCUAXILITECLK_delay;
  wire PLVCUAXIMCUCLK_delay;
  wire PLVCUBREADYAXILITEAPB_delay;
  wire PLVCUDECARREADY0_delay;
  wire PLVCUDECARREADY1_delay;
  wire PLVCUDECAWREADY0_delay;
  wire PLVCUDECAWREADY1_delay;
  wire PLVCUDECBVALID0_delay;
  wire PLVCUDECBVALID1_delay;
  wire PLVCUDECRLAST0_delay;
  wire PLVCUDECRLAST1_delay;
  wire PLVCUDECRVALID0_delay;
  wire PLVCUDECRVALID1_delay;
  wire PLVCUDECWREADY0_delay;
  wire PLVCUDECWREADY1_delay;
  wire PLVCUENCALL2CRREADY_delay;
  wire PLVCUENCARREADY0_delay;
  wire PLVCUENCARREADY1_delay;
  wire PLVCUENCAWREADY0_delay;
  wire PLVCUENCAWREADY1_delay;
  wire PLVCUENCBVALID0_delay;
  wire PLVCUENCBVALID1_delay;
  wire PLVCUENCL2CCLK_delay;
  wire PLVCUENCRLAST0_delay;
  wire PLVCUENCRLAST1_delay;
  wire PLVCUENCRVALID0_delay;
  wire PLVCUENCRVALID1_delay;
  wire PLVCUENCWREADY0_delay;
  wire PLVCUENCWREADY1_delay;
  wire PLVCUMCUMAXIICDCARREADY_delay;
  wire PLVCUMCUMAXIICDCAWREADY_delay;
  wire PLVCUMCUMAXIICDCBVALID_delay;
  wire PLVCUMCUMAXIICDCRLAST_delay;
  wire PLVCUMCUMAXIICDCRVALID_delay;
  wire PLVCUMCUMAXIICDCWREADY_delay;
  wire PLVCURREADYAXILITEAPB_delay;
  wire PLVCUWVALIDAXILITEAPB_delay;
  wire [127:0] PLVCUDECRDATA0_delay;
  wire [127:0] PLVCUDECRDATA1_delay;
  wire [127:0] PLVCUENCRDATA0_delay;
  wire [127:0] PLVCUENCRDATA1_delay;
  wire [19:0] PLVCUARADDRAXILITEAPB_delay;
  wire [19:0] PLVCUAWADDRAXILITEAPB_delay;
  wire [1:0] PLVCUDECBRESP0_delay;
  wire [1:0] PLVCUDECBRESP1_delay;
  wire [1:0] PLVCUDECRRESP0_delay;
  wire [1:0] PLVCUDECRRESP1_delay;
  wire [1:0] PLVCUENCBRESP0_delay;
  wire [1:0] PLVCUENCBRESP1_delay;
  wire [1:0] PLVCUENCRRESP0_delay;
  wire [1:0] PLVCUENCRRESP1_delay;
  wire [1:0] PLVCUMCUMAXIICDCBRESP_delay;
  wire [1:0] PLVCUMCUMAXIICDCRRESP_delay;
  wire [2:0] PLVCUARPROTAXILITEAPB_delay;
  wire [2:0] PLVCUAWPROTAXILITEAPB_delay;
  wire [2:0] PLVCUMCUMAXIICDCBID_delay;
  wire [2:0] PLVCUMCUMAXIICDCRID_delay;
  wire [319:0] PLVCUENCALL2CRDATA_delay;
  wire [31:0] PLVCUMCUMAXIICDCRDATA_delay;
  wire [31:0] PLVCUWDATAAXILITEAPB_delay;
  wire [3:0] PLVCUDECBID0_delay;
  wire [3:0] PLVCUDECBID1_delay;
  wire [3:0] PLVCUDECRID0_delay;
  wire [3:0] PLVCUDECRID1_delay;
  wire [3:0] PLVCUENCBID0_delay;
  wire [3:0] PLVCUENCBID1_delay;
  wire [3:0] PLVCUENCRID0_delay;
  wire [3:0] PLVCUENCRID1_delay;
  wire [3:0] PLVCUWSTRBAXILITEAPB_delay;
`endif
//  assign VCUPLCORESTATUSCLKPLL = VCUPLCORESTATUSCLKPLL_out;
//  assign VCUPLMCUSTATUSCLKPLL = VCUPLMCUSTATUSCLKPLL_out;
  assign VCUPLARREADYAXILITEAPB = VCUPLARREADYAXILITEAPB_out;
  assign VCUPLAWREADYAXILITEAPB = VCUPLAWREADYAXILITEAPB_out;
  assign VCUPLBRESPAXILITEAPB = VCUPLBRESPAXILITEAPB_out;
  assign VCUPLBVALIDAXILITEAPB = VCUPLBVALIDAXILITEAPB_out;
  assign VCUPLCORESTATUSCLKPLL = VCUPLCORESTATUSCLKPLL_out;
  assign VCUPLDECARADDR0 = VCUPLDECARADDR0_out;
  assign VCUPLDECARADDR1 = VCUPLDECARADDR1_out;
  assign VCUPLDECARBURST0 = VCUPLDECARBURST0_out;
  assign VCUPLDECARBURST1 = VCUPLDECARBURST1_out;
  assign VCUPLDECARCACHE0 = VCUPLDECARCACHE0_out;
  assign VCUPLDECARCACHE1 = VCUPLDECARCACHE1_out;
  assign VCUPLDECARID0 = VCUPLDECARID0_out;
  assign VCUPLDECARID1 = VCUPLDECARID1_out;
  assign VCUPLDECARLEN0 = VCUPLDECARLEN0_out;
  assign VCUPLDECARLEN1 = VCUPLDECARLEN1_out;
  assign VCUPLDECARPROT0 = VCUPLDECARPROT0_out;
  assign VCUPLDECARPROT1 = VCUPLDECARPROT1_out;
  assign VCUPLDECARQOS0 = VCUPLDECARQOS0_out;
  assign VCUPLDECARQOS1 = VCUPLDECARQOS1_out;
  assign VCUPLDECARSIZE0 = VCUPLDECARSIZE0_out;
  assign VCUPLDECARSIZE1 = VCUPLDECARSIZE1_out;
  assign VCUPLDECARVALID0 = VCUPLDECARVALID0_out;
  assign VCUPLDECARVALID1 = VCUPLDECARVALID1_out;
  assign VCUPLDECAWADDR0 = VCUPLDECAWADDR0_out;
  assign VCUPLDECAWADDR1 = VCUPLDECAWADDR1_out;
  assign VCUPLDECAWBURST0 = VCUPLDECAWBURST0_out;
  assign VCUPLDECAWBURST1 = VCUPLDECAWBURST1_out;
  assign VCUPLDECAWCACHE0 = VCUPLDECAWCACHE0_out;
  assign VCUPLDECAWCACHE1 = VCUPLDECAWCACHE1_out;
  assign VCUPLDECAWID0 = VCUPLDECAWID0_out;
  assign VCUPLDECAWID1 = VCUPLDECAWID1_out;
  assign VCUPLDECAWLEN0 = VCUPLDECAWLEN0_out;
  assign VCUPLDECAWLEN1 = VCUPLDECAWLEN1_out;
  assign VCUPLDECAWPROT0 = VCUPLDECAWPROT0_out;
  assign VCUPLDECAWPROT1 = VCUPLDECAWPROT1_out;
  assign VCUPLDECAWQOS0 = VCUPLDECAWQOS0_out;
  assign VCUPLDECAWQOS1 = VCUPLDECAWQOS1_out;
  assign VCUPLDECAWSIZE0 = VCUPLDECAWSIZE0_out;
  assign VCUPLDECAWSIZE1 = VCUPLDECAWSIZE1_out;
  assign VCUPLDECAWVALID0 = VCUPLDECAWVALID0_out;
  assign VCUPLDECAWVALID1 = VCUPLDECAWVALID1_out;
  assign VCUPLDECBREADY0 = VCUPLDECBREADY0_out;
  assign VCUPLDECBREADY1 = VCUPLDECBREADY1_out;
  assign VCUPLDECRREADY0 = VCUPLDECRREADY0_out;
  assign VCUPLDECRREADY1 = VCUPLDECRREADY1_out;
  assign VCUPLDECWDATA0 = VCUPLDECWDATA0_out;
  assign VCUPLDECWDATA1 = VCUPLDECWDATA1_out;
  assign VCUPLDECWLAST0 = VCUPLDECWLAST0_out;
  assign VCUPLDECWLAST1 = VCUPLDECWLAST1_out;
  assign VCUPLDECWVALID0 = VCUPLDECWVALID0_out;
  assign VCUPLDECWVALID1 = VCUPLDECWVALID1_out;
  assign VCUPLENCALL2CADDR = VCUPLENCALL2CADDR_out;
  assign VCUPLENCALL2CRVALID = VCUPLENCALL2CRVALID_out;
  assign VCUPLENCALL2CWDATA = VCUPLENCALL2CWDATA_out;
  assign VCUPLENCALL2CWVALID = VCUPLENCALL2CWVALID_out;
  assign VCUPLENCARADDR0 = VCUPLENCARADDR0_out;
  assign VCUPLENCARADDR1 = VCUPLENCARADDR1_out;
  assign VCUPLENCARBURST0 = VCUPLENCARBURST0_out;
  assign VCUPLENCARBURST1 = VCUPLENCARBURST1_out;
  assign VCUPLENCARCACHE0 = VCUPLENCARCACHE0_out;
  assign VCUPLENCARCACHE1 = VCUPLENCARCACHE1_out;
  assign VCUPLENCARID0 = VCUPLENCARID0_out;
  assign VCUPLENCARID1 = VCUPLENCARID1_out;
  assign VCUPLENCARLEN0 = VCUPLENCARLEN0_out;
  assign VCUPLENCARLEN1 = VCUPLENCARLEN1_out;
  assign VCUPLENCARPROT0 = VCUPLENCARPROT0_out;
  assign VCUPLENCARPROT1 = VCUPLENCARPROT1_out;
  assign VCUPLENCARQOS0 = VCUPLENCARQOS0_out;
  assign VCUPLENCARQOS1 = VCUPLENCARQOS1_out;
  assign VCUPLENCARSIZE0 = VCUPLENCARSIZE0_out;
  assign VCUPLENCARSIZE1 = VCUPLENCARSIZE1_out;
  assign VCUPLENCARVALID0 = VCUPLENCARVALID0_out;
  assign VCUPLENCARVALID1 = VCUPLENCARVALID1_out;
  assign VCUPLENCAWADDR0 = VCUPLENCAWADDR0_out;
  assign VCUPLENCAWADDR1 = VCUPLENCAWADDR1_out;
  assign VCUPLENCAWBURST0 = VCUPLENCAWBURST0_out;
  assign VCUPLENCAWBURST1 = VCUPLENCAWBURST1_out;
  assign VCUPLENCAWCACHE0 = VCUPLENCAWCACHE0_out;
  assign VCUPLENCAWCACHE1 = VCUPLENCAWCACHE1_out;
  assign VCUPLENCAWID0 = VCUPLENCAWID0_out;
  assign VCUPLENCAWID1 = VCUPLENCAWID1_out;
  assign VCUPLENCAWLEN0 = VCUPLENCAWLEN0_out;
  assign VCUPLENCAWLEN1 = VCUPLENCAWLEN1_out;
  assign VCUPLENCAWPROT0 = VCUPLENCAWPROT0_out;
  assign VCUPLENCAWPROT1 = VCUPLENCAWPROT1_out;
  assign VCUPLENCAWQOS0 = VCUPLENCAWQOS0_out;
  assign VCUPLENCAWQOS1 = VCUPLENCAWQOS1_out;
  assign VCUPLENCAWSIZE0 = VCUPLENCAWSIZE0_out;
  assign VCUPLENCAWSIZE1 = VCUPLENCAWSIZE1_out;
  assign VCUPLENCAWVALID0 = VCUPLENCAWVALID0_out;
  assign VCUPLENCAWVALID1 = VCUPLENCAWVALID1_out;
  assign VCUPLENCBREADY0 = VCUPLENCBREADY0_out;
  assign VCUPLENCBREADY1 = VCUPLENCBREADY1_out;
  assign VCUPLENCRREADY0 = VCUPLENCRREADY0_out;
  assign VCUPLENCRREADY1 = VCUPLENCRREADY1_out;
  assign VCUPLENCWDATA0 = VCUPLENCWDATA0_out;
  assign VCUPLENCWDATA1 = VCUPLENCWDATA1_out;
  assign VCUPLENCWLAST0 = VCUPLENCWLAST0_out;
  assign VCUPLENCWLAST1 = VCUPLENCWLAST1_out;
  assign VCUPLENCWVALID0 = VCUPLENCWVALID0_out;
  assign VCUPLENCWVALID1 = VCUPLENCWVALID1_out;
  assign VCUPLMCUMAXIICDCARADDR = VCUPLMCUMAXIICDCARADDR_out;
  assign VCUPLMCUMAXIICDCARBURST = VCUPLMCUMAXIICDCARBURST_out;
  assign VCUPLMCUMAXIICDCARCACHE = VCUPLMCUMAXIICDCARCACHE_out;
  assign VCUPLMCUMAXIICDCARID = VCUPLMCUMAXIICDCARID_out;
  assign VCUPLMCUMAXIICDCARLEN = VCUPLMCUMAXIICDCARLEN_out;
  assign VCUPLMCUMAXIICDCARLOCK = VCUPLMCUMAXIICDCARLOCK_out;
  assign VCUPLMCUMAXIICDCARPROT = VCUPLMCUMAXIICDCARPROT_out;
  assign VCUPLMCUMAXIICDCARQOS = VCUPLMCUMAXIICDCARQOS_out;
  assign VCUPLMCUMAXIICDCARSIZE = VCUPLMCUMAXIICDCARSIZE_out;
  assign VCUPLMCUMAXIICDCARVALID = VCUPLMCUMAXIICDCARVALID_out;
  assign VCUPLMCUMAXIICDCAWADDR = VCUPLMCUMAXIICDCAWADDR_out;
  assign VCUPLMCUMAXIICDCAWBURST = VCUPLMCUMAXIICDCAWBURST_out;
  assign VCUPLMCUMAXIICDCAWCACHE = VCUPLMCUMAXIICDCAWCACHE_out;
  assign VCUPLMCUMAXIICDCAWID = VCUPLMCUMAXIICDCAWID_out;
  assign VCUPLMCUMAXIICDCAWLEN = VCUPLMCUMAXIICDCAWLEN_out;
  assign VCUPLMCUMAXIICDCAWLOCK = VCUPLMCUMAXIICDCAWLOCK_out;
  assign VCUPLMCUMAXIICDCAWPROT = VCUPLMCUMAXIICDCAWPROT_out;
  assign VCUPLMCUMAXIICDCAWQOS = VCUPLMCUMAXIICDCAWQOS_out;
  assign VCUPLMCUMAXIICDCAWSIZE = VCUPLMCUMAXIICDCAWSIZE_out;
  assign VCUPLMCUMAXIICDCAWVALID = VCUPLMCUMAXIICDCAWVALID_out;
  assign VCUPLMCUMAXIICDCBREADY = VCUPLMCUMAXIICDCBREADY_out;
  assign VCUPLMCUMAXIICDCRREADY = VCUPLMCUMAXIICDCRREADY_out;
  assign VCUPLMCUMAXIICDCWDATA = VCUPLMCUMAXIICDCWDATA_out;
  assign VCUPLMCUMAXIICDCWLAST = VCUPLMCUMAXIICDCWLAST_out;
  assign VCUPLMCUMAXIICDCWSTRB = VCUPLMCUMAXIICDCWSTRB_out;
  assign VCUPLMCUMAXIICDCWVALID = VCUPLMCUMAXIICDCWVALID_out;
  assign VCUPLMCUSTATUSCLKPLL = VCUPLMCUSTATUSCLKPLL_out;
  assign VCUPLPINTREQ = VCUPLPINTREQ_out;
  assign VCUPLPLLSTATUSPLLLOCK = VCUPLPLLSTATUSPLLLOCK_out;
  assign VCUPLPWRSUPPLYSTATUSVCCAUX = VCUPLPWRSUPPLYSTATUSVCCAUX_out;
  assign VCUPLPWRSUPPLYSTATUSVCUINT = VCUPLPWRSUPPLYSTATUSVCUINT_out;
  assign VCUPLRDATAAXILITEAPB = VCUPLRDATAAXILITEAPB_out;
  assign VCUPLRRESPAXILITEAPB = VCUPLRRESPAXILITEAPB_out;
  assign VCUPLRVALIDAXILITEAPB = VCUPLRVALIDAXILITEAPB_out;
  assign VCUPLWREADYAXILITEAPB = VCUPLWREADYAXILITEAPB_out;
`ifdef XIL_TIMING
  assign PLVCUARADDRAXILITEAPB_in = PLVCUARADDRAXILITEAPB_delay;
  assign PLVCUARPROTAXILITEAPB_in = PLVCUARPROTAXILITEAPB_delay;
  assign PLVCUARVALIDAXILITEAPB_in = PLVCUARVALIDAXILITEAPB_delay;
  assign PLVCUAWADDRAXILITEAPB_in = PLVCUAWADDRAXILITEAPB_delay;
  assign PLVCUAWPROTAXILITEAPB_in = PLVCUAWPROTAXILITEAPB_delay;
  assign PLVCUAWVALIDAXILITEAPB_in = PLVCUAWVALIDAXILITEAPB_delay;
  assign PLVCUAXIDECCLK_in = PLVCUAXIDECCLK_delay;
  assign PLVCUAXIENCCLK_in = PLVCUAXIENCCLK_delay;
  assign PLVCUAXILITECLK_in = PLVCUAXILITECLK_delay;
  assign PLVCUAXIMCUCLK_in = PLVCUAXIMCUCLK_delay;
  assign PLVCUBREADYAXILITEAPB_in = PLVCUBREADYAXILITEAPB_delay;
  assign PLVCUDECARREADY0_in = PLVCUDECARREADY0_delay;
  assign PLVCUDECARREADY1_in = PLVCUDECARREADY1_delay;
  assign PLVCUDECAWREADY0_in = PLVCUDECAWREADY0_delay;
  assign PLVCUDECAWREADY1_in = PLVCUDECAWREADY1_delay;
  assign PLVCUDECBID0_in = PLVCUDECBID0_delay;
  assign PLVCUDECBID1_in = PLVCUDECBID1_delay;
  assign PLVCUDECBRESP0_in = PLVCUDECBRESP0_delay;
  assign PLVCUDECBRESP1_in = PLVCUDECBRESP1_delay;
  assign PLVCUDECBVALID0_in = PLVCUDECBVALID0_delay;
  assign PLVCUDECBVALID1_in = PLVCUDECBVALID1_delay;
  assign PLVCUDECRDATA0_in = PLVCUDECRDATA0_delay;
  assign PLVCUDECRDATA1_in = PLVCUDECRDATA1_delay;
  assign PLVCUDECRID0_in = PLVCUDECRID0_delay;
  assign PLVCUDECRID1_in = PLVCUDECRID1_delay;
  assign PLVCUDECRLAST0_in = PLVCUDECRLAST0_delay;
  assign PLVCUDECRLAST1_in = PLVCUDECRLAST1_delay;
  assign PLVCUDECRRESP0_in = PLVCUDECRRESP0_delay;
  assign PLVCUDECRRESP1_in = PLVCUDECRRESP1_delay;
  assign PLVCUDECRVALID0_in = PLVCUDECRVALID0_delay;
  assign PLVCUDECRVALID1_in = PLVCUDECRVALID1_delay;
  assign PLVCUDECWREADY0_in = PLVCUDECWREADY0_delay;
  assign PLVCUDECWREADY1_in = PLVCUDECWREADY1_delay;
  assign PLVCUENCALL2CRDATA_in = PLVCUENCALL2CRDATA_delay;
  assign PLVCUENCALL2CRREADY_in = (PLVCUENCALL2CRREADY === 1'bz) || PLVCUENCALL2CRREADY_delay; // rv 1
  assign PLVCUENCARREADY0_in = PLVCUENCARREADY0_delay;
  assign PLVCUENCARREADY1_in = PLVCUENCARREADY1_delay;
  assign PLVCUENCAWREADY0_in = PLVCUENCAWREADY0_delay;
  assign PLVCUENCAWREADY1_in = PLVCUENCAWREADY1_delay;
  assign PLVCUENCBID0_in = PLVCUENCBID0_delay;
  assign PLVCUENCBID1_in = PLVCUENCBID1_delay;
  assign PLVCUENCBRESP0_in = PLVCUENCBRESP0_delay;
  assign PLVCUENCBRESP1_in = PLVCUENCBRESP1_delay;
  assign PLVCUENCBVALID0_in = PLVCUENCBVALID0_delay;
  assign PLVCUENCBVALID1_in = PLVCUENCBVALID1_delay;
  assign PLVCUENCL2CCLK_in = PLVCUENCL2CCLK_delay;
  assign PLVCUENCRDATA0_in = PLVCUENCRDATA0_delay;
  assign PLVCUENCRDATA1_in = PLVCUENCRDATA1_delay;
  assign PLVCUENCRID0_in = PLVCUENCRID0_delay;
  assign PLVCUENCRID1_in = PLVCUENCRID1_delay;
  assign PLVCUENCRLAST0_in = PLVCUENCRLAST0_delay;
  assign PLVCUENCRLAST1_in = PLVCUENCRLAST1_delay;
  assign PLVCUENCRRESP0_in = PLVCUENCRRESP0_delay;
  assign PLVCUENCRRESP1_in = PLVCUENCRRESP1_delay;
  assign PLVCUENCRVALID0_in = PLVCUENCRVALID0_delay;
  assign PLVCUENCRVALID1_in = PLVCUENCRVALID1_delay;
  assign PLVCUENCWREADY0_in = PLVCUENCWREADY0_delay;
  assign PLVCUENCWREADY1_in = PLVCUENCWREADY1_delay;
  assign PLVCUMCUMAXIICDCARREADY_in = PLVCUMCUMAXIICDCARREADY_delay;
  assign PLVCUMCUMAXIICDCAWREADY_in = PLVCUMCUMAXIICDCAWREADY_delay;
  assign PLVCUMCUMAXIICDCBID_in = PLVCUMCUMAXIICDCBID_delay;
  assign PLVCUMCUMAXIICDCBRESP_in = PLVCUMCUMAXIICDCBRESP_delay;
  assign PLVCUMCUMAXIICDCBVALID_in = PLVCUMCUMAXIICDCBVALID_delay;
  assign PLVCUMCUMAXIICDCRDATA_in = PLVCUMCUMAXIICDCRDATA_delay;
  assign PLVCUMCUMAXIICDCRID_in = PLVCUMCUMAXIICDCRID_delay;
  assign PLVCUMCUMAXIICDCRLAST_in = PLVCUMCUMAXIICDCRLAST_delay;
  assign PLVCUMCUMAXIICDCRRESP_in = PLVCUMCUMAXIICDCRRESP_delay;
  assign PLVCUMCUMAXIICDCRVALID_in = PLVCUMCUMAXIICDCRVALID_delay;
  assign PLVCUMCUMAXIICDCWREADY_in = PLVCUMCUMAXIICDCWREADY_delay;
  assign PLVCURREADYAXILITEAPB_in = PLVCURREADYAXILITEAPB_delay;
  assign PLVCUWDATAAXILITEAPB_in = PLVCUWDATAAXILITEAPB_delay;
  assign PLVCUWSTRBAXILITEAPB_in = PLVCUWSTRBAXILITEAPB_delay;
  assign PLVCUWVALIDAXILITEAPB_in = PLVCUWVALIDAXILITEAPB_delay;
`else
  assign PLVCUARADDRAXILITEAPB_in = PLVCUARADDRAXILITEAPB;
  assign PLVCUARPROTAXILITEAPB_in = PLVCUARPROTAXILITEAPB;
  assign PLVCUARVALIDAXILITEAPB_in = PLVCUARVALIDAXILITEAPB;
  assign PLVCUAWADDRAXILITEAPB_in = PLVCUAWADDRAXILITEAPB;
  assign PLVCUAWPROTAXILITEAPB_in = PLVCUAWPROTAXILITEAPB;
  assign PLVCUAWVALIDAXILITEAPB_in = PLVCUAWVALIDAXILITEAPB;
  assign PLVCUAXIDECCLK_in = PLVCUAXIDECCLK;
  assign PLVCUAXIENCCLK_in = PLVCUAXIENCCLK;
  assign PLVCUAXILITECLK_in = PLVCUAXILITECLK;
  assign PLVCUAXIMCUCLK_in = PLVCUAXIMCUCLK;
  assign PLVCUBREADYAXILITEAPB_in = PLVCUBREADYAXILITEAPB;
  assign PLVCUDECARREADY0_in = PLVCUDECARREADY0;
  assign PLVCUDECARREADY1_in = PLVCUDECARREADY1;
  assign PLVCUDECAWREADY0_in = PLVCUDECAWREADY0;
  assign PLVCUDECAWREADY1_in = PLVCUDECAWREADY1;
  assign PLVCUDECBID0_in = PLVCUDECBID0;
  assign PLVCUDECBID1_in = PLVCUDECBID1;
  assign PLVCUDECBRESP0_in = PLVCUDECBRESP0;
  assign PLVCUDECBRESP1_in = PLVCUDECBRESP1;
  assign PLVCUDECBVALID0_in = PLVCUDECBVALID0;
  assign PLVCUDECBVALID1_in = PLVCUDECBVALID1;
  assign PLVCUDECRDATA0_in = PLVCUDECRDATA0;
  assign PLVCUDECRDATA1_in = PLVCUDECRDATA1;
  assign PLVCUDECRID0_in = PLVCUDECRID0;
  assign PLVCUDECRID1_in = PLVCUDECRID1;
  assign PLVCUDECRLAST0_in = PLVCUDECRLAST0;
  assign PLVCUDECRLAST1_in = PLVCUDECRLAST1;
  assign PLVCUDECRRESP0_in = PLVCUDECRRESP0;
  assign PLVCUDECRRESP1_in = PLVCUDECRRESP1;
  assign PLVCUDECRVALID0_in = PLVCUDECRVALID0;
  assign PLVCUDECRVALID1_in = PLVCUDECRVALID1;
  assign PLVCUDECWREADY0_in = PLVCUDECWREADY0;
  assign PLVCUDECWREADY1_in = PLVCUDECWREADY1;
  assign PLVCUENCALL2CRDATA_in = PLVCUENCALL2CRDATA;
  assign PLVCUENCALL2CRREADY_in = (PLVCUENCALL2CRREADY === 1'bz) || PLVCUENCALL2CRREADY; // rv 1
  assign PLVCUENCARREADY0_in = PLVCUENCARREADY0;
  assign PLVCUENCARREADY1_in = PLVCUENCARREADY1;
  assign PLVCUENCAWREADY0_in = PLVCUENCAWREADY0;
  assign PLVCUENCAWREADY1_in = PLVCUENCAWREADY1;
  assign PLVCUENCBID0_in = PLVCUENCBID0;
  assign PLVCUENCBID1_in = PLVCUENCBID1;
  assign PLVCUENCBRESP0_in = PLVCUENCBRESP0;
  assign PLVCUENCBRESP1_in = PLVCUENCBRESP1;
  assign PLVCUENCBVALID0_in = PLVCUENCBVALID0;
  assign PLVCUENCBVALID1_in = PLVCUENCBVALID1;
  assign PLVCUENCL2CCLK_in = PLVCUENCL2CCLK;
  assign PLVCUENCRDATA0_in = PLVCUENCRDATA0;
  assign PLVCUENCRDATA1_in = PLVCUENCRDATA1;
  assign PLVCUENCRID0_in = PLVCUENCRID0;
  assign PLVCUENCRID1_in = PLVCUENCRID1;
  assign PLVCUENCRLAST0_in = PLVCUENCRLAST0;
  assign PLVCUENCRLAST1_in = PLVCUENCRLAST1;
  assign PLVCUENCRRESP0_in = PLVCUENCRRESP0;
  assign PLVCUENCRRESP1_in = PLVCUENCRRESP1;
  assign PLVCUENCRVALID0_in = PLVCUENCRVALID0;
  assign PLVCUENCRVALID1_in = PLVCUENCRVALID1;
  assign PLVCUENCWREADY0_in = PLVCUENCWREADY0;
  assign PLVCUENCWREADY1_in = PLVCUENCWREADY1;
  assign PLVCUMCUMAXIICDCARREADY_in = PLVCUMCUMAXIICDCARREADY;
  assign PLVCUMCUMAXIICDCAWREADY_in = PLVCUMCUMAXIICDCAWREADY;
  assign PLVCUMCUMAXIICDCBID_in = PLVCUMCUMAXIICDCBID;
  assign PLVCUMCUMAXIICDCBRESP_in = PLVCUMCUMAXIICDCBRESP;
  assign PLVCUMCUMAXIICDCBVALID_in = PLVCUMCUMAXIICDCBVALID;
  assign PLVCUMCUMAXIICDCRDATA_in = PLVCUMCUMAXIICDCRDATA;
  assign PLVCUMCUMAXIICDCRID_in = PLVCUMCUMAXIICDCRID;
  assign PLVCUMCUMAXIICDCRLAST_in = PLVCUMCUMAXIICDCRLAST;
  assign PLVCUMCUMAXIICDCRRESP_in = PLVCUMCUMAXIICDCRRESP;
  assign PLVCUMCUMAXIICDCRVALID_in = PLVCUMCUMAXIICDCRVALID;
  assign PLVCUMCUMAXIICDCWREADY_in = PLVCUMCUMAXIICDCWREADY;
  assign PLVCURREADYAXILITEAPB_in = PLVCURREADYAXILITEAPB;
  assign PLVCUWDATAAXILITEAPB_in = PLVCUWDATAAXILITEAPB;
  assign PLVCUWSTRBAXILITEAPB_in = PLVCUWSTRBAXILITEAPB;
  assign PLVCUWVALIDAXILITEAPB_in = PLVCUWVALIDAXILITEAPB;
`endif
  assign INITPLVCUGASKETCLAMPCONTROLLVLSHVCCINTD_in = INITPLVCUGASKETCLAMPCONTROLLVLSHVCCINTD;
  assign PLVCUCORECLK_in = PLVCUCORECLK;
  assign PLVCUMCUCLK_in = PLVCUMCUCLK;
  assign PLVCUPLLREFCLKPL_in = PLVCUPLLREFCLKPL;
  assign PLVCURAWRSTN_in = PLVCURAWRSTN;
`ifndef XIL_XECLIB
  initial begin
    #1;
    trig_attr = ~trig_attr;
  end
`endif
`ifdef XIL_XECLIB
  assign CORECLKREQ_BIN = CORECLKREQ_REG[9:0];
  assign DECHORRESOLUTION_BIN = DECHORRESOLUTION_REG[13:0];
  assign DECODERCHROMAFORMAT_BIN =
      (DECODERCHROMAFORMAT_REG == "4_2_2") ? DECODERCHROMAFORMAT_4_2_2 :
      (DECODERCHROMAFORMAT_REG == "4_2_0") ? DECODERCHROMAFORMAT_4_2_0 :
       DECODERCHROMAFORMAT_4_2_2;
  assign DECODERCODING_BIN =
      (DECODERCODING_REG == "H.265") ? DECODERCODING_H_265 :
      (DECODERCODING_REG == "H.264") ? DECODERCODING_H_264 :
       DECODERCODING_H_265;
  assign DECODERCOLORDEPTH_BIN = DECODERCOLORDEPTH_REG[3:0];
  assign DECODERNUMCORES_BIN = DECODERNUMCORES_REG[1:0];
  assign DECVERTRESOLUTION_BIN = DECVERTRESOLUTION_REG[12:0];
  assign ENABLEDECODER_BIN =
      (ENABLEDECODER_REG == "TRUE") ? ENABLEDECODER_TRUE :
      (ENABLEDECODER_REG == "FALSE") ? ENABLEDECODER_FALSE :
       ENABLEDECODER_TRUE;
  assign ENABLEENCODER_BIN =
      (ENABLEENCODER_REG == "TRUE") ? ENABLEENCODER_TRUE :
      (ENABLEENCODER_REG == "FALSE") ? ENABLEENCODER_FALSE :
       ENABLEENCODER_TRUE;
  assign ENCHORRESOLUTION_BIN = ENCHORRESOLUTION_REG[13:0];
  assign ENCODERCHROMAFORMAT_BIN =
      (ENCODERCHROMAFORMAT_REG == "4_2_2") ? ENCODERCHROMAFORMAT_4_2_2 :
      (ENCODERCHROMAFORMAT_REG == "4_2_0") ? ENCODERCHROMAFORMAT_4_2_0 :
       ENCODERCHROMAFORMAT_4_2_2;
  assign ENCODERCODING_BIN =
      (ENCODERCODING_REG == "H.265") ? ENCODERCODING_H_265 :
      (ENCODERCODING_REG == "H.264") ? ENCODERCODING_H_264 :
       ENCODERCODING_H_265;
  assign ENCODERCOLORDEPTH_BIN = ENCODERCOLORDEPTH_REG[3:0];
  assign ENCODERNUMCORES_BIN = ENCODERNUMCORES_REG[2:0];
  assign ENCVERTRESOLUTION_BIN = ENCVERTRESOLUTION_REG[12:0];
`else
  always @ (trig_attr) begin
  #1;
  CORECLKREQ_BIN = CORECLKREQ_REG[9:0];
  DECHORRESOLUTION_BIN = DECHORRESOLUTION_REG[13:0];
  DECODERCHROMAFORMAT_BIN =
      (DECODERCHROMAFORMAT_REG == "4_2_2") ? DECODERCHROMAFORMAT_4_2_2 :
      (DECODERCHROMAFORMAT_REG == "4_2_0") ? DECODERCHROMAFORMAT_4_2_0 :
       DECODERCHROMAFORMAT_4_2_2;
  DECODERCODING_BIN =
      (DECODERCODING_REG == "H.265") ? DECODERCODING_H_265 :
      (DECODERCODING_REG == "H.264") ? DECODERCODING_H_264 :
       DECODERCODING_H_265;
  DECODERCOLORDEPTH_BIN = DECODERCOLORDEPTH_REG[3:0];
  DECODERNUMCORES_BIN = DECODERNUMCORES_REG[1:0];
  DECVERTRESOLUTION_BIN = DECVERTRESOLUTION_REG[12:0];
  ENABLEDECODER_BIN =
      (ENABLEDECODER_REG == "TRUE") ? ENABLEDECODER_TRUE :
      (ENABLEDECODER_REG == "FALSE") ? ENABLEDECODER_FALSE :
       ENABLEDECODER_TRUE;
  ENABLEENCODER_BIN =
      (ENABLEENCODER_REG == "TRUE") ? ENABLEENCODER_TRUE :
      (ENABLEENCODER_REG == "FALSE") ? ENABLEENCODER_FALSE :
       ENABLEENCODER_TRUE;
  ENCHORRESOLUTION_BIN = ENCHORRESOLUTION_REG[13:0];
  ENCODERCHROMAFORMAT_BIN =
      (ENCODERCHROMAFORMAT_REG == "4_2_2") ? ENCODERCHROMAFORMAT_4_2_2 :
      (ENCODERCHROMAFORMAT_REG == "4_2_0") ? ENCODERCHROMAFORMAT_4_2_0 :
       ENCODERCHROMAFORMAT_4_2_2;
  ENCODERCODING_BIN =
      (ENCODERCODING_REG == "H.265") ? ENCODERCODING_H_265 :
      (ENCODERCODING_REG == "H.264") ? ENCODERCODING_H_264 :
       ENCODERCODING_H_265;
  ENCODERCOLORDEPTH_BIN = ENCODERCOLORDEPTH_REG[3:0];
  ENCODERNUMCORES_BIN = ENCODERNUMCORES_REG[2:0];
  ENCVERTRESOLUTION_BIN = ENCVERTRESOLUTION_REG[12:0];
  end
`endif
`ifndef XIL_XECLIB
always @ (trig_attr) begin
  #1;
  if ((attr_test == 1'b1) ||
      ((CORECLKREQ_REG < 0) || (CORECLKREQ_REG > 667))) begin
    $display("Error: [Unisim %s-101] CORECLKREQ attribute is set to %d.  Legal values for this attribute are 0 to 667. Instance: %m", MODULE_NAME, CORECLKREQ_REG);
    attr_err = 1'b1;
  end
  if ((attr_test == 1'b1) ||
      ((DECHORRESOLUTION_REG < 320) || (DECHORRESOLUTION_REG > 8192))) begin
    $display("Error: [Unisim %s-102] DECHORRESOLUTION attribute is set to %d.  Legal values for this attribute are 320 to 8192. Instance: %m", MODULE_NAME, DECHORRESOLUTION_REG);
    attr_err = 1'b1;
  end
  if ((attr_test == 1'b1) ||
      ((DECODERCHROMAFORMAT_REG != "4_2_2") &&
       (DECODERCHROMAFORMAT_REG != "4_2_0"))) begin
    $display("Error: [Unisim %s-103] DECODERCHROMAFORMAT attribute is set to %s.  Legal values for this attribute are 4_2_2 or 4_2_0. Instance: %m", MODULE_NAME, DECODERCHROMAFORMAT_REG);
    attr_err = 1'b1;
  end
  if ((attr_test == 1'b1) ||
      ((DECODERCODING_REG != "H.265") &&
       (DECODERCODING_REG != "H.264"))) begin
    $display("Error: [Unisim %s-104] DECODERCODING attribute is set to %s.  Legal values for this attribute are H.265 or H.264. Instance: %m", MODULE_NAME, DECODERCODING_REG);
    attr_err = 1'b1;
  end
  if ((attr_test == 1'b1) ||
      ((DECODERCOLORDEPTH_REG != 10) &&
       (DECODERCOLORDEPTH_REG != 8))) begin
    $display("Error: [Unisim %s-105] DECODERCOLORDEPTH attribute is set to %d.  Legal values for this attribute are 10 or 8. Instance: %m", MODULE_NAME, DECODERCOLORDEPTH_REG);
    attr_err = 1'b1;
  end
  if ((attr_test == 1'b1) ||
      ((DECODERNUMCORES_REG < 1) || (DECODERNUMCORES_REG > 2))) begin
    $display("Error: [Unisim %s-106] DECODERNUMCORES attribute is set to %d.  Legal values for this attribute are 1 to 2. Instance: %m", MODULE_NAME, DECODERNUMCORES_REG);
    attr_err = 1'b1;
  end
  if ((attr_test == 1'b1) ||
      ((DECVERTRESOLUTION_REG < 240) || (DECVERTRESOLUTION_REG > 4352))) begin
    $display("Error: [Unisim %s-107] DECVERTRESOLUTION attribute is set to %d.  Legal values for this attribute are 240 to 4352. Instance: %m", MODULE_NAME, DECVERTRESOLUTION_REG);
    attr_err = 1'b1;
  end
  if ((attr_test == 1'b1) ||
      ((ENABLEDECODER_REG != "TRUE") &&
       (ENABLEDECODER_REG != "FALSE"))) begin
    $display("Error: [Unisim %s-108] ENABLEDECODER attribute is set to %s.  Legal values for this attribute are TRUE or FALSE. Instance: %m", MODULE_NAME, ENABLEDECODER_REG);
    attr_err = 1'b1;
  end
  if ((attr_test == 1'b1) ||
      ((ENABLEENCODER_REG != "TRUE") &&
       (ENABLEENCODER_REG != "FALSE"))) begin
    $display("Error: [Unisim %s-109] ENABLEENCODER attribute is set to %s.  Legal values for this attribute are TRUE or FALSE. Instance: %m", MODULE_NAME, ENABLEENCODER_REG);
    attr_err = 1'b1;
  end
  if ((attr_test == 1'b1) ||
      ((ENCHORRESOLUTION_REG < 320) || (ENCHORRESOLUTION_REG > 8192))) begin
    $display("Error: [Unisim %s-110] ENCHORRESOLUTION attribute is set to %d.  Legal values for this attribute are 320 to 8192. Instance: %m", MODULE_NAME, ENCHORRESOLUTION_REG);
    attr_err = 1'b1;
  end
  if ((attr_test == 1'b1) ||
      ((ENCODERCHROMAFORMAT_REG != "4_2_2") &&
       (ENCODERCHROMAFORMAT_REG != "4_2_0"))) begin
    $display("Error: [Unisim %s-111] ENCODERCHROMAFORMAT attribute is set to %s.  Legal values for this attribute are 4_2_2 or 4_2_0. Instance: %m", MODULE_NAME, ENCODERCHROMAFORMAT_REG);
    attr_err = 1'b1;
  end
  if ((attr_test == 1'b1) ||
      ((ENCODERCODING_REG != "H.265") &&
       (ENCODERCODING_REG != "H.264"))) begin
    $display("Error: [Unisim %s-112] ENCODERCODING attribute is set to %s.  Legal values for this attribute are H.265 or H.264. Instance: %m", MODULE_NAME, ENCODERCODING_REG);
    attr_err = 1'b1;
  end
  if ((attr_test == 1'b1) ||
      ((ENCODERCOLORDEPTH_REG != 10) &&
       (ENCODERCOLORDEPTH_REG != 8))) begin
    $display("Error: [Unisim %s-113] ENCODERCOLORDEPTH attribute is set to %d.  Legal values for this attribute are 10 or 8. Instance: %m", MODULE_NAME, ENCODERCOLORDEPTH_REG);
    attr_err = 1'b1;
  end
  if ((attr_test == 1'b1) ||
      ((ENCODERNUMCORES_REG < 1) || (ENCODERNUMCORES_REG > 4))) begin
    $display("Error: [Unisim %s-114] ENCODERNUMCORES attribute is set to %d.  Legal values for this attribute are 1 to 4. Instance: %m", MODULE_NAME, ENCODERNUMCORES_REG);
    attr_err = 1'b1;
  end
  if ((attr_test == 1'b1) ||
      ((ENCVERTRESOLUTION_REG < 240) || (ENCVERTRESOLUTION_REG > 4352))) begin
    $display("Error: [Unisim %s-115] ENCVERTRESOLUTION attribute is set to %d.  Legal values for this attribute are 240 to 4352. Instance: %m", MODULE_NAME, ENCVERTRESOLUTION_REG);
    attr_err = 1'b1;
  end
  if (attr_err == 1'b1) #1 $finish;
end
`endif
`ifndef XIL_XECLIB
`ifdef XIL_TIMING
  reg notifier;
`endif
  specify
    (PLVCUAXIDECCLK => VCUPLDECARADDR0[0]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARADDR0[10]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARADDR0[11]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARADDR0[12]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARADDR0[13]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARADDR0[14]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARADDR0[15]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARADDR0[16]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARADDR0[17]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARADDR0[18]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARADDR0[19]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARADDR0[1]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARADDR0[20]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARADDR0[21]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARADDR0[22]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARADDR0[23]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARADDR0[24]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARADDR0[25]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARADDR0[26]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARADDR0[27]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARADDR0[28]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARADDR0[29]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARADDR0[2]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARADDR0[30]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARADDR0[31]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARADDR0[32]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARADDR0[33]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARADDR0[34]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARADDR0[35]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARADDR0[36]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARADDR0[37]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARADDR0[38]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARADDR0[39]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARADDR0[3]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARADDR0[40]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARADDR0[41]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARADDR0[42]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARADDR0[43]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARADDR0[4]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARADDR0[5]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARADDR0[6]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARADDR0[7]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARADDR0[8]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARADDR0[9]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARADDR1[0]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARADDR1[10]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARADDR1[11]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARADDR1[12]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARADDR1[13]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARADDR1[14]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARADDR1[15]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARADDR1[16]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARADDR1[17]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARADDR1[18]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARADDR1[19]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARADDR1[1]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARADDR1[20]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARADDR1[21]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARADDR1[22]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARADDR1[23]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARADDR1[24]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARADDR1[25]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARADDR1[26]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARADDR1[27]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARADDR1[28]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARADDR1[29]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARADDR1[2]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARADDR1[30]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARADDR1[31]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARADDR1[32]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARADDR1[33]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARADDR1[34]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARADDR1[35]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARADDR1[36]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARADDR1[37]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARADDR1[38]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARADDR1[39]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARADDR1[3]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARADDR1[40]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARADDR1[41]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARADDR1[42]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARADDR1[43]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARADDR1[4]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARADDR1[5]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARADDR1[6]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARADDR1[7]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARADDR1[8]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARADDR1[9]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARBURST0[0]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARBURST0[1]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARBURST1[0]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARBURST1[1]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARCACHE0[0]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARCACHE0[1]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARCACHE0[2]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARCACHE0[3]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARCACHE1[0]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARCACHE1[1]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARCACHE1[2]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARCACHE1[3]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARID0[0]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARID0[1]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARID0[2]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARID0[3]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARID1[0]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARID1[1]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARID1[2]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARID1[3]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARLEN0[0]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARLEN0[1]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARLEN0[2]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARLEN0[3]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARLEN0[4]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARLEN0[5]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARLEN0[6]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARLEN0[7]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARLEN1[0]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARLEN1[1]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARLEN1[2]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARLEN1[3]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARLEN1[4]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARLEN1[5]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARLEN1[6]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARLEN1[7]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARPROT0) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARPROT1) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARQOS0[0]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARQOS0[1]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARQOS0[2]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARQOS0[3]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARQOS1[0]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARQOS1[1]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARQOS1[2]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARQOS1[3]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARSIZE0[0]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARSIZE0[1]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARSIZE0[2]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARSIZE1[0]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARSIZE1[1]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARSIZE1[2]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARVALID0) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECARVALID1) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWADDR0[0]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWADDR0[10]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWADDR0[11]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWADDR0[12]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWADDR0[13]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWADDR0[14]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWADDR0[15]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWADDR0[16]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWADDR0[17]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWADDR0[18]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWADDR0[19]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWADDR0[1]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWADDR0[20]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWADDR0[21]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWADDR0[22]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWADDR0[23]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWADDR0[24]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWADDR0[25]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWADDR0[26]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWADDR0[27]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWADDR0[28]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWADDR0[29]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWADDR0[2]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWADDR0[30]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWADDR0[31]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWADDR0[32]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWADDR0[33]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWADDR0[34]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWADDR0[35]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWADDR0[36]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWADDR0[37]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWADDR0[38]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWADDR0[39]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWADDR0[3]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWADDR0[40]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWADDR0[41]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWADDR0[42]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWADDR0[43]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWADDR0[4]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWADDR0[5]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWADDR0[6]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWADDR0[7]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWADDR0[8]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWADDR0[9]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWADDR1[0]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWADDR1[10]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWADDR1[11]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWADDR1[12]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWADDR1[13]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWADDR1[14]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWADDR1[15]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWADDR1[16]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWADDR1[17]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWADDR1[18]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWADDR1[19]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWADDR1[1]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWADDR1[20]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWADDR1[21]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWADDR1[22]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWADDR1[23]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWADDR1[24]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWADDR1[25]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWADDR1[26]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWADDR1[27]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWADDR1[28]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWADDR1[29]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWADDR1[2]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWADDR1[30]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWADDR1[31]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWADDR1[32]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWADDR1[33]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWADDR1[34]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWADDR1[35]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWADDR1[36]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWADDR1[37]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWADDR1[38]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWADDR1[39]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWADDR1[3]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWADDR1[40]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWADDR1[41]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWADDR1[42]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWADDR1[43]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWADDR1[4]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWADDR1[5]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWADDR1[6]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWADDR1[7]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWADDR1[8]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWADDR1[9]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWBURST0[0]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWBURST0[1]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWBURST1[0]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWBURST1[1]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWCACHE0[0]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWCACHE0[1]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWCACHE0[2]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWCACHE0[3]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWCACHE1[0]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWCACHE1[1]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWCACHE1[2]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWCACHE1[3]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWID0[0]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWID0[1]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWID0[2]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWID0[3]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWID1[0]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWID1[1]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWID1[2]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWID1[3]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWLEN0[0]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWLEN0[1]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWLEN0[2]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWLEN0[3]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWLEN0[4]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWLEN0[5]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWLEN0[6]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWLEN0[7]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWLEN1[0]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWLEN1[1]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWLEN1[2]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWLEN1[3]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWLEN1[4]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWLEN1[5]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWLEN1[6]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWLEN1[7]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWPROT0) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWPROT1) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWQOS0[0]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWQOS0[1]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWQOS0[2]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWQOS0[3]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWQOS1[0]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWQOS1[1]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWQOS1[2]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWQOS1[3]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWSIZE0[0]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWSIZE0[1]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWSIZE0[2]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWSIZE1[0]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWSIZE1[1]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWSIZE1[2]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWVALID0) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECAWVALID1) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECBREADY0) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECBREADY1) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECRREADY0) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECRREADY1) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[0]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[100]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[101]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[102]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[103]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[104]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[105]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[106]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[107]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[108]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[109]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[10]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[110]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[111]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[112]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[113]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[114]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[115]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[116]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[117]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[118]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[119]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[11]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[120]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[121]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[122]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[123]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[124]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[125]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[126]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[127]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[12]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[13]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[14]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[15]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[16]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[17]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[18]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[19]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[1]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[20]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[21]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[22]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[23]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[24]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[25]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[26]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[27]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[28]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[29]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[2]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[30]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[31]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[32]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[33]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[34]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[35]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[36]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[37]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[38]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[39]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[3]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[40]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[41]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[42]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[43]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[44]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[45]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[46]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[47]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[48]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[49]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[4]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[50]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[51]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[52]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[53]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[54]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[55]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[56]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[57]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[58]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[59]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[5]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[60]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[61]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[62]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[63]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[64]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[65]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[66]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[67]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[68]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[69]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[6]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[70]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[71]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[72]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[73]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[74]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[75]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[76]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[77]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[78]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[79]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[7]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[80]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[81]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[82]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[83]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[84]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[85]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[86]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[87]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[88]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[89]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[8]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[90]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[91]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[92]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[93]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[94]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[95]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[96]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[97]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[98]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[99]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA0[9]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[0]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[100]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[101]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[102]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[103]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[104]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[105]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[106]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[107]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[108]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[109]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[10]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[110]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[111]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[112]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[113]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[114]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[115]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[116]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[117]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[118]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[119]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[11]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[120]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[121]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[122]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[123]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[124]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[125]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[126]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[127]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[12]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[13]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[14]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[15]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[16]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[17]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[18]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[19]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[1]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[20]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[21]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[22]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[23]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[24]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[25]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[26]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[27]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[28]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[29]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[2]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[30]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[31]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[32]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[33]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[34]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[35]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[36]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[37]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[38]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[39]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[3]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[40]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[41]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[42]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[43]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[44]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[45]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[46]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[47]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[48]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[49]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[4]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[50]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[51]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[52]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[53]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[54]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[55]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[56]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[57]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[58]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[59]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[5]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[60]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[61]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[62]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[63]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[64]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[65]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[66]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[67]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[68]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[69]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[6]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[70]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[71]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[72]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[73]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[74]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[75]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[76]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[77]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[78]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[79]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[7]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[80]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[81]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[82]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[83]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[84]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[85]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[86]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[87]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[88]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[89]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[8]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[90]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[91]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[92]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[93]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[94]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[95]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[96]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[97]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[98]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[99]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWDATA1[9]) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWLAST0) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWLAST1) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWVALID0) = (100:100:100, 100:100:100);
    (PLVCUAXIDECCLK => VCUPLDECWVALID1) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARADDR0[0]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARADDR0[10]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARADDR0[11]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARADDR0[12]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARADDR0[13]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARADDR0[14]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARADDR0[15]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARADDR0[16]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARADDR0[17]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARADDR0[18]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARADDR0[19]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARADDR0[1]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARADDR0[20]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARADDR0[21]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARADDR0[22]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARADDR0[23]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARADDR0[24]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARADDR0[25]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARADDR0[26]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARADDR0[27]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARADDR0[28]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARADDR0[29]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARADDR0[2]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARADDR0[30]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARADDR0[31]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARADDR0[32]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARADDR0[33]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARADDR0[34]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARADDR0[35]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARADDR0[36]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARADDR0[37]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARADDR0[38]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARADDR0[39]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARADDR0[3]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARADDR0[40]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARADDR0[41]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARADDR0[42]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARADDR0[43]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARADDR0[4]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARADDR0[5]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARADDR0[6]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARADDR0[7]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARADDR0[8]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARADDR0[9]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARADDR1[0]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARADDR1[10]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARADDR1[11]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARADDR1[12]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARADDR1[13]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARADDR1[14]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARADDR1[15]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARADDR1[16]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARADDR1[17]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARADDR1[18]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARADDR1[19]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARADDR1[1]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARADDR1[20]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARADDR1[21]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARADDR1[22]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARADDR1[23]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARADDR1[24]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARADDR1[25]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARADDR1[26]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARADDR1[27]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARADDR1[28]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARADDR1[29]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARADDR1[2]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARADDR1[30]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARADDR1[31]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARADDR1[32]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARADDR1[33]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARADDR1[34]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARADDR1[35]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARADDR1[36]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARADDR1[37]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARADDR1[38]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARADDR1[39]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARADDR1[3]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARADDR1[40]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARADDR1[41]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARADDR1[42]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARADDR1[43]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARADDR1[4]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARADDR1[5]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARADDR1[6]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARADDR1[7]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARADDR1[8]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARADDR1[9]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARBURST0[0]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARBURST0[1]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARBURST1[0]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARBURST1[1]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARCACHE0[0]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARCACHE0[1]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARCACHE0[2]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARCACHE0[3]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARCACHE1[0]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARCACHE1[1]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARCACHE1[2]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARCACHE1[3]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARID0[0]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARID0[1]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARID0[2]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARID0[3]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARID1[0]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARID1[1]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARID1[2]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARID1[3]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARLEN0[0]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARLEN0[1]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARLEN0[2]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARLEN0[3]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARLEN0[4]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARLEN0[5]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARLEN0[6]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARLEN0[7]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARLEN1[0]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARLEN1[1]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARLEN1[2]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARLEN1[3]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARLEN1[4]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARLEN1[5]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARLEN1[6]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARLEN1[7]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARPROT0) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARPROT1) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARQOS0[0]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARQOS0[1]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARQOS0[2]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARQOS0[3]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARQOS1[0]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARQOS1[1]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARQOS1[2]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARQOS1[3]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARSIZE0[0]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARSIZE0[1]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARSIZE0[2]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARSIZE1[0]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARSIZE1[1]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARSIZE1[2]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARVALID0) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCARVALID1) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWADDR0[0]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWADDR0[10]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWADDR0[11]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWADDR0[12]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWADDR0[13]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWADDR0[14]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWADDR0[15]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWADDR0[16]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWADDR0[17]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWADDR0[18]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWADDR0[19]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWADDR0[1]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWADDR0[20]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWADDR0[21]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWADDR0[22]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWADDR0[23]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWADDR0[24]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWADDR0[25]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWADDR0[26]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWADDR0[27]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWADDR0[28]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWADDR0[29]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWADDR0[2]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWADDR0[30]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWADDR0[31]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWADDR0[32]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWADDR0[33]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWADDR0[34]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWADDR0[35]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWADDR0[36]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWADDR0[37]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWADDR0[38]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWADDR0[39]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWADDR0[3]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWADDR0[40]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWADDR0[41]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWADDR0[42]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWADDR0[43]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWADDR0[4]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWADDR0[5]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWADDR0[6]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWADDR0[7]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWADDR0[8]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWADDR0[9]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWADDR1[0]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWADDR1[10]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWADDR1[11]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWADDR1[12]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWADDR1[13]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWADDR1[14]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWADDR1[15]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWADDR1[16]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWADDR1[17]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWADDR1[18]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWADDR1[19]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWADDR1[1]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWADDR1[20]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWADDR1[21]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWADDR1[22]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWADDR1[23]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWADDR1[24]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWADDR1[25]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWADDR1[26]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWADDR1[27]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWADDR1[28]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWADDR1[29]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWADDR1[2]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWADDR1[30]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWADDR1[31]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWADDR1[32]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWADDR1[33]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWADDR1[34]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWADDR1[35]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWADDR1[36]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWADDR1[37]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWADDR1[38]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWADDR1[39]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWADDR1[3]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWADDR1[40]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWADDR1[41]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWADDR1[42]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWADDR1[43]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWADDR1[4]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWADDR1[5]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWADDR1[6]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWADDR1[7]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWADDR1[8]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWADDR1[9]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWBURST0[0]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWBURST0[1]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWBURST1[0]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWBURST1[1]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWCACHE0[0]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWCACHE0[1]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWCACHE0[2]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWCACHE0[3]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWCACHE1[0]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWCACHE1[1]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWCACHE1[2]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWCACHE1[3]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWID0[0]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWID0[1]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWID0[2]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWID0[3]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWID1[0]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWID1[1]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWID1[2]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWID1[3]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWLEN0[0]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWLEN0[1]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWLEN0[2]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWLEN0[3]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWLEN0[4]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWLEN0[5]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWLEN0[6]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWLEN0[7]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWLEN1[0]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWLEN1[1]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWLEN1[2]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWLEN1[3]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWLEN1[4]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWLEN1[5]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWLEN1[6]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWLEN1[7]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWPROT0) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWPROT1) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWQOS0[0]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWQOS0[1]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWQOS0[2]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWQOS0[3]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWQOS1[0]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWQOS1[1]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWQOS1[2]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWQOS1[3]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWSIZE0[0]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWSIZE0[1]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWSIZE0[2]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWSIZE1[0]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWSIZE1[1]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWSIZE1[2]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWVALID0) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCAWVALID1) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCBREADY0) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCBREADY1) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCRREADY0) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCRREADY1) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[0]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[100]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[101]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[102]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[103]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[104]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[105]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[106]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[107]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[108]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[109]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[10]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[110]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[111]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[112]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[113]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[114]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[115]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[116]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[117]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[118]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[119]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[11]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[120]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[121]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[122]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[123]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[124]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[125]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[126]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[127]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[12]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[13]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[14]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[15]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[16]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[17]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[18]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[19]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[1]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[20]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[21]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[22]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[23]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[24]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[25]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[26]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[27]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[28]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[29]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[2]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[30]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[31]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[32]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[33]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[34]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[35]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[36]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[37]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[38]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[39]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[3]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[40]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[41]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[42]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[43]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[44]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[45]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[46]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[47]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[48]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[49]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[4]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[50]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[51]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[52]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[53]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[54]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[55]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[56]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[57]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[58]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[59]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[5]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[60]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[61]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[62]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[63]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[64]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[65]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[66]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[67]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[68]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[69]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[6]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[70]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[71]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[72]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[73]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[74]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[75]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[76]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[77]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[78]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[79]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[7]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[80]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[81]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[82]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[83]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[84]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[85]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[86]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[87]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[88]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[89]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[8]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[90]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[91]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[92]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[93]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[94]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[95]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[96]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[97]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[98]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[99]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA0[9]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[0]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[100]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[101]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[102]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[103]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[104]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[105]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[106]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[107]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[108]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[109]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[10]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[110]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[111]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[112]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[113]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[114]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[115]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[116]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[117]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[118]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[119]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[11]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[120]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[121]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[122]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[123]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[124]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[125]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[126]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[127]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[12]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[13]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[14]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[15]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[16]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[17]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[18]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[19]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[1]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[20]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[21]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[22]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[23]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[24]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[25]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[26]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[27]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[28]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[29]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[2]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[30]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[31]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[32]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[33]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[34]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[35]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[36]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[37]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[38]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[39]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[3]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[40]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[41]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[42]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[43]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[44]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[45]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[46]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[47]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[48]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[49]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[4]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[50]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[51]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[52]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[53]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[54]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[55]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[56]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[57]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[58]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[59]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[5]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[60]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[61]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[62]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[63]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[64]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[65]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[66]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[67]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[68]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[69]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[6]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[70]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[71]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[72]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[73]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[74]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[75]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[76]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[77]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[78]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[79]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[7]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[80]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[81]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[82]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[83]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[84]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[85]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[86]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[87]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[88]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[89]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[8]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[90]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[91]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[92]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[93]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[94]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[95]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[96]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[97]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[98]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[99]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWDATA1[9]) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWLAST0) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWLAST1) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWVALID0) = (100:100:100, 100:100:100);
    (PLVCUAXIENCCLK => VCUPLENCWVALID1) = (100:100:100, 100:100:100);
    (PLVCUAXILITECLK => VCUPLARREADYAXILITEAPB) = (100:100:100, 100:100:100);
    (PLVCUAXILITECLK => VCUPLAWREADYAXILITEAPB) = (100:100:100, 100:100:100);
    (PLVCUAXILITECLK => VCUPLBRESPAXILITEAPB[0]) = (100:100:100, 100:100:100);
    (PLVCUAXILITECLK => VCUPLBRESPAXILITEAPB[1]) = (100:100:100, 100:100:100);
    (PLVCUAXILITECLK => VCUPLBVALIDAXILITEAPB) = (100:100:100, 100:100:100);
    (PLVCUAXILITECLK => VCUPLPINTREQ) = (100:100:100, 100:100:100);
    (PLVCUAXILITECLK => VCUPLRDATAAXILITEAPB[0]) = (100:100:100, 100:100:100);
    (PLVCUAXILITECLK => VCUPLRDATAAXILITEAPB[10]) = (100:100:100, 100:100:100);
    (PLVCUAXILITECLK => VCUPLRDATAAXILITEAPB[11]) = (100:100:100, 100:100:100);
    (PLVCUAXILITECLK => VCUPLRDATAAXILITEAPB[12]) = (100:100:100, 100:100:100);
    (PLVCUAXILITECLK => VCUPLRDATAAXILITEAPB[13]) = (100:100:100, 100:100:100);
    (PLVCUAXILITECLK => VCUPLRDATAAXILITEAPB[14]) = (100:100:100, 100:100:100);
    (PLVCUAXILITECLK => VCUPLRDATAAXILITEAPB[15]) = (100:100:100, 100:100:100);
    (PLVCUAXILITECLK => VCUPLRDATAAXILITEAPB[16]) = (100:100:100, 100:100:100);
    (PLVCUAXILITECLK => VCUPLRDATAAXILITEAPB[17]) = (100:100:100, 100:100:100);
    (PLVCUAXILITECLK => VCUPLRDATAAXILITEAPB[18]) = (100:100:100, 100:100:100);
    (PLVCUAXILITECLK => VCUPLRDATAAXILITEAPB[19]) = (100:100:100, 100:100:100);
    (PLVCUAXILITECLK => VCUPLRDATAAXILITEAPB[1]) = (100:100:100, 100:100:100);
    (PLVCUAXILITECLK => VCUPLRDATAAXILITEAPB[20]) = (100:100:100, 100:100:100);
    (PLVCUAXILITECLK => VCUPLRDATAAXILITEAPB[21]) = (100:100:100, 100:100:100);
    (PLVCUAXILITECLK => VCUPLRDATAAXILITEAPB[22]) = (100:100:100, 100:100:100);
    (PLVCUAXILITECLK => VCUPLRDATAAXILITEAPB[23]) = (100:100:100, 100:100:100);
    (PLVCUAXILITECLK => VCUPLRDATAAXILITEAPB[24]) = (100:100:100, 100:100:100);
    (PLVCUAXILITECLK => VCUPLRDATAAXILITEAPB[25]) = (100:100:100, 100:100:100);
    (PLVCUAXILITECLK => VCUPLRDATAAXILITEAPB[26]) = (100:100:100, 100:100:100);
    (PLVCUAXILITECLK => VCUPLRDATAAXILITEAPB[27]) = (100:100:100, 100:100:100);
    (PLVCUAXILITECLK => VCUPLRDATAAXILITEAPB[28]) = (100:100:100, 100:100:100);
    (PLVCUAXILITECLK => VCUPLRDATAAXILITEAPB[29]) = (100:100:100, 100:100:100);
    (PLVCUAXILITECLK => VCUPLRDATAAXILITEAPB[2]) = (100:100:100, 100:100:100);
    (PLVCUAXILITECLK => VCUPLRDATAAXILITEAPB[30]) = (100:100:100, 100:100:100);
    (PLVCUAXILITECLK => VCUPLRDATAAXILITEAPB[31]) = (100:100:100, 100:100:100);
    (PLVCUAXILITECLK => VCUPLRDATAAXILITEAPB[3]) = (100:100:100, 100:100:100);
    (PLVCUAXILITECLK => VCUPLRDATAAXILITEAPB[4]) = (100:100:100, 100:100:100);
    (PLVCUAXILITECLK => VCUPLRDATAAXILITEAPB[5]) = (100:100:100, 100:100:100);
    (PLVCUAXILITECLK => VCUPLRDATAAXILITEAPB[6]) = (100:100:100, 100:100:100);
    (PLVCUAXILITECLK => VCUPLRDATAAXILITEAPB[7]) = (100:100:100, 100:100:100);
    (PLVCUAXILITECLK => VCUPLRDATAAXILITEAPB[8]) = (100:100:100, 100:100:100);
    (PLVCUAXILITECLK => VCUPLRDATAAXILITEAPB[9]) = (100:100:100, 100:100:100);
    (PLVCUAXILITECLK => VCUPLRRESPAXILITEAPB[0]) = (100:100:100, 100:100:100);
    (PLVCUAXILITECLK => VCUPLRRESPAXILITEAPB[1]) = (100:100:100, 100:100:100);
    (PLVCUAXILITECLK => VCUPLRVALIDAXILITEAPB) = (100:100:100, 100:100:100);
    (PLVCUAXILITECLK => VCUPLWREADYAXILITEAPB) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCARADDR[0]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCARADDR[10]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCARADDR[11]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCARADDR[12]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCARADDR[13]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCARADDR[14]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCARADDR[15]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCARADDR[16]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCARADDR[17]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCARADDR[18]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCARADDR[19]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCARADDR[1]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCARADDR[20]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCARADDR[21]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCARADDR[22]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCARADDR[23]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCARADDR[24]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCARADDR[25]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCARADDR[26]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCARADDR[27]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCARADDR[28]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCARADDR[29]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCARADDR[2]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCARADDR[30]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCARADDR[31]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCARADDR[32]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCARADDR[33]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCARADDR[34]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCARADDR[35]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCARADDR[36]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCARADDR[37]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCARADDR[38]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCARADDR[39]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCARADDR[3]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCARADDR[40]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCARADDR[41]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCARADDR[42]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCARADDR[43]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCARADDR[4]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCARADDR[5]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCARADDR[6]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCARADDR[7]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCARADDR[8]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCARADDR[9]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCARBURST[0]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCARBURST[1]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCARCACHE[0]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCARCACHE[1]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCARCACHE[2]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCARCACHE[3]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCARID[0]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCARID[1]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCARID[2]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCARLEN[0]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCARLEN[1]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCARLEN[2]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCARLEN[3]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCARLEN[4]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCARLEN[5]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCARLEN[6]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCARLEN[7]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCARLOCK) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCARPROT[0]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCARPROT[1]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCARPROT[2]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCARQOS[0]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCARQOS[1]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCARQOS[2]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCARQOS[3]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCARSIZE[0]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCARSIZE[1]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCARSIZE[2]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCARVALID) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCAWADDR[0]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCAWADDR[10]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCAWADDR[11]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCAWADDR[12]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCAWADDR[13]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCAWADDR[14]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCAWADDR[15]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCAWADDR[16]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCAWADDR[17]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCAWADDR[18]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCAWADDR[19]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCAWADDR[1]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCAWADDR[20]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCAWADDR[21]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCAWADDR[22]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCAWADDR[23]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCAWADDR[24]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCAWADDR[25]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCAWADDR[26]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCAWADDR[27]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCAWADDR[28]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCAWADDR[29]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCAWADDR[2]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCAWADDR[30]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCAWADDR[31]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCAWADDR[32]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCAWADDR[33]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCAWADDR[34]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCAWADDR[35]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCAWADDR[36]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCAWADDR[37]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCAWADDR[38]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCAWADDR[39]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCAWADDR[3]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCAWADDR[40]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCAWADDR[41]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCAWADDR[42]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCAWADDR[43]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCAWADDR[4]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCAWADDR[5]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCAWADDR[6]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCAWADDR[7]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCAWADDR[8]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCAWADDR[9]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCAWBURST[0]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCAWBURST[1]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCAWCACHE[0]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCAWCACHE[1]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCAWCACHE[2]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCAWCACHE[3]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCAWID[0]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCAWID[1]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCAWID[2]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCAWLEN[0]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCAWLEN[1]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCAWLEN[2]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCAWLEN[3]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCAWLEN[4]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCAWLEN[5]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCAWLEN[6]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCAWLEN[7]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCAWLOCK) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCAWPROT[0]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCAWPROT[1]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCAWPROT[2]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCAWQOS[0]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCAWQOS[1]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCAWQOS[2]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCAWQOS[3]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCAWSIZE[0]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCAWSIZE[1]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCAWSIZE[2]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCAWVALID) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCBREADY) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCRREADY) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCWDATA[0]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCWDATA[10]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCWDATA[11]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCWDATA[12]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCWDATA[13]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCWDATA[14]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCWDATA[15]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCWDATA[16]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCWDATA[17]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCWDATA[18]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCWDATA[19]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCWDATA[1]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCWDATA[20]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCWDATA[21]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCWDATA[22]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCWDATA[23]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCWDATA[24]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCWDATA[25]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCWDATA[26]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCWDATA[27]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCWDATA[28]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCWDATA[29]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCWDATA[2]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCWDATA[30]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCWDATA[31]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCWDATA[3]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCWDATA[4]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCWDATA[5]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCWDATA[6]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCWDATA[7]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCWDATA[8]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCWDATA[9]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCWLAST) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCWSTRB[0]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCWSTRB[1]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCWSTRB[2]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCWSTRB[3]) = (100:100:100, 100:100:100);
    (PLVCUAXIMCUCLK => VCUPLMCUMAXIICDCWVALID) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CADDR[0]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CADDR[10]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CADDR[11]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CADDR[12]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CADDR[13]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CADDR[14]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CADDR[15]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CADDR[16]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CADDR[1]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CADDR[2]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CADDR[3]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CADDR[4]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CADDR[5]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CADDR[6]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CADDR[7]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CADDR[8]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CADDR[9]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CRVALID) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[0]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[100]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[101]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[102]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[103]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[104]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[105]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[106]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[107]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[108]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[109]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[10]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[110]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[111]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[112]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[113]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[114]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[115]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[116]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[117]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[118]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[119]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[11]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[120]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[121]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[122]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[123]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[124]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[125]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[126]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[127]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[128]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[129]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[12]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[130]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[131]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[132]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[133]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[134]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[135]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[136]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[137]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[138]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[139]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[13]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[140]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[141]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[142]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[143]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[144]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[145]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[146]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[147]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[148]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[149]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[14]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[150]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[151]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[152]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[153]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[154]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[155]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[156]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[157]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[158]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[159]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[15]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[160]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[161]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[162]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[163]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[164]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[165]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[166]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[167]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[168]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[169]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[16]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[170]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[171]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[172]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[173]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[174]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[175]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[176]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[177]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[178]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[179]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[17]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[180]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[181]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[182]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[183]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[184]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[185]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[186]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[187]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[188]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[189]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[18]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[190]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[191]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[192]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[193]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[194]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[195]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[196]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[197]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[198]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[199]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[19]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[1]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[200]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[201]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[202]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[203]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[204]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[205]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[206]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[207]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[208]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[209]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[20]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[210]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[211]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[212]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[213]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[214]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[215]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[216]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[217]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[218]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[219]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[21]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[220]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[221]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[222]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[223]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[224]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[225]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[226]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[227]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[228]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[229]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[22]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[230]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[231]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[232]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[233]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[234]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[235]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[236]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[237]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[238]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[239]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[23]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[240]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[241]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[242]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[243]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[244]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[245]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[246]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[247]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[248]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[249]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[24]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[250]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[251]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[252]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[253]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[254]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[255]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[256]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[257]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[258]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[259]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[25]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[260]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[261]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[262]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[263]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[264]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[265]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[266]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[267]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[268]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[269]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[26]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[270]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[271]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[272]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[273]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[274]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[275]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[276]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[277]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[278]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[279]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[27]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[280]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[281]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[282]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[283]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[284]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[285]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[286]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[287]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[288]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[289]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[28]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[290]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[291]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[292]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[293]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[294]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[295]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[296]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[297]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[298]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[299]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[29]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[2]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[300]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[301]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[302]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[303]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[304]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[305]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[306]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[307]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[308]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[309]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[30]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[310]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[311]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[312]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[313]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[314]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[315]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[316]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[317]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[318]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[319]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[31]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[32]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[33]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[34]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[35]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[36]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[37]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[38]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[39]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[3]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[40]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[41]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[42]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[43]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[44]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[45]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[46]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[47]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[48]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[49]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[4]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[50]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[51]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[52]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[53]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[54]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[55]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[56]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[57]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[58]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[59]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[5]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[60]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[61]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[62]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[63]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[64]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[65]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[66]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[67]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[68]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[69]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[6]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[70]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[71]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[72]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[73]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[74]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[75]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[76]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[77]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[78]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[79]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[7]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[80]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[81]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[82]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[83]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[84]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[85]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[86]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[87]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[88]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[89]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[8]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[90]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[91]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[92]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[93]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[94]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[95]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[96]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[97]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[98]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[99]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWDATA[9]) = (100:100:100, 100:100:100);
    (PLVCUENCL2CCLK => VCUPLENCALL2CWVALID) = (100:100:100, 100:100:100);
`ifdef XIL_TIMING
    $period (negedge PLVCUAXIDECCLK, 0:0:0, notifier);
    $period (negedge PLVCUAXIENCCLK, 0:0:0, notifier);
    $period (negedge PLVCUAXILITECLK, 0:0:0, notifier);
    $period (negedge PLVCUAXIMCUCLK, 0:0:0, notifier);
    $period (negedge PLVCUCORECLK, 0:0:0, notifier);
    $period (negedge PLVCUENCL2CCLK, 0:0:0, notifier);
    $period (negedge PLVCUMCUCLK, 0:0:0, notifier);
    $period (negedge PLVCUPLLREFCLKPL, 0:0:0, notifier);
    $period (negedge VCUPLCORESTATUSCLKPLL, 0:0:0, notifier);
    $period (negedge VCUPLMCUSTATUSCLKPLL, 0:0:0, notifier);
    $period (posedge PLVCUAXIDECCLK, 0:0:0, notifier);
    $period (posedge PLVCUAXIENCCLK, 0:0:0, notifier);
    $period (posedge PLVCUAXILITECLK, 0:0:0, notifier);
    $period (posedge PLVCUAXIMCUCLK, 0:0:0, notifier);
    $period (posedge PLVCUCORECLK, 0:0:0, notifier);
    $period (posedge PLVCUENCL2CCLK, 0:0:0, notifier);
    $period (posedge PLVCUMCUCLK, 0:0:0, notifier);
    $period (posedge PLVCUPLLREFCLKPL, 0:0:0, notifier);
    $period (posedge VCUPLCORESTATUSCLKPLL, 0:0:0, notifier);
    $period (posedge VCUPLMCUSTATUSCLKPLL, 0:0:0, notifier);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECARREADY0, 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECARREADY0_delay);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECARREADY1, 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECARREADY1_delay);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECAWREADY0, 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECAWREADY0_delay);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECAWREADY1, 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECAWREADY1_delay);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECBID0[0], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECBID0_delay[0]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECBID0[1], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECBID0_delay[1]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECBID0[2], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECBID0_delay[2]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECBID0[3], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECBID0_delay[3]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECBID1[0], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECBID1_delay[0]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECBID1[1], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECBID1_delay[1]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECBID1[2], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECBID1_delay[2]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECBID1[3], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECBID1_delay[3]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECBRESP0[1], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECBRESP0_delay[1]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECBRESP1[1], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECBRESP1_delay[1]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECBVALID0, 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECBVALID0_delay);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECBVALID1, 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECBVALID1_delay);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[0], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[0]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[100], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[100]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[101], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[101]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[102], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[102]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[103], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[103]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[104], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[104]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[105], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[105]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[106], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[106]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[107], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[107]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[108], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[108]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[109], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[109]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[10], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[10]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[110], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[110]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[111], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[111]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[112], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[112]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[113], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[113]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[114], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[114]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[115], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[115]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[116], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[116]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[117], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[117]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[118], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[118]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[119], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[119]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[11], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[11]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[120], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[120]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[121], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[121]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[122], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[122]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[123], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[123]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[124], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[124]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[125], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[125]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[126], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[126]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[127], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[127]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[12], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[12]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[13], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[13]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[14], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[14]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[15], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[15]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[16], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[16]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[17], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[17]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[18], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[18]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[19], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[19]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[1], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[1]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[20], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[20]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[21], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[21]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[22], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[22]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[23], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[23]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[24], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[24]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[25], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[25]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[26], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[26]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[27], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[27]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[28], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[28]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[29], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[29]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[2], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[2]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[30], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[30]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[31], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[31]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[32], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[32]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[33], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[33]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[34], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[34]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[35], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[35]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[36], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[36]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[37], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[37]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[38], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[38]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[39], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[39]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[3], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[3]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[40], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[40]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[41], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[41]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[42], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[42]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[43], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[43]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[44], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[44]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[45], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[45]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[46], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[46]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[47], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[47]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[48], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[48]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[49], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[49]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[4], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[4]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[50], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[50]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[51], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[51]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[52], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[52]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[53], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[53]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[54], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[54]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[55], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[55]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[56], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[56]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[57], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[57]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[58], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[58]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[59], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[59]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[5], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[5]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[60], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[60]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[61], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[61]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[62], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[62]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[63], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[63]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[64], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[64]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[65], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[65]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[66], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[66]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[67], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[67]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[68], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[68]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[69], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[69]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[6], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[6]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[70], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[70]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[71], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[71]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[72], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[72]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[73], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[73]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[74], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[74]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[75], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[75]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[76], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[76]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[77], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[77]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[78], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[78]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[79], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[79]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[7], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[7]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[80], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[80]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[81], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[81]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[82], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[82]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[83], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[83]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[84], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[84]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[85], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[85]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[86], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[86]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[87], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[87]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[88], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[88]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[89], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[89]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[8], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[8]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[90], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[90]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[91], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[91]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[92], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[92]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[93], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[93]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[94], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[94]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[95], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[95]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[96], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[96]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[97], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[97]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[98], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[98]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[99], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[99]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA0[9], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[9]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[0], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[0]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[100], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[100]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[101], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[101]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[102], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[102]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[103], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[103]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[104], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[104]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[105], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[105]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[106], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[106]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[107], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[107]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[108], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[108]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[109], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[109]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[10], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[10]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[110], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[110]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[111], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[111]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[112], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[112]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[113], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[113]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[114], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[114]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[115], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[115]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[116], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[116]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[117], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[117]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[118], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[118]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[119], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[119]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[11], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[11]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[120], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[120]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[121], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[121]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[122], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[122]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[123], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[123]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[124], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[124]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[125], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[125]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[126], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[126]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[127], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[127]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[12], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[12]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[13], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[13]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[14], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[14]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[15], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[15]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[16], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[16]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[17], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[17]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[18], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[18]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[19], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[19]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[1], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[1]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[20], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[20]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[21], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[21]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[22], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[22]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[23], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[23]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[24], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[24]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[25], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[25]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[26], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[26]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[27], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[27]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[28], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[28]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[29], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[29]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[2], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[2]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[30], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[30]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[31], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[31]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[32], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[32]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[33], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[33]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[34], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[34]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[35], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[35]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[36], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[36]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[37], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[37]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[38], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[38]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[39], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[39]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[3], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[3]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[40], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[40]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[41], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[41]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[42], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[42]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[43], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[43]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[44], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[44]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[45], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[45]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[46], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[46]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[47], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[47]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[48], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[48]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[49], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[49]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[4], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[4]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[50], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[50]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[51], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[51]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[52], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[52]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[53], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[53]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[54], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[54]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[55], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[55]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[56], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[56]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[57], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[57]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[58], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[58]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[59], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[59]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[5], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[5]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[60], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[60]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[61], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[61]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[62], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[62]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[63], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[63]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[64], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[64]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[65], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[65]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[66], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[66]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[67], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[67]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[68], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[68]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[69], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[69]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[6], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[6]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[70], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[70]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[71], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[71]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[72], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[72]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[73], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[73]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[74], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[74]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[75], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[75]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[76], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[76]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[77], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[77]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[78], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[78]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[79], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[79]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[7], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[7]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[80], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[80]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[81], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[81]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[82], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[82]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[83], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[83]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[84], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[84]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[85], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[85]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[86], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[86]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[87], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[87]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[88], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[88]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[89], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[89]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[8], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[8]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[90], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[90]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[91], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[91]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[92], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[92]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[93], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[93]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[94], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[94]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[95], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[95]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[96], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[96]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[97], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[97]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[98], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[98]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[99], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[99]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRDATA1[9], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[9]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRID0[0], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRID0_delay[0]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRID0[1], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRID0_delay[1]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRID0[2], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRID0_delay[2]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRID0[3], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRID0_delay[3]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRID1[0], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRID1_delay[0]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRID1[1], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRID1_delay[1]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRID1[2], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRID1_delay[2]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRID1[3], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRID1_delay[3]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRLAST0, 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRLAST0_delay);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRLAST1, 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRLAST1_delay);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRRESP0[1], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRRESP0_delay[1]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRRESP1[1], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRRESP1_delay[1]);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRVALID0, 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRVALID0_delay);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECRVALID1, 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRVALID1_delay);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECWREADY0, 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECWREADY0_delay);
    $setuphold (posedge PLVCUAXIDECCLK, negedge PLVCUDECWREADY1, 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECWREADY1_delay);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECARREADY0, 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECARREADY0_delay);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECARREADY1, 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECARREADY1_delay);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECAWREADY0, 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECAWREADY0_delay);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECAWREADY1, 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECAWREADY1_delay);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECBID0[0], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECBID0_delay[0]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECBID0[1], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECBID0_delay[1]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECBID0[2], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECBID0_delay[2]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECBID0[3], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECBID0_delay[3]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECBID1[0], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECBID1_delay[0]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECBID1[1], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECBID1_delay[1]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECBID1[2], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECBID1_delay[2]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECBID1[3], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECBID1_delay[3]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECBRESP0[1], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECBRESP0_delay[1]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECBRESP1[1], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECBRESP1_delay[1]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECBVALID0, 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECBVALID0_delay);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECBVALID1, 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECBVALID1_delay);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[0], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[0]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[100], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[100]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[101], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[101]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[102], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[102]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[103], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[103]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[104], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[104]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[105], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[105]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[106], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[106]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[107], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[107]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[108], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[108]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[109], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[109]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[10], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[10]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[110], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[110]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[111], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[111]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[112], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[112]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[113], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[113]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[114], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[114]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[115], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[115]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[116], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[116]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[117], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[117]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[118], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[118]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[119], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[119]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[11], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[11]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[120], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[120]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[121], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[121]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[122], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[122]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[123], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[123]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[124], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[124]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[125], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[125]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[126], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[126]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[127], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[127]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[12], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[12]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[13], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[13]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[14], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[14]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[15], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[15]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[16], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[16]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[17], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[17]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[18], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[18]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[19], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[19]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[1], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[1]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[20], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[20]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[21], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[21]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[22], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[22]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[23], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[23]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[24], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[24]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[25], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[25]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[26], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[26]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[27], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[27]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[28], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[28]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[29], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[29]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[2], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[2]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[30], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[30]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[31], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[31]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[32], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[32]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[33], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[33]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[34], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[34]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[35], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[35]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[36], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[36]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[37], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[37]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[38], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[38]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[39], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[39]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[3], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[3]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[40], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[40]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[41], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[41]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[42], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[42]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[43], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[43]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[44], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[44]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[45], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[45]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[46], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[46]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[47], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[47]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[48], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[48]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[49], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[49]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[4], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[4]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[50], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[50]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[51], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[51]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[52], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[52]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[53], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[53]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[54], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[54]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[55], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[55]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[56], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[56]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[57], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[57]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[58], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[58]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[59], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[59]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[5], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[5]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[60], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[60]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[61], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[61]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[62], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[62]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[63], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[63]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[64], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[64]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[65], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[65]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[66], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[66]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[67], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[67]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[68], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[68]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[69], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[69]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[6], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[6]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[70], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[70]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[71], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[71]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[72], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[72]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[73], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[73]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[74], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[74]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[75], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[75]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[76], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[76]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[77], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[77]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[78], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[78]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[79], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[79]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[7], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[7]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[80], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[80]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[81], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[81]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[82], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[82]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[83], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[83]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[84], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[84]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[85], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[85]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[86], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[86]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[87], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[87]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[88], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[88]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[89], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[89]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[8], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[8]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[90], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[90]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[91], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[91]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[92], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[92]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[93], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[93]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[94], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[94]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[95], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[95]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[96], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[96]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[97], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[97]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[98], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[98]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[99], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[99]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA0[9], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA0_delay[9]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[0], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[0]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[100], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[100]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[101], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[101]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[102], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[102]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[103], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[103]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[104], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[104]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[105], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[105]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[106], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[106]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[107], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[107]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[108], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[108]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[109], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[109]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[10], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[10]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[110], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[110]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[111], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[111]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[112], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[112]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[113], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[113]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[114], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[114]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[115], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[115]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[116], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[116]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[117], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[117]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[118], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[118]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[119], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[119]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[11], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[11]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[120], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[120]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[121], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[121]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[122], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[122]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[123], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[123]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[124], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[124]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[125], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[125]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[126], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[126]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[127], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[127]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[12], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[12]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[13], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[13]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[14], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[14]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[15], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[15]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[16], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[16]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[17], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[17]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[18], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[18]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[19], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[19]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[1], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[1]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[20], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[20]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[21], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[21]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[22], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[22]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[23], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[23]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[24], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[24]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[25], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[25]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[26], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[26]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[27], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[27]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[28], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[28]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[29], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[29]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[2], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[2]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[30], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[30]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[31], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[31]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[32], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[32]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[33], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[33]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[34], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[34]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[35], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[35]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[36], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[36]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[37], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[37]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[38], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[38]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[39], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[39]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[3], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[3]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[40], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[40]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[41], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[41]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[42], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[42]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[43], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[43]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[44], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[44]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[45], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[45]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[46], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[46]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[47], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[47]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[48], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[48]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[49], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[49]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[4], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[4]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[50], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[50]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[51], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[51]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[52], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[52]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[53], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[53]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[54], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[54]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[55], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[55]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[56], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[56]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[57], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[57]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[58], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[58]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[59], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[59]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[5], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[5]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[60], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[60]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[61], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[61]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[62], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[62]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[63], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[63]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[64], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[64]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[65], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[65]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[66], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[66]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[67], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[67]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[68], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[68]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[69], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[69]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[6], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[6]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[70], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[70]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[71], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[71]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[72], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[72]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[73], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[73]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[74], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[74]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[75], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[75]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[76], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[76]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[77], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[77]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[78], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[78]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[79], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[79]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[7], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[7]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[80], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[80]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[81], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[81]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[82], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[82]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[83], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[83]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[84], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[84]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[85], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[85]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[86], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[86]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[87], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[87]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[88], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[88]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[89], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[89]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[8], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[8]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[90], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[90]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[91], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[91]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[92], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[92]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[93], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[93]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[94], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[94]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[95], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[95]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[96], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[96]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[97], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[97]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[98], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[98]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[99], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[99]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRDATA1[9], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRDATA1_delay[9]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRID0[0], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRID0_delay[0]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRID0[1], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRID0_delay[1]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRID0[2], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRID0_delay[2]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRID0[3], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRID0_delay[3]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRID1[0], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRID1_delay[0]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRID1[1], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRID1_delay[1]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRID1[2], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRID1_delay[2]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRID1[3], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRID1_delay[3]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRLAST0, 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRLAST0_delay);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRLAST1, 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRLAST1_delay);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRRESP0[1], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRRESP0_delay[1]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRRESP1[1], 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRRESP1_delay[1]);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRVALID0, 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRVALID0_delay);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECRVALID1, 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECRVALID1_delay);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECWREADY0, 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECWREADY0_delay);
    $setuphold (posedge PLVCUAXIDECCLK, posedge PLVCUDECWREADY1, 0:0:0, 0:0:0, notifier, , , PLVCUAXIDECCLK_delay, PLVCUDECWREADY1_delay);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCARREADY0, 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCARREADY0_delay);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCARREADY1, 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCARREADY1_delay);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCAWREADY0, 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCAWREADY0_delay);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCAWREADY1, 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCAWREADY1_delay);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCBID0[0], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCBID0_delay[0]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCBID0[1], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCBID0_delay[1]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCBID0[2], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCBID0_delay[2]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCBID0[3], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCBID0_delay[3]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCBID1[0], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCBID1_delay[0]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCBID1[1], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCBID1_delay[1]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCBID1[2], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCBID1_delay[2]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCBID1[3], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCBID1_delay[3]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCBRESP0[1], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCBRESP0_delay[1]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCBRESP1[1], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCBRESP1_delay[1]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCBVALID0, 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCBVALID0_delay);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCBVALID1, 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCBVALID1_delay);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[0], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[0]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[100], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[100]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[101], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[101]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[102], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[102]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[103], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[103]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[104], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[104]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[105], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[105]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[106], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[106]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[107], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[107]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[108], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[108]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[109], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[109]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[10], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[10]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[110], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[110]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[111], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[111]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[112], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[112]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[113], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[113]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[114], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[114]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[115], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[115]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[116], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[116]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[117], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[117]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[118], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[118]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[119], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[119]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[11], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[11]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[120], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[120]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[121], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[121]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[122], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[122]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[123], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[123]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[124], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[124]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[125], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[125]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[126], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[126]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[127], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[127]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[12], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[12]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[13], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[13]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[14], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[14]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[15], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[15]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[16], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[16]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[17], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[17]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[18], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[18]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[19], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[19]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[1], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[1]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[20], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[20]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[21], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[21]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[22], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[22]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[23], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[23]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[24], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[24]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[25], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[25]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[26], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[26]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[27], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[27]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[28], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[28]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[29], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[29]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[2], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[2]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[30], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[30]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[31], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[31]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[32], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[32]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[33], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[33]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[34], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[34]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[35], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[35]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[36], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[36]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[37], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[37]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[38], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[38]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[39], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[39]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[3], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[3]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[40], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[40]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[41], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[41]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[42], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[42]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[43], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[43]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[44], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[44]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[45], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[45]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[46], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[46]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[47], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[47]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[48], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[48]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[49], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[49]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[4], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[4]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[50], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[50]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[51], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[51]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[52], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[52]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[53], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[53]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[54], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[54]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[55], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[55]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[56], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[56]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[57], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[57]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[58], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[58]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[59], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[59]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[5], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[5]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[60], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[60]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[61], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[61]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[62], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[62]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[63], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[63]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[64], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[64]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[65], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[65]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[66], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[66]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[67], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[67]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[68], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[68]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[69], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[69]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[6], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[6]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[70], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[70]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[71], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[71]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[72], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[72]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[73], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[73]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[74], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[74]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[75], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[75]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[76], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[76]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[77], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[77]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[78], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[78]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[79], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[79]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[7], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[7]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[80], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[80]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[81], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[81]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[82], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[82]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[83], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[83]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[84], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[84]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[85], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[85]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[86], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[86]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[87], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[87]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[88], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[88]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[89], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[89]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[8], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[8]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[90], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[90]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[91], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[91]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[92], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[92]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[93], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[93]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[94], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[94]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[95], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[95]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[96], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[96]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[97], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[97]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[98], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[98]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[99], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[99]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA0[9], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[9]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[0], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[0]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[100], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[100]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[101], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[101]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[102], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[102]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[103], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[103]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[104], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[104]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[105], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[105]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[106], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[106]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[107], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[107]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[108], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[108]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[109], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[109]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[10], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[10]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[110], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[110]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[111], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[111]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[112], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[112]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[113], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[113]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[114], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[114]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[115], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[115]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[116], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[116]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[117], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[117]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[118], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[118]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[119], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[119]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[11], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[11]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[120], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[120]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[121], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[121]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[122], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[122]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[123], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[123]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[124], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[124]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[125], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[125]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[126], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[126]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[127], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[127]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[12], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[12]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[13], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[13]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[14], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[14]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[15], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[15]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[16], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[16]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[17], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[17]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[18], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[18]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[19], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[19]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[1], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[1]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[20], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[20]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[21], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[21]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[22], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[22]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[23], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[23]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[24], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[24]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[25], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[25]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[26], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[26]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[27], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[27]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[28], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[28]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[29], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[29]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[2], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[2]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[30], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[30]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[31], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[31]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[32], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[32]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[33], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[33]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[34], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[34]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[35], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[35]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[36], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[36]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[37], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[37]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[38], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[38]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[39], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[39]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[3], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[3]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[40], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[40]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[41], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[41]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[42], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[42]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[43], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[43]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[44], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[44]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[45], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[45]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[46], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[46]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[47], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[47]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[48], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[48]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[49], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[49]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[4], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[4]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[50], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[50]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[51], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[51]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[52], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[52]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[53], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[53]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[54], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[54]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[55], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[55]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[56], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[56]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[57], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[57]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[58], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[58]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[59], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[59]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[5], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[5]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[60], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[60]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[61], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[61]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[62], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[62]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[63], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[63]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[64], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[64]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[65], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[65]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[66], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[66]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[67], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[67]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[68], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[68]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[69], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[69]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[6], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[6]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[70], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[70]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[71], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[71]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[72], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[72]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[73], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[73]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[74], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[74]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[75], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[75]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[76], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[76]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[77], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[77]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[78], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[78]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[79], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[79]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[7], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[7]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[80], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[80]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[81], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[81]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[82], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[82]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[83], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[83]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[84], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[84]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[85], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[85]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[86], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[86]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[87], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[87]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[88], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[88]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[89], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[89]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[8], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[8]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[90], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[90]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[91], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[91]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[92], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[92]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[93], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[93]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[94], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[94]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[95], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[95]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[96], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[96]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[97], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[97]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[98], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[98]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[99], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[99]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRDATA1[9], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[9]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRID0[0], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRID0_delay[0]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRID0[1], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRID0_delay[1]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRID0[2], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRID0_delay[2]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRID0[3], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRID0_delay[3]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRID1[0], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRID1_delay[0]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRID1[1], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRID1_delay[1]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRID1[2], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRID1_delay[2]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRID1[3], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRID1_delay[3]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRLAST0, 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRLAST0_delay);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRLAST1, 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRLAST1_delay);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRRESP0[1], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRRESP0_delay[1]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRRESP1[1], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRRESP1_delay[1]);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRVALID0, 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRVALID0_delay);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCRVALID1, 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRVALID1_delay);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCWREADY0, 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCWREADY0_delay);
    $setuphold (posedge PLVCUAXIENCCLK, negedge PLVCUENCWREADY1, 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCWREADY1_delay);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCARREADY0, 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCARREADY0_delay);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCARREADY1, 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCARREADY1_delay);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCAWREADY0, 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCAWREADY0_delay);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCAWREADY1, 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCAWREADY1_delay);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCBID0[0], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCBID0_delay[0]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCBID0[1], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCBID0_delay[1]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCBID0[2], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCBID0_delay[2]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCBID0[3], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCBID0_delay[3]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCBID1[0], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCBID1_delay[0]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCBID1[1], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCBID1_delay[1]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCBID1[2], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCBID1_delay[2]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCBID1[3], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCBID1_delay[3]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCBRESP0[1], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCBRESP0_delay[1]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCBRESP1[1], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCBRESP1_delay[1]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCBVALID0, 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCBVALID0_delay);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCBVALID1, 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCBVALID1_delay);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[0], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[0]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[100], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[100]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[101], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[101]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[102], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[102]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[103], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[103]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[104], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[104]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[105], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[105]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[106], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[106]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[107], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[107]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[108], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[108]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[109], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[109]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[10], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[10]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[110], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[110]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[111], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[111]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[112], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[112]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[113], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[113]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[114], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[114]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[115], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[115]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[116], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[116]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[117], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[117]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[118], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[118]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[119], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[119]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[11], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[11]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[120], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[120]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[121], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[121]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[122], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[122]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[123], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[123]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[124], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[124]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[125], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[125]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[126], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[126]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[127], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[127]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[12], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[12]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[13], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[13]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[14], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[14]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[15], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[15]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[16], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[16]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[17], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[17]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[18], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[18]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[19], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[19]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[1], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[1]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[20], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[20]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[21], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[21]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[22], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[22]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[23], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[23]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[24], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[24]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[25], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[25]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[26], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[26]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[27], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[27]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[28], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[28]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[29], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[29]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[2], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[2]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[30], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[30]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[31], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[31]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[32], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[32]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[33], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[33]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[34], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[34]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[35], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[35]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[36], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[36]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[37], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[37]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[38], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[38]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[39], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[39]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[3], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[3]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[40], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[40]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[41], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[41]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[42], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[42]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[43], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[43]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[44], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[44]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[45], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[45]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[46], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[46]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[47], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[47]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[48], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[48]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[49], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[49]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[4], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[4]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[50], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[50]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[51], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[51]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[52], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[52]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[53], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[53]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[54], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[54]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[55], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[55]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[56], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[56]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[57], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[57]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[58], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[58]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[59], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[59]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[5], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[5]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[60], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[60]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[61], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[61]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[62], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[62]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[63], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[63]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[64], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[64]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[65], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[65]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[66], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[66]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[67], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[67]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[68], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[68]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[69], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[69]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[6], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[6]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[70], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[70]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[71], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[71]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[72], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[72]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[73], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[73]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[74], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[74]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[75], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[75]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[76], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[76]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[77], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[77]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[78], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[78]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[79], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[79]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[7], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[7]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[80], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[80]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[81], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[81]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[82], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[82]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[83], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[83]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[84], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[84]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[85], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[85]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[86], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[86]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[87], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[87]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[88], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[88]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[89], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[89]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[8], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[8]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[90], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[90]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[91], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[91]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[92], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[92]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[93], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[93]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[94], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[94]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[95], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[95]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[96], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[96]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[97], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[97]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[98], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[98]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[99], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[99]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA0[9], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA0_delay[9]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[0], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[0]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[100], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[100]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[101], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[101]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[102], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[102]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[103], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[103]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[104], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[104]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[105], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[105]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[106], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[106]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[107], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[107]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[108], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[108]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[109], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[109]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[10], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[10]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[110], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[110]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[111], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[111]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[112], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[112]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[113], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[113]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[114], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[114]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[115], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[115]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[116], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[116]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[117], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[117]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[118], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[118]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[119], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[119]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[11], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[11]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[120], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[120]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[121], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[121]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[122], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[122]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[123], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[123]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[124], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[124]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[125], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[125]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[126], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[126]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[127], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[127]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[12], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[12]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[13], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[13]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[14], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[14]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[15], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[15]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[16], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[16]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[17], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[17]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[18], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[18]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[19], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[19]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[1], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[1]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[20], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[20]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[21], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[21]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[22], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[22]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[23], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[23]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[24], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[24]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[25], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[25]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[26], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[26]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[27], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[27]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[28], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[28]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[29], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[29]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[2], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[2]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[30], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[30]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[31], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[31]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[32], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[32]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[33], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[33]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[34], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[34]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[35], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[35]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[36], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[36]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[37], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[37]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[38], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[38]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[39], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[39]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[3], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[3]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[40], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[40]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[41], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[41]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[42], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[42]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[43], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[43]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[44], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[44]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[45], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[45]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[46], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[46]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[47], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[47]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[48], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[48]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[49], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[49]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[4], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[4]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[50], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[50]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[51], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[51]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[52], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[52]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[53], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[53]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[54], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[54]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[55], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[55]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[56], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[56]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[57], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[57]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[58], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[58]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[59], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[59]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[5], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[5]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[60], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[60]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[61], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[61]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[62], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[62]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[63], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[63]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[64], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[64]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[65], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[65]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[66], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[66]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[67], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[67]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[68], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[68]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[69], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[69]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[6], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[6]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[70], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[70]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[71], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[71]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[72], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[72]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[73], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[73]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[74], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[74]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[75], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[75]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[76], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[76]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[77], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[77]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[78], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[78]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[79], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[79]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[7], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[7]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[80], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[80]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[81], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[81]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[82], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[82]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[83], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[83]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[84], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[84]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[85], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[85]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[86], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[86]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[87], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[87]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[88], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[88]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[89], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[89]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[8], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[8]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[90], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[90]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[91], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[91]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[92], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[92]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[93], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[93]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[94], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[94]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[95], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[95]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[96], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[96]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[97], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[97]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[98], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[98]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[99], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[99]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRDATA1[9], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRDATA1_delay[9]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRID0[0], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRID0_delay[0]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRID0[1], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRID0_delay[1]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRID0[2], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRID0_delay[2]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRID0[3], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRID0_delay[3]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRID1[0], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRID1_delay[0]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRID1[1], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRID1_delay[1]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRID1[2], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRID1_delay[2]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRID1[3], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRID1_delay[3]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRLAST0, 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRLAST0_delay);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRLAST1, 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRLAST1_delay);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRRESP0[1], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRRESP0_delay[1]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRRESP1[1], 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRRESP1_delay[1]);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRVALID0, 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRVALID0_delay);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCRVALID1, 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCRVALID1_delay);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCWREADY0, 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCWREADY0_delay);
    $setuphold (posedge PLVCUAXIENCCLK, posedge PLVCUENCWREADY1, 0:0:0, 0:0:0, notifier, , , PLVCUAXIENCCLK_delay, PLVCUENCWREADY1_delay);
    $setuphold (posedge PLVCUAXILITECLK, negedge PLVCUARADDRAXILITEAPB[0], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUARADDRAXILITEAPB_delay[0]);
    $setuphold (posedge PLVCUAXILITECLK, negedge PLVCUARADDRAXILITEAPB[10], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUARADDRAXILITEAPB_delay[10]);
    $setuphold (posedge PLVCUAXILITECLK, negedge PLVCUARADDRAXILITEAPB[11], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUARADDRAXILITEAPB_delay[11]);
    $setuphold (posedge PLVCUAXILITECLK, negedge PLVCUARADDRAXILITEAPB[12], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUARADDRAXILITEAPB_delay[12]);
    $setuphold (posedge PLVCUAXILITECLK, negedge PLVCUARADDRAXILITEAPB[13], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUARADDRAXILITEAPB_delay[13]);
    $setuphold (posedge PLVCUAXILITECLK, negedge PLVCUARADDRAXILITEAPB[14], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUARADDRAXILITEAPB_delay[14]);
    $setuphold (posedge PLVCUAXILITECLK, negedge PLVCUARADDRAXILITEAPB[15], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUARADDRAXILITEAPB_delay[15]);
    $setuphold (posedge PLVCUAXILITECLK, negedge PLVCUARADDRAXILITEAPB[16], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUARADDRAXILITEAPB_delay[16]);
    $setuphold (posedge PLVCUAXILITECLK, negedge PLVCUARADDRAXILITEAPB[17], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUARADDRAXILITEAPB_delay[17]);
    $setuphold (posedge PLVCUAXILITECLK, negedge PLVCUARADDRAXILITEAPB[18], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUARADDRAXILITEAPB_delay[18]);
    $setuphold (posedge PLVCUAXILITECLK, negedge PLVCUARADDRAXILITEAPB[19], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUARADDRAXILITEAPB_delay[19]);
    $setuphold (posedge PLVCUAXILITECLK, negedge PLVCUARADDRAXILITEAPB[1], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUARADDRAXILITEAPB_delay[1]);
    $setuphold (posedge PLVCUAXILITECLK, negedge PLVCUARADDRAXILITEAPB[2], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUARADDRAXILITEAPB_delay[2]);
    $setuphold (posedge PLVCUAXILITECLK, negedge PLVCUARADDRAXILITEAPB[3], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUARADDRAXILITEAPB_delay[3]);
    $setuphold (posedge PLVCUAXILITECLK, negedge PLVCUARADDRAXILITEAPB[4], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUARADDRAXILITEAPB_delay[4]);
    $setuphold (posedge PLVCUAXILITECLK, negedge PLVCUARADDRAXILITEAPB[5], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUARADDRAXILITEAPB_delay[5]);
    $setuphold (posedge PLVCUAXILITECLK, negedge PLVCUARADDRAXILITEAPB[6], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUARADDRAXILITEAPB_delay[6]);
    $setuphold (posedge PLVCUAXILITECLK, negedge PLVCUARADDRAXILITEAPB[7], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUARADDRAXILITEAPB_delay[7]);
    $setuphold (posedge PLVCUAXILITECLK, negedge PLVCUARADDRAXILITEAPB[8], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUARADDRAXILITEAPB_delay[8]);
    $setuphold (posedge PLVCUAXILITECLK, negedge PLVCUARADDRAXILITEAPB[9], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUARADDRAXILITEAPB_delay[9]);
    $setuphold (posedge PLVCUAXILITECLK, negedge PLVCUARPROTAXILITEAPB[0], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUARPROTAXILITEAPB_delay[0]);
    $setuphold (posedge PLVCUAXILITECLK, negedge PLVCUARPROTAXILITEAPB[1], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUARPROTAXILITEAPB_delay[1]);
    $setuphold (posedge PLVCUAXILITECLK, negedge PLVCUARPROTAXILITEAPB[2], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUARPROTAXILITEAPB_delay[2]);
    $setuphold (posedge PLVCUAXILITECLK, negedge PLVCUARVALIDAXILITEAPB, 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUARVALIDAXILITEAPB_delay);
    $setuphold (posedge PLVCUAXILITECLK, negedge PLVCUAWADDRAXILITEAPB[0], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUAWADDRAXILITEAPB_delay[0]);
    $setuphold (posedge PLVCUAXILITECLK, negedge PLVCUAWADDRAXILITEAPB[10], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUAWADDRAXILITEAPB_delay[10]);
    $setuphold (posedge PLVCUAXILITECLK, negedge PLVCUAWADDRAXILITEAPB[11], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUAWADDRAXILITEAPB_delay[11]);
    $setuphold (posedge PLVCUAXILITECLK, negedge PLVCUAWADDRAXILITEAPB[12], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUAWADDRAXILITEAPB_delay[12]);
    $setuphold (posedge PLVCUAXILITECLK, negedge PLVCUAWADDRAXILITEAPB[13], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUAWADDRAXILITEAPB_delay[13]);
    $setuphold (posedge PLVCUAXILITECLK, negedge PLVCUAWADDRAXILITEAPB[14], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUAWADDRAXILITEAPB_delay[14]);
    $setuphold (posedge PLVCUAXILITECLK, negedge PLVCUAWADDRAXILITEAPB[15], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUAWADDRAXILITEAPB_delay[15]);
    $setuphold (posedge PLVCUAXILITECLK, negedge PLVCUAWADDRAXILITEAPB[16], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUAWADDRAXILITEAPB_delay[16]);
    $setuphold (posedge PLVCUAXILITECLK, negedge PLVCUAWADDRAXILITEAPB[17], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUAWADDRAXILITEAPB_delay[17]);
    $setuphold (posedge PLVCUAXILITECLK, negedge PLVCUAWADDRAXILITEAPB[18], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUAWADDRAXILITEAPB_delay[18]);
    $setuphold (posedge PLVCUAXILITECLK, negedge PLVCUAWADDRAXILITEAPB[19], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUAWADDRAXILITEAPB_delay[19]);
    $setuphold (posedge PLVCUAXILITECLK, negedge PLVCUAWADDRAXILITEAPB[1], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUAWADDRAXILITEAPB_delay[1]);
    $setuphold (posedge PLVCUAXILITECLK, negedge PLVCUAWADDRAXILITEAPB[2], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUAWADDRAXILITEAPB_delay[2]);
    $setuphold (posedge PLVCUAXILITECLK, negedge PLVCUAWADDRAXILITEAPB[3], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUAWADDRAXILITEAPB_delay[3]);
    $setuphold (posedge PLVCUAXILITECLK, negedge PLVCUAWADDRAXILITEAPB[4], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUAWADDRAXILITEAPB_delay[4]);
    $setuphold (posedge PLVCUAXILITECLK, negedge PLVCUAWADDRAXILITEAPB[5], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUAWADDRAXILITEAPB_delay[5]);
    $setuphold (posedge PLVCUAXILITECLK, negedge PLVCUAWADDRAXILITEAPB[6], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUAWADDRAXILITEAPB_delay[6]);
    $setuphold (posedge PLVCUAXILITECLK, negedge PLVCUAWADDRAXILITEAPB[7], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUAWADDRAXILITEAPB_delay[7]);
    $setuphold (posedge PLVCUAXILITECLK, negedge PLVCUAWADDRAXILITEAPB[8], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUAWADDRAXILITEAPB_delay[8]);
    $setuphold (posedge PLVCUAXILITECLK, negedge PLVCUAWADDRAXILITEAPB[9], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUAWADDRAXILITEAPB_delay[9]);
    $setuphold (posedge PLVCUAXILITECLK, negedge PLVCUAWPROTAXILITEAPB[0], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUAWPROTAXILITEAPB_delay[0]);
    $setuphold (posedge PLVCUAXILITECLK, negedge PLVCUAWPROTAXILITEAPB[1], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUAWPROTAXILITEAPB_delay[1]);
    $setuphold (posedge PLVCUAXILITECLK, negedge PLVCUAWPROTAXILITEAPB[2], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUAWPROTAXILITEAPB_delay[2]);
    $setuphold (posedge PLVCUAXILITECLK, negedge PLVCUAWVALIDAXILITEAPB, 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUAWVALIDAXILITEAPB_delay);
    $setuphold (posedge PLVCUAXILITECLK, negedge PLVCUBREADYAXILITEAPB, 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUBREADYAXILITEAPB_delay);
    $setuphold (posedge PLVCUAXILITECLK, negedge PLVCURREADYAXILITEAPB, 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCURREADYAXILITEAPB_delay);
    $setuphold (posedge PLVCUAXILITECLK, negedge PLVCUWDATAAXILITEAPB[0], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUWDATAAXILITEAPB_delay[0]);
    $setuphold (posedge PLVCUAXILITECLK, negedge PLVCUWDATAAXILITEAPB[10], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUWDATAAXILITEAPB_delay[10]);
    $setuphold (posedge PLVCUAXILITECLK, negedge PLVCUWDATAAXILITEAPB[11], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUWDATAAXILITEAPB_delay[11]);
    $setuphold (posedge PLVCUAXILITECLK, negedge PLVCUWDATAAXILITEAPB[12], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUWDATAAXILITEAPB_delay[12]);
    $setuphold (posedge PLVCUAXILITECLK, negedge PLVCUWDATAAXILITEAPB[13], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUWDATAAXILITEAPB_delay[13]);
    $setuphold (posedge PLVCUAXILITECLK, negedge PLVCUWDATAAXILITEAPB[14], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUWDATAAXILITEAPB_delay[14]);
    $setuphold (posedge PLVCUAXILITECLK, negedge PLVCUWDATAAXILITEAPB[15], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUWDATAAXILITEAPB_delay[15]);
    $setuphold (posedge PLVCUAXILITECLK, negedge PLVCUWDATAAXILITEAPB[16], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUWDATAAXILITEAPB_delay[16]);
    $setuphold (posedge PLVCUAXILITECLK, negedge PLVCUWDATAAXILITEAPB[17], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUWDATAAXILITEAPB_delay[17]);
    $setuphold (posedge PLVCUAXILITECLK, negedge PLVCUWDATAAXILITEAPB[18], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUWDATAAXILITEAPB_delay[18]);
    $setuphold (posedge PLVCUAXILITECLK, negedge PLVCUWDATAAXILITEAPB[19], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUWDATAAXILITEAPB_delay[19]);
    $setuphold (posedge PLVCUAXILITECLK, negedge PLVCUWDATAAXILITEAPB[1], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUWDATAAXILITEAPB_delay[1]);
    $setuphold (posedge PLVCUAXILITECLK, negedge PLVCUWDATAAXILITEAPB[20], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUWDATAAXILITEAPB_delay[20]);
    $setuphold (posedge PLVCUAXILITECLK, negedge PLVCUWDATAAXILITEAPB[21], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUWDATAAXILITEAPB_delay[21]);
    $setuphold (posedge PLVCUAXILITECLK, negedge PLVCUWDATAAXILITEAPB[22], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUWDATAAXILITEAPB_delay[22]);
    $setuphold (posedge PLVCUAXILITECLK, negedge PLVCUWDATAAXILITEAPB[23], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUWDATAAXILITEAPB_delay[23]);
    $setuphold (posedge PLVCUAXILITECLK, negedge PLVCUWDATAAXILITEAPB[24], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUWDATAAXILITEAPB_delay[24]);
    $setuphold (posedge PLVCUAXILITECLK, negedge PLVCUWDATAAXILITEAPB[25], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUWDATAAXILITEAPB_delay[25]);
    $setuphold (posedge PLVCUAXILITECLK, negedge PLVCUWDATAAXILITEAPB[26], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUWDATAAXILITEAPB_delay[26]);
    $setuphold (posedge PLVCUAXILITECLK, negedge PLVCUWDATAAXILITEAPB[27], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUWDATAAXILITEAPB_delay[27]);
    $setuphold (posedge PLVCUAXILITECLK, negedge PLVCUWDATAAXILITEAPB[28], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUWDATAAXILITEAPB_delay[28]);
    $setuphold (posedge PLVCUAXILITECLK, negedge PLVCUWDATAAXILITEAPB[29], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUWDATAAXILITEAPB_delay[29]);
    $setuphold (posedge PLVCUAXILITECLK, negedge PLVCUWDATAAXILITEAPB[2], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUWDATAAXILITEAPB_delay[2]);
    $setuphold (posedge PLVCUAXILITECLK, negedge PLVCUWDATAAXILITEAPB[30], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUWDATAAXILITEAPB_delay[30]);
    $setuphold (posedge PLVCUAXILITECLK, negedge PLVCUWDATAAXILITEAPB[31], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUWDATAAXILITEAPB_delay[31]);
    $setuphold (posedge PLVCUAXILITECLK, negedge PLVCUWDATAAXILITEAPB[3], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUWDATAAXILITEAPB_delay[3]);
    $setuphold (posedge PLVCUAXILITECLK, negedge PLVCUWDATAAXILITEAPB[4], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUWDATAAXILITEAPB_delay[4]);
    $setuphold (posedge PLVCUAXILITECLK, negedge PLVCUWDATAAXILITEAPB[5], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUWDATAAXILITEAPB_delay[5]);
    $setuphold (posedge PLVCUAXILITECLK, negedge PLVCUWDATAAXILITEAPB[6], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUWDATAAXILITEAPB_delay[6]);
    $setuphold (posedge PLVCUAXILITECLK, negedge PLVCUWDATAAXILITEAPB[7], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUWDATAAXILITEAPB_delay[7]);
    $setuphold (posedge PLVCUAXILITECLK, negedge PLVCUWDATAAXILITEAPB[8], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUWDATAAXILITEAPB_delay[8]);
    $setuphold (posedge PLVCUAXILITECLK, negedge PLVCUWDATAAXILITEAPB[9], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUWDATAAXILITEAPB_delay[9]);
    $setuphold (posedge PLVCUAXILITECLK, negedge PLVCUWSTRBAXILITEAPB[0], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUWSTRBAXILITEAPB_delay[0]);
    $setuphold (posedge PLVCUAXILITECLK, negedge PLVCUWSTRBAXILITEAPB[1], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUWSTRBAXILITEAPB_delay[1]);
    $setuphold (posedge PLVCUAXILITECLK, negedge PLVCUWSTRBAXILITEAPB[2], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUWSTRBAXILITEAPB_delay[2]);
    $setuphold (posedge PLVCUAXILITECLK, negedge PLVCUWSTRBAXILITEAPB[3], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUWSTRBAXILITEAPB_delay[3]);
    $setuphold (posedge PLVCUAXILITECLK, negedge PLVCUWVALIDAXILITEAPB, 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUWVALIDAXILITEAPB_delay);
    $setuphold (posedge PLVCUAXILITECLK, posedge PLVCUARADDRAXILITEAPB[0], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUARADDRAXILITEAPB_delay[0]);
    $setuphold (posedge PLVCUAXILITECLK, posedge PLVCUARADDRAXILITEAPB[10], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUARADDRAXILITEAPB_delay[10]);
    $setuphold (posedge PLVCUAXILITECLK, posedge PLVCUARADDRAXILITEAPB[11], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUARADDRAXILITEAPB_delay[11]);
    $setuphold (posedge PLVCUAXILITECLK, posedge PLVCUARADDRAXILITEAPB[12], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUARADDRAXILITEAPB_delay[12]);
    $setuphold (posedge PLVCUAXILITECLK, posedge PLVCUARADDRAXILITEAPB[13], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUARADDRAXILITEAPB_delay[13]);
    $setuphold (posedge PLVCUAXILITECLK, posedge PLVCUARADDRAXILITEAPB[14], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUARADDRAXILITEAPB_delay[14]);
    $setuphold (posedge PLVCUAXILITECLK, posedge PLVCUARADDRAXILITEAPB[15], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUARADDRAXILITEAPB_delay[15]);
    $setuphold (posedge PLVCUAXILITECLK, posedge PLVCUARADDRAXILITEAPB[16], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUARADDRAXILITEAPB_delay[16]);
    $setuphold (posedge PLVCUAXILITECLK, posedge PLVCUARADDRAXILITEAPB[17], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUARADDRAXILITEAPB_delay[17]);
    $setuphold (posedge PLVCUAXILITECLK, posedge PLVCUARADDRAXILITEAPB[18], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUARADDRAXILITEAPB_delay[18]);
    $setuphold (posedge PLVCUAXILITECLK, posedge PLVCUARADDRAXILITEAPB[19], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUARADDRAXILITEAPB_delay[19]);
    $setuphold (posedge PLVCUAXILITECLK, posedge PLVCUARADDRAXILITEAPB[1], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUARADDRAXILITEAPB_delay[1]);
    $setuphold (posedge PLVCUAXILITECLK, posedge PLVCUARADDRAXILITEAPB[2], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUARADDRAXILITEAPB_delay[2]);
    $setuphold (posedge PLVCUAXILITECLK, posedge PLVCUARADDRAXILITEAPB[3], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUARADDRAXILITEAPB_delay[3]);
    $setuphold (posedge PLVCUAXILITECLK, posedge PLVCUARADDRAXILITEAPB[4], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUARADDRAXILITEAPB_delay[4]);
    $setuphold (posedge PLVCUAXILITECLK, posedge PLVCUARADDRAXILITEAPB[5], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUARADDRAXILITEAPB_delay[5]);
    $setuphold (posedge PLVCUAXILITECLK, posedge PLVCUARADDRAXILITEAPB[6], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUARADDRAXILITEAPB_delay[6]);
    $setuphold (posedge PLVCUAXILITECLK, posedge PLVCUARADDRAXILITEAPB[7], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUARADDRAXILITEAPB_delay[7]);
    $setuphold (posedge PLVCUAXILITECLK, posedge PLVCUARADDRAXILITEAPB[8], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUARADDRAXILITEAPB_delay[8]);
    $setuphold (posedge PLVCUAXILITECLK, posedge PLVCUARADDRAXILITEAPB[9], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUARADDRAXILITEAPB_delay[9]);
    $setuphold (posedge PLVCUAXILITECLK, posedge PLVCUARPROTAXILITEAPB[0], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUARPROTAXILITEAPB_delay[0]);
    $setuphold (posedge PLVCUAXILITECLK, posedge PLVCUARPROTAXILITEAPB[1], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUARPROTAXILITEAPB_delay[1]);
    $setuphold (posedge PLVCUAXILITECLK, posedge PLVCUARPROTAXILITEAPB[2], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUARPROTAXILITEAPB_delay[2]);
    $setuphold (posedge PLVCUAXILITECLK, posedge PLVCUARVALIDAXILITEAPB, 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUARVALIDAXILITEAPB_delay);
    $setuphold (posedge PLVCUAXILITECLK, posedge PLVCUAWADDRAXILITEAPB[0], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUAWADDRAXILITEAPB_delay[0]);
    $setuphold (posedge PLVCUAXILITECLK, posedge PLVCUAWADDRAXILITEAPB[10], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUAWADDRAXILITEAPB_delay[10]);
    $setuphold (posedge PLVCUAXILITECLK, posedge PLVCUAWADDRAXILITEAPB[11], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUAWADDRAXILITEAPB_delay[11]);
    $setuphold (posedge PLVCUAXILITECLK, posedge PLVCUAWADDRAXILITEAPB[12], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUAWADDRAXILITEAPB_delay[12]);
    $setuphold (posedge PLVCUAXILITECLK, posedge PLVCUAWADDRAXILITEAPB[13], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUAWADDRAXILITEAPB_delay[13]);
    $setuphold (posedge PLVCUAXILITECLK, posedge PLVCUAWADDRAXILITEAPB[14], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUAWADDRAXILITEAPB_delay[14]);
    $setuphold (posedge PLVCUAXILITECLK, posedge PLVCUAWADDRAXILITEAPB[15], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUAWADDRAXILITEAPB_delay[15]);
    $setuphold (posedge PLVCUAXILITECLK, posedge PLVCUAWADDRAXILITEAPB[16], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUAWADDRAXILITEAPB_delay[16]);
    $setuphold (posedge PLVCUAXILITECLK, posedge PLVCUAWADDRAXILITEAPB[17], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUAWADDRAXILITEAPB_delay[17]);
    $setuphold (posedge PLVCUAXILITECLK, posedge PLVCUAWADDRAXILITEAPB[18], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUAWADDRAXILITEAPB_delay[18]);
    $setuphold (posedge PLVCUAXILITECLK, posedge PLVCUAWADDRAXILITEAPB[19], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUAWADDRAXILITEAPB_delay[19]);
    $setuphold (posedge PLVCUAXILITECLK, posedge PLVCUAWADDRAXILITEAPB[1], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUAWADDRAXILITEAPB_delay[1]);
    $setuphold (posedge PLVCUAXILITECLK, posedge PLVCUAWADDRAXILITEAPB[2], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUAWADDRAXILITEAPB_delay[2]);
    $setuphold (posedge PLVCUAXILITECLK, posedge PLVCUAWADDRAXILITEAPB[3], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUAWADDRAXILITEAPB_delay[3]);
    $setuphold (posedge PLVCUAXILITECLK, posedge PLVCUAWADDRAXILITEAPB[4], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUAWADDRAXILITEAPB_delay[4]);
    $setuphold (posedge PLVCUAXILITECLK, posedge PLVCUAWADDRAXILITEAPB[5], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUAWADDRAXILITEAPB_delay[5]);
    $setuphold (posedge PLVCUAXILITECLK, posedge PLVCUAWADDRAXILITEAPB[6], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUAWADDRAXILITEAPB_delay[6]);
    $setuphold (posedge PLVCUAXILITECLK, posedge PLVCUAWADDRAXILITEAPB[7], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUAWADDRAXILITEAPB_delay[7]);
    $setuphold (posedge PLVCUAXILITECLK, posedge PLVCUAWADDRAXILITEAPB[8], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUAWADDRAXILITEAPB_delay[8]);
    $setuphold (posedge PLVCUAXILITECLK, posedge PLVCUAWADDRAXILITEAPB[9], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUAWADDRAXILITEAPB_delay[9]);
    $setuphold (posedge PLVCUAXILITECLK, posedge PLVCUAWPROTAXILITEAPB[0], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUAWPROTAXILITEAPB_delay[0]);
    $setuphold (posedge PLVCUAXILITECLK, posedge PLVCUAWPROTAXILITEAPB[1], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUAWPROTAXILITEAPB_delay[1]);
    $setuphold (posedge PLVCUAXILITECLK, posedge PLVCUAWPROTAXILITEAPB[2], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUAWPROTAXILITEAPB_delay[2]);
    $setuphold (posedge PLVCUAXILITECLK, posedge PLVCUAWVALIDAXILITEAPB, 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUAWVALIDAXILITEAPB_delay);
    $setuphold (posedge PLVCUAXILITECLK, posedge PLVCUBREADYAXILITEAPB, 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUBREADYAXILITEAPB_delay);
    $setuphold (posedge PLVCUAXILITECLK, posedge PLVCURREADYAXILITEAPB, 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCURREADYAXILITEAPB_delay);
    $setuphold (posedge PLVCUAXILITECLK, posedge PLVCUWDATAAXILITEAPB[0], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUWDATAAXILITEAPB_delay[0]);
    $setuphold (posedge PLVCUAXILITECLK, posedge PLVCUWDATAAXILITEAPB[10], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUWDATAAXILITEAPB_delay[10]);
    $setuphold (posedge PLVCUAXILITECLK, posedge PLVCUWDATAAXILITEAPB[11], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUWDATAAXILITEAPB_delay[11]);
    $setuphold (posedge PLVCUAXILITECLK, posedge PLVCUWDATAAXILITEAPB[12], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUWDATAAXILITEAPB_delay[12]);
    $setuphold (posedge PLVCUAXILITECLK, posedge PLVCUWDATAAXILITEAPB[13], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUWDATAAXILITEAPB_delay[13]);
    $setuphold (posedge PLVCUAXILITECLK, posedge PLVCUWDATAAXILITEAPB[14], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUWDATAAXILITEAPB_delay[14]);
    $setuphold (posedge PLVCUAXILITECLK, posedge PLVCUWDATAAXILITEAPB[15], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUWDATAAXILITEAPB_delay[15]);
    $setuphold (posedge PLVCUAXILITECLK, posedge PLVCUWDATAAXILITEAPB[16], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUWDATAAXILITEAPB_delay[16]);
    $setuphold (posedge PLVCUAXILITECLK, posedge PLVCUWDATAAXILITEAPB[17], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUWDATAAXILITEAPB_delay[17]);
    $setuphold (posedge PLVCUAXILITECLK, posedge PLVCUWDATAAXILITEAPB[18], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUWDATAAXILITEAPB_delay[18]);
    $setuphold (posedge PLVCUAXILITECLK, posedge PLVCUWDATAAXILITEAPB[19], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUWDATAAXILITEAPB_delay[19]);
    $setuphold (posedge PLVCUAXILITECLK, posedge PLVCUWDATAAXILITEAPB[1], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUWDATAAXILITEAPB_delay[1]);
    $setuphold (posedge PLVCUAXILITECLK, posedge PLVCUWDATAAXILITEAPB[20], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUWDATAAXILITEAPB_delay[20]);
    $setuphold (posedge PLVCUAXILITECLK, posedge PLVCUWDATAAXILITEAPB[21], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUWDATAAXILITEAPB_delay[21]);
    $setuphold (posedge PLVCUAXILITECLK, posedge PLVCUWDATAAXILITEAPB[22], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUWDATAAXILITEAPB_delay[22]);
    $setuphold (posedge PLVCUAXILITECLK, posedge PLVCUWDATAAXILITEAPB[23], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUWDATAAXILITEAPB_delay[23]);
    $setuphold (posedge PLVCUAXILITECLK, posedge PLVCUWDATAAXILITEAPB[24], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUWDATAAXILITEAPB_delay[24]);
    $setuphold (posedge PLVCUAXILITECLK, posedge PLVCUWDATAAXILITEAPB[25], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUWDATAAXILITEAPB_delay[25]);
    $setuphold (posedge PLVCUAXILITECLK, posedge PLVCUWDATAAXILITEAPB[26], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUWDATAAXILITEAPB_delay[26]);
    $setuphold (posedge PLVCUAXILITECLK, posedge PLVCUWDATAAXILITEAPB[27], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUWDATAAXILITEAPB_delay[27]);
    $setuphold (posedge PLVCUAXILITECLK, posedge PLVCUWDATAAXILITEAPB[28], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUWDATAAXILITEAPB_delay[28]);
    $setuphold (posedge PLVCUAXILITECLK, posedge PLVCUWDATAAXILITEAPB[29], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUWDATAAXILITEAPB_delay[29]);
    $setuphold (posedge PLVCUAXILITECLK, posedge PLVCUWDATAAXILITEAPB[2], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUWDATAAXILITEAPB_delay[2]);
    $setuphold (posedge PLVCUAXILITECLK, posedge PLVCUWDATAAXILITEAPB[30], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUWDATAAXILITEAPB_delay[30]);
    $setuphold (posedge PLVCUAXILITECLK, posedge PLVCUWDATAAXILITEAPB[31], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUWDATAAXILITEAPB_delay[31]);
    $setuphold (posedge PLVCUAXILITECLK, posedge PLVCUWDATAAXILITEAPB[3], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUWDATAAXILITEAPB_delay[3]);
    $setuphold (posedge PLVCUAXILITECLK, posedge PLVCUWDATAAXILITEAPB[4], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUWDATAAXILITEAPB_delay[4]);
    $setuphold (posedge PLVCUAXILITECLK, posedge PLVCUWDATAAXILITEAPB[5], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUWDATAAXILITEAPB_delay[5]);
    $setuphold (posedge PLVCUAXILITECLK, posedge PLVCUWDATAAXILITEAPB[6], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUWDATAAXILITEAPB_delay[6]);
    $setuphold (posedge PLVCUAXILITECLK, posedge PLVCUWDATAAXILITEAPB[7], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUWDATAAXILITEAPB_delay[7]);
    $setuphold (posedge PLVCUAXILITECLK, posedge PLVCUWDATAAXILITEAPB[8], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUWDATAAXILITEAPB_delay[8]);
    $setuphold (posedge PLVCUAXILITECLK, posedge PLVCUWDATAAXILITEAPB[9], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUWDATAAXILITEAPB_delay[9]);
    $setuphold (posedge PLVCUAXILITECLK, posedge PLVCUWSTRBAXILITEAPB[0], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUWSTRBAXILITEAPB_delay[0]);
    $setuphold (posedge PLVCUAXILITECLK, posedge PLVCUWSTRBAXILITEAPB[1], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUWSTRBAXILITEAPB_delay[1]);
    $setuphold (posedge PLVCUAXILITECLK, posedge PLVCUWSTRBAXILITEAPB[2], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUWSTRBAXILITEAPB_delay[2]);
    $setuphold (posedge PLVCUAXILITECLK, posedge PLVCUWSTRBAXILITEAPB[3], 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUWSTRBAXILITEAPB_delay[3]);
    $setuphold (posedge PLVCUAXILITECLK, posedge PLVCUWVALIDAXILITEAPB, 0:0:0, 0:0:0, notifier, , , PLVCUAXILITECLK_delay, PLVCUWVALIDAXILITEAPB_delay);
    $setuphold (posedge PLVCUAXIMCUCLK, negedge PLVCUMCUMAXIICDCARREADY, 0:0:0, 0:0:0, notifier, , , PLVCUAXIMCUCLK_delay, PLVCUMCUMAXIICDCARREADY_delay);
    $setuphold (posedge PLVCUAXIMCUCLK, negedge PLVCUMCUMAXIICDCAWREADY, 0:0:0, 0:0:0, notifier, , , PLVCUAXIMCUCLK_delay, PLVCUMCUMAXIICDCAWREADY_delay);
    $setuphold (posedge PLVCUAXIMCUCLK, negedge PLVCUMCUMAXIICDCBID[0], 0:0:0, 0:0:0, notifier, , , PLVCUAXIMCUCLK_delay, PLVCUMCUMAXIICDCBID_delay[0]);
    $setuphold (posedge PLVCUAXIMCUCLK, negedge PLVCUMCUMAXIICDCBID[1], 0:0:0, 0:0:0, notifier, , , PLVCUAXIMCUCLK_delay, PLVCUMCUMAXIICDCBID_delay[1]);
    $setuphold (posedge PLVCUAXIMCUCLK, negedge PLVCUMCUMAXIICDCBID[2], 0:0:0, 0:0:0, notifier, , , PLVCUAXIMCUCLK_delay, PLVCUMCUMAXIICDCBID_delay[2]);
    $setuphold (posedge PLVCUAXIMCUCLK, negedge PLVCUMCUMAXIICDCBRESP[0], 0:0:0, 0:0:0, notifier, , , PLVCUAXIMCUCLK_delay, PLVCUMCUMAXIICDCBRESP_delay[0]);
    $setuphold (posedge PLVCUAXIMCUCLK, negedge PLVCUMCUMAXIICDCBRESP[1], 0:0:0, 0:0:0, notifier, , , PLVCUAXIMCUCLK_delay, PLVCUMCUMAXIICDCBRESP_delay[1]);
    $setuphold (posedge PLVCUAXIMCUCLK, negedge PLVCUMCUMAXIICDCBVALID, 0:0:0, 0:0:0, notifier, , , PLVCUAXIMCUCLK_delay, PLVCUMCUMAXIICDCBVALID_delay);
    $setuphold (posedge PLVCUAXIMCUCLK, negedge PLVCUMCUMAXIICDCRDATA[0], 0:0:0, 0:0:0, notifier, , , PLVCUAXIMCUCLK_delay, PLVCUMCUMAXIICDCRDATA_delay[0]);
    $setuphold (posedge PLVCUAXIMCUCLK, negedge PLVCUMCUMAXIICDCRDATA[10], 0:0:0, 0:0:0, notifier, , , PLVCUAXIMCUCLK_delay, PLVCUMCUMAXIICDCRDATA_delay[10]);
    $setuphold (posedge PLVCUAXIMCUCLK, negedge PLVCUMCUMAXIICDCRDATA[11], 0:0:0, 0:0:0, notifier, , , PLVCUAXIMCUCLK_delay, PLVCUMCUMAXIICDCRDATA_delay[11]);
    $setuphold (posedge PLVCUAXIMCUCLK, negedge PLVCUMCUMAXIICDCRDATA[12], 0:0:0, 0:0:0, notifier, , , PLVCUAXIMCUCLK_delay, PLVCUMCUMAXIICDCRDATA_delay[12]);
    $setuphold (posedge PLVCUAXIMCUCLK, negedge PLVCUMCUMAXIICDCRDATA[13], 0:0:0, 0:0:0, notifier, , , PLVCUAXIMCUCLK_delay, PLVCUMCUMAXIICDCRDATA_delay[13]);
    $setuphold (posedge PLVCUAXIMCUCLK, negedge PLVCUMCUMAXIICDCRDATA[14], 0:0:0, 0:0:0, notifier, , , PLVCUAXIMCUCLK_delay, PLVCUMCUMAXIICDCRDATA_delay[14]);
    $setuphold (posedge PLVCUAXIMCUCLK, negedge PLVCUMCUMAXIICDCRDATA[15], 0:0:0, 0:0:0, notifier, , , PLVCUAXIMCUCLK_delay, PLVCUMCUMAXIICDCRDATA_delay[15]);
    $setuphold (posedge PLVCUAXIMCUCLK, negedge PLVCUMCUMAXIICDCRDATA[16], 0:0:0, 0:0:0, notifier, , , PLVCUAXIMCUCLK_delay, PLVCUMCUMAXIICDCRDATA_delay[16]);
    $setuphold (posedge PLVCUAXIMCUCLK, negedge PLVCUMCUMAXIICDCRDATA[17], 0:0:0, 0:0:0, notifier, , , PLVCUAXIMCUCLK_delay, PLVCUMCUMAXIICDCRDATA_delay[17]);
    $setuphold (posedge PLVCUAXIMCUCLK, negedge PLVCUMCUMAXIICDCRDATA[18], 0:0:0, 0:0:0, notifier, , , PLVCUAXIMCUCLK_delay, PLVCUMCUMAXIICDCRDATA_delay[18]);
    $setuphold (posedge PLVCUAXIMCUCLK, negedge PLVCUMCUMAXIICDCRDATA[19], 0:0:0, 0:0:0, notifier, , , PLVCUAXIMCUCLK_delay, PLVCUMCUMAXIICDCRDATA_delay[19]);
    $setuphold (posedge PLVCUAXIMCUCLK, negedge PLVCUMCUMAXIICDCRDATA[1], 0:0:0, 0:0:0, notifier, , , PLVCUAXIMCUCLK_delay, PLVCUMCUMAXIICDCRDATA_delay[1]);
    $setuphold (posedge PLVCUAXIMCUCLK, negedge PLVCUMCUMAXIICDCRDATA[20], 0:0:0, 0:0:0, notifier, , , PLVCUAXIMCUCLK_delay, PLVCUMCUMAXIICDCRDATA_delay[20]);
    $setuphold (posedge PLVCUAXIMCUCLK, negedge PLVCUMCUMAXIICDCRDATA[21], 0:0:0, 0:0:0, notifier, , , PLVCUAXIMCUCLK_delay, PLVCUMCUMAXIICDCRDATA_delay[21]);
    $setuphold (posedge PLVCUAXIMCUCLK, negedge PLVCUMCUMAXIICDCRDATA[22], 0:0:0, 0:0:0, notifier, , , PLVCUAXIMCUCLK_delay, PLVCUMCUMAXIICDCRDATA_delay[22]);
    $setuphold (posedge PLVCUAXIMCUCLK, negedge PLVCUMCUMAXIICDCRDATA[23], 0:0:0, 0:0:0, notifier, , , PLVCUAXIMCUCLK_delay, PLVCUMCUMAXIICDCRDATA_delay[23]);
    $setuphold (posedge PLVCUAXIMCUCLK, negedge PLVCUMCUMAXIICDCRDATA[24], 0:0:0, 0:0:0, notifier, , , PLVCUAXIMCUCLK_delay, PLVCUMCUMAXIICDCRDATA_delay[24]);
    $setuphold (posedge PLVCUAXIMCUCLK, negedge PLVCUMCUMAXIICDCRDATA[25], 0:0:0, 0:0:0, notifier, , , PLVCUAXIMCUCLK_delay, PLVCUMCUMAXIICDCRDATA_delay[25]);
    $setuphold (posedge PLVCUAXIMCUCLK, negedge PLVCUMCUMAXIICDCRDATA[26], 0:0:0, 0:0:0, notifier, , , PLVCUAXIMCUCLK_delay, PLVCUMCUMAXIICDCRDATA_delay[26]);
    $setuphold (posedge PLVCUAXIMCUCLK, negedge PLVCUMCUMAXIICDCRDATA[27], 0:0:0, 0:0:0, notifier, , , PLVCUAXIMCUCLK_delay, PLVCUMCUMAXIICDCRDATA_delay[27]);
    $setuphold (posedge PLVCUAXIMCUCLK, negedge PLVCUMCUMAXIICDCRDATA[28], 0:0:0, 0:0:0, notifier, , , PLVCUAXIMCUCLK_delay, PLVCUMCUMAXIICDCRDATA_delay[28]);
    $setuphold (posedge PLVCUAXIMCUCLK, negedge PLVCUMCUMAXIICDCRDATA[29], 0:0:0, 0:0:0, notifier, , , PLVCUAXIMCUCLK_delay, PLVCUMCUMAXIICDCRDATA_delay[29]);
    $setuphold (posedge PLVCUAXIMCUCLK, negedge PLVCUMCUMAXIICDCRDATA[2], 0:0:0, 0:0:0, notifier, , , PLVCUAXIMCUCLK_delay, PLVCUMCUMAXIICDCRDATA_delay[2]);
    $setuphold (posedge PLVCUAXIMCUCLK, negedge PLVCUMCUMAXIICDCRDATA[30], 0:0:0, 0:0:0, notifier, , , PLVCUAXIMCUCLK_delay, PLVCUMCUMAXIICDCRDATA_delay[30]);
    $setuphold (posedge PLVCUAXIMCUCLK, negedge PLVCUMCUMAXIICDCRDATA[31], 0:0:0, 0:0:0, notifier, , , PLVCUAXIMCUCLK_delay, PLVCUMCUMAXIICDCRDATA_delay[31]);
    $setuphold (posedge PLVCUAXIMCUCLK, negedge PLVCUMCUMAXIICDCRDATA[3], 0:0:0, 0:0:0, notifier, , , PLVCUAXIMCUCLK_delay, PLVCUMCUMAXIICDCRDATA_delay[3]);
    $setuphold (posedge PLVCUAXIMCUCLK, negedge PLVCUMCUMAXIICDCRDATA[4], 0:0:0, 0:0:0, notifier, , , PLVCUAXIMCUCLK_delay, PLVCUMCUMAXIICDCRDATA_delay[4]);
    $setuphold (posedge PLVCUAXIMCUCLK, negedge PLVCUMCUMAXIICDCRDATA[5], 0:0:0, 0:0:0, notifier, , , PLVCUAXIMCUCLK_delay, PLVCUMCUMAXIICDCRDATA_delay[5]);
    $setuphold (posedge PLVCUAXIMCUCLK, negedge PLVCUMCUMAXIICDCRDATA[6], 0:0:0, 0:0:0, notifier, , , PLVCUAXIMCUCLK_delay, PLVCUMCUMAXIICDCRDATA_delay[6]);
    $setuphold (posedge PLVCUAXIMCUCLK, negedge PLVCUMCUMAXIICDCRDATA[7], 0:0:0, 0:0:0, notifier, , , PLVCUAXIMCUCLK_delay, PLVCUMCUMAXIICDCRDATA_delay[7]);
    $setuphold (posedge PLVCUAXIMCUCLK, negedge PLVCUMCUMAXIICDCRDATA[8], 0:0:0, 0:0:0, notifier, , , PLVCUAXIMCUCLK_delay, PLVCUMCUMAXIICDCRDATA_delay[8]);
    $setuphold (posedge PLVCUAXIMCUCLK, negedge PLVCUMCUMAXIICDCRDATA[9], 0:0:0, 0:0:0, notifier, , , PLVCUAXIMCUCLK_delay, PLVCUMCUMAXIICDCRDATA_delay[9]);
    $setuphold (posedge PLVCUAXIMCUCLK, negedge PLVCUMCUMAXIICDCRID[0], 0:0:0, 0:0:0, notifier, , , PLVCUAXIMCUCLK_delay, PLVCUMCUMAXIICDCRID_delay[0]);
    $setuphold (posedge PLVCUAXIMCUCLK, negedge PLVCUMCUMAXIICDCRID[1], 0:0:0, 0:0:0, notifier, , , PLVCUAXIMCUCLK_delay, PLVCUMCUMAXIICDCRID_delay[1]);
    $setuphold (posedge PLVCUAXIMCUCLK, negedge PLVCUMCUMAXIICDCRID[2], 0:0:0, 0:0:0, notifier, , , PLVCUAXIMCUCLK_delay, PLVCUMCUMAXIICDCRID_delay[2]);
    $setuphold (posedge PLVCUAXIMCUCLK, negedge PLVCUMCUMAXIICDCRLAST, 0:0:0, 0:0:0, notifier, , , PLVCUAXIMCUCLK_delay, PLVCUMCUMAXIICDCRLAST_delay);
    $setuphold (posedge PLVCUAXIMCUCLK, negedge PLVCUMCUMAXIICDCRRESP[0], 0:0:0, 0:0:0, notifier, , , PLVCUAXIMCUCLK_delay, PLVCUMCUMAXIICDCRRESP_delay[0]);
    $setuphold (posedge PLVCUAXIMCUCLK, negedge PLVCUMCUMAXIICDCRRESP[1], 0:0:0, 0:0:0, notifier, , , PLVCUAXIMCUCLK_delay, PLVCUMCUMAXIICDCRRESP_delay[1]);
    $setuphold (posedge PLVCUAXIMCUCLK, negedge PLVCUMCUMAXIICDCRVALID, 0:0:0, 0:0:0, notifier, , , PLVCUAXIMCUCLK_delay, PLVCUMCUMAXIICDCRVALID_delay);
    $setuphold (posedge PLVCUAXIMCUCLK, negedge PLVCUMCUMAXIICDCWREADY, 0:0:0, 0:0:0, notifier, , , PLVCUAXIMCUCLK_delay, PLVCUMCUMAXIICDCWREADY_delay);
    $setuphold (posedge PLVCUAXIMCUCLK, posedge PLVCUMCUMAXIICDCARREADY, 0:0:0, 0:0:0, notifier, , , PLVCUAXIMCUCLK_delay, PLVCUMCUMAXIICDCARREADY_delay);
    $setuphold (posedge PLVCUAXIMCUCLK, posedge PLVCUMCUMAXIICDCAWREADY, 0:0:0, 0:0:0, notifier, , , PLVCUAXIMCUCLK_delay, PLVCUMCUMAXIICDCAWREADY_delay);
    $setuphold (posedge PLVCUAXIMCUCLK, posedge PLVCUMCUMAXIICDCBID[0], 0:0:0, 0:0:0, notifier, , , PLVCUAXIMCUCLK_delay, PLVCUMCUMAXIICDCBID_delay[0]);
    $setuphold (posedge PLVCUAXIMCUCLK, posedge PLVCUMCUMAXIICDCBID[1], 0:0:0, 0:0:0, notifier, , , PLVCUAXIMCUCLK_delay, PLVCUMCUMAXIICDCBID_delay[1]);
    $setuphold (posedge PLVCUAXIMCUCLK, posedge PLVCUMCUMAXIICDCBID[2], 0:0:0, 0:0:0, notifier, , , PLVCUAXIMCUCLK_delay, PLVCUMCUMAXIICDCBID_delay[2]);
    $setuphold (posedge PLVCUAXIMCUCLK, posedge PLVCUMCUMAXIICDCBRESP[0], 0:0:0, 0:0:0, notifier, , , PLVCUAXIMCUCLK_delay, PLVCUMCUMAXIICDCBRESP_delay[0]);
    $setuphold (posedge PLVCUAXIMCUCLK, posedge PLVCUMCUMAXIICDCBRESP[1], 0:0:0, 0:0:0, notifier, , , PLVCUAXIMCUCLK_delay, PLVCUMCUMAXIICDCBRESP_delay[1]);
    $setuphold (posedge PLVCUAXIMCUCLK, posedge PLVCUMCUMAXIICDCBVALID, 0:0:0, 0:0:0, notifier, , , PLVCUAXIMCUCLK_delay, PLVCUMCUMAXIICDCBVALID_delay);
    $setuphold (posedge PLVCUAXIMCUCLK, posedge PLVCUMCUMAXIICDCRDATA[0], 0:0:0, 0:0:0, notifier, , , PLVCUAXIMCUCLK_delay, PLVCUMCUMAXIICDCRDATA_delay[0]);
    $setuphold (posedge PLVCUAXIMCUCLK, posedge PLVCUMCUMAXIICDCRDATA[10], 0:0:0, 0:0:0, notifier, , , PLVCUAXIMCUCLK_delay, PLVCUMCUMAXIICDCRDATA_delay[10]);
    $setuphold (posedge PLVCUAXIMCUCLK, posedge PLVCUMCUMAXIICDCRDATA[11], 0:0:0, 0:0:0, notifier, , , PLVCUAXIMCUCLK_delay, PLVCUMCUMAXIICDCRDATA_delay[11]);
    $setuphold (posedge PLVCUAXIMCUCLK, posedge PLVCUMCUMAXIICDCRDATA[12], 0:0:0, 0:0:0, notifier, , , PLVCUAXIMCUCLK_delay, PLVCUMCUMAXIICDCRDATA_delay[12]);
    $setuphold (posedge PLVCUAXIMCUCLK, posedge PLVCUMCUMAXIICDCRDATA[13], 0:0:0, 0:0:0, notifier, , , PLVCUAXIMCUCLK_delay, PLVCUMCUMAXIICDCRDATA_delay[13]);
    $setuphold (posedge PLVCUAXIMCUCLK, posedge PLVCUMCUMAXIICDCRDATA[14], 0:0:0, 0:0:0, notifier, , , PLVCUAXIMCUCLK_delay, PLVCUMCUMAXIICDCRDATA_delay[14]);
    $setuphold (posedge PLVCUAXIMCUCLK, posedge PLVCUMCUMAXIICDCRDATA[15], 0:0:0, 0:0:0, notifier, , , PLVCUAXIMCUCLK_delay, PLVCUMCUMAXIICDCRDATA_delay[15]);
    $setuphold (posedge PLVCUAXIMCUCLK, posedge PLVCUMCUMAXIICDCRDATA[16], 0:0:0, 0:0:0, notifier, , , PLVCUAXIMCUCLK_delay, PLVCUMCUMAXIICDCRDATA_delay[16]);
    $setuphold (posedge PLVCUAXIMCUCLK, posedge PLVCUMCUMAXIICDCRDATA[17], 0:0:0, 0:0:0, notifier, , , PLVCUAXIMCUCLK_delay, PLVCUMCUMAXIICDCRDATA_delay[17]);
    $setuphold (posedge PLVCUAXIMCUCLK, posedge PLVCUMCUMAXIICDCRDATA[18], 0:0:0, 0:0:0, notifier, , , PLVCUAXIMCUCLK_delay, PLVCUMCUMAXIICDCRDATA_delay[18]);
    $setuphold (posedge PLVCUAXIMCUCLK, posedge PLVCUMCUMAXIICDCRDATA[19], 0:0:0, 0:0:0, notifier, , , PLVCUAXIMCUCLK_delay, PLVCUMCUMAXIICDCRDATA_delay[19]);
    $setuphold (posedge PLVCUAXIMCUCLK, posedge PLVCUMCUMAXIICDCRDATA[1], 0:0:0, 0:0:0, notifier, , , PLVCUAXIMCUCLK_delay, PLVCUMCUMAXIICDCRDATA_delay[1]);
    $setuphold (posedge PLVCUAXIMCUCLK, posedge PLVCUMCUMAXIICDCRDATA[20], 0:0:0, 0:0:0, notifier, , , PLVCUAXIMCUCLK_delay, PLVCUMCUMAXIICDCRDATA_delay[20]);
    $setuphold (posedge PLVCUAXIMCUCLK, posedge PLVCUMCUMAXIICDCRDATA[21], 0:0:0, 0:0:0, notifier, , , PLVCUAXIMCUCLK_delay, PLVCUMCUMAXIICDCRDATA_delay[21]);
    $setuphold (posedge PLVCUAXIMCUCLK, posedge PLVCUMCUMAXIICDCRDATA[22], 0:0:0, 0:0:0, notifier, , , PLVCUAXIMCUCLK_delay, PLVCUMCUMAXIICDCRDATA_delay[22]);
    $setuphold (posedge PLVCUAXIMCUCLK, posedge PLVCUMCUMAXIICDCRDATA[23], 0:0:0, 0:0:0, notifier, , , PLVCUAXIMCUCLK_delay, PLVCUMCUMAXIICDCRDATA_delay[23]);
    $setuphold (posedge PLVCUAXIMCUCLK, posedge PLVCUMCUMAXIICDCRDATA[24], 0:0:0, 0:0:0, notifier, , , PLVCUAXIMCUCLK_delay, PLVCUMCUMAXIICDCRDATA_delay[24]);
    $setuphold (posedge PLVCUAXIMCUCLK, posedge PLVCUMCUMAXIICDCRDATA[25], 0:0:0, 0:0:0, notifier, , , PLVCUAXIMCUCLK_delay, PLVCUMCUMAXIICDCRDATA_delay[25]);
    $setuphold (posedge PLVCUAXIMCUCLK, posedge PLVCUMCUMAXIICDCRDATA[26], 0:0:0, 0:0:0, notifier, , , PLVCUAXIMCUCLK_delay, PLVCUMCUMAXIICDCRDATA_delay[26]);
    $setuphold (posedge PLVCUAXIMCUCLK, posedge PLVCUMCUMAXIICDCRDATA[27], 0:0:0, 0:0:0, notifier, , , PLVCUAXIMCUCLK_delay, PLVCUMCUMAXIICDCRDATA_delay[27]);
    $setuphold (posedge PLVCUAXIMCUCLK, posedge PLVCUMCUMAXIICDCRDATA[28], 0:0:0, 0:0:0, notifier, , , PLVCUAXIMCUCLK_delay, PLVCUMCUMAXIICDCRDATA_delay[28]);
    $setuphold (posedge PLVCUAXIMCUCLK, posedge PLVCUMCUMAXIICDCRDATA[29], 0:0:0, 0:0:0, notifier, , , PLVCUAXIMCUCLK_delay, PLVCUMCUMAXIICDCRDATA_delay[29]);
    $setuphold (posedge PLVCUAXIMCUCLK, posedge PLVCUMCUMAXIICDCRDATA[2], 0:0:0, 0:0:0, notifier, , , PLVCUAXIMCUCLK_delay, PLVCUMCUMAXIICDCRDATA_delay[2]);
    $setuphold (posedge PLVCUAXIMCUCLK, posedge PLVCUMCUMAXIICDCRDATA[30], 0:0:0, 0:0:0, notifier, , , PLVCUAXIMCUCLK_delay, PLVCUMCUMAXIICDCRDATA_delay[30]);
    $setuphold (posedge PLVCUAXIMCUCLK, posedge PLVCUMCUMAXIICDCRDATA[31], 0:0:0, 0:0:0, notifier, , , PLVCUAXIMCUCLK_delay, PLVCUMCUMAXIICDCRDATA_delay[31]);
    $setuphold (posedge PLVCUAXIMCUCLK, posedge PLVCUMCUMAXIICDCRDATA[3], 0:0:0, 0:0:0, notifier, , , PLVCUAXIMCUCLK_delay, PLVCUMCUMAXIICDCRDATA_delay[3]);
    $setuphold (posedge PLVCUAXIMCUCLK, posedge PLVCUMCUMAXIICDCRDATA[4], 0:0:0, 0:0:0, notifier, , , PLVCUAXIMCUCLK_delay, PLVCUMCUMAXIICDCRDATA_delay[4]);
    $setuphold (posedge PLVCUAXIMCUCLK, posedge PLVCUMCUMAXIICDCRDATA[5], 0:0:0, 0:0:0, notifier, , , PLVCUAXIMCUCLK_delay, PLVCUMCUMAXIICDCRDATA_delay[5]);
    $setuphold (posedge PLVCUAXIMCUCLK, posedge PLVCUMCUMAXIICDCRDATA[6], 0:0:0, 0:0:0, notifier, , , PLVCUAXIMCUCLK_delay, PLVCUMCUMAXIICDCRDATA_delay[6]);
    $setuphold (posedge PLVCUAXIMCUCLK, posedge PLVCUMCUMAXIICDCRDATA[7], 0:0:0, 0:0:0, notifier, , , PLVCUAXIMCUCLK_delay, PLVCUMCUMAXIICDCRDATA_delay[7]);
    $setuphold (posedge PLVCUAXIMCUCLK, posedge PLVCUMCUMAXIICDCRDATA[8], 0:0:0, 0:0:0, notifier, , , PLVCUAXIMCUCLK_delay, PLVCUMCUMAXIICDCRDATA_delay[8]);
    $setuphold (posedge PLVCUAXIMCUCLK, posedge PLVCUMCUMAXIICDCRDATA[9], 0:0:0, 0:0:0, notifier, , , PLVCUAXIMCUCLK_delay, PLVCUMCUMAXIICDCRDATA_delay[9]);
    $setuphold (posedge PLVCUAXIMCUCLK, posedge PLVCUMCUMAXIICDCRID[0], 0:0:0, 0:0:0, notifier, , , PLVCUAXIMCUCLK_delay, PLVCUMCUMAXIICDCRID_delay[0]);
    $setuphold (posedge PLVCUAXIMCUCLK, posedge PLVCUMCUMAXIICDCRID[1], 0:0:0, 0:0:0, notifier, , , PLVCUAXIMCUCLK_delay, PLVCUMCUMAXIICDCRID_delay[1]);
    $setuphold (posedge PLVCUAXIMCUCLK, posedge PLVCUMCUMAXIICDCRID[2], 0:0:0, 0:0:0, notifier, , , PLVCUAXIMCUCLK_delay, PLVCUMCUMAXIICDCRID_delay[2]);
    $setuphold (posedge PLVCUAXIMCUCLK, posedge PLVCUMCUMAXIICDCRLAST, 0:0:0, 0:0:0, notifier, , , PLVCUAXIMCUCLK_delay, PLVCUMCUMAXIICDCRLAST_delay);
    $setuphold (posedge PLVCUAXIMCUCLK, posedge PLVCUMCUMAXIICDCRRESP[0], 0:0:0, 0:0:0, notifier, , , PLVCUAXIMCUCLK_delay, PLVCUMCUMAXIICDCRRESP_delay[0]);
    $setuphold (posedge PLVCUAXIMCUCLK, posedge PLVCUMCUMAXIICDCRRESP[1], 0:0:0, 0:0:0, notifier, , , PLVCUAXIMCUCLK_delay, PLVCUMCUMAXIICDCRRESP_delay[1]);
    $setuphold (posedge PLVCUAXIMCUCLK, posedge PLVCUMCUMAXIICDCRVALID, 0:0:0, 0:0:0, notifier, , , PLVCUAXIMCUCLK_delay, PLVCUMCUMAXIICDCRVALID_delay);
    $setuphold (posedge PLVCUAXIMCUCLK, posedge PLVCUMCUMAXIICDCWREADY, 0:0:0, 0:0:0, notifier, , , PLVCUAXIMCUCLK_delay, PLVCUMCUMAXIICDCWREADY_delay);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[0], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[0]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[100], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[100]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[101], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[101]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[102], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[102]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[103], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[103]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[104], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[104]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[105], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[105]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[106], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[106]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[107], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[107]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[108], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[108]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[109], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[109]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[10], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[10]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[110], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[110]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[111], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[111]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[112], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[112]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[113], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[113]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[114], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[114]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[115], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[115]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[116], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[116]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[117], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[117]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[118], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[118]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[119], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[119]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[11], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[11]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[120], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[120]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[121], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[121]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[122], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[122]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[123], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[123]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[124], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[124]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[125], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[125]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[126], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[126]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[127], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[127]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[128], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[128]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[129], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[129]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[12], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[12]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[130], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[130]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[131], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[131]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[132], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[132]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[133], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[133]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[134], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[134]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[135], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[135]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[136], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[136]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[137], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[137]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[138], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[138]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[139], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[139]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[13], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[13]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[140], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[140]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[141], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[141]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[142], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[142]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[143], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[143]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[144], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[144]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[145], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[145]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[146], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[146]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[147], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[147]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[148], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[148]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[149], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[149]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[14], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[14]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[150], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[150]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[151], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[151]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[152], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[152]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[153], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[153]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[154], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[154]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[155], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[155]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[156], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[156]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[157], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[157]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[158], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[158]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[159], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[159]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[15], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[15]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[160], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[160]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[161], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[161]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[162], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[162]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[163], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[163]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[164], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[164]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[165], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[165]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[166], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[166]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[167], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[167]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[168], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[168]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[169], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[169]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[16], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[16]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[170], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[170]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[171], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[171]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[172], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[172]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[173], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[173]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[174], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[174]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[175], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[175]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[176], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[176]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[177], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[177]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[178], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[178]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[179], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[179]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[17], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[17]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[180], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[180]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[181], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[181]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[182], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[182]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[183], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[183]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[184], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[184]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[185], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[185]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[186], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[186]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[187], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[187]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[188], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[188]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[189], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[189]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[18], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[18]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[190], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[190]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[191], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[191]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[192], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[192]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[193], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[193]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[194], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[194]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[195], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[195]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[196], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[196]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[197], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[197]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[198], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[198]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[199], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[199]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[19], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[19]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[1], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[1]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[200], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[200]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[201], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[201]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[202], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[202]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[203], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[203]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[204], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[204]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[205], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[205]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[206], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[206]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[207], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[207]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[208], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[208]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[209], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[209]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[20], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[20]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[210], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[210]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[211], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[211]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[212], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[212]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[213], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[213]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[214], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[214]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[215], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[215]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[216], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[216]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[217], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[217]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[218], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[218]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[219], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[219]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[21], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[21]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[220], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[220]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[221], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[221]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[222], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[222]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[223], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[223]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[224], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[224]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[225], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[225]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[226], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[226]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[227], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[227]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[228], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[228]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[229], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[229]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[22], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[22]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[230], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[230]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[231], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[231]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[232], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[232]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[233], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[233]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[234], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[234]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[235], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[235]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[236], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[236]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[237], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[237]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[238], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[238]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[239], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[239]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[23], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[23]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[240], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[240]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[241], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[241]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[242], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[242]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[243], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[243]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[244], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[244]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[245], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[245]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[246], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[246]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[247], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[247]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[248], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[248]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[249], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[249]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[24], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[24]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[250], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[250]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[251], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[251]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[252], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[252]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[253], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[253]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[254], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[254]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[255], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[255]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[256], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[256]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[257], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[257]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[258], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[258]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[259], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[259]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[25], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[25]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[260], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[260]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[261], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[261]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[262], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[262]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[263], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[263]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[264], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[264]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[265], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[265]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[266], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[266]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[267], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[267]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[268], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[268]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[269], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[269]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[26], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[26]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[270], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[270]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[271], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[271]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[272], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[272]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[273], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[273]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[274], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[274]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[275], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[275]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[276], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[276]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[277], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[277]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[278], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[278]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[279], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[279]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[27], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[27]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[280], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[280]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[281], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[281]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[282], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[282]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[283], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[283]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[284], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[284]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[285], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[285]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[286], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[286]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[287], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[287]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[288], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[288]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[289], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[289]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[28], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[28]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[290], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[290]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[291], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[291]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[292], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[292]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[293], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[293]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[294], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[294]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[295], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[295]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[296], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[296]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[297], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[297]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[298], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[298]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[299], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[299]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[29], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[29]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[2], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[2]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[300], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[300]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[301], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[301]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[302], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[302]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[303], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[303]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[304], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[304]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[305], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[305]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[306], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[306]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[307], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[307]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[308], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[308]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[309], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[309]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[30], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[30]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[310], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[310]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[311], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[311]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[312], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[312]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[313], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[313]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[314], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[314]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[315], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[315]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[316], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[316]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[317], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[317]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[318], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[318]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[319], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[319]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[31], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[31]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[32], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[32]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[33], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[33]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[34], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[34]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[35], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[35]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[36], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[36]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[37], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[37]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[38], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[38]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[39], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[39]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[3], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[3]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[40], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[40]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[41], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[41]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[42], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[42]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[43], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[43]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[44], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[44]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[45], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[45]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[46], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[46]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[47], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[47]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[48], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[48]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[49], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[49]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[4], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[4]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[50], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[50]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[51], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[51]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[52], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[52]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[53], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[53]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[54], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[54]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[55], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[55]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[56], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[56]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[57], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[57]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[58], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[58]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[59], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[59]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[5], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[5]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[60], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[60]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[61], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[61]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[62], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[62]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[63], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[63]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[64], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[64]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[65], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[65]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[66], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[66]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[67], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[67]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[68], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[68]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[69], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[69]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[6], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[6]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[70], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[70]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[71], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[71]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[72], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[72]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[73], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[73]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[74], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[74]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[75], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[75]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[76], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[76]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[77], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[77]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[78], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[78]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[79], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[79]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[7], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[7]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[80], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[80]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[81], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[81]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[82], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[82]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[83], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[83]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[84], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[84]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[85], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[85]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[86], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[86]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[87], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[87]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[88], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[88]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[89], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[89]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[8], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[8]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[90], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[90]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[91], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[91]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[92], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[92]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[93], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[93]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[94], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[94]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[95], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[95]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[96], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[96]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[97], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[97]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[98], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[98]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[99], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[99]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRDATA[9], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[9]);
    $setuphold (posedge PLVCUENCL2CCLK, negedge PLVCUENCALL2CRREADY, 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRREADY_delay);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[0], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[0]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[100], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[100]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[101], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[101]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[102], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[102]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[103], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[103]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[104], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[104]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[105], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[105]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[106], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[106]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[107], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[107]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[108], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[108]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[109], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[109]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[10], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[10]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[110], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[110]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[111], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[111]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[112], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[112]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[113], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[113]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[114], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[114]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[115], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[115]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[116], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[116]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[117], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[117]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[118], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[118]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[119], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[119]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[11], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[11]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[120], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[120]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[121], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[121]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[122], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[122]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[123], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[123]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[124], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[124]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[125], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[125]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[126], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[126]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[127], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[127]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[128], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[128]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[129], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[129]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[12], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[12]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[130], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[130]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[131], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[131]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[132], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[132]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[133], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[133]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[134], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[134]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[135], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[135]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[136], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[136]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[137], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[137]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[138], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[138]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[139], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[139]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[13], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[13]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[140], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[140]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[141], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[141]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[142], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[142]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[143], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[143]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[144], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[144]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[145], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[145]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[146], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[146]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[147], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[147]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[148], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[148]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[149], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[149]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[14], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[14]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[150], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[150]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[151], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[151]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[152], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[152]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[153], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[153]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[154], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[154]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[155], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[155]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[156], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[156]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[157], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[157]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[158], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[158]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[159], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[159]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[15], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[15]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[160], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[160]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[161], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[161]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[162], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[162]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[163], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[163]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[164], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[164]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[165], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[165]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[166], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[166]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[167], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[167]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[168], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[168]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[169], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[169]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[16], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[16]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[170], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[170]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[171], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[171]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[172], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[172]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[173], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[173]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[174], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[174]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[175], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[175]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[176], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[176]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[177], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[177]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[178], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[178]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[179], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[179]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[17], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[17]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[180], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[180]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[181], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[181]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[182], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[182]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[183], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[183]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[184], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[184]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[185], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[185]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[186], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[186]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[187], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[187]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[188], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[188]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[189], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[189]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[18], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[18]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[190], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[190]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[191], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[191]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[192], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[192]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[193], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[193]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[194], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[194]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[195], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[195]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[196], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[196]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[197], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[197]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[198], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[198]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[199], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[199]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[19], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[19]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[1], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[1]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[200], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[200]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[201], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[201]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[202], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[202]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[203], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[203]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[204], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[204]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[205], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[205]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[206], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[206]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[207], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[207]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[208], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[208]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[209], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[209]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[20], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[20]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[210], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[210]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[211], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[211]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[212], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[212]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[213], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[213]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[214], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[214]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[215], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[215]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[216], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[216]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[217], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[217]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[218], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[218]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[219], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[219]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[21], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[21]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[220], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[220]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[221], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[221]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[222], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[222]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[223], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[223]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[224], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[224]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[225], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[225]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[226], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[226]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[227], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[227]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[228], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[228]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[229], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[229]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[22], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[22]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[230], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[230]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[231], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[231]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[232], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[232]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[233], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[233]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[234], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[234]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[235], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[235]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[236], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[236]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[237], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[237]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[238], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[238]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[239], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[239]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[23], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[23]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[240], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[240]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[241], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[241]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[242], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[242]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[243], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[243]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[244], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[244]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[245], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[245]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[246], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[246]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[247], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[247]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[248], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[248]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[249], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[249]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[24], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[24]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[250], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[250]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[251], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[251]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[252], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[252]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[253], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[253]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[254], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[254]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[255], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[255]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[256], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[256]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[257], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[257]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[258], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[258]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[259], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[259]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[25], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[25]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[260], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[260]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[261], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[261]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[262], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[262]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[263], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[263]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[264], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[264]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[265], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[265]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[266], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[266]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[267], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[267]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[268], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[268]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[269], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[269]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[26], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[26]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[270], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[270]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[271], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[271]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[272], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[272]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[273], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[273]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[274], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[274]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[275], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[275]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[276], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[276]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[277], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[277]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[278], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[278]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[279], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[279]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[27], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[27]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[280], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[280]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[281], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[281]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[282], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[282]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[283], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[283]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[284], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[284]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[285], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[285]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[286], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[286]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[287], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[287]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[288], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[288]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[289], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[289]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[28], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[28]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[290], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[290]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[291], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[291]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[292], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[292]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[293], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[293]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[294], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[294]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[295], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[295]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[296], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[296]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[297], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[297]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[298], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[298]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[299], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[299]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[29], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[29]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[2], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[2]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[300], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[300]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[301], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[301]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[302], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[302]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[303], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[303]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[304], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[304]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[305], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[305]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[306], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[306]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[307], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[307]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[308], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[308]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[309], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[309]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[30], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[30]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[310], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[310]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[311], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[311]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[312], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[312]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[313], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[313]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[314], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[314]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[315], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[315]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[316], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[316]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[317], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[317]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[318], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[318]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[319], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[319]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[31], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[31]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[32], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[32]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[33], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[33]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[34], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[34]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[35], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[35]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[36], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[36]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[37], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[37]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[38], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[38]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[39], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[39]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[3], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[3]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[40], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[40]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[41], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[41]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[42], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[42]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[43], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[43]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[44], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[44]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[45], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[45]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[46], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[46]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[47], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[47]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[48], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[48]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[49], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[49]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[4], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[4]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[50], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[50]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[51], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[51]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[52], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[52]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[53], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[53]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[54], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[54]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[55], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[55]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[56], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[56]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[57], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[57]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[58], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[58]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[59], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[59]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[5], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[5]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[60], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[60]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[61], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[61]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[62], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[62]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[63], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[63]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[64], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[64]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[65], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[65]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[66], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[66]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[67], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[67]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[68], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[68]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[69], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[69]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[6], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[6]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[70], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[70]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[71], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[71]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[72], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[72]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[73], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[73]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[74], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[74]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[75], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[75]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[76], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[76]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[77], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[77]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[78], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[78]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[79], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[79]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[7], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[7]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[80], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[80]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[81], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[81]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[82], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[82]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[83], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[83]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[84], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[84]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[85], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[85]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[86], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[86]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[87], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[87]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[88], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[88]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[89], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[89]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[8], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[8]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[90], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[90]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[91], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[91]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[92], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[92]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[93], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[93]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[94], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[94]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[95], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[95]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[96], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[96]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[97], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[97]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[98], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[98]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[99], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[99]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRDATA[9], 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRDATA_delay[9]);
    $setuphold (posedge PLVCUENCL2CCLK, posedge PLVCUENCALL2CRREADY, 0:0:0, 0:0:0, notifier, , , PLVCUENCL2CCLK_delay, PLVCUENCALL2CRREADY_delay);
    $width (negedge PLVCUAXIDECCLK, 0:0:0, 0, notifier);
    $width (negedge PLVCUAXIENCCLK, 0:0:0, 0, notifier);
    $width (negedge PLVCUAXILITECLK, 0:0:0, 0, notifier);
    $width (negedge PLVCUAXIMCUCLK, 0:0:0, 0, notifier);
    $width (negedge PLVCUCORECLK, 0:0:0, 0, notifier);
    $width (negedge PLVCUENCL2CCLK, 0:0:0, 0, notifier);
    $width (negedge PLVCUMCUCLK, 0:0:0, 0, notifier);
    $width (negedge PLVCUPLLREFCLKPL, 0:0:0, 0, notifier);
    $width (posedge PLVCUAXIDECCLK, 0:0:0, 0, notifier);
    $width (posedge PLVCUAXIENCCLK, 0:0:0, 0, notifier);
    $width (posedge PLVCUAXILITECLK, 0:0:0, 0, notifier);
    $width (posedge PLVCUAXIMCUCLK, 0:0:0, 0, notifier);
    $width (posedge PLVCUCORECLK, 0:0:0, 0, notifier);
    $width (posedge PLVCUENCL2CCLK, 0:0:0, 0, notifier);
    $width (posedge PLVCUMCUCLK, 0:0:0, 0, notifier);
    $width (posedge PLVCUPLLREFCLKPL, 0:0:0, 0, notifier);
`endif
    specparam PATHPULSE$ = 0;
  endspecify
`endif
endmodule