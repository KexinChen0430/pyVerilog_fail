module outputs
  wire [63 : 0] slave_rdata;
  wire [15 : 0] slave_bid, slave_rid;
  wire [1 : 0] slave_bresp, slave_rresp;
  wire RDY_set_addr_map,
       slave_arready,
       slave_awready,
       slave_bvalid,
       slave_rlast,
       slave_rvalid,
       slave_wready;
  // register rg_addr_base
  reg [63 : 0] rg_addr_base;
  wire [63 : 0] rg_addr_base$D_IN;
  wire rg_addr_base$EN;
  // register rg_addr_lim
  reg [63 : 0] rg_addr_lim;
  wire [63 : 0] rg_addr_lim$D_IN;
  wire rg_addr_lim$EN;
  // register rg_module_ready
  reg rg_module_ready;
  wire rg_module_ready$D_IN, rg_module_ready$EN;
  // ports of submodule slave_xactor_f_rd_addr
  wire [108 : 0] slave_xactor_f_rd_addr$D_IN, slave_xactor_f_rd_addr$D_OUT;
  wire slave_xactor_f_rd_addr$CLR,
       slave_xactor_f_rd_addr$DEQ,
       slave_xactor_f_rd_addr$EMPTY_N,
       slave_xactor_f_rd_addr$ENQ,
       slave_xactor_f_rd_addr$FULL_N;
  // ports of submodule slave_xactor_f_rd_data
  wire [82 : 0] slave_xactor_f_rd_data$D_IN, slave_xactor_f_rd_data$D_OUT;
  wire slave_xactor_f_rd_data$CLR,
       slave_xactor_f_rd_data$DEQ,
       slave_xactor_f_rd_data$EMPTY_N,
       slave_xactor_f_rd_data$ENQ,
       slave_xactor_f_rd_data$FULL_N;
  // ports of submodule slave_xactor_f_wr_addr
  wire [108 : 0] slave_xactor_f_wr_addr$D_IN, slave_xactor_f_wr_addr$D_OUT;
  wire slave_xactor_f_wr_addr$CLR,
       slave_xactor_f_wr_addr$DEQ,
       slave_xactor_f_wr_addr$EMPTY_N,
       slave_xactor_f_wr_addr$ENQ,
       slave_xactor_f_wr_addr$FULL_N;
  // ports of submodule slave_xactor_f_wr_data
  wire [72 : 0] slave_xactor_f_wr_data$D_IN;
  wire slave_xactor_f_wr_data$CLR,
       slave_xactor_f_wr_data$DEQ,
       slave_xactor_f_wr_data$EMPTY_N,
       slave_xactor_f_wr_data$ENQ,
       slave_xactor_f_wr_data$FULL_N;
  // ports of submodule slave_xactor_f_wr_resp
  wire [17 : 0] slave_xactor_f_wr_resp$D_IN, slave_xactor_f_wr_resp$D_OUT;
  wire slave_xactor_f_wr_resp$CLR,
       slave_xactor_f_wr_resp$DEQ,
       slave_xactor_f_wr_resp$EMPTY_N,
       slave_xactor_f_wr_resp$ENQ,
       slave_xactor_f_wr_resp$FULL_N;
  // rule scheduling signals
  wire CAN_FIRE_RL_rl_process_rd_req,
       CAN_FIRE_RL_rl_process_wr_req,
       CAN_FIRE_set_addr_map,
       CAN_FIRE_slave_m_arvalid,
       CAN_FIRE_slave_m_awvalid,
       CAN_FIRE_slave_m_bready,
       CAN_FIRE_slave_m_rready,
       CAN_FIRE_slave_m_wvalid,
       WILL_FIRE_RL_rl_process_rd_req,
       WILL_FIRE_RL_rl_process_wr_req,
       WILL_FIRE_set_addr_map,
       WILL_FIRE_slave_m_arvalid,
       WILL_FIRE_slave_m_awvalid,
       WILL_FIRE_slave_m_bready,
       WILL_FIRE_slave_m_rready,
       WILL_FIRE_slave_m_wvalid;
  // declarations used by system tasks
  // synopsys translate_off
  reg [31 : 0] v__h889;
  reg [31 : 0] v__h6517;
  reg [31 : 0] v__h6810;
  reg [31 : 0] v__h6916;
  reg [31 : 0] v__h883;
  reg [31 : 0] v__h6511;
  reg [31 : 0] v__h6804;
  reg [31 : 0] v__h6910;
  // synopsys translate_on
  // remaining internal signals
  reg [63 : 0] data64__h1057;
  reg [31 : 0] CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q2,
	       CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q3;
  reg CASE_slave_xactor_f_rd_addrD_OUT_BITS_20_TO_1_ETC__q4,
      CASE_slave_xactor_f_wr_addrD_OUT_BITS_20_TO_1_ETC__q5;
  wire [63 : 0] rdata__h1019,
		slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_MIN_ETC__q1;
  wire [1 : 0] rdr_rresp__h1046;
  wire NOT_slave_xactor_f_rd_addr_first_BITS_20_TO_18_ETC___d33,
       NOT_slave_xactor_f_wr_addr_first__223_BITS_20__ETC___d1248;
  // action method set_addr_map
  assign RDY_set_addr_map = 1'd1 ;
  assign CAN_FIRE_set_addr_map = 1'd1 ;
  assign WILL_FIRE_set_addr_map = EN_set_addr_map ;
  // action method slave_m_awvalid
  assign CAN_FIRE_slave_m_awvalid = 1'd1 ;
  assign WILL_FIRE_slave_m_awvalid = 1'd1 ;
  // value method slave_m_awready
  assign slave_awready = slave_xactor_f_wr_addr$FULL_N ;
  // action method slave_m_wvalid
  assign CAN_FIRE_slave_m_wvalid = 1'd1 ;
  assign WILL_FIRE_slave_m_wvalid = 1'd1 ;
  // value method slave_m_wready
  assign slave_wready = slave_xactor_f_wr_data$FULL_N ;
  // value method slave_m_bvalid
  assign slave_bvalid = slave_xactor_f_wr_resp$EMPTY_N ;
  // value method slave_m_bid
  assign slave_bid = slave_xactor_f_wr_resp$D_OUT[17:2] ;
  // value method slave_m_bresp
  assign slave_bresp = slave_xactor_f_wr_resp$D_OUT[1:0] ;
  // action method slave_m_bready
  assign CAN_FIRE_slave_m_bready = 1'd1 ;
  assign WILL_FIRE_slave_m_bready = 1'd1 ;
  // action method slave_m_arvalid
  assign CAN_FIRE_slave_m_arvalid = 1'd1 ;
  assign WILL_FIRE_slave_m_arvalid = 1'd1 ;
  // value method slave_m_arready
  assign slave_arready = slave_xactor_f_rd_addr$FULL_N ;
  // value method slave_m_rvalid
  assign slave_rvalid = slave_xactor_f_rd_data$EMPTY_N ;
  // value method slave_m_rid
  assign slave_rid = slave_xactor_f_rd_data$D_OUT[82:67] ;
  // value method slave_m_rdata
  assign slave_rdata = slave_xactor_f_rd_data$D_OUT[66:3] ;
  // value method slave_m_rresp
  assign slave_rresp = slave_xactor_f_rd_data$D_OUT[2:1] ;
  // value method slave_m_rlast
  assign slave_rlast = slave_xactor_f_rd_data$D_OUT[0] ;
  // action method slave_m_rready
  assign CAN_FIRE_slave_m_rready = 1'd1 ;
  assign WILL_FIRE_slave_m_rready = 1'd1 ;
  // submodule slave_xactor_f_rd_addr
  FIFO2 #(.width(32'd109), .guarded(1'd1)) slave_xactor_f_rd_addr(.RST(RST_N),
								  .CLK(CLK),
								  .D_IN(slave_xactor_f_rd_addr$D_IN),
								  .ENQ(slave_xactor_f_rd_addr$ENQ),
								  .DEQ(slave_xactor_f_rd_addr$DEQ),
								  .CLR(slave_xactor_f_rd_addr$CLR),
								  .D_OUT(slave_xactor_f_rd_addr$D_OUT),
								  .FULL_N(slave_xactor_f_rd_addr$FULL_N),
								  .EMPTY_N(slave_xactor_f_rd_addr$EMPTY_N));
  // submodule slave_xactor_f_rd_data
  FIFO2 #(.width(32'd83), .guarded(1'd1)) slave_xactor_f_rd_data(.RST(RST_N),
								 .CLK(CLK),
								 .D_IN(slave_xactor_f_rd_data$D_IN),
								 .ENQ(slave_xactor_f_rd_data$ENQ),
								 .DEQ(slave_xactor_f_rd_data$DEQ),
								 .CLR(slave_xactor_f_rd_data$CLR),
								 .D_OUT(slave_xactor_f_rd_data$D_OUT),
								 .FULL_N(slave_xactor_f_rd_data$FULL_N),
								 .EMPTY_N(slave_xactor_f_rd_data$EMPTY_N));
  // submodule slave_xactor_f_wr_addr
  FIFO2 #(.width(32'd109), .guarded(1'd1)) slave_xactor_f_wr_addr(.RST(RST_N),
								  .CLK(CLK),
								  .D_IN(slave_xactor_f_wr_addr$D_IN),
								  .ENQ(slave_xactor_f_wr_addr$ENQ),
								  .DEQ(slave_xactor_f_wr_addr$DEQ),
								  .CLR(slave_xactor_f_wr_addr$CLR),
								  .D_OUT(slave_xactor_f_wr_addr$D_OUT),
								  .FULL_N(slave_xactor_f_wr_addr$FULL_N),
								  .EMPTY_N(slave_xactor_f_wr_addr$EMPTY_N));
  // submodule slave_xactor_f_wr_data
  FIFO2 #(.width(32'd73), .guarded(1'd1)) slave_xactor_f_wr_data(.RST(RST_N),
								 .CLK(CLK),
								 .D_IN(slave_xactor_f_wr_data$D_IN),
								 .ENQ(slave_xactor_f_wr_data$ENQ),
								 .DEQ(slave_xactor_f_wr_data$DEQ),
								 .CLR(slave_xactor_f_wr_data$CLR),
								 .D_OUT(),
								 .FULL_N(slave_xactor_f_wr_data$FULL_N),
								 .EMPTY_N(slave_xactor_f_wr_data$EMPTY_N));
  // submodule slave_xactor_f_wr_resp
  FIFO2 #(.width(32'd18), .guarded(1'd1)) slave_xactor_f_wr_resp(.RST(RST_N),
								 .CLK(CLK),
								 .D_IN(slave_xactor_f_wr_resp$D_IN),
								 .ENQ(slave_xactor_f_wr_resp$ENQ),
								 .DEQ(slave_xactor_f_wr_resp$DEQ),
								 .CLR(slave_xactor_f_wr_resp$CLR),
								 .D_OUT(slave_xactor_f_wr_resp$D_OUT),
								 .FULL_N(slave_xactor_f_wr_resp$FULL_N),
								 .EMPTY_N(slave_xactor_f_wr_resp$EMPTY_N));
  // rule RL_rl_process_rd_req
  assign CAN_FIRE_RL_rl_process_rd_req =
	     slave_xactor_f_rd_addr$EMPTY_N &&
	     slave_xactor_f_rd_data$FULL_N &&
	     rg_module_ready ;
  assign WILL_FIRE_RL_rl_process_rd_req = CAN_FIRE_RL_rl_process_rd_req ;
  // rule RL_rl_process_wr_req
  assign CAN_FIRE_RL_rl_process_wr_req =
	     slave_xactor_f_wr_addr$EMPTY_N &&
	     slave_xactor_f_wr_data$EMPTY_N &&
	     slave_xactor_f_wr_resp$FULL_N &&
	     rg_module_ready ;
  assign WILL_FIRE_RL_rl_process_wr_req = CAN_FIRE_RL_rl_process_wr_req ;
  // register rg_addr_base
  assign rg_addr_base$D_IN = set_addr_map_addr_base ;
  assign rg_addr_base$EN = EN_set_addr_map ;
  // register rg_addr_lim
  assign rg_addr_lim$D_IN = set_addr_map_addr_lim ;
  assign rg_addr_lim$EN = EN_set_addr_map ;
  // register rg_module_ready
  assign rg_module_ready$D_IN = 1'd1 ;
  assign rg_module_ready$EN = EN_set_addr_map ;
  // submodule slave_xactor_f_rd_addr
  assign slave_xactor_f_rd_addr$D_IN =
	     { slave_arid,
	       slave_araddr,
	       slave_arlen,
	       slave_arsize,
	       slave_arburst,
	       slave_arlock,
	       slave_arcache,
	       slave_arprot,
	       slave_arqos,
	       slave_arregion } ;
  assign slave_xactor_f_rd_addr$ENQ =
	     slave_arvalid && slave_xactor_f_rd_addr$FULL_N ;
  assign slave_xactor_f_rd_addr$DEQ = CAN_FIRE_RL_rl_process_rd_req ;
  assign slave_xactor_f_rd_addr$CLR = 1'b0 ;
  // submodule slave_xactor_f_rd_data
  assign slave_xactor_f_rd_data$D_IN =
	     { slave_xactor_f_rd_addr$D_OUT[108:93],
	       rdata__h1019,
	       rdr_rresp__h1046,
	       1'd1 } ;
  assign slave_xactor_f_rd_data$ENQ = CAN_FIRE_RL_rl_process_rd_req ;
  assign slave_xactor_f_rd_data$DEQ =
	     slave_rready && slave_xactor_f_rd_data$EMPTY_N ;
  assign slave_xactor_f_rd_data$CLR = 1'b0 ;
  // submodule slave_xactor_f_wr_addr
  assign slave_xactor_f_wr_addr$D_IN =
	     { slave_awid,
	       slave_awaddr,
	       slave_awlen,
	       slave_awsize,
	       slave_awburst,
	       slave_awlock,
	       slave_awcache,
	       slave_awprot,
	       slave_awqos,
	       slave_awregion } ;
  assign slave_xactor_f_wr_addr$ENQ =
	     slave_awvalid && slave_xactor_f_wr_addr$FULL_N ;
  assign slave_xactor_f_wr_addr$DEQ = CAN_FIRE_RL_rl_process_wr_req ;
  assign slave_xactor_f_wr_addr$CLR = 1'b0 ;
  // submodule slave_xactor_f_wr_data
  assign slave_xactor_f_wr_data$D_IN =
	     { slave_wdata, slave_wstrb, slave_wlast } ;
  assign slave_xactor_f_wr_data$ENQ =
	     slave_wvalid && slave_xactor_f_wr_data$FULL_N ;
  assign slave_xactor_f_wr_data$DEQ = CAN_FIRE_RL_rl_process_wr_req ;
  assign slave_xactor_f_wr_data$CLR = 1'b0 ;
  // submodule slave_xactor_f_wr_resp
  assign slave_xactor_f_wr_resp$D_IN =
	     { slave_xactor_f_wr_addr$D_OUT[108:93],
	       NOT_slave_xactor_f_wr_addr_first__223_BITS_20__ETC___d1248 ?
		 2'b10 :
		 2'b0 } ;
  assign slave_xactor_f_wr_resp$ENQ = CAN_FIRE_RL_rl_process_wr_req ;
  assign slave_xactor_f_wr_resp$DEQ =
	     slave_bready && slave_xactor_f_wr_resp$EMPTY_N ;
  assign slave_xactor_f_wr_resp$CLR = 1'b0 ;
  // remaining internal signals
  assign NOT_slave_xactor_f_rd_addr_first_BITS_20_TO_18_ETC___d33 =
	     slave_xactor_f_rd_addr$D_OUT[20:18] != 3'b0 &&
	     CASE_slave_xactor_f_rd_addrD_OUT_BITS_20_TO_1_ETC__q4 ||
	     rg_addr_base > slave_xactor_f_rd_addr$D_OUT[92:29] ||
	     slave_xactor_f_rd_addr$D_OUT[92:29] >= rg_addr_lim ;
  assign NOT_slave_xactor_f_wr_addr_first__223_BITS_20__ETC___d1248 =
	     slave_xactor_f_wr_addr$D_OUT[20:18] != 3'b0 &&
	     CASE_slave_xactor_f_wr_addrD_OUT_BITS_20_TO_1_ETC__q5 ||
	     rg_addr_base > slave_xactor_f_wr_addr$D_OUT[92:29] ||
	     slave_xactor_f_wr_addr$D_OUT[92:29] >= rg_addr_lim ;
  assign rdata__h1019 =
	     NOT_slave_xactor_f_rd_addr_first_BITS_20_TO_18_ETC___d33 ?
	       64'd0 :
	       data64__h1057 ;
  assign rdr_rresp__h1046 =
	     NOT_slave_xactor_f_rd_addr_first_BITS_20_TO_18_ETC___d33 ?
	       2'b10 :
	       2'b0 ;
  assign slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_MIN_ETC__q1 =
	     slave_xactor_f_rd_addr$D_OUT[92:29] - rg_addr_base ;
  always@(slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_MIN_ETC__q1)
  begin
    case (slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_MIN_ETC__q1[63:3])
      61'd2,
      61'd3,
      61'd7,
      61'd9,
      61'd10,
      61'd11,
      61'd25,
      61'd29,
      61'd39,
      61'd53,
      61'd56,
      61'd75,
      61'd91,
      61'd142,
      61'd143,
      61'd144,
      61'd145,
      61'd146,
      61'd147,
      61'd148,
      61'd149,
      61'd150,
      61'd151,
      61'd152,
      61'd153,
      61'd154,
      61'd155,
      61'd156,
      61'd157,
      61'd158,
      61'd159,
      61'd160,
      61'd161,
      61'd162,
      61'd163,
      61'd164,
      61'd165,
      61'd166,
      61'd167,
      61'd168,
      61'd169,
      61'd170,
      61'd171,
      61'd172,
      61'd173,
      61'd174,
      61'd175,
      61'd176,
      61'd177,
      61'd178,
      61'd179,
      61'd180,
      61'd181,
      61'd182,
      61'd183,
      61'd184,
      61'd185,
      61'd186,
      61'd187,
      61'd188,
      61'd189,
      61'd190,
      61'd191,
      61'd192,
      61'd193,
      61'd194,
      61'd195,
      61'd196,
      61'd197,
      61'd198,
      61'd199,
      61'd200,
      61'd201,
      61'd202,
      61'd203,
      61'd204,
      61'd205,
      61'd206,
      61'd207,
      61'd208,
      61'd209,
      61'd210,
      61'd211,
      61'd212,
      61'd213,
      61'd214,
      61'd215,
      61'd216,
      61'd217,
      61'd218,
      61'd219,
      61'd220,
      61'd221,
      61'd222,
      61'd223,
      61'd224,
      61'd225,
      61'd226,
      61'd227,
      61'd228,
      61'd229,
      61'd230,
      61'd231,
      61'd232,
      61'd233,
      61'd234,
      61'd235,
      61'd236,
      61'd237,
      61'd238,
      61'd239,
      61'd240,
      61'd241,
      61'd242,
      61'd243,
      61'd244,
      61'd245,
      61'd246,
      61'd247,
      61'd248,
      61'd249,
      61'd250,
      61'd251,
      61'd252,
      61'd253,
      61'd254,
      61'd255,
      61'd256,
      61'd257,
      61'd258,
      61'd259,
      61'd260,
      61'd261,
      61'd262,
      61'd263,
      61'd264,
      61'd265,
      61'd266,
      61'd267,
      61'd268,
      61'd269,
      61'd270,
      61'd271,
      61'd272,
      61'd273,
      61'd274,
      61'd275,
      61'd276,
      61'd277,
      61'd278,
      61'd279,
      61'd280,
      61'd281,
      61'd282,
      61'd283,
      61'd284,
      61'd285,
      61'd286,
      61'd287,
      61'd288,
      61'd289,
      61'd290,
      61'd291,
      61'd292,
      61'd293,
      61'd294,
      61'd295,
      61'd296,
      61'd297,
      61'd298,
      61'd299,
      61'd300,
      61'd301,
      61'd302,
      61'd303,
      61'd304,
      61'd305,
      61'd306,
      61'd307,
      61'd308,
      61'd309,
      61'd310,
      61'd311,
      61'd312,
      61'd313,
      61'd314,
      61'd315,
      61'd316,
      61'd317,
      61'd318,
      61'd319,
      61'd320,
      61'd321,
      61'd322,
      61'd323,
      61'd324,
      61'd325,
      61'd326,
      61'd327,
      61'd328,
      61'd329,
      61'd330,
      61'd331,
      61'd332,
      61'd333,
      61'd334,
      61'd335,
      61'd336,
      61'd337,
      61'd338,
      61'd339,
      61'd340,
      61'd341,
      61'd342,
      61'd343,
      61'd344,
      61'd345,
      61'd346,
      61'd347,
      61'd348,
      61'd349,
      61'd350,
      61'd351,
      61'd352,
      61'd353,
      61'd354,
      61'd355,
      61'd356,
      61'd357,
      61'd358,
      61'd359,
      61'd360,
      61'd361,
      61'd362,
      61'd363,
      61'd364,
      61'd365,
      61'd366,
      61'd367,
      61'd368,
      61'd369,
      61'd370,
      61'd371,
      61'd372,
      61'd373,
      61'd374,
      61'd375,
      61'd376,
      61'd377,
      61'd378,
      61'd379,
      61'd380,
      61'd381,
      61'd382,
      61'd383,
      61'd384,
      61'd385,
      61'd386,
      61'd387,
      61'd388,
      61'd389,
      61'd390,
      61'd391,
      61'd392,
      61'd393,
      61'd394,
      61'd395,
      61'd396,
      61'd397,
      61'd398,
      61'd399,
      61'd400,
      61'd401,
      61'd402,
      61'd403,
      61'd404,
      61'd405,
      61'd406,
      61'd407,
      61'd408,
      61'd409,
      61'd410,
      61'd411,
      61'd412,
      61'd413,
      61'd414,
      61'd415,
      61'd416,
      61'd417,
      61'd418,
      61'd419,
      61'd420,
      61'd421,
      61'd422,
      61'd423,
      61'd424,
      61'd425,
      61'd426,
      61'd427,
      61'd428,
      61'd429,
      61'd430,
      61'd431,
      61'd432,
      61'd433,
      61'd434,
      61'd435,
      61'd436,
      61'd437,
      61'd438,
      61'd439,
      61'd440,
      61'd441,
      61'd442,
      61'd443,
      61'd444,
      61'd445,
      61'd446,
      61'd447,
      61'd448,
      61'd449,
      61'd450,
      61'd451,
      61'd452,
      61'd453,
      61'd454,
      61'd455,
      61'd456,
      61'd457,
      61'd458,
      61'd459,
      61'd460,
      61'd461,
      61'd462,
      61'd463,
      61'd464,
      61'd465,
      61'd466,
      61'd467,
      61'd468,
      61'd469,
      61'd470,
      61'd471,
      61'd472,
      61'd473,
      61'd474,
      61'd475,
      61'd476,
      61'd477,
      61'd478,
      61'd479,
      61'd480,
      61'd481,
      61'd482,
      61'd483,
      61'd484,
      61'd485,
      61'd486,
      61'd487,
      61'd488,
      61'd489,
      61'd490,
      61'd491,
      61'd492,
      61'd493,
      61'd494,
      61'd495,
      61'd496,
      61'd497,
      61'd498,
      61'd499,
      61'd500,
      61'd501,
      61'd502,
      61'd503,
      61'd504,
      61'd505,
      61'd506,
      61'd507,
      61'd508,
      61'd509,
      61'd510,
      61'd511:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q2 = 32'h0;
      61'd4:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q2 =
	      32'h54040000;
      61'd5:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q2 =
	      32'h88030000;
      61'd6:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q2 =
	      32'h11000000;
      61'd8:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q2 =
	      32'h50030000;
      61'd12,
      61'd14,
      61'd26,
      61'd28,
      61'd30,
      61'd54,
      61'd61,
      61'd109,
      61'd111:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q2 =
	      32'h04000000;
      61'd13, 61'd15, 61'd63, 61'd99, 61'd115:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q2 =
	      32'h02000000;
      61'd16:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q2 =
	      32'h16000000;
      61'd17:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q2 =
	      32'h62626375;
      61'd18:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q2 =
	      32'h656B6970;
      61'd19:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q2 =
	      32'h65642D65;
      61'd20,
      61'd33,
      61'd35,
      61'd37,
      61'd42,
      61'd45,
      61'd48,
      61'd57,
      61'd69,
      61'd74,
      61'd76,
      61'd78,
      61'd84,
      61'd88,
      61'd95,
      61'd102,
      61'd105,
      61'd110:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q2 =
	      32'h03000000;
      61'd21:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q2 =
	      32'h26000000;
      61'd22, 61'd80:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q2 =
	      32'h732C7261;
      61'd23, 61'd81:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q2 =
	      32'h7261622D;
      61'd24,
      61'd27,
      61'd50,
      61'd55,
      61'd62,
      61'd64,
      61'd73,
      61'd93,
      61'd94,
      61'd114:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q2 =
	      32'h01000000;
      61'd31, 61'd112:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q2 =
	      32'h80969800;
      61'd32:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q2 =
	      32'h40757063;
      61'd34:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q2 =
	      32'h3F000000;
      61'd36, 61'd70, 61'd96, 61'd106:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q2 =
	      32'h4B000000;
      61'd38:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q2 =
	      32'h4F000000;
      61'd40:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q2 =
	      32'h06000000;
      61'd41:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q2 =
	      32'h63736972;
      61'd43:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q2 =
	      32'h56000000;
      61'd44:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q2 =
	      32'h75616D69;
      61'd46:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q2 =
	      32'h60000000;
      61'd47:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q2 =
	      32'h76732C76;
      61'd49:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q2 =
	      32'h69000000;
      61'd51:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q2 =
	      32'h70757272;
      61'd52:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q2 =
	      32'h6F72746E;
      61'd58, 61'd79, 61'd89, 61'd103:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q2 =
	      32'h1B000000;
      61'd59:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q2 =
	      32'h70632C76;
      61'd60:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q2 =
	      32'h00006374;
      61'd65:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q2 =
	      32'h38407972;
      61'd66:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q2 =
	      32'h00303030;
      61'd67:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q2 =
	      32'h07000000;
      61'd68:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q2 =
	      32'h6F6D656D;
      61'd71:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q2 =
	      32'h00000080;
      61'd72:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q2 =
	      32'h00000010;
      61'd77:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q2 =
	      32'h0F000000;
      61'd82:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q2 =
	      32'h69730063;
      61'd83:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q2 =
	      32'h7375622D;
      61'd85:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q2 =
	      32'hA7000000;
      61'd86:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q2 =
	      32'h6E696C63;
      61'd87, 61'd101:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q2 =
	      32'h30303030;
      61'd90:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q2 =
	      32'h6C632C76;
      61'd92:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q2 =
	      32'h10000000;
      61'd97:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q2 =
	      32'h00000002;
      61'd98:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q2 =
	      32'h00000C00;
      61'd100:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q2 =
	      32'h74726175;
      61'd104:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q2 =
	      32'h61303535;
      61'd107:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q2 =
	      32'h000000C0;
      61'd108:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q2 =
	      32'h40000000;
      61'd113:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q2 =
	      32'h08000000;
      61'd116:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q2 =
	      32'h09000000;
      61'd117:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q2 =
	      32'h73736572;
      61'd118:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q2 =
	      32'h2300736C;
      61'd119:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q2 =
	      32'h6C65632D;
      61'd120:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q2 =
	      32'h61706D6F;
      61'd121:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q2 =
	      32'h6F6D0065;
      61'd122:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q2 =
	      32'h656D6974;
      61'd123:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q2 =
	      32'h6572662D;
      61'd124:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q2 =
	      32'h64007963;
      61'd125:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q2 =
	      32'h79745F65;
      61'd126:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q2 =
	      32'h73006765;
      61'd127:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q2 =
	      32'h69720073;
      61'd128:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q2 =
	      32'h00617369;
      61'd129:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q2 =
	      32'h65707974;
      61'd130:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q2 =
	      32'h662D6B63;
      61'd131:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q2 =
	      32'h79636E65;
      61'd132, 61'd134:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q2 =
	      32'h72726574;
      61'd133:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q2 =
	      32'h6C6C6563;
      61'd135:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q2 =
	      32'h746E6F63;
      61'd136:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q2 =
	      32'h70007265;
      61'd137:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q2 =
	      32'h7200656C;
      61'd138:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q2 =
	      32'h6E690073;
      61'd139:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q2 =
	      32'h73747075;
      61'd140:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q2 =
	      32'h65646E65;
      61'd141:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q2 =
	      32'h68732D67;
      default: CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q2 =
		   32'hAAAAAAAA;
    endcase
  end
  always@(slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_MIN_ETC__q1)
  begin
    case (slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_MIN_ETC__q1[63:3])
      61'd2:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q3 =
	      32'h00028067;
      61'd3:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q3 =
	      32'h80000000;
      61'd4:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q3 =
	      32'hEDFE0DD0;
      61'd5:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q3 =
	      32'h38000000;
      61'd6:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q3 =
	      32'h28000000;
      61'd7, 61'd70, 61'd96, 61'd106:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q3 =
	      32'h10000000;
      61'd8:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q3 =
	      32'hCC000000;
      61'd9,
      61'd10,
      61'd13,
      61'd27,
      61'd37,
      61'd71,
      61'd72,
      61'd84,
      61'd85,
      61'd97,
      61'd98,
      61'd105,
      61'd107,
      61'd108,
      61'd143,
      61'd144,
      61'd145,
      61'd146,
      61'd147,
      61'd148,
      61'd149,
      61'd150,
      61'd151,
      61'd152,
      61'd153,
      61'd154,
      61'd155,
      61'd156,
      61'd157,
      61'd158,
      61'd159,
      61'd160,
      61'd161,
      61'd162,
      61'd163,
      61'd164,
      61'd165,
      61'd166,
      61'd167,
      61'd168,
      61'd169,
      61'd170,
      61'd171,
      61'd172,
      61'd173,
      61'd174,
      61'd175,
      61'd176,
      61'd177,
      61'd178,
      61'd179,
      61'd180,
      61'd181,
      61'd182,
      61'd183,
      61'd184,
      61'd185,
      61'd186,
      61'd187,
      61'd188,
      61'd189,
      61'd190,
      61'd191,
      61'd192,
      61'd193,
      61'd194,
      61'd195,
      61'd196,
      61'd197,
      61'd198,
      61'd199,
      61'd200,
      61'd201,
      61'd202,
      61'd203,
      61'd204,
      61'd205,
      61'd206,
      61'd207,
      61'd208,
      61'd209,
      61'd210,
      61'd211,
      61'd212,
      61'd213,
      61'd214,
      61'd215,
      61'd216,
      61'd217,
      61'd218,
      61'd219,
      61'd220,
      61'd221,
      61'd222,
      61'd223,
      61'd224,
      61'd225,
      61'd226,
      61'd227,
      61'd228,
      61'd229,
      61'd230,
      61'd231,
      61'd232,
      61'd233,
      61'd234,
      61'd235,
      61'd236,
      61'd237,
      61'd238,
      61'd239,
      61'd240,
      61'd241,
      61'd242,
      61'd243,
      61'd244,
      61'd245,
      61'd246,
      61'd247,
      61'd248,
      61'd249,
      61'd250,
      61'd251,
      61'd252,
      61'd253,
      61'd254,
      61'd255,
      61'd256,
      61'd257,
      61'd258,
      61'd259,
      61'd260,
      61'd261,
      61'd262,
      61'd263,
      61'd264,
      61'd265,
      61'd266,
      61'd267,
      61'd268,
      61'd269,
      61'd270,
      61'd271,
      61'd272,
      61'd273,
      61'd274,
      61'd275,
      61'd276,
      61'd277,
      61'd278,
      61'd279,
      61'd280,
      61'd281,
      61'd282,
      61'd283,
      61'd284,
      61'd285,
      61'd286,
      61'd287,
      61'd288,
      61'd289,
      61'd290,
      61'd291,
      61'd292,
      61'd293,
      61'd294,
      61'd295,
      61'd296,
      61'd297,
      61'd298,
      61'd299,
      61'd300,
      61'd301,
      61'd302,
      61'd303,
      61'd304,
      61'd305,
      61'd306,
      61'd307,
      61'd308,
      61'd309,
      61'd310,
      61'd311,
      61'd312,
      61'd313,
      61'd314,
      61'd315,
      61'd316,
      61'd317,
      61'd318,
      61'd319,
      61'd320,
      61'd321,
      61'd322,
      61'd323,
      61'd324,
      61'd325,
      61'd326,
      61'd327,
      61'd328,
      61'd329,
      61'd330,
      61'd331,
      61'd332,
      61'd333,
      61'd334,
      61'd335,
      61'd336,
      61'd337,
      61'd338,
      61'd339,
      61'd340,
      61'd341,
      61'd342,
      61'd343,
      61'd344,
      61'd345,
      61'd346,
      61'd347,
      61'd348,
      61'd349,
      61'd350,
      61'd351,
      61'd352,
      61'd353,
      61'd354,
      61'd355,
      61'd356,
      61'd357,
      61'd358,
      61'd359,
      61'd360,
      61'd361,
      61'd362,
      61'd363,
      61'd364,
      61'd365,
      61'd366,
      61'd367,
      61'd368,
      61'd369,
      61'd370,
      61'd371,
      61'd372,
      61'd373,
      61'd374,
      61'd375,
      61'd376,
      61'd377,
      61'd378,
      61'd379,
      61'd380,
      61'd381,
      61'd382,
      61'd383,
      61'd384,
      61'd385,
      61'd386,
      61'd387,
      61'd388,
      61'd389,
      61'd390,
      61'd391,
      61'd392,
      61'd393,
      61'd394,
      61'd395,
      61'd396,
      61'd397,
      61'd398,
      61'd399,
      61'd400,
      61'd401,
      61'd402,
      61'd403,
      61'd404,
      61'd405,
      61'd406,
      61'd407,
      61'd408,
      61'd409,
      61'd410,
      61'd411,
      61'd412,
      61'd413,
      61'd414,
      61'd415,
      61'd416,
      61'd417,
      61'd418,
      61'd419,
      61'd420,
      61'd421,
      61'd422,
      61'd423,
      61'd424,
      61'd425,
      61'd426,
      61'd427,
      61'd428,
      61'd429,
      61'd430,
      61'd431,
      61'd432,
      61'd433,
      61'd434,
      61'd435,
      61'd436,
      61'd437,
      61'd438,
      61'd439,
      61'd440,
      61'd441,
      61'd442,
      61'd443,
      61'd444,
      61'd445,
      61'd446,
      61'd447,
      61'd448,
      61'd449,
      61'd450,
      61'd451,
      61'd452,
      61'd453,
      61'd454,
      61'd455,
      61'd456,
      61'd457,
      61'd458,
      61'd459,
      61'd460,
      61'd461,
      61'd462,
      61'd463,
      61'd464,
      61'd465,
      61'd466,
      61'd467,
      61'd468,
      61'd469,
      61'd470,
      61'd471,
      61'd472,
      61'd473,
      61'd474,
      61'd475,
      61'd476,
      61'd477,
      61'd478,
      61'd479,
      61'd480,
      61'd481,
      61'd482,
      61'd483,
      61'd484,
      61'd485,
      61'd486,
      61'd487,
      61'd488,
      61'd489,
      61'd490,
      61'd491,
      61'd492,
      61'd493,
      61'd494,
      61'd495,
      61'd496,
      61'd497,
      61'd498,
      61'd499,
      61'd500,
      61'd501,
      61'd502,
      61'd503,
      61'd504,
      61'd505,
      61'd506,
      61'd507,
      61'd508,
      61'd509,
      61'd510,
      61'd511:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q3 = 32'h0;
      61'd11, 61'd32, 61'd86, 61'd100:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q3 =
	      32'h01000000;
      61'd12,
      61'd14,
      61'd16,
      61'd26,
      61'd28,
      61'd30,
      61'd40,
      61'd54,
      61'd56,
      61'd61,
      61'd67,
      61'd92,
      61'd94,
      61'd109,
      61'd111,
      61'd113:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q3 =
	      32'h03000000;
      61'd15, 61'd29, 61'd58:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q3 =
	      32'h0F000000;
      61'd17, 61'd41:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q3 =
	      32'h1B000000;
      61'd18:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q3 =
	      32'h732C7261;
      61'd19:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q3 =
	      32'h7261622D;
      61'd20, 61'd42:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q3 =
	      32'h00000076;
      61'd21:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q3 =
	      32'h12000000;
      61'd22, 61'd80:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q3 =
	      32'h62626375;
      61'd23, 61'd81:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q3 =
	      32'h656B6970;
      61'd24:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q3 =
	      32'h00000065;
      61'd25:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q3 =
	      32'h73757063;
      61'd31:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q3 =
	      32'h2C000000;
      61'd33, 61'd88, 61'd102:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q3 =
	      32'h00000030;
      61'd34, 61'd36, 61'd49, 61'd75, 61'd77:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q3 =
	      32'h04000000;
      61'd35:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q3 =
	      32'h00757063;
      61'd38:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q3 =
	      32'h05000000;
      61'd39:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q3 =
	      32'h79616B6F;
      61'd43:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q3 =
	      32'h0A000000;
      61'd44:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q3 =
	      32'h34367672;
      61'd45:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q3 =
	      32'h00000073;
      61'd46, 61'd115:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q3 =
	      32'h0B000000;
      61'd47, 61'd59, 61'd90:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q3 =
	      32'h63736972;
      61'd48:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q3 =
	      32'h00003933;
      61'd50:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q3 =
	      32'h80969800;
      61'd51:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q3 =
	      32'h65746E69;
      61'd52:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q3 =
	      32'h6F632D74;
      61'd53:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q3 =
	      32'h72656C6C;
      61'd55:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q3 =
	      32'h79000000;
      61'd57:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q3 =
	      32'h8A000000;
      61'd60:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q3 =
	      32'h6E692D75;
      61'd62:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q3 =
	      32'h9F000000;
      61'd63, 61'd64, 61'd73, 61'd76, 61'd78, 61'd99, 61'd116:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q3 =
	      32'h02000000;
      61'd65:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q3 =
	      32'h6F6D656D;
      61'd66:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q3 =
	      32'h30303030;
      61'd68:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q3 =
	      32'h3F000000;
      61'd69:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q3 =
	      32'h00007972;
      61'd74:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q3 =
	      32'h00636F73;
      61'd79:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q3 =
	      32'h21000000;
      61'd82:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q3 =
	      32'h6F732D65;
      61'd83:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q3 =
	      32'h656C706D;
      61'd87:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q3 =
	      32'h30324074;
      61'd89:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q3 =
	      32'h0D000000;
      61'd91:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q3 =
	      32'h30746E69;
      61'd93, 61'd114:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q3 =
	      32'hAE000000;
      61'd95:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q3 =
	      32'h07000000;
      61'd101:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q3 =
	      32'h30306340;
      61'd103:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q3 =
	      32'h09000000;
      61'd104:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q3 =
	      32'h3631736E;
      61'd110:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q3 =
	      32'hC2000000;
      61'd112:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q3 =
	      32'h69000000;
      61'd117:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q3 =
	      32'h64646123;
      61'd118:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q3 =
	      32'h6C65632D;
      61'd119:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q3 =
	      32'h657A6973;
      61'd120:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q3 =
	      32'h6300736C;
      61'd121:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q3 =
	      32'h6C626974;
      61'd122:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q3 =
	      32'h006C6564;
      61'd123:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q3 =
	      32'h65736162;
      61'd124:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q3 =
	      32'h6E657571;
      61'd125:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q3 =
	      32'h63697665;
      61'd126:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q3 =
	      32'h72006570;
      61'd127:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q3 =
	      32'h75746174;
      61'd128:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q3 =
	      32'h2C766373;
      61'd129:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q3 =
	      32'h2D756D6D;
      61'd130:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q3 =
	      32'h6F6C6300;
      61'd131:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q3 =
	      32'h75716572;
      61'd132:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q3 =
	      32'h6E692300;
      61'd133, 61'd135:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q3 =
	      32'h2D747075;
      61'd134:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q3 =
	      32'h6E690073;
      61'd136:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q3 =
	      32'h6C6C6F72;
      61'd137:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q3 =
	      32'h646E6168;
      61'd138:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q3 =
	      32'h65676E61;
      61'd139:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q3 =
	      32'h72726574;
      61'd140:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q3 =
	      32'h7478652D;
      61'd141:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q3 =
	      32'h65720064;
      61'd142:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q3 =
	      32'h00746669;
      default: CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q3 =
		   32'hAAAAAAAA;
    endcase
  end
  always@(slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_MIN_ETC__q1 or
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q2 or
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q3)
  begin
    case (slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_MIN_ETC__q1[63:3])
      61'd0: data64__h1057 = 64'h0202859300000297;
      61'd1: data64__h1057 = 64'h0182B283F1402573;
      default: data64__h1057 =
		   { CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q2,
		     CASE_slave_xactor_f_rd_addrD_OUT_BITS_92_TO_29_ETC__q3 };
    endcase
  end
  always@(slave_xactor_f_rd_addr$D_OUT)
  begin
    case (slave_xactor_f_rd_addr$D_OUT[20:18])
      3'b001:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_20_TO_1_ETC__q4 =
	      slave_xactor_f_rd_addr$D_OUT[29];
      3'b010:
	  CASE_slave_xactor_f_rd_addrD_OUT_BITS_20_TO_1_ETC__q4 =
	      slave_xactor_f_rd_addr$D_OUT[30:29] != 2'b0;
      default: CASE_slave_xactor_f_rd_addrD_OUT_BITS_20_TO_1_ETC__q4 =
		   slave_xactor_f_rd_addr$D_OUT[20:18] != 3'b011 ||
		   slave_xactor_f_rd_addr$D_OUT[31:29] != 3'b0;
    endcase
  end
  always@(slave_xactor_f_wr_addr$D_OUT)
  begin
    case (slave_xactor_f_wr_addr$D_OUT[20:18])
      3'b001:
	  CASE_slave_xactor_f_wr_addrD_OUT_BITS_20_TO_1_ETC__q5 =
	      slave_xactor_f_wr_addr$D_OUT[29];
      3'b010:
	  CASE_slave_xactor_f_wr_addrD_OUT_BITS_20_TO_1_ETC__q5 =
	      slave_xactor_f_wr_addr$D_OUT[30:29] != 2'b0;
      default: CASE_slave_xactor_f_wr_addrD_OUT_BITS_20_TO_1_ETC__q5 =
		   slave_xactor_f_wr_addr$D_OUT[20:18] != 3'b011 ||
		   slave_xactor_f_wr_addr$D_OUT[31:29] != 3'b0;
    endcase
  end
  // handling of inlined registers
  always@(posedge CLK)
  begin
    if (RST_N == `BSV_RESET_VALUE)
      begin
        rg_module_ready <= `BSV_ASSIGNMENT_DELAY 1'd0;
      end
    else
      begin
        if (rg_module_ready$EN)
	  rg_module_ready <= `BSV_ASSIGNMENT_DELAY rg_module_ready$D_IN;
      end
    if (rg_addr_base$EN)
      rg_addr_base <= `BSV_ASSIGNMENT_DELAY rg_addr_base$D_IN;
    if (rg_addr_lim$EN) rg_addr_lim <= `BSV_ASSIGNMENT_DELAY rg_addr_lim$D_IN;
  end
  // synopsys translate_off
  `ifdef BSV_NO_INITIAL_BLOCKS
  `else // not BSV_NO_INITIAL_BLOCKS
  initial
  begin
    rg_addr_base = 64'hAAAAAAAAAAAAAAAA;
    rg_addr_lim = 64'hAAAAAAAAAAAAAAAA;
    rg_module_ready = 1'h0;
  end
  `endif // BSV_NO_INITIAL_BLOCKS
  // synopsys translate_on
  // handling of system tasks
  // synopsys translate_off
  always@(negedge CLK)
  begin
    #0;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_rd_req &&
	  NOT_slave_xactor_f_rd_addr_first_BITS_20_TO_18_ETC___d33)
	begin
	  v__h889 = $stime;
	  #0;
	end
    v__h883 = v__h889 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_rd_req &&
	  NOT_slave_xactor_f_rd_addr_first_BITS_20_TO_18_ETC___d33)
	$display("%0d: ERROR: Boot_ROM.rl_process_rd_req: unrecognized or misaligned addr",
		 v__h883);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_rd_req &&
	  NOT_slave_xactor_f_rd_addr_first_BITS_20_TO_18_ETC___d33)
	$write("    ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_rd_req &&
	  NOT_slave_xactor_f_rd_addr_first_BITS_20_TO_18_ETC___d33)
	$write("AXI4_Rd_Addr { ", "arid: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_rd_req &&
	  NOT_slave_xactor_f_rd_addr_first_BITS_20_TO_18_ETC___d33)
	$write("'h%h", slave_xactor_f_rd_addr$D_OUT[108:93]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_rd_req &&
	  NOT_slave_xactor_f_rd_addr_first_BITS_20_TO_18_ETC___d33)
	$write(", ", "araddr: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_rd_req &&
	  NOT_slave_xactor_f_rd_addr_first_BITS_20_TO_18_ETC___d33)
	$write("'h%h", slave_xactor_f_rd_addr$D_OUT[92:29]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_rd_req &&
	  NOT_slave_xactor_f_rd_addr_first_BITS_20_TO_18_ETC___d33)
	$write(", ", "arlen: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_rd_req &&
	  NOT_slave_xactor_f_rd_addr_first_BITS_20_TO_18_ETC___d33)
	$write("'h%h", slave_xactor_f_rd_addr$D_OUT[28:21]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_rd_req &&
	  NOT_slave_xactor_f_rd_addr_first_BITS_20_TO_18_ETC___d33)
	$write(", ", "arsize: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_rd_req &&
	  NOT_slave_xactor_f_rd_addr_first_BITS_20_TO_18_ETC___d33)
	$write("'h%h", slave_xactor_f_rd_addr$D_OUT[20:18]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_rd_req &&
	  NOT_slave_xactor_f_rd_addr_first_BITS_20_TO_18_ETC___d33)
	$write(", ", "arburst: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_rd_req &&
	  NOT_slave_xactor_f_rd_addr_first_BITS_20_TO_18_ETC___d33)
	$write("'h%h", slave_xactor_f_rd_addr$D_OUT[17:16]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_rd_req &&
	  NOT_slave_xactor_f_rd_addr_first_BITS_20_TO_18_ETC___d33)
	$write(", ", "arlock: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_rd_req &&
	  NOT_slave_xactor_f_rd_addr_first_BITS_20_TO_18_ETC___d33)
	$write("'h%h", slave_xactor_f_rd_addr$D_OUT[15]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_rd_req &&
	  NOT_slave_xactor_f_rd_addr_first_BITS_20_TO_18_ETC___d33)
	$write(", ", "arcache: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_rd_req &&
	  NOT_slave_xactor_f_rd_addr_first_BITS_20_TO_18_ETC___d33)
	$write("'h%h", slave_xactor_f_rd_addr$D_OUT[14:11]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_rd_req &&
	  NOT_slave_xactor_f_rd_addr_first_BITS_20_TO_18_ETC___d33)
	$write(", ", "arprot: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_rd_req &&
	  NOT_slave_xactor_f_rd_addr_first_BITS_20_TO_18_ETC___d33)
	$write("'h%h", slave_xactor_f_rd_addr$D_OUT[10:8]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_rd_req &&
	  NOT_slave_xactor_f_rd_addr_first_BITS_20_TO_18_ETC___d33)
	$write(", ", "arqos: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_rd_req &&
	  NOT_slave_xactor_f_rd_addr_first_BITS_20_TO_18_ETC___d33)
	$write("'h%h", slave_xactor_f_rd_addr$D_OUT[7:4]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_rd_req &&
	  NOT_slave_xactor_f_rd_addr_first_BITS_20_TO_18_ETC___d33)
	$write(", ", "arregion: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_rd_req &&
	  NOT_slave_xactor_f_rd_addr_first_BITS_20_TO_18_ETC___d33)
	$write("'h%h", slave_xactor_f_rd_addr$D_OUT[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_rd_req &&
	  NOT_slave_xactor_f_rd_addr_first_BITS_20_TO_18_ETC___d33)
	$write(", ", "aruser: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_rd_req &&
	  NOT_slave_xactor_f_rd_addr_first_BITS_20_TO_18_ETC___d33)
	$write("'h%h", 1'd0, " }");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_rd_req &&
	  NOT_slave_xactor_f_rd_addr_first_BITS_20_TO_18_ETC___d33)
	$write("\n");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_wr_req &&
	  NOT_slave_xactor_f_wr_addr_first__223_BITS_20__ETC___d1248)
	begin
	  v__h6517 = $stime;
	  #0;
	end
    v__h6511 = v__h6517 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_wr_req &&
	  NOT_slave_xactor_f_wr_addr_first__223_BITS_20__ETC___d1248)
	$display("%0d: ERROR: Boot_ROM.rl_process_wr_req: unrecognized or misaligned addr",
		 v__h6511);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_wr_req &&
	  NOT_slave_xactor_f_wr_addr_first__223_BITS_20__ETC___d1248)
	$write("    ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_wr_req &&
	  NOT_slave_xactor_f_wr_addr_first__223_BITS_20__ETC___d1248)
	$write("AXI4_Wr_Addr { ", "awid: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_wr_req &&
	  NOT_slave_xactor_f_wr_addr_first__223_BITS_20__ETC___d1248)
	$write("'h%h", slave_xactor_f_wr_addr$D_OUT[108:93]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_wr_req &&
	  NOT_slave_xactor_f_wr_addr_first__223_BITS_20__ETC___d1248)
	$write(", ", "awaddr: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_wr_req &&
	  NOT_slave_xactor_f_wr_addr_first__223_BITS_20__ETC___d1248)
	$write("'h%h", slave_xactor_f_wr_addr$D_OUT[92:29]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_wr_req &&
	  NOT_slave_xactor_f_wr_addr_first__223_BITS_20__ETC___d1248)
	$write(", ", "awlen: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_wr_req &&
	  NOT_slave_xactor_f_wr_addr_first__223_BITS_20__ETC___d1248)
	$write("'h%h", slave_xactor_f_wr_addr$D_OUT[28:21]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_wr_req &&
	  NOT_slave_xactor_f_wr_addr_first__223_BITS_20__ETC___d1248)
	$write(", ", "awsize: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_wr_req &&
	  NOT_slave_xactor_f_wr_addr_first__223_BITS_20__ETC___d1248)
	$write("'h%h", slave_xactor_f_wr_addr$D_OUT[20:18]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_wr_req &&
	  NOT_slave_xactor_f_wr_addr_first__223_BITS_20__ETC___d1248)
	$write(", ", "awburst: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_wr_req &&
	  NOT_slave_xactor_f_wr_addr_first__223_BITS_20__ETC___d1248)
	$write("'h%h", slave_xactor_f_wr_addr$D_OUT[17:16]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_wr_req &&
	  NOT_slave_xactor_f_wr_addr_first__223_BITS_20__ETC___d1248)
	$write(", ", "awlock: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_wr_req &&
	  NOT_slave_xactor_f_wr_addr_first__223_BITS_20__ETC___d1248)
	$write("'h%h", slave_xactor_f_wr_addr$D_OUT[15]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_wr_req &&
	  NOT_slave_xactor_f_wr_addr_first__223_BITS_20__ETC___d1248)
	$write(", ", "awcache: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_wr_req &&
	  NOT_slave_xactor_f_wr_addr_first__223_BITS_20__ETC___d1248)
	$write("'h%h", slave_xactor_f_wr_addr$D_OUT[14:11]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_wr_req &&
	  NOT_slave_xactor_f_wr_addr_first__223_BITS_20__ETC___d1248)
	$write(", ", "awprot: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_wr_req &&
	  NOT_slave_xactor_f_wr_addr_first__223_BITS_20__ETC___d1248)
	$write("'h%h", slave_xactor_f_wr_addr$D_OUT[10:8]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_wr_req &&
	  NOT_slave_xactor_f_wr_addr_first__223_BITS_20__ETC___d1248)
	$write(", ", "awqos: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_wr_req &&
	  NOT_slave_xactor_f_wr_addr_first__223_BITS_20__ETC___d1248)
	$write("'h%h", slave_xactor_f_wr_addr$D_OUT[7:4]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_wr_req &&
	  NOT_slave_xactor_f_wr_addr_first__223_BITS_20__ETC___d1248)
	$write(", ", "awregion: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_wr_req &&
	  NOT_slave_xactor_f_wr_addr_first__223_BITS_20__ETC___d1248)
	$write("'h%h", slave_xactor_f_wr_addr$D_OUT[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_wr_req &&
	  NOT_slave_xactor_f_wr_addr_first__223_BITS_20__ETC___d1248)
	$write(", ", "awuser: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_wr_req &&
	  NOT_slave_xactor_f_wr_addr_first__223_BITS_20__ETC___d1248)
	$write("'h%h", 1'd0, " }");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_rl_process_wr_req &&
	  NOT_slave_xactor_f_wr_addr_first__223_BITS_20__ETC___d1248)
	$write("\n");
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_set_addr_map && set_addr_map_addr_base[2:0] != 3'd0)
	begin
	  v__h6810 = $stime;
	  #0;
	end
    v__h6804 = v__h6810 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_set_addr_map && set_addr_map_addr_base[2:0] != 3'd0)
	$display("%0d: WARNING: Boot_ROM.set_addr_map: addr_base 0x%0h is not 4-Byte-aligned",
		 v__h6804,
		 set_addr_map_addr_base);
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_set_addr_map && set_addr_map_addr_lim[2:0] != 3'd0)
	begin
	  v__h6916 = $stime;
	  #0;
	end
    v__h6910 = v__h6916 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_set_addr_map && set_addr_map_addr_lim[2:0] != 3'd0)
	$display("%0d: WARNING: Boot_ROM.set_addr_map: addr_lim 0x%0h is not 4-Byte-aligned",
		 v__h6910,
		 set_addr_map_addr_lim);
  end
  // synopsys translate_on
endmodule