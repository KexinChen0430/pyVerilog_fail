module. As an alternative,
// a standard cell from the library could also be directly instanciated here
// (don't forget the "dont_touch" attribute)
//=============================================================================
// 2)  AND GATE
//=============================================================================
assign  y  =  a & b;
endmodule