module cycloneiiils_mux21 (MO, A, B, S);
   input A, B, S;
   output MO;
   wire A_in;
   wire B_in;
   wire S_in;
   buf(A_in, A);
   buf(B_in, B);
   buf(S_in, S);
   wire   tmp_MO;
   specify
      (A => MO) = (0, 0);
      (B => MO) = (0, 0);
      (S => MO) = (0, 0);
   endspecify
   assign tmp_MO = (S_in == 1) ? B_in : A_in;
   buf (MO, tmp_MO);
endmodule