module  al7af2f(
   sys_clk,
   rst_n,
   ofc3555,
   mg1aaad,
   jcd5569,
   jraab4b,
   vv55a5f,
   vkad2fe,
   lq697f3,
   kd4bf9b,
   jp5fcdc,
   lqfe6e7,
   thf373b,
   bn9b9df,
   nt8b8a0,
   ls1e282,
   yxe2831,
   ym3bfe4,
   rib82be,
   icc15f2,
   jpd27c8,
   do93e46,
   mt9f233,
   mt18edf,
   hbc76fc,
   ie3b7e7,
   sudbf39,
   fadf9c9,
   hbfce4b,
   mre725f,
   kf392fc,
   gbc97e4,
   cz4bf24,
   xj5f924,
   vvfc927,
   fp27e80,
   je3f407,
   ayfa03b,
   tue493f,
   mg249fa,
   ie24fd0,
`ifdef AER
   hod01d9,
   sj80ecb,
   ux765d,
   ie3b2ed,
   uvd9769 ,
   uicbb4d,
   jc5da68,
   iped342,
   lq69a15,
   fa4d0aa,
`endif
   lf198b2,
   yxcc596,
   os62cb4,
   fp165a1,
   xyb2d0e,
   ba96872,
   wlb4393,
   uxa1c9c,
   vke4e4,
`ifdef AER
   kd54529,
`endif
   me6705e,
   lf382f0,
   mec1786
   );
parameter uvc3724   = 2'b00;
parameter je1b925  = 2'b01;
parameter mrdc92b = 2'b10;
input                     sys_clk;
input                     rst_n;
input [(8*`NUM_VC)-1:0]  ofc3555;
input [(8*`NUM_VC)-1:0]  mg1aaad;
input [(8*`NUM_VC)-1:0]  jcd5569;
input [(12*`NUM_VC)-1:0] jraab4b;
input [(12*`NUM_VC)-1:0] vv55a5f;
input [(12*`NUM_VC)-1:0] vkad2fe;
input  [6:0]             lq697f3;
input  [10:0]            kd4bf9b;
input  [6:0]             jp5fcdc;
input  [10:0]            lqfe6e7;
input  [6:0]             thf373b;
input  [10:0]            bn9b9df;
input  [11:0]            nt8b8a0;
input [`NUM_VC-1:0]       ls1e282;
input                     yxe2831;
input                     ym3bfe4;
input                     rib82be;
input                     icc15f2;
input [`NUM_VC-1:0]       jpd27c8;
input [`NUM_VC-1:0]       do93e46;
input [`NUM_VC-1:0]       mt9f233;
input [`NUM_VC-1:0]       mt18edf;
input [`NUM_VC-1:0]       hbc76fc;
input [`NUM_VC-1:0]       ie3b7e7;
input [`NUM_VC-1:0]       sudbf39;
input [`NUM_VC-1:0]       fadf9c9;
input [`NUM_VC-1:0]       hbfce4b;
input [`NUM_VC-1:0]       mre725f;
input [`NUM_VC-1:0]       kf392fc;
input [`NUM_VC-1:0]       gbc97e4;
input [`NUM_VC-1:0]       cz4bf24;
input [`NUM_VC-1:0]       xj5f924;
input [`NUM_VC-1:0]       vvfc927;
input                     fp27e80;
input                     je3f407;
input                     ayfa03b;
input [(8*`NUM_VC)-1:0]   tue493f;
input [(8*`NUM_VC)-1:0]   mg249fa;
input [(8*`NUM_VC)-1:0]   ie24fd0;
`ifdef AER
input   [`NUM_VC-1:0]     hod01d9;
input                     sj80ecb;
input                     ux765d;
input                     ie3b2ed;
input                     uvd9769;
input  [8:0]              uicbb4d;
input                     jc5da68;
input                     iped342;
input                     lq69a15;
input                     fa4d0aa;
`endif
output                    lf198b2;
output   [2:0]            yxcc596;
output   [1:0]            os62cb4;
output                    fp165a1;
output   [2:0]            xyb2d0e;
output   [1:0]            ba96872;
output  [`NUM_VC-1:0]     wlb4393;
output  [`NUM_VC-1:0]     uxa1c9c;
output  [`NUM_VC-1:0]     vke4e4;
output [(24*`NUM_VC)-1:0] me6705e;
output [(24*`NUM_VC)-1:0] lf382f0;
output [(24*`NUM_VC)-1:0] mec1786;
`ifdef AER
output                    kd54529;
`endif
integer                     ir85a38;
wire  [`NUM_VC-1:0]         ym1549d;
wire  [`NUM_VC-1:0]         zzaa4e9;
wire  [`NUM_VC-1:0]         ne5274e;
wire  [`NUM_VC-1:0]         je93a72;
wire  [`NUM_VC-1:0]         gq9d393;
wire  [`NUM_VC-1:0]         pfe9c99;
wire  [`NUM_VC-1:0]         mr4e4ce;
wire  [`NUM_VC-1:0]         ay72675;
wire  [`NUM_VC-1:0]         do933a9;
wire  [`NUM_VC-1:0]         hq99d4a;
wire  [`NUM_VC-1:0]         qgcea52;
wire  [`NUM_VC-1:0]         en75290;
wire                        ofe77fc;
wire  [13:0]                ykfa0d0;
reg   [13:0]                rgd0681;
wire  [`NUM_VC -1:0]        tw8340b;
wire  [`NUM_VC -1:0]        aa1a05b;
wire  [`NUM_VC -1:0]        ned02d8;
wire  [`NUM_VC -1:0]        ph816c3;
`ifdef VC1
`else
`endif
`ifdef AER
`endif
`ifdef AER
`endif
reg [(8 * `NUM_VC) - 1 : 0] hq83f1a;
reg [(8 * `NUM_VC) - 1 : 0] ec1f8d2;
reg [(8 * `NUM_VC) - 1 : 0] zxfc691;
reg [(12 * `NUM_VC) - 1 : 0] xje348e;
reg [(12 * `NUM_VC) - 1 : 0] sw1a476;
reg [(12 * `NUM_VC) - 1 : 0] dzd23b0;
reg [6 : 0] jr91d86;
reg [10 : 0] fp8ec36;
reg [6 : 0] tu761b6;
reg [10 : 0] bnb0db3;
reg [6 : 0] ls86d9f;
reg [10 : 0] mt36cfa;
reg [11 : 0] ir95972;
reg [`NUM_VC - 1 : 0] vv7e6c2;
reg al65ca0;
reg an9f508;
reg ofc3f97;
reg ie1fcbc;
reg [`NUM_VC - 1 : 0] mefa844;
reg [`NUM_VC - 1 : 0] uid4220;
reg [`NUM_VC - 1 : 0] sja1101;
reg [`NUM_VC - 1 : 0] ri1b63;
reg [`NUM_VC - 1 : 0] mtdb1b;
reg [`NUM_VC - 1 : 0] ay6d8dd;
reg [`NUM_VC - 1 : 0] vi6c6e8;
reg [`NUM_VC - 1 : 0] lq63743;
reg [`NUM_VC - 1 : 0] ba1ba1a;
reg [`NUM_VC - 1 : 0] bldd0d3;
reg [`NUM_VC - 1 : 0] ale869f;
reg [`NUM_VC - 1 : 0] yk434fd;
reg [`NUM_VC - 1 : 0] ou1a7e9;
reg [`NUM_VC - 1 : 0] wjd3f48;
reg [`NUM_VC - 1 : 0] ir9fa45;
reg fn45b3b;
reg vx2d9df;
reg ho6cefe;
reg [(8 * `NUM_VC) - 1 : 0] enfd22d;
reg [(8 * `NUM_VC) - 1 : 0] lde916c;
reg [(8 * `NUM_VC) - 1 : 0] jc48b67;
reg [`NUM_VC - 1 : 0] dmfe5e1;
reg [`NUM_VC - 1 : 0] gbf2f0b;
reg [`NUM_VC - 1 : 0] uk9785c;
reg [`NUM_VC - 1 : 0] qibc2e1;
reg [`NUM_VC - 1 : 0] bye1708;
reg [`NUM_VC - 1 : 0] dob843;
reg [`NUM_VC - 1 : 0] cm5c21a;
reg [`NUM_VC - 1 : 0] hoe10d1;
reg [`NUM_VC - 1 : 0] an868b;
reg [`NUM_VC - 1 : 0] kf880d;
reg [`NUM_VC - 1 : 0] mr4406d;
reg [`NUM_VC - 1 : 0] tw2036c;
reg aab3ea1;
reg [13 : 0] ira415d;
reg [13 : 0] hq20aed;
reg [`NUM_VC - 1 : 0] uk576a;
reg [`NUM_VC - 1 : 0] ec2bb50;
reg [`NUM_VC - 1 : 0] fa5da81;
reg [`NUM_VC - 1 : 0] czed40a;
reg [2047:0] necf6c2;
wire [57:0] ld7b613;
`ifdef AER
`endif
`ifdef AER
`endif
`ifdef VC1
`else
`endif
`ifdef AER
`endif
`ifdef AER
`endif
localparam qgdb09f = 58,nrd84f8 = 32'hfdffc68b;
localparam [31:0] thc27c7 = nrd84f8;
localparam mt9f1ff = nrd84f8 & 4'hf;
localparam [11:0] fnc7fe5 = 'h7ff;
wire  [(1 << mt9f1ff)  -1:0] suff972;
reg    [qgdb09f-1:0] cme5c87;
reg [mt9f1ff-1:0] qg721c0 [0:1];
reg [mt9f1ff-1:0] ym8700c;
reg rv38061;
integer jcc030e;
integer vk1872;
`ifdef AER
`endif
`ifdef AER
`endif
`ifdef VC1
`else
`endif
`ifdef AER
`endif
`ifdef AER
`endif
`ifdef AER
`endif
`ifdef AER
`endif
`ifdef VC1
   assign tw8340b = fn45b3b;   assign aa1a05b = vx2d9df;   assign ned02d8  = ho6cefe;
`else
   assign tw8340b = {{`NUM_VC -1{1'b0}},fn45b3b};   assign aa1a05b = {{`NUM_VC -1{1'b0}},vx2d9df};   assign ned02d8  = {{`NUM_VC -1{1'b0}},ho6cefe};
`endif
assign kd54529 = |czed40a;
assign ykfa0d0 = (al65ca0) ? {ir95972, 2'b00} : {2'b00, ir95972};
always @(posedge sys_clk or negedge rst_n) begin   if (rst_n == 1'b0)      rgd0681 <= 14'h0;   else if (aab3ea1)      rgd0681 <= 14'h0;   else      rgd0681 <= hq20aed + 14'h1;
end
assign ofe77fc = (hq20aed == ira415d) ? 1'b1  : 1'b0;
   wjfdce2 qi97de4(            .sys_clk                  (sys_clk),      .rst_n                    (rst_n),      .rib82be               (ofc3f97),      .icc15f2               (ie1fcbc),      .ym1549d                (dmfe5e1),      .zzaa4e9               (gbf2f0b),      .ne5274e              (uk9785c),      .je93a72               (qibc2e1),      .gq9d393              (bye1708),      .pfe9c99             (dob843),      .mr4e4ce                 (cm5c21a),      .ay72675                (hoe10d1),      .do933a9               (an868b),            .lf198b2               (lf198b2),      .yxcc596                 (yxcc596),      .os62cb4                 (os62cb4),      .fp165a1               (fp165a1),      .xyb2d0e                 (xyb2d0e),      .ba96872                 (ba96872),      .hq99d4a               (hq99d4a),      .qgcea52              (qgcea52),      .en75290             (en75290)      );
ep2c61a rv322e4 [`NUM_VC-1:0] (            .sys_clk                  (sys_clk),      .rst_n                    (rst_n),            .ofc3555               (hq83f1a),      .mg1aaad              (ec1f8d2),      .jcd5569             (zxfc691),      .jraab4b               (xje348e),      .vv55a5f              (sw1a476),      .vkad2fe             (dzd23b0),      .lq697f3           (jr91d86),      .kd4bf9b           (fp8ec36),      .jp5fcdc          (tu761b6),      .lqfe6e7          (bnb0db3),      .thf373b         (ls86d9f),      .bn9b9df         (mt36cfa),      .aldceff                  (vv7e6c2),      .ofe77fc              (aab3ea1),      .ym3bfe4               (an9f508),      .jpd27c8              (mefa844),      .do93e46             (uid4220),      .mt9f233            (sja1101),      .hq99d4a               (kf880d),      .qgcea52              (mr4406d),      .en75290             (tw2036c),      .mt18edf            (ri1b63),      .hbc76fc            (mtdb1b),      .ie3b7e7           (ay6d8dd),      .sudbf39           (vi6c6e8),      .fadf9c9          (lq63743),      .hbfce4b          (ba1ba1a),      .mre725f             (bldd0d3),      .kf392fc             (ale869f),      .gbc97e4            (yk434fd),      .cz4bf24            (ou1a7e9),      .xj5f924           (wjd3f48),      .vvfc927           (ir9fa45),      .fp27e80        (uk576a),      .je3f407        (ec2bb50),      .ayfa03b         (fa5da81),      .tue493f                   (enfd22d),      .mg249fa                  (lde916c),      .ie24fd0                 (jc48b67),
`ifdef AER
            .hod01d9                  (hod01d9),      .sj80ecb                  (sj80ecb),      .ux765d                  (ux765d),      .ie3b2ed                 (ie3b2ed),      .uvd9769                 (uvd9769),      .uicbb4d             (uicbb4d),      .jc5da68              (jc5da68),      .iped342              (iped342),      .lq69a15             (lq69a15),      .fa4d0aa             (fa4d0aa),
`endif
            .ym1549d                (ym1549d),      .zzaa4e9               (zzaa4e9),      .ne5274e              (ne5274e),      .je93a72               (je93a72),      .gq9d393              (gq9d393),      .pfe9c99             (pfe9c99),      .mr4e4ce                 (mr4e4ce),      .ay72675                (ay72675),      .do933a9               (do933a9),
      .wlb4393            (wlb4393),      .uxa1c9c           (uxa1c9c),      .vke4e4          (vke4e4),
`ifdef AER
      .zxece0b                 (ph816c3),
`endif
      .me6705e                     (me6705e),      .lf382f0                    (lf382f0),      .mec1786                   (mec1786)
      );
always@* begin hq83f1a<={ofc3555>>1,ld7b613[0]};ec1f8d2<={mg1aaad>>1,ld7b613[1]};zxfc691<={jcd5569>>1,ld7b613[2]};xje348e<={jraab4b>>1,ld7b613[3]};sw1a476<={vv55a5f>>1,ld7b613[4]};dzd23b0<={vkad2fe>>1,ld7b613[5]};jr91d86<={lq697f3>>1,ld7b613[6]};fp8ec36<={kd4bf9b>>1,ld7b613[7]};tu761b6<={jp5fcdc>>1,ld7b613[8]};bnb0db3<={lqfe6e7>>1,ld7b613[9]};ls86d9f<={thf373b>>1,ld7b613[10]};mt36cfa<={bn9b9df>>1,ld7b613[11]};ir95972<={nt8b8a0>>1,ld7b613[12]};vv7e6c2<={ls1e282>>1,ld7b613[13]};al65ca0<=ld7b613[14];an9f508<=ld7b613[15];ofc3f97<=ld7b613[16];ie1fcbc<=ld7b613[17];mefa844<={jpd27c8>>1,ld7b613[18]};uid4220<={do93e46>>1,ld7b613[19]};sja1101<={mt9f233>>1,ld7b613[20]};ri1b63<={mt18edf>>1,ld7b613[21]};mtdb1b<={hbc76fc>>1,ld7b613[22]};ay6d8dd<={ie3b7e7>>1,ld7b613[23]};vi6c6e8<={sudbf39>>1,ld7b613[24]};lq63743<={fadf9c9>>1,ld7b613[25]};ba1ba1a<={hbfce4b>>1,ld7b613[26]};bldd0d3<={mre725f>>1,ld7b613[27]};ale869f<={kf392fc>>1,ld7b613[28]};yk434fd<={gbc97e4>>1,ld7b613[29]};ou1a7e9<={cz4bf24>>1,ld7b613[30]};wjd3f48<={xj5f924>>1,ld7b613[31]};ir9fa45<={vvfc927>>1,ld7b613[32]};fn45b3b<=ld7b613[33];vx2d9df<=ld7b613[34];ho6cefe<=ld7b613[35];enfd22d<={tue493f>>1,ld7b613[36]};lde916c<={mg249fa>>1,ld7b613[37]};jc48b67<={ie24fd0>>1,ld7b613[38]};dmfe5e1<={ym1549d>>1,ld7b613[39]};gbf2f0b<={zzaa4e9>>1,ld7b613[40]};uk9785c<={ne5274e>>1,ld7b613[41]};qibc2e1<={je93a72>>1,ld7b613[42]};bye1708<={gq9d393>>1,ld7b613[43]};dob843<={pfe9c99>>1,ld7b613[44]};cm5c21a<={mr4e4ce>>1,ld7b613[45]};hoe10d1<={ay72675>>1,ld7b613[46]};an868b<={do933a9>>1,ld7b613[47]};kf880d<={hq99d4a>>1,ld7b613[48]};mr4406d<={qgcea52>>1,ld7b613[49]};tw2036c<={en75290>>1,ld7b613[50]};aab3ea1<=ld7b613[51];ira415d<={ykfa0d0>>1,ld7b613[52]};hq20aed<={rgd0681>>1,ld7b613[53]};uk576a<={tw8340b>>1,ld7b613[54]};ec2bb50<={aa1a05b>>1,ld7b613[55]};fa5da81<={ned02d8>>1,ld7b613[56]};czed40a<={ph816c3>>1,ld7b613[57]};end
always@* begin necf6c2[2047]<=mg1aaad[0];necf6c2[2046]<=jcd5569[0];necf6c2[2044]<=jraab4b[0];necf6c2[2040]<=vv55a5f[0];necf6c2[2032]<=vkad2fe[0];necf6c2[2017]<=lq697f3[0];necf6c2[1987]<=kd4bf9b[0];necf6c2[1980]<=qgcea52[0];necf6c2[1963]<=fp27e80;necf6c2[1942]<=tw8340b[0];necf6c2[1926]<=jp5fcdc[0];necf6c2[1921]<=ie3b7e7[0];necf6c2[1913]<=en75290[0];necf6c2[1903]<=je93a72[0];necf6c2[1879]<=je3f407;necf6c2[1837]<=aa1a05b[0];necf6c2[1805]<=lqfe6e7[0];necf6c2[1795]<=sudbf39[0];necf6c2[1783]<=ay72675[0];necf6c2[1778]<=ofe77fc;necf6c2[1758]<=gq9d393[0];necf6c2[1710]<=ayfa03b;necf6c2[1679]<=rib82be;necf6c2[1627]<=ned02d8[0];necf6c2[1562]<=thf373b[0];necf6c2[1543]<=fadf9c9[0];necf6c2[1519]<=do933a9[0];necf6c2[1509]<=ykfa0d0[0];necf6c2[1499]<=zzaa4e9[0];necf6c2[1469]<=pfe9c99[0];necf6c2[1398]<=ie24fd0[0];necf6c2[1373]<=tue493f[0];necf6c2[1310]<=icc15f2;necf6c2[1207]<=ph816c3[0];necf6c2[1144]<=do93e46[0];necf6c2[1076]<=bn9b9df[0];necf6c2[1039]<=hbfce4b[0];necf6c2[1023]<=ofc3555[0];necf6c2[990]<=hq99d4a[0];necf6c2[981]<=vvfc927[0];necf6c2[971]<=rgd0681[0];necf6c2[960]<=hbc76fc[0];necf6c2[951]<=ne5274e[0];necf6c2[891]<=mr4e4ce[0];necf6c2[839]<=ym3bfe4;necf6c2[749]<=ym1549d[0];necf6c2[699]<=mg249fa[0];necf6c2[572]<=jpd27c8[0];necf6c2[490]<=xj5f924[0];necf6c2[480]<=mt18edf[0];necf6c2[419]<=yxe2831;necf6c2[245]<=cz4bf24[0];necf6c2[240]<=mt9f233[0];necf6c2[209]<=ls1e282[0];necf6c2[122]<=gbc97e4[0];necf6c2[104]<=nt8b8a0[0];necf6c2[61]<=kf392fc[0];necf6c2[30]<=mre725f[0];end         assign suff972 = necf6c2,ld7b613 = cme5c87;   initial begin   jcc030e = $fopen(".fred");   $fdisplay( jcc030e, "%3h\n%3h", (thc27c7 >> 4) & fnc7fe5, (thc27c7 >> (mt9f1ff+4)) & fnc7fe5 );   $fclose(jcc030e);   $readmemh(".fred", qg721c0);   end   always @ (suff972) begin   ym8700c = qg721c0[1];       for (vk1872=0; vk1872<qgdb09f; vk1872=vk1872+1) begin           cme5c87[vk1872] = suff972[ym8700c];       rv38061  = ^(ym8700c & qg721c0[0]);       ym8700c =  {ym8700c, rv38061};       end   end
endmodule