module above.
  cf_adc_wr #(.C_CF_BUFTYPE(C_CF_BUFTYPE), .C_IODELAY_GROUP(C_IODELAY_GROUP)) i_adc_wr (
    .adc_clk_in_p (adc_clk_in_p),
    .adc_clk_in_n (adc_clk_in_n),
    .adc_data_in_p (adc_data_in_p),
    .adc_data_in_n (adc_data_in_n),
    .adc_data_or_p (adc_data_or_p),
    .adc_data_or_n (adc_data_or_n),
    .adc_clk (adc_clk),
    .adc_valid (adc_valid_s),
    .adc_data (adc_data_s),
    .adc_or (adc_or_s),
    .adc_pn_oos (adc_pn_oos_s),
    .adc_pn_err (adc_pn_err_s),
    .up_signext_enable (up_signext_enable),
    .up_muladd_enable (up_muladd_enable),
    .up_muladd_offbin (up_muladd_offbin),
    .up_muladd_scale_a (up_muladd_scale_a),
    .up_muladd_offset_a (up_muladd_offset_a),
    .up_muladd_scale_b (up_muladd_scale_b),
    .up_muladd_offset_b (up_muladd_offset_b),
    .up_pn_type (up_pn_type),
    .up_dmode (up_dmode),
    .up_ch_sel (up_ch_sel),
    .up_usr_sel (up_usr_sel),
    .up_delay_sel (up_delay_sel),
    .up_delay_rwn (up_delay_rwn),
    .up_delay_addr (up_delay_addr),
    .up_delay_wdata (up_delay_wdata),
    .up_decimation_m (up_decimation_m),
    .up_decimation_n (up_decimation_n),
    .up_data_type (up_data_type),
    .up_dcfilter_coeff_a (up_dcfilter_coeff_a),
    .up_dcfilter_coeff_b (up_dcfilter_coeff_b),
    .usr_decimation_m (usr_decimation_m_s),
    .usr_decimation_n (usr_decimation_n_s),
    .usr_data_type (usr_data_type_s),
    .usr_max_channels (usr_max_channels_s),
    .delay_clk (delay_clk),
    .delay_ack (delay_ack_s),
    .delay_rdata (delay_rdata_s),
    .delay_locked (delay_locked_s),
    .debug_data (),
    .debug_trigger (),
    .adc_mon_valid (adc_mon_valid),
    .adc_mon_data (adc_mon_data));
endmodule