module header
	// Internal signals
	// Generated Signal List
	// End of Generated Signal List
	// %COMPILER_OPTS%
	// Generated Signal Assignments
	// Generated Instances and Port Mappings
		// Generated Instance Port Map for pad_data9
		IO60DRV1 pad_data9 (
			.pad(data9)	// From TopLevel Boundary
		);
		// End of Generated Instance Port Map for pad_data9
endmodule