module test_pe;
	// Inputs
	reg clk;
	reg reset;
	reg [10:0] ctrl;
	reg [`WIDTH_D0:0] d0;
	reg [`WIDTH:0] d1;
	reg [`WIDTH:0] d2;
    reg [`WIDTH:0] wish;
	// Outputs
	wire [`WIDTH:0] out;
	// Instantiate the Unit Under Test (UUT)
	PE uut (
		.clk(clk),
		.reset(reset),
		.ctrl(ctrl),
		.d0(d0),
		.d1(d1),
        .d2(d2),
		.out(out)
	);
	initial begin
		// Initialize Inputs
		clk = 0;
		reset = 0;
		ctrl = 0;
		d0 = 0;
		d1 = 0;
        d2 = 0;
		// Wait 100 ns for global reset to finish
		#100;
		// Add stimulus here
        // test mult
        d0 = 1186'h245958540550916859984664a9559916599551944415826a8429555562950a5555a9661855015655694448585615852515916545158595955690a96a566591598660556a61880a410615585525454612010662a4a9116906410014611105015955161455804415166155815941116592650115564164556112804292528419450a45840158a926588250411118055565654556964;
        d1 = 1186'h212291922556595445146a555159a2414515699455212899424869242411a459a6a96954461552562556a11694912451a058440646451050819559181a546891566865542169546869551654262068564119555949915194580525869959a159444051555a01a11509919294620158600555158520569556a514684225201a255a586294585262195922250514115a05542946299;
        d2 = d1;
        wish = 1186'h21a0004a5961412a2068488080020408114aa1aa6296a615418a9a22220948905a4a119849a541100016a14141625a21a906a05024001559086584205a1241804215518688468146052485a40581824a1146915164288a904150960222022aa49555608086151504905a68065906122568a2188a22aa09004451464946201a689926105411588591198551a1085145a6846196910;
        @(negedge clk);
        reset=1;#`P reset=0;
        ctrl=11'b11111_000000; #`P;
        ctrl=11'b00000_111111; #(198*`P);
        check;
        // test cubic
        d0 = {6'b10101, 1182'd0};
        d1 = 1186'h198565655595622106a15596a98a5186101959554541466581244585515555665552584505511552650944484555052655692189595619806549462551a56051552069242a6555542014551599866559955466a604511499554654119144668125851211419566a645856592a55865458582952556a916189591194655519664218a5a9a64990415a516a5169865415a912605951;
        d2 = d1;
        wish = 1186'h01a1425a929600890401891a44129844120112246215a566842954a605aaa8aa08588091659481a062a8519a868aa1548569a18a642222490a80aa8026a22501a8492a10555158491155025a84686680984852046a88a1008249008541a550556181952208252029264a0a4151045415450886854129a9658608684901089910281a22a46262a18108451120145a2625904921a96;
        @(negedge clk);
        reset=1;#`P reset=0;
        ctrl=11'b11111_000000; #`P;
        ctrl=1; #(`P);
        check;
        // test add
        d0 = {6'b000101, 1182'd0};
        d1 = 1186'h00a6540512a166a914956a65149495511551891946505601545514458a955815a5596918a2195a565906902549a4954419294a5045199954951561555804612a6655256899454941a51a590259466611545a628496596845046015584a4455a5aa69858911112a9666549561252a156559564966195415951a41226620598145a0441915951185246145aa55615556585564965a5;
        d2 = 1186'h219146612691209655566446a585291504580155555689915a555564404562896415518a65915062459564695665590a11465845a6659441a515a50a656a0a809016195545425645a509895161841616a665599585a0115416a8952185954555564146a56025559466a85a098a68584564969965441822018992901511a954664a90555414555114149641a811854525452a65612;
        wish = 1186'h21449a6605425640692892a88959826619a98a6298a61092a2aa69a90a1a8a9219628a9614aaaa8592980452901922422a609695284261954a2a1650816268aa06680281128490865a1416508a0a49240a808859580949991a18aa4900199a0a01aa08624106406a9900206aa05661aa812916985160049694108248010615a82a146269a966160845182801421a98419a5208884;
        @(negedge clk);
        reset=1;#`P reset=0;
        ctrl=11'b11111_000000; #`P;
        ctrl=11'b10001; #(`P);
        check;
        // test sub
        d0 = {6'b001001, 1182'd0};
        d1 = 1186'h00a6540512a166a914956a65149495511551891946505601545514458a955815a5596918a2195a565906902549a4954419294a5045199954951561555804612a6655256899454941a51a590259466611545a628496596845046015584a4455a5aa69858911112a9666549561252a156559564966195415951a41226620598145a0441915951185246145aa55615556585564965a5;
        d2 = 1186'h219146612691209655566446a585291504580155555689915a555564404562896415518a65915062459564695665590a11465845a6659441a515a50a656a0a809016195545425645a509895161841616a665599585a0115416a8952185954555564146a56025559466a85a098a68584564969965441822018992901511a954664a90555414555114149641a811854525452a65612;
        wish = 1186'h1215119428104616824206226212a8481105888421099960090082114a5029584144185149480a24146168882642484908a6221a92a405162000885a2699666a9642181654062608001190a12882500aa125152211a95a212184406a85a2105054284214a128950200a84a646a8289202580a0019548269451a2525112a0691265a484818188641059a269a950901166104961296;
        @(negedge clk);
        reset=1;#`P reset=0;
        ctrl=11'b11111_000000; #`P;
        ctrl=11'b10001; #(`P);
        check;
        $display("Good!");
        $finish;
	end
    initial #100 forever #(`P/2) clk = ~clk;
    task check;
        begin
          if (out !== wish)
            begin $display("E %h %h", out, wish); $finish; end
        end
    endtask
endmodule