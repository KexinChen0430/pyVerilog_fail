module imp_test_mod;
   import imp_test_pkg::byte_t;
   byte_t some_byte;
endmodule