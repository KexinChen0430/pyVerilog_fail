module outputs)
   wire [31:0]		outp;			// From test of Test.v
   // End of automatics
   Test test (/*AUTOINST*/
	      // Outputs
	      .outp			(outp[31:0]),
	      // Inputs
	      .reset			(reset),
	      .clk			(clk),
	      .inp			(inp[31:0]));
   // Aggregate outputs into a single result vector
   wire [63:0] result = {32'h0, outp};
   // What checksum will we end up with
`define EXPECTED_SUM 64'ha7f0a34f9cf56ccb
   // Test loop
   always @ (posedge clk) begin
`ifdef TEST_VERBOSE
      $write("[%0t] cyc==%0d crc=%x result=%x\n",$time, cyc, crc, result);
`endif
      cyc <= cyc + 1;
      crc <= {crc[62:0], crc[63]^crc[2]^crc[0]};
      sum <= result ^ {sum[62:0],sum[63]^sum[2]^sum[0]};
      if (cyc==0) begin
	 // Setup
	 crc <= 64'h5aef0c8d_d70a4497;
      end
      else if (cyc<10) begin
	 sum <= 64'h0;
      end
      else if (cyc<90) begin
      end
      else if (cyc==99) begin
	 $write("[%0t] cyc==%0d crc=%x sum=%x\n",$time, cyc, crc, sum);
	 if (crc !== 64'hc77bb9b3784ea091) $stop;
	 if (sum !== `EXPECTED_SUM) $stop;
	 $write("*-* All Finished *-*\n");
	 $finish;
      end
   end
endmodule