module FFT (
  aclk, s_axis_config_tvalid, s_axis_data_tvalid, s_axis_data_tlast, s_axis_config_tready, s_axis_data_tready, m_axis_data_tvalid, m_axis_data_tlast,
event_frame_started, event_tlast_unexpected, event_tlast_missing, event_data_in_channel_halt, s_axis_config_tdata, s_axis_data_tdata,
m_axis_data_tdata, m_axis_data_tuser
)/* synthesis syn_black_box syn_noprune=1 */;
  input aclk;
  input s_axis_config_tvalid;
  input s_axis_data_tvalid;
  input s_axis_data_tlast;
  output s_axis_config_tready;
  output s_axis_data_tready;
  output m_axis_data_tvalid;
  output m_axis_data_tlast;
  output event_frame_started;
  output event_tlast_unexpected;
  output event_tlast_missing;
  output event_data_in_channel_halt;
  input [7 : 0] s_axis_config_tdata;
  input [31 : 0] s_axis_data_tdata;
  output [31 : 0] m_axis_data_tdata;
  output [7 : 0] m_axis_data_tuser;
  // synthesis translate_off
  wire \U0/i_synth/axi_wrapper/event_frame_started ;
  wire \U0/i_synth/axi_wrapper/event_tlast_missing ;
  wire \U0/i_synth/axi_wrapper/event_data_in_channel_halt_int ;
  wire sig00000001;
  wire sig00000002;
  wire sig00000003;
  wire sig00000004;
  wire sig00000005;
  wire sig00000006;
  wire sig00000007;
  wire sig00000008;
  wire sig00000009;
  wire sig0000000a;
  wire sig0000000b;
  wire sig0000000c;
  wire sig0000000d;
  wire sig0000000e;
  wire sig0000000f;
  wire sig00000010;
  wire sig00000011;
  wire sig00000012;
  wire sig00000013;
  wire sig00000014;
  wire sig00000015;
  wire sig00000016;
  wire sig00000017;
  wire sig00000018;
  wire sig00000019;
  wire sig0000001a;
  wire sig0000001b;
  wire sig0000001c;
  wire sig0000001d;
  wire sig0000001e;
  wire sig0000001f;
  wire sig00000020;
  wire sig00000021;
  wire sig00000022;
  wire sig00000023;
  wire sig00000024;
  wire sig00000025;
  wire sig00000026;
  wire sig00000027;
  wire sig00000028;
  wire sig00000029;
  wire sig0000002a;
  wire sig0000002b;
  wire sig0000002c;
  wire sig0000002d;
  wire sig0000002e;
  wire sig0000002f;
  wire sig00000030;
  wire sig00000031;
  wire sig00000032;
  wire sig00000033;
  wire sig00000034;
  wire sig00000035;
  wire sig00000036;
  wire sig00000037;
  wire sig00000038;
  wire sig00000039;
  wire sig0000003a;
  wire sig0000003b;
  wire sig0000003c;
  wire sig0000003d;
  wire sig0000003e;
  wire sig0000003f;
  wire sig00000040;
  wire sig00000041;
  wire sig00000042;
  wire sig00000043;
  wire sig00000044;
  wire sig00000045;
  wire sig00000046;
  wire sig00000047;
  wire sig00000048;
  wire sig00000049;
  wire sig0000004a;
  wire sig0000004b;
  wire sig0000004c;
  wire sig0000004d;
  wire sig0000004e;
  wire sig0000004f;
  wire sig00000050;
  wire sig00000051;
  wire sig00000052;
  wire sig00000053;
  wire sig00000054;
  wire sig00000055;
  wire sig00000056;
  wire sig00000057;
  wire sig00000058;
  wire sig00000059;
  wire sig0000005a;
  wire sig0000005b;
  wire sig0000005c;
  wire sig0000005d;
  wire sig0000005e;
  wire sig0000005f;
  wire sig00000060;
  wire sig00000061;
  wire sig00000062;
  wire sig00000063;
  wire sig00000064;
  wire sig00000065;
  wire sig00000066;
  wire sig00000067;
  wire sig00000068;
  wire \NlwRenamedSig_OI_U0/i_synth/axi_wrapper/dv_resolved_prev ;
  wire sig00000069;
  wire sig0000006a;
  wire sig0000006b;
  wire sig0000006c;
  wire sig0000006d;
  wire sig0000006e;
  wire sig0000006f;
  wire sig00000070;
  wire sig00000071;
  wire sig00000072;
  wire sig00000073;
  wire sig00000074;
  wire sig00000075;
  wire sig00000076;
  wire sig00000077;
  wire sig00000078;
  wire sig00000079;
  wire sig0000007a;
  wire sig0000007b;
  wire sig0000007c;
  wire sig0000007d;
  wire sig0000007e;
  wire sig0000007f;
  wire sig00000080;
  wire sig00000081;
  wire sig00000082;
  wire sig00000083;
  wire sig00000084;
  wire sig00000085;
  wire sig00000086;
  wire sig00000087;
  wire sig00000088;
  wire sig00000089;
  wire sig0000008a;
  wire sig0000008b;
  wire sig0000008c;
  wire sig0000008d;
  wire sig0000008e;
  wire sig0000008f;
  wire sig00000090;
  wire sig00000091;
  wire sig00000092;
  wire sig00000093;
  wire sig00000094;
  wire sig00000095;
  wire sig00000096;
  wire sig00000097;
  wire sig00000098;
  wire sig00000099;
  wire sig0000009a;
  wire sig0000009b;
  wire sig0000009c;
  wire sig0000009d;
  wire sig0000009e;
  wire sig0000009f;
  wire sig000000a0;
  wire sig000000a1;
  wire sig000000a2;
  wire sig000000a3;
  wire sig000000a4;
  wire sig000000a5;
  wire sig000000a6;
  wire sig000000a7;
  wire sig000000a8;
  wire sig000000a9;
  wire sig000000aa;
  wire sig000000ab;
  wire sig000000ac;
  wire sig000000ad;
  wire sig000000ae;
  wire sig000000af;
  wire sig000000b0;
  wire sig000000b1;
  wire sig000000b2;
  wire sig000000b3;
  wire sig000000b4;
  wire sig000000b5;
  wire sig000000b6;
  wire sig000000b7;
  wire sig000000b8;
  wire sig000000b9;
  wire sig000000ba;
  wire sig000000bb;
  wire sig000000bc;
  wire sig000000bd;
  wire sig000000be;
  wire sig000000bf;
  wire sig000000c0;
  wire sig000000c1;
  wire sig000000c2;
  wire sig000000c3;
  wire sig000000c4;
  wire sig000000c5;
  wire sig000000c6;
  wire sig000000c7;
  wire sig000000c8;
  wire sig000000c9;
  wire sig000000ca;
  wire sig000000cb;
  wire sig000000cc;
  wire sig000000cd;
  wire sig000000ce;
  wire sig000000cf;
  wire sig000000d0;
  wire sig000000d1;
  wire sig000000d2;
  wire sig000000d3;
  wire sig000000d4;
  wire sig000000d5;
  wire sig000000d6;
  wire sig000000d7;
  wire sig000000d8;
  wire sig000000d9;
  wire sig000000da;
  wire sig000000db;
  wire sig000000dc;
  wire sig000000dd;
  wire sig000000de;
  wire sig000000df;
  wire sig000000e0;
  wire sig000000e1;
  wire sig000000e2;
  wire sig000000e3;
  wire sig000000e4;
  wire sig000000e5;
  wire sig000000e6;
  wire sig000000e7;
  wire sig000000e8;
  wire sig000000e9;
  wire sig000000ea;
  wire sig000000eb;
  wire sig000000ec;
  wire sig000000ed;
  wire sig000000ee;
  wire sig000000ef;
  wire sig000000f0;
  wire sig000000f1;
  wire sig000000f2;
  wire sig000000f3;
  wire sig000000f4;
  wire sig000000f5;
  wire sig000000f6;
  wire sig000000f7;
  wire sig000000f8;
  wire sig000000f9;
  wire sig000000fa;
  wire sig000000fb;
  wire sig000000fc;
  wire sig000000fd;
  wire sig000000fe;
  wire sig000000ff;
  wire sig00000100;
  wire sig00000101;
  wire sig00000102;
  wire sig00000103;
  wire sig00000104;
  wire sig00000105;
  wire sig00000106;
  wire sig00000107;
  wire sig00000108;
  wire sig00000109;
  wire sig0000010a;
  wire sig0000010b;
  wire sig0000010c;
  wire sig0000010d;
  wire sig0000010e;
  wire sig0000010f;
  wire sig00000110;
  wire sig00000111;
  wire sig00000112;
  wire sig00000113;
  wire sig00000114;
  wire sig00000115;
  wire sig00000116;
  wire sig00000117;
  wire sig00000118;
  wire sig00000119;
  wire sig0000011a;
  wire sig0000011b;
  wire sig0000011c;
  wire sig0000011d;
  wire sig0000011e;
  wire sig0000011f;
  wire sig00000120;
  wire sig00000121;
  wire sig00000122;
  wire sig00000123;
  wire sig00000124;
  wire sig00000125;
  wire sig00000126;
  wire sig00000127;
  wire sig00000128;
  wire sig00000129;
  wire sig0000012a;
  wire sig0000012b;
  wire sig0000012c;
  wire sig0000012d;
  wire sig0000012e;
  wire sig0000012f;
  wire sig00000130;
  wire sig00000131;
  wire sig00000132;
  wire sig00000133;
  wire sig00000134;
  wire sig00000135;
  wire sig00000136;
  wire sig00000137;
  wire sig00000138;
  wire sig00000139;
  wire sig0000013a;
  wire sig0000013b;
  wire sig0000013c;
  wire sig0000013d;
  wire sig0000013e;
  wire sig0000013f;
  wire sig00000140;
  wire sig00000141;
  wire sig00000142;
  wire sig00000143;
  wire sig00000144;
  wire sig00000145;
  wire sig00000146;
  wire sig00000147;
  wire sig00000148;
  wire sig00000149;
  wire sig0000014a;
  wire sig0000014b;
  wire sig0000014c;
  wire sig0000014d;
  wire sig0000014e;
  wire sig0000014f;
  wire sig00000150;
  wire sig00000151;
  wire sig00000152;
  wire sig00000153;
  wire sig00000154;
  wire sig00000155;
  wire sig00000156;
  wire sig00000157;
  wire sig00000158;
  wire sig00000159;
  wire sig0000015a;
  wire sig0000015b;
  wire sig0000015c;
  wire sig0000015d;
  wire sig0000015e;
  wire sig0000015f;
  wire sig00000160;
  wire sig00000161;
  wire sig00000162;
  wire sig00000163;
  wire sig00000164;
  wire sig00000165;
  wire sig00000166;
  wire sig00000167;
  wire sig00000168;
  wire sig00000169;
  wire sig0000016a;
  wire sig0000016b;
  wire sig0000016c;
  wire sig0000016d;
  wire sig0000016e;
  wire sig0000016f;
  wire sig00000170;
  wire sig00000171;
  wire sig00000172;
  wire sig00000173;
  wire sig00000174;
  wire sig00000175;
  wire sig00000176;
  wire sig00000177;
  wire sig00000178;
  wire sig00000179;
  wire sig0000017a;
  wire sig0000017b;
  wire sig0000017c;
  wire sig0000017d;
  wire sig0000017e;
  wire sig0000017f;
  wire sig00000180;
  wire sig00000181;
  wire sig00000182;
  wire sig00000183;
  wire sig00000184;
  wire sig00000185;
  wire sig00000186;
  wire sig00000187;
  wire sig00000188;
  wire sig00000189;
  wire sig0000018a;
  wire sig0000018b;
  wire sig0000018c;
  wire sig0000018d;
  wire sig0000018e;
  wire sig0000018f;
  wire sig00000190;
  wire sig00000191;
  wire sig00000192;
  wire sig00000193;
  wire sig00000194;
  wire sig00000198;
  wire sig00000199;
  wire sig0000019b;
  wire sig0000019c;
  wire sig0000019d;
  wire sig000001a0;
  wire sig000001ae;
  wire sig000001af;
  wire sig000001b0;
  wire sig000001b1;
  wire sig000001b2;
  wire sig000001b3;
  wire sig000001b4;
  wire sig000001b5;
  wire sig000001b6;
  wire sig000001b7;
  wire sig000001b8;
  wire sig000001b9;
  wire sig000001ba;
  wire sig000001bb;
  wire sig000001bc;
  wire sig000001bd;
  wire sig000001be;
  wire sig000001bf;
  wire sig000001c0;
  wire sig000001c1;
  wire sig000001c2;
  wire sig000001c3;
  wire sig000001c4;
  wire sig000001c5;
  wire sig000001c6;
  wire sig000001c7;
  wire sig000001c8;
  wire sig000001c9;
  wire sig000001ca;
  wire sig000001cb;
  wire sig000001cc;
  wire sig000001cd;
  wire sig000001ce;
  wire sig000001cf;
  wire sig000001d0;
  wire sig000001d1;
  wire sig000001d2;
  wire sig000001d3;
  wire sig000001d4;
  wire sig000001d5;
  wire sig000001d6;
  wire sig000001d7;
  wire sig000001d8;
  wire sig000001d9;
  wire sig000001da;
  wire sig000001db;
  wire sig000001dc;
  wire sig000001dd;
  wire sig000001de;
  wire sig000001df;
  wire sig000001e0;
  wire sig000001e1;
  wire sig000001e2;
  wire sig000001e3;
  wire sig000001e4;
  wire sig000001e5;
  wire sig000001e6;
  wire sig000001e7;
  wire sig000001e8;
  wire sig000001e9;
  wire sig000001ea;
  wire sig000001eb;
  wire sig000001ec;
  wire sig000001ed;
  wire sig000001ee;
  wire sig000001ef;
  wire sig000001f0;
  wire sig000001f1;
  wire sig000001f2;
  wire sig000001f3;
  wire sig000001f4;
  wire sig000001f5;
  wire sig000001f6;
  wire sig000001f7;
  wire sig000001f8;
  wire sig000001f9;
  wire sig000001fa;
  wire sig000001fb;
  wire sig000001fc;
  wire sig000001fd;
  wire sig000001fe;
  wire sig000001ff;
  wire sig00000200;
  wire sig00000201;
  wire sig00000202;
  wire sig00000203;
  wire sig00000204;
  wire sig00000205;
  wire sig00000206;
  wire sig00000207;
  wire sig00000208;
  wire sig00000209;
  wire sig0000020a;
  wire sig0000020b;
  wire sig0000020c;
  wire sig0000020d;
  wire sig0000020e;
  wire sig0000020f;
  wire sig00000210;
  wire sig00000211;
  wire sig00000212;
  wire sig00000213;
  wire sig00000214;
  wire sig00000215;
  wire sig00000216;
  wire sig00000217;
  wire sig00000218;
  wire sig00000219;
  wire sig0000021a;
  wire sig0000021b;
  wire sig0000021c;
  wire sig0000021d;
  wire sig0000021e;
  wire sig0000021f;
  wire sig00000220;
  wire sig00000221;
  wire sig00000222;
  wire sig00000223;
  wire sig00000224;
  wire sig00000225;
  wire sig00000226;
  wire sig00000227;
  wire sig00000228;
  wire sig00000229;
  wire sig0000022a;
  wire sig0000022b;
  wire sig0000022c;
  wire sig0000022d;
  wire sig0000022e;
  wire sig0000022f;
  wire sig00000230;
  wire sig00000231;
  wire sig00000232;
  wire sig00000233;
  wire sig00000234;
  wire sig00000235;
  wire sig00000236;
  wire sig00000237;
  wire sig00000238;
  wire sig00000239;
  wire sig0000023a;
  wire sig0000023b;
  wire sig0000023c;
  wire sig0000023d;
  wire sig0000023e;
  wire sig0000023f;
  wire sig00000240;
  wire sig00000241;
  wire sig00000242;
  wire sig00000243;
  wire sig00000244;
  wire sig00000245;
  wire sig00000246;
  wire sig00000247;
  wire sig00000248;
  wire sig00000249;
  wire sig0000024a;
  wire sig0000024b;
  wire sig0000024c;
  wire sig0000024d;
  wire sig0000024e;
  wire sig0000024f;
  wire sig00000250;
  wire sig00000251;
  wire sig00000252;
  wire sig00000253;
  wire sig00000254;
  wire sig00000255;
  wire sig00000256;
  wire sig00000257;
  wire sig00000258;
  wire sig00000259;
  wire sig0000025a;
  wire sig0000025b;
  wire sig0000025c;
  wire sig0000025d;
  wire sig0000025e;
  wire sig0000025f;
  wire sig00000260;
  wire sig00000261;
  wire sig00000262;
  wire sig00000263;
  wire sig00000264;
  wire sig00000265;
  wire sig00000266;
  wire sig00000267;
  wire sig00000268;
  wire sig00000269;
  wire sig0000026a;
  wire sig0000026b;
  wire sig0000026c;
  wire sig0000026d;
  wire sig0000026e;
  wire sig0000026f;
  wire sig00000270;
  wire sig00000271;
  wire sig00000272;
  wire sig00000273;
  wire sig00000274;
  wire sig00000275;
  wire sig00000276;
  wire sig00000277;
  wire sig00000278;
  wire sig00000279;
  wire sig0000027a;
  wire sig0000027b;
  wire sig0000027c;
  wire sig0000027d;
  wire sig0000027e;
  wire sig0000027f;
  wire sig00000280;
  wire sig00000281;
  wire sig00000282;
  wire sig00000283;
  wire sig00000284;
  wire sig00000285;
  wire sig00000286;
  wire sig00000287;
  wire sig00000288;
  wire sig00000289;
  wire sig0000028a;
  wire sig0000028b;
  wire sig0000028c;
  wire sig0000028d;
  wire sig0000028e;
  wire sig0000028f;
  wire sig00000290;
  wire sig00000291;
  wire sig00000292;
  wire sig00000293;
  wire sig00000294;
  wire sig00000295;
  wire sig00000296;
  wire sig00000297;
  wire sig00000298;
  wire sig00000299;
  wire sig0000029a;
  wire sig0000029b;
  wire sig0000029c;
  wire sig0000029d;
  wire sig0000029e;
  wire sig0000029f;
  wire sig000002a0;
  wire sig000002a1;
  wire sig000002a2;
  wire sig000002a3;
  wire sig000002a4;
  wire sig000002a5;
  wire sig000002a6;
  wire sig000002a7;
  wire sig000002a8;
  wire sig000002a9;
  wire sig000002aa;
  wire sig000002ab;
  wire sig000002ac;
  wire sig000002ad;
  wire sig000002ae;
  wire sig000002af;
  wire sig000002b0;
  wire sig000002b1;
  wire sig000002b2;
  wire sig000002b3;
  wire sig000002b4;
  wire sig000002b5;
  wire sig000002b6;
  wire sig000002b7;
  wire sig000002b8;
  wire sig000002b9;
  wire sig000002ba;
  wire sig000002bb;
  wire sig000002bc;
  wire sig000002bd;
  wire sig000002be;
  wire sig000002bf;
  wire sig000002c0;
  wire sig000002c1;
  wire sig000002c2;
  wire sig000002c3;
  wire sig000002c4;
  wire sig000002c5;
  wire sig000002c6;
  wire sig000002c7;
  wire sig000002c8;
  wire sig000002c9;
  wire sig000002ca;
  wire sig000002cb;
  wire sig000002cc;
  wire sig000002cd;
  wire sig000002ce;
  wire sig000002cf;
  wire sig000002d0;
  wire sig000002d1;
  wire sig000002d2;
  wire sig000002d3;
  wire sig000002d4;
  wire sig000002d5;
  wire sig000002d6;
  wire sig000002d7;
  wire sig000002d8;
  wire sig000002d9;
  wire sig000002da;
  wire sig000002db;
  wire sig000002dc;
  wire sig000002dd;
  wire sig000002de;
  wire sig000002df;
  wire sig000002e0;
  wire sig000002e1;
  wire sig000002e2;
  wire sig000002e3;
  wire sig000002e4;
  wire sig000002e5;
  wire sig000002e6;
  wire sig000002e7;
  wire sig000002e8;
  wire sig000002e9;
  wire sig000002ea;
  wire sig000002eb;
  wire sig000002ec;
  wire sig000002ed;
  wire sig000002ee;
  wire sig000002ef;
  wire sig000002f0;
  wire sig000002f1;
  wire sig000002f2;
  wire sig000002f3;
  wire sig000002f4;
  wire sig000002f5;
  wire sig000002f6;
  wire sig000002f7;
  wire sig000002f8;
  wire sig000002f9;
  wire sig000002fa;
  wire sig000002fb;
  wire sig000002fc;
  wire sig000002fd;
  wire sig000002fe;
  wire sig000002ff;
  wire sig00000300;
  wire sig00000301;
  wire sig00000302;
  wire sig00000303;
  wire sig00000304;
  wire sig00000305;
  wire sig00000306;
  wire sig00000307;
  wire sig00000308;
  wire sig00000309;
  wire sig0000030a;
  wire sig0000030b;
  wire sig0000030c;
  wire sig0000030d;
  wire sig0000030e;
  wire sig0000030f;
  wire sig00000310;
  wire sig00000311;
  wire sig00000312;
  wire sig00000313;
  wire sig00000314;
  wire sig00000315;
  wire sig00000316;
  wire sig00000317;
  wire sig00000318;
  wire sig00000319;
  wire sig0000031a;
  wire sig0000031b;
  wire sig0000031c;
  wire sig0000031d;
  wire sig0000031e;
  wire sig0000031f;
  wire sig00000320;
  wire sig00000321;
  wire sig00000322;
  wire sig00000323;
  wire sig00000324;
  wire sig00000325;
  wire sig00000326;
  wire sig00000327;
  wire sig00000328;
  wire sig00000329;
  wire sig0000032a;
  wire sig0000032b;
  wire sig0000032c;
  wire sig0000032d;
  wire sig0000032e;
  wire sig0000032f;
  wire sig00000330;
  wire sig00000331;
  wire sig00000332;
  wire sig00000333;
  wire sig00000334;
  wire sig00000335;
  wire sig00000336;
  wire sig00000337;
  wire sig00000338;
  wire sig00000339;
  wire sig0000033a;
  wire sig0000033b;
  wire sig0000033c;
  wire sig0000033d;
  wire sig0000033e;
  wire sig0000033f;
  wire sig00000340;
  wire sig00000341;
  wire sig00000342;
  wire sig00000343;
  wire sig00000344;
  wire sig00000345;
  wire sig00000346;
  wire sig00000347;
  wire sig00000348;
  wire sig00000349;
  wire sig0000034a;
  wire sig0000034b;
  wire sig0000034c;
  wire sig0000034d;
  wire sig0000034e;
  wire sig0000034f;
  wire sig00000350;
  wire sig00000351;
  wire sig00000352;
  wire sig00000353;
  wire sig00000354;
  wire sig00000355;
  wire sig00000356;
  wire sig00000357;
  wire sig00000358;
  wire sig00000359;
  wire sig0000035a;
  wire sig0000035b;
  wire sig0000035c;
  wire sig0000035d;
  wire sig0000035e;
  wire sig0000035f;
  wire sig00000360;
  wire sig00000361;
  wire sig00000362;
  wire sig00000363;
  wire sig00000364;
  wire sig00000365;
  wire sig00000366;
  wire sig00000367;
  wire sig00000368;
  wire sig00000369;
  wire sig0000036a;
  wire sig0000036b;
  wire sig0000036c;
  wire sig0000036d;
  wire sig0000036e;
  wire sig0000036f;
  wire sig00000370;
  wire sig00000371;
  wire sig00000372;
  wire sig00000373;
  wire sig00000374;
  wire sig00000375;
  wire sig00000376;
  wire sig00000377;
  wire sig00000378;
  wire sig00000379;
  wire sig0000037a;
  wire sig0000037b;
  wire sig0000037c;
  wire sig0000037d;
  wire sig0000037e;
  wire sig0000037f;
  wire sig00000380;
  wire sig00000381;
  wire sig00000382;
  wire sig00000383;
  wire sig00000384;
  wire sig00000385;
  wire sig00000386;
  wire sig00000387;
  wire sig00000388;
  wire sig00000389;
  wire sig0000038a;
  wire sig0000038b;
  wire sig0000038c;
  wire sig0000038d;
  wire sig0000038e;
  wire sig0000038f;
  wire sig00000390;
  wire sig00000391;
  wire sig00000392;
  wire sig00000393;
  wire sig00000394;
  wire sig00000395;
  wire sig00000396;
  wire sig00000397;
  wire sig00000398;
  wire sig00000399;
  wire sig0000039a;
  wire sig0000039b;
  wire sig0000039c;
  wire sig0000039d;
  wire sig0000039e;
  wire sig0000039f;
  wire sig000003a0;
  wire sig000003a1;
  wire sig000003a2;
  wire sig000003a3;
  wire sig000003a4;
  wire sig000003a5;
  wire sig000003a6;
  wire sig000003a7;
  wire sig000003a8;
  wire sig000003a9;
  wire sig000003aa;
  wire sig000003ab;
  wire sig000003ac;
  wire sig000003ad;
  wire sig000003ae;
  wire sig000003af;
  wire sig000003b0;
  wire sig000003b1;
  wire sig000003b2;
  wire sig000003b3;
  wire sig000003b4;
  wire sig000003b5;
  wire sig000003b6;
  wire sig000003b7;
  wire sig000003b8;
  wire sig000003b9;
  wire sig000003ba;
  wire sig000003bb;
  wire sig000003bc;
  wire sig000003bd;
  wire sig000003be;
  wire sig000003bf;
  wire sig000003c0;
  wire sig000003c1;
  wire sig000003c2;
  wire sig000003c3;
  wire sig000003c4;
  wire sig000003c5;
  wire sig000003c6;
  wire sig000003c7;
  wire sig000003c8;
  wire sig000003c9;
  wire sig000003ca;
  wire sig000003cb;
  wire sig000003cc;
  wire sig000003cd;
  wire sig000003ce;
  wire sig000003cf;
  wire sig000003d0;
  wire sig000003d1;
  wire sig000003d2;
  wire sig000003d3;
  wire sig000003d4;
  wire sig000003d5;
  wire sig000003d6;
  wire sig000003d7;
  wire sig000003d8;
  wire sig000003d9;
  wire sig000003da;
  wire sig000003db;
  wire sig000003dc;
  wire sig000003dd;
  wire sig000003de;
  wire sig000003df;
  wire sig000003e0;
  wire sig000003e1;
  wire sig000003e2;
  wire sig000003e3;
  wire sig000003e4;
  wire sig000003e5;
  wire sig000003e6;
  wire sig000003e7;
  wire sig000003e8;
  wire sig000003e9;
  wire sig000003ea;
  wire sig000003eb;
  wire sig000003ec;
  wire sig000003ed;
  wire sig000003ee;
  wire sig000003ef;
  wire sig000003f0;
  wire sig000003f1;
  wire sig000003f2;
  wire sig000003f3;
  wire sig000003f4;
  wire sig000003f5;
  wire sig000003f6;
  wire sig000003f7;
  wire sig000003f8;
  wire sig000003f9;
  wire sig000003fa;
  wire sig000003fb;
  wire sig000003fc;
  wire sig000003fd;
  wire sig000003fe;
  wire sig000003ff;
  wire sig00000400;
  wire sig00000401;
  wire sig00000402;
  wire sig00000403;
  wire sig00000404;
  wire sig00000405;
  wire sig00000406;
  wire sig00000407;
  wire sig00000408;
  wire sig00000409;
  wire sig0000040a;
  wire sig0000040b;
  wire sig0000040c;
  wire sig0000040d;
  wire sig0000040e;
  wire sig0000040f;
  wire sig00000410;
  wire sig00000411;
  wire sig00000412;
  wire sig00000413;
  wire sig00000414;
  wire sig00000415;
  wire sig00000416;
  wire sig00000417;
  wire sig00000418;
  wire sig00000419;
  wire sig0000041a;
  wire sig0000041b;
  wire sig0000041c;
  wire sig0000041d;
  wire sig0000041e;
  wire sig0000041f;
  wire sig00000420;
  wire sig00000421;
  wire sig00000422;
  wire sig00000423;
  wire sig00000424;
  wire sig00000425;
  wire sig00000426;
  wire sig00000427;
  wire sig00000428;
  wire sig00000429;
  wire sig0000042a;
  wire sig0000042b;
  wire sig0000042c;
  wire sig0000042d;
  wire sig0000042e;
  wire sig0000042f;
  wire sig00000430;
  wire sig00000431;
  wire sig00000432;
  wire sig00000433;
  wire sig00000434;
  wire sig00000435;
  wire sig00000436;
  wire sig00000437;
  wire sig00000438;
  wire sig00000439;
  wire sig0000043a;
  wire sig0000043b;
  wire sig0000043c;
  wire sig0000043d;
  wire sig0000043e;
  wire sig0000043f;
  wire sig00000440;
  wire sig00000441;
  wire sig00000442;
  wire sig00000443;
  wire sig00000444;
  wire sig00000445;
  wire sig00000446;
  wire sig00000447;
  wire sig00000448;
  wire sig00000449;
  wire sig0000044a;
  wire sig0000044b;
  wire sig0000044c;
  wire sig0000044d;
  wire sig0000044e;
  wire sig0000044f;
  wire sig00000450;
  wire sig00000451;
  wire sig00000452;
  wire sig00000453;
  wire sig00000454;
  wire sig00000455;
  wire sig00000456;
  wire sig00000457;
  wire sig00000458;
  wire sig00000459;
  wire sig0000045a;
  wire sig0000045b;
  wire sig0000045c;
  wire sig0000045d;
  wire sig0000045e;
  wire sig0000045f;
  wire sig00000460;
  wire sig00000461;
  wire sig00000462;
  wire sig00000463;
  wire sig00000464;
  wire sig00000465;
  wire sig00000466;
  wire sig00000467;
  wire sig00000468;
  wire sig00000469;
  wire sig0000046a;
  wire sig0000046b;
  wire sig0000046c;
  wire sig0000046d;
  wire sig0000046e;
  wire sig0000046f;
  wire sig00000470;
  wire sig00000471;
  wire sig00000472;
  wire sig00000473;
  wire sig00000474;
  wire sig00000475;
  wire sig00000476;
  wire sig00000477;
  wire sig00000478;
  wire sig00000479;
  wire sig0000047a;
  wire sig0000047b;
  wire sig0000047c;
  wire sig0000047d;
  wire sig0000047e;
  wire sig0000047f;
  wire sig00000480;
  wire sig00000481;
  wire sig00000482;
  wire sig00000483;
  wire sig00000484;
  wire sig00000485;
  wire sig00000486;
  wire sig00000487;
  wire sig00000488;
  wire sig00000489;
  wire sig0000048a;
  wire sig0000048b;
  wire sig0000048c;
  wire sig0000048d;
  wire sig0000048e;
  wire sig0000048f;
  wire sig00000490;
  wire sig00000491;
  wire sig00000492;
  wire sig00000493;
  wire sig00000494;
  wire sig00000495;
  wire sig00000496;
  wire sig00000497;
  wire sig00000498;
  wire sig00000499;
  wire sig0000049a;
  wire sig0000049b;
  wire sig0000049c;
  wire sig0000049d;
  wire sig0000049e;
  wire sig0000049f;
  wire sig000004a0;
  wire sig000004a1;
  wire sig000004a2;
  wire sig000004a3;
  wire sig000004a4;
  wire sig000004a5;
  wire sig000004a6;
  wire sig000004a7;
  wire sig000004a8;
  wire sig000004a9;
  wire sig000004aa;
  wire sig000004ab;
  wire sig000004ac;
  wire sig000004ad;
  wire sig000004ae;
  wire sig000004af;
  wire sig000004b0;
  wire sig000004b1;
  wire sig000004b2;
  wire sig000004b3;
  wire sig000004b4;
  wire sig000004b5;
  wire sig000004b6;
  wire sig000004b7;
  wire sig000004b8;
  wire sig000004b9;
  wire sig000004ba;
  wire sig000004bb;
  wire sig000004bc;
  wire sig000004bd;
  wire sig000004be;
  wire sig000004bf;
  wire sig000004c0;
  wire sig000004c1;
  wire sig000004c2;
  wire sig000004c3;
  wire sig000004c4;
  wire sig000004c5;
  wire sig000004c6;
  wire sig000004c7;
  wire sig000004c8;
  wire sig000004c9;
  wire sig000004ca;
  wire sig000004cb;
  wire sig000004cc;
  wire sig000004cd;
  wire sig000004ce;
  wire sig000004cf;
  wire sig000004d0;
  wire sig000004d1;
  wire sig000004d2;
  wire sig000004d3;
  wire sig000004d4;
  wire sig000004d5;
  wire sig000004d6;
  wire sig000004d7;
  wire sig000004d8;
  wire sig000004d9;
  wire sig000004da;
  wire sig000004db;
  wire sig000004dc;
  wire sig000004dd;
  wire sig000004de;
  wire sig000004df;
  wire sig000004e0;
  wire sig000004e1;
  wire sig000004e2;
  wire sig000004e3;
  wire sig000004e4;
  wire sig000004e5;
  wire sig000004e6;
  wire sig000004e7;
  wire sig000004e8;
  wire sig000004e9;
  wire sig000004ea;
  wire sig000004eb;
  wire sig000004ec;
  wire sig000004ed;
  wire sig000004ee;
  wire sig000004ef;
  wire sig000004f0;
  wire sig000004f1;
  wire sig000004f2;
  wire sig000004f3;
  wire sig000004f4;
  wire sig000004f5;
  wire sig000004f6;
  wire sig000004f7;
  wire sig000004f8;
  wire sig000004f9;
  wire sig000004fa;
  wire sig000004fb;
  wire sig000004fc;
  wire sig000004fd;
  wire sig000004fe;
  wire sig000004ff;
  wire sig00000500;
  wire sig00000501;
  wire sig00000502;
  wire sig00000503;
  wire sig00000504;
  wire sig00000505;
  wire sig00000506;
  wire sig00000507;
  wire sig00000508;
  wire sig00000509;
  wire sig0000050a;
  wire sig0000050b;
  wire sig0000050c;
  wire sig0000050d;
  wire sig0000050e;
  wire sig0000050f;
  wire sig00000510;
  wire sig00000511;
  wire sig00000512;
  wire sig00000513;
  wire sig00000514;
  wire sig00000515;
  wire sig00000516;
  wire sig00000517;
  wire sig00000518;
  wire sig00000519;
  wire sig0000051a;
  wire sig0000051b;
  wire sig0000051c;
  wire sig0000051d;
  wire sig0000051e;
  wire sig0000051f;
  wire sig00000520;
  wire sig00000521;
  wire sig00000522;
  wire sig00000523;
  wire sig00000524;
  wire sig00000525;
  wire sig00000526;
  wire sig00000527;
  wire sig00000528;
  wire sig00000529;
  wire sig0000052a;
  wire sig0000052b;
  wire sig0000052c;
  wire sig0000052d;
  wire sig0000052e;
  wire sig0000052f;
  wire sig00000530;
  wire sig00000531;
  wire sig00000532;
  wire sig00000533;
  wire sig00000534;
  wire sig00000535;
  wire sig00000536;
  wire sig00000537;
  wire sig00000538;
  wire sig00000539;
  wire sig0000053a;
  wire sig0000053b;
  wire sig0000053c;
  wire sig0000053d;
  wire sig0000053e;
  wire sig0000053f;
  wire sig00000540;
  wire sig00000541;
  wire sig00000542;
  wire sig00000543;
  wire sig00000544;
  wire sig00000545;
  wire sig00000546;
  wire sig00000547;
  wire sig00000548;
  wire sig00000549;
  wire sig0000054a;
  wire sig0000054b;
  wire sig0000054c;
  wire sig0000054d;
  wire sig0000054e;
  wire sig0000054f;
  wire sig00000550;
  wire sig00000551;
  wire sig00000552;
  wire sig00000553;
  wire sig00000554;
  wire sig00000555;
  wire sig00000556;
  wire sig00000557;
  wire sig00000558;
  wire sig00000559;
  wire sig0000055a;
  wire sig0000055b;
  wire sig0000055c;
  wire sig0000055d;
  wire sig0000055e;
  wire sig0000055f;
  wire sig00000560;
  wire sig00000561;
  wire sig00000562;
  wire sig00000563;
  wire sig00000564;
  wire sig00000565;
  wire sig00000566;
  wire sig00000567;
  wire sig00000568;
  wire sig00000569;
  wire sig0000056a;
  wire sig0000056b;
  wire sig0000056c;
  wire sig0000056d;
  wire sig0000056e;
  wire sig0000056f;
  wire sig00000570;
  wire sig00000571;
  wire sig00000572;
  wire sig00000573;
  wire sig00000574;
  wire sig00000575;
  wire sig00000576;
  wire sig00000577;
  wire sig00000578;
  wire sig00000579;
  wire sig0000057a;
  wire sig0000057b;
  wire sig0000057c;
  wire sig0000057d;
  wire sig0000057e;
  wire sig0000057f;
  wire sig00000580;
  wire sig00000581;
  wire sig00000582;
  wire sig00000583;
  wire sig00000584;
  wire sig00000585;
  wire sig00000586;
  wire sig00000587;
  wire sig00000588;
  wire sig00000589;
  wire sig0000058a;
  wire sig0000058b;
  wire sig0000058c;
  wire sig0000058d;
  wire sig0000058e;
  wire sig0000058f;
  wire sig00000590;
  wire sig00000591;
  wire sig00000592;
  wire sig00000593;
  wire sig00000594;
  wire sig00000595;
  wire sig00000596;
  wire sig00000597;
  wire sig00000598;
  wire sig00000599;
  wire sig0000059a;
  wire sig0000059b;
  wire sig0000059c;
  wire sig0000059d;
  wire sig0000059e;
  wire sig0000059f;
  wire sig000005a0;
  wire sig000005a1;
  wire sig000005a2;
  wire sig000005a3;
  wire sig000005a4;
  wire sig000005a5;
  wire sig000005a6;
  wire sig000005a7;
  wire sig000005a8;
  wire sig000005a9;
  wire sig000005aa;
  wire sig000005ab;
  wire sig000005ac;
  wire sig000005ad;
  wire sig000005ae;
  wire sig000005af;
  wire sig000005b0;
  wire sig000005b1;
  wire sig000005b2;
  wire sig000005b3;
  wire sig000005b4;
  wire sig000005b5;
  wire sig000005b6;
  wire sig000005b7;
  wire sig000005b8;
  wire sig000005b9;
  wire sig000005ba;
  wire sig000005bb;
  wire sig000005bc;
  wire sig000005bd;
  wire sig000005be;
  wire sig000005bf;
  wire sig000005c0;
  wire sig000005c1;
  wire sig000005c2;
  wire sig000005c3;
  wire sig000005c4;
  wire sig000005c5;
  wire sig000005c6;
  wire sig000005c7;
  wire sig000005c8;
  wire sig000005c9;
  wire sig000005ca;
  wire sig000005cb;
  wire sig000005cc;
  wire sig000005cd;
  wire sig000005ce;
  wire sig000005cf;
  wire sig000005d0;
  wire sig000005d1;
  wire sig000005d2;
  wire sig000005d3;
  wire sig000005d4;
  wire sig000005d5;
  wire sig000005d6;
  wire sig000005d7;
  wire sig000005d8;
  wire sig000005d9;
  wire sig000005da;
  wire sig000005db;
  wire sig000005dc;
  wire sig000005dd;
  wire sig000005de;
  wire sig000005df;
  wire sig000005e0;
  wire sig000005e1;
  wire sig000005e2;
  wire sig000005e3;
  wire sig000005e4;
  wire sig000005e5;
  wire sig000005e6;
  wire sig000005e7;
  wire sig000005e8;
  wire sig000005e9;
  wire sig000005ea;
  wire sig000005eb;
  wire sig000005ec;
  wire sig000005ed;
  wire sig000005ee;
  wire sig000005ef;
  wire sig000005f0;
  wire sig000005f1;
  wire sig000005f2;
  wire sig000005f3;
  wire sig000005f4;
  wire sig000005f5;
  wire sig000005f6;
  wire sig000005f7;
  wire sig000005f8;
  wire sig000005f9;
  wire sig000005fa;
  wire sig000005fb;
  wire sig000005fc;
  wire sig000005fd;
  wire sig000005fe;
  wire sig000005ff;
  wire sig00000600;
  wire sig00000601;
  wire sig00000602;
  wire sig00000603;
  wire sig00000604;
  wire sig00000605;
  wire sig00000606;
  wire sig00000607;
  wire sig00000620;
  wire sig00000621;
  wire sig00000622;
  wire sig00000623;
  wire sig00000624;
  wire sig00000625;
  wire sig00000626;
  wire sig00000627;
  wire sig00000628;
  wire sig00000629;
  wire sig0000062a;
  wire sig00000633;
  wire sig00000634;
  wire sig00000635;
  wire sig00000636;
  wire sig00000637;
  wire sig00000638;
  wire sig00000639;
  wire sig0000063a;
  wire sig0000063b;
  wire sig0000063c;
  wire sig0000063d;
  wire sig0000063e;
  wire sig0000063f;
  wire sig00000640;
  wire sig00000641;
  wire sig00000643;
  wire sig00000644;
  wire sig00000645;
  wire sig00000646;
  wire sig00000647;
  wire sig00000648;
  wire sig00000649;
  wire sig0000064a;
  wire sig0000064b;
  wire sig0000064c;
  wire sig0000064d;
  wire sig0000064e;
  wire sig0000064f;
  wire sig00000650;
  wire sig00000651;
  wire sig00000652;
  wire sig00000653;
  wire sig00000654;
  wire sig00000655;
  wire sig00000656;
  wire sig00000657;
  wire sig00000658;
  wire sig00000659;
  wire sig0000065a;
  wire sig0000065b;
  wire sig0000065c;
  wire sig0000065d;
  wire sig0000065e;
  wire sig0000065f;
  wire sig00000660;
  wire sig00000661;
  wire sig00000662;
  wire sig00000663;
  wire sig00000664;
  wire sig00000665;
  wire sig00000666;
  wire sig00000667;
  wire sig00000668;
  wire sig00000669;
  wire sig0000066a;
  wire sig0000066b;
  wire sig0000066c;
  wire sig0000066d;
  wire sig0000066e;
  wire sig0000066f;
  wire sig00000670;
  wire sig00000671;
  wire sig00000672;
  wire sig00000673;
  wire sig00000674;
  wire sig00000675;
  wire sig00000676;
  wire sig00000677;
  wire sig00000678;
  wire sig00000679;
  wire sig0000067a;
  wire sig0000067b;
  wire sig0000067c;
  wire sig0000067d;
  wire sig0000067e;
  wire sig0000067f;
  wire sig00000680;
  wire sig00000688;
  wire sig00000689;
  wire sig0000068a;
  wire sig0000068b;
  wire sig0000068c;
  wire sig0000068d;
  wire sig0000068e;
  wire sig0000068f;
  wire sig00000690;
  wire sig00000691;
  wire sig00000692;
  wire sig00000693;
  wire sig00000694;
  wire sig00000695;
  wire sig00000696;
  wire sig00000697;
  wire sig00000698;
  wire sig00000699;
  wire sig0000069b;
  wire sig0000069c;
  wire sig0000069d;
  wire sig0000069e;
  wire sig0000069f;
  wire sig000006a0;
  wire sig000006a1;
  wire sig000006a2;
  wire sig000006a3;
  wire sig000006a4;
  wire sig000006a5;
  wire sig000006a6;
  wire sig000006a7;
  wire sig000006a8;
  wire sig000006a9;
  wire sig000006ab;
  wire sig000006ac;
  wire sig000006ad;
  wire sig000006ae;
  wire sig000006af;
  wire sig000006b0;
  wire sig000006b1;
  wire sig000006b2;
  wire sig000006b3;
  wire sig000006cc;
  wire sig000006cd;
  wire sig000006ce;
  wire sig000006cf;
  wire sig000006d0;
  wire sig000006d1;
  wire sig000006d2;
  wire sig000006d3;
  wire sig000006d4;
  wire sig000006d5;
  wire sig000006ef;
  wire sig000006f0;
  wire sig000006f1;
  wire sig000006f2;
  wire sig000006f3;
  wire sig000006f4;
  wire sig000006f5;
  wire sig000006f6;
  wire sig000006f7;
  wire sig000006f8;
  wire sig000006f9;
  wire sig000006fa;
  wire sig000006fb;
  wire sig000006fc;
  wire sig000006fd;
  wire sig000006fe;
  wire sig000006ff;
  wire sig00000700;
  wire sig00000749;
  wire sig0000074a;
  wire sig0000074b;
  wire sig0000074c;
  wire sig0000074d;
  wire sig0000074e;
  wire sig0000074f;
  wire sig00000750;
  wire sig00000751;
  wire sig00000752;
  wire sig00000753;
  wire sig00000754;
  wire sig00000755;
  wire sig00000756;
  wire sig00000757;
  wire sig00000758;
  wire sig00000769;
  wire sig0000076a;
  wire sig0000076b;
  wire sig0000076c;
  wire sig0000076d;
  wire sig0000076e;
  wire sig0000076f;
  wire sig00000770;
  wire sig00000771;
  wire sig00000772;
  wire sig00000773;
  wire sig00000774;
  wire sig00000775;
  wire sig00000776;
  wire sig00000777;
  wire sig00000778;
  wire sig00000789;
  wire sig0000078a;
  wire sig0000078b;
  wire sig0000078c;
  wire sig0000078d;
  wire sig0000078e;
  wire sig0000078f;
  wire sig00000790;
  wire sig00000791;
  wire sig00000792;
  wire sig00000793;
  wire sig00000794;
  wire sig00000795;
  wire sig00000796;
  wire sig00000797;
  wire sig00000798;
  wire sig00000799;
  wire sig0000079a;
  wire sig000007ad;
  wire sig000007ae;
  wire sig000007af;
  wire sig000007b0;
  wire sig000007b1;
  wire sig000007b2;
  wire sig000007b3;
  wire sig000007b4;
  wire sig000007b5;
  wire sig000007b6;
  wire sig000007b7;
  wire sig000007b8;
  wire sig000007b9;
  wire sig000007ba;
  wire sig000007bb;
  wire sig000007bc;
  wire sig000007bd;
  wire sig000007be;
  wire sig000007bf;
  wire sig000007c0;
  wire sig000007c1;
  wire sig000007c2;
  wire sig000007c3;
  wire sig000007c4;
  wire sig000007c5;
  wire sig000007c6;
  wire sig000007c7;
  wire sig000007c8;
  wire sig000007c9;
  wire sig000007ca;
  wire sig000007cb;
  wire sig000007cc;
  wire sig000007cd;
  wire sig000007ce;
  wire sig000007cf;
  wire sig000007d0;
  wire sig000007d1;
  wire sig000007d2;
  wire sig000007d3;
  wire sig000007d4;
  wire sig000007d5;
  wire sig000007d6;
  wire sig000007d7;
  wire sig000007d8;
  wire sig000007d9;
  wire sig000007da;
  wire sig000007db;
  wire sig000007dc;
  wire sig000007dd;
  wire sig000007de;
  wire sig000007df;
  wire sig000007e0;
  wire sig000007e1;
  wire sig000007e2;
  wire sig000007e3;
  wire sig000007e4;
  wire sig000007e5;
  wire sig000007e6;
  wire sig000007e7;
  wire sig000007e8;
  wire sig000007e9;
  wire sig000007ea;
  wire sig000007eb;
  wire sig000007ec;
  wire sig000007ed;
  wire sig000007ee;
  wire sig000007ef;
  wire sig000007f0;
  wire sig000007f1;
  wire sig000007f2;
  wire sig000007f3;
  wire sig000007f4;
  wire sig000007f5;
  wire sig000007f6;
  wire sig000007f7;
  wire sig000007f8;
  wire sig000007f9;
  wire sig000007fa;
  wire sig000007fb;
  wire sig000007fc;
  wire sig000007fd;
  wire sig000007fe;
  wire sig000007ff;
  wire sig00000800;
  wire sig00000801;
  wire sig00000802;
  wire sig00000803;
  wire sig00000804;
  wire sig00000805;
  wire sig00000806;
  wire sig00000807;
  wire sig00000808;
  wire sig00000809;
  wire sig0000080a;
  wire sig0000080b;
  wire sig0000080c;
  wire sig0000080d;
  wire sig0000080e;
  wire sig0000080f;
  wire sig00000810;
  wire sig00000811;
  wire sig00000812;
  wire sig00000813;
  wire sig00000814;
  wire sig00000815;
  wire sig00000816;
  wire sig00000817;
  wire sig00000818;
  wire sig00000819;
  wire sig0000081a;
  wire sig0000081b;
  wire sig0000081c;
  wire sig0000081d;
  wire sig0000081e;
  wire sig0000081f;
  wire sig00000820;
  wire sig00000821;
  wire sig00000822;
  wire sig00000823;
  wire sig00000824;
  wire sig00000825;
  wire sig00000826;
  wire sig00000827;
  wire sig00000828;
  wire sig00000829;
  wire sig0000082a;
  wire sig0000082b;
  wire sig0000082c;
  wire sig0000082d;
  wire sig0000082e;
  wire sig0000082f;
  wire sig00000830;
  wire sig00000831;
  wire sig00000832;
  wire sig00000833;
  wire sig00000834;
  wire sig00000835;
  wire sig00000836;
  wire sig00000837;
  wire sig00000838;
  wire sig00000839;
  wire sig0000083a;
  wire sig0000083b;
  wire sig0000083c;
  wire sig0000083d;
  wire sig0000083e;
  wire sig0000083f;
  wire sig00000840;
  wire sig00000841;
  wire sig00000842;
  wire sig00000843;
  wire sig00000844;
  wire sig00000845;
  wire sig00000846;
  wire sig00000847;
  wire sig00000848;
  wire sig00000849;
  wire sig0000084a;
  wire sig0000084b;
  wire sig0000084c;
  wire sig0000084d;
  wire sig0000084e;
  wire sig0000084f;
  wire sig00000850;
  wire sig00000851;
  wire sig00000852;
  wire sig00000853;
  wire sig00000854;
  wire sig00000855;
  wire sig00000856;
  wire sig00000857;
  wire sig00000858;
  wire sig00000859;
  wire sig0000085a;
  wire sig0000085b;
  wire sig0000085c;
  wire sig0000085d;
  wire sig0000085e;
  wire sig0000085f;
  wire sig00000860;
  wire sig00000861;
  wire sig00000862;
  wire sig00000863;
  wire sig00000864;
  wire sig00000865;
  wire sig00000866;
  wire sig00000867;
  wire sig00000868;
  wire sig00000869;
  wire sig0000086a;
  wire sig0000086b;
  wire sig0000086c;
  wire sig0000086d;
  wire sig0000086e;
  wire sig0000086f;
  wire sig00000870;
  wire sig00000871;
  wire sig00000872;
  wire sig00000873;
  wire sig00000874;
  wire sig00000875;
  wire sig00000876;
  wire sig00000877;
  wire sig00000878;
  wire sig00000879;
  wire sig0000087a;
  wire sig0000087b;
  wire sig0000087c;
  wire sig0000087d;
  wire sig0000087e;
  wire sig0000087f;
  wire sig00000880;
  wire sig00000881;
  wire sig00000882;
  wire sig00000883;
  wire sig00000884;
  wire sig00000885;
  wire sig00000886;
  wire sig00000887;
  wire sig00000888;
  wire sig00000889;
  wire sig0000088a;
  wire sig0000088b;
  wire sig0000088c;
  wire sig0000088d;
  wire sig0000088e;
  wire sig0000088f;
  wire sig00000890;
  wire sig00000891;
  wire sig00000892;
  wire sig00000893;
  wire sig00000894;
  wire sig00000895;
  wire sig00000896;
  wire sig00000897;
  wire sig00000898;
  wire sig00000899;
  wire sig0000089a;
  wire sig0000089b;
  wire sig0000089c;
  wire sig0000089d;
  wire sig0000089e;
  wire sig0000089f;
  wire sig000008a0;
  wire sig000008a1;
  wire sig000008a2;
  wire sig000008a3;
  wire sig000008a4;
  wire sig000008a5;
  wire sig000008a6;
  wire sig000008a7;
  wire sig000008a8;
  wire sig000008a9;
  wire sig000008aa;
  wire sig000008ab;
  wire sig000008ac;
  wire sig000008ad;
  wire sig000008ae;
  wire sig000008af;
  wire sig000008b0;
  wire sig000008b1;
  wire sig000008b2;
  wire sig000008b3;
  wire sig000008b4;
  wire sig000008b5;
  wire sig000008b6;
  wire sig000008b7;
  wire sig000008b8;
  wire sig000008b9;
  wire sig000008ba;
  wire sig000008bb;
  wire sig000008bc;
  wire sig000008bd;
  wire sig000008be;
  wire sig000008bf;
  wire sig000008c0;
  wire sig000008c1;
  wire sig000008c2;
  wire sig000008c3;
  wire sig000008c4;
  wire sig000008c5;
  wire sig000008c6;
  wire sig000008c7;
  wire sig000008c8;
  wire sig000008c9;
  wire sig000008ca;
  wire sig000008cb;
  wire sig000008cc;
  wire sig000008cd;
  wire sig000008ce;
  wire sig000008cf;
  wire sig000008d0;
  wire sig000008d1;
  wire sig000008d2;
  wire sig000008d3;
  wire sig000008d4;
  wire sig000008d5;
  wire sig000008d6;
  wire sig000008d7;
  wire sig000008d8;
  wire sig000008d9;
  wire sig000008da;
  wire sig000008db;
  wire sig000008dc;
  wire sig000008dd;
  wire sig000008de;
  wire sig000008df;
  wire sig000008e0;
  wire sig000008e1;
  wire sig000008e2;
  wire sig000008e3;
  wire sig000008e4;
  wire sig000008e5;
  wire sig000008e6;
  wire sig000008e7;
  wire sig000008e8;
  wire sig000008e9;
  wire sig000008ea;
  wire sig000008eb;
  wire sig000008ec;
  wire sig000008ed;
  wire sig000008ee;
  wire sig000008ef;
  wire sig000008f0;
  wire sig000008f1;
  wire sig000008f2;
  wire sig000008f3;
  wire sig000008f4;
  wire sig000008f5;
  wire sig000008f6;
  wire sig000008f7;
  wire sig000008f8;
  wire sig000008f9;
  wire sig000008fa;
  wire sig000008fb;
  wire sig000008fc;
  wire sig000008fd;
  wire sig000008fe;
  wire sig000008ff;
  wire sig00000900;
  wire sig00000901;
  wire sig00000902;
  wire sig00000903;
  wire sig00000904;
  wire sig00000905;
  wire sig00000906;
  wire sig00000907;
  wire sig00000908;
  wire sig00000909;
  wire sig0000090a;
  wire sig0000090b;
  wire sig0000090c;
  wire sig0000090d;
  wire sig0000090e;
  wire sig0000090f;
  wire sig00000910;
  wire sig00000911;
  wire sig00000912;
  wire sig00000913;
  wire sig00000914;
  wire sig00000915;
  wire sig00000916;
  wire sig00000917;
  wire sig00000918;
  wire sig00000919;
  wire sig0000091a;
  wire sig0000091b;
  wire sig0000091c;
  wire sig0000091d;
  wire sig0000091e;
  wire sig0000091f;
  wire sig00000920;
  wire sig00000921;
  wire sig00000922;
  wire sig00000923;
  wire sig00000924;
  wire sig00000925;
  wire sig00000926;
  wire sig00000927;
  wire sig00000928;
  wire sig00000929;
  wire sig0000092a;
  wire sig0000092b;
  wire sig0000092c;
  wire sig0000092d;
  wire sig0000092e;
  wire sig0000092f;
  wire sig00000930;
  wire sig00000931;
  wire sig00000932;
  wire sig00000933;
  wire sig00000934;
  wire sig00000935;
  wire sig00000936;
  wire sig00000937;
  wire sig00000938;
  wire sig00000939;
  wire sig0000093a;
  wire sig0000093b;
  wire sig0000093c;
  wire sig0000093d;
  wire sig0000093e;
  wire sig0000093f;
  wire sig00000940;
  wire sig00000941;
  wire sig00000942;
  wire sig00000943;
  wire sig00000944;
  wire sig00000945;
  wire sig00000946;
  wire sig00000947;
  wire sig00000948;
  wire sig00000949;
  wire sig0000094a;
  wire sig0000094b;
  wire sig0000094c;
  wire sig0000094d;
  wire sig0000094e;
  wire sig0000094f;
  wire sig00000950;
  wire sig00000951;
  wire sig00000952;
  wire sig00000953;
  wire sig00000954;
  wire sig00000955;
  wire sig00000956;
  wire sig00000957;
  wire sig00000958;
  wire sig00000959;
  wire sig0000095a;
  wire sig0000095b;
  wire sig0000095c;
  wire sig0000095d;
  wire sig0000095e;
  wire sig0000095f;
  wire sig00000960;
  wire sig00000961;
  wire sig00000962;
  wire sig00000963;
  wire sig00000964;
  wire sig00000965;
  wire sig00000966;
  wire sig00000967;
  wire sig00000968;
  wire sig00000969;
  wire sig0000096a;
  wire sig0000096b;
  wire sig0000096c;
  wire sig0000096d;
  wire sig0000096e;
  wire sig0000096f;
  wire sig00000970;
  wire sig00000971;
  wire sig00000972;
  wire sig00000973;
  wire sig00000974;
  wire sig00000975;
  wire sig00000976;
  wire sig00000977;
  wire sig00000978;
  wire sig00000979;
  wire sig0000097a;
  wire sig0000097b;
  wire sig0000097c;
  wire sig0000097d;
  wire sig0000097e;
  wire sig0000097f;
  wire sig00000980;
  wire sig00000981;
  wire sig00000982;
  wire sig00000983;
  wire sig00000984;
  wire sig00000985;
  wire sig00000986;
  wire sig00000987;
  wire sig00000988;
  wire sig00000989;
  wire sig0000098a;
  wire sig0000098b;
  wire sig0000098c;
  wire sig0000098d;
  wire sig0000098e;
  wire sig0000098f;
  wire sig00000990;
  wire sig00000991;
  wire sig00000992;
  wire sig00000993;
  wire sig00000994;
  wire sig00000995;
  wire sig00000996;
  wire sig00000997;
  wire sig00000998;
  wire sig00000999;
  wire sig0000099a;
  wire sig0000099b;
  wire sig0000099c;
  wire sig0000099d;
  wire sig0000099e;
  wire sig0000099f;
  wire sig000009a0;
  wire sig000009a1;
  wire sig000009a2;
  wire sig000009a3;
  wire sig000009a4;
  wire sig000009a5;
  wire sig000009a6;
  wire sig000009a7;
  wire sig000009a8;
  wire sig000009a9;
  wire sig000009aa;
  wire sig000009ab;
  wire sig000009ac;
  wire sig000009ad;
  wire sig000009ae;
  wire sig000009af;
  wire sig000009b0;
  wire sig000009b1;
  wire sig000009b2;
  wire sig000009b3;
  wire sig000009b4;
  wire sig000009b5;
  wire sig000009b6;
  wire sig000009b7;
  wire sig000009b8;
  wire sig000009b9;
  wire sig000009ba;
  wire sig000009bb;
  wire sig000009bc;
  wire sig000009bd;
  wire sig000009be;
  wire sig000009bf;
  wire sig000009c0;
  wire sig000009c1;
  wire sig000009c2;
  wire sig000009c3;
  wire sig000009c4;
  wire sig000009c5;
  wire sig000009c6;
  wire sig000009c7;
  wire sig000009c8;
  wire sig000009c9;
  wire sig000009ca;
  wire sig000009cb;
  wire sig000009cc;
  wire sig000009cd;
  wire sig000009ce;
  wire sig000009cf;
  wire sig000009d0;
  wire sig000009d1;
  wire sig000009d2;
  wire sig000009d3;
  wire sig000009d4;
  wire sig000009d5;
  wire sig000009d6;
  wire sig000009d7;
  wire sig000009d8;
  wire sig000009d9;
  wire sig000009da;
  wire sig000009db;
  wire sig000009dc;
  wire sig000009dd;
  wire sig000009de;
  wire sig000009df;
  wire sig000009e0;
  wire sig000009e1;
  wire sig000009e2;
  wire sig000009e3;
  wire sig000009e4;
  wire sig000009e5;
  wire sig000009e6;
  wire sig000009e7;
  wire sig000009e8;
  wire sig000009e9;
  wire sig000009ea;
  wire sig000009eb;
  wire sig000009ec;
  wire sig000009ed;
  wire sig000009ee;
  wire sig000009ef;
  wire sig000009f0;
  wire sig000009f1;
  wire sig000009f2;
  wire sig000009f3;
  wire sig000009f4;
  wire sig000009f5;
  wire sig000009f6;
  wire sig000009f7;
  wire sig000009f8;
  wire sig000009f9;
  wire sig000009fa;
  wire sig000009fb;
  wire sig000009fc;
  wire sig000009fd;
  wire sig000009fe;
  wire sig000009ff;
  wire sig00000a00;
  wire sig00000a01;
  wire sig00000a02;
  wire sig00000a03;
  wire sig00000a04;
  wire sig00000a05;
  wire sig00000a06;
  wire sig00000a07;
  wire sig00000a08;
  wire sig00000a09;
  wire sig00000a0a;
  wire sig00000a0b;
  wire sig00000a0c;
  wire sig00000a0d;
  wire sig00000a0e;
  wire sig00000a0f;
  wire sig00000a10;
  wire sig00000a11;
  wire sig00000a12;
  wire sig00000a13;
  wire sig00000a14;
  wire sig00000a15;
  wire sig00000a16;
  wire sig00000a17;
  wire sig00000a18;
  wire sig00000a19;
  wire sig00000a1a;
  wire sig00000a1b;
  wire sig00000a1c;
  wire sig00000a1d;
  wire sig00000a1e;
  wire sig00000a1f;
  wire sig00000a20;
  wire sig00000a21;
  wire sig00000a22;
  wire sig00000a23;
  wire sig00000a24;
  wire sig00000a25;
  wire sig00000a26;
  wire sig00000a27;
  wire sig00000a28;
  wire sig00000a29;
  wire sig00000a2a;
  wire sig00000a2b;
  wire sig00000a2c;
  wire sig00000a2d;
  wire sig00000a2e;
  wire sig00000a2f;
  wire sig00000a30;
  wire sig00000a31;
  wire sig00000a32;
  wire sig00000a33;
  wire sig00000a34;
  wire sig00000a35;
  wire sig00000a36;
  wire sig00000a37;
  wire sig00000a38;
  wire sig00000a39;
  wire sig00000a3a;
  wire sig00000a3b;
  wire sig00000a3c;
  wire sig00000a3d;
  wire sig00000a3e;
  wire sig00000a3f;
  wire sig00000a40;
  wire sig00000a41;
  wire sig00000a42;
  wire sig00000a43;
  wire sig00000a44;
  wire sig00000a45;
  wire sig00000a46;
  wire sig00000a47;
  wire sig00000a48;
  wire sig00000a49;
  wire sig00000a4a;
  wire sig00000a4b;
  wire sig00000a4c;
  wire sig00000a4d;
  wire sig00000a4e;
  wire sig00000a4f;
  wire sig00000a50;
  wire sig00000a51;
  wire sig00000a52;
  wire sig00000a53;
  wire sig00000a54;
  wire sig00000a55;
  wire sig00000a56;
  wire sig00000a57;
  wire sig00000a58;
  wire sig00000a59;
  wire sig00000a5a;
  wire sig00000a5b;
  wire sig00000a5c;
  wire sig00000a5d;
  wire sig00000a5e;
  wire sig00000a5f;
  wire sig00000a60;
  wire sig00000a61;
  wire sig00000a62;
  wire sig00000a63;
  wire sig00000a64;
  wire sig00000a65;
  wire sig00000a66;
  wire sig00000a67;
  wire sig00000a68;
  wire sig00000a69;
  wire sig00000a6a;
  wire sig00000a6b;
  wire sig00000a6c;
  wire sig00000a6d;
  wire sig00000a6e;
  wire sig00000a6f;
  wire sig00000a70;
  wire sig00000a71;
  wire sig00000a72;
  wire sig00000a73;
  wire sig00000a74;
  wire sig00000a75;
  wire sig00000a76;
  wire sig00000a77;
  wire sig00000a78;
  wire sig00000a79;
  wire sig00000a7a;
  wire sig00000a7b;
  wire sig00000a7c;
  wire sig00000a7d;
  wire sig00000a7e;
  wire sig00000a7f;
  wire sig00000a80;
  wire sig00000a81;
  wire sig00000a82;
  wire sig00000a83;
  wire sig00000a84;
  wire sig00000a85;
  wire sig00000a86;
  wire sig00000a87;
  wire sig00000a88;
  wire sig00000a89;
  wire sig00000a8a;
  wire sig00000a8b;
  wire sig00000a8c;
  wire sig00000a8d;
  wire sig00000a8e;
  wire sig00000a8f;
  wire sig00000a90;
  wire sig00000a91;
  wire sig00000a92;
  wire sig00000a93;
  wire sig00000a94;
  wire sig00000a95;
  wire sig00000a96;
  wire sig00000a97;
  wire sig00000a98;
  wire sig00000a99;
  wire sig00000a9a;
  wire sig00000a9b;
  wire sig00000a9c;
  wire sig00000a9d;
  wire sig00000a9e;
  wire sig00000a9f;
  wire sig00000aa0;
  wire sig00000aa1;
  wire sig00000aa2;
  wire sig00000aa3;
  wire sig00000aa4;
  wire sig00000aa5;
  wire sig00000aa6;
  wire sig00000aa7;
  wire sig00000aa8;
  wire sig00000aa9;
  wire sig00000aaa;
  wire sig00000aab;
  wire sig00000aac;
  wire sig00000aad;
  wire sig00000aae;
  wire sig00000aaf;
  wire sig00000ab0;
  wire sig00000ab1;
  wire sig00000ab2;
  wire sig00000ab3;
  wire sig00000ab4;
  wire sig00000ab5;
  wire sig00000ab6;
  wire sig00000ab7;
  wire sig00000ab8;
  wire sig00000ab9;
  wire sig00000aba;
  wire sig00000abb;
  wire sig00000abc;
  wire sig00000abd;
  wire sig00000abe;
  wire sig00000abf;
  wire sig00000ac0;
  wire sig00000ac1;
  wire sig00000ac2;
  wire sig00000ac3;
  wire sig00000ac4;
  wire sig00000ac5;
  wire sig00000ac6;
  wire sig00000ac7;
  wire sig00000ac8;
  wire sig00000ac9;
  wire sig00000aca;
  wire sig00000acb;
  wire sig00000acc;
  wire sig00000acd;
  wire sig00000ace;
  wire sig00000acf;
  wire sig00000ad0;
  wire sig00000ad1;
  wire sig00000ad2;
  wire sig00000ad3;
  wire sig00000ad4;
  wire sig00000ad5;
  wire sig00000ad6;
  wire sig00000ad7;
  wire sig00000ad8;
  wire sig00000ad9;
  wire sig00000ada;
  wire sig00000adb;
  wire sig00000adc;
  wire sig00000add;
  wire sig00000ade;
  wire sig00000adf;
  wire sig00000ae0;
  wire sig00000ae1;
  wire sig00000ae2;
  wire sig00000ae3;
  wire sig00000ae4;
  wire sig00000ae5;
  wire sig00000ae6;
  wire sig00000ae7;
  wire sig00000ae8;
  wire sig00000ae9;
  wire sig00000aea;
  wire sig00000aeb;
  wire sig00000aec;
  wire sig00000aed;
  wire sig00000aee;
  wire sig00000aef;
  wire sig00000af0;
  wire sig00000af1;
  wire sig00000af2;
  wire sig00000af3;
  wire sig00000af4;
  wire sig00000af5;
  wire sig00000af6;
  wire sig00000af7;
  wire sig00000af8;
  wire sig00000af9;
  wire sig00000afa;
  wire sig00000afb;
  wire sig00000afc;
  wire sig00000afd;
  wire sig00000afe;
  wire sig00000aff;
  wire sig00000b00;
  wire sig00000b01;
  wire sig00000b02;
  wire sig00000b03;
  wire sig00000b04;
  wire sig00000b05;
  wire sig00000b06;
  wire sig00000b07;
  wire sig00000b08;
  wire sig00000b09;
  wire sig00000b0a;
  wire sig00000b0b;
  wire sig00000b0c;
  wire sig00000b0d;
  wire sig00000b0e;
  wire sig00000b0f;
  wire sig00000b10;
  wire sig00000b11;
  wire sig00000b12;
  wire sig00000b13;
  wire sig00000b14;
  wire sig00000b15;
  wire sig00000b16;
  wire sig00000b17;
  wire sig00000b18;
  wire sig00000b19;
  wire sig00000b1a;
  wire sig00000b1b;
  wire sig00000b1c;
  wire sig00000b1d;
  wire sig00000b1e;
  wire sig00000b1f;
  wire sig00000b20;
  wire sig00000b21;
  wire sig00000b22;
  wire sig00000b23;
  wire sig00000b24;
  wire sig00000b25;
  wire sig00000b26;
  wire sig00000b27;
  wire sig00000b28;
  wire sig00000b29;
  wire sig00000b2a;
  wire sig00000b2b;
  wire sig00000b2c;
  wire sig00000b2d;
  wire sig00000b2e;
  wire sig00000b2f;
  wire sig00000b30;
  wire sig00000b31;
  wire sig00000b32;
  wire sig00000b33;
  wire sig00000b34;
  wire sig00000b35;
  wire sig00000b36;
  wire sig00000b37;
  wire sig00000b38;
  wire sig00000b39;
  wire sig00000b3a;
  wire sig00000b3b;
  wire sig00000b3c;
  wire sig00000b3d;
  wire sig00000b3e;
  wire sig00000b3f;
  wire sig00000b40;
  wire sig00000b41;
  wire sig00000b42;
  wire sig00000b43;
  wire sig00000b44;
  wire sig00000b45;
  wire sig00000b46;
  wire sig00000b47;
  wire sig00000b48;
  wire sig00000b49;
  wire sig00000b4a;
  wire sig00000b4b;
  wire sig00000b4c;
  wire sig00000b4d;
  wire sig00000b4e;
  wire sig00000b4f;
  wire sig00000b50;
  wire sig00000b51;
  wire sig00000b52;
  wire sig00000b53;
  wire sig00000b54;
  wire sig00000b55;
  wire sig00000b56;
  wire sig00000b57;
  wire sig00000b58;
  wire sig00000b59;
  wire sig00000b5a;
  wire sig00000b5b;
  wire sig00000b5c;
  wire sig00000b5d;
  wire sig00000b5e;
  wire sig00000b5f;
  wire sig00000b60;
  wire sig00000b61;
  wire sig00000b62;
  wire sig00000b63;
  wire sig00000b64;
  wire sig00000b65;
  wire sig00000b66;
  wire sig00000b67;
  wire sig00000b68;
  wire sig00000b69;
  wire sig00000b6a;
  wire sig00000b6b;
  wire sig00000b6c;
  wire sig00000b6d;
  wire sig00000b6e;
  wire sig00000b6f;
  wire sig00000b70;
  wire sig00000b71;
  wire sig00000b72;
  wire sig00000b73;
  wire sig00000b74;
  wire sig00000b75;
  wire sig00000b76;
  wire sig00000b77;
  wire sig00000b78;
  wire sig00000b79;
  wire sig00000b7a;
  wire sig00000b7b;
  wire sig00000b7c;
  wire sig00000b7d;
  wire sig00000b7e;
  wire sig00000b7f;
  wire sig00000b80;
  wire sig00000b81;
  wire sig00000b82;
  wire sig00000b83;
  wire sig00000b84;
  wire sig00000b85;
  wire sig00000b86;
  wire sig00000b87;
  wire sig00000b88;
  wire sig00000b89;
  wire sig00000b8a;
  wire sig00000b8b;
  wire sig00000b8c;
  wire sig00000b8d;
  wire sig00000b8e;
  wire sig00000b8f;
  wire sig00000b90;
  wire sig00000b91;
  wire sig00000b92;
  wire sig00000b93;
  wire sig00000b94;
  wire sig00000b95;
  wire sig00000b96;
  wire sig00000b97;
  wire sig00000b98;
  wire sig00000b99;
  wire sig00000b9a;
  wire sig00000b9b;
  wire sig00000b9c;
  wire sig00000b9d;
  wire sig00000b9e;
  wire sig00000b9f;
  wire sig00000ba0;
  wire sig00000ba1;
  wire sig00000ba2;
  wire sig00000ba3;
  wire sig00000ba4;
  wire sig00000ba5;
  wire sig00000ba6;
  wire sig00000ba7;
  wire sig00000ba8;
  wire sig00000ba9;
  wire sig00000baa;
  wire sig00000bab;
  wire sig00000bac;
  wire sig00000bad;
  wire sig00000bae;
  wire sig00000baf;
  wire sig00000bb0;
  wire sig00000bb1;
  wire sig00000bb2;
  wire sig00000bb3;
  wire sig00000bb4;
  wire sig00000bb5;
  wire sig00000bb6;
  wire sig00000bb7;
  wire sig00000bb8;
  wire sig00000bb9;
  wire sig00000bba;
  wire sig00000bbb;
  wire sig00000bbc;
  wire sig00000bbd;
  wire sig00000bbe;
  wire sig00000bbf;
  wire sig00000bc0;
  wire sig00000bc1;
  wire sig00000bc2;
  wire sig00000bc3;
  wire sig00000bc4;
  wire sig00000bc5;
  wire sig00000bc6;
  wire sig00000bc7;
  wire sig00000bc8;
  wire sig00000bc9;
  wire sig00000bca;
  wire sig00000bcb;
  wire sig00000bcc;
  wire sig00000bcd;
  wire sig00000bce;
  wire sig00000bcf;
  wire sig00000bd0;
  wire sig00000bd1;
  wire sig00000bd2;
  wire sig00000bd3;
  wire sig00000bd4;
  wire sig00000bd5;
  wire sig00000bd6;
  wire sig00000bd7;
  wire sig00000bd8;
  wire sig00000bd9;
  wire sig00000bda;
  wire sig00000bdb;
  wire sig00000bdc;
  wire sig00000bdd;
  wire sig00000bde;
  wire sig00000bdf;
  wire sig00000be0;
  wire sig00000be1;
  wire sig00000be2;
  wire sig00000be3;
  wire sig00000be4;
  wire sig00000be5;
  wire sig00000be6;
  wire sig00000be7;
  wire sig00000be8;
  wire sig00000be9;
  wire sig00000bea;
  wire sig00000beb;
  wire sig00000bec;
  wire sig00000bed;
  wire sig00000bee;
  wire sig00000bef;
  wire sig00000bf0;
  wire sig00000bf1;
  wire sig00000bf2;
  wire sig00000bf3;
  wire sig00000bf4;
  wire sig00000bf5;
  wire sig00000bf6;
  wire sig00000bf7;
  wire sig00000bf8;
  wire sig00000bf9;
  wire sig00000bfa;
  wire sig00000bfb;
  wire sig00000bfc;
  wire sig00000bfd;
  wire sig00000bfe;
  wire sig00000bff;
  wire sig00000c00;
  wire sig00000c01;
  wire sig00000c02;
  wire sig00000c03;
  wire sig00000c04;
  wire sig00000c05;
  wire sig00000c06;
  wire sig00000c07;
  wire sig00000c08;
  wire sig00000c09;
  wire sig00000c0a;
  wire sig00000c0b;
  wire sig00000c0c;
  wire sig00000c0d;
  wire sig00000c0e;
  wire sig00000c0f;
  wire sig00000c10;
  wire sig00000c11;
  wire sig00000c12;
  wire sig00000c13;
  wire sig00000c14;
  wire sig00000c15;
  wire sig00000c16;
  wire sig00000c17;
  wire sig00000c18;
  wire sig00000c19;
  wire sig00000c1a;
  wire sig00000c1b;
  wire sig00000c1c;
  wire sig00000c1d;
  wire sig00000c1e;
  wire sig00000c1f;
  wire sig00000c20;
  wire sig00000c21;
  wire sig00000c22;
  wire sig00000c23;
  wire sig00000c24;
  wire sig00000c25;
  wire sig00000c26;
  wire sig00000c27;
  wire sig00000c28;
  wire sig00000c29;
  wire sig00000c2a;
  wire sig00000c2b;
  wire sig00000c2c;
  wire sig00000c2d;
  wire sig00000c2e;
  wire sig00000c2f;
  wire sig00000c30;
  wire sig00000c31;
  wire sig00000c32;
  wire sig00000c33;
  wire sig00000c34;
  wire sig00000c35;
  wire sig00000c36;
  wire sig00000c37;
  wire sig00000c38;
  wire sig00000c39;
  wire sig00000c3a;
  wire sig00000c3b;
  wire sig00000c3c;
  wire sig00000c3d;
  wire sig00000c3e;
  wire sig00000c3f;
  wire sig00000c40;
  wire sig00000c41;
  wire sig00000c42;
  wire sig00000c43;
  wire sig00000c44;
  wire sig00000c45;
  wire sig00000c46;
  wire sig00000c47;
  wire sig00000c48;
  wire sig00000c49;
  wire sig00000c4a;
  wire sig00000c4b;
  wire sig00000c4c;
  wire sig00000c4d;
  wire sig00000c4e;
  wire sig00000c4f;
  wire sig00000c50;
  wire sig00000c51;
  wire sig00000c52;
  wire sig00000c53;
  wire sig00000c54;
  wire sig00000c55;
  wire sig00000c56;
  wire sig00000c57;
  wire sig00000c58;
  wire sig00000c59;
  wire sig00000c5a;
  wire sig00000c5b;
  wire sig00000c5c;
  wire sig00000c5d;
  wire sig00000c5e;
  wire sig00000c5f;
  wire sig00000c60;
  wire sig00000c61;
  wire sig00000c62;
  wire sig00000c63;
  wire sig00000c64;
  wire sig00000c65;
  wire sig00000c66;
  wire sig00000c67;
  wire sig00000c68;
  wire sig00000c69;
  wire sig00000c6a;
  wire sig00000c6b;
  wire sig00000c6c;
  wire sig00000c6d;
  wire sig00000c6e;
  wire sig00000c6f;
  wire sig00000c70;
  wire sig00000c71;
  wire sig00000c72;
  wire sig00000c73;
  wire sig00000c74;
  wire sig00000c75;
  wire sig00000c76;
  wire sig00000c77;
  wire sig00000c78;
  wire sig00000c79;
  wire sig00000c7a;
  wire sig00000c7b;
  wire sig00000c7c;
  wire sig00000c7d;
  wire sig00000c7e;
  wire sig00000c7f;
  wire sig00000c80;
  wire sig00000c81;
  wire sig00000c82;
  wire sig00000c83;
  wire sig00000c84;
  wire sig00000c85;
  wire sig00000c86;
  wire sig00000c87;
  wire sig00000c88;
  wire sig00000c89;
  wire sig00000c8a;
  wire sig00000c8b;
  wire sig00000c8c;
  wire sig00000c8d;
  wire sig00000c8e;
  wire sig00000c8f;
  wire sig00000c90;
  wire sig00000c91;
  wire sig00000c92;
  wire sig00000c93;
  wire sig00000c94;
  wire sig00000c95;
  wire sig00000c96;
  wire sig00000c97;
  wire sig00000c98;
  wire sig00000c99;
  wire sig00000c9a;
  wire sig00000c9b;
  wire sig00000c9c;
  wire sig00000c9d;
  wire sig00000c9e;
  wire sig00000c9f;
  wire sig00000ca0;
  wire sig00000ca1;
  wire sig00000ca2;
  wire sig00000ca3;
  wire sig00000ca4;
  wire sig00000ca5;
  wire sig00000ca6;
  wire sig00000ca7;
  wire sig00000ca8;
  wire sig00000ca9;
  wire sig00000caa;
  wire sig00000cab;
  wire sig00000cac;
  wire sig00000cad;
  wire \blk000000dc/sig00000cb4 ;
  wire \blk000000dc/sig00000cb3 ;
  wire \blk000000dc/sig00000cb2 ;
  wire \blk000001f6/sig00000cba ;
  wire \blk000001f6/sig00000cb9 ;
  wire \blk000001f6/sig00000cb8 ;
  wire \blk000002a3/sig00000cc3 ;
  wire \blk000002a3/sig00000cc2 ;
  wire \blk000002a3/sig00000cc1 ;
  wire \blk000002a3/sig00000cc0 ;
  wire \blk000002aa/sig00000cc9 ;
  wire \blk000002aa/sig00000cc8 ;
  wire \blk000002aa/sig00000cc7 ;
  wire \blk000002af/sig00000ccf ;
  wire \blk000002af/sig00000cce ;
  wire \blk000002af/sig00000ccd ;
  wire \blk000002b4/sig00000cd5 ;
  wire \blk000002b4/sig00000cd4 ;
  wire \blk000002b4/sig00000cd3 ;
  wire \blk000002b9/sig00000cde ;
  wire \blk000002b9/sig00000cdd ;
  wire \blk000002b9/sig00000cdc ;
  wire \blk000002b9/sig00000cdb ;
  wire \blk000002c0/sig00000ce7 ;
  wire \blk000002c0/sig00000ce6 ;
  wire \blk000002c0/sig00000ce5 ;
  wire \blk000002c0/sig00000ce4 ;
  wire \blk000003fc/sig00000ced ;
  wire \blk000003fc/sig00000cec ;
  wire \blk00000400/sig00000cf3 ;
  wire \blk00000400/sig00000cf2 ;
  wire \blk00000404/sig00000cf9 ;
  wire \blk00000404/sig00000cf8 ;
  wire \blk00000404/sig00000cf7 ;
  wire \blk00000503/sig00000cff ;
  wire \blk00000503/sig00000cfe ;
  wire \blk00000503/sig00000cfd ;
  wire \blk00000508/sig00000d05 ;
  wire \blk00000508/sig00000d04 ;
  wire \blk00000522/sig00000d2d ;
  wire \blk00000522/sig00000d2c ;
  wire \blk00000522/sig00000d2b ;
  wire \blk00000522/sig00000d2a ;
  wire \blk00000522/sig00000d29 ;
  wire \blk00000522/sig00000d27 ;
  wire \blk00000522/sig00000d26 ;
  wire \blk00000522/sig00000d25 ;
  wire \blk00000522/sig00000d24 ;
  wire \blk00000522/sig00000d23 ;
  wire \blk00000522/sig00000d21 ;
  wire \blk00000522/sig00000d20 ;
  wire \blk00000522/sig00000d1f ;
  wire \blk00000522/sig00000d1e ;
  wire \blk00000522/sig00000d1d ;
  wire \blk00000522/sig00000d1c ;
  wire \blk00000522/sig00000d1b ;
  wire \blk00000522/sig00000d1a ;
  wire \blk00000522/sig00000d19 ;
  wire \blk00000522/sig00000d18 ;
  wire \blk00000522/sig00000d17 ;
  wire \blk00000522/sig00000d16 ;
  wire \blk00000522/sig00000d0a ;
  wire \blk00000522/sig00000d09 ;
  wire \blk00000640/sig00000e36 ;
  wire \blk00000640/sig00000e35 ;
  wire \blk00000640/sig00000e34 ;
  wire \blk00000659/sig00000e3c ;
  wire \blk00000659/sig00000e3b ;
  wire \blk000007cb/sig00000e42 ;
  wire \blk000007cb/sig00000e41 ;
  wire \blk000007cb/sig00000e40 ;
  wire \blk0000083a/sig00000e48 ;
  wire \blk0000083a/sig00000e47 ;
  wire \blk0000083e/sig00000e4e ;
  wire \blk0000083e/sig00000e4d ;
  wire NLW_blk00000062_Q_UNCONNECTED;
  wire NLW_blk000000e6_Q_UNCONNECTED;
  wire NLW_blk000000e7_Q_UNCONNECTED;
  wire NLW_blk000000e8_Q_UNCONNECTED;
  wire NLW_blk000002cb_Q_UNCONNECTED;
  wire NLW_blk000002cc_Q_UNCONNECTED;
  wire NLW_blk000002cd_Q_UNCONNECTED;
  wire NLW_blk000002ce_Q_UNCONNECTED;
  wire NLW_blk000002d5_Q_UNCONNECTED;
  wire NLW_blk000002d6_Q_UNCONNECTED;
  wire NLW_blk00000341_O_UNCONNECTED;
  wire NLW_blk00000366_O_UNCONNECTED;
  wire NLW_blk00000510_O_UNCONNECTED;
  wire NLW_blk00000546_PATTERNBDETECT_UNCONNECTED;
  wire NLW_blk00000546_MULTSIGNOUT_UNCONNECTED;
  wire NLW_blk00000546_CARRYCASCOUT_UNCONNECTED;
  wire NLW_blk00000546_UNDERFLOW_UNCONNECTED;
  wire NLW_blk00000546_PATTERNDETECT_UNCONNECTED;
  wire NLW_blk00000546_OVERFLOW_UNCONNECTED;
  wire \NLW_blk00000546_ACOUT<29>_UNCONNECTED ;
  wire \NLW_blk00000546_ACOUT<28>_UNCONNECTED ;
  wire \NLW_blk00000546_ACOUT<27>_UNCONNECTED ;
  wire \NLW_blk00000546_ACOUT<26>_UNCONNECTED ;
  wire \NLW_blk00000546_ACOUT<25>_UNCONNECTED ;
  wire \NLW_blk00000546_ACOUT<24>_UNCONNECTED ;
  wire \NLW_blk00000546_ACOUT<23>_UNCONNECTED ;
  wire \NLW_blk00000546_ACOUT<22>_UNCONNECTED ;
  wire \NLW_blk00000546_ACOUT<21>_UNCONNECTED ;
  wire \NLW_blk00000546_ACOUT<20>_UNCONNECTED ;
  wire \NLW_blk00000546_ACOUT<19>_UNCONNECTED ;
  wire \NLW_blk00000546_ACOUT<18>_UNCONNECTED ;
  wire \NLW_blk00000546_ACOUT<17>_UNCONNECTED ;
  wire \NLW_blk00000546_ACOUT<16>_UNCONNECTED ;
  wire \NLW_blk00000546_ACOUT<15>_UNCONNECTED ;
  wire \NLW_blk00000546_ACOUT<14>_UNCONNECTED ;
  wire \NLW_blk00000546_ACOUT<13>_UNCONNECTED ;
  wire \NLW_blk00000546_ACOUT<12>_UNCONNECTED ;
  wire \NLW_blk00000546_ACOUT<11>_UNCONNECTED ;
  wire \NLW_blk00000546_ACOUT<10>_UNCONNECTED ;
  wire \NLW_blk00000546_ACOUT<9>_UNCONNECTED ;
  wire \NLW_blk00000546_ACOUT<8>_UNCONNECTED ;
  wire \NLW_blk00000546_ACOUT<7>_UNCONNECTED ;
  wire \NLW_blk00000546_ACOUT<6>_UNCONNECTED ;
  wire \NLW_blk00000546_ACOUT<5>_UNCONNECTED ;
  wire \NLW_blk00000546_ACOUT<4>_UNCONNECTED ;
  wire \NLW_blk00000546_ACOUT<3>_UNCONNECTED ;
  wire \NLW_blk00000546_ACOUT<2>_UNCONNECTED ;
  wire \NLW_blk00000546_ACOUT<1>_UNCONNECTED ;
  wire \NLW_blk00000546_ACOUT<0>_UNCONNECTED ;
  wire \NLW_blk00000546_CARRYOUT<3>_UNCONNECTED ;
  wire \NLW_blk00000546_CARRYOUT<2>_UNCONNECTED ;
  wire \NLW_blk00000546_CARRYOUT<1>_UNCONNECTED ;
  wire \NLW_blk00000546_CARRYOUT<0>_UNCONNECTED ;
  wire \NLW_blk00000546_BCOUT<17>_UNCONNECTED ;
  wire \NLW_blk00000546_BCOUT<16>_UNCONNECTED ;
  wire \NLW_blk00000546_BCOUT<15>_UNCONNECTED ;
  wire \NLW_blk00000546_BCOUT<14>_UNCONNECTED ;
  wire \NLW_blk00000546_BCOUT<13>_UNCONNECTED ;
  wire \NLW_blk00000546_BCOUT<12>_UNCONNECTED ;
  wire \NLW_blk00000546_BCOUT<11>_UNCONNECTED ;
  wire \NLW_blk00000546_BCOUT<10>_UNCONNECTED ;
  wire \NLW_blk00000546_BCOUT<9>_UNCONNECTED ;
  wire \NLW_blk00000546_BCOUT<8>_UNCONNECTED ;
  wire \NLW_blk00000546_BCOUT<7>_UNCONNECTED ;
  wire \NLW_blk00000546_BCOUT<6>_UNCONNECTED ;
  wire \NLW_blk00000546_BCOUT<5>_UNCONNECTED ;
  wire \NLW_blk00000546_BCOUT<4>_UNCONNECTED ;
  wire \NLW_blk00000546_BCOUT<3>_UNCONNECTED ;
  wire \NLW_blk00000546_BCOUT<2>_UNCONNECTED ;
  wire \NLW_blk00000546_BCOUT<1>_UNCONNECTED ;
  wire \NLW_blk00000546_BCOUT<0>_UNCONNECTED ;
  wire \NLW_blk00000546_P<47>_UNCONNECTED ;
  wire \NLW_blk00000546_P<46>_UNCONNECTED ;
  wire \NLW_blk00000546_P<45>_UNCONNECTED ;
  wire \NLW_blk00000546_P<44>_UNCONNECTED ;
  wire \NLW_blk00000546_P<43>_UNCONNECTED ;
  wire \NLW_blk00000546_PCOUT<47>_UNCONNECTED ;
  wire \NLW_blk00000546_PCOUT<46>_UNCONNECTED ;
  wire \NLW_blk00000546_PCOUT<45>_UNCONNECTED ;
  wire \NLW_blk00000546_PCOUT<44>_UNCONNECTED ;
  wire \NLW_blk00000546_PCOUT<43>_UNCONNECTED ;
  wire \NLW_blk00000546_PCOUT<42>_UNCONNECTED ;
  wire \NLW_blk00000546_PCOUT<41>_UNCONNECTED ;
  wire \NLW_blk00000546_PCOUT<40>_UNCONNECTED ;
  wire \NLW_blk00000546_PCOUT<39>_UNCONNECTED ;
  wire \NLW_blk00000546_PCOUT<38>_UNCONNECTED ;
  wire \NLW_blk00000546_PCOUT<37>_UNCONNECTED ;
  wire \NLW_blk00000546_PCOUT<36>_UNCONNECTED ;
  wire \NLW_blk00000546_PCOUT<35>_UNCONNECTED ;
  wire \NLW_blk00000546_PCOUT<34>_UNCONNECTED ;
  wire \NLW_blk00000546_PCOUT<33>_UNCONNECTED ;
  wire \NLW_blk00000546_PCOUT<32>_UNCONNECTED ;
  wire \NLW_blk00000546_PCOUT<31>_UNCONNECTED ;
  wire \NLW_blk00000546_PCOUT<30>_UNCONNECTED ;
  wire \NLW_blk00000546_PCOUT<29>_UNCONNECTED ;
  wire \NLW_blk00000546_PCOUT<28>_UNCONNECTED ;
  wire \NLW_blk00000546_PCOUT<27>_UNCONNECTED ;
  wire \NLW_blk00000546_PCOUT<26>_UNCONNECTED ;
  wire \NLW_blk00000546_PCOUT<25>_UNCONNECTED ;
  wire \NLW_blk00000546_PCOUT<24>_UNCONNECTED ;
  wire \NLW_blk00000546_PCOUT<23>_UNCONNECTED ;
  wire \NLW_blk00000546_PCOUT<22>_UNCONNECTED ;
  wire \NLW_blk00000546_PCOUT<21>_UNCONNECTED ;
  wire \NLW_blk00000546_PCOUT<20>_UNCONNECTED ;
  wire \NLW_blk00000546_PCOUT<19>_UNCONNECTED ;
  wire \NLW_blk00000546_PCOUT<18>_UNCONNECTED ;
  wire \NLW_blk00000546_PCOUT<17>_UNCONNECTED ;
  wire \NLW_blk00000546_PCOUT<16>_UNCONNECTED ;
  wire \NLW_blk00000546_PCOUT<15>_UNCONNECTED ;
  wire \NLW_blk00000546_PCOUT<14>_UNCONNECTED ;
  wire \NLW_blk00000546_PCOUT<13>_UNCONNECTED ;
  wire \NLW_blk00000546_PCOUT<12>_UNCONNECTED ;
  wire \NLW_blk00000546_PCOUT<11>_UNCONNECTED ;
  wire \NLW_blk00000546_PCOUT<10>_UNCONNECTED ;
  wire \NLW_blk00000546_PCOUT<9>_UNCONNECTED ;
  wire \NLW_blk00000546_PCOUT<8>_UNCONNECTED ;
  wire \NLW_blk00000546_PCOUT<7>_UNCONNECTED ;
  wire \NLW_blk00000546_PCOUT<6>_UNCONNECTED ;
  wire \NLW_blk00000546_PCOUT<5>_UNCONNECTED ;
  wire \NLW_blk00000546_PCOUT<4>_UNCONNECTED ;
  wire \NLW_blk00000546_PCOUT<3>_UNCONNECTED ;
  wire \NLW_blk00000546_PCOUT<2>_UNCONNECTED ;
  wire \NLW_blk00000546_PCOUT<1>_UNCONNECTED ;
  wire \NLW_blk00000546_PCOUT<0>_UNCONNECTED ;
  wire NLW_blk00000547_PATTERNBDETECT_UNCONNECTED;
  wire NLW_blk00000547_MULTSIGNOUT_UNCONNECTED;
  wire NLW_blk00000547_CARRYCASCOUT_UNCONNECTED;
  wire NLW_blk00000547_UNDERFLOW_UNCONNECTED;
  wire NLW_blk00000547_PATTERNDETECT_UNCONNECTED;
  wire NLW_blk00000547_OVERFLOW_UNCONNECTED;
  wire \NLW_blk00000547_ACOUT<29>_UNCONNECTED ;
  wire \NLW_blk00000547_ACOUT<28>_UNCONNECTED ;
  wire \NLW_blk00000547_ACOUT<27>_UNCONNECTED ;
  wire \NLW_blk00000547_ACOUT<26>_UNCONNECTED ;
  wire \NLW_blk00000547_ACOUT<25>_UNCONNECTED ;
  wire \NLW_blk00000547_ACOUT<24>_UNCONNECTED ;
  wire \NLW_blk00000547_ACOUT<23>_UNCONNECTED ;
  wire \NLW_blk00000547_ACOUT<22>_UNCONNECTED ;
  wire \NLW_blk00000547_ACOUT<21>_UNCONNECTED ;
  wire \NLW_blk00000547_ACOUT<20>_UNCONNECTED ;
  wire \NLW_blk00000547_ACOUT<19>_UNCONNECTED ;
  wire \NLW_blk00000547_ACOUT<18>_UNCONNECTED ;
  wire \NLW_blk00000547_ACOUT<17>_UNCONNECTED ;
  wire \NLW_blk00000547_ACOUT<16>_UNCONNECTED ;
  wire \NLW_blk00000547_ACOUT<15>_UNCONNECTED ;
  wire \NLW_blk00000547_ACOUT<14>_UNCONNECTED ;
  wire \NLW_blk00000547_ACOUT<13>_UNCONNECTED ;
  wire \NLW_blk00000547_ACOUT<12>_UNCONNECTED ;
  wire \NLW_blk00000547_ACOUT<11>_UNCONNECTED ;
  wire \NLW_blk00000547_ACOUT<10>_UNCONNECTED ;
  wire \NLW_blk00000547_ACOUT<9>_UNCONNECTED ;
  wire \NLW_blk00000547_ACOUT<8>_UNCONNECTED ;
  wire \NLW_blk00000547_ACOUT<7>_UNCONNECTED ;
  wire \NLW_blk00000547_ACOUT<6>_UNCONNECTED ;
  wire \NLW_blk00000547_ACOUT<5>_UNCONNECTED ;
  wire \NLW_blk00000547_ACOUT<4>_UNCONNECTED ;
  wire \NLW_blk00000547_ACOUT<3>_UNCONNECTED ;
  wire \NLW_blk00000547_ACOUT<2>_UNCONNECTED ;
  wire \NLW_blk00000547_ACOUT<1>_UNCONNECTED ;
  wire \NLW_blk00000547_ACOUT<0>_UNCONNECTED ;
  wire \NLW_blk00000547_CARRYOUT<3>_UNCONNECTED ;
  wire \NLW_blk00000547_CARRYOUT<2>_UNCONNECTED ;
  wire \NLW_blk00000547_CARRYOUT<1>_UNCONNECTED ;
  wire \NLW_blk00000547_CARRYOUT<0>_UNCONNECTED ;
  wire \NLW_blk00000547_BCOUT<17>_UNCONNECTED ;
  wire \NLW_blk00000547_BCOUT<16>_UNCONNECTED ;
  wire \NLW_blk00000547_BCOUT<15>_UNCONNECTED ;
  wire \NLW_blk00000547_BCOUT<14>_UNCONNECTED ;
  wire \NLW_blk00000547_BCOUT<13>_UNCONNECTED ;
  wire \NLW_blk00000547_BCOUT<12>_UNCONNECTED ;
  wire \NLW_blk00000547_BCOUT<11>_UNCONNECTED ;
  wire \NLW_blk00000547_BCOUT<10>_UNCONNECTED ;
  wire \NLW_blk00000547_BCOUT<9>_UNCONNECTED ;
  wire \NLW_blk00000547_BCOUT<8>_UNCONNECTED ;
  wire \NLW_blk00000547_BCOUT<7>_UNCONNECTED ;
  wire \NLW_blk00000547_BCOUT<6>_UNCONNECTED ;
  wire \NLW_blk00000547_BCOUT<5>_UNCONNECTED ;
  wire \NLW_blk00000547_BCOUT<4>_UNCONNECTED ;
  wire \NLW_blk00000547_BCOUT<3>_UNCONNECTED ;
  wire \NLW_blk00000547_BCOUT<2>_UNCONNECTED ;
  wire \NLW_blk00000547_BCOUT<1>_UNCONNECTED ;
  wire \NLW_blk00000547_BCOUT<0>_UNCONNECTED ;
  wire \NLW_blk00000547_P<47>_UNCONNECTED ;
  wire \NLW_blk00000547_P<46>_UNCONNECTED ;
  wire \NLW_blk00000547_P<45>_UNCONNECTED ;
  wire \NLW_blk00000547_P<44>_UNCONNECTED ;
  wire \NLW_blk00000547_P<43>_UNCONNECTED ;
  wire \NLW_blk00000547_PCOUT<47>_UNCONNECTED ;
  wire \NLW_blk00000547_PCOUT<46>_UNCONNECTED ;
  wire \NLW_blk00000547_PCOUT<45>_UNCONNECTED ;
  wire \NLW_blk00000547_PCOUT<44>_UNCONNECTED ;
  wire \NLW_blk00000547_PCOUT<43>_UNCONNECTED ;
  wire \NLW_blk00000547_PCOUT<42>_UNCONNECTED ;
  wire \NLW_blk00000547_PCOUT<41>_UNCONNECTED ;
  wire \NLW_blk00000547_PCOUT<40>_UNCONNECTED ;
  wire \NLW_blk00000547_PCOUT<39>_UNCONNECTED ;
  wire \NLW_blk00000547_PCOUT<38>_UNCONNECTED ;
  wire \NLW_blk00000547_PCOUT<37>_UNCONNECTED ;
  wire \NLW_blk00000547_PCOUT<36>_UNCONNECTED ;
  wire \NLW_blk00000547_PCOUT<35>_UNCONNECTED ;
  wire \NLW_blk00000547_PCOUT<34>_UNCONNECTED ;
  wire \NLW_blk00000547_PCOUT<33>_UNCONNECTED ;
  wire \NLW_blk00000547_PCOUT<32>_UNCONNECTED ;
  wire \NLW_blk00000547_PCOUT<31>_UNCONNECTED ;
  wire \NLW_blk00000547_PCOUT<30>_UNCONNECTED ;
  wire \NLW_blk00000547_PCOUT<29>_UNCONNECTED ;
  wire \NLW_blk00000547_PCOUT<28>_UNCONNECTED ;
  wire \NLW_blk00000547_PCOUT<27>_UNCONNECTED ;
  wire \NLW_blk00000547_PCOUT<26>_UNCONNECTED ;
  wire \NLW_blk00000547_PCOUT<25>_UNCONNECTED ;
  wire \NLW_blk00000547_PCOUT<24>_UNCONNECTED ;
  wire \NLW_blk00000547_PCOUT<23>_UNCONNECTED ;
  wire \NLW_blk00000547_PCOUT<22>_UNCONNECTED ;
  wire \NLW_blk00000547_PCOUT<21>_UNCONNECTED ;
  wire \NLW_blk00000547_PCOUT<20>_UNCONNECTED ;
  wire \NLW_blk00000547_PCOUT<19>_UNCONNECTED ;
  wire \NLW_blk00000547_PCOUT<18>_UNCONNECTED ;
  wire \NLW_blk00000547_PCOUT<17>_UNCONNECTED ;
  wire \NLW_blk00000547_PCOUT<16>_UNCONNECTED ;
  wire \NLW_blk00000547_PCOUT<15>_UNCONNECTED ;
  wire \NLW_blk00000547_PCOUT<14>_UNCONNECTED ;
  wire \NLW_blk00000547_PCOUT<13>_UNCONNECTED ;
  wire \NLW_blk00000547_PCOUT<12>_UNCONNECTED ;
  wire \NLW_blk00000547_PCOUT<11>_UNCONNECTED ;
  wire \NLW_blk00000547_PCOUT<10>_UNCONNECTED ;
  wire \NLW_blk00000547_PCOUT<9>_UNCONNECTED ;
  wire \NLW_blk00000547_PCOUT<8>_UNCONNECTED ;
  wire \NLW_blk00000547_PCOUT<7>_UNCONNECTED ;
  wire \NLW_blk00000547_PCOUT<6>_UNCONNECTED ;
  wire \NLW_blk00000547_PCOUT<5>_UNCONNECTED ;
  wire \NLW_blk00000547_PCOUT<4>_UNCONNECTED ;
  wire \NLW_blk00000547_PCOUT<3>_UNCONNECTED ;
  wire \NLW_blk00000547_PCOUT<2>_UNCONNECTED ;
  wire \NLW_blk00000547_PCOUT<1>_UNCONNECTED ;
  wire \NLW_blk00000547_PCOUT<0>_UNCONNECTED ;
  wire NLW_blk00000548_PATTERNBDETECT_UNCONNECTED;
  wire NLW_blk00000548_MULTSIGNOUT_UNCONNECTED;
  wire NLW_blk00000548_CARRYCASCOUT_UNCONNECTED;
  wire NLW_blk00000548_UNDERFLOW_UNCONNECTED;
  wire NLW_blk00000548_PATTERNDETECT_UNCONNECTED;
  wire NLW_blk00000548_OVERFLOW_UNCONNECTED;
  wire \NLW_blk00000548_ACOUT<29>_UNCONNECTED ;
  wire \NLW_blk00000548_ACOUT<28>_UNCONNECTED ;
  wire \NLW_blk00000548_ACOUT<27>_UNCONNECTED ;
  wire \NLW_blk00000548_ACOUT<26>_UNCONNECTED ;
  wire \NLW_blk00000548_ACOUT<25>_UNCONNECTED ;
  wire \NLW_blk00000548_ACOUT<24>_UNCONNECTED ;
  wire \NLW_blk00000548_ACOUT<23>_UNCONNECTED ;
  wire \NLW_blk00000548_ACOUT<22>_UNCONNECTED ;
  wire \NLW_blk00000548_ACOUT<21>_UNCONNECTED ;
  wire \NLW_blk00000548_ACOUT<20>_UNCONNECTED ;
  wire \NLW_blk00000548_ACOUT<19>_UNCONNECTED ;
  wire \NLW_blk00000548_ACOUT<18>_UNCONNECTED ;
  wire \NLW_blk00000548_ACOUT<17>_UNCONNECTED ;
  wire \NLW_blk00000548_ACOUT<16>_UNCONNECTED ;
  wire \NLW_blk00000548_ACOUT<15>_UNCONNECTED ;
  wire \NLW_blk00000548_ACOUT<14>_UNCONNECTED ;
  wire \NLW_blk00000548_ACOUT<13>_UNCONNECTED ;
  wire \NLW_blk00000548_ACOUT<12>_UNCONNECTED ;
  wire \NLW_blk00000548_ACOUT<11>_UNCONNECTED ;
  wire \NLW_blk00000548_ACOUT<10>_UNCONNECTED ;
  wire \NLW_blk00000548_ACOUT<9>_UNCONNECTED ;
  wire \NLW_blk00000548_ACOUT<8>_UNCONNECTED ;
  wire \NLW_blk00000548_ACOUT<7>_UNCONNECTED ;
  wire \NLW_blk00000548_ACOUT<6>_UNCONNECTED ;
  wire \NLW_blk00000548_ACOUT<5>_UNCONNECTED ;
  wire \NLW_blk00000548_ACOUT<4>_UNCONNECTED ;
  wire \NLW_blk00000548_ACOUT<3>_UNCONNECTED ;
  wire \NLW_blk00000548_ACOUT<2>_UNCONNECTED ;
  wire \NLW_blk00000548_ACOUT<1>_UNCONNECTED ;
  wire \NLW_blk00000548_ACOUT<0>_UNCONNECTED ;
  wire \NLW_blk00000548_CARRYOUT<3>_UNCONNECTED ;
  wire \NLW_blk00000548_CARRYOUT<2>_UNCONNECTED ;
  wire \NLW_blk00000548_CARRYOUT<1>_UNCONNECTED ;
  wire \NLW_blk00000548_CARRYOUT<0>_UNCONNECTED ;
  wire \NLW_blk00000548_BCOUT<17>_UNCONNECTED ;
  wire \NLW_blk00000548_BCOUT<16>_UNCONNECTED ;
  wire \NLW_blk00000548_BCOUT<15>_UNCONNECTED ;
  wire \NLW_blk00000548_BCOUT<14>_UNCONNECTED ;
  wire \NLW_blk00000548_BCOUT<13>_UNCONNECTED ;
  wire \NLW_blk00000548_BCOUT<12>_UNCONNECTED ;
  wire \NLW_blk00000548_BCOUT<11>_UNCONNECTED ;
  wire \NLW_blk00000548_BCOUT<10>_UNCONNECTED ;
  wire \NLW_blk00000548_BCOUT<9>_UNCONNECTED ;
  wire \NLW_blk00000548_BCOUT<8>_UNCONNECTED ;
  wire \NLW_blk00000548_BCOUT<7>_UNCONNECTED ;
  wire \NLW_blk00000548_BCOUT<6>_UNCONNECTED ;
  wire \NLW_blk00000548_BCOUT<5>_UNCONNECTED ;
  wire \NLW_blk00000548_BCOUT<4>_UNCONNECTED ;
  wire \NLW_blk00000548_BCOUT<3>_UNCONNECTED ;
  wire \NLW_blk00000548_BCOUT<2>_UNCONNECTED ;
  wire \NLW_blk00000548_BCOUT<1>_UNCONNECTED ;
  wire \NLW_blk00000548_BCOUT<0>_UNCONNECTED ;
  wire \NLW_blk00000548_P<47>_UNCONNECTED ;
  wire \NLW_blk00000548_P<46>_UNCONNECTED ;
  wire \NLW_blk00000548_P<45>_UNCONNECTED ;
  wire \NLW_blk00000548_P<44>_UNCONNECTED ;
  wire \NLW_blk00000548_P<43>_UNCONNECTED ;
  wire \NLW_blk00000548_PCOUT<47>_UNCONNECTED ;
  wire \NLW_blk00000548_PCOUT<46>_UNCONNECTED ;
  wire \NLW_blk00000548_PCOUT<45>_UNCONNECTED ;
  wire \NLW_blk00000548_PCOUT<44>_UNCONNECTED ;
  wire \NLW_blk00000548_PCOUT<43>_UNCONNECTED ;
  wire \NLW_blk00000548_PCOUT<42>_UNCONNECTED ;
  wire \NLW_blk00000548_PCOUT<41>_UNCONNECTED ;
  wire \NLW_blk00000548_PCOUT<40>_UNCONNECTED ;
  wire \NLW_blk00000548_PCOUT<39>_UNCONNECTED ;
  wire \NLW_blk00000548_PCOUT<38>_UNCONNECTED ;
  wire \NLW_blk00000548_PCOUT<37>_UNCONNECTED ;
  wire \NLW_blk00000548_PCOUT<36>_UNCONNECTED ;
  wire \NLW_blk00000548_PCOUT<35>_UNCONNECTED ;
  wire \NLW_blk00000548_PCOUT<34>_UNCONNECTED ;
  wire \NLW_blk00000548_PCOUT<33>_UNCONNECTED ;
  wire \NLW_blk00000548_PCOUT<32>_UNCONNECTED ;
  wire \NLW_blk00000548_PCOUT<31>_UNCONNECTED ;
  wire \NLW_blk00000548_PCOUT<30>_UNCONNECTED ;
  wire \NLW_blk00000548_PCOUT<29>_UNCONNECTED ;
  wire \NLW_blk00000548_PCOUT<28>_UNCONNECTED ;
  wire \NLW_blk00000548_PCOUT<27>_UNCONNECTED ;
  wire \NLW_blk00000548_PCOUT<26>_UNCONNECTED ;
  wire \NLW_blk00000548_PCOUT<25>_UNCONNECTED ;
  wire \NLW_blk00000548_PCOUT<24>_UNCONNECTED ;
  wire \NLW_blk00000548_PCOUT<23>_UNCONNECTED ;
  wire \NLW_blk00000548_PCOUT<22>_UNCONNECTED ;
  wire \NLW_blk00000548_PCOUT<21>_UNCONNECTED ;
  wire \NLW_blk00000548_PCOUT<20>_UNCONNECTED ;
  wire \NLW_blk00000548_PCOUT<19>_UNCONNECTED ;
  wire \NLW_blk00000548_PCOUT<18>_UNCONNECTED ;
  wire \NLW_blk00000548_PCOUT<17>_UNCONNECTED ;
  wire \NLW_blk00000548_PCOUT<16>_UNCONNECTED ;
  wire \NLW_blk00000548_PCOUT<15>_UNCONNECTED ;
  wire \NLW_blk00000548_PCOUT<14>_UNCONNECTED ;
  wire \NLW_blk00000548_PCOUT<13>_UNCONNECTED ;
  wire \NLW_blk00000548_PCOUT<12>_UNCONNECTED ;
  wire \NLW_blk00000548_PCOUT<11>_UNCONNECTED ;
  wire \NLW_blk00000548_PCOUT<10>_UNCONNECTED ;
  wire \NLW_blk00000548_PCOUT<9>_UNCONNECTED ;
  wire \NLW_blk00000548_PCOUT<8>_UNCONNECTED ;
  wire \NLW_blk00000548_PCOUT<7>_UNCONNECTED ;
  wire \NLW_blk00000548_PCOUT<6>_UNCONNECTED ;
  wire \NLW_blk00000548_PCOUT<5>_UNCONNECTED ;
  wire \NLW_blk00000548_PCOUT<4>_UNCONNECTED ;
  wire \NLW_blk00000548_PCOUT<3>_UNCONNECTED ;
  wire \NLW_blk00000548_PCOUT<2>_UNCONNECTED ;
  wire \NLW_blk00000548_PCOUT<1>_UNCONNECTED ;
  wire \NLW_blk00000548_PCOUT<0>_UNCONNECTED ;
  wire NLW_blk000005ef_Q_UNCONNECTED;
  wire NLW_blk000005f0_Q_UNCONNECTED;
  wire NLW_blk000005f1_Q_UNCONNECTED;
  wire NLW_blk000005f2_Q_UNCONNECTED;
  wire NLW_blk000005f3_Q_UNCONNECTED;
  wire NLW_blk000005f4_Q_UNCONNECTED;
  wire NLW_blk000005f5_Q_UNCONNECTED;
  wire NLW_blk000005f6_Q_UNCONNECTED;
  wire NLW_blk00000607_Q_UNCONNECTED;
  wire NLW_blk00000608_Q_UNCONNECTED;
  wire NLW_blk00000609_Q_UNCONNECTED;
  wire NLW_blk00000625_Q_UNCONNECTED;
  wire NLW_blk00000626_Q_UNCONNECTED;
  wire NLW_blk00000627_Q_UNCONNECTED;
  wire NLW_blk00000628_Q_UNCONNECTED;
  wire NLW_blk00000629_Q_UNCONNECTED;
  wire NLW_blk0000062a_Q_UNCONNECTED;
  wire NLW_blk0000062b_Q_UNCONNECTED;
  wire NLW_blk0000062c_Q_UNCONNECTED;
  wire NLW_blk0000063d_Q_UNCONNECTED;
  wire NLW_blk0000063e_Q_UNCONNECTED;
  wire NLW_blk0000063f_Q_UNCONNECTED;
  wire NLW_blk0000064e_Q_UNCONNECTED;
  wire NLW_blk0000064f_Q_UNCONNECTED;
  wire NLW_blk00000652_R_UNCONNECTED;
  wire NLW_blk000008ac_O_UNCONNECTED;
  wire NLW_blk000008d1_O_UNCONNECTED;
  wire NLW_blk000009c5_Q_UNCONNECTED;
  wire NLW_blk000009c6_Q_UNCONNECTED;
  wire NLW_blk000009c7_Q_UNCONNECTED;
  wire NLW_blk000009d8_Q_UNCONNECTED;
  wire NLW_blk000009d9_Q_UNCONNECTED;
  wire NLW_blk000009ef_Q_UNCONNECTED;
  wire NLW_blk000009f0_Q_UNCONNECTED;
  wire NLW_blk000009f1_Q_UNCONNECTED;
  wire NLW_blk00000a02_Q_UNCONNECTED;
  wire NLW_blk00000a03_Q_UNCONNECTED;
  wire NLW_blk00000a25_R_UNCONNECTED;
  wire NLW_blk00000a26_Q_UNCONNECTED;
  wire NLW_blk00000b84_Q15_UNCONNECTED;
  wire NLW_blk00000b86_Q15_UNCONNECTED;
  wire NLW_blk00000b88_Q15_UNCONNECTED;
  wire NLW_blk00000b8a_Q15_UNCONNECTED;
  wire NLW_blk00000b8c_Q15_UNCONNECTED;
  wire NLW_blk00000b8e_Q15_UNCONNECTED;
  wire NLW_blk00000b90_Q15_UNCONNECTED;
  wire NLW_blk00000b92_Q15_UNCONNECTED;
  wire NLW_blk00000b94_Q15_UNCONNECTED;
  wire NLW_blk00000b96_Q15_UNCONNECTED;
  wire NLW_blk00000b98_Q15_UNCONNECTED;
  wire NLW_blk00000b9a_Q15_UNCONNECTED;
  wire NLW_blk00000b9c_Q15_UNCONNECTED;
  wire NLW_blk00000b9e_Q15_UNCONNECTED;
  wire NLW_blk00000ba0_Q15_UNCONNECTED;
  wire NLW_blk00000ba2_Q15_UNCONNECTED;
  wire NLW_blk00000ba4_Q15_UNCONNECTED;
  wire NLW_blk00000ba6_Q15_UNCONNECTED;
  wire NLW_blk00000ba8_Q15_UNCONNECTED;
  wire NLW_blk00000baa_Q15_UNCONNECTED;
  wire NLW_blk00000bac_Q15_UNCONNECTED;
  wire NLW_blk00000bae_Q15_UNCONNECTED;
  wire NLW_blk00000bb0_Q15_UNCONNECTED;
  wire NLW_blk00000bb2_Q15_UNCONNECTED;
  wire NLW_blk00000bb4_Q15_UNCONNECTED;
  wire NLW_blk00000bb6_Q15_UNCONNECTED;
  wire NLW_blk00000bb8_Q15_UNCONNECTED;
  wire NLW_blk00000bba_Q15_UNCONNECTED;
  wire NLW_blk00000bbc_Q15_UNCONNECTED;
  wire NLW_blk00000bbe_Q15_UNCONNECTED;
  wire NLW_blk00000bc0_Q15_UNCONNECTED;
  wire NLW_blk00000bc2_Q15_UNCONNECTED;
  wire NLW_blk00000bc4_Q15_UNCONNECTED;
  wire NLW_blk00000bc6_Q15_UNCONNECTED;
  wire NLW_blk00000bc8_Q15_UNCONNECTED;
  wire NLW_blk00000bca_Q15_UNCONNECTED;
  wire NLW_blk00000bcc_Q15_UNCONNECTED;
  wire NLW_blk00000bce_Q15_UNCONNECTED;
  wire NLW_blk00000bd0_Q15_UNCONNECTED;
  wire NLW_blk00000bd2_Q15_UNCONNECTED;
  wire NLW_blk00000bd4_Q15_UNCONNECTED;
  wire NLW_blk00000bd6_Q15_UNCONNECTED;
  wire NLW_blk00000bd8_Q15_UNCONNECTED;
  wire NLW_blk00000bda_Q15_UNCONNECTED;
  wire NLW_blk00000bdc_Q15_UNCONNECTED;
  wire NLW_blk00000bde_Q15_UNCONNECTED;
  wire NLW_blk00000be0_Q15_UNCONNECTED;
  wire NLW_blk00000be2_Q15_UNCONNECTED;
  wire NLW_blk00000be4_Q15_UNCONNECTED;
  wire NLW_blk00000be6_Q15_UNCONNECTED;
  wire NLW_blk00000be8_Q15_UNCONNECTED;
  wire NLW_blk00000bea_Q15_UNCONNECTED;
  wire NLW_blk00000bec_Q15_UNCONNECTED;
  wire NLW_blk00000bee_Q15_UNCONNECTED;
  wire NLW_blk00000bf0_Q15_UNCONNECTED;
  wire NLW_blk00000bf2_Q15_UNCONNECTED;
  wire NLW_blk00000bf4_Q15_UNCONNECTED;
  wire NLW_blk00000bf6_Q15_UNCONNECTED;
  wire NLW_blk00000bf8_Q15_UNCONNECTED;
  wire NLW_blk00000bfa_Q15_UNCONNECTED;
  wire NLW_blk00000bfc_Q15_UNCONNECTED;
  wire NLW_blk00000bfe_Q15_UNCONNECTED;
  wire NLW_blk00000c00_Q15_UNCONNECTED;
  wire NLW_blk00000c02_Q15_UNCONNECTED;
  wire NLW_blk00000c04_Q15_UNCONNECTED;
  wire NLW_blk00000c06_Q15_UNCONNECTED;
  wire NLW_blk00000c08_Q15_UNCONNECTED;
  wire NLW_blk00000c0a_Q15_UNCONNECTED;
  wire NLW_blk00000c0c_Q15_UNCONNECTED;
  wire \NLW_blk000000dc/blk000000df_Q15_UNCONNECTED ;
  wire \NLW_blk000001f6/blk000001f9_Q15_UNCONNECTED ;
  wire \NLW_blk000002a3/blk000002a8_Q31_UNCONNECTED ;
  wire \NLW_blk000002a3/blk000002a6_Q31_UNCONNECTED ;
  wire \NLW_blk000002aa/blk000002ad_Q31_UNCONNECTED ;
  wire \NLW_blk000002af/blk000002b2_Q15_UNCONNECTED ;
  wire \NLW_blk000002b4/blk000002b7_Q31_UNCONNECTED ;
  wire \NLW_blk000002b9/blk000002be_Q31_UNCONNECTED ;
  wire \NLW_blk000002b9/blk000002bc_Q31_UNCONNECTED ;
  wire \NLW_blk000002c0/blk000002c5_Q31_UNCONNECTED ;
  wire \NLW_blk000002c0/blk000002c3_Q31_UNCONNECTED ;
  wire \NLW_blk000003fc/blk000003fe_Q15_UNCONNECTED ;
  wire \NLW_blk00000400/blk00000402_Q15_UNCONNECTED ;
  wire \NLW_blk00000404/blk00000407_Q15_UNCONNECTED ;
  wire \NLW_blk00000503/blk00000506_Q15_UNCONNECTED ;
  wire \NLW_blk00000508/blk0000050a_Q15_UNCONNECTED ;
  wire \NLW_blk00000522/blk00000544_Q15_UNCONNECTED ;
  wire \NLW_blk00000522/blk00000542_Q15_UNCONNECTED ;
  wire \NLW_blk00000640/blk00000643_Q15_UNCONNECTED ;
  wire \NLW_blk00000659/blk0000065b_Q15_UNCONNECTED ;
  wire \NLW_blk000007cb/blk000007ce_Q15_UNCONNECTED ;
  wire \NLW_blk0000083a/blk0000083c_Q15_UNCONNECTED ;
  wire \NLW_blk0000083e/blk00000840_Q15_UNCONNECTED ;
  wire [36 : 0] \U0/i_synth/axi_wrapper/data_out_channel/data_out ;
  wire [0 : 0] \U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer ;
  wire [1 : 1] \NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer ;
  assign
    m_axis_data_tdata[31] = \U0/i_synth/axi_wrapper/data_out_channel/data_out [32],
    m_axis_data_tdata[30] = \U0/i_synth/axi_wrapper/data_out_channel/data_out [31],
    m_axis_data_tdata[29] = \U0/i_synth/axi_wrapper/data_out_channel/data_out [30],
    m_axis_data_tdata[28] = \U0/i_synth/axi_wrapper/data_out_channel/data_out [29],
    m_axis_data_tdata[27] = \U0/i_synth/axi_wrapper/data_out_channel/data_out [28],
    m_axis_data_tdata[26] = \U0/i_synth/axi_wrapper/data_out_channel/data_out [27],
    m_axis_data_tdata[25] = \U0/i_synth/axi_wrapper/data_out_channel/data_out [26],
    m_axis_data_tdata[24] = \U0/i_synth/axi_wrapper/data_out_channel/data_out [25],
    m_axis_data_tdata[23] = \U0/i_synth/axi_wrapper/data_out_channel/data_out [24],
    m_axis_data_tdata[22] = \U0/i_synth/axi_wrapper/data_out_channel/data_out [23],
    m_axis_data_tdata[21] = \U0/i_synth/axi_wrapper/data_out_channel/data_out [22],
    m_axis_data_tdata[20] = \U0/i_synth/axi_wrapper/data_out_channel/data_out [21],
    m_axis_data_tdata[19] = \U0/i_synth/axi_wrapper/data_out_channel/data_out [20],
    m_axis_data_tdata[18] = \U0/i_synth/axi_wrapper/data_out_channel/data_out [19],
    m_axis_data_tdata[17] = \U0/i_synth/axi_wrapper/data_out_channel/data_out [18],
    m_axis_data_tdata[16] = \U0/i_synth/axi_wrapper/data_out_channel/data_out [17],
    m_axis_data_tdata[15] = \U0/i_synth/axi_wrapper/data_out_channel/data_out [16],
    m_axis_data_tdata[14] = \U0/i_synth/axi_wrapper/data_out_channel/data_out [15],
    m_axis_data_tdata[13] = \U0/i_synth/axi_wrapper/data_out_channel/data_out [14],
    m_axis_data_tdata[12] = \U0/i_synth/axi_wrapper/data_out_channel/data_out [13],
    m_axis_data_tdata[11] = \U0/i_synth/axi_wrapper/data_out_channel/data_out [12],
    m_axis_data_tdata[10] = \U0/i_synth/axi_wrapper/data_out_channel/data_out [11],
    m_axis_data_tdata[9] = \U0/i_synth/axi_wrapper/data_out_channel/data_out [10],
    m_axis_data_tdata[8] = \U0/i_synth/axi_wrapper/data_out_channel/data_out [9],
    m_axis_data_tdata[7] = \U0/i_synth/axi_wrapper/data_out_channel/data_out [8],
    m_axis_data_tdata[6] = \U0/i_synth/axi_wrapper/data_out_channel/data_out [7],
    m_axis_data_tdata[5] = \U0/i_synth/axi_wrapper/data_out_channel/data_out [6],
    m_axis_data_tdata[4] = \U0/i_synth/axi_wrapper/data_out_channel/data_out [5],
    m_axis_data_tdata[3] = \U0/i_synth/axi_wrapper/data_out_channel/data_out [4],
    m_axis_data_tdata[2] = \U0/i_synth/axi_wrapper/data_out_channel/data_out [3],
    m_axis_data_tdata[1] = \U0/i_synth/axi_wrapper/data_out_channel/data_out [2],
    m_axis_data_tdata[0] = \U0/i_synth/axi_wrapper/data_out_channel/data_out [1],
    m_axis_data_tuser[7] = \NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
    m_axis_data_tuser[6] = \NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
    m_axis_data_tuser[5] = \NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
    m_axis_data_tuser[4] = \NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
    m_axis_data_tuser[3] = \U0/i_synth/axi_wrapper/data_out_channel/data_out [36],
    m_axis_data_tuser[2] = \U0/i_synth/axi_wrapper/data_out_channel/data_out [35],
    m_axis_data_tuser[1] = \U0/i_synth/axi_wrapper/data_out_channel/data_out [34],
    m_axis_data_tuser[0] = \U0/i_synth/axi_wrapper/data_out_channel/data_out [33],
    m_axis_data_tvalid = \NlwRenamedSig_OI_U0/i_synth/axi_wrapper/dv_resolved_prev ,
    m_axis_data_tlast = \U0/i_synth/axi_wrapper/data_out_channel/data_out [0],
    event_frame_started = \U0/i_synth/axi_wrapper/event_frame_started ,
    event_tlast_unexpected = \U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [0],
    event_tlast_missing = \U0/i_synth/axi_wrapper/event_tlast_missing ,
    event_data_in_channel_halt = \U0/i_synth/axi_wrapper/event_data_in_channel_halt_int ;
  VCC   blk00000001 (
    .P(sig00000344)
  );
  GND   blk00000002 (
    .G(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1])
  );
  FDR #(
    .INIT ( 1'b0 ))
  blk00000003 (
    .C(aclk),
    .D(sig00000054),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(\U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [0])
  );
  FDR   blk00000004 (
    .C(aclk),
    .D(sig0000006d),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig0000006a)
  );
  FDR   blk00000005 (
    .C(aclk),
    .D(sig0000002c),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000069)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000006 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000005e),
    .Q(sig00000065)
  );
  FDR #(
    .INIT ( 1'b0 ))
  blk00000007 (
    .C(aclk),
    .D(sig00000061),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(\U0/i_synth/axi_wrapper/event_data_in_channel_halt_int )
  );
  FDR #(
    .INIT ( 1'b0 ))
  blk00000008 (
    .C(aclk),
    .D(sig0000005d),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000066)
  );
  FDR #(
    .INIT ( 1'b0 ))
  blk00000009 (
    .C(aclk),
    .D(sig0000002d),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000067)
  );
  FDS #(
    .INIT ( 1'b1 ))
  blk0000000a (
    .C(aclk),
    .D(sig0000005a),
    .S(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000068)
  );
  FDR #(
    .INIT ( 1'b0 ))
  blk0000000b (
    .C(aclk),
    .D(sig0000005b),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(\U0/i_synth/axi_wrapper/event_tlast_missing )
  );
  FDR #(
    .INIT ( 1'b0 ))
  blk0000000c (
    .C(aclk),
    .D(sig00000059),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(\U0/i_synth/axi_wrapper/event_frame_started )
  );
  FDR #(
    .INIT ( 1'b0 ))
  blk0000000d (
    .C(aclk),
    .D(sig00000001),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/dv_resolved_prev )
  );
  FDR #(
    .INIT ( 1'b0 ))
  blk0000000e (
    .C(aclk),
    .D(sig0000005f),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig0000002c)
  );
  FDE   blk0000000f (
    .C(aclk),
    .CE(sig0000006c),
    .D(s_axis_config_tdata[4]),
    .Q(sig00000031)
  );
  FDE   blk00000010 (
    .C(aclk),
    .CE(sig0000006c),
    .D(s_axis_config_tdata[3]),
    .Q(sig00000030)
  );
  FDE   blk00000011 (
    .C(aclk),
    .CE(sig0000006c),
    .D(s_axis_config_tdata[2]),
    .Q(sig0000002f)
  );
  FDE   blk00000012 (
    .C(aclk),
    .CE(sig0000006c),
    .D(s_axis_config_tdata[1]),
    .Q(sig0000002e)
  );
  FDE   blk00000013 (
    .C(aclk),
    .CE(sig0000006c),
    .D(s_axis_config_tdata[0]),
    .Q(sig0000002b)
  );
  FDE   blk00000014 (
    .C(aclk),
    .CE(sig0000006e),
    .D(s_axis_data_tdata[31]),
    .Q(sig00000041)
  );
  FDE   blk00000015 (
    .C(aclk),
    .CE(sig0000006e),
    .D(s_axis_data_tdata[30]),
    .Q(sig00000040)
  );
  FDE   blk00000016 (
    .C(aclk),
    .CE(sig0000006e),
    .D(s_axis_data_tdata[29]),
    .Q(sig0000003f)
  );
  FDE   blk00000017 (
    .C(aclk),
    .CE(sig0000006e),
    .D(s_axis_data_tdata[28]),
    .Q(sig0000003e)
  );
  FDE   blk00000018 (
    .C(aclk),
    .CE(sig0000006e),
    .D(s_axis_data_tdata[27]),
    .Q(sig0000003d)
  );
  FDE   blk00000019 (
    .C(aclk),
    .CE(sig0000006e),
    .D(s_axis_data_tdata[26]),
    .Q(sig0000003c)
  );
  FDE   blk0000001a (
    .C(aclk),
    .CE(sig0000006e),
    .D(s_axis_data_tdata[25]),
    .Q(sig0000003b)
  );
  FDE   blk0000001b (
    .C(aclk),
    .CE(sig0000006e),
    .D(s_axis_data_tdata[24]),
    .Q(sig0000003a)
  );
  FDE   blk0000001c (
    .C(aclk),
    .CE(sig0000006e),
    .D(s_axis_data_tdata[23]),
    .Q(sig00000039)
  );
  FDE   blk0000001d (
    .C(aclk),
    .CE(sig0000006e),
    .D(s_axis_data_tdata[22]),
    .Q(sig00000038)
  );
  FDE   blk0000001e (
    .C(aclk),
    .CE(sig0000006e),
    .D(s_axis_data_tdata[21]),
    .Q(sig00000037)
  );
  FDE   blk0000001f (
    .C(aclk),
    .CE(sig0000006e),
    .D(s_axis_data_tdata[20]),
    .Q(sig00000036)
  );
  FDE   blk00000020 (
    .C(aclk),
    .CE(sig0000006e),
    .D(s_axis_data_tdata[19]),
    .Q(sig00000035)
  );
  FDE   blk00000021 (
    .C(aclk),
    .CE(sig0000006e),
    .D(s_axis_data_tdata[18]),
    .Q(sig00000034)
  );
  FDE   blk00000022 (
    .C(aclk),
    .CE(sig0000006e),
    .D(s_axis_data_tdata[17]),
    .Q(sig00000033)
  );
  FDE   blk00000023 (
    .C(aclk),
    .CE(sig0000006e),
    .D(s_axis_data_tdata[16]),
    .Q(sig00000032)
  );
  FDE   blk00000024 (
    .C(aclk),
    .CE(sig0000006e),
    .D(s_axis_data_tdata[15]),
    .Q(sig00000051)
  );
  FDE   blk00000025 (
    .C(aclk),
    .CE(sig0000006e),
    .D(s_axis_data_tdata[14]),
    .Q(sig00000050)
  );
  FDE   blk00000026 (
    .C(aclk),
    .CE(sig0000006e),
    .D(s_axis_data_tdata[13]),
    .Q(sig0000004f)
  );
  FDE   blk00000027 (
    .C(aclk),
    .CE(sig0000006e),
    .D(s_axis_data_tdata[12]),
    .Q(sig0000004e)
  );
  FDE   blk00000028 (
    .C(aclk),
    .CE(sig0000006e),
    .D(s_axis_data_tdata[11]),
    .Q(sig0000004d)
  );
  FDE   blk00000029 (
    .C(aclk),
    .CE(sig0000006e),
    .D(s_axis_data_tdata[10]),
    .Q(sig0000004c)
  );
  FDE   blk0000002a (
    .C(aclk),
    .CE(sig0000006e),
    .D(s_axis_data_tdata[9]),
    .Q(sig0000004b)
  );
  FDE   blk0000002b (
    .C(aclk),
    .CE(sig0000006e),
    .D(s_axis_data_tdata[8]),
    .Q(sig0000004a)
  );
  FDE   blk0000002c (
    .C(aclk),
    .CE(sig0000006e),
    .D(s_axis_data_tdata[7]),
    .Q(sig00000049)
  );
  FDE   blk0000002d (
    .C(aclk),
    .CE(sig0000006e),
    .D(s_axis_data_tdata[6]),
    .Q(sig00000048)
  );
  FDE   blk0000002e (
    .C(aclk),
    .CE(sig0000006e),
    .D(s_axis_data_tdata[5]),
    .Q(sig00000047)
  );
  FDE   blk0000002f (
    .C(aclk),
    .CE(sig0000006e),
    .D(s_axis_data_tdata[4]),
    .Q(sig00000046)
  );
  FDE   blk00000030 (
    .C(aclk),
    .CE(sig0000006e),
    .D(s_axis_data_tdata[3]),
    .Q(sig00000045)
  );
  FDE   blk00000031 (
    .C(aclk),
    .CE(sig0000006e),
    .D(s_axis_data_tdata[2]),
    .Q(sig00000044)
  );
  FDE   blk00000032 (
    .C(aclk),
    .CE(sig0000006e),
    .D(s_axis_data_tdata[1]),
    .Q(sig00000043)
  );
  FDE   blk00000033 (
    .C(aclk),
    .CE(sig0000006e),
    .D(s_axis_data_tdata[0]),
    .Q(sig00000042)
  );
  FDE   blk00000034 (
    .C(aclk),
    .CE(sig0000006e),
    .D(s_axis_data_tlast),
    .Q(sig0000006b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000035 (
    .C(aclk),
    .CE(sig00000001),
    .D(sig00000026),
    .Q(\U0/i_synth/axi_wrapper/data_out_channel/data_out [36])
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000036 (
    .C(aclk),
    .CE(sig00000001),
    .D(sig00000025),
    .Q(\U0/i_synth/axi_wrapper/data_out_channel/data_out [35])
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000037 (
    .C(aclk),
    .CE(sig00000001),
    .D(sig00000024),
    .Q(\U0/i_synth/axi_wrapper/data_out_channel/data_out [34])
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000038 (
    .C(aclk),
    .CE(sig00000001),
    .D(sig00000023),
    .Q(\U0/i_synth/axi_wrapper/data_out_channel/data_out [33])
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000039 (
    .C(aclk),
    .CE(sig00000001),
    .D(sig00000012),
    .Q(\U0/i_synth/axi_wrapper/data_out_channel/data_out [32])
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000003a (
    .C(aclk),
    .CE(sig00000001),
    .D(sig00000011),
    .Q(\U0/i_synth/axi_wrapper/data_out_channel/data_out [31])
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000003b (
    .C(aclk),
    .CE(sig00000001),
    .D(sig00000010),
    .Q(\U0/i_synth/axi_wrapper/data_out_channel/data_out [30])
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000003c (
    .C(aclk),
    .CE(sig00000001),
    .D(sig0000000f),
    .Q(\U0/i_synth/axi_wrapper/data_out_channel/data_out [29])
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000003d (
    .C(aclk),
    .CE(sig00000001),
    .D(sig0000000e),
    .Q(\U0/i_synth/axi_wrapper/data_out_channel/data_out [28])
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000003e (
    .C(aclk),
    .CE(sig00000001),
    .D(sig0000000d),
    .Q(\U0/i_synth/axi_wrapper/data_out_channel/data_out [27])
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000003f (
    .C(aclk),
    .CE(sig00000001),
    .D(sig0000000c),
    .Q(\U0/i_synth/axi_wrapper/data_out_channel/data_out [26])
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000040 (
    .C(aclk),
    .CE(sig00000001),
    .D(sig0000000b),
    .Q(\U0/i_synth/axi_wrapper/data_out_channel/data_out [25])
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000041 (
    .C(aclk),
    .CE(sig00000001),
    .D(sig0000000a),
    .Q(\U0/i_synth/axi_wrapper/data_out_channel/data_out [24])
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000042 (
    .C(aclk),
    .CE(sig00000001),
    .D(sig00000009),
    .Q(\U0/i_synth/axi_wrapper/data_out_channel/data_out [23])
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000043 (
    .C(aclk),
    .CE(sig00000001),
    .D(sig00000008),
    .Q(\U0/i_synth/axi_wrapper/data_out_channel/data_out [22])
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000044 (
    .C(aclk),
    .CE(sig00000001),
    .D(sig00000007),
    .Q(\U0/i_synth/axi_wrapper/data_out_channel/data_out [21])
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000045 (
    .C(aclk),
    .CE(sig00000001),
    .D(sig00000006),
    .Q(\U0/i_synth/axi_wrapper/data_out_channel/data_out [20])
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000046 (
    .C(aclk),
    .CE(sig00000001),
    .D(sig00000005),
    .Q(\U0/i_synth/axi_wrapper/data_out_channel/data_out [19])
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000047 (
    .C(aclk),
    .CE(sig00000001),
    .D(sig00000004),
    .Q(\U0/i_synth/axi_wrapper/data_out_channel/data_out [18])
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000048 (
    .C(aclk),
    .CE(sig00000001),
    .D(sig00000003),
    .Q(\U0/i_synth/axi_wrapper/data_out_channel/data_out [17])
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000049 (
    .C(aclk),
    .CE(sig00000001),
    .D(sig00000022),
    .Q(\U0/i_synth/axi_wrapper/data_out_channel/data_out [16])
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000004a (
    .C(aclk),
    .CE(sig00000001),
    .D(sig00000021),
    .Q(\U0/i_synth/axi_wrapper/data_out_channel/data_out [15])
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000004b (
    .C(aclk),
    .CE(sig00000001),
    .D(sig00000020),
    .Q(\U0/i_synth/axi_wrapper/data_out_channel/data_out [14])
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000004c (
    .C(aclk),
    .CE(sig00000001),
    .D(sig0000001f),
    .Q(\U0/i_synth/axi_wrapper/data_out_channel/data_out [13])
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000004d (
    .C(aclk),
    .CE(sig00000001),
    .D(sig0000001e),
    .Q(\U0/i_synth/axi_wrapper/data_out_channel/data_out [12])
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000004e (
    .C(aclk),
    .CE(sig00000001),
    .D(sig0000001d),
    .Q(\U0/i_synth/axi_wrapper/data_out_channel/data_out [11])
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000004f (
    .C(aclk),
    .CE(sig00000001),
    .D(sig0000001c),
    .Q(\U0/i_synth/axi_wrapper/data_out_channel/data_out [10])
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000050 (
    .C(aclk),
    .CE(sig00000001),
    .D(sig0000001b),
    .Q(\U0/i_synth/axi_wrapper/data_out_channel/data_out [9])
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000051 (
    .C(aclk),
    .CE(sig00000001),
    .D(sig0000001a),
    .Q(\U0/i_synth/axi_wrapper/data_out_channel/data_out [8])
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000052 (
    .C(aclk),
    .CE(sig00000001),
    .D(sig00000019),
    .Q(\U0/i_synth/axi_wrapper/data_out_channel/data_out [7])
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000053 (
    .C(aclk),
    .CE(sig00000001),
    .D(sig00000018),
    .Q(\U0/i_synth/axi_wrapper/data_out_channel/data_out [6])
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000054 (
    .C(aclk),
    .CE(sig00000001),
    .D(sig00000017),
    .Q(\U0/i_synth/axi_wrapper/data_out_channel/data_out [5])
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000055 (
    .C(aclk),
    .CE(sig00000001),
    .D(sig00000016),
    .Q(\U0/i_synth/axi_wrapper/data_out_channel/data_out [4])
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000056 (
    .C(aclk),
    .CE(sig00000001),
    .D(sig00000015),
    .Q(\U0/i_synth/axi_wrapper/data_out_channel/data_out [3])
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000057 (
    .C(aclk),
    .CE(sig00000001),
    .D(sig00000014),
    .Q(\U0/i_synth/axi_wrapper/data_out_channel/data_out [2])
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000058 (
    .C(aclk),
    .CE(sig00000001),
    .D(sig00000013),
    .Q(\U0/i_synth/axi_wrapper/data_out_channel/data_out [1])
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000059 (
    .C(aclk),
    .CE(sig00000001),
    .D(sig00000060),
    .Q(\U0/i_synth/axi_wrapper/data_out_channel/data_out [0])
  );
  LUT3 #(
    .INIT ( 8'hAE ))
  blk0000005a (
    .I0(sig00000070),
    .I1(sig000000c4),
    .I2(sig00000072),
    .O(sig00000073)
  );
  MUXCY   blk0000005b (
    .CI(sig00000344),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig00000075),
    .O(sig00000074)
  );
  XORCY   blk0000005c (
    .CI(sig00000079),
    .LI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .O(sig00000077)
  );
  MUXCY   blk0000005d (
    .CI(sig00000344),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig0000007a),
    .O(sig00000078)
  );
  MUXCY   blk0000005e (
    .CI(sig00000078),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig0000007b),
    .O(sig00000079)
  );
  LUT6 #(
    .INIT ( 64'h9009000000009009 ))
  blk0000005f (
    .I0(sig000000c8),
    .I1(sig00000344),
    .I2(sig000000c7),
    .I3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .I4(sig000000c6),
    .I5(sig00000344),
    .O(sig0000007a)
  );
  LUT6 #(
    .INIT ( 64'h9009000000009009 ))
  blk00000060 (
    .I0(sig000000c5),
    .I1(sig00000344),
    .I2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .I3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .I4(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .I5(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .O(sig0000007b)
  );
  FDR #(
    .INIT ( 1'b0 ))
  blk00000061 (
    .C(aclk),
    .D(sig000000c4),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000001)
  );
  FDR #(
    .INIT ( 1'b0 ))
  blk00000062 (
    .C(aclk),
    .D(sig00000070),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(NLW_blk00000062_Q_UNCONNECTED)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000063 (
    .C(aclk),
    .D(sig000000ca),
    .Q(sig00000071)
  );
  FDR #(
    .INIT ( 1'b0 ))
  blk00000064 (
    .C(aclk),
    .D(sig00000071),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000000c2)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000065 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000073),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000000c4)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000066 (
    .C(aclk),
    .CE(sig000000c4),
    .D(sig00000077),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000076)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000067 (
    .C(aclk),
    .CE(sig000000c4),
    .D(sig00000076),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000072)
  );
  FDR #(
    .INIT ( 1'b0 ))
  blk00000068 (
    .C(aclk),
    .D(sig000000c8),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000026)
  );
  FDR #(
    .INIT ( 1'b0 ))
  blk00000069 (
    .C(aclk),
    .D(sig000000c7),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000025)
  );
  FDR #(
    .INIT ( 1'b0 ))
  blk0000006a (
    .C(aclk),
    .D(sig000000c6),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000024)
  );
  FDR #(
    .INIT ( 1'b0 ))
  blk0000006b (
    .C(aclk),
    .D(sig000000c5),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000023)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000006c (
    .A0(sig00000344),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000041),
    .Q(sig000000ef)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000006d (
    .A0(sig00000344),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000040),
    .Q(sig000000f0)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000006e (
    .A0(sig00000344),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig0000003f),
    .Q(sig000000f1)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000006f (
    .A0(sig00000344),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig0000003e),
    .Q(sig000000f2)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000070 (
    .A0(sig00000344),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig0000003d),
    .Q(sig000000f3)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000071 (
    .A0(sig00000344),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig0000003c),
    .Q(sig000000f4)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000072 (
    .A0(sig00000344),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig0000003b),
    .Q(sig000000f5)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000073 (
    .A0(sig00000344),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig0000003a),
    .Q(sig000000f6)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000074 (
    .A0(sig00000344),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000039),
    .Q(sig000000f7)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000075 (
    .A0(sig00000344),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000038),
    .Q(sig000000f8)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000076 (
    .A0(sig00000344),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000037),
    .Q(sig000000f9)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000077 (
    .A0(sig00000344),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000036),
    .Q(sig000000fa)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000078 (
    .A0(sig00000344),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000035),
    .Q(sig000000fb)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000079 (
    .A0(sig00000344),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000034),
    .Q(sig000000fc)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000007a (
    .A0(sig00000344),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000033),
    .Q(sig000000fd)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000007b (
    .A0(sig00000344),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000032),
    .Q(sig000000fe)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000007c (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000000ef),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000000de)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000007d (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000000f0),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000000dd)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000007e (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000000f1),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000000dc)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000007f (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000000f2),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000000db)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000080 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000000f3),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000000da)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000081 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000000f4),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000000d9)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000082 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000000f5),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000000d8)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000083 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000000f6),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000000d7)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000084 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000000f7),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000000d6)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000085 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000000f8),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000000d5)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000086 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000000f9),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000000d4)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000087 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000000fa),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000000d3)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000088 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000000fb),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000000d2)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000089 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000000fc),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000000d1)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000008a (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000000fd),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000000d0)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000008b (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000000fe),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000000cf)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000008c (
    .A0(sig00000344),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000051),
    .Q(sig000000ff)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000008d (
    .A0(sig00000344),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000050),
    .Q(sig00000100)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000008e (
    .A0(sig00000344),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig0000004f),
    .Q(sig00000101)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000008f (
    .A0(sig00000344),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig0000004e),
    .Q(sig00000102)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000090 (
    .A0(sig00000344),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig0000004d),
    .Q(sig00000103)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000091 (
    .A0(sig00000344),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig0000004c),
    .Q(sig00000104)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000092 (
    .A0(sig00000344),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig0000004b),
    .Q(sig00000105)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000093 (
    .A0(sig00000344),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig0000004a),
    .Q(sig00000106)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000094 (
    .A0(sig00000344),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000049),
    .Q(sig00000107)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000095 (
    .A0(sig00000344),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000048),
    .Q(sig00000108)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000096 (
    .A0(sig00000344),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000047),
    .Q(sig00000109)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000097 (
    .A0(sig00000344),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000046),
    .Q(sig0000010a)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000098 (
    .A0(sig00000344),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000045),
    .Q(sig0000010b)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000099 (
    .A0(sig00000344),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000044),
    .Q(sig0000010c)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000009a (
    .A0(sig00000344),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000043),
    .Q(sig0000010d)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000009b (
    .A0(sig00000344),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000042),
    .Q(sig0000010e)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000009c (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000000ff),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000000ee)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000009d (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000100),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000000ed)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000009e (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000101),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000000ec)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000009f (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000102),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000000eb)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000000a0 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000103),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000000ea)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000000a1 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000104),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000000e9)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000000a2 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000105),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000000e8)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000000a3 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000106),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000000e7)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000000a4 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000107),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000000e6)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000000a5 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000108),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000000e5)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000000a6 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000109),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000000e4)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000000a7 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000010a),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000000e3)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000000a8 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000010b),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000000e2)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000000a9 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000010c),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000000e1)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000000aa (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000010d),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000000e0)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000000ab (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000010e),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000000df)
  );
  LUT6 #(
    .INIT ( 64'h9009000000009009 ))
  blk000000ac (
    .I0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .I1(sig0000002a),
    .I2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .I3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .I4(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .I5(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .O(sig0000010f)
  );
  LUT6 #(
    .INIT ( 64'h9009000000009009 ))
  blk000000ad (
    .I0(sig00000344),
    .I1(sig00000027),
    .I2(sig00000344),
    .I3(sig00000028),
    .I4(sig00000344),
    .I5(sig00000029),
    .O(sig00000110)
  );
  MUXCY   blk000000ae (
    .CI(sig00000112),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig0000010f),
    .O(sig00000111)
  );
  MUXCY   blk000000af (
    .CI(sig00000344),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig00000110),
    .O(sig00000112)
  );
  XORCY   blk000000b0 (
    .CI(sig00000111),
    .LI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .O(sig0000011b)
  );
  LUT6 #(
    .INIT ( 64'h9009000000009009 ))
  blk000000b1 (
    .I0(sig0000002a),
    .I1(sig00000344),
    .I2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .I3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .I4(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .I5(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .O(sig00000113)
  );
  LUT6 #(
    .INIT ( 64'h9009000000009009 ))
  blk000000b2 (
    .I0(sig00000027),
    .I1(sig00000344),
    .I2(sig00000028),
    .I3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .I4(sig00000029),
    .I5(sig00000344),
    .O(sig00000114)
  );
  MUXCY   blk000000b3 (
    .CI(sig00000116),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig00000113),
    .O(sig00000115)
  );
  MUXCY   blk000000b4 (
    .CI(sig00000344),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig00000114),
    .O(sig00000116)
  );
  XORCY   blk000000b5 (
    .CI(sig00000115),
    .LI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .O(sig00000117)
  );
  MUXCY   blk000000b6 (
    .CI(sig00000344),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig00000119),
    .O(sig0000011a)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000000b7 (
    .C(aclk),
    .CE(sig00000002),
    .D(sig00000118),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000121)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000000b8 (
    .C(aclk),
    .CE(sig00000002),
    .D(sig00000117),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000118)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000000b9 (
    .C(aclk),
    .D(sig0000011b),
    .Q(sig000000ca)
  );
  FDE #(
    .INIT ( 1'b1 ))
  blk000000ba (
    .C(aclk),
    .CE(sig00000120),
    .D(sig0000011e),
    .Q(sig000000c9)
  );
  FDE #(
    .INIT ( 1'b1 ))
  blk000000bb (
    .C(aclk),
    .CE(sig00000120),
    .D(sig00000125),
    .Q(sig000000ce)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000bc (
    .C(aclk),
    .CE(sig00000120),
    .D(sig00000124),
    .Q(sig000000cd)
  );
  FDE #(
    .INIT ( 1'b1 ))
  blk000000bd (
    .C(aclk),
    .CE(sig00000120),
    .D(sig00000123),
    .Q(sig000000cc)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000be (
    .C(aclk),
    .CE(sig00000120),
    .D(sig00000122),
    .Q(sig000000cb)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000bf (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000011c),
    .Q(sig00000002)
  );
  FDE #(
    .INIT ( 1'b1 ))
  blk000000c0 (
    .C(aclk),
    .CE(sig0000002c),
    .D(sig0000002b),
    .Q(sig0000011e)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000000c1 (
    .C(aclk),
    .D(sig0000011d),
    .Q(sig0000011f)
  );
  FDE #(
    .INIT ( 1'b1 ))
  blk000000c2 (
    .C(aclk),
    .CE(sig0000002c),
    .D(sig00000031),
    .Q(sig00000125)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000c3 (
    .C(aclk),
    .CE(sig0000002c),
    .D(sig00000030),
    .Q(sig00000124)
  );
  FDE #(
    .INIT ( 1'b1 ))
  blk000000c4 (
    .C(aclk),
    .CE(sig0000002c),
    .D(sig0000002f),
    .Q(sig00000123)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000c5 (
    .C(aclk),
    .CE(sig0000002c),
    .D(sig0000002e),
    .Q(sig00000122)
  );
  XORCY   blk000000c6 (
    .CI(sig0000012d),
    .LI(sig0000012b),
    .O(sig00000126)
  );
  XORCY   blk000000c7 (
    .CI(sig0000012e),
    .LI(sig00000c4f),
    .O(sig00000127)
  );
  XORCY   blk000000c8 (
    .CI(sig00000130),
    .LI(sig00000c50),
    .O(sig00000128)
  );
  MUXCY   blk000000c9 (
    .CI(sig0000012e),
    .DI(sig00000129),
    .S(sig00000c4f),
    .O(sig0000012d)
  );
  MUXCY   blk000000ca (
    .CI(sig00000130),
    .DI(sig0000012a),
    .S(sig00000c50),
    .O(sig0000012e)
  );
  XORCY   blk000000cb (
    .CI(sig0000011a),
    .LI(sig00000c51),
    .O(sig0000012f)
  );
  MUXCY   blk000000cc (
    .CI(sig0000011a),
    .DI(sig0000012c),
    .S(sig00000c51),
    .O(sig00000130)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000000cd (
    .C(aclk),
    .CE(sig00000002),
    .D(sig0000012f),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000027)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000000ce (
    .C(aclk),
    .CE(sig00000002),
    .D(sig00000128),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000028)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000000cf (
    .C(aclk),
    .CE(sig00000002),
    .D(sig00000127),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000029)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000000d0 (
    .C(aclk),
    .CE(sig00000002),
    .D(sig00000126),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig0000002a)
  );
  XORCY   blk000000d1 (
    .CI(sig00000138),
    .LI(sig00000136),
    .O(sig00000131)
  );
  XORCY   blk000000d2 (
    .CI(sig00000139),
    .LI(sig00000c52),
    .O(sig00000132)
  );
  XORCY   blk000000d3 (
    .CI(sig0000013b),
    .LI(sig00000c53),
    .O(sig00000133)
  );
  MUXCY   blk000000d4 (
    .CI(sig00000139),
    .DI(sig00000134),
    .S(sig00000c52),
    .O(sig00000138)
  );
  MUXCY   blk000000d5 (
    .CI(sig0000013b),
    .DI(sig00000135),
    .S(sig00000c53),
    .O(sig00000139)
  );
  XORCY   blk000000d6 (
    .CI(sig00000074),
    .LI(sig00000c54),
    .O(sig0000013a)
  );
  MUXCY   blk000000d7 (
    .CI(sig00000074),
    .DI(sig00000137),
    .S(sig00000c54),
    .O(sig0000013b)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000000d8 (
    .C(aclk),
    .CE(sig000000c4),
    .D(sig0000013a),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000000c8)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000000d9 (
    .C(aclk),
    .CE(sig000000c4),
    .D(sig00000133),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000000c7)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000000da (
    .C(aclk),
    .CE(sig000000c4),
    .D(sig00000132),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000000c6)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000000db (
    .C(aclk),
    .CE(sig000000c4),
    .D(sig00000131),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000000c5)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000000e1 (
    .A0(sig00000344),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig0000002a),
    .Q(sig0000013c)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000000e2 (
    .A0(sig00000344),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000029),
    .Q(sig0000013d)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000000e3 (
    .A0(sig00000344),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000028),
    .Q(sig0000013e)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000000e4 (
    .A0(sig00000344),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000027),
    .Q(sig0000013f)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000000e5 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000013c),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000000c3)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000000e6 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000013d),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(NLW_blk000000e6_Q_UNCONNECTED)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000000e7 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000013e),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(NLW_blk000000e7_Q_UNCONNECTED)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000000e8 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000013f),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(NLW_blk000000e8_Q_UNCONNECTED)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000000e9 (
    .C(aclk),
    .CE(sig00000151),
    .D(sig0000014a),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000208)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000000ea (
    .C(aclk),
    .CE(sig00000151),
    .D(sig00000149),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000207)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000000eb (
    .C(aclk),
    .CE(sig00000151),
    .D(sig00000148),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000206)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000000ec (
    .C(aclk),
    .CE(sig00000151),
    .D(sig00000141),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000205)
  );
  MUXCY   blk000000ed (
    .CI(sig00000156),
    .DI(sig00000144),
    .S(sig00000c55),
    .O(sig00000140)
  );
  XORCY   blk000000ee (
    .CI(sig00000156),
    .LI(sig00000c55),
    .O(sig00000141)
  );
  MUXCY   blk000000ef (
    .CI(sig00000140),
    .DI(sig00000146),
    .S(sig00000c56),
    .O(sig00000142)
  );
  MUXCY   blk000000f0 (
    .CI(sig00000142),
    .DI(sig00000147),
    .S(sig00000c57),
    .O(sig00000143)
  );
  XORCY   blk000000f1 (
    .CI(sig00000140),
    .LI(sig00000c56),
    .O(sig00000148)
  );
  XORCY   blk000000f2 (
    .CI(sig00000142),
    .LI(sig00000c57),
    .O(sig00000149)
  );
  XORCY   blk000000f3 (
    .CI(sig00000143),
    .LI(sig00000145),
    .O(sig0000014a)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000000f4 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(sig00000344),
    .A3(sig00000344),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000205),
    .Q(sig0000014b)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000000f5 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(sig00000344),
    .A3(sig00000344),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000206),
    .Q(sig0000014c)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000000f6 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(sig00000344),
    .A3(sig00000344),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000207),
    .Q(sig0000014d)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000000f7 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(sig00000344),
    .A3(sig00000344),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000208),
    .Q(sig0000014e)
  );
  LUT3 #(
    .INIT ( 8'hAE ))
  blk000000f8 (
    .I0(sig00000209),
    .I1(sig00000151),
    .I2(sig00000150),
    .O(sig00000152)
  );
  MUXCY   blk000000f9 (
    .CI(sig00000153),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig00000c58),
    .O(sig00000154)
  );
  XORCY   blk000000fa (
    .CI(sig00000154),
    .LI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .O(sig00000155)
  );
  MUXCY   blk000000fb (
    .CI(sig00000344),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig00000157),
    .O(sig00000156)
  );
  XORCY   blk000000fc (
    .CI(sig0000015b),
    .LI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .O(sig00000159)
  );
  MUXCY   blk000000fd (
    .CI(sig00000344),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig0000015c),
    .O(sig0000015a)
  );
  MUXCY   blk000000fe (
    .CI(sig0000015a),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig0000015d),
    .O(sig0000015b)
  );
  LUT6 #(
    .INIT ( 64'h9009000000009009 ))
  blk000000ff (
    .I0(sig00000205),
    .I1(sig00000344),
    .I2(sig00000206),
    .I3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .I4(sig00000207),
    .I5(sig00000344),
    .O(sig0000015c)
  );
  LUT6 #(
    .INIT ( 64'h9009000000009009 ))
  blk00000100 (
    .I0(sig00000208),
    .I1(sig00000344),
    .I2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .I3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .I4(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .I5(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .O(sig0000015d)
  );
  MUXCY   blk00000101 (
    .CI(sig00000344),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig0000015f),
    .O(sig0000015e)
  );
  MUXCY   blk00000102 (
    .CI(sig0000015e),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig00000160),
    .O(sig00000153)
  );
  LUT6 #(
    .INIT ( 64'h9009000000009009 ))
  blk00000103 (
    .I0(sig00000205),
    .I1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .I2(sig00000206),
    .I3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .I4(sig00000207),
    .I5(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .O(sig0000015f)
  );
  LUT6 #(
    .INIT ( 64'h9009000000009009 ))
  blk00000104 (
    .I0(sig00000208),
    .I1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .I2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .I3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .I4(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .I5(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .O(sig00000160)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000105 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000014b),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000001b2)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000106 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000014c),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000001b3)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000107 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000014d),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000001b0)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000108 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000014e),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000001b1)
  );
  FDR #(
    .INIT ( 1'b0 ))
  blk00000109 (
    .C(aclk),
    .D(sig0000014f),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig0000009d)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000010a (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000152),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000151)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000010b (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000155),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000204)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000010c (
    .C(aclk),
    .CE(sig00000151),
    .D(sig00000159),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000158)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000010d (
    .C(aclk),
    .CE(sig00000151),
    .D(sig00000158),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000150)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000010e (
    .C(aclk),
    .CE(sig00000209),
    .D(sig000000cb),
    .Q(sig000001dc)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000010f (
    .C(aclk),
    .CE(sig00000209),
    .D(sig000000cc),
    .Q(sig000001dd)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000110 (
    .C(aclk),
    .CE(sig00000209),
    .D(sig000000cd),
    .Q(sig000001de)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000111 (
    .C(aclk),
    .CE(sig00000209),
    .D(sig000000ce),
    .Q(sig000001df)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000112 (
    .C(aclk),
    .D(sig00000161),
    .Q(sig000001e1)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000113 (
    .C(aclk),
    .CE(sig00000209),
    .D(sig000001e1),
    .Q(sig00000162)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000114 (
    .C(aclk),
    .CE(sig00000228),
    .D(sig00000218),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig0000020d)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000115 (
    .C(aclk),
    .CE(sig00000228),
    .D(sig00000217),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig0000020c)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000116 (
    .C(aclk),
    .CE(sig00000228),
    .D(sig00000216),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig0000020b)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000117 (
    .C(aclk),
    .CE(sig00000228),
    .D(sig0000020f),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig0000020a)
  );
  MUXCY   blk00000118 (
    .CI(sig00000223),
    .DI(sig00000212),
    .S(sig00000c59),
    .O(sig0000020e)
  );
  XORCY   blk00000119 (
    .CI(sig00000223),
    .LI(sig00000c59),
    .O(sig0000020f)
  );
  MUXCY   blk0000011a (
    .CI(sig0000020e),
    .DI(sig00000214),
    .S(sig00000c5a),
    .O(sig00000210)
  );
  MUXCY   blk0000011b (
    .CI(sig00000210),
    .DI(sig00000215),
    .S(sig00000c5b),
    .O(sig00000211)
  );
  XORCY   blk0000011c (
    .CI(sig0000020e),
    .LI(sig00000c5a),
    .O(sig00000216)
  );
  XORCY   blk0000011d (
    .CI(sig00000210),
    .LI(sig00000c5b),
    .O(sig00000217)
  );
  XORCY   blk0000011e (
    .CI(sig00000211),
    .LI(sig00000213),
    .O(sig00000218)
  );
  LUT6 #(
    .INIT ( 64'h9009000000009009 ))
  blk0000011f (
    .I0(sig0000020d),
    .I1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .I2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .I3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .I4(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .I5(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .O(sig00000219)
  );
  LUT6 #(
    .INIT ( 64'h9009000000009009 ))
  blk00000120 (
    .I0(sig0000020a),
    .I1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .I2(sig0000020b),
    .I3(sig00000344),
    .I4(sig0000020c),
    .I5(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .O(sig0000021a)
  );
  MUXCY   blk00000121 (
    .CI(sig0000021b),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig00000219),
    .O(sig00000226)
  );
  MUXCY   blk00000122 (
    .CI(sig00000344),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig0000021a),
    .O(sig0000021b)
  );
  LUT6 #(
    .INIT ( 64'h9009000000009009 ))
  blk00000123 (
    .I0(sig0000020d),
    .I1(sig00000344),
    .I2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .I3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .I4(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .I5(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .O(sig0000021c)
  );
  LUT6 #(
    .INIT ( 64'h9009000000009009 ))
  blk00000124 (
    .I0(sig0000020a),
    .I1(sig00000344),
    .I2(sig0000020b),
    .I3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .I4(sig0000020c),
    .I5(sig00000344),
    .O(sig0000021d)
  );
  MUXCY   blk00000125 (
    .CI(sig0000021f),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig0000021c),
    .O(sig0000021e)
  );
  MUXCY   blk00000126 (
    .CI(sig00000344),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig0000021d),
    .O(sig0000021f)
  );
  XORCY   blk00000127 (
    .CI(sig0000021e),
    .LI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .O(sig00000220)
  );
  MUXCY   blk00000128 (
    .CI(sig00000344),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig00000222),
    .O(sig00000223)
  );
  XORCY   blk00000129 (
    .CI(sig00000225),
    .LI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .O(sig00000224)
  );
  MUXCY   blk0000012a (
    .CI(sig00000226),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig00000c5c),
    .O(sig00000225)
  );
  LUT3 #(
    .INIT ( 8'hAE ))
  blk0000012b (
    .I0(sig000000c2),
    .I1(sig00000228),
    .I2(sig00000229),
    .O(sig00000227)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000012c (
    .C(aclk),
    .CE(sig00000228),
    .D(sig00000221),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000229)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000012d (
    .C(aclk),
    .CE(sig00000228),
    .D(sig00000220),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000221)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000012e (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000224),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000209)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000012f (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000227),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000228)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000130 (
    .I0(sig0000029f),
    .I1(sig0000027d),
    .I2(sig000002c0),
    .O(sig0000022a)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000131 (
    .I0(sig000002a0),
    .I1(sig0000027e),
    .I2(sig000002c0),
    .O(sig0000022b)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000132 (
    .I0(sig000002a1),
    .I1(sig0000027f),
    .I2(sig000002c0),
    .O(sig0000022c)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000133 (
    .I0(sig000002a2),
    .I1(sig00000280),
    .I2(sig000002c0),
    .O(sig0000022d)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000134 (
    .I0(sig000002a3),
    .I1(sig00000281),
    .I2(sig000002c0),
    .O(sig0000022e)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000135 (
    .I0(sig000002a4),
    .I1(sig00000282),
    .I2(sig000002c0),
    .O(sig0000022f)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000136 (
    .I0(sig000002a5),
    .I1(sig00000283),
    .I2(sig000002c0),
    .O(sig00000230)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000137 (
    .I0(sig000002a6),
    .I1(sig00000284),
    .I2(sig000002c0),
    .O(sig00000231)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000138 (
    .I0(sig000002a7),
    .I1(sig00000285),
    .I2(sig000002c0),
    .O(sig00000232)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000139 (
    .I0(sig000002a8),
    .I1(sig00000286),
    .I2(sig000002c0),
    .O(sig00000233)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk0000013a (
    .I0(sig000002a9),
    .I1(sig00000287),
    .I2(sig000002c0),
    .O(sig00000234)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk0000013b (
    .I0(sig000002aa),
    .I1(sig00000288),
    .I2(sig000002c0),
    .O(sig00000235)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk0000013c (
    .I0(sig000002ab),
    .I1(sig00000289),
    .I2(sig000002c0),
    .O(sig00000236)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk0000013d (
    .I0(sig000002ac),
    .I1(sig0000028a),
    .I2(sig000002c0),
    .O(sig00000237)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk0000013e (
    .I0(sig000002ad),
    .I1(sig0000028b),
    .I2(sig000002c0),
    .O(sig00000238)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk0000013f (
    .I0(sig000002ae),
    .I1(sig0000028c),
    .I2(sig000002c0),
    .O(sig00000239)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000140 (
    .I0(sig000002af),
    .I1(sig0000028d),
    .I2(sig000002c0),
    .O(sig0000023a)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000141 (
    .I0(sig0000027d),
    .I1(sig0000029f),
    .I2(sig000002c0),
    .O(sig0000023b)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000142 (
    .I0(sig0000027e),
    .I1(sig000002a0),
    .I2(sig000002c0),
    .O(sig0000023c)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000143 (
    .I0(sig0000027f),
    .I1(sig000002a1),
    .I2(sig000002c0),
    .O(sig0000023d)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000144 (
    .I0(sig00000280),
    .I1(sig000002a2),
    .I2(sig000002c0),
    .O(sig0000023e)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000145 (
    .I0(sig00000281),
    .I1(sig000002a3),
    .I2(sig000002c0),
    .O(sig0000023f)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000146 (
    .I0(sig00000282),
    .I1(sig000002a4),
    .I2(sig000002c0),
    .O(sig00000240)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000147 (
    .I0(sig00000283),
    .I1(sig000002a5),
    .I2(sig000002c0),
    .O(sig00000241)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000148 (
    .I0(sig00000284),
    .I1(sig000002a6),
    .I2(sig000002c0),
    .O(sig00000242)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000149 (
    .I0(sig00000285),
    .I1(sig000002a7),
    .I2(sig000002c0),
    .O(sig00000243)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk0000014a (
    .I0(sig00000286),
    .I1(sig000002a8),
    .I2(sig000002c0),
    .O(sig00000244)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk0000014b (
    .I0(sig00000287),
    .I1(sig000002a9),
    .I2(sig000002c0),
    .O(sig00000245)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk0000014c (
    .I0(sig00000288),
    .I1(sig000002aa),
    .I2(sig000002c0),
    .O(sig00000246)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk0000014d (
    .I0(sig00000289),
    .I1(sig000002ab),
    .I2(sig000002c0),
    .O(sig00000247)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk0000014e (
    .I0(sig0000028a),
    .I1(sig000002ac),
    .I2(sig000002c0),
    .O(sig00000248)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk0000014f (
    .I0(sig0000028b),
    .I1(sig000002ad),
    .I2(sig000002c0),
    .O(sig00000249)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000150 (
    .I0(sig0000028c),
    .I1(sig000002ae),
    .I2(sig000002c0),
    .O(sig0000024a)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000151 (
    .I0(sig0000028d),
    .I1(sig000002af),
    .I2(sig000002c0),
    .O(sig0000024b)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000152 (
    .I0(sig000000df),
    .I1(sig000002c3),
    .I2(sig000000c3),
    .O(sig0000024c)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000153 (
    .I0(sig000000e0),
    .I1(sig000002c4),
    .I2(sig000000c3),
    .O(sig0000024d)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000154 (
    .I0(sig000000e1),
    .I1(sig000002c5),
    .I2(sig000000c3),
    .O(sig0000024e)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000155 (
    .I0(sig000000e2),
    .I1(sig000002c6),
    .I2(sig000000c3),
    .O(sig0000024f)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000156 (
    .I0(sig000000e3),
    .I1(sig000002c7),
    .I2(sig000000c3),
    .O(sig00000250)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000157 (
    .I0(sig000000e4),
    .I1(sig000002c8),
    .I2(sig000000c3),
    .O(sig00000251)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000158 (
    .I0(sig000000e5),
    .I1(sig000002c9),
    .I2(sig000000c3),
    .O(sig00000252)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000159 (
    .I0(sig000000e6),
    .I1(sig000002ca),
    .I2(sig000000c3),
    .O(sig00000253)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk0000015a (
    .I0(sig000000e7),
    .I1(sig000002cb),
    .I2(sig000000c3),
    .O(sig00000254)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk0000015b (
    .I0(sig000000e8),
    .I1(sig000002cc),
    .I2(sig000000c3),
    .O(sig00000255)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk0000015c (
    .I0(sig000000e9),
    .I1(sig000002cd),
    .I2(sig000000c3),
    .O(sig00000256)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk0000015d (
    .I0(sig000000ea),
    .I1(sig000002ce),
    .I2(sig000000c3),
    .O(sig00000257)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk0000015e (
    .I0(sig000000eb),
    .I1(sig000002cf),
    .I2(sig000000c3),
    .O(sig00000258)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk0000015f (
    .I0(sig000000ec),
    .I1(sig000002d0),
    .I2(sig000000c3),
    .O(sig00000259)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000160 (
    .I0(sig000000ed),
    .I1(sig000002d1),
    .I2(sig000000c3),
    .O(sig0000025a)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000161 (
    .I0(sig000000ee),
    .I1(sig000002d2),
    .I2(sig000000c3),
    .O(sig0000025b)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000162 (
    .I0(sig000002c3),
    .I1(sig000000df),
    .I2(sig000000c3),
    .O(sig0000025c)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000163 (
    .I0(sig000002c4),
    .I1(sig000000e0),
    .I2(sig000000c3),
    .O(sig0000025d)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000164 (
    .I0(sig000002c5),
    .I1(sig000000e1),
    .I2(sig000000c3),
    .O(sig0000025e)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000165 (
    .I0(sig000002c6),
    .I1(sig000000e2),
    .I2(sig000000c3),
    .O(sig0000025f)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000166 (
    .I0(sig000002c7),
    .I1(sig000000e3),
    .I2(sig000000c3),
    .O(sig00000260)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000167 (
    .I0(sig000002c8),
    .I1(sig000000e4),
    .I2(sig000000c3),
    .O(sig00000261)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000168 (
    .I0(sig000002c9),
    .I1(sig000000e5),
    .I2(sig000000c3),
    .O(sig00000262)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000169 (
    .I0(sig000002ca),
    .I1(sig000000e6),
    .I2(sig000000c3),
    .O(sig00000263)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk0000016a (
    .I0(sig000002cb),
    .I1(sig000000e7),
    .I2(sig000000c3),
    .O(sig00000264)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk0000016b (
    .I0(sig000002cc),
    .I1(sig000000e8),
    .I2(sig000000c3),
    .O(sig00000265)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk0000016c (
    .I0(sig000002cd),
    .I1(sig000000e9),
    .I2(sig000000c3),
    .O(sig00000266)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk0000016d (
    .I0(sig000002ce),
    .I1(sig000000ea),
    .I2(sig000000c3),
    .O(sig00000267)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk0000016e (
    .I0(sig000002cf),
    .I1(sig000000eb),
    .I2(sig000000c3),
    .O(sig00000268)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk0000016f (
    .I0(sig000002d0),
    .I1(sig000000ec),
    .I2(sig000000c3),
    .O(sig00000269)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000170 (
    .I0(sig000002d1),
    .I1(sig000000ed),
    .I2(sig000000c3),
    .O(sig0000026a)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000171 (
    .I0(sig000002d2),
    .I1(sig000000ee),
    .I2(sig000000c3),
    .O(sig0000026b)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000172 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000022a),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig0000026c)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000173 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000022b),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig0000026d)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000174 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000022c),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig0000026e)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000175 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000022d),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig0000026f)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000176 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000022e),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000270)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000177 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000022f),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000271)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000178 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000230),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000272)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000179 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000231),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000273)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000017a (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000232),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000274)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000017b (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000233),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000275)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000017c (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000234),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000276)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000017d (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000235),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000277)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000017e (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000236),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000278)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000017f (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000237),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000279)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000180 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000238),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig0000027a)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000181 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000239),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig0000027b)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000182 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000023a),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig0000027c)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000183 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000023b),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000001e2)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000184 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000023c),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000001e3)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000185 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000023d),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000001e4)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000186 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000023e),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000001e5)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000187 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000023f),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000001e6)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000188 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000240),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000001e7)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000189 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000241),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000001e8)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000018a (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000242),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000001e9)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000018b (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000243),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000001ea)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000018c (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000244),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000001eb)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000018d (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000245),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000001ec)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000018e (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000246),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000001ed)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000018f (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000247),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000001ee)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000190 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000248),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000001ef)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000191 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000249),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000001f0)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000192 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000024a),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000001f1)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000193 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000024b),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000001f2)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000194 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000002c2),
    .Q(sig000002c1)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000195 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000024c),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000002e3)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000196 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000024d),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000002e4)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000197 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000024e),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000002e5)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000198 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000024f),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000002e6)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000199 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000250),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000002e7)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000019a (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000251),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000002e8)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000019b (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000252),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000002e9)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000019c (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000253),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000002ea)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000019d (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000254),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000002eb)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000019e (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000255),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000002ec)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000019f (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000256),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000002ed)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000001a0 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000257),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000002ee)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000001a1 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000258),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000002ef)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000001a2 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000259),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000002f0)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000001a3 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000025a),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000002f1)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000001a4 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000025b),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000002f2)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000001a5 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000025c),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000002d3)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000001a6 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000025d),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000002d4)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000001a7 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000025e),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000002d5)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000001a8 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000025f),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000002d6)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000001a9 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000260),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000002d7)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000001aa (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000261),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000002d8)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000001ab (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000262),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000002d9)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000001ac (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000263),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000002da)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000001ad (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000264),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000002db)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000001ae (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000265),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000002dc)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000001af (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000266),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000002dd)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000001b0 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000267),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000002de)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000001b1 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000268),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000002df)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000001b2 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000269),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000002e0)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000001b3 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000026a),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000002e1)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000001b4 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000026b),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000002e2)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001b5 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000000c3),
    .Q(sig000002c2)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000001b6 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(sig00000344),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000002f2),
    .Q(sig000002f3)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000001b7 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(sig00000344),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000002f1),
    .Q(sig000002f4)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000001b8 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(sig00000344),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000002f0),
    .Q(sig000002f5)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000001b9 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(sig00000344),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000002ef),
    .Q(sig000002f6)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000001ba (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(sig00000344),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000002ee),
    .Q(sig000002f7)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000001bb (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(sig00000344),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000002ed),
    .Q(sig000002f8)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000001bc (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(sig00000344),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000002ec),
    .Q(sig000002f9)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000001bd (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(sig00000344),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000002eb),
    .Q(sig000002fa)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000001be (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(sig00000344),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000002ea),
    .Q(sig000002fb)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000001bf (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(sig00000344),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000002e9),
    .Q(sig000002fc)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000001c0 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(sig00000344),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000002e8),
    .Q(sig000002fd)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000001c1 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(sig00000344),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000002e7),
    .Q(sig000002fe)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000001c2 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(sig00000344),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000002e6),
    .Q(sig000002ff)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000001c3 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(sig00000344),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000002e5),
    .Q(sig00000300)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000001c4 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(sig00000344),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000002e4),
    .Q(sig00000301)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000001c5 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(sig00000344),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000002e3),
    .Q(sig00000302)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000001c6 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000002f3),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000002bf)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000001c7 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000002f4),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000002be)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000001c8 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000002f5),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000002bd)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000001c9 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000002f6),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000002bc)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000001ca (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000002f7),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000002bb)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000001cb (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000002f8),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000002ba)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000001cc (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000002f9),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000002b9)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000001cd (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000002fa),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000002b8)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000001ce (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000002fb),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000002b7)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000001cf (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000002fc),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000002b6)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000001d0 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000002fd),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000002b5)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000001d1 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000002fe),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000002b4)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000001d2 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000002ff),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000002b3)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000001d3 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000300),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000002b2)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000001d4 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000301),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000002b1)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000001d5 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000302),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000002b0)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000001d6 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(sig00000344),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000000de),
    .Q(sig00000303)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000001d7 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(sig00000344),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000000dd),
    .Q(sig00000304)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000001d8 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(sig00000344),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000000dc),
    .Q(sig00000305)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000001d9 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(sig00000344),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000000db),
    .Q(sig00000306)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000001da (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(sig00000344),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000000da),
    .Q(sig00000307)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000001db (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(sig00000344),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000000d9),
    .Q(sig00000308)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000001dc (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(sig00000344),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000000d8),
    .Q(sig00000309)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000001dd (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(sig00000344),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000000d7),
    .Q(sig0000030a)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000001de (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(sig00000344),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000000d6),
    .Q(sig0000030b)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000001df (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(sig00000344),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000000d5),
    .Q(sig0000030c)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000001e0 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(sig00000344),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000000d4),
    .Q(sig0000030d)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000001e1 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(sig00000344),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000000d3),
    .Q(sig0000030e)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000001e2 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(sig00000344),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000000d2),
    .Q(sig0000030f)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000001e3 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(sig00000344),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000000d1),
    .Q(sig00000310)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000001e4 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(sig00000344),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000000d0),
    .Q(sig00000311)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000001e5 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(sig00000344),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000000cf),
    .Q(sig00000312)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000001e6 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000303),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000002d2)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000001e7 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000304),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000002d1)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000001e8 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000305),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000002d0)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000001e9 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000306),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000002cf)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000001ea (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000307),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000002ce)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000001eb (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000308),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000002cd)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000001ec (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000309),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000002cc)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000001ed (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000030a),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000002cb)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000001ee (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000030b),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000002ca)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000001ef (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000030c),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000002c9)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000001f0 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000030d),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000002c8)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000001f1 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000030e),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000002c7)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000001f2 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000030f),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000002c6)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000001f3 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000310),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000002c5)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000001f4 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000311),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000002c4)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000001f5 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000312),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000002c3)
  );
  XORCY   blk000001fb (
    .CI(sig00000334),
    .LI(sig00000324),
    .O(sig00000313)
  );
  XORCY   blk000001fc (
    .CI(sig00000335),
    .LI(sig00000c5d),
    .O(sig00000314)
  );
  XORCY   blk000001fd (
    .CI(sig00000336),
    .LI(sig00000325),
    .O(sig00000315)
  );
  XORCY   blk000001fe (
    .CI(sig00000337),
    .LI(sig00000326),
    .O(sig00000316)
  );
  XORCY   blk000001ff (
    .CI(sig00000338),
    .LI(sig00000327),
    .O(sig00000317)
  );
  XORCY   blk00000200 (
    .CI(sig00000339),
    .LI(sig00000328),
    .O(sig00000318)
  );
  XORCY   blk00000201 (
    .CI(sig0000033a),
    .LI(sig00000329),
    .O(sig00000319)
  );
  XORCY   blk00000202 (
    .CI(sig0000033b),
    .LI(sig0000032a),
    .O(sig0000031a)
  );
  XORCY   blk00000203 (
    .CI(sig0000033c),
    .LI(sig0000032b),
    .O(sig0000031b)
  );
  XORCY   blk00000204 (
    .CI(sig0000033d),
    .LI(sig0000032c),
    .O(sig0000031c)
  );
  XORCY   blk00000205 (
    .CI(sig0000033e),
    .LI(sig0000032d),
    .O(sig0000031d)
  );
  XORCY   blk00000206 (
    .CI(sig0000033f),
    .LI(sig0000032e),
    .O(sig0000031e)
  );
  XORCY   blk00000207 (
    .CI(sig00000340),
    .LI(sig0000032f),
    .O(sig0000031f)
  );
  XORCY   blk00000208 (
    .CI(sig00000341),
    .LI(sig00000330),
    .O(sig00000320)
  );
  XORCY   blk00000209 (
    .CI(sig00000342),
    .LI(sig00000331),
    .O(sig00000321)
  );
  XORCY   blk0000020a (
    .CI(sig00000343),
    .LI(sig00000332),
    .O(sig00000322)
  );
  XORCY   blk0000020b (
    .CI(sig00000344),
    .LI(sig00000333),
    .O(sig00000323)
  );
  MUXCY   blk0000020c (
    .CI(sig00000335),
    .DI(sig000002bf),
    .S(sig00000c5d),
    .O(sig00000334)
  );
  MUXCY   blk0000020d (
    .CI(sig00000336),
    .DI(sig000002be),
    .S(sig00000325),
    .O(sig00000335)
  );
  MUXCY   blk0000020e (
    .CI(sig00000337),
    .DI(sig000002bd),
    .S(sig00000326),
    .O(sig00000336)
  );
  MUXCY   blk0000020f (
    .CI(sig00000338),
    .DI(sig000002bc),
    .S(sig00000327),
    .O(sig00000337)
  );
  MUXCY   blk00000210 (
    .CI(sig00000339),
    .DI(sig000002bb),
    .S(sig00000328),
    .O(sig00000338)
  );
  MUXCY   blk00000211 (
    .CI(sig0000033a),
    .DI(sig000002ba),
    .S(sig00000329),
    .O(sig00000339)
  );
  MUXCY   blk00000212 (
    .CI(sig0000033b),
    .DI(sig000002b9),
    .S(sig0000032a),
    .O(sig0000033a)
  );
  MUXCY   blk00000213 (
    .CI(sig0000033c),
    .DI(sig000002b8),
    .S(sig0000032b),
    .O(sig0000033b)
  );
  MUXCY   blk00000214 (
    .CI(sig0000033d),
    .DI(sig000002b7),
    .S(sig0000032c),
    .O(sig0000033c)
  );
  MUXCY   blk00000215 (
    .CI(sig0000033e),
    .DI(sig000002b6),
    .S(sig0000032d),
    .O(sig0000033d)
  );
  MUXCY   blk00000216 (
    .CI(sig0000033f),
    .DI(sig000002b5),
    .S(sig0000032e),
    .O(sig0000033e)
  );
  MUXCY   blk00000217 (
    .CI(sig00000340),
    .DI(sig000002b4),
    .S(sig0000032f),
    .O(sig0000033f)
  );
  MUXCY   blk00000218 (
    .CI(sig00000341),
    .DI(sig000002b3),
    .S(sig00000330),
    .O(sig00000340)
  );
  MUXCY   blk00000219 (
    .CI(sig00000342),
    .DI(sig000002b2),
    .S(sig00000331),
    .O(sig00000341)
  );
  MUXCY   blk0000021a (
    .CI(sig00000343),
    .DI(sig000002b1),
    .S(sig00000332),
    .O(sig00000342)
  );
  MUXCY   blk0000021b (
    .CI(sig00000344),
    .DI(sig000002b0),
    .S(sig00000333),
    .O(sig00000343)
  );
  XORCY   blk0000021c (
    .CI(sig00000366),
    .LI(sig00000356),
    .O(sig00000345)
  );
  XORCY   blk0000021d (
    .CI(sig00000367),
    .LI(sig00000c5e),
    .O(sig00000346)
  );
  XORCY   blk0000021e (
    .CI(sig00000368),
    .LI(sig00000357),
    .O(sig00000347)
  );
  XORCY   blk0000021f (
    .CI(sig00000369),
    .LI(sig00000358),
    .O(sig00000348)
  );
  XORCY   blk00000220 (
    .CI(sig0000036a),
    .LI(sig00000359),
    .O(sig00000349)
  );
  XORCY   blk00000221 (
    .CI(sig0000036b),
    .LI(sig0000035a),
    .O(sig0000034a)
  );
  XORCY   blk00000222 (
    .CI(sig0000036c),
    .LI(sig0000035b),
    .O(sig0000034b)
  );
  XORCY   blk00000223 (
    .CI(sig0000036d),
    .LI(sig0000035c),
    .O(sig0000034c)
  );
  XORCY   blk00000224 (
    .CI(sig0000036e),
    .LI(sig0000035d),
    .O(sig0000034d)
  );
  XORCY   blk00000225 (
    .CI(sig0000036f),
    .LI(sig0000035e),
    .O(sig0000034e)
  );
  XORCY   blk00000226 (
    .CI(sig00000370),
    .LI(sig0000035f),
    .O(sig0000034f)
  );
  XORCY   blk00000227 (
    .CI(sig00000371),
    .LI(sig00000360),
    .O(sig00000350)
  );
  XORCY   blk00000228 (
    .CI(sig00000372),
    .LI(sig00000361),
    .O(sig00000351)
  );
  XORCY   blk00000229 (
    .CI(sig00000373),
    .LI(sig00000362),
    .O(sig00000352)
  );
  XORCY   blk0000022a (
    .CI(sig00000374),
    .LI(sig00000363),
    .O(sig00000353)
  );
  XORCY   blk0000022b (
    .CI(sig00000375),
    .LI(sig00000364),
    .O(sig00000354)
  );
  XORCY   blk0000022c (
    .CI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .LI(sig00000365),
    .O(sig00000355)
  );
  MUXCY   blk0000022d (
    .CI(sig00000367),
    .DI(sig000002bf),
    .S(sig00000c5e),
    .O(sig00000366)
  );
  MUXCY   blk0000022e (
    .CI(sig00000368),
    .DI(sig000002be),
    .S(sig00000357),
    .O(sig00000367)
  );
  MUXCY   blk0000022f (
    .CI(sig00000369),
    .DI(sig000002bd),
    .S(sig00000358),
    .O(sig00000368)
  );
  MUXCY   blk00000230 (
    .CI(sig0000036a),
    .DI(sig000002bc),
    .S(sig00000359),
    .O(sig00000369)
  );
  MUXCY   blk00000231 (
    .CI(sig0000036b),
    .DI(sig000002bb),
    .S(sig0000035a),
    .O(sig0000036a)
  );
  MUXCY   blk00000232 (
    .CI(sig0000036c),
    .DI(sig000002ba),
    .S(sig0000035b),
    .O(sig0000036b)
  );
  MUXCY   blk00000233 (
    .CI(sig0000036d),
    .DI(sig000002b9),
    .S(sig0000035c),
    .O(sig0000036c)
  );
  MUXCY   blk00000234 (
    .CI(sig0000036e),
    .DI(sig000002b8),
    .S(sig0000035d),
    .O(sig0000036d)
  );
  MUXCY   blk00000235 (
    .CI(sig0000036f),
    .DI(sig000002b7),
    .S(sig0000035e),
    .O(sig0000036e)
  );
  MUXCY   blk00000236 (
    .CI(sig00000370),
    .DI(sig000002b6),
    .S(sig0000035f),
    .O(sig0000036f)
  );
  MUXCY   blk00000237 (
    .CI(sig00000371),
    .DI(sig000002b5),
    .S(sig00000360),
    .O(sig00000370)
  );
  MUXCY   blk00000238 (
    .CI(sig00000372),
    .DI(sig000002b4),
    .S(sig00000361),
    .O(sig00000371)
  );
  MUXCY   blk00000239 (
    .CI(sig00000373),
    .DI(sig000002b3),
    .S(sig00000362),
    .O(sig00000372)
  );
  MUXCY   blk0000023a (
    .CI(sig00000374),
    .DI(sig000002b2),
    .S(sig00000363),
    .O(sig00000373)
  );
  MUXCY   blk0000023b (
    .CI(sig00000375),
    .DI(sig000002b1),
    .S(sig00000364),
    .O(sig00000374)
  );
  MUXCY   blk0000023c (
    .CI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .DI(sig000002b0),
    .S(sig00000365),
    .O(sig00000375)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000023d (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000345),
    .Q(sig000002af)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000023e (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000346),
    .Q(sig000002ae)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000023f (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000347),
    .Q(sig000002ad)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000240 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000348),
    .Q(sig000002ac)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000241 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000349),
    .Q(sig000002ab)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000242 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000034a),
    .Q(sig000002aa)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000243 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000034b),
    .Q(sig000002a9)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000244 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000034c),
    .Q(sig000002a8)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000245 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000034d),
    .Q(sig000002a7)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000246 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000034e),
    .Q(sig000002a6)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000247 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000034f),
    .Q(sig000002a5)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000248 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000350),
    .Q(sig000002a4)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000249 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000351),
    .Q(sig000002a3)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000024a (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000352),
    .Q(sig000002a2)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000024b (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000353),
    .Q(sig000002a1)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000024c (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000354),
    .Q(sig000002a0)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000024d (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000355),
    .Q(sig0000029f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000024e (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000313),
    .Q(sig0000029e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000024f (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000314),
    .Q(sig0000029d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000250 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000315),
    .Q(sig0000029c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000251 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000316),
    .Q(sig0000029b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000252 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000317),
    .Q(sig0000029a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000253 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000318),
    .Q(sig00000299)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000254 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000319),
    .Q(sig00000298)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000255 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000031a),
    .Q(sig00000297)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000256 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000031b),
    .Q(sig00000296)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000257 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000031c),
    .Q(sig00000295)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000258 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000031d),
    .Q(sig00000294)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000259 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000031e),
    .Q(sig00000293)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000025a (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000031f),
    .Q(sig00000292)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000025b (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000320),
    .Q(sig00000291)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000025c (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000321),
    .Q(sig00000290)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000025d (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000322),
    .Q(sig0000028f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000025e (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000323),
    .Q(sig0000028e)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000025f (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(sig00000344),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig0000027c),
    .Q(sig00000376)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000260 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(sig00000344),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig0000027b),
    .Q(sig00000377)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000261 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(sig00000344),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig0000027a),
    .Q(sig00000378)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000262 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(sig00000344),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000279),
    .Q(sig00000379)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000263 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(sig00000344),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000278),
    .Q(sig0000037a)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000264 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(sig00000344),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000277),
    .Q(sig0000037b)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000265 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(sig00000344),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000276),
    .Q(sig0000037c)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000266 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(sig00000344),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000275),
    .Q(sig0000037d)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000267 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(sig00000344),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000274),
    .Q(sig0000037e)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000268 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(sig00000344),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000273),
    .Q(sig0000037f)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000269 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(sig00000344),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000272),
    .Q(sig00000380)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000026a (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(sig00000344),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000271),
    .Q(sig00000381)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000026b (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(sig00000344),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000270),
    .Q(sig00000382)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000026c (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(sig00000344),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig0000026f),
    .Q(sig00000383)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000026d (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(sig00000344),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig0000026e),
    .Q(sig00000384)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000026e (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(sig00000344),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig0000026d),
    .Q(sig00000385)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000026f (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(sig00000344),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig0000026c),
    .Q(sig00000386)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000270 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000376),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000203)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000271 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000377),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000202)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000272 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000378),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000201)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000273 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000379),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000200)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000274 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000037a),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000001ff)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000275 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000037b),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000001fe)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000276 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000037c),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000001fd)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000277 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000037d),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000001fc)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000278 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000037e),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000001fb)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000279 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000037f),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000001fa)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000027a (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000380),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000001f9)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000027b (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000381),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000001f8)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000027c (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000382),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000001f7)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000027d (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000383),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000001f6)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000027e (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000384),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000001f5)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000027f (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000385),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000001f4)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000280 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000386),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000001f3)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000281 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(sig00000344),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig0000029e),
    .Q(sig00000387)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000282 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(sig00000344),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig0000029d),
    .Q(sig00000388)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000283 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(sig00000344),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig0000029c),
    .Q(sig00000389)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000284 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(sig00000344),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig0000029b),
    .Q(sig0000038a)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000285 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(sig00000344),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig0000029a),
    .Q(sig0000038b)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000286 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(sig00000344),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000299),
    .Q(sig0000038c)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000287 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(sig00000344),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000298),
    .Q(sig0000038d)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000288 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(sig00000344),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000297),
    .Q(sig0000038e)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000289 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(sig00000344),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000296),
    .Q(sig0000038f)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000028a (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(sig00000344),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000295),
    .Q(sig00000390)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000028b (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(sig00000344),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000294),
    .Q(sig00000391)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000028c (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(sig00000344),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000293),
    .Q(sig00000392)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000028d (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(sig00000344),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000292),
    .Q(sig00000393)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000028e (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(sig00000344),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000291),
    .Q(sig00000394)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000028f (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(sig00000344),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000290),
    .Q(sig00000395)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000290 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(sig00000344),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig0000028f),
    .Q(sig00000396)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000291 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(sig00000344),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig0000028e),
    .Q(sig00000397)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000292 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000387),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig0000028d)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000293 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000388),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig0000028c)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000294 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000389),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig0000028b)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000295 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000038a),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig0000028a)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000296 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000038b),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000289)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000297 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000038c),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000288)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000298 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000038d),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000287)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000299 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000038e),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000286)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000029a (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000038f),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000285)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000029b (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000390),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000284)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000029c (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000391),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000283)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000029d (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000392),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000282)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000029e (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000393),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000281)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000029f (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000394),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000280)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000002a0 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000395),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig0000027f)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000002a1 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000396),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig0000027e)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000002a2 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000397),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig0000027d)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000002c7 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(sig00000344),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000208),
    .Q(sig00000398)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000002c8 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(sig00000344),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000207),
    .Q(sig00000399)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000002c9 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(sig00000344),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000206),
    .Q(sig0000039a)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000002ca (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(sig00000344),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000205),
    .Q(sig0000039b)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000002cb (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000398),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(NLW_blk000002cb_Q_UNCONNECTED)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000002cc (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000399),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(NLW_blk000002cc_Q_UNCONNECTED)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000002cd (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000039a),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(NLW_blk000002cd_Q_UNCONNECTED)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000002ce (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000039b),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(NLW_blk000002ce_Q_UNCONNECTED)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000002cf (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(sig00000344),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig0000020d),
    .Q(sig0000039c)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000002d0 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(sig00000344),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig0000020c),
    .Q(sig0000039d)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000002d1 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(sig00000344),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig0000020b),
    .Q(sig0000039e)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000002d2 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(sig00000344),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig0000020a),
    .Q(sig0000039f)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000002d3 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000039c),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000001d9)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000002d4 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000039d),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000001d8)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000002d5 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000039e),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(NLW_blk000002d5_Q_UNCONNECTED)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000002d6 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000039f),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(NLW_blk000002d6_Q_UNCONNECTED)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000002d7 (
    .I0(sig00000455),
    .I1(sig000004e5),
    .I2(sig00000530),
    .O(sig000003a0)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000002d8 (
    .I0(sig00000456),
    .I1(sig000004e6),
    .I2(sig00000530),
    .O(sig000003a1)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000002d9 (
    .I0(sig00000457),
    .I1(sig000004e7),
    .I2(sig00000530),
    .O(sig000003a2)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000002da (
    .I0(sig00000458),
    .I1(sig000004e8),
    .I2(sig00000530),
    .O(sig000003a3)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000002db (
    .I0(sig00000459),
    .I1(sig000004e9),
    .I2(sig00000530),
    .O(sig000003a4)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000002dc (
    .I0(sig0000045a),
    .I1(sig000004ea),
    .I2(sig00000530),
    .O(sig000003a5)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000002dd (
    .I0(sig0000045b),
    .I1(sig000004eb),
    .I2(sig00000530),
    .O(sig000003a6)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000002de (
    .I0(sig0000045c),
    .I1(sig000004ec),
    .I2(sig00000530),
    .O(sig000003a7)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000002df (
    .I0(sig0000045d),
    .I1(sig000004ed),
    .I2(sig00000530),
    .O(sig000003a8)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000002e0 (
    .I0(sig0000045e),
    .I1(sig000004ee),
    .I2(sig00000530),
    .O(sig000003a9)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000002e1 (
    .I0(sig0000045f),
    .I1(sig000004ef),
    .I2(sig00000530),
    .O(sig000003aa)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000002e2 (
    .I0(sig00000460),
    .I1(sig000004f0),
    .I2(sig00000530),
    .O(sig000003ab)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000002e3 (
    .I0(sig00000461),
    .I1(sig000004f1),
    .I2(sig00000530),
    .O(sig000003ac)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000002e4 (
    .I0(sig00000462),
    .I1(sig000004f2),
    .I2(sig00000530),
    .O(sig000003ad)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000002e5 (
    .I0(sig00000463),
    .I1(sig000004f3),
    .I2(sig00000530),
    .O(sig000003ae)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000002e6 (
    .I0(sig00000464),
    .I1(sig000004f4),
    .I2(sig00000530),
    .O(sig000003af)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000002e7 (
    .I0(sig00000465),
    .I1(sig000004f5),
    .I2(sig00000530),
    .O(sig000003b0)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000002e8 (
    .I0(sig00000466),
    .I1(sig000004f6),
    .I2(sig00000530),
    .O(sig000003b1)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000002e9 (
    .I0(sig000004e5),
    .I1(sig00000455),
    .I2(sig00000530),
    .O(sig000003b2)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000002ea (
    .I0(sig000004e6),
    .I1(sig00000456),
    .I2(sig00000530),
    .O(sig000003b3)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000002eb (
    .I0(sig000004e7),
    .I1(sig00000457),
    .I2(sig00000530),
    .O(sig000003b4)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000002ec (
    .I0(sig000004e8),
    .I1(sig00000458),
    .I2(sig00000530),
    .O(sig000003b5)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000002ed (
    .I0(sig000004e9),
    .I1(sig00000459),
    .I2(sig00000530),
    .O(sig000003b6)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000002ee (
    .I0(sig000004ea),
    .I1(sig0000045a),
    .I2(sig00000530),
    .O(sig000003b7)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000002ef (
    .I0(sig000004eb),
    .I1(sig0000045b),
    .I2(sig00000530),
    .O(sig000003b8)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000002f0 (
    .I0(sig000004ec),
    .I1(sig0000045c),
    .I2(sig00000530),
    .O(sig000003b9)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000002f1 (
    .I0(sig000004ed),
    .I1(sig0000045d),
    .I2(sig00000530),
    .O(sig000003ba)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000002f2 (
    .I0(sig000004ee),
    .I1(sig0000045e),
    .I2(sig00000530),
    .O(sig000003bb)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000002f3 (
    .I0(sig000004ef),
    .I1(sig0000045f),
    .I2(sig00000530),
    .O(sig000003bc)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000002f4 (
    .I0(sig000004f0),
    .I1(sig00000460),
    .I2(sig00000530),
    .O(sig000003bd)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000002f5 (
    .I0(sig000004f1),
    .I1(sig00000461),
    .I2(sig00000530),
    .O(sig000003be)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000002f6 (
    .I0(sig000004f2),
    .I1(sig00000462),
    .I2(sig00000530),
    .O(sig000003bf)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000002f7 (
    .I0(sig000004f3),
    .I1(sig00000463),
    .I2(sig00000530),
    .O(sig000003c0)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000002f8 (
    .I0(sig000004f4),
    .I1(sig00000464),
    .I2(sig00000530),
    .O(sig000003c1)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000002f9 (
    .I0(sig000004f5),
    .I1(sig00000465),
    .I2(sig00000530),
    .O(sig000003c2)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000002fa (
    .I0(sig000004f6),
    .I1(sig00000466),
    .I2(sig00000530),
    .O(sig000003c3)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000002fb (
    .I0(sig000004af),
    .I1(sig0000048b),
    .I2(sig0000052e),
    .O(sig000003c4)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000002fc (
    .I0(sig000004b0),
    .I1(sig0000048c),
    .I2(sig0000052e),
    .O(sig000003c5)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000002fd (
    .I0(sig000004b1),
    .I1(sig0000048d),
    .I2(sig0000052e),
    .O(sig000003c6)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000002fe (
    .I0(sig000004b2),
    .I1(sig0000048e),
    .I2(sig0000052e),
    .O(sig000003c7)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000002ff (
    .I0(sig000004b3),
    .I1(sig0000048f),
    .I2(sig0000052e),
    .O(sig000003c8)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000300 (
    .I0(sig000004b4),
    .I1(sig00000490),
    .I2(sig0000052e),
    .O(sig000003c9)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000301 (
    .I0(sig000004b5),
    .I1(sig00000491),
    .I2(sig0000052e),
    .O(sig000003ca)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000302 (
    .I0(sig000004b6),
    .I1(sig00000492),
    .I2(sig0000052e),
    .O(sig000003cb)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000303 (
    .I0(sig000004b7),
    .I1(sig00000493),
    .I2(sig0000052e),
    .O(sig000003cc)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000304 (
    .I0(sig000004b8),
    .I1(sig00000494),
    .I2(sig0000052e),
    .O(sig000003cd)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000305 (
    .I0(sig000004b9),
    .I1(sig00000495),
    .I2(sig0000052e),
    .O(sig000003ce)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000306 (
    .I0(sig000004ba),
    .I1(sig00000496),
    .I2(sig0000052e),
    .O(sig000003cf)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000307 (
    .I0(sig000004bb),
    .I1(sig00000497),
    .I2(sig0000052e),
    .O(sig000003d0)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000308 (
    .I0(sig000004bc),
    .I1(sig00000498),
    .I2(sig0000052e),
    .O(sig000003d1)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000309 (
    .I0(sig000004bd),
    .I1(sig00000499),
    .I2(sig0000052e),
    .O(sig000003d2)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk0000030a (
    .I0(sig000004be),
    .I1(sig0000049a),
    .I2(sig0000052e),
    .O(sig000003d3)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk0000030b (
    .I0(sig000004bf),
    .I1(sig0000049b),
    .I2(sig0000052e),
    .O(sig000003d4)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk0000030c (
    .I0(sig000004c0),
    .I1(sig0000049c),
    .I2(sig0000052e),
    .O(sig000003d5)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk0000030d (
    .I0(sig0000048b),
    .I1(sig000004af),
    .I2(sig0000052e),
    .O(sig000003d6)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk0000030e (
    .I0(sig0000048c),
    .I1(sig000004b0),
    .I2(sig0000052e),
    .O(sig000003d7)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk0000030f (
    .I0(sig0000048d),
    .I1(sig000004b1),
    .I2(sig0000052e),
    .O(sig000003d8)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000310 (
    .I0(sig0000048e),
    .I1(sig000004b2),
    .I2(sig0000052e),
    .O(sig000003d9)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000311 (
    .I0(sig0000048f),
    .I1(sig000004b3),
    .I2(sig0000052e),
    .O(sig000003da)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000312 (
    .I0(sig00000490),
    .I1(sig000004b4),
    .I2(sig0000052e),
    .O(sig000003db)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000313 (
    .I0(sig00000491),
    .I1(sig000004b5),
    .I2(sig0000052e),
    .O(sig000003dc)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000314 (
    .I0(sig00000492),
    .I1(sig000004b6),
    .I2(sig0000052e),
    .O(sig000003dd)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000315 (
    .I0(sig00000493),
    .I1(sig000004b7),
    .I2(sig0000052e),
    .O(sig000003de)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000316 (
    .I0(sig00000494),
    .I1(sig000004b8),
    .I2(sig0000052e),
    .O(sig000003df)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000317 (
    .I0(sig00000495),
    .I1(sig000004b9),
    .I2(sig0000052e),
    .O(sig000003e0)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000318 (
    .I0(sig00000496),
    .I1(sig000004ba),
    .I2(sig0000052e),
    .O(sig000003e1)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000319 (
    .I0(sig00000497),
    .I1(sig000004bb),
    .I2(sig0000052e),
    .O(sig000003e2)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk0000031a (
    .I0(sig00000498),
    .I1(sig000004bc),
    .I2(sig0000052e),
    .O(sig000003e3)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk0000031b (
    .I0(sig00000499),
    .I1(sig000004bd),
    .I2(sig0000052e),
    .O(sig000003e4)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk0000031c (
    .I0(sig0000049a),
    .I1(sig000004be),
    .I2(sig0000052e),
    .O(sig000003e5)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk0000031d (
    .I0(sig0000049b),
    .I1(sig000004bf),
    .I2(sig0000052e),
    .O(sig000003e6)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk0000031e (
    .I0(sig0000049c),
    .I1(sig000004c0),
    .I2(sig0000052e),
    .O(sig000003e7)
  );
  MUXCY   blk0000031f (
    .CI(sig0000041d),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig000003e8),
    .O(sig000003fa)
  );
  XORCY   blk00000320 (
    .CI(sig0000041d),
    .LI(sig000003e8),
    .O(sig000003fb)
  );
  MUXCY   blk00000321 (
    .CI(sig000003fa),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig000003e9),
    .O(sig000003fc)
  );
  XORCY   blk00000322 (
    .CI(sig000003fa),
    .LI(sig000003e9),
    .O(sig000003fd)
  );
  MUXCY   blk00000323 (
    .CI(sig000003fc),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig000003ea),
    .O(sig000003fe)
  );
  XORCY   blk00000324 (
    .CI(sig000003fc),
    .LI(sig000003ea),
    .O(sig000003ff)
  );
  MUXCY   blk00000325 (
    .CI(sig000003fe),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig000003eb),
    .O(sig00000400)
  );
  XORCY   blk00000326 (
    .CI(sig000003fe),
    .LI(sig000003eb),
    .O(sig00000401)
  );
  MUXCY   blk00000327 (
    .CI(sig00000400),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig000003ec),
    .O(sig00000402)
  );
  XORCY   blk00000328 (
    .CI(sig00000400),
    .LI(sig000003ec),
    .O(sig00000403)
  );
  MUXCY   blk00000329 (
    .CI(sig00000402),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig000003ed),
    .O(sig00000404)
  );
  XORCY   blk0000032a (
    .CI(sig00000402),
    .LI(sig000003ed),
    .O(sig00000405)
  );
  MUXCY   blk0000032b (
    .CI(sig00000404),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig000003ee),
    .O(sig00000406)
  );
  XORCY   blk0000032c (
    .CI(sig00000404),
    .LI(sig000003ee),
    .O(sig00000407)
  );
  MUXCY   blk0000032d (
    .CI(sig00000406),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig000003ef),
    .O(sig00000408)
  );
  XORCY   blk0000032e (
    .CI(sig00000406),
    .LI(sig000003ef),
    .O(sig00000409)
  );
  MUXCY   blk0000032f (
    .CI(sig00000408),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig000003f0),
    .O(sig0000040a)
  );
  XORCY   blk00000330 (
    .CI(sig00000408),
    .LI(sig000003f0),
    .O(sig0000040b)
  );
  MUXCY   blk00000331 (
    .CI(sig0000040a),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig000003f1),
    .O(sig0000040c)
  );
  XORCY   blk00000332 (
    .CI(sig0000040a),
    .LI(sig000003f1),
    .O(sig0000040d)
  );
  MUXCY   blk00000333 (
    .CI(sig0000040c),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig000003f2),
    .O(sig0000040e)
  );
  XORCY   blk00000334 (
    .CI(sig0000040c),
    .LI(sig000003f2),
    .O(sig0000040f)
  );
  MUXCY   blk00000335 (
    .CI(sig0000040e),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig000003f3),
    .O(sig00000410)
  );
  XORCY   blk00000336 (
    .CI(sig0000040e),
    .LI(sig000003f3),
    .O(sig00000411)
  );
  MUXCY   blk00000337 (
    .CI(sig00000410),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig000003f4),
    .O(sig00000412)
  );
  XORCY   blk00000338 (
    .CI(sig00000410),
    .LI(sig000003f4),
    .O(sig00000413)
  );
  MUXCY   blk00000339 (
    .CI(sig00000412),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig000003f5),
    .O(sig00000414)
  );
  XORCY   blk0000033a (
    .CI(sig00000412),
    .LI(sig000003f5),
    .O(sig00000415)
  );
  MUXCY   blk0000033b (
    .CI(sig00000414),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig000003f6),
    .O(sig00000416)
  );
  XORCY   blk0000033c (
    .CI(sig00000414),
    .LI(sig000003f6),
    .O(sig00000417)
  );
  MUXCY   blk0000033d (
    .CI(sig00000416),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig000003f7),
    .O(sig00000418)
  );
  XORCY   blk0000033e (
    .CI(sig00000416),
    .LI(sig000003f7),
    .O(sig00000419)
  );
  MUXCY   blk0000033f (
    .CI(sig00000418),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig00000c5f),
    .O(sig0000041a)
  );
  XORCY   blk00000340 (
    .CI(sig00000418),
    .LI(sig00000c5f),
    .O(sig0000041b)
  );
  MUXCY   blk00000341 (
    .CI(sig0000041a),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig000003f8),
    .O(NLW_blk00000341_O_UNCONNECTED)
  );
  XORCY   blk00000342 (
    .CI(sig0000041a),
    .LI(sig000003f8),
    .O(sig0000041c)
  );
  MUXCY   blk00000343 (
    .CI(sig00000344),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig000003f9),
    .O(sig0000041d)
  );
  MUXCY   blk00000344 (
    .CI(sig00000453),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig0000041e),
    .O(sig00000430)
  );
  XORCY   blk00000345 (
    .CI(sig00000453),
    .LI(sig0000041e),
    .O(sig00000431)
  );
  MUXCY   blk00000346 (
    .CI(sig00000430),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig0000041f),
    .O(sig00000432)
  );
  XORCY   blk00000347 (
    .CI(sig00000430),
    .LI(sig0000041f),
    .O(sig00000433)
  );
  MUXCY   blk00000348 (
    .CI(sig00000432),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig00000420),
    .O(sig00000434)
  );
  XORCY   blk00000349 (
    .CI(sig00000432),
    .LI(sig00000420),
    .O(sig00000435)
  );
  MUXCY   blk0000034a (
    .CI(sig00000434),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig00000421),
    .O(sig00000436)
  );
  XORCY   blk0000034b (
    .CI(sig00000434),
    .LI(sig00000421),
    .O(sig00000437)
  );
  MUXCY   blk0000034c (
    .CI(sig00000436),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig00000422),
    .O(sig00000438)
  );
  XORCY   blk0000034d (
    .CI(sig00000436),
    .LI(sig00000422),
    .O(sig00000439)
  );
  MUXCY   blk0000034e (
    .CI(sig00000438),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig00000423),
    .O(sig0000043a)
  );
  XORCY   blk0000034f (
    .CI(sig00000438),
    .LI(sig00000423),
    .O(sig0000043b)
  );
  MUXCY   blk00000350 (
    .CI(sig0000043a),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig00000424),
    .O(sig0000043c)
  );
  XORCY   blk00000351 (
    .CI(sig0000043a),
    .LI(sig00000424),
    .O(sig0000043d)
  );
  MUXCY   blk00000352 (
    .CI(sig0000043c),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig00000425),
    .O(sig0000043e)
  );
  XORCY   blk00000353 (
    .CI(sig0000043c),
    .LI(sig00000425),
    .O(sig0000043f)
  );
  MUXCY   blk00000354 (
    .CI(sig0000043e),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig00000426),
    .O(sig00000440)
  );
  XORCY   blk00000355 (
    .CI(sig0000043e),
    .LI(sig00000426),
    .O(sig00000441)
  );
  MUXCY   blk00000356 (
    .CI(sig00000440),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig00000427),
    .O(sig00000442)
  );
  XORCY   blk00000357 (
    .CI(sig00000440),
    .LI(sig00000427),
    .O(sig00000443)
  );
  MUXCY   blk00000358 (
    .CI(sig00000442),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig00000428),
    .O(sig00000444)
  );
  XORCY   blk00000359 (
    .CI(sig00000442),
    .LI(sig00000428),
    .O(sig00000445)
  );
  MUXCY   blk0000035a (
    .CI(sig00000444),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig00000429),
    .O(sig00000446)
  );
  XORCY   blk0000035b (
    .CI(sig00000444),
    .LI(sig00000429),
    .O(sig00000447)
  );
  MUXCY   blk0000035c (
    .CI(sig00000446),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig0000042a),
    .O(sig00000448)
  );
  XORCY   blk0000035d (
    .CI(sig00000446),
    .LI(sig0000042a),
    .O(sig00000449)
  );
  MUXCY   blk0000035e (
    .CI(sig00000448),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig0000042b),
    .O(sig0000044a)
  );
  XORCY   blk0000035f (
    .CI(sig00000448),
    .LI(sig0000042b),
    .O(sig0000044b)
  );
  MUXCY   blk00000360 (
    .CI(sig0000044a),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig0000042c),
    .O(sig0000044c)
  );
  XORCY   blk00000361 (
    .CI(sig0000044a),
    .LI(sig0000042c),
    .O(sig0000044d)
  );
  MUXCY   blk00000362 (
    .CI(sig0000044c),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig0000042d),
    .O(sig0000044e)
  );
  XORCY   blk00000363 (
    .CI(sig0000044c),
    .LI(sig0000042d),
    .O(sig0000044f)
  );
  MUXCY   blk00000364 (
    .CI(sig0000044e),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig00000c60),
    .O(sig00000450)
  );
  XORCY   blk00000365 (
    .CI(sig0000044e),
    .LI(sig00000c60),
    .O(sig00000451)
  );
  MUXCY   blk00000366 (
    .CI(sig00000450),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig0000042e),
    .O(NLW_blk00000366_O_UNCONNECTED)
  );
  XORCY   blk00000367 (
    .CI(sig00000450),
    .LI(sig0000042e),
    .O(sig00000452)
  );
  MUXCY   blk00000368 (
    .CI(sig00000344),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig0000042f),
    .O(sig00000453)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000369 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000003a0),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000004d3)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000036a (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000003a1),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000004d4)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000036b (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000003a2),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000004d5)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000036c (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000003a3),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000004d6)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000036d (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000003a4),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000004d7)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000036e (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000003a5),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000004d8)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000036f (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000003a6),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000004d9)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000370 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000003a7),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000004da)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000371 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000003a8),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000004db)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000372 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000003a9),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000004dc)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000373 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000003aa),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000004dd)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000374 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000003ab),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000004de)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000375 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000003ac),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000004df)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000376 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000003ad),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000004e0)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000377 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000003ae),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000004e1)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000378 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000003af),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000004e2)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000379 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000003b0),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000004e3)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000037a (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000003b1),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000004e4)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000037b (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000003b2),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000004c1)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000037c (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000003b3),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000004c2)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000037d (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000003b4),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000004c3)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000037e (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000003b5),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000004c4)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000037f (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000003b6),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000004c5)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000380 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000003b7),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000004c6)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000381 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000003b8),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000004c7)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000382 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000003b9),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000004c8)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000383 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000003ba),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000004c9)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000384 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000003bb),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000004ca)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000385 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000003bc),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000004cb)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000386 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000003bd),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000004cc)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000387 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000003be),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000004cd)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000388 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000003bf),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000004ce)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000389 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000003c0),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000004cf)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000038a (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000003c1),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000004d0)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000038b (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000003c2),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000004d1)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000038c (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000003c3),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000004d2)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000038d (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000003c4),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000479)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000038e (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000003c5),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig0000047a)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000038f (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000003c6),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig0000047b)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000390 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000003c7),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig0000047c)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000391 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000003c8),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig0000047d)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000392 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000003c9),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig0000047e)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000393 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000003ca),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig0000047f)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000394 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000003cb),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000480)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000395 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000003cc),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000481)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000396 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000003cd),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000482)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000397 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000003ce),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000483)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000398 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000003cf),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000484)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000399 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000003d0),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000485)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000039a (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000003d1),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000486)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000039b (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000003d2),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000487)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000039c (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000003d3),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000488)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000039d (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000003d4),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000489)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000039e (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000003d5),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig0000048a)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000039f (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000003d6),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000001b4)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000003a0 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000003d7),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000001b5)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000003a1 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000003d8),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000001b6)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000003a2 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000003d9),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000001b7)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000003a3 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000003da),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000001b8)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000003a4 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000003db),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000001b9)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000003a5 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000003dc),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000001ba)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000003a6 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000003dd),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000001bb)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000003a7 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000003de),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000001bc)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000003a8 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000003df),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000001bd)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000003a9 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000003e0),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000001be)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000003aa (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000003e1),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000001bf)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000003ab (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000003e2),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000001c0)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000003ac (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000003e3),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000001c1)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000003ad (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000003e4),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000001c2)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000003ae (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000003e5),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000001c3)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000003af (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000003e6),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000001c4)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000003b0 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000003e7),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000001c5)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003b1 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000003fb),
    .Q(sig00000509)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003b2 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000003fd),
    .Q(sig0000050a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003b3 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000003ff),
    .Q(sig0000050b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003b4 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000401),
    .Q(sig0000050c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003b5 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000403),
    .Q(sig0000050d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003b6 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000405),
    .Q(sig0000050e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003b7 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000407),
    .Q(sig0000050f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003b8 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000409),
    .Q(sig00000510)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003b9 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000040b),
    .Q(sig00000511)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003ba (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000040d),
    .Q(sig00000512)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003bb (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000040f),
    .Q(sig00000513)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003bc (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000411),
    .Q(sig00000514)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003bd (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000413),
    .Q(sig00000515)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003be (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000415),
    .Q(sig00000516)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003bf (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000417),
    .Q(sig00000517)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003c0 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000419),
    .Q(sig00000518)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003c1 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000041b),
    .Q(sig00000519)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003c2 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000041c),
    .Q(sig0000051a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003c3 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000431),
    .Q(sig0000051b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003c4 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000433),
    .Q(sig0000051c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003c5 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000435),
    .Q(sig0000051d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003c6 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000437),
    .Q(sig0000051e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003c7 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000439),
    .Q(sig0000051f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003c8 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000043b),
    .Q(sig00000520)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003c9 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000043d),
    .Q(sig00000521)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003ca (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000043f),
    .Q(sig00000522)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003cb (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000441),
    .Q(sig00000523)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003cc (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000443),
    .Q(sig00000524)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003cd (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000445),
    .Q(sig00000525)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003ce (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000447),
    .Q(sig00000526)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003cf (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000449),
    .Q(sig00000527)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003d0 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000044b),
    .Q(sig00000528)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003d1 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000044d),
    .Q(sig00000529)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003d2 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000044f),
    .Q(sig0000052a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003d3 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000451),
    .Q(sig0000052b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003d4 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000452),
    .Q(sig0000052c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003d5 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000001e0),
    .Q(sig00000532)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003d6 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000454),
    .Q(sig0000052d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003d7 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000001d8),
    .Q(sig00000531)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000003d8 (
    .C(aclk),
    .D(sig0000052c),
    .Q(sig00000466)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000003d9 (
    .C(aclk),
    .D(sig0000052b),
    .Q(sig00000465)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000003da (
    .C(aclk),
    .D(sig0000052a),
    .Q(sig00000464)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000003db (
    .C(aclk),
    .D(sig00000529),
    .Q(sig00000463)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000003dc (
    .C(aclk),
    .D(sig00000528),
    .Q(sig00000462)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000003dd (
    .C(aclk),
    .D(sig00000527),
    .Q(sig00000461)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000003de (
    .C(aclk),
    .D(sig00000526),
    .Q(sig00000460)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000003df (
    .C(aclk),
    .D(sig00000525),
    .Q(sig0000045f)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000003e0 (
    .C(aclk),
    .D(sig00000524),
    .Q(sig0000045e)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000003e1 (
    .C(aclk),
    .D(sig00000523),
    .Q(sig0000045d)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000003e2 (
    .C(aclk),
    .D(sig00000522),
    .Q(sig0000045c)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000003e3 (
    .C(aclk),
    .D(sig00000521),
    .Q(sig0000045b)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000003e4 (
    .C(aclk),
    .D(sig00000520),
    .Q(sig0000045a)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000003e5 (
    .C(aclk),
    .D(sig0000051f),
    .Q(sig00000459)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000003e6 (
    .C(aclk),
    .D(sig0000051e),
    .Q(sig00000458)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000003e7 (
    .C(aclk),
    .D(sig0000051d),
    .Q(sig00000457)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000003e8 (
    .C(aclk),
    .D(sig0000051c),
    .Q(sig00000456)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000003e9 (
    .C(aclk),
    .D(sig0000051b),
    .Q(sig00000455)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000003ea (
    .C(aclk),
    .D(sig0000051a),
    .Q(sig00000478)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000003eb (
    .C(aclk),
    .D(sig00000519),
    .Q(sig00000477)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000003ec (
    .C(aclk),
    .D(sig00000518),
    .Q(sig00000476)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000003ed (
    .C(aclk),
    .D(sig00000517),
    .Q(sig00000475)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000003ee (
    .C(aclk),
    .D(sig00000516),
    .Q(sig00000474)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000003ef (
    .C(aclk),
    .D(sig00000515),
    .Q(sig00000473)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000003f0 (
    .C(aclk),
    .D(sig00000514),
    .Q(sig00000472)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000003f1 (
    .C(aclk),
    .D(sig00000513),
    .Q(sig00000471)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000003f2 (
    .C(aclk),
    .D(sig00000512),
    .Q(sig00000470)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000003f3 (
    .C(aclk),
    .D(sig00000511),
    .Q(sig0000046f)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000003f4 (
    .C(aclk),
    .D(sig00000510),
    .Q(sig0000046e)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000003f5 (
    .C(aclk),
    .D(sig0000050f),
    .Q(sig0000046d)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000003f6 (
    .C(aclk),
    .D(sig0000050e),
    .Q(sig0000046c)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000003f7 (
    .C(aclk),
    .D(sig0000050d),
    .Q(sig0000046b)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000003f8 (
    .C(aclk),
    .D(sig0000050c),
    .Q(sig0000046a)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000003f9 (
    .C(aclk),
    .D(sig0000050b),
    .Q(sig00000469)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000003fa (
    .C(aclk),
    .D(sig0000050a),
    .Q(sig00000468)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000003fb (
    .C(aclk),
    .D(sig00000509),
    .Q(sig00000467)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000409 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig0000048a),
    .Q(sig00000533)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000040a (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000489),
    .Q(sig00000534)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000040b (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000488),
    .Q(sig00000535)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000040c (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000487),
    .Q(sig00000536)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000040d (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000486),
    .Q(sig00000537)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000040e (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000485),
    .Q(sig00000538)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000040f (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000484),
    .Q(sig00000539)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000410 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000483),
    .Q(sig0000053a)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000411 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000482),
    .Q(sig0000053b)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000412 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000481),
    .Q(sig0000053c)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000413 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000480),
    .Q(sig0000053d)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000414 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig0000047f),
    .Q(sig0000053e)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000415 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig0000047e),
    .Q(sig0000053f)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000416 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig0000047d),
    .Q(sig00000540)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000417 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig0000047c),
    .Q(sig00000541)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000418 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig0000047b),
    .Q(sig00000542)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000419 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig0000047a),
    .Q(sig00000543)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000041a (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000479),
    .Q(sig00000544)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000041b (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000533),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000001d7)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000041c (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000534),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000001d6)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000041d (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000535),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000001d5)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000041e (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000536),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000001d4)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000041f (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000537),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000001d3)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000420 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000538),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000001d2)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000421 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000539),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000001d1)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000422 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000053a),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000001d0)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000423 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000053b),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000001cf)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000424 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000053c),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000001ce)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000425 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000053d),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000001cd)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000426 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000053e),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000001cc)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000427 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000053f),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000001cb)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000428 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000540),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000001ca)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000429 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000541),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000001c9)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000042a (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000542),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000001c8)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000042b (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000543),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000001c7)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000042c (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000544),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000001c6)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000042d (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000004ae),
    .Q(sig00000545)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000042e (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000004ad),
    .Q(sig00000546)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000042f (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000004ac),
    .Q(sig00000547)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000430 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000004ab),
    .Q(sig00000548)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000431 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000004aa),
    .Q(sig00000549)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000432 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000004a9),
    .Q(sig0000054a)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000433 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000004a8),
    .Q(sig0000054b)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000434 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000004a7),
    .Q(sig0000054c)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000435 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000004a6),
    .Q(sig0000054d)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000436 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000004a5),
    .Q(sig0000054e)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000437 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000004a4),
    .Q(sig0000054f)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000438 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000004a3),
    .Q(sig00000550)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000439 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000004a2),
    .Q(sig00000551)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000043a (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000004a1),
    .Q(sig00000552)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000043b (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000004a0),
    .Q(sig00000553)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000043c (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig0000049f),
    .Q(sig00000554)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000043d (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig0000049e),
    .Q(sig00000555)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000043e (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig0000049d),
    .Q(sig00000556)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000043f (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000545),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig0000049c)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000440 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000546),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig0000049b)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000441 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000547),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig0000049a)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000442 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000548),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000499)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000443 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000549),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000498)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000444 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000054a),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000497)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000445 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000054b),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000496)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000446 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000054c),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000495)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000447 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000054d),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000494)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000448 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000054e),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000493)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000449 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000054f),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000492)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000044a (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000550),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000491)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000044b (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000551),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000490)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000044c (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000552),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig0000048f)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000044d (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000553),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig0000048e)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000044e (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000554),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig0000048d)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000044f (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000555),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig0000048c)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000450 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000556),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig0000048b)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000451 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000478),
    .Q(sig00000557)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000452 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000477),
    .Q(sig00000558)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000453 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000476),
    .Q(sig00000559)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000454 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000475),
    .Q(sig0000055a)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000455 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000474),
    .Q(sig0000055b)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000456 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000473),
    .Q(sig0000055c)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000457 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000472),
    .Q(sig0000055d)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000458 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000471),
    .Q(sig0000055e)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000459 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000470),
    .Q(sig0000055f)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000045a (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig0000046f),
    .Q(sig00000560)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000045b (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig0000046e),
    .Q(sig00000561)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000045c (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig0000046d),
    .Q(sig00000562)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000045d (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig0000046c),
    .Q(sig00000563)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000045e (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig0000046b),
    .Q(sig00000564)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000045f (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig0000046a),
    .Q(sig00000565)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000460 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000469),
    .Q(sig00000566)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000461 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000468),
    .Q(sig00000567)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000462 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000467),
    .Q(sig00000568)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000463 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000557),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000004f6)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000464 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000558),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000004f5)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000465 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000559),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000004f4)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000466 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000055a),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000004f3)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000467 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000055b),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000004f2)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000468 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000055c),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000004f1)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000469 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000055d),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000004f0)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000046a (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000055e),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000004ef)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000046b (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000055f),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000004ee)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000046c (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000560),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000004ed)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000046d (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000561),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000004ec)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000046e (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000562),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000004eb)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000046f (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000563),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000004ea)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000470 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000564),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000004e9)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000471 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000565),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000004e8)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000472 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000566),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000004e7)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000473 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000567),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000004e6)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000474 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000568),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000004e5)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000475 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000004e4),
    .Q(sig00000569)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000476 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000004e3),
    .Q(sig0000056a)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000477 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000004e2),
    .Q(sig0000056b)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000478 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000004e1),
    .Q(sig0000056c)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000479 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000004e0),
    .Q(sig0000056d)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000047a (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000004df),
    .Q(sig0000056e)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000047b (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000004de),
    .Q(sig0000056f)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000047c (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000004dd),
    .Q(sig00000570)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000047d (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000004dc),
    .Q(sig00000571)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000047e (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000004db),
    .Q(sig00000572)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000047f (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000004da),
    .Q(sig00000573)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000480 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000004d9),
    .Q(sig00000574)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000481 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000004d8),
    .Q(sig00000575)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000482 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000004d7),
    .Q(sig00000576)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000483 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000004d6),
    .Q(sig00000577)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000484 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000004d5),
    .Q(sig00000578)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000485 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000004d4),
    .Q(sig00000579)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000486 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000004d3),
    .Q(sig0000057a)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000487 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000569),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000508)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000488 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000056a),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000507)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000489 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000056b),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000506)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000048a (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000056c),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000505)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000048b (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000056d),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000504)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000048c (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000056e),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000503)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000048d (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000056f),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000502)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000048e (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000570),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000501)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000048f (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000571),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000500)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000490 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000572),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000004ff)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000491 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000573),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000004fe)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000492 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000574),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000004fd)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000493 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000575),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000004fc)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000494 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000576),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000004fb)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000495 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000577),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000004fa)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000496 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000578),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000004f9)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000497 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000579),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000004f8)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000498 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000057a),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000004f7)
  );
  XORCY   blk00000499 (
    .CI(sig0000059f),
    .LI(sig0000059d),
    .O(sig0000057b)
  );
  XORCY   blk0000049a (
    .CI(sig000005a0),
    .LI(sig0000058d),
    .O(sig0000057c)
  );
  XORCY   blk0000049b (
    .CI(sig000005a1),
    .LI(sig0000058e),
    .O(sig0000057d)
  );
  XORCY   blk0000049c (
    .CI(sig000005a2),
    .LI(sig0000058f),
    .O(sig0000057e)
  );
  XORCY   blk0000049d (
    .CI(sig000005a3),
    .LI(sig00000590),
    .O(sig0000057f)
  );
  XORCY   blk0000049e (
    .CI(sig000005a4),
    .LI(sig00000591),
    .O(sig00000580)
  );
  XORCY   blk0000049f (
    .CI(sig000005a5),
    .LI(sig00000592),
    .O(sig00000581)
  );
  XORCY   blk000004a0 (
    .CI(sig000005a6),
    .LI(sig00000593),
    .O(sig00000582)
  );
  XORCY   blk000004a1 (
    .CI(sig000005a7),
    .LI(sig00000594),
    .O(sig00000583)
  );
  XORCY   blk000004a2 (
    .CI(sig000005a8),
    .LI(sig00000595),
    .O(sig00000584)
  );
  XORCY   blk000004a3 (
    .CI(sig000005a9),
    .LI(sig00000596),
    .O(sig00000585)
  );
  XORCY   blk000004a4 (
    .CI(sig000005aa),
    .LI(sig00000597),
    .O(sig00000586)
  );
  XORCY   blk000004a5 (
    .CI(sig000005ab),
    .LI(sig00000598),
    .O(sig00000587)
  );
  XORCY   blk000004a6 (
    .CI(sig000005ac),
    .LI(sig00000599),
    .O(sig00000588)
  );
  XORCY   blk000004a7 (
    .CI(sig000005ad),
    .LI(sig0000059a),
    .O(sig00000589)
  );
  XORCY   blk000004a8 (
    .CI(sig000005ae),
    .LI(sig0000059b),
    .O(sig0000058a)
  );
  XORCY   blk000004a9 (
    .CI(sig000005af),
    .LI(sig0000059c),
    .O(sig0000058b)
  );
  XORCY   blk000004aa (
    .CI(sig00000344),
    .LI(sig0000059e),
    .O(sig0000058c)
  );
  MUXCY   blk000004ab (
    .CI(sig000005a0),
    .DI(sig00000507),
    .S(sig0000058d),
    .O(sig0000059f)
  );
  MUXCY   blk000004ac (
    .CI(sig000005a1),
    .DI(sig00000506),
    .S(sig0000058e),
    .O(sig000005a0)
  );
  MUXCY   blk000004ad (
    .CI(sig000005a2),
    .DI(sig00000505),
    .S(sig0000058f),
    .O(sig000005a1)
  );
  MUXCY   blk000004ae (
    .CI(sig000005a3),
    .DI(sig00000504),
    .S(sig00000590),
    .O(sig000005a2)
  );
  MUXCY   blk000004af (
    .CI(sig000005a4),
    .DI(sig00000503),
    .S(sig00000591),
    .O(sig000005a3)
  );
  MUXCY   blk000004b0 (
    .CI(sig000005a5),
    .DI(sig00000502),
    .S(sig00000592),
    .O(sig000005a4)
  );
  MUXCY   blk000004b1 (
    .CI(sig000005a6),
    .DI(sig00000501),
    .S(sig00000593),
    .O(sig000005a5)
  );
  MUXCY   blk000004b2 (
    .CI(sig000005a7),
    .DI(sig00000500),
    .S(sig00000594),
    .O(sig000005a6)
  );
  MUXCY   blk000004b3 (
    .CI(sig000005a8),
    .DI(sig000004ff),
    .S(sig00000595),
    .O(sig000005a7)
  );
  MUXCY   blk000004b4 (
    .CI(sig000005a9),
    .DI(sig000004fe),
    .S(sig00000596),
    .O(sig000005a8)
  );
  MUXCY   blk000004b5 (
    .CI(sig000005aa),
    .DI(sig000004fd),
    .S(sig00000597),
    .O(sig000005a9)
  );
  MUXCY   blk000004b6 (
    .CI(sig000005ab),
    .DI(sig000004fc),
    .S(sig00000598),
    .O(sig000005aa)
  );
  MUXCY   blk000004b7 (
    .CI(sig000005ac),
    .DI(sig000004fb),
    .S(sig00000599),
    .O(sig000005ab)
  );
  MUXCY   blk000004b8 (
    .CI(sig000005ad),
    .DI(sig000004fa),
    .S(sig0000059a),
    .O(sig000005ac)
  );
  MUXCY   blk000004b9 (
    .CI(sig000005ae),
    .DI(sig000004f9),
    .S(sig0000059b),
    .O(sig000005ad)
  );
  MUXCY   blk000004ba (
    .CI(sig000005af),
    .DI(sig000004f8),
    .S(sig0000059c),
    .O(sig000005ae)
  );
  MUXCY   blk000004bb (
    .CI(sig00000344),
    .DI(sig000004f7),
    .S(sig0000059e),
    .O(sig000005af)
  );
  XORCY   blk000004bc (
    .CI(sig000005d4),
    .LI(sig000005d2),
    .O(sig000005b0)
  );
  XORCY   blk000004bd (
    .CI(sig000005d5),
    .LI(sig000005c2),
    .O(sig000005b1)
  );
  XORCY   blk000004be (
    .CI(sig000005d6),
    .LI(sig000005c3),
    .O(sig000005b2)
  );
  XORCY   blk000004bf (
    .CI(sig000005d7),
    .LI(sig000005c4),
    .O(sig000005b3)
  );
  XORCY   blk000004c0 (
    .CI(sig000005d8),
    .LI(sig000005c5),
    .O(sig000005b4)
  );
  XORCY   blk000004c1 (
    .CI(sig000005d9),
    .LI(sig000005c6),
    .O(sig000005b5)
  );
  XORCY   blk000004c2 (
    .CI(sig000005da),
    .LI(sig000005c7),
    .O(sig000005b6)
  );
  XORCY   blk000004c3 (
    .CI(sig000005db),
    .LI(sig000005c8),
    .O(sig000005b7)
  );
  XORCY   blk000004c4 (
    .CI(sig000005dc),
    .LI(sig000005c9),
    .O(sig000005b8)
  );
  XORCY   blk000004c5 (
    .CI(sig000005dd),
    .LI(sig000005ca),
    .O(sig000005b9)
  );
  XORCY   blk000004c6 (
    .CI(sig000005de),
    .LI(sig000005cb),
    .O(sig000005ba)
  );
  XORCY   blk000004c7 (
    .CI(sig000005df),
    .LI(sig000005cc),
    .O(sig000005bb)
  );
  XORCY   blk000004c8 (
    .CI(sig000005e0),
    .LI(sig000005cd),
    .O(sig000005bc)
  );
  XORCY   blk000004c9 (
    .CI(sig000005e1),
    .LI(sig000005ce),
    .O(sig000005bd)
  );
  XORCY   blk000004ca (
    .CI(sig000005e2),
    .LI(sig000005cf),
    .O(sig000005be)
  );
  XORCY   blk000004cb (
    .CI(sig000005e3),
    .LI(sig000005d0),
    .O(sig000005bf)
  );
  XORCY   blk000004cc (
    .CI(sig000005e4),
    .LI(sig000005d1),
    .O(sig000005c0)
  );
  XORCY   blk000004cd (
    .CI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .LI(sig000005d3),
    .O(sig000005c1)
  );
  MUXCY   blk000004ce (
    .CI(sig000005d5),
    .DI(sig00000507),
    .S(sig000005c2),
    .O(sig000005d4)
  );
  MUXCY   blk000004cf (
    .CI(sig000005d6),
    .DI(sig00000506),
    .S(sig000005c3),
    .O(sig000005d5)
  );
  MUXCY   blk000004d0 (
    .CI(sig000005d7),
    .DI(sig00000505),
    .S(sig000005c4),
    .O(sig000005d6)
  );
  MUXCY   blk000004d1 (
    .CI(sig000005d8),
    .DI(sig00000504),
    .S(sig000005c5),
    .O(sig000005d7)
  );
  MUXCY   blk000004d2 (
    .CI(sig000005d9),
    .DI(sig00000503),
    .S(sig000005c6),
    .O(sig000005d8)
  );
  MUXCY   blk000004d3 (
    .CI(sig000005da),
    .DI(sig00000502),
    .S(sig000005c7),
    .O(sig000005d9)
  );
  MUXCY   blk000004d4 (
    .CI(sig000005db),
    .DI(sig00000501),
    .S(sig000005c8),
    .O(sig000005da)
  );
  MUXCY   blk000004d5 (
    .CI(sig000005dc),
    .DI(sig00000500),
    .S(sig000005c9),
    .O(sig000005db)
  );
  MUXCY   blk000004d6 (
    .CI(sig000005dd),
    .DI(sig000004ff),
    .S(sig000005ca),
    .O(sig000005dc)
  );
  MUXCY   blk000004d7 (
    .CI(sig000005de),
    .DI(sig000004fe),
    .S(sig000005cb),
    .O(sig000005dd)
  );
  MUXCY   blk000004d8 (
    .CI(sig000005df),
    .DI(sig000004fd),
    .S(sig000005cc),
    .O(sig000005de)
  );
  MUXCY   blk000004d9 (
    .CI(sig000005e0),
    .DI(sig000004fc),
    .S(sig000005cd),
    .O(sig000005df)
  );
  MUXCY   blk000004da (
    .CI(sig000005e1),
    .DI(sig000004fb),
    .S(sig000005ce),
    .O(sig000005e0)
  );
  MUXCY   blk000004db (
    .CI(sig000005e2),
    .DI(sig000004fa),
    .S(sig000005cf),
    .O(sig000005e1)
  );
  MUXCY   blk000004dc (
    .CI(sig000005e3),
    .DI(sig000004f9),
    .S(sig000005d0),
    .O(sig000005e2)
  );
  MUXCY   blk000004dd (
    .CI(sig000005e4),
    .DI(sig000004f8),
    .S(sig000005d1),
    .O(sig000005e3)
  );
  MUXCY   blk000004de (
    .CI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .DI(sig000004f7),
    .S(sig000005d3),
    .O(sig000005e4)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000004df (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000005b0),
    .Q(sig000004c0)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000004e0 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000005b1),
    .Q(sig000004bf)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000004e1 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000005b2),
    .Q(sig000004be)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000004e2 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000005b3),
    .Q(sig000004bd)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000004e3 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000005b4),
    .Q(sig000004bc)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000004e4 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000005b5),
    .Q(sig000004bb)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000004e5 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000005b6),
    .Q(sig000004ba)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000004e6 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000005b7),
    .Q(sig000004b9)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000004e7 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000005b8),
    .Q(sig000004b8)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000004e8 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000005b9),
    .Q(sig000004b7)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000004e9 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000005ba),
    .Q(sig000004b6)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000004ea (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000005bb),
    .Q(sig000004b5)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000004eb (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000005bc),
    .Q(sig000004b4)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000004ec (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000005bd),
    .Q(sig000004b3)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000004ed (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000005be),
    .Q(sig000004b2)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000004ee (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000005bf),
    .Q(sig000004b1)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000004ef (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000005c0),
    .Q(sig000004b0)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000004f0 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000005c1),
    .Q(sig000004af)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000004f1 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000057b),
    .Q(sig000004ae)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000004f2 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000057c),
    .Q(sig000004ad)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000004f3 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000057d),
    .Q(sig000004ac)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000004f4 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000057e),
    .Q(sig000004ab)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000004f5 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000057f),
    .Q(sig000004aa)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000004f6 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000580),
    .Q(sig000004a9)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000004f7 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000581),
    .Q(sig000004a8)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000004f8 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000582),
    .Q(sig000004a7)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000004f9 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000583),
    .Q(sig000004a6)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000004fa (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000584),
    .Q(sig000004a5)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000004fb (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000585),
    .Q(sig000004a4)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000004fc (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000586),
    .Q(sig000004a3)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000004fd (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000587),
    .Q(sig000004a2)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000004fe (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000588),
    .Q(sig000004a1)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000004ff (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000589),
    .Q(sig000004a0)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000500 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000058a),
    .Q(sig0000049f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000501 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000058b),
    .Q(sig0000049e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000502 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000058c),
    .Q(sig0000049d)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000050c (
    .C(aclk),
    .D(sig000001b1),
    .Q(sig000005f1)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000050d (
    .C(aclk),
    .D(sig000001b0),
    .Q(sig000005f0)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000050e (
    .C(aclk),
    .D(sig000001b3),
    .Q(sig000005f3)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000050f (
    .C(aclk),
    .D(sig000001b2),
    .Q(sig000005f2)
  );
  XORCY   blk00000510 (
    .CI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .LI(sig00000c62),
    .O(NLW_blk00000510_O_UNCONNECTED)
  );
  XORCY   blk00000511 (
    .CI(sig000005f8),
    .LI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .O(sig000005f4)
  );
  XORCY   blk00000512 (
    .CI(sig000005f9),
    .LI(sig00000c61),
    .O(sig000005f5)
  );
  XORCY   blk00000513 (
    .CI(sig000005fa),
    .LI(sig000005f7),
    .O(sig000005f6)
  );
  MUXCY   blk00000514 (
    .CI(sig000005f9),
    .DI(sig000001b3),
    .S(sig00000c61),
    .O(sig000005f8)
  );
  MUXCY   blk00000515 (
    .CI(sig000005fa),
    .DI(sig000001b2),
    .S(sig000005f7),
    .O(sig000005f9)
  );
  MUXCY   blk00000516 (
    .CI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig00000c62),
    .O(sig000005fa)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000517 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000005f6),
    .Q(sig000005ed)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000518 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000005f5),
    .Q(sig000005ee)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000519 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000005f4),
    .Q(sig000005ef)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk0000051a (
    .I0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .I1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .I2(sig000005f2),
    .I3(sig000005f2),
    .I4(sig000005f0),
    .I5(sig000005f1),
    .O(sig000005fb)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk0000051b (
    .I0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .I1(sig000005f2),
    .I2(sig000005f3),
    .I3(sig000005ed),
    .I4(sig000005f0),
    .I5(sig000005f1),
    .O(sig000005fc)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk0000051c (
    .I0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .I1(sig000005f3),
    .I2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .I3(sig000005ee),
    .I4(sig000005f0),
    .I5(sig000005f1),
    .O(sig000005fd)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk0000051d (
    .I0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .I1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .I2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .I3(sig000005ef),
    .I4(sig000005f0),
    .I5(sig000005f1),
    .O(sig000005fe)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000051e (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000005fb),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000005ea)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000051f (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000005fc),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000005eb)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000520 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000005fd),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000005ec)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000521 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000005fe),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000005e9)
  );
  DSP48E1 #(
    .ACASCREG ( 1 ),
    .ADREG ( 1 ),
    .ALUMODEREG ( 0 ),
    .AREG ( 1 ),
    .AUTORESET_PATDET ( "NO_RESET" ),
    .A_INPUT ( "DIRECT" ),
    .BCASCREG ( 2 ),
    .BREG ( 2 ),
    .B_INPUT ( "DIRECT" ),
    .CARRYINREG ( 0 ),
    .CARRYINSELREG ( 0 ),
    .CREG ( 1 ),
    .DREG ( 1 ),
    .INMODEREG ( 0 ),
    .MASK ( 48'h000000000000 ),
    .MREG ( 1 ),
    .OPMODEREG ( 0 ),
    .PATTERN ( 48'h000000000000 ),
    .PREG ( 1 ),
    .SEL_MASK ( "MASK" ),
    .SEL_PATTERN ( "PATTERN" ),
    .USE_DPORT ( "TRUE" ),
    .USE_MULT ( "MULTIPLY" ),
    .USE_PATTERN_DETECT ( "NO_PATDET" ),
    .USE_SIMD ( "ONE48" ))
  blk00000546 (
    .PATTERNBDETECT(NLW_blk00000546_PATTERNBDETECT_UNCONNECTED),
    .RSTC(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CEB1(sig00000344),
    .CEAD(sig00000344),
    .MULTSIGNOUT(NLW_blk00000546_MULTSIGNOUT_UNCONNECTED),
    .CEC(sig00000344),
    .RSTM(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .MULTSIGNIN(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CEB2(sig00000344),
    .RSTCTRL(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CEP(sig00000344),
    .CARRYCASCOUT(NLW_blk00000546_CARRYCASCOUT_UNCONNECTED),
    .RSTA(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CECARRYIN(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .UNDERFLOW(NLW_blk00000546_UNDERFLOW_UNCONNECTED),
    .PATTERNDETECT(NLW_blk00000546_PATTERNDETECT_UNCONNECTED),
    .RSTALUMODE(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .RSTALLCARRYIN(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CED(sig00000344),
    .RSTD(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CEALUMODE(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CEA2(sig00000344),
    .CLK(aclk),
    .CEA1(sig00000344),
    .RSTB(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .OVERFLOW(NLW_blk00000546_OVERFLOW_UNCONNECTED),
    .CECTRL(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CEM(sig00000344),
    .CARRYIN(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CARRYCASCIN(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .RSTINMODE(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CEINMODE(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .RSTP(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .ACOUT({\NLW_blk00000546_ACOUT<29>_UNCONNECTED , \NLW_blk00000546_ACOUT<28>_UNCONNECTED , \NLW_blk00000546_ACOUT<27>_UNCONNECTED ,
\NLW_blk00000546_ACOUT<26>_UNCONNECTED , \NLW_blk00000546_ACOUT<25>_UNCONNECTED , \NLW_blk00000546_ACOUT<24>_UNCONNECTED ,
\NLW_blk00000546_ACOUT<23>_UNCONNECTED , \NLW_blk00000546_ACOUT<22>_UNCONNECTED , \NLW_blk00000546_ACOUT<21>_UNCONNECTED ,
\NLW_blk00000546_ACOUT<20>_UNCONNECTED , \NLW_blk00000546_ACOUT<19>_UNCONNECTED , \NLW_blk00000546_ACOUT<18>_UNCONNECTED ,
\NLW_blk00000546_ACOUT<17>_UNCONNECTED , \NLW_blk00000546_ACOUT<16>_UNCONNECTED , \NLW_blk00000546_ACOUT<15>_UNCONNECTED ,
\NLW_blk00000546_ACOUT<14>_UNCONNECTED , \NLW_blk00000546_ACOUT<13>_UNCONNECTED , \NLW_blk00000546_ACOUT<12>_UNCONNECTED ,
\NLW_blk00000546_ACOUT<11>_UNCONNECTED , \NLW_blk00000546_ACOUT<10>_UNCONNECTED , \NLW_blk00000546_ACOUT<9>_UNCONNECTED ,
\NLW_blk00000546_ACOUT<8>_UNCONNECTED , \NLW_blk00000546_ACOUT<7>_UNCONNECTED , \NLW_blk00000546_ACOUT<6>_UNCONNECTED ,
\NLW_blk00000546_ACOUT<5>_UNCONNECTED , \NLW_blk00000546_ACOUT<4>_UNCONNECTED , \NLW_blk00000546_ACOUT<3>_UNCONNECTED ,
\NLW_blk00000546_ACOUT<2>_UNCONNECTED , \NLW_blk00000546_ACOUT<1>_UNCONNECTED , \NLW_blk00000546_ACOUT<0>_UNCONNECTED }),
    .OPMODE({\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1], sig00000344, sig00000344,
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1], sig00000344,
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1], sig00000344}),
    .PCIN({\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]}),
    .ALUMODE({\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]}),
    .C({sig0000065c, sig0000065c, sig0000065c, sig0000065c, sig0000065c, sig0000065c, sig0000065c, sig0000065c, sig0000065c, sig0000065c, sig0000065c
, sig0000065c, sig0000065c, sig0000065d, sig0000065e, sig0000065f, sig00000660, sig00000661, sig00000662, sig00000663, sig00000664, sig00000665,
sig00000666, sig00000667, sig00000668, sig00000669, sig0000066a, sig0000066b, sig0000066c, sig0000066d, sig0000066e, sig0000066f, sig00000670,
sig00000671, sig00000672, sig00000673, sig00000674, sig00000675, sig00000676, sig00000677, sig00000678, sig00000679, sig0000067a, sig0000067b,
sig0000067c, sig0000067d, sig0000067e, sig0000067f}),
    .CARRYOUT({\NLW_blk00000546_CARRYOUT<3>_UNCONNECTED , \NLW_blk00000546_CARRYOUT<2>_UNCONNECTED , \NLW_blk00000546_CARRYOUT<1>_UNCONNECTED ,
\NLW_blk00000546_CARRYOUT<0>_UNCONNECTED }),
    .INMODE({\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1], sig00000344, sig00000344,
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]}),
    .BCIN({\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]}),
    .B({sig00000643, sig00000644, sig00000645, sig00000646, sig00000647, sig00000648, sig00000649, sig0000064a, sig0000064b, sig0000064c, sig0000064d
, sig0000064e, sig0000064f, sig00000650, sig00000651, sig00000652, sig00000653, sig00000654}),
    .BCOUT({\NLW_blk00000546_BCOUT<17>_UNCONNECTED , \NLW_blk00000546_BCOUT<16>_UNCONNECTED , \NLW_blk00000546_BCOUT<15>_UNCONNECTED ,
\NLW_blk00000546_BCOUT<14>_UNCONNECTED , \NLW_blk00000546_BCOUT<13>_UNCONNECTED , \NLW_blk00000546_BCOUT<12>_UNCONNECTED ,
\NLW_blk00000546_BCOUT<11>_UNCONNECTED , \NLW_blk00000546_BCOUT<10>_UNCONNECTED , \NLW_blk00000546_BCOUT<9>_UNCONNECTED ,
\NLW_blk00000546_BCOUT<8>_UNCONNECTED , \NLW_blk00000546_BCOUT<7>_UNCONNECTED , \NLW_blk00000546_BCOUT<6>_UNCONNECTED ,
\NLW_blk00000546_BCOUT<5>_UNCONNECTED , \NLW_blk00000546_BCOUT<4>_UNCONNECTED , \NLW_blk00000546_BCOUT<3>_UNCONNECTED ,
\NLW_blk00000546_BCOUT<2>_UNCONNECTED , \NLW_blk00000546_BCOUT<1>_UNCONNECTED , \NLW_blk00000546_BCOUT<0>_UNCONNECTED }),
    .D({sig00000758, sig00000758, sig00000758, sig00000758, sig00000758, sig00000758, sig00000758, sig00000758, sig00000758, sig00000757, sig00000756
, sig00000755, sig00000754, sig00000753, sig00000752, sig00000751, sig00000750, sig0000074f, sig0000074e, sig0000074d, sig0000074c, sig0000074b,
sig0000074a, sig00000749, \NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]}),
    .P({\NLW_blk00000546_P<47>_UNCONNECTED , \NLW_blk00000546_P<46>_UNCONNECTED , \NLW_blk00000546_P<45>_UNCONNECTED ,
\NLW_blk00000546_P<44>_UNCONNECTED , \NLW_blk00000546_P<43>_UNCONNECTED , sig000005ff, sig00000600, sig00000601, sig00000602, sig00000603, sig00000604
, sig00000605, sig00000606, sig00000607, sig0000017a, sig00000179, sig00000178, sig00000177, sig00000176, sig00000175, sig00000174, sig00000173,
sig00000172, sig00000171, sig00000170, sig0000016f, sig0000016e, sig0000016d, sig0000016c, sig0000016b, sig0000016a, sig00000169, sig00000168,
sig00000167, sig00000166, sig00000165, sig00000164, sig00000163, sig00000620, sig00000621, sig00000622, sig00000623, sig00000624, sig00000625,
sig00000626, sig00000627, sig00000628, sig00000629}),
    .A({\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1], sig0000062a, sig0000062a, sig0000062a, sig0000062a,
sig0000062a, sig0000062a, sig0000062a, sig0000062a, sig0000062a, sig00000633, sig00000634, sig00000635, sig00000636, sig00000637, sig00000638,
sig00000639, sig0000063a, sig0000063b, sig0000063c, sig0000063d, sig0000063e, sig0000063f, sig00000640, sig00000641,
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]}),
    .PCOUT({\NLW_blk00000546_PCOUT<47>_UNCONNECTED , \NLW_blk00000546_PCOUT<46>_UNCONNECTED , \NLW_blk00000546_PCOUT<45>_UNCONNECTED ,
\NLW_blk00000546_PCOUT<44>_UNCONNECTED , \NLW_blk00000546_PCOUT<43>_UNCONNECTED , \NLW_blk00000546_PCOUT<42>_UNCONNECTED ,
\NLW_blk00000546_PCOUT<41>_UNCONNECTED , \NLW_blk00000546_PCOUT<40>_UNCONNECTED , \NLW_blk00000546_PCOUT<39>_UNCONNECTED ,
\NLW_blk00000546_PCOUT<38>_UNCONNECTED , \NLW_blk00000546_PCOUT<37>_UNCONNECTED , \NLW_blk00000546_PCOUT<36>_UNCONNECTED ,
\NLW_blk00000546_PCOUT<35>_UNCONNECTED , \NLW_blk00000546_PCOUT<34>_UNCONNECTED , \NLW_blk00000546_PCOUT<33>_UNCONNECTED ,
\NLW_blk00000546_PCOUT<32>_UNCONNECTED , \NLW_blk00000546_PCOUT<31>_UNCONNECTED , \NLW_blk00000546_PCOUT<30>_UNCONNECTED ,
\NLW_blk00000546_PCOUT<29>_UNCONNECTED , \NLW_blk00000546_PCOUT<28>_UNCONNECTED , \NLW_blk00000546_PCOUT<27>_UNCONNECTED ,
\NLW_blk00000546_PCOUT<26>_UNCONNECTED , \NLW_blk00000546_PCOUT<25>_UNCONNECTED , \NLW_blk00000546_PCOUT<24>_UNCONNECTED ,
\NLW_blk00000546_PCOUT<23>_UNCONNECTED , \NLW_blk00000546_PCOUT<22>_UNCONNECTED , \NLW_blk00000546_PCOUT<21>_UNCONNECTED ,
\NLW_blk00000546_PCOUT<20>_UNCONNECTED , \NLW_blk00000546_PCOUT<19>_UNCONNECTED , \NLW_blk00000546_PCOUT<18>_UNCONNECTED ,
\NLW_blk00000546_PCOUT<17>_UNCONNECTED , \NLW_blk00000546_PCOUT<16>_UNCONNECTED , \NLW_blk00000546_PCOUT<15>_UNCONNECTED ,
\NLW_blk00000546_PCOUT<14>_UNCONNECTED , \NLW_blk00000546_PCOUT<13>_UNCONNECTED , \NLW_blk00000546_PCOUT<12>_UNCONNECTED ,
\NLW_blk00000546_PCOUT<11>_UNCONNECTED , \NLW_blk00000546_PCOUT<10>_UNCONNECTED , \NLW_blk00000546_PCOUT<9>_UNCONNECTED ,
\NLW_blk00000546_PCOUT<8>_UNCONNECTED , \NLW_blk00000546_PCOUT<7>_UNCONNECTED , \NLW_blk00000546_PCOUT<6>_UNCONNECTED ,
\NLW_blk00000546_PCOUT<5>_UNCONNECTED , \NLW_blk00000546_PCOUT<4>_UNCONNECTED , \NLW_blk00000546_PCOUT<3>_UNCONNECTED ,
\NLW_blk00000546_PCOUT<2>_UNCONNECTED , \NLW_blk00000546_PCOUT<1>_UNCONNECTED , \NLW_blk00000546_PCOUT<0>_UNCONNECTED }),
    .ACIN({\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]}),
    .CARRYINSEL({\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]})
  );
  DSP48E1 #(
    .ACASCREG ( 1 ),
    .ADREG ( 1 ),
    .ALUMODEREG ( 0 ),
    .AREG ( 1 ),
    .AUTORESET_PATDET ( "NO_RESET" ),
    .A_INPUT ( "DIRECT" ),
    .BCASCREG ( 2 ),
    .BREG ( 2 ),
    .B_INPUT ( "DIRECT" ),
    .CARRYINREG ( 0 ),
    .CARRYINSELREG ( 0 ),
    .CREG ( 0 ),
    .DREG ( 1 ),
    .INMODEREG ( 0 ),
    .MASK ( 48'h000000000000 ),
    .MREG ( 1 ),
    .OPMODEREG ( 0 ),
    .PATTERN ( 48'h000000000000 ),
    .PREG ( 1 ),
    .SEL_MASK ( "MASK" ),
    .SEL_PATTERN ( "PATTERN" ),
    .USE_DPORT ( "TRUE" ),
    .USE_MULT ( "MULTIPLY" ),
    .USE_PATTERN_DETECT ( "NO_PATDET" ),
    .USE_SIMD ( "ONE48" ))
  blk00000547 (
    .PATTERNBDETECT(NLW_blk00000547_PATTERNBDETECT_UNCONNECTED),
    .RSTC(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CEB1(sig00000344),
    .CEAD(sig00000344),
    .MULTSIGNOUT(NLW_blk00000547_MULTSIGNOUT_UNCONNECTED),
    .CEC(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .RSTM(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .MULTSIGNIN(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CEB2(sig00000344),
    .RSTCTRL(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CEP(sig00000344),
    .CARRYCASCOUT(NLW_blk00000547_CARRYCASCOUT_UNCONNECTED),
    .RSTA(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CECARRYIN(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .UNDERFLOW(NLW_blk00000547_UNDERFLOW_UNCONNECTED),
    .PATTERNDETECT(NLW_blk00000547_PATTERNDETECT_UNCONNECTED),
    .RSTALUMODE(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .RSTALLCARRYIN(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CED(sig00000344),
    .RSTD(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CEALUMODE(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CEA2(sig00000344),
    .CLK(aclk),
    .CEA1(sig00000344),
    .RSTB(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .OVERFLOW(NLW_blk00000547_OVERFLOW_UNCONNECTED),
    .CECTRL(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CEM(sig00000344),
    .CARRYIN(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CARRYCASCIN(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .RSTINMODE(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CEINMODE(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .RSTP(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .ACOUT({\NLW_blk00000547_ACOUT<29>_UNCONNECTED , \NLW_blk00000547_ACOUT<28>_UNCONNECTED , \NLW_blk00000547_ACOUT<27>_UNCONNECTED ,
\NLW_blk00000547_ACOUT<26>_UNCONNECTED , \NLW_blk00000547_ACOUT<25>_UNCONNECTED , \NLW_blk00000547_ACOUT<24>_UNCONNECTED ,
\NLW_blk00000547_ACOUT<23>_UNCONNECTED , \NLW_blk00000547_ACOUT<22>_UNCONNECTED , \NLW_blk00000547_ACOUT<21>_UNCONNECTED ,
\NLW_blk00000547_ACOUT<20>_UNCONNECTED , \NLW_blk00000547_ACOUT<19>_UNCONNECTED , \NLW_blk00000547_ACOUT<18>_UNCONNECTED ,
\NLW_blk00000547_ACOUT<17>_UNCONNECTED , \NLW_blk00000547_ACOUT<16>_UNCONNECTED , \NLW_blk00000547_ACOUT<15>_UNCONNECTED ,
\NLW_blk00000547_ACOUT<14>_UNCONNECTED , \NLW_blk00000547_ACOUT<13>_UNCONNECTED , \NLW_blk00000547_ACOUT<12>_UNCONNECTED ,
\NLW_blk00000547_ACOUT<11>_UNCONNECTED , \NLW_blk00000547_ACOUT<10>_UNCONNECTED , \NLW_blk00000547_ACOUT<9>_UNCONNECTED ,
\NLW_blk00000547_ACOUT<8>_UNCONNECTED , \NLW_blk00000547_ACOUT<7>_UNCONNECTED , \NLW_blk00000547_ACOUT<6>_UNCONNECTED ,
\NLW_blk00000547_ACOUT<5>_UNCONNECTED , \NLW_blk00000547_ACOUT<4>_UNCONNECTED , \NLW_blk00000547_ACOUT<3>_UNCONNECTED ,
\NLW_blk00000547_ACOUT<2>_UNCONNECTED , \NLW_blk00000547_ACOUT<1>_UNCONNECTED , \NLW_blk00000547_ACOUT<0>_UNCONNECTED }),
    .OPMODE({\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1], sig00000344, sig00000344,
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1], sig00000344,
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1], sig00000344}),
    .PCIN({\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]}),
    .ALUMODE({\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]}),
    .C({\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1], sig00000344, sig00000344, sig00000344, sig00000344,
sig00000344, sig00000344, sig00000344, sig00000344, sig00000344}),
    .CARRYOUT({\NLW_blk00000547_CARRYOUT<3>_UNCONNECTED , \NLW_blk00000547_CARRYOUT<2>_UNCONNECTED , \NLW_blk00000547_CARRYOUT<1>_UNCONNECTED ,
\NLW_blk00000547_CARRYOUT<0>_UNCONNECTED }),
    .INMODE({\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1], sig00000344,
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]}),
    .BCIN({\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]}),
    .B({sig00000699, sig00000699, sig0000069b, sig0000069c, sig0000069d, sig0000069e, sig0000069f, sig000006a0, sig000006a1, sig000006a2, sig000006a3
, sig000006a4, sig000006a5, sig000006a6, sig000006a7, sig000006a8, sig000006a9,
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]}),
    .BCOUT({\NLW_blk00000547_BCOUT<17>_UNCONNECTED , \NLW_blk00000547_BCOUT<16>_UNCONNECTED , \NLW_blk00000547_BCOUT<15>_UNCONNECTED ,
\NLW_blk00000547_BCOUT<14>_UNCONNECTED , \NLW_blk00000547_BCOUT<13>_UNCONNECTED , \NLW_blk00000547_BCOUT<12>_UNCONNECTED ,
\NLW_blk00000547_BCOUT<11>_UNCONNECTED , \NLW_blk00000547_BCOUT<10>_UNCONNECTED , \NLW_blk00000547_BCOUT<9>_UNCONNECTED ,
\NLW_blk00000547_BCOUT<8>_UNCONNECTED , \NLW_blk00000547_BCOUT<7>_UNCONNECTED , \NLW_blk00000547_BCOUT<6>_UNCONNECTED ,
\NLW_blk00000547_BCOUT<5>_UNCONNECTED , \NLW_blk00000547_BCOUT<4>_UNCONNECTED , \NLW_blk00000547_BCOUT<3>_UNCONNECTED ,
\NLW_blk00000547_BCOUT<2>_UNCONNECTED , \NLW_blk00000547_BCOUT<1>_UNCONNECTED , \NLW_blk00000547_BCOUT<0>_UNCONNECTED }),
    .D({sig0000079a, sig0000079a, sig0000079a, sig0000079a, sig0000079a, sig0000079a, sig0000079a, sig0000079a, sig00000799, sig00000798, sig00000797
, sig00000796, sig00000795, sig00000794, sig00000793, sig00000792, sig00000791, sig00000790, sig0000078f, sig0000078e, sig0000078d, sig0000078c,
sig0000078b, sig0000078a, sig00000789}),
    .P({\NLW_blk00000547_P<47>_UNCONNECTED , \NLW_blk00000547_P<46>_UNCONNECTED , \NLW_blk00000547_P<45>_UNCONNECTED ,
\NLW_blk00000547_P<44>_UNCONNECTED , \NLW_blk00000547_P<43>_UNCONNECTED , sig00000655, sig00000656, sig00000657, sig00000658, sig00000659, sig0000065a
, sig0000065b, sig0000065c, sig0000065d, sig0000065e, sig0000065f, sig00000660, sig00000661, sig00000662, sig00000663, sig00000664, sig00000665,
sig00000666, sig00000667, sig00000668, sig00000669, sig0000066a, sig0000066b, sig0000066c, sig0000066d, sig0000066e, sig0000066f, sig00000670,
sig00000671, sig00000672, sig00000673, sig00000674, sig00000675, sig00000676, sig00000677, sig00000678, sig00000679, sig0000067a, sig0000067b,
sig0000067c, sig0000067d, sig0000067e, sig0000067f}),
    .A({\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1], sig00000680, sig00000680, sig00000680, sig00000680,
sig00000680, sig00000680, sig00000680, sig00000680, sig00000688, sig00000689, sig0000068a, sig0000068b, sig0000068c, sig0000068d, sig0000068e,
sig0000068f, sig00000690, sig00000691, sig00000692, sig00000693, sig00000694, sig00000695, sig00000696, sig00000697, sig00000698}),
    .PCOUT({\NLW_blk00000547_PCOUT<47>_UNCONNECTED , \NLW_blk00000547_PCOUT<46>_UNCONNECTED , \NLW_blk00000547_PCOUT<45>_UNCONNECTED ,
\NLW_blk00000547_PCOUT<44>_UNCONNECTED , \NLW_blk00000547_PCOUT<43>_UNCONNECTED , \NLW_blk00000547_PCOUT<42>_UNCONNECTED ,
\NLW_blk00000547_PCOUT<41>_UNCONNECTED , \NLW_blk00000547_PCOUT<40>_UNCONNECTED , \NLW_blk00000547_PCOUT<39>_UNCONNECTED ,
\NLW_blk00000547_PCOUT<38>_UNCONNECTED , \NLW_blk00000547_PCOUT<37>_UNCONNECTED , \NLW_blk00000547_PCOUT<36>_UNCONNECTED ,
\NLW_blk00000547_PCOUT<35>_UNCONNECTED , \NLW_blk00000547_PCOUT<34>_UNCONNECTED , \NLW_blk00000547_PCOUT<33>_UNCONNECTED ,
\NLW_blk00000547_PCOUT<32>_UNCONNECTED , \NLW_blk00000547_PCOUT<31>_UNCONNECTED , \NLW_blk00000547_PCOUT<30>_UNCONNECTED ,
\NLW_blk00000547_PCOUT<29>_UNCONNECTED , \NLW_blk00000547_PCOUT<28>_UNCONNECTED , \NLW_blk00000547_PCOUT<27>_UNCONNECTED ,
\NLW_blk00000547_PCOUT<26>_UNCONNECTED , \NLW_blk00000547_PCOUT<25>_UNCONNECTED , \NLW_blk00000547_PCOUT<24>_UNCONNECTED ,
\NLW_blk00000547_PCOUT<23>_UNCONNECTED , \NLW_blk00000547_PCOUT<22>_UNCONNECTED , \NLW_blk00000547_PCOUT<21>_UNCONNECTED ,
\NLW_blk00000547_PCOUT<20>_UNCONNECTED , \NLW_blk00000547_PCOUT<19>_UNCONNECTED , \NLW_blk00000547_PCOUT<18>_UNCONNECTED ,
\NLW_blk00000547_PCOUT<17>_UNCONNECTED , \NLW_blk00000547_PCOUT<16>_UNCONNECTED , \NLW_blk00000547_PCOUT<15>_UNCONNECTED ,
\NLW_blk00000547_PCOUT<14>_UNCONNECTED , \NLW_blk00000547_PCOUT<13>_UNCONNECTED , \NLW_blk00000547_PCOUT<12>_UNCONNECTED ,
\NLW_blk00000547_PCOUT<11>_UNCONNECTED , \NLW_blk00000547_PCOUT<10>_UNCONNECTED , \NLW_blk00000547_PCOUT<9>_UNCONNECTED ,
\NLW_blk00000547_PCOUT<8>_UNCONNECTED , \NLW_blk00000547_PCOUT<7>_UNCONNECTED , \NLW_blk00000547_PCOUT<6>_UNCONNECTED ,
\NLW_blk00000547_PCOUT<5>_UNCONNECTED , \NLW_blk00000547_PCOUT<4>_UNCONNECTED , \NLW_blk00000547_PCOUT<3>_UNCONNECTED ,
\NLW_blk00000547_PCOUT<2>_UNCONNECTED , \NLW_blk00000547_PCOUT<1>_UNCONNECTED , \NLW_blk00000547_PCOUT<0>_UNCONNECTED }),
    .ACIN({\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]}),
    .CARRYINSEL({\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]})
  );
  DSP48E1 #(
    .ACASCREG ( 1 ),
    .ADREG ( 1 ),
    .ALUMODEREG ( 0 ),
    .AREG ( 1 ),
    .AUTORESET_PATDET ( "NO_RESET" ),
    .A_INPUT ( "DIRECT" ),
    .BCASCREG ( 2 ),
    .BREG ( 2 ),
    .B_INPUT ( "DIRECT" ),
    .CARRYINREG ( 0 ),
    .CARRYINSELREG ( 0 ),
    .CREG ( 1 ),
    .DREG ( 1 ),
    .INMODEREG ( 0 ),
    .MASK ( 48'h000000000000 ),
    .MREG ( 1 ),
    .OPMODEREG ( 0 ),
    .PATTERN ( 48'h000000000000 ),
    .PREG ( 1 ),
    .SEL_MASK ( "MASK" ),
    .SEL_PATTERN ( "PATTERN" ),
    .USE_DPORT ( "TRUE" ),
    .USE_MULT ( "MULTIPLY" ),
    .USE_PATTERN_DETECT ( "NO_PATDET" ),
    .USE_SIMD ( "ONE48" ))
  blk00000548 (
    .PATTERNBDETECT(NLW_blk00000548_PATTERNBDETECT_UNCONNECTED),
    .RSTC(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CEB1(sig00000344),
    .CEAD(sig00000344),
    .MULTSIGNOUT(NLW_blk00000548_MULTSIGNOUT_UNCONNECTED),
    .CEC(sig00000344),
    .RSTM(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .MULTSIGNIN(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CEB2(sig00000344),
    .RSTCTRL(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CEP(sig00000344),
    .CARRYCASCOUT(NLW_blk00000548_CARRYCASCOUT_UNCONNECTED),
    .RSTA(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CECARRYIN(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .UNDERFLOW(NLW_blk00000548_UNDERFLOW_UNCONNECTED),
    .PATTERNDETECT(NLW_blk00000548_PATTERNDETECT_UNCONNECTED),
    .RSTALUMODE(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .RSTALLCARRYIN(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CED(sig00000344),
    .RSTD(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CEALUMODE(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CEA2(sig00000344),
    .CLK(aclk),
    .CEA1(sig00000344),
    .RSTB(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .OVERFLOW(NLW_blk00000548_OVERFLOW_UNCONNECTED),
    .CECTRL(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CEM(sig00000344),
    .CARRYIN(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CARRYCASCIN(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .RSTINMODE(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CEINMODE(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .RSTP(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .ACOUT({\NLW_blk00000548_ACOUT<29>_UNCONNECTED , \NLW_blk00000548_ACOUT<28>_UNCONNECTED , \NLW_blk00000548_ACOUT<27>_UNCONNECTED ,
\NLW_blk00000548_ACOUT<26>_UNCONNECTED , \NLW_blk00000548_ACOUT<25>_UNCONNECTED , \NLW_blk00000548_ACOUT<24>_UNCONNECTED ,
\NLW_blk00000548_ACOUT<23>_UNCONNECTED , \NLW_blk00000548_ACOUT<22>_UNCONNECTED , \NLW_blk00000548_ACOUT<21>_UNCONNECTED ,
\NLW_blk00000548_ACOUT<20>_UNCONNECTED , \NLW_blk00000548_ACOUT<19>_UNCONNECTED , \NLW_blk00000548_ACOUT<18>_UNCONNECTED ,
\NLW_blk00000548_ACOUT<17>_UNCONNECTED , \NLW_blk00000548_ACOUT<16>_UNCONNECTED , \NLW_blk00000548_ACOUT<15>_UNCONNECTED ,
\NLW_blk00000548_ACOUT<14>_UNCONNECTED , \NLW_blk00000548_ACOUT<13>_UNCONNECTED , \NLW_blk00000548_ACOUT<12>_UNCONNECTED ,
\NLW_blk00000548_ACOUT<11>_UNCONNECTED , \NLW_blk00000548_ACOUT<10>_UNCONNECTED , \NLW_blk00000548_ACOUT<9>_UNCONNECTED ,
\NLW_blk00000548_ACOUT<8>_UNCONNECTED , \NLW_blk00000548_ACOUT<7>_UNCONNECTED , \NLW_blk00000548_ACOUT<6>_UNCONNECTED ,
\NLW_blk00000548_ACOUT<5>_UNCONNECTED , \NLW_blk00000548_ACOUT<4>_UNCONNECTED , \NLW_blk00000548_ACOUT<3>_UNCONNECTED ,
\NLW_blk00000548_ACOUT<2>_UNCONNECTED , \NLW_blk00000548_ACOUT<1>_UNCONNECTED , \NLW_blk00000548_ACOUT<0>_UNCONNECTED }),
    .OPMODE({\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1], sig00000344, sig00000344,
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1], sig00000344,
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1], sig00000344}),
    .PCIN({\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]}),
    .ALUMODE({\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1], sig00000344, sig00000344}),
    .C({sig0000065c, sig0000065c, sig0000065c, sig0000065c, sig0000065c, sig0000065c, sig0000065c, sig0000065c, sig0000065c, sig0000065c, sig0000065c
, sig0000065c, sig0000065c, sig0000065d, sig0000065e, sig0000065f, sig00000660, sig00000661, sig00000662, sig00000663, sig00000664, sig00000665,
sig00000666, sig00000667, sig00000668, sig00000669, sig0000066a, sig0000066b, sig0000066c, sig0000066d, sig0000066e, sig0000066f, sig00000670,
sig00000671, sig00000672, sig00000673, sig00000674, sig00000675, sig00000676, sig00000677, sig00000678, sig00000679, sig0000067a, sig0000067b,
sig0000067c, sig0000067d, sig0000067e, sig0000067f}),
    .CARRYOUT({\NLW_blk00000548_CARRYOUT<3>_UNCONNECTED , \NLW_blk00000548_CARRYOUT<2>_UNCONNECTED , \NLW_blk00000548_CARRYOUT<1>_UNCONNECTED ,
\NLW_blk00000548_CARRYOUT<0>_UNCONNECTED }),
    .INMODE({\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1], sig00000344,
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]}),
    .BCIN({\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]}),
    .B({sig000006ef, sig000006f0, sig000006f1, sig000006f2, sig000006f3, sig000006f4, sig000006f5, sig000006f6, sig000006f7, sig000006f8, sig000006f9
, sig000006fa, sig000006fb, sig000006fc, sig000006fd, sig000006fe, sig000006ff, sig00000700}),
    .BCOUT({\NLW_blk00000548_BCOUT<17>_UNCONNECTED , \NLW_blk00000548_BCOUT<16>_UNCONNECTED , \NLW_blk00000548_BCOUT<15>_UNCONNECTED ,
\NLW_blk00000548_BCOUT<14>_UNCONNECTED , \NLW_blk00000548_BCOUT<13>_UNCONNECTED , \NLW_blk00000548_BCOUT<12>_UNCONNECTED ,
\NLW_blk00000548_BCOUT<11>_UNCONNECTED , \NLW_blk00000548_BCOUT<10>_UNCONNECTED , \NLW_blk00000548_BCOUT<9>_UNCONNECTED ,
\NLW_blk00000548_BCOUT<8>_UNCONNECTED , \NLW_blk00000548_BCOUT<7>_UNCONNECTED , \NLW_blk00000548_BCOUT<6>_UNCONNECTED ,
\NLW_blk00000548_BCOUT<5>_UNCONNECTED , \NLW_blk00000548_BCOUT<4>_UNCONNECTED , \NLW_blk00000548_BCOUT<3>_UNCONNECTED ,
\NLW_blk00000548_BCOUT<2>_UNCONNECTED , \NLW_blk00000548_BCOUT<1>_UNCONNECTED , \NLW_blk00000548_BCOUT<0>_UNCONNECTED }),
    .D({sig00000758, sig00000758, sig00000758, sig00000758, sig00000758, sig00000758, sig00000758, sig00000758, sig00000758, sig00000757, sig00000756
, sig00000755, sig00000754, sig00000753, sig00000752, sig00000751, sig00000750, sig0000074f, sig0000074e, sig0000074d, sig0000074c, sig0000074b,
sig0000074a, sig00000749, \NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]}),
    .P({\NLW_blk00000548_P<47>_UNCONNECTED , \NLW_blk00000548_P<46>_UNCONNECTED , \NLW_blk00000548_P<45>_UNCONNECTED ,
\NLW_blk00000548_P<44>_UNCONNECTED , \NLW_blk00000548_P<43>_UNCONNECTED , sig000006ab, sig000006ac, sig000006ad, sig000006ae, sig000006af, sig000006b0
, sig000006b1, sig000006b2, sig000006b3, sig00000192, sig00000191, sig00000190, sig0000018f, sig0000018e, sig0000018d, sig0000018c, sig0000018b,
sig0000018a, sig00000189, sig00000188, sig00000187, sig00000186, sig00000185, sig00000184, sig00000183, sig00000182, sig00000181, sig00000180,
sig0000017f, sig0000017e, sig0000017d, sig0000017c, sig0000017b, sig000006cc, sig000006cd, sig000006ce, sig000006cf, sig000006d0, sig000006d1,
sig000006d2, sig000006d3, sig000006d4, sig000006d5}),
    .A({\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1], sig0000062a, sig0000062a, sig0000062a, sig0000062a,
sig0000062a, sig0000062a, sig0000062a, sig0000062a, sig0000062a, sig00000633, sig00000634, sig00000635, sig00000636, sig00000637, sig00000638,
sig00000639, sig0000063a, sig0000063b, sig0000063c, sig0000063d, sig0000063e, sig0000063f, sig00000640, sig00000641,
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]}),
    .PCOUT({\NLW_blk00000548_PCOUT<47>_UNCONNECTED , \NLW_blk00000548_PCOUT<46>_UNCONNECTED , \NLW_blk00000548_PCOUT<45>_UNCONNECTED ,
\NLW_blk00000548_PCOUT<44>_UNCONNECTED , \NLW_blk00000548_PCOUT<43>_UNCONNECTED , \NLW_blk00000548_PCOUT<42>_UNCONNECTED ,
\NLW_blk00000548_PCOUT<41>_UNCONNECTED , \NLW_blk00000548_PCOUT<40>_UNCONNECTED , \NLW_blk00000548_PCOUT<39>_UNCONNECTED ,
\NLW_blk00000548_PCOUT<38>_UNCONNECTED , \NLW_blk00000548_PCOUT<37>_UNCONNECTED , \NLW_blk00000548_PCOUT<36>_UNCONNECTED ,
\NLW_blk00000548_PCOUT<35>_UNCONNECTED , \NLW_blk00000548_PCOUT<34>_UNCONNECTED , \NLW_blk00000548_PCOUT<33>_UNCONNECTED ,
\NLW_blk00000548_PCOUT<32>_UNCONNECTED , \NLW_blk00000548_PCOUT<31>_UNCONNECTED , \NLW_blk00000548_PCOUT<30>_UNCONNECTED ,
\NLW_blk00000548_PCOUT<29>_UNCONNECTED , \NLW_blk00000548_PCOUT<28>_UNCONNECTED , \NLW_blk00000548_PCOUT<27>_UNCONNECTED ,
\NLW_blk00000548_PCOUT<26>_UNCONNECTED , \NLW_blk00000548_PCOUT<25>_UNCONNECTED , \NLW_blk00000548_PCOUT<24>_UNCONNECTED ,
\NLW_blk00000548_PCOUT<23>_UNCONNECTED , \NLW_blk00000548_PCOUT<22>_UNCONNECTED , \NLW_blk00000548_PCOUT<21>_UNCONNECTED ,
\NLW_blk00000548_PCOUT<20>_UNCONNECTED , \NLW_blk00000548_PCOUT<19>_UNCONNECTED , \NLW_blk00000548_PCOUT<18>_UNCONNECTED ,
\NLW_blk00000548_PCOUT<17>_UNCONNECTED , \NLW_blk00000548_PCOUT<16>_UNCONNECTED , \NLW_blk00000548_PCOUT<15>_UNCONNECTED ,
\NLW_blk00000548_PCOUT<14>_UNCONNECTED , \NLW_blk00000548_PCOUT<13>_UNCONNECTED , \NLW_blk00000548_PCOUT<12>_UNCONNECTED ,
\NLW_blk00000548_PCOUT<11>_UNCONNECTED , \NLW_blk00000548_PCOUT<10>_UNCONNECTED , \NLW_blk00000548_PCOUT<9>_UNCONNECTED ,
\NLW_blk00000548_PCOUT<8>_UNCONNECTED , \NLW_blk00000548_PCOUT<7>_UNCONNECTED , \NLW_blk00000548_PCOUT<6>_UNCONNECTED ,
\NLW_blk00000548_PCOUT<5>_UNCONNECTED , \NLW_blk00000548_PCOUT<4>_UNCONNECTED , \NLW_blk00000548_PCOUT<3>_UNCONNECTED ,
\NLW_blk00000548_PCOUT<2>_UNCONNECTED , \NLW_blk00000548_PCOUT<1>_UNCONNECTED , \NLW_blk00000548_PCOUT<0>_UNCONNECTED }),
    .ACIN({\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]}),
    .CARRYINSEL({\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1],
\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]})
  );
  XORCY   blk00000549 (
    .CI(sig000007ad),
    .LI(sig00000344),
    .O(sig00000806)
  );
  XORCY   blk0000054a (
    .CI(sig000007af),
    .LI(sig000007ae),
    .O(sig00000805)
  );
  MUXCY   blk0000054b (
    .CI(sig000007af),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig000007ae),
    .O(sig000007ad)
  );
  XORCY   blk0000054c (
    .CI(sig000007b1),
    .LI(sig000007b0),
    .O(sig00000804)
  );
  MUXCY   blk0000054d (
    .CI(sig000007b1),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig000007b0),
    .O(sig000007af)
  );
  XORCY   blk0000054e (
    .CI(sig000007b3),
    .LI(sig000007b2),
    .O(sig00000803)
  );
  MUXCY   blk0000054f (
    .CI(sig000007b3),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig000007b2),
    .O(sig000007b1)
  );
  XORCY   blk00000550 (
    .CI(sig000007b5),
    .LI(sig000007b4),
    .O(sig00000802)
  );
  MUXCY   blk00000551 (
    .CI(sig000007b5),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig000007b4),
    .O(sig000007b3)
  );
  XORCY   blk00000552 (
    .CI(sig000007b7),
    .LI(sig000007b6),
    .O(sig00000801)
  );
  MUXCY   blk00000553 (
    .CI(sig000007b7),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig000007b6),
    .O(sig000007b5)
  );
  XORCY   blk00000554 (
    .CI(sig000007b9),
    .LI(sig000007b8),
    .O(sig00000800)
  );
  MUXCY   blk00000555 (
    .CI(sig000007b9),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig000007b8),
    .O(sig000007b7)
  );
  XORCY   blk00000556 (
    .CI(sig000007bb),
    .LI(sig000007ba),
    .O(sig000007ff)
  );
  MUXCY   blk00000557 (
    .CI(sig000007bb),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig000007ba),
    .O(sig000007b9)
  );
  XORCY   blk00000558 (
    .CI(sig000007bc),
    .LI(sig00000344),
    .O(sig000007fe)
  );
  MUXCY   blk00000559 (
    .CI(sig000007bc),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig00000344),
    .O(sig000007bb)
  );
  XORCY   blk0000055a (
    .CI(sig000007be),
    .LI(sig000007bd),
    .O(sig000007fd)
  );
  MUXCY   blk0000055b (
    .CI(sig000007be),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig000007bd),
    .O(sig000007bc)
  );
  XORCY   blk0000055c (
    .CI(sig000007c0),
    .LI(sig000007bf),
    .O(sig000007fc)
  );
  MUXCY   blk0000055d (
    .CI(sig000007c0),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig000007bf),
    .O(sig000007be)
  );
  XORCY   blk0000055e (
    .CI(sig000007c2),
    .LI(sig000007c1),
    .O(sig000007fb)
  );
  MUXCY   blk0000055f (
    .CI(sig000007c2),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig000007c1),
    .O(sig000007c0)
  );
  XORCY   blk00000560 (
    .CI(sig000007c4),
    .LI(sig000007c3),
    .O(sig000007fa)
  );
  MUXCY   blk00000561 (
    .CI(sig000007c4),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig000007c3),
    .O(sig000007c2)
  );
  XORCY   blk00000562 (
    .CI(sig000007c6),
    .LI(sig000007c5),
    .O(sig000007f9)
  );
  MUXCY   blk00000563 (
    .CI(sig000007c6),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig000007c5),
    .O(sig000007c4)
  );
  XORCY   blk00000564 (
    .CI(sig000007c8),
    .LI(sig000007c7),
    .O(sig000007f8)
  );
  MUXCY   blk00000565 (
    .CI(sig000007c8),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig000007c7),
    .O(sig000007c6)
  );
  XORCY   blk00000566 (
    .CI(sig00000344),
    .LI(sig000007c9),
    .O(sig000007f7)
  );
  MUXCY   blk00000567 (
    .CI(sig00000344),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig000007c9),
    .O(sig000007c8)
  );
  XORCY   blk00000568 (
    .CI(sig000007ca),
    .LI(sig00000344),
    .O(sig00000826)
  );
  XORCY   blk00000569 (
    .CI(sig000007cc),
    .LI(sig000007cb),
    .O(sig00000825)
  );
  MUXCY   blk0000056a (
    .CI(sig000007cc),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig000007cb),
    .O(sig000007ca)
  );
  XORCY   blk0000056b (
    .CI(sig000007ce),
    .LI(sig000007cd),
    .O(sig00000824)
  );
  MUXCY   blk0000056c (
    .CI(sig000007ce),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig000007cd),
    .O(sig000007cc)
  );
  XORCY   blk0000056d (
    .CI(sig000007d0),
    .LI(sig000007cf),
    .O(sig00000823)
  );
  MUXCY   blk0000056e (
    .CI(sig000007d0),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig000007cf),
    .O(sig000007ce)
  );
  XORCY   blk0000056f (
    .CI(sig000007d2),
    .LI(sig000007d1),
    .O(sig00000822)
  );
  MUXCY   blk00000570 (
    .CI(sig000007d2),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig000007d1),
    .O(sig000007d0)
  );
  XORCY   blk00000571 (
    .CI(sig000007d4),
    .LI(sig000007d3),
    .O(sig00000821)
  );
  MUXCY   blk00000572 (
    .CI(sig000007d4),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig000007d3),
    .O(sig000007d2)
  );
  XORCY   blk00000573 (
    .CI(sig000007d6),
    .LI(sig000007d5),
    .O(sig00000820)
  );
  MUXCY   blk00000574 (
    .CI(sig000007d6),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig000007d5),
    .O(sig000007d4)
  );
  XORCY   blk00000575 (
    .CI(sig000007d8),
    .LI(sig000007d7),
    .O(sig0000081f)
  );
  MUXCY   blk00000576 (
    .CI(sig000007d8),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig000007d7),
    .O(sig000007d6)
  );
  XORCY   blk00000577 (
    .CI(sig000007d9),
    .LI(sig00000344),
    .O(sig0000081e)
  );
  MUXCY   blk00000578 (
    .CI(sig000007d9),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig00000344),
    .O(sig000007d8)
  );
  XORCY   blk00000579 (
    .CI(sig000007db),
    .LI(sig000007da),
    .O(sig0000081d)
  );
  MUXCY   blk0000057a (
    .CI(sig000007db),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig000007da),
    .O(sig000007d9)
  );
  XORCY   blk0000057b (
    .CI(sig000007dd),
    .LI(sig000007dc),
    .O(sig0000081c)
  );
  MUXCY   blk0000057c (
    .CI(sig000007dd),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig000007dc),
    .O(sig000007db)
  );
  XORCY   blk0000057d (
    .CI(sig000007df),
    .LI(sig000007de),
    .O(sig0000081b)
  );
  MUXCY   blk0000057e (
    .CI(sig000007df),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig000007de),
    .O(sig000007dd)
  );
  XORCY   blk0000057f (
    .CI(sig000007e1),
    .LI(sig000007e0),
    .O(sig0000081a)
  );
  MUXCY   blk00000580 (
    .CI(sig000007e1),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig000007e0),
    .O(sig000007df)
  );
  XORCY   blk00000581 (
    .CI(sig000007e3),
    .LI(sig000007e2),
    .O(sig00000819)
  );
  MUXCY   blk00000582 (
    .CI(sig000007e3),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig000007e2),
    .O(sig000007e1)
  );
  XORCY   blk00000583 (
    .CI(sig000007e5),
    .LI(sig000007e4),
    .O(sig00000818)
  );
  MUXCY   blk00000584 (
    .CI(sig000007e5),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig000007e4),
    .O(sig000007e3)
  );
  XORCY   blk00000585 (
    .CI(sig00000344),
    .LI(sig000007e6),
    .O(sig00000817)
  );
  MUXCY   blk00000586 (
    .CI(sig00000344),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig000007e6),
    .O(sig000007e5)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000587 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000816),
    .Q(sig00000699)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000588 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000815),
    .Q(sig0000069b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000589 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000814),
    .Q(sig0000069c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000058a (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000813),
    .Q(sig0000069d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000058b (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000812),
    .Q(sig0000069e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000058c (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000811),
    .Q(sig0000069f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000058d (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000810),
    .Q(sig000006a0)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000058e (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000080f),
    .Q(sig000006a1)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000058f (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000080e),
    .Q(sig000006a2)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000590 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000080d),
    .Q(sig000006a3)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000591 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000080c),
    .Q(sig000006a4)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000592 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000080b),
    .Q(sig000006a5)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000593 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000080a),
    .Q(sig000006a6)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000594 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000809),
    .Q(sig000006a7)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000595 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000808),
    .Q(sig000006a8)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000596 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000807),
    .Q(sig000006a9)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000597 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000007f6),
    .Q(sig00000778)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000598 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000007f5),
    .Q(sig00000777)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000599 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000007f4),
    .Q(sig00000776)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000059a (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000007f3),
    .Q(sig00000775)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000059b (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000007f2),
    .Q(sig00000774)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000059c (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000007f1),
    .Q(sig00000773)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000059d (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000007f0),
    .Q(sig00000772)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000059e (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000007ef),
    .Q(sig00000771)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000059f (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000007ee),
    .Q(sig00000770)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000005a0 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000007ed),
    .Q(sig0000076f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000005a1 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000007ec),
    .Q(sig0000076e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000005a2 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000007eb),
    .Q(sig0000076d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000005a3 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000007ea),
    .Q(sig0000076c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000005a4 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000007e9),
    .Q(sig0000076b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000005a5 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000007e8),
    .Q(sig0000076a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000005a6 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000007e7),
    .Q(sig00000769)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000005a7 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000001c5),
    .Q(sig0000079a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000005a8 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000001c4),
    .Q(sig00000799)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000005a9 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000001c3),
    .Q(sig00000798)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000005aa (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000001c2),
    .Q(sig00000797)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000005ab (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000001c1),
    .Q(sig00000796)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000005ac (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000001c0),
    .Q(sig00000795)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000005ad (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000001bf),
    .Q(sig00000794)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000005ae (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000001be),
    .Q(sig00000793)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000005af (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000001bd),
    .Q(sig00000792)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000005b0 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000001bc),
    .Q(sig00000791)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000005b1 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000001bb),
    .Q(sig00000790)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000005b2 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000001ba),
    .Q(sig0000078f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000005b3 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000001b9),
    .Q(sig0000078e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000005b4 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000001b8),
    .Q(sig0000078d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000005b5 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000001b7),
    .Q(sig0000078c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000005b6 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000001b6),
    .Q(sig0000078b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000005b7 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000001b5),
    .Q(sig0000078a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000005b8 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000001b4),
    .Q(sig00000789)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000005b9 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000001d7),
    .Q(sig00000680)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000005ba (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000001d6),
    .Q(sig00000688)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000005bb (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000001d5),
    .Q(sig00000689)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000005bc (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000001d4),
    .Q(sig0000068a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000005bd (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000001d3),
    .Q(sig0000068b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000005be (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000001d2),
    .Q(sig0000068c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000005bf (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000001d1),
    .Q(sig0000068d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000005c0 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000001d0),
    .Q(sig0000068e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000005c1 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000001cf),
    .Q(sig0000068f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000005c2 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000001ce),
    .Q(sig00000690)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000005c3 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000001cd),
    .Q(sig00000691)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000005c4 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000001cc),
    .Q(sig00000692)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000005c5 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000001cb),
    .Q(sig00000693)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000005c6 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000001ca),
    .Q(sig00000694)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000005c7 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000001c9),
    .Q(sig00000695)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000005c8 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000001c8),
    .Q(sig00000696)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000005c9 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000001c7),
    .Q(sig00000697)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000005ca (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000001c6),
    .Q(sig00000698)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000005d4 (
    .I0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .I1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .I2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .I3(sig0000017b),
    .I4(sig000001da),
    .I5(sig000001db),
    .O(sig00000827)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000005d5 (
    .I0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .I1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .I2(sig0000017b),
    .I3(sig0000017c),
    .I4(sig000001da),
    .I5(sig000001db),
    .O(sig00000828)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000005d6 (
    .I0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .I1(sig0000017b),
    .I2(sig0000017c),
    .I3(sig0000017d),
    .I4(sig000001da),
    .I5(sig000001db),
    .O(sig00000829)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000005d7 (
    .I0(sig0000017b),
    .I1(sig0000017c),
    .I2(sig0000017d),
    .I3(sig0000017e),
    .I4(sig000001da),
    .I5(sig000001db),
    .O(sig0000082a)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000005d8 (
    .I0(sig0000017c),
    .I1(sig0000017d),
    .I2(sig0000017e),
    .I3(sig0000017f),
    .I4(sig000001da),
    .I5(sig000001db),
    .O(sig0000082b)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000005d9 (
    .I0(sig0000017d),
    .I1(sig0000017e),
    .I2(sig0000017f),
    .I3(sig00000180),
    .I4(sig000001da),
    .I5(sig000001db),
    .O(sig0000082c)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000005da (
    .I0(sig0000017e),
    .I1(sig0000017f),
    .I2(sig00000180),
    .I3(sig00000181),
    .I4(sig000001da),
    .I5(sig000001db),
    .O(sig0000082d)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000005db (
    .I0(sig0000017f),
    .I1(sig00000180),
    .I2(sig00000181),
    .I3(sig00000182),
    .I4(sig000001da),
    .I5(sig000001db),
    .O(sig0000082e)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000005dc (
    .I0(sig00000180),
    .I1(sig00000181),
    .I2(sig00000182),
    .I3(sig00000183),
    .I4(sig000001da),
    .I5(sig000001db),
    .O(sig0000082f)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000005dd (
    .I0(sig00000181),
    .I1(sig00000182),
    .I2(sig00000183),
    .I3(sig00000184),
    .I4(sig000001da),
    .I5(sig000001db),
    .O(sig00000830)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000005de (
    .I0(sig00000182),
    .I1(sig00000183),
    .I2(sig00000184),
    .I3(sig00000185),
    .I4(sig000001da),
    .I5(sig000001db),
    .O(sig00000831)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000005df (
    .I0(sig00000183),
    .I1(sig00000184),
    .I2(sig00000185),
    .I3(sig00000186),
    .I4(sig000001da),
    .I5(sig000001db),
    .O(sig00000832)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000005e0 (
    .I0(sig00000184),
    .I1(sig00000185),
    .I2(sig00000186),
    .I3(sig00000187),
    .I4(sig000001da),
    .I5(sig000001db),
    .O(sig00000833)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000005e1 (
    .I0(sig00000185),
    .I1(sig00000186),
    .I2(sig00000187),
    .I3(sig00000188),
    .I4(sig000001da),
    .I5(sig000001db),
    .O(sig00000834)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000005e2 (
    .I0(sig00000186),
    .I1(sig00000187),
    .I2(sig00000188),
    .I3(sig00000189),
    .I4(sig000001da),
    .I5(sig000001db),
    .O(sig00000835)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000005e3 (
    .I0(sig00000187),
    .I1(sig00000188),
    .I2(sig00000189),
    .I3(sig0000018a),
    .I4(sig000001da),
    .I5(sig000001db),
    .O(sig00000836)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000005e4 (
    .I0(sig00000188),
    .I1(sig00000189),
    .I2(sig0000018a),
    .I3(sig0000018b),
    .I4(sig000001da),
    .I5(sig000001db),
    .O(sig00000837)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000005e5 (
    .I0(sig00000189),
    .I1(sig0000018a),
    .I2(sig0000018b),
    .I3(sig0000018c),
    .I4(sig000001da),
    .I5(sig000001db),
    .O(sig00000838)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000005e6 (
    .I0(sig0000018a),
    .I1(sig0000018b),
    .I2(sig0000018c),
    .I3(sig0000018d),
    .I4(sig000001da),
    .I5(sig000001db),
    .O(sig00000839)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000005e7 (
    .I0(sig0000018b),
    .I1(sig0000018c),
    .I2(sig0000018d),
    .I3(sig0000018e),
    .I4(sig000001da),
    .I5(sig000001db),
    .O(sig0000083a)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000005e8 (
    .I0(sig0000018c),
    .I1(sig0000018d),
    .I2(sig0000018e),
    .I3(sig0000018f),
    .I4(sig000001da),
    .I5(sig000001db),
    .O(sig0000083b)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000005e9 (
    .I0(sig0000018d),
    .I1(sig0000018e),
    .I2(sig0000018f),
    .I3(sig00000190),
    .I4(sig000001da),
    .I5(sig000001db),
    .O(sig0000083c)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000005ea (
    .I0(sig0000018e),
    .I1(sig0000018f),
    .I2(sig00000190),
    .I3(sig00000191),
    .I4(sig000001da),
    .I5(sig000001db),
    .O(sig0000083d)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000005eb (
    .I0(sig0000018f),
    .I1(sig00000190),
    .I2(sig00000191),
    .I3(sig00000192),
    .I4(sig000001da),
    .I5(sig000001db),
    .O(sig0000083e)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000005ec (
    .I0(sig00000190),
    .I1(sig00000191),
    .I2(sig00000192),
    .I3(sig00000192),
    .I4(sig000001da),
    .I5(sig000001db),
    .O(sig0000083f)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000005ed (
    .I0(sig00000191),
    .I1(sig00000192),
    .I2(sig00000192),
    .I3(sig00000192),
    .I4(sig000001da),
    .I5(sig000001db),
    .O(sig00000840)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000005ee (
    .I0(sig00000192),
    .I1(sig00000192),
    .I2(sig00000192),
    .I3(sig00000192),
    .I4(sig000001da),
    .I5(sig000001db),
    .O(sig00000841)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000005ef (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000827),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(NLW_blk000005ef_Q_UNCONNECTED)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000005f0 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000828),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(NLW_blk000005f0_Q_UNCONNECTED)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000005f1 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000829),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(NLW_blk000005f1_Q_UNCONNECTED)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000005f2 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000082a),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(NLW_blk000005f2_Q_UNCONNECTED)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000005f3 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000082b),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(NLW_blk000005f3_Q_UNCONNECTED)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000005f4 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000082c),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(NLW_blk000005f4_Q_UNCONNECTED)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000005f5 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000082d),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(NLW_blk000005f5_Q_UNCONNECTED)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000005f6 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000082e),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(NLW_blk000005f6_Q_UNCONNECTED)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000005f7 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000082f),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000000ae)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000005f8 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000830),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000000af)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000005f9 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000831),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000000b0)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000005fa (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000832),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000000b1)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000005fb (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000833),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000000b2)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000005fc (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000834),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000000b3)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000005fd (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000835),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000000b4)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000005fe (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000836),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000000b5)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000005ff (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000837),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000000b6)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000600 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000838),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000000b7)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000601 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000839),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000000b8)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000602 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000083a),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000000b9)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000603 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000083b),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000000ba)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000604 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000083c),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000000bb)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000605 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000083d),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000000bc)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000606 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000083e),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000000bd)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000607 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000083f),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(NLW_blk00000607_Q_UNCONNECTED)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000608 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000840),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(NLW_blk00000608_Q_UNCONNECTED)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000609 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000841),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(NLW_blk00000609_Q_UNCONNECTED)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk0000060a (
    .I0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .I1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .I2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .I3(sig00000163),
    .I4(sig000001da),
    .I5(sig000001db),
    .O(sig00000842)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk0000060b (
    .I0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .I1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .I2(sig00000163),
    .I3(sig00000164),
    .I4(sig000001da),
    .I5(sig000001db),
    .O(sig00000843)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk0000060c (
    .I0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .I1(sig00000163),
    .I2(sig00000164),
    .I3(sig00000165),
    .I4(sig000001da),
    .I5(sig000001db),
    .O(sig00000844)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk0000060d (
    .I0(sig00000163),
    .I1(sig00000164),
    .I2(sig00000165),
    .I3(sig00000166),
    .I4(sig000001da),
    .I5(sig000001db),
    .O(sig00000845)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk0000060e (
    .I0(sig00000164),
    .I1(sig00000165),
    .I2(sig00000166),
    .I3(sig00000167),
    .I4(sig000001da),
    .I5(sig000001db),
    .O(sig00000846)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk0000060f (
    .I0(sig00000165),
    .I1(sig00000166),
    .I2(sig00000167),
    .I3(sig00000168),
    .I4(sig000001da),
    .I5(sig000001db),
    .O(sig00000847)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk00000610 (
    .I0(sig00000166),
    .I1(sig00000167),
    .I2(sig00000168),
    .I3(sig00000169),
    .I4(sig000001da),
    .I5(sig000001db),
    .O(sig00000848)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk00000611 (
    .I0(sig00000167),
    .I1(sig00000168),
    .I2(sig00000169),
    .I3(sig0000016a),
    .I4(sig000001da),
    .I5(sig000001db),
    .O(sig00000849)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk00000612 (
    .I0(sig00000168),
    .I1(sig00000169),
    .I2(sig0000016a),
    .I3(sig0000016b),
    .I4(sig000001da),
    .I5(sig000001db),
    .O(sig0000084a)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk00000613 (
    .I0(sig00000169),
    .I1(sig0000016a),
    .I2(sig0000016b),
    .I3(sig0000016c),
    .I4(sig000001da),
    .I5(sig000001db),
    .O(sig0000084b)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk00000614 (
    .I0(sig0000016a),
    .I1(sig0000016b),
    .I2(sig0000016c),
    .I3(sig0000016d),
    .I4(sig000001da),
    .I5(sig000001db),
    .O(sig0000084c)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk00000615 (
    .I0(sig0000016b),
    .I1(sig0000016c),
    .I2(sig0000016d),
    .I3(sig0000016e),
    .I4(sig000001da),
    .I5(sig000001db),
    .O(sig0000084d)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk00000616 (
    .I0(sig0000016c),
    .I1(sig0000016d),
    .I2(sig0000016e),
    .I3(sig0000016f),
    .I4(sig000001da),
    .I5(sig000001db),
    .O(sig0000084e)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk00000617 (
    .I0(sig0000016d),
    .I1(sig0000016e),
    .I2(sig0000016f),
    .I3(sig00000170),
    .I4(sig000001da),
    .I5(sig000001db),
    .O(sig0000084f)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk00000618 (
    .I0(sig0000016e),
    .I1(sig0000016f),
    .I2(sig00000170),
    .I3(sig00000171),
    .I4(sig000001da),
    .I5(sig000001db),
    .O(sig00000850)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk00000619 (
    .I0(sig0000016f),
    .I1(sig00000170),
    .I2(sig00000171),
    .I3(sig00000172),
    .I4(sig000001da),
    .I5(sig000001db),
    .O(sig00000851)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk0000061a (
    .I0(sig00000170),
    .I1(sig00000171),
    .I2(sig00000172),
    .I3(sig00000173),
    .I4(sig000001da),
    .I5(sig000001db),
    .O(sig00000852)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk0000061b (
    .I0(sig00000171),
    .I1(sig00000172),
    .I2(sig00000173),
    .I3(sig00000174),
    .I4(sig000001da),
    .I5(sig000001db),
    .O(sig00000853)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk0000061c (
    .I0(sig00000172),
    .I1(sig00000173),
    .I2(sig00000174),
    .I3(sig00000175),
    .I4(sig000001da),
    .I5(sig000001db),
    .O(sig00000854)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk0000061d (
    .I0(sig00000173),
    .I1(sig00000174),
    .I2(sig00000175),
    .I3(sig00000176),
    .I4(sig000001da),
    .I5(sig000001db),
    .O(sig00000855)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk0000061e (
    .I0(sig00000174),
    .I1(sig00000175),
    .I2(sig00000176),
    .I3(sig00000177),
    .I4(sig000001da),
    .I5(sig000001db),
    .O(sig00000856)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk0000061f (
    .I0(sig00000175),
    .I1(sig00000176),
    .I2(sig00000177),
    .I3(sig00000178),
    .I4(sig000001da),
    .I5(sig000001db),
    .O(sig00000857)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk00000620 (
    .I0(sig00000176),
    .I1(sig00000177),
    .I2(sig00000178),
    .I3(sig00000179),
    .I4(sig000001da),
    .I5(sig000001db),
    .O(sig00000858)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk00000621 (
    .I0(sig00000177),
    .I1(sig00000178),
    .I2(sig00000179),
    .I3(sig0000017a),
    .I4(sig000001da),
    .I5(sig000001db),
    .O(sig00000859)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk00000622 (
    .I0(sig00000178),
    .I1(sig00000179),
    .I2(sig0000017a),
    .I3(sig0000017a),
    .I4(sig000001da),
    .I5(sig000001db),
    .O(sig0000085a)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk00000623 (
    .I0(sig00000179),
    .I1(sig0000017a),
    .I2(sig0000017a),
    .I3(sig0000017a),
    .I4(sig000001da),
    .I5(sig000001db),
    .O(sig0000085b)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk00000624 (
    .I0(sig0000017a),
    .I1(sig0000017a),
    .I2(sig0000017a),
    .I3(sig0000017a),
    .I4(sig000001da),
    .I5(sig000001db),
    .O(sig0000085c)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000625 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000842),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(NLW_blk00000625_Q_UNCONNECTED)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000626 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000843),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(NLW_blk00000626_Q_UNCONNECTED)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000627 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000844),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(NLW_blk00000627_Q_UNCONNECTED)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000628 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000845),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(NLW_blk00000628_Q_UNCONNECTED)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000629 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000846),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(NLW_blk00000629_Q_UNCONNECTED)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000062a (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000847),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(NLW_blk0000062a_Q_UNCONNECTED)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000062b (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000848),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(NLW_blk0000062b_Q_UNCONNECTED)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000062c (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000849),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(NLW_blk0000062c_Q_UNCONNECTED)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000062d (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000084a),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig0000009e)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000062e (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000084b),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig0000009f)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000062f (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000084c),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000000a0)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000630 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000084d),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000000a1)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000631 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000084e),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000000a2)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000632 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000084f),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000000a3)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000633 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000850),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000000a4)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000634 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000851),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000000a5)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000635 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000852),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000000a6)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000636 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000853),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000000a7)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000637 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000854),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000000a8)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000638 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000855),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000000a9)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000639 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000856),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000000aa)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000063a (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000857),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000000ab)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000063b (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000858),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000000ac)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000063c (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000859),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000000ad)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000063d (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000085a),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(NLW_blk0000063d_Q_UNCONNECTED)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000063e (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000085b),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(NLW_blk0000063e_Q_UNCONNECTED)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000063f (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000085c),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(NLW_blk0000063f_Q_UNCONNECTED)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000645 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig0000085d)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000646 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(sig00000344),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig0000085e)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000647 (
    .A0(sig00000344),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(sig00000344),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000891),
    .Q(sig0000085f)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000648 (
    .A0(sig00000344),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(sig00000344),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000892),
    .Q(sig00000860)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000649 (
    .A0(sig00000344),
    .A1(sig00000344),
    .A2(sig00000344),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000890),
    .Q(sig00000861)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000064a (
    .A0(sig00000344),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000000be),
    .Q(sig00000863)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000064b (
    .A0(sig00000344),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000000bf),
    .Q(sig00000864)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000064c (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(sig00000344),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000000c0),
    .Q(sig00000865)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000064d (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(sig00000344),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000000c1),
    .Q(sig00000866)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000064e (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000085d),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(NLW_blk0000064e_Q_UNCONNECTED)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000064f (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000085e),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(NLW_blk0000064f_Q_UNCONNECTED)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000650 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000085f),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig0000088c)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000651 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000860),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig0000088d)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000652 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000861),
    .R(NLW_blk00000652_R_UNCONNECTED),
    .Q(sig00000862)
  );
  FDR #(
    .INIT ( 1'b0 ))
  blk00000653 (
    .C(aclk),
    .D(sig00000862),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000070)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000654 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000863),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000891)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000655 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000864),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000892)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000656 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000865),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000893)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000657 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000866),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000894)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000658 (
    .C(aclk),
    .D(sig00000867),
    .Q(sig0000088f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000065d (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000090a),
    .Q(sig0000097f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000065e (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000090b),
    .Q(sig00000980)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000065f (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000090c),
    .Q(sig00000981)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000660 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000090d),
    .Q(sig00000982)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000661 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000090e),
    .Q(sig00000983)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000662 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000090f),
    .Q(sig00000984)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000663 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000910),
    .Q(sig00000985)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000664 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000911),
    .Q(sig00000986)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000665 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000912),
    .Q(sig00000987)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000666 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000913),
    .Q(sig00000988)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000667 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000914),
    .Q(sig00000989)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000668 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000915),
    .Q(sig0000098a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000669 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000916),
    .Q(sig0000098b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000066a (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000917),
    .Q(sig0000098c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000066b (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000918),
    .Q(sig0000098d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000066c (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000919),
    .Q(sig0000098e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000066d (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000091a),
    .Q(sig0000098f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000066e (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000008d8),
    .Q(sig00000990)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000066f (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000008d9),
    .Q(sig00000991)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000670 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000008da),
    .Q(sig00000992)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000671 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000008db),
    .Q(sig00000993)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000672 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000008dc),
    .Q(sig00000994)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000673 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000008dd),
    .Q(sig00000995)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000674 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000008de),
    .Q(sig00000996)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000675 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000008df),
    .Q(sig00000997)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000676 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000008e0),
    .Q(sig00000998)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000677 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000008e1),
    .Q(sig00000999)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000678 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000008e2),
    .Q(sig0000099a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000679 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000008e3),
    .Q(sig0000099b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000067a (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000008e4),
    .Q(sig0000099c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000067b (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000008e5),
    .Q(sig0000099d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000067c (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000008e6),
    .Q(sig0000099e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000067d (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000008e7),
    .Q(sig0000099f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000067e (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000008e8),
    .Q(sig000009a0)
  );
  MUXCY   blk0000067f (
    .CI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .DI(sig000009a1),
    .S(sig000008c7),
    .O(sig000008b7)
  );
  MUXCY   blk00000680 (
    .CI(sig000008b7),
    .DI(sig000009a2),
    .S(sig000008c9),
    .O(sig000008b8)
  );
  MUXCY   blk00000681 (
    .CI(sig000008b8),
    .DI(sig000009a3),
    .S(sig000008ca),
    .O(sig000008b9)
  );
  MUXCY   blk00000682 (
    .CI(sig000008b9),
    .DI(sig000009a4),
    .S(sig000008cb),
    .O(sig000008ba)
  );
  MUXCY   blk00000683 (
    .CI(sig000008ba),
    .DI(sig000009a5),
    .S(sig000008cc),
    .O(sig000008bb)
  );
  MUXCY   blk00000684 (
    .CI(sig000008bb),
    .DI(sig000009a6),
    .S(sig000008cd),
    .O(sig000008bc)
  );
  MUXCY   blk00000685 (
    .CI(sig000008bc),
    .DI(sig000009a7),
    .S(sig000008ce),
    .O(sig000008bd)
  );
  MUXCY   blk00000686 (
    .CI(sig000008bd),
    .DI(sig000009a8),
    .S(sig000008cf),
    .O(sig000008be)
  );
  MUXCY   blk00000687 (
    .CI(sig000008be),
    .DI(sig000009a9),
    .S(sig000008d0),
    .O(sig000008bf)
  );
  MUXCY   blk00000688 (
    .CI(sig000008bf),
    .DI(sig000009aa),
    .S(sig000008d1),
    .O(sig000008c0)
  );
  MUXCY   blk00000689 (
    .CI(sig000008c0),
    .DI(sig000009ab),
    .S(sig000008d2),
    .O(sig000008c1)
  );
  MUXCY   blk0000068a (
    .CI(sig000008c1),
    .DI(sig000009ac),
    .S(sig000008d3),
    .O(sig000008c2)
  );
  MUXCY   blk0000068b (
    .CI(sig000008c2),
    .DI(sig000009ad),
    .S(sig000008d4),
    .O(sig000008c3)
  );
  MUXCY   blk0000068c (
    .CI(sig000008c3),
    .DI(sig000009ae),
    .S(sig000008d5),
    .O(sig000008c4)
  );
  MUXCY   blk0000068d (
    .CI(sig000008c4),
    .DI(sig000009af),
    .S(sig000008d6),
    .O(sig000008c5)
  );
  MUXCY   blk0000068e (
    .CI(sig000008c5),
    .DI(sig000009b0),
    .S(sig000008d7),
    .O(sig000008c6)
  );
  XORCY   blk0000068f (
    .CI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .LI(sig000008c7),
    .O(sig000008d8)
  );
  XORCY   blk00000690 (
    .CI(sig000008b7),
    .LI(sig000008c9),
    .O(sig000008d9)
  );
  XORCY   blk00000691 (
    .CI(sig000008b8),
    .LI(sig000008ca),
    .O(sig000008da)
  );
  XORCY   blk00000692 (
    .CI(sig000008b9),
    .LI(sig000008cb),
    .O(sig000008db)
  );
  XORCY   blk00000693 (
    .CI(sig000008ba),
    .LI(sig000008cc),
    .O(sig000008dc)
  );
  XORCY   blk00000694 (
    .CI(sig000008bb),
    .LI(sig000008cd),
    .O(sig000008dd)
  );
  XORCY   blk00000695 (
    .CI(sig000008bc),
    .LI(sig000008ce),
    .O(sig000008de)
  );
  XORCY   blk00000696 (
    .CI(sig000008bd),
    .LI(sig000008cf),
    .O(sig000008df)
  );
  XORCY   blk00000697 (
    .CI(sig000008be),
    .LI(sig000008d0),
    .O(sig000008e0)
  );
  XORCY   blk00000698 (
    .CI(sig000008bf),
    .LI(sig000008d1),
    .O(sig000008e1)
  );
  XORCY   blk00000699 (
    .CI(sig000008c0),
    .LI(sig000008d2),
    .O(sig000008e2)
  );
  XORCY   blk0000069a (
    .CI(sig000008c1),
    .LI(sig000008d3),
    .O(sig000008e3)
  );
  XORCY   blk0000069b (
    .CI(sig000008c2),
    .LI(sig000008d4),
    .O(sig000008e4)
  );
  XORCY   blk0000069c (
    .CI(sig000008c3),
    .LI(sig000008d5),
    .O(sig000008e5)
  );
  XORCY   blk0000069d (
    .CI(sig000008c4),
    .LI(sig000008d6),
    .O(sig000008e6)
  );
  XORCY   blk0000069e (
    .CI(sig000008c5),
    .LI(sig000008d7),
    .O(sig000008e7)
  );
  XORCY   blk0000069f (
    .CI(sig000008c6),
    .LI(sig000008c8),
    .O(sig000008e8)
  );
  MUXCY   blk000006a0 (
    .CI(sig00000344),
    .DI(sig000009a1),
    .S(sig000008f9),
    .O(sig000008e9)
  );
  MUXCY   blk000006a1 (
    .CI(sig000008e9),
    .DI(sig000009a2),
    .S(sig000008fb),
    .O(sig000008ea)
  );
  MUXCY   blk000006a2 (
    .CI(sig000008ea),
    .DI(sig000009a3),
    .S(sig000008fc),
    .O(sig000008eb)
  );
  MUXCY   blk000006a3 (
    .CI(sig000008eb),
    .DI(sig000009a4),
    .S(sig000008fd),
    .O(sig000008ec)
  );
  MUXCY   blk000006a4 (
    .CI(sig000008ec),
    .DI(sig000009a5),
    .S(sig000008fe),
    .O(sig000008ed)
  );
  MUXCY   blk000006a5 (
    .CI(sig000008ed),
    .DI(sig000009a6),
    .S(sig000008ff),
    .O(sig000008ee)
  );
  MUXCY   blk000006a6 (
    .CI(sig000008ee),
    .DI(sig000009a7),
    .S(sig00000900),
    .O(sig000008ef)
  );
  MUXCY   blk000006a7 (
    .CI(sig000008ef),
    .DI(sig000009a8),
    .S(sig00000901),
    .O(sig000008f0)
  );
  MUXCY   blk000006a8 (
    .CI(sig000008f0),
    .DI(sig000009a9),
    .S(sig00000902),
    .O(sig000008f1)
  );
  MUXCY   blk000006a9 (
    .CI(sig000008f1),
    .DI(sig000009aa),
    .S(sig00000903),
    .O(sig000008f2)
  );
  MUXCY   blk000006aa (
    .CI(sig000008f2),
    .DI(sig000009ab),
    .S(sig00000904),
    .O(sig000008f3)
  );
  MUXCY   blk000006ab (
    .CI(sig000008f3),
    .DI(sig000009ac),
    .S(sig00000905),
    .O(sig000008f4)
  );
  MUXCY   blk000006ac (
    .CI(sig000008f4),
    .DI(sig000009ad),
    .S(sig00000906),
    .O(sig000008f5)
  );
  MUXCY   blk000006ad (
    .CI(sig000008f5),
    .DI(sig000009ae),
    .S(sig00000907),
    .O(sig000008f6)
  );
  MUXCY   blk000006ae (
    .CI(sig000008f6),
    .DI(sig000009af),
    .S(sig00000908),
    .O(sig000008f7)
  );
  MUXCY   blk000006af (
    .CI(sig000008f7),
    .DI(sig000009b0),
    .S(sig00000909),
    .O(sig000008f8)
  );
  XORCY   blk000006b0 (
    .CI(sig00000344),
    .LI(sig000008f9),
    .O(sig0000090a)
  );
  XORCY   blk000006b1 (
    .CI(sig000008e9),
    .LI(sig000008fb),
    .O(sig0000090b)
  );
  XORCY   blk000006b2 (
    .CI(sig000008ea),
    .LI(sig000008fc),
    .O(sig0000090c)
  );
  XORCY   blk000006b3 (
    .CI(sig000008eb),
    .LI(sig000008fd),
    .O(sig0000090d)
  );
  XORCY   blk000006b4 (
    .CI(sig000008ec),
    .LI(sig000008fe),
    .O(sig0000090e)
  );
  XORCY   blk000006b5 (
    .CI(sig000008ed),
    .LI(sig000008ff),
    .O(sig0000090f)
  );
  XORCY   blk000006b6 (
    .CI(sig000008ee),
    .LI(sig00000900),
    .O(sig00000910)
  );
  XORCY   blk000006b7 (
    .CI(sig000008ef),
    .LI(sig00000901),
    .O(sig00000911)
  );
  XORCY   blk000006b8 (
    .CI(sig000008f0),
    .LI(sig00000902),
    .O(sig00000912)
  );
  XORCY   blk000006b9 (
    .CI(sig000008f1),
    .LI(sig00000903),
    .O(sig00000913)
  );
  XORCY   blk000006ba (
    .CI(sig000008f2),
    .LI(sig00000904),
    .O(sig00000914)
  );
  XORCY   blk000006bb (
    .CI(sig000008f3),
    .LI(sig00000905),
    .O(sig00000915)
  );
  XORCY   blk000006bc (
    .CI(sig000008f4),
    .LI(sig00000906),
    .O(sig00000916)
  );
  XORCY   blk000006bd (
    .CI(sig000008f5),
    .LI(sig00000907),
    .O(sig00000917)
  );
  XORCY   blk000006be (
    .CI(sig000008f6),
    .LI(sig00000908),
    .O(sig00000918)
  );
  XORCY   blk000006bf (
    .CI(sig000008f7),
    .LI(sig00000909),
    .O(sig00000919)
  );
  XORCY   blk000006c0 (
    .CI(sig000008f8),
    .LI(sig000008fa),
    .O(sig0000091a)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000006c1 (
    .I0(sig00000990),
    .I1(sig0000096e),
    .I2(sig000009b1),
    .O(sig0000091b)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000006c2 (
    .I0(sig00000991),
    .I1(sig0000096f),
    .I2(sig000009b1),
    .O(sig0000091c)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000006c3 (
    .I0(sig00000992),
    .I1(sig00000970),
    .I2(sig000009b1),
    .O(sig0000091d)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000006c4 (
    .I0(sig00000993),
    .I1(sig00000971),
    .I2(sig000009b1),
    .O(sig0000091e)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000006c5 (
    .I0(sig00000994),
    .I1(sig00000972),
    .I2(sig000009b1),
    .O(sig0000091f)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000006c6 (
    .I0(sig00000995),
    .I1(sig00000973),
    .I2(sig000009b1),
    .O(sig00000920)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000006c7 (
    .I0(sig00000996),
    .I1(sig00000974),
    .I2(sig000009b1),
    .O(sig00000921)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000006c8 (
    .I0(sig00000997),
    .I1(sig00000975),
    .I2(sig000009b1),
    .O(sig00000922)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000006c9 (
    .I0(sig00000998),
    .I1(sig00000976),
    .I2(sig000009b1),
    .O(sig00000923)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000006ca (
    .I0(sig00000999),
    .I1(sig00000977),
    .I2(sig000009b1),
    .O(sig00000924)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000006cb (
    .I0(sig0000099a),
    .I1(sig00000978),
    .I2(sig000009b1),
    .O(sig00000925)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000006cc (
    .I0(sig0000099b),
    .I1(sig00000979),
    .I2(sig000009b1),
    .O(sig00000926)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000006cd (
    .I0(sig0000099c),
    .I1(sig0000097a),
    .I2(sig000009b1),
    .O(sig00000927)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000006ce (
    .I0(sig0000099d),
    .I1(sig0000097b),
    .I2(sig000009b1),
    .O(sig00000928)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000006cf (
    .I0(sig0000099e),
    .I1(sig0000097c),
    .I2(sig000009b1),
    .O(sig00000929)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000006d0 (
    .I0(sig0000099f),
    .I1(sig0000097d),
    .I2(sig000009b1),
    .O(sig0000092a)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000006d1 (
    .I0(sig000009a0),
    .I1(sig0000097e),
    .I2(sig000009b1),
    .O(sig0000092b)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000006d2 (
    .I0(sig0000096e),
    .I1(sig00000990),
    .I2(sig000009b1),
    .O(sig0000092c)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000006d3 (
    .I0(sig0000096f),
    .I1(sig00000991),
    .I2(sig000009b1),
    .O(sig0000092d)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000006d4 (
    .I0(sig00000970),
    .I1(sig00000992),
    .I2(sig000009b1),
    .O(sig0000092e)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000006d5 (
    .I0(sig00000971),
    .I1(sig00000993),
    .I2(sig000009b1),
    .O(sig0000092f)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000006d6 (
    .I0(sig00000972),
    .I1(sig00000994),
    .I2(sig000009b1),
    .O(sig00000930)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000006d7 (
    .I0(sig00000973),
    .I1(sig00000995),
    .I2(sig000009b1),
    .O(sig00000931)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000006d8 (
    .I0(sig00000974),
    .I1(sig00000996),
    .I2(sig000009b1),
    .O(sig00000932)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000006d9 (
    .I0(sig00000975),
    .I1(sig00000997),
    .I2(sig000009b1),
    .O(sig00000933)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000006da (
    .I0(sig00000976),
    .I1(sig00000998),
    .I2(sig000009b1),
    .O(sig00000934)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000006db (
    .I0(sig00000977),
    .I1(sig00000999),
    .I2(sig000009b1),
    .O(sig00000935)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000006dc (
    .I0(sig00000978),
    .I1(sig0000099a),
    .I2(sig000009b1),
    .O(sig00000936)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000006dd (
    .I0(sig00000979),
    .I1(sig0000099b),
    .I2(sig000009b1),
    .O(sig00000937)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000006de (
    .I0(sig0000097a),
    .I1(sig0000099c),
    .I2(sig000009b1),
    .O(sig00000938)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000006df (
    .I0(sig0000097b),
    .I1(sig0000099d),
    .I2(sig000009b1),
    .O(sig00000939)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000006e0 (
    .I0(sig0000097c),
    .I1(sig0000099e),
    .I2(sig000009b1),
    .O(sig0000093a)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000006e1 (
    .I0(sig0000097d),
    .I1(sig0000099f),
    .I2(sig000009b1),
    .O(sig0000093b)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000006e2 (
    .I0(sig0000097e),
    .I1(sig000009a0),
    .I2(sig000009b1),
    .O(sig0000093c)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000006e3 (
    .I0(sig000000ae),
    .I1(sig000009b4),
    .I2(sig000000c1),
    .O(sig0000093d)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000006e4 (
    .I0(sig000000af),
    .I1(sig000009b5),
    .I2(sig000000c1),
    .O(sig0000093e)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000006e5 (
    .I0(sig000000b0),
    .I1(sig000009b6),
    .I2(sig000000c1),
    .O(sig0000093f)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000006e6 (
    .I0(sig000000b1),
    .I1(sig000009b7),
    .I2(sig000000c1),
    .O(sig00000940)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000006e7 (
    .I0(sig000000b2),
    .I1(sig000009b8),
    .I2(sig000000c1),
    .O(sig00000941)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000006e8 (
    .I0(sig000000b3),
    .I1(sig000009b9),
    .I2(sig000000c1),
    .O(sig00000942)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000006e9 (
    .I0(sig000000b4),
    .I1(sig000009ba),
    .I2(sig000000c1),
    .O(sig00000943)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000006ea (
    .I0(sig000000b5),
    .I1(sig000009bb),
    .I2(sig000000c1),
    .O(sig00000944)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000006eb (
    .I0(sig000000b6),
    .I1(sig000009bc),
    .I2(sig000000c1),
    .O(sig00000945)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000006ec (
    .I0(sig000000b7),
    .I1(sig000009bd),
    .I2(sig000000c1),
    .O(sig00000946)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000006ed (
    .I0(sig000000b8),
    .I1(sig000009be),
    .I2(sig000000c1),
    .O(sig00000947)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000006ee (
    .I0(sig000000b9),
    .I1(sig000009bf),
    .I2(sig000000c1),
    .O(sig00000948)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000006ef (
    .I0(sig000000ba),
    .I1(sig000009c0),
    .I2(sig000000c1),
    .O(sig00000949)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000006f0 (
    .I0(sig000000bb),
    .I1(sig000009c1),
    .I2(sig000000c1),
    .O(sig0000094a)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000006f1 (
    .I0(sig000000bc),
    .I1(sig000009c2),
    .I2(sig000000c1),
    .O(sig0000094b)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000006f2 (
    .I0(sig000000bd),
    .I1(sig000009c3),
    .I2(sig000000c1),
    .O(sig0000094c)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000006f3 (
    .I0(sig000009b4),
    .I1(sig000000ae),
    .I2(sig000000c1),
    .O(sig0000094d)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000006f4 (
    .I0(sig000009b5),
    .I1(sig000000af),
    .I2(sig000000c1),
    .O(sig0000094e)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000006f5 (
    .I0(sig000009b6),
    .I1(sig000000b0),
    .I2(sig000000c1),
    .O(sig0000094f)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000006f6 (
    .I0(sig000009b7),
    .I1(sig000000b1),
    .I2(sig000000c1),
    .O(sig00000950)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000006f7 (
    .I0(sig000009b8),
    .I1(sig000000b2),
    .I2(sig000000c1),
    .O(sig00000951)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000006f8 (
    .I0(sig000009b9),
    .I1(sig000000b3),
    .I2(sig000000c1),
    .O(sig00000952)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000006f9 (
    .I0(sig000009ba),
    .I1(sig000000b4),
    .I2(sig000000c1),
    .O(sig00000953)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000006fa (
    .I0(sig000009bb),
    .I1(sig000000b5),
    .I2(sig000000c1),
    .O(sig00000954)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000006fb (
    .I0(sig000009bc),
    .I1(sig000000b6),
    .I2(sig000000c1),
    .O(sig00000955)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000006fc (
    .I0(sig000009bd),
    .I1(sig000000b7),
    .I2(sig000000c1),
    .O(sig00000956)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000006fd (
    .I0(sig000009be),
    .I1(sig000000b8),
    .I2(sig000000c1),
    .O(sig00000957)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000006fe (
    .I0(sig000009bf),
    .I1(sig000000b9),
    .I2(sig000000c1),
    .O(sig00000958)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000006ff (
    .I0(sig000009c0),
    .I1(sig000000ba),
    .I2(sig000000c1),
    .O(sig00000959)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000700 (
    .I0(sig000009c1),
    .I1(sig000000bb),
    .I2(sig000000c1),
    .O(sig0000095a)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000701 (
    .I0(sig000009c2),
    .I1(sig000000bc),
    .I2(sig000000c1),
    .O(sig0000095b)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000702 (
    .I0(sig000009c3),
    .I1(sig000000bd),
    .I2(sig000000c1),
    .O(sig0000095c)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000703 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000091b),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig0000095d)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000704 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000091c),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig0000095e)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000705 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000091d),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig0000095f)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000706 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000091e),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000960)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000707 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000091f),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000961)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000708 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000920),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000962)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000709 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000921),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000963)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000070a (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000922),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000964)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000070b (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000923),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000965)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000070c (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000924),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000966)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000070d (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000925),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000967)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000070e (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000926),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000968)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000070f (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000927),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000969)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000710 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000928),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig0000096a)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000711 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000929),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig0000096b)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000712 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000092a),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig0000096c)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000713 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000092b),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig0000096d)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000714 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000092c),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000895)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000715 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000092d),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000896)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000716 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000092e),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000897)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000717 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000092f),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000898)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000718 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000930),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000899)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000719 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000931),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig0000089a)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000071a (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000932),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig0000089b)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000071b (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000933),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig0000089c)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000071c (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000934),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig0000089d)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000071d (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000935),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig0000089e)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000071e (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000936),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig0000089f)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000071f (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000937),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000008a0)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000720 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000938),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000008a1)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000721 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000939),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000008a2)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000722 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000093a),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000008a3)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000723 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000093b),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000008a4)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000724 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000093c),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000008a5)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000725 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000009b3),
    .Q(sig000009b2)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000726 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000093d),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000009d4)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000727 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000093e),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000009d5)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000728 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000093f),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000009d6)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000729 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000940),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000009d7)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000072a (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000941),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000009d8)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000072b (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000942),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000009d9)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000072c (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000943),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000009da)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000072d (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000944),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000009db)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000072e (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000945),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000009dc)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000072f (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000946),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000009dd)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000730 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000947),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000009de)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000731 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000948),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000009df)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000732 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000949),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000009e0)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000733 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000094a),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000009e1)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000734 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000094b),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000009e2)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000735 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000094c),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000009e3)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000736 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000094d),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000009c4)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000737 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000094e),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000009c5)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000738 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000094f),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000009c6)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000739 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000950),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000009c7)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000073a (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000951),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000009c8)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000073b (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000952),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000009c9)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000073c (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000953),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000009ca)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000073d (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000954),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000009cb)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000073e (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000955),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000009cc)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000073f (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000956),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000009cd)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000740 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000957),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000009ce)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000741 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000958),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000009cf)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000742 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000959),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000009d0)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000743 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000095a),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000009d1)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000744 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000095b),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000009d2)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000745 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000095c),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000009d3)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000746 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000000c1),
    .Q(sig000009b3)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000747 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000009e3),
    .Q(sig000009e4)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000748 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000009e2),
    .Q(sig000009e5)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000749 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000009e1),
    .Q(sig000009e6)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000074a (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000009e0),
    .Q(sig000009e7)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000074b (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000009df),
    .Q(sig000009e8)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000074c (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000009de),
    .Q(sig000009e9)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000074d (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000009dd),
    .Q(sig000009ea)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000074e (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000009dc),
    .Q(sig000009eb)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000074f (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000009db),
    .Q(sig000009ec)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000750 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000009da),
    .Q(sig000009ed)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000751 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000009d9),
    .Q(sig000009ee)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000752 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000009d8),
    .Q(sig000009ef)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000753 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000009d7),
    .Q(sig000009f0)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000754 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000009d6),
    .Q(sig000009f1)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000755 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000009d5),
    .Q(sig000009f2)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000756 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000009d4),
    .Q(sig000009f3)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000757 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000009e4),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000009b0)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000758 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000009e5),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000009af)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000759 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000009e6),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000009ae)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000075a (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000009e7),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000009ad)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000075b (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000009e8),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000009ac)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000075c (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000009e9),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000009ab)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000075d (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000009ea),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000009aa)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000075e (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000009eb),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000009a9)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000075f (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000009ec),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000009a8)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000760 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000009ed),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000009a7)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000761 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000009ee),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000009a6)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000762 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000009ef),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000009a5)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000763 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000009f0),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000009a4)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000764 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000009f1),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000009a3)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000765 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000009f2),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000009a2)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000766 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000009f3),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000009a1)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000767 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000000ad),
    .Q(sig000009f4)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000768 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000000ac),
    .Q(sig000009f5)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000769 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000000ab),
    .Q(sig000009f6)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000076a (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000000aa),
    .Q(sig000009f7)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000076b (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000000a9),
    .Q(sig000009f8)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000076c (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000000a8),
    .Q(sig000009f9)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000076d (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000000a7),
    .Q(sig000009fa)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000076e (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000000a6),
    .Q(sig000009fb)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000076f (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000000a5),
    .Q(sig000009fc)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000770 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000000a4),
    .Q(sig000009fd)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000771 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000000a3),
    .Q(sig000009fe)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000772 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000000a2),
    .Q(sig000009ff)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000773 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000000a1),
    .Q(sig00000a00)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000774 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000000a0),
    .Q(sig00000a01)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000775 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig0000009f),
    .Q(sig00000a02)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000776 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig0000009e),
    .Q(sig00000a03)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000777 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000009f4),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000009c3)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000778 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000009f5),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000009c2)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000779 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000009f6),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000009c1)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000077a (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000009f7),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000009c0)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000077b (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000009f8),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000009bf)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000077c (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000009f9),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000009be)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000077d (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000009fa),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000009bd)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000077e (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000009fb),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000009bc)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000077f (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000009fc),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000009bb)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000780 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000009fd),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000009ba)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000781 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000009fe),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000009b9)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000782 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig000009ff),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000009b8)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000783 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000a00),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000009b7)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000784 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000a01),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000009b6)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000785 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000a02),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000009b5)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000786 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000a03),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000009b4)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000787 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig0000096d),
    .Q(sig00000a04)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000788 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig0000096c),
    .Q(sig00000a05)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000789 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig0000096b),
    .Q(sig00000a06)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000078a (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig0000096a),
    .Q(sig00000a07)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000078b (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000969),
    .Q(sig00000a08)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000078c (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000968),
    .Q(sig00000a09)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000078d (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000967),
    .Q(sig00000a0a)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000078e (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000966),
    .Q(sig00000a0b)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000078f (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000965),
    .Q(sig00000a0c)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000790 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000964),
    .Q(sig00000a0d)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000791 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000963),
    .Q(sig00000a0e)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000792 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000962),
    .Q(sig00000a0f)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000793 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000961),
    .Q(sig00000a10)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000794 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000960),
    .Q(sig00000a11)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000795 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig0000095f),
    .Q(sig00000a12)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000796 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig0000095e),
    .Q(sig00000a13)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000797 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig0000095d),
    .Q(sig00000a14)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000798 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000a04),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000008b6)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000799 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000a05),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000008b5)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000079a (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000a06),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000008b4)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000079b (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000a07),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000008b3)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000079c (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000a08),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000008b2)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000079d (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000a09),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000008b1)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000079e (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000a0a),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000008b0)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000079f (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000a0b),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000008af)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000007a0 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000a0c),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000008ae)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000007a1 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000a0d),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000008ad)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000007a2 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000a0e),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000008ac)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000007a3 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000a0f),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000008ab)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000007a4 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000a10),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000008aa)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000007a5 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000a11),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000008a9)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000007a6 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000a12),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000008a8)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000007a7 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000a13),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000008a7)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000007a8 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000a14),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig000008a6)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000007a9 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig0000098f),
    .Q(sig00000a15)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000007aa (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig0000098e),
    .Q(sig00000a16)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000007ab (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig0000098d),
    .Q(sig00000a17)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000007ac (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig0000098c),
    .Q(sig00000a18)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000007ad (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig0000098b),
    .Q(sig00000a19)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000007ae (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig0000098a),
    .Q(sig00000a1a)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000007af (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000989),
    .Q(sig00000a1b)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000007b0 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000988),
    .Q(sig00000a1c)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000007b1 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000987),
    .Q(sig00000a1d)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000007b2 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000986),
    .Q(sig00000a1e)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000007b3 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000985),
    .Q(sig00000a1f)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000007b4 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000984),
    .Q(sig00000a20)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000007b5 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000983),
    .Q(sig00000a21)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000007b6 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000982),
    .Q(sig00000a22)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000007b7 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000981),
    .Q(sig00000a23)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000007b8 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000980),
    .Q(sig00000a24)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000007b9 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig0000097f),
    .Q(sig00000a25)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000007ba (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000a15),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig0000097e)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000007bb (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000a16),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig0000097d)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000007bc (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000a17),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig0000097c)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000007bd (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000a18),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig0000097b)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000007be (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000a19),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig0000097a)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000007bf (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000a1a),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000979)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000007c0 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000a1b),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000978)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000007c1 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000a1c),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000977)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000007c2 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000a1d),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000976)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000007c3 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000a1e),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000975)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000007c4 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000a1f),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000974)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000007c5 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000a20),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000973)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000007c6 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000a21),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000972)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000007c7 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000a22),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000971)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000007c8 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000a23),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000970)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000007c9 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000a24),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig0000096f)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000007ca (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000a25),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig0000096e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000007d0 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000a7e),
    .Q(sig00000b8d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000007d1 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000a7f),
    .Q(sig00000b8e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000007d2 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000a80),
    .Q(sig00000b8f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000007d3 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000a81),
    .Q(sig00000b90)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000007d4 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000a82),
    .Q(sig00000b91)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000007d5 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000a83),
    .Q(sig00000b92)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000007d6 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000a84),
    .Q(sig00000b93)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000007d7 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000a85),
    .Q(sig00000b94)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000007d8 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000a86),
    .Q(sig00000b95)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000007d9 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000a87),
    .Q(sig00000b96)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000007da (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000a88),
    .Q(sig00000b97)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000007db (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000a89),
    .Q(sig00000b98)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000007dc (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000a8a),
    .Q(sig00000b99)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000007dd (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000a8b),
    .Q(sig00000b9a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000007de (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000a8c),
    .Q(sig00000b9b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000007df (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000a8d),
    .Q(sig00000b9c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000007e0 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000a8e),
    .Q(sig00000b9d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000007e1 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000a8f),
    .Q(sig00000b9e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000007e2 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000a49),
    .Q(sig00000b9f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000007e3 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000a4a),
    .Q(sig00000ba0)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000007e4 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000a4b),
    .Q(sig00000ba1)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000007e5 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000a4c),
    .Q(sig00000ba2)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000007e6 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000a4d),
    .Q(sig00000ba3)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000007e7 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000a4e),
    .Q(sig00000ba4)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000007e8 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000a4f),
    .Q(sig00000ba5)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000007e9 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000a50),
    .Q(sig00000ba6)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000007ea (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000a51),
    .Q(sig00000ba7)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000007eb (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000a52),
    .Q(sig00000ba8)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000007ec (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000a53),
    .Q(sig00000ba9)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000007ed (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000a54),
    .Q(sig00000baa)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000007ee (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000a55),
    .Q(sig00000bab)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000007ef (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000a56),
    .Q(sig00000bac)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000007f0 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000a57),
    .Q(sig00000bad)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000007f1 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000a58),
    .Q(sig00000bae)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000007f2 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000a59),
    .Q(sig00000baf)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000007f3 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000a5a),
    .Q(sig00000bb0)
  );
  MUXCY   blk000007f4 (
    .CI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .DI(sig00000be7),
    .S(sig00000a37),
    .O(sig00000a26)
  );
  MUXCY   blk000007f5 (
    .CI(sig00000a26),
    .DI(sig00000be8),
    .S(sig00000a39),
    .O(sig00000a27)
  );
  MUXCY   blk000007f6 (
    .CI(sig00000a27),
    .DI(sig00000be9),
    .S(sig00000a3a),
    .O(sig00000a28)
  );
  MUXCY   blk000007f7 (
    .CI(sig00000a28),
    .DI(sig00000bea),
    .S(sig00000a3b),
    .O(sig00000a29)
  );
  MUXCY   blk000007f8 (
    .CI(sig00000a29),
    .DI(sig00000beb),
    .S(sig00000a3c),
    .O(sig00000a2a)
  );
  MUXCY   blk000007f9 (
    .CI(sig00000a2a),
    .DI(sig00000bec),
    .S(sig00000a3d),
    .O(sig00000a2b)
  );
  MUXCY   blk000007fa (
    .CI(sig00000a2b),
    .DI(sig00000bed),
    .S(sig00000a3e),
    .O(sig00000a2c)
  );
  MUXCY   blk000007fb (
    .CI(sig00000a2c),
    .DI(sig00000bee),
    .S(sig00000a3f),
    .O(sig00000a2d)
  );
  MUXCY   blk000007fc (
    .CI(sig00000a2d),
    .DI(sig00000bef),
    .S(sig00000a40),
    .O(sig00000a2e)
  );
  MUXCY   blk000007fd (
    .CI(sig00000a2e),
    .DI(sig00000bf0),
    .S(sig00000a41),
    .O(sig00000a2f)
  );
  MUXCY   blk000007fe (
    .CI(sig00000a2f),
    .DI(sig00000bf1),
    .S(sig00000a42),
    .O(sig00000a30)
  );
  MUXCY   blk000007ff (
    .CI(sig00000a30),
    .DI(sig00000bf2),
    .S(sig00000a43),
    .O(sig00000a31)
  );
  MUXCY   blk00000800 (
    .CI(sig00000a31),
    .DI(sig00000bf3),
    .S(sig00000a44),
    .O(sig00000a32)
  );
  MUXCY   blk00000801 (
    .CI(sig00000a32),
    .DI(sig00000bf4),
    .S(sig00000a45),
    .O(sig00000a33)
  );
  MUXCY   blk00000802 (
    .CI(sig00000a33),
    .DI(sig00000bf5),
    .S(sig00000a46),
    .O(sig00000a34)
  );
  MUXCY   blk00000803 (
    .CI(sig00000a34),
    .DI(sig00000bf6),
    .S(sig00000a47),
    .O(sig00000a35)
  );
  MUXCY   blk00000804 (
    .CI(sig00000a35),
    .DI(sig00000bf7),
    .S(sig00000a48),
    .O(sig00000a36)
  );
  XORCY   blk00000805 (
    .CI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .LI(sig00000a37),
    .O(sig00000a49)
  );
  XORCY   blk00000806 (
    .CI(sig00000a26),
    .LI(sig00000a39),
    .O(sig00000a4a)
  );
  XORCY   blk00000807 (
    .CI(sig00000a27),
    .LI(sig00000a3a),
    .O(sig00000a4b)
  );
  XORCY   blk00000808 (
    .CI(sig00000a28),
    .LI(sig00000a3b),
    .O(sig00000a4c)
  );
  XORCY   blk00000809 (
    .CI(sig00000a29),
    .LI(sig00000a3c),
    .O(sig00000a4d)
  );
  XORCY   blk0000080a (
    .CI(sig00000a2a),
    .LI(sig00000a3d),
    .O(sig00000a4e)
  );
  XORCY   blk0000080b (
    .CI(sig00000a2b),
    .LI(sig00000a3e),
    .O(sig00000a4f)
  );
  XORCY   blk0000080c (
    .CI(sig00000a2c),
    .LI(sig00000a3f),
    .O(sig00000a50)
  );
  XORCY   blk0000080d (
    .CI(sig00000a2d),
    .LI(sig00000a40),
    .O(sig00000a51)
  );
  XORCY   blk0000080e (
    .CI(sig00000a2e),
    .LI(sig00000a41),
    .O(sig00000a52)
  );
  XORCY   blk0000080f (
    .CI(sig00000a2f),
    .LI(sig00000a42),
    .O(sig00000a53)
  );
  XORCY   blk00000810 (
    .CI(sig00000a30),
    .LI(sig00000a43),
    .O(sig00000a54)
  );
  XORCY   blk00000811 (
    .CI(sig00000a31),
    .LI(sig00000a44),
    .O(sig00000a55)
  );
  XORCY   blk00000812 (
    .CI(sig00000a32),
    .LI(sig00000a45),
    .O(sig00000a56)
  );
  XORCY   blk00000813 (
    .CI(sig00000a33),
    .LI(sig00000a46),
    .O(sig00000a57)
  );
  XORCY   blk00000814 (
    .CI(sig00000a34),
    .LI(sig00000a47),
    .O(sig00000a58)
  );
  XORCY   blk00000815 (
    .CI(sig00000a35),
    .LI(sig00000a48),
    .O(sig00000a59)
  );
  XORCY   blk00000816 (
    .CI(sig00000a36),
    .LI(sig00000a38),
    .O(sig00000a5a)
  );
  MUXCY   blk00000817 (
    .CI(sig00000344),
    .DI(sig00000be7),
    .S(sig00000a6c),
    .O(sig00000a5b)
  );
  MUXCY   blk00000818 (
    .CI(sig00000a5b),
    .DI(sig00000be8),
    .S(sig00000a6e),
    .O(sig00000a5c)
  );
  MUXCY   blk00000819 (
    .CI(sig00000a5c),
    .DI(sig00000be9),
    .S(sig00000a6f),
    .O(sig00000a5d)
  );
  MUXCY   blk0000081a (
    .CI(sig00000a5d),
    .DI(sig00000bea),
    .S(sig00000a70),
    .O(sig00000a5e)
  );
  MUXCY   blk0000081b (
    .CI(sig00000a5e),
    .DI(sig00000beb),
    .S(sig00000a71),
    .O(sig00000a5f)
  );
  MUXCY   blk0000081c (
    .CI(sig00000a5f),
    .DI(sig00000bec),
    .S(sig00000a72),
    .O(sig00000a60)
  );
  MUXCY   blk0000081d (
    .CI(sig00000a60),
    .DI(sig00000bed),
    .S(sig00000a73),
    .O(sig00000a61)
  );
  MUXCY   blk0000081e (
    .CI(sig00000a61),
    .DI(sig00000bee),
    .S(sig00000a74),
    .O(sig00000a62)
  );
  MUXCY   blk0000081f (
    .CI(sig00000a62),
    .DI(sig00000bef),
    .S(sig00000a75),
    .O(sig00000a63)
  );
  MUXCY   blk00000820 (
    .CI(sig00000a63),
    .DI(sig00000bf0),
    .S(sig00000a76),
    .O(sig00000a64)
  );
  MUXCY   blk00000821 (
    .CI(sig00000a64),
    .DI(sig00000bf1),
    .S(sig00000a77),
    .O(sig00000a65)
  );
  MUXCY   blk00000822 (
    .CI(sig00000a65),
    .DI(sig00000bf2),
    .S(sig00000a78),
    .O(sig00000a66)
  );
  MUXCY   blk00000823 (
    .CI(sig00000a66),
    .DI(sig00000bf3),
    .S(sig00000a79),
    .O(sig00000a67)
  );
  MUXCY   blk00000824 (
    .CI(sig00000a67),
    .DI(sig00000bf4),
    .S(sig00000a7a),
    .O(sig00000a68)
  );
  MUXCY   blk00000825 (
    .CI(sig00000a68),
    .DI(sig00000bf5),
    .S(sig00000a7b),
    .O(sig00000a69)
  );
  MUXCY   blk00000826 (
    .CI(sig00000a69),
    .DI(sig00000bf6),
    .S(sig00000a7c),
    .O(sig00000a6a)
  );
  MUXCY   blk00000827 (
    .CI(sig00000a6a),
    .DI(sig00000bf7),
    .S(sig00000a7d),
    .O(sig00000a6b)
  );
  XORCY   blk00000828 (
    .CI(sig00000344),
    .LI(sig00000a6c),
    .O(sig00000a7e)
  );
  XORCY   blk00000829 (
    .CI(sig00000a5b),
    .LI(sig00000a6e),
    .O(sig00000a7f)
  );
  XORCY   blk0000082a (
    .CI(sig00000a5c),
    .LI(sig00000a6f),
    .O(sig00000a80)
  );
  XORCY   blk0000082b (
    .CI(sig00000a5d),
    .LI(sig00000a70),
    .O(sig00000a81)
  );
  XORCY   blk0000082c (
    .CI(sig00000a5e),
    .LI(sig00000a71),
    .O(sig00000a82)
  );
  XORCY   blk0000082d (
    .CI(sig00000a5f),
    .LI(sig00000a72),
    .O(sig00000a83)
  );
  XORCY   blk0000082e (
    .CI(sig00000a60),
    .LI(sig00000a73),
    .O(sig00000a84)
  );
  XORCY   blk0000082f (
    .CI(sig00000a61),
    .LI(sig00000a74),
    .O(sig00000a85)
  );
  XORCY   blk00000830 (
    .CI(sig00000a62),
    .LI(sig00000a75),
    .O(sig00000a86)
  );
  XORCY   blk00000831 (
    .CI(sig00000a63),
    .LI(sig00000a76),
    .O(sig00000a87)
  );
  XORCY   blk00000832 (
    .CI(sig00000a64),
    .LI(sig00000a77),
    .O(sig00000a88)
  );
  XORCY   blk00000833 (
    .CI(sig00000a65),
    .LI(sig00000a78),
    .O(sig00000a89)
  );
  XORCY   blk00000834 (
    .CI(sig00000a66),
    .LI(sig00000a79),
    .O(sig00000a8a)
  );
  XORCY   blk00000835 (
    .CI(sig00000a67),
    .LI(sig00000a7a),
    .O(sig00000a8b)
  );
  XORCY   blk00000836 (
    .CI(sig00000a68),
    .LI(sig00000a7b),
    .O(sig00000a8c)
  );
  XORCY   blk00000837 (
    .CI(sig00000a69),
    .LI(sig00000a7c),
    .O(sig00000a8d)
  );
  XORCY   blk00000838 (
    .CI(sig00000a6a),
    .LI(sig00000a7d),
    .O(sig00000a8e)
  );
  XORCY   blk00000839 (
    .CI(sig00000a6b),
    .LI(sig00000a6d),
    .O(sig00000a8f)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000842 (
    .I0(sig00000b45),
    .I1(sig00000bd5),
    .I2(sig00000c20),
    .O(sig00000a90)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000843 (
    .I0(sig00000b46),
    .I1(sig00000bd6),
    .I2(sig00000c20),
    .O(sig00000a91)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000844 (
    .I0(sig00000b47),
    .I1(sig00000bd7),
    .I2(sig00000c20),
    .O(sig00000a92)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000845 (
    .I0(sig00000b48),
    .I1(sig00000bd8),
    .I2(sig00000c20),
    .O(sig00000a93)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000846 (
    .I0(sig00000b49),
    .I1(sig00000bd9),
    .I2(sig00000c20),
    .O(sig00000a94)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000847 (
    .I0(sig00000b4a),
    .I1(sig00000bda),
    .I2(sig00000c20),
    .O(sig00000a95)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000848 (
    .I0(sig00000b4b),
    .I1(sig00000bdb),
    .I2(sig00000c20),
    .O(sig00000a96)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000849 (
    .I0(sig00000b4c),
    .I1(sig00000bdc),
    .I2(sig00000c20),
    .O(sig00000a97)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk0000084a (
    .I0(sig00000b4d),
    .I1(sig00000bdd),
    .I2(sig00000c20),
    .O(sig00000a98)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk0000084b (
    .I0(sig00000b4e),
    .I1(sig00000bde),
    .I2(sig00000c20),
    .O(sig00000a99)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk0000084c (
    .I0(sig00000b4f),
    .I1(sig00000bdf),
    .I2(sig00000c20),
    .O(sig00000a9a)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk0000084d (
    .I0(sig00000b50),
    .I1(sig00000be0),
    .I2(sig00000c20),
    .O(sig00000a9b)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk0000084e (
    .I0(sig00000b51),
    .I1(sig00000be1),
    .I2(sig00000c20),
    .O(sig00000a9c)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk0000084f (
    .I0(sig00000b52),
    .I1(sig00000be2),
    .I2(sig00000c20),
    .O(sig00000a9d)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000850 (
    .I0(sig00000b53),
    .I1(sig00000be3),
    .I2(sig00000c20),
    .O(sig00000a9e)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000851 (
    .I0(sig00000b54),
    .I1(sig00000be4),
    .I2(sig00000c20),
    .O(sig00000a9f)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000852 (
    .I0(sig00000b55),
    .I1(sig00000be5),
    .I2(sig00000c20),
    .O(sig00000aa0)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000853 (
    .I0(sig00000b56),
    .I1(sig00000be6),
    .I2(sig00000c20),
    .O(sig00000aa1)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000854 (
    .I0(sig00000bd5),
    .I1(sig00000b45),
    .I2(sig00000c20),
    .O(sig00000aa2)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000855 (
    .I0(sig00000bd6),
    .I1(sig00000b46),
    .I2(sig00000c20),
    .O(sig00000aa3)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000856 (
    .I0(sig00000bd7),
    .I1(sig00000b47),
    .I2(sig00000c20),
    .O(sig00000aa4)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000857 (
    .I0(sig00000bd8),
    .I1(sig00000b48),
    .I2(sig00000c20),
    .O(sig00000aa5)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000858 (
    .I0(sig00000bd9),
    .I1(sig00000b49),
    .I2(sig00000c20),
    .O(sig00000aa6)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000859 (
    .I0(sig00000bda),
    .I1(sig00000b4a),
    .I2(sig00000c20),
    .O(sig00000aa7)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk0000085a (
    .I0(sig00000bdb),
    .I1(sig00000b4b),
    .I2(sig00000c20),
    .O(sig00000aa8)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk0000085b (
    .I0(sig00000bdc),
    .I1(sig00000b4c),
    .I2(sig00000c20),
    .O(sig00000aa9)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk0000085c (
    .I0(sig00000bdd),
    .I1(sig00000b4d),
    .I2(sig00000c20),
    .O(sig00000aaa)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk0000085d (
    .I0(sig00000bde),
    .I1(sig00000b4e),
    .I2(sig00000c20),
    .O(sig00000aab)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk0000085e (
    .I0(sig00000bdf),
    .I1(sig00000b4f),
    .I2(sig00000c20),
    .O(sig00000aac)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk0000085f (
    .I0(sig00000be0),
    .I1(sig00000b50),
    .I2(sig00000c20),
    .O(sig00000aad)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000860 (
    .I0(sig00000be1),
    .I1(sig00000b51),
    .I2(sig00000c20),
    .O(sig00000aae)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000861 (
    .I0(sig00000be2),
    .I1(sig00000b52),
    .I2(sig00000c20),
    .O(sig00000aaf)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000862 (
    .I0(sig00000be3),
    .I1(sig00000b53),
    .I2(sig00000c20),
    .O(sig00000ab0)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000863 (
    .I0(sig00000be4),
    .I1(sig00000b54),
    .I2(sig00000c20),
    .O(sig00000ab1)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000864 (
    .I0(sig00000be5),
    .I1(sig00000b55),
    .I2(sig00000c20),
    .O(sig00000ab2)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000865 (
    .I0(sig00000be6),
    .I1(sig00000b56),
    .I2(sig00000c20),
    .O(sig00000ab3)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000866 (
    .I0(sig00000b9f),
    .I1(sig00000b7b),
    .I2(sig00000c1e),
    .O(sig00000ab4)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000867 (
    .I0(sig00000ba0),
    .I1(sig00000b7c),
    .I2(sig00000c1e),
    .O(sig00000ab5)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000868 (
    .I0(sig00000ba1),
    .I1(sig00000b7d),
    .I2(sig00000c1e),
    .O(sig00000ab6)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000869 (
    .I0(sig00000ba2),
    .I1(sig00000b7e),
    .I2(sig00000c1e),
    .O(sig00000ab7)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk0000086a (
    .I0(sig00000ba3),
    .I1(sig00000b7f),
    .I2(sig00000c1e),
    .O(sig00000ab8)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk0000086b (
    .I0(sig00000ba4),
    .I1(sig00000b80),
    .I2(sig00000c1e),
    .O(sig00000ab9)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk0000086c (
    .I0(sig00000ba5),
    .I1(sig00000b81),
    .I2(sig00000c1e),
    .O(sig00000aba)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk0000086d (
    .I0(sig00000ba6),
    .I1(sig00000b82),
    .I2(sig00000c1e),
    .O(sig00000abb)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk0000086e (
    .I0(sig00000ba7),
    .I1(sig00000b83),
    .I2(sig00000c1e),
    .O(sig00000abc)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk0000086f (
    .I0(sig00000ba8),
    .I1(sig00000b84),
    .I2(sig00000c1e),
    .O(sig00000abd)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000870 (
    .I0(sig00000ba9),
    .I1(sig00000b85),
    .I2(sig00000c1e),
    .O(sig00000abe)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000871 (
    .I0(sig00000baa),
    .I1(sig00000b86),
    .I2(sig00000c1e),
    .O(sig00000abf)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000872 (
    .I0(sig00000bab),
    .I1(sig00000b87),
    .I2(sig00000c1e),
    .O(sig00000ac0)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000873 (
    .I0(sig00000bac),
    .I1(sig00000b88),
    .I2(sig00000c1e),
    .O(sig00000ac1)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000874 (
    .I0(sig00000bad),
    .I1(sig00000b89),
    .I2(sig00000c1e),
    .O(sig00000ac2)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000875 (
    .I0(sig00000bae),
    .I1(sig00000b8a),
    .I2(sig00000c1e),
    .O(sig00000ac3)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000876 (
    .I0(sig00000baf),
    .I1(sig00000b8b),
    .I2(sig00000c1e),
    .O(sig00000ac4)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000877 (
    .I0(sig00000bb0),
    .I1(sig00000b8c),
    .I2(sig00000c1e),
    .O(sig00000ac5)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000878 (
    .I0(sig00000b7b),
    .I1(sig00000b9f),
    .I2(sig00000c1e),
    .O(sig00000ac6)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000879 (
    .I0(sig00000b7c),
    .I1(sig00000ba0),
    .I2(sig00000c1e),
    .O(sig00000ac7)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk0000087a (
    .I0(sig00000b7d),
    .I1(sig00000ba1),
    .I2(sig00000c1e),
    .O(sig00000ac8)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk0000087b (
    .I0(sig00000b7e),
    .I1(sig00000ba2),
    .I2(sig00000c1e),
    .O(sig00000ac9)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk0000087c (
    .I0(sig00000b7f),
    .I1(sig00000ba3),
    .I2(sig00000c1e),
    .O(sig00000aca)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk0000087d (
    .I0(sig00000b80),
    .I1(sig00000ba4),
    .I2(sig00000c1e),
    .O(sig00000acb)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk0000087e (
    .I0(sig00000b81),
    .I1(sig00000ba5),
    .I2(sig00000c1e),
    .O(sig00000acc)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk0000087f (
    .I0(sig00000b82),
    .I1(sig00000ba6),
    .I2(sig00000c1e),
    .O(sig00000acd)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000880 (
    .I0(sig00000b83),
    .I1(sig00000ba7),
    .I2(sig00000c1e),
    .O(sig00000ace)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000881 (
    .I0(sig00000b84),
    .I1(sig00000ba8),
    .I2(sig00000c1e),
    .O(sig00000acf)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000882 (
    .I0(sig00000b85),
    .I1(sig00000ba9),
    .I2(sig00000c1e),
    .O(sig00000ad0)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000883 (
    .I0(sig00000b86),
    .I1(sig00000baa),
    .I2(sig00000c1e),
    .O(sig00000ad1)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000884 (
    .I0(sig00000b87),
    .I1(sig00000bab),
    .I2(sig00000c1e),
    .O(sig00000ad2)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000885 (
    .I0(sig00000b88),
    .I1(sig00000bac),
    .I2(sig00000c1e),
    .O(sig00000ad3)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000886 (
    .I0(sig00000b89),
    .I1(sig00000bad),
    .I2(sig00000c1e),
    .O(sig00000ad4)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000887 (
    .I0(sig00000b8a),
    .I1(sig00000bae),
    .I2(sig00000c1e),
    .O(sig00000ad5)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000888 (
    .I0(sig00000b8b),
    .I1(sig00000baf),
    .I2(sig00000c1e),
    .O(sig00000ad6)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000889 (
    .I0(sig00000b8c),
    .I1(sig00000bb0),
    .I2(sig00000c1e),
    .O(sig00000ad7)
  );
  MUXCY   blk0000088a (
    .CI(sig00000b0d),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig00000ad8),
    .O(sig00000aea)
  );
  XORCY   blk0000088b (
    .CI(sig00000b0d),
    .LI(sig00000ad8),
    .O(sig00000aeb)
  );
  MUXCY   blk0000088c (
    .CI(sig00000aea),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig00000ad9),
    .O(sig00000aec)
  );
  XORCY   blk0000088d (
    .CI(sig00000aea),
    .LI(sig00000ad9),
    .O(sig00000aed)
  );
  MUXCY   blk0000088e (
    .CI(sig00000aec),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig00000ada),
    .O(sig00000aee)
  );
  XORCY   blk0000088f (
    .CI(sig00000aec),
    .LI(sig00000ada),
    .O(sig00000aef)
  );
  MUXCY   blk00000890 (
    .CI(sig00000aee),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig00000adb),
    .O(sig00000af0)
  );
  XORCY   blk00000891 (
    .CI(sig00000aee),
    .LI(sig00000adb),
    .O(sig00000af1)
  );
  MUXCY   blk00000892 (
    .CI(sig00000af0),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig00000adc),
    .O(sig00000af2)
  );
  XORCY   blk00000893 (
    .CI(sig00000af0),
    .LI(sig00000adc),
    .O(sig00000af3)
  );
  MUXCY   blk00000894 (
    .CI(sig00000af2),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig00000add),
    .O(sig00000af4)
  );
  XORCY   blk00000895 (
    .CI(sig00000af2),
    .LI(sig00000add),
    .O(sig00000af5)
  );
  MUXCY   blk00000896 (
    .CI(sig00000af4),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig00000ade),
    .O(sig00000af6)
  );
  XORCY   blk00000897 (
    .CI(sig00000af4),
    .LI(sig00000ade),
    .O(sig00000af7)
  );
  MUXCY   blk00000898 (
    .CI(sig00000af6),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig00000adf),
    .O(sig00000af8)
  );
  XORCY   blk00000899 (
    .CI(sig00000af6),
    .LI(sig00000adf),
    .O(sig00000af9)
  );
  MUXCY   blk0000089a (
    .CI(sig00000af8),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig00000ae0),
    .O(sig00000afa)
  );
  XORCY   blk0000089b (
    .CI(sig00000af8),
    .LI(sig00000ae0),
    .O(sig00000afb)
  );
  MUXCY   blk0000089c (
    .CI(sig00000afa),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig00000ae1),
    .O(sig00000afc)
  );
  XORCY   blk0000089d (
    .CI(sig00000afa),
    .LI(sig00000ae1),
    .O(sig00000afd)
  );
  MUXCY   blk0000089e (
    .CI(sig00000afc),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig00000ae2),
    .O(sig00000afe)
  );
  XORCY   blk0000089f (
    .CI(sig00000afc),
    .LI(sig00000ae2),
    .O(sig00000aff)
  );
  MUXCY   blk000008a0 (
    .CI(sig00000afe),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig00000ae3),
    .O(sig00000b00)
  );
  XORCY   blk000008a1 (
    .CI(sig00000afe),
    .LI(sig00000ae3),
    .O(sig00000b01)
  );
  MUXCY   blk000008a2 (
    .CI(sig00000b00),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig00000ae4),
    .O(sig00000b02)
  );
  XORCY   blk000008a3 (
    .CI(sig00000b00),
    .LI(sig00000ae4),
    .O(sig00000b03)
  );
  MUXCY   blk000008a4 (
    .CI(sig00000b02),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig00000ae5),
    .O(sig00000b04)
  );
  XORCY   blk000008a5 (
    .CI(sig00000b02),
    .LI(sig00000ae5),
    .O(sig00000b05)
  );
  MUXCY   blk000008a6 (
    .CI(sig00000b04),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig00000ae6),
    .O(sig00000b06)
  );
  XORCY   blk000008a7 (
    .CI(sig00000b04),
    .LI(sig00000ae6),
    .O(sig00000b07)
  );
  MUXCY   blk000008a8 (
    .CI(sig00000b06),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig00000ae7),
    .O(sig00000b08)
  );
  XORCY   blk000008a9 (
    .CI(sig00000b06),
    .LI(sig00000ae7),
    .O(sig00000b09)
  );
  MUXCY   blk000008aa (
    .CI(sig00000b08),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig00000c63),
    .O(sig00000b0a)
  );
  XORCY   blk000008ab (
    .CI(sig00000b08),
    .LI(sig00000c63),
    .O(sig00000b0b)
  );
  MUXCY   blk000008ac (
    .CI(sig00000b0a),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig00000ae8),
    .O(NLW_blk000008ac_O_UNCONNECTED)
  );
  XORCY   blk000008ad (
    .CI(sig00000b0a),
    .LI(sig00000ae8),
    .O(sig00000b0c)
  );
  MUXCY   blk000008ae (
    .CI(sig00000344),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig00000ae9),
    .O(sig00000b0d)
  );
  MUXCY   blk000008af (
    .CI(sig00000b43),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig00000b0e),
    .O(sig00000b20)
  );
  XORCY   blk000008b0 (
    .CI(sig00000b43),
    .LI(sig00000b0e),
    .O(sig00000b21)
  );
  MUXCY   blk000008b1 (
    .CI(sig00000b20),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig00000b0f),
    .O(sig00000b22)
  );
  XORCY   blk000008b2 (
    .CI(sig00000b20),
    .LI(sig00000b0f),
    .O(sig00000b23)
  );
  MUXCY   blk000008b3 (
    .CI(sig00000b22),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig00000b10),
    .O(sig00000b24)
  );
  XORCY   blk000008b4 (
    .CI(sig00000b22),
    .LI(sig00000b10),
    .O(sig00000b25)
  );
  MUXCY   blk000008b5 (
    .CI(sig00000b24),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig00000b11),
    .O(sig00000b26)
  );
  XORCY   blk000008b6 (
    .CI(sig00000b24),
    .LI(sig00000b11),
    .O(sig00000b27)
  );
  MUXCY   blk000008b7 (
    .CI(sig00000b26),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig00000b12),
    .O(sig00000b28)
  );
  XORCY   blk000008b8 (
    .CI(sig00000b26),
    .LI(sig00000b12),
    .O(sig00000b29)
  );
  MUXCY   blk000008b9 (
    .CI(sig00000b28),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig00000b13),
    .O(sig00000b2a)
  );
  XORCY   blk000008ba (
    .CI(sig00000b28),
    .LI(sig00000b13),
    .O(sig00000b2b)
  );
  MUXCY   blk000008bb (
    .CI(sig00000b2a),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig00000b14),
    .O(sig00000b2c)
  );
  XORCY   blk000008bc (
    .CI(sig00000b2a),
    .LI(sig00000b14),
    .O(sig00000b2d)
  );
  MUXCY   blk000008bd (
    .CI(sig00000b2c),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig00000b15),
    .O(sig00000b2e)
  );
  XORCY   blk000008be (
    .CI(sig00000b2c),
    .LI(sig00000b15),
    .O(sig00000b2f)
  );
  MUXCY   blk000008bf (
    .CI(sig00000b2e),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig00000b16),
    .O(sig00000b30)
  );
  XORCY   blk000008c0 (
    .CI(sig00000b2e),
    .LI(sig00000b16),
    .O(sig00000b31)
  );
  MUXCY   blk000008c1 (
    .CI(sig00000b30),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig00000b17),
    .O(sig00000b32)
  );
  XORCY   blk000008c2 (
    .CI(sig00000b30),
    .LI(sig00000b17),
    .O(sig00000b33)
  );
  MUXCY   blk000008c3 (
    .CI(sig00000b32),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig00000b18),
    .O(sig00000b34)
  );
  XORCY   blk000008c4 (
    .CI(sig00000b32),
    .LI(sig00000b18),
    .O(sig00000b35)
  );
  MUXCY   blk000008c5 (
    .CI(sig00000b34),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig00000b19),
    .O(sig00000b36)
  );
  XORCY   blk000008c6 (
    .CI(sig00000b34),
    .LI(sig00000b19),
    .O(sig00000b37)
  );
  MUXCY   blk000008c7 (
    .CI(sig00000b36),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig00000b1a),
    .O(sig00000b38)
  );
  XORCY   blk000008c8 (
    .CI(sig00000b36),
    .LI(sig00000b1a),
    .O(sig00000b39)
  );
  MUXCY   blk000008c9 (
    .CI(sig00000b38),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig00000b1b),
    .O(sig00000b3a)
  );
  XORCY   blk000008ca (
    .CI(sig00000b38),
    .LI(sig00000b1b),
    .O(sig00000b3b)
  );
  MUXCY   blk000008cb (
    .CI(sig00000b3a),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig00000b1c),
    .O(sig00000b3c)
  );
  XORCY   blk000008cc (
    .CI(sig00000b3a),
    .LI(sig00000b1c),
    .O(sig00000b3d)
  );
  MUXCY   blk000008cd (
    .CI(sig00000b3c),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig00000b1d),
    .O(sig00000b3e)
  );
  XORCY   blk000008ce (
    .CI(sig00000b3c),
    .LI(sig00000b1d),
    .O(sig00000b3f)
  );
  MUXCY   blk000008cf (
    .CI(sig00000b3e),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig00000c64),
    .O(sig00000b40)
  );
  XORCY   blk000008d0 (
    .CI(sig00000b3e),
    .LI(sig00000c64),
    .O(sig00000b41)
  );
  MUXCY   blk000008d1 (
    .CI(sig00000b40),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig00000b1e),
    .O(NLW_blk000008d1_O_UNCONNECTED)
  );
  XORCY   blk000008d2 (
    .CI(sig00000b40),
    .LI(sig00000b1e),
    .O(sig00000b42)
  );
  MUXCY   blk000008d3 (
    .CI(sig00000344),
    .DI(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .S(sig00000b1f),
    .O(sig00000b43)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000008d4 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000a90),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000bc3)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000008d5 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000a91),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000bc4)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000008d6 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000a92),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000bc5)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000008d7 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000a93),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000bc6)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000008d8 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000a94),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000bc7)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000008d9 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000a95),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000bc8)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000008da (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000a96),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000bc9)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000008db (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000a97),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000bca)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000008dc (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000a98),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000bcb)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000008dd (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000a99),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000bcc)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000008de (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000a9a),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000bcd)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000008df (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000a9b),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000bce)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000008e0 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000a9c),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000bcf)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000008e1 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000a9d),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000bd0)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000008e2 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000a9e),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000bd1)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000008e3 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000a9f),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000bd2)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000008e4 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000aa0),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000bd3)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000008e5 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000aa1),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000bd4)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000008e6 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000aa2),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000bb1)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000008e7 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000aa3),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000bb2)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000008e8 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000aa4),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000bb3)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000008e9 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000aa5),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000bb4)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000008ea (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000aa6),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000bb5)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000008eb (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000aa7),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000bb6)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000008ec (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000aa8),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000bb7)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000008ed (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000aa9),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000bb8)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000008ee (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000aaa),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000bb9)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000008ef (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000aab),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000bba)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000008f0 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000aac),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000bbb)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000008f1 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000aad),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000bbc)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000008f2 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000aae),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000bbd)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000008f3 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000aaf),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000bbe)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000008f4 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000ab0),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000bbf)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000008f5 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000ab1),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000bc0)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000008f6 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000ab2),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000bc1)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000008f7 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000ab3),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000bc2)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000008f8 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000ab4),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000b69)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000008f9 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000ab5),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000b6a)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000008fa (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000ab6),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000b6b)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000008fb (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000ab7),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000b6c)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000008fc (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000ab8),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000b6d)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000008fd (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000ab9),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000b6e)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000008fe (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000aba),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000b6f)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000008ff (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000abb),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000b70)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000900 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000abc),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000b71)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000901 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000abd),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000b72)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000902 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000abe),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000b73)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000903 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000abf),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000b74)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000904 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000ac0),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000b75)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000905 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000ac1),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000b76)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000906 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000ac2),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000b77)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000907 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000ac3),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000b78)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000908 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000ac4),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000b79)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000909 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000ac5),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000b7a)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000090a (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000ac6),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000868)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000090b (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000ac7),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000869)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000090c (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000ac8),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig0000086a)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000090d (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000ac9),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig0000086b)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000090e (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000aca),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig0000086c)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000090f (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000acb),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig0000086d)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000910 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000acc),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig0000086e)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000911 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000acd),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig0000086f)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000912 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000ace),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000870)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000913 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000acf),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000871)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000914 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000ad0),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000872)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000915 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000ad1),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000873)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000916 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000ad2),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000874)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000917 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000ad3),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000875)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000918 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000ad4),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000876)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000919 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000ad5),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000877)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000091a (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000ad6),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000878)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000091b (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000ad7),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000879)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000091c (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000aeb),
    .Q(sig00000bf9)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000091d (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000aed),
    .Q(sig00000bfa)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000091e (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000aef),
    .Q(sig00000bfb)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000091f (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000af1),
    .Q(sig00000bfc)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000920 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000af3),
    .Q(sig00000bfd)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000921 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000af5),
    .Q(sig00000bfe)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000922 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000af7),
    .Q(sig00000bff)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000923 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000af9),
    .Q(sig00000c00)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000924 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000afb),
    .Q(sig00000c01)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000925 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000afd),
    .Q(sig00000c02)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000926 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000aff),
    .Q(sig00000c03)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000927 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000b01),
    .Q(sig00000c04)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000928 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000b03),
    .Q(sig00000c05)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000929 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000b05),
    .Q(sig00000c06)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000092a (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000b07),
    .Q(sig00000c07)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000092b (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000b09),
    .Q(sig00000c08)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000092c (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000b0b),
    .Q(sig00000c09)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000092d (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000b0c),
    .Q(sig00000c0a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000092e (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000b21),
    .Q(sig00000c0b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000092f (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000b23),
    .Q(sig00000c0c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000930 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000b25),
    .Q(sig00000c0d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000931 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000b27),
    .Q(sig00000c0e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000932 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000b29),
    .Q(sig00000c0f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000933 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000b2b),
    .Q(sig00000c10)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000934 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000b2d),
    .Q(sig00000c11)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000935 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000b2f),
    .Q(sig00000c12)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000936 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000b31),
    .Q(sig00000c13)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000937 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000b33),
    .Q(sig00000c14)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000938 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000b35),
    .Q(sig00000c15)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000939 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000b37),
    .Q(sig00000c16)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000093a (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000b39),
    .Q(sig00000c17)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000093b (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000b3b),
    .Q(sig00000c18)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000093c (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000b3d),
    .Q(sig00000c19)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000093d (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000b3f),
    .Q(sig00000c1a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000093e (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000b41),
    .Q(sig00000c1b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000093f (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000b42),
    .Q(sig00000c1c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000940 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000088e),
    .Q(sig00000c22)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000941 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000c1f),
    .Q(sig00000c1e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000942 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000b44),
    .Q(sig00000c1d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000943 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000893),
    .Q(sig00000c21)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000944 (
    .C(aclk),
    .D(sig00000c1c),
    .Q(sig00000b56)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000945 (
    .C(aclk),
    .D(sig00000c1b),
    .Q(sig00000b55)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000946 (
    .C(aclk),
    .D(sig00000c1a),
    .Q(sig00000b54)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000947 (
    .C(aclk),
    .D(sig00000c19),
    .Q(sig00000b53)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000948 (
    .C(aclk),
    .D(sig00000c18),
    .Q(sig00000b52)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000949 (
    .C(aclk),
    .D(sig00000c17),
    .Q(sig00000b51)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000094a (
    .C(aclk),
    .D(sig00000c16),
    .Q(sig00000b50)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000094b (
    .C(aclk),
    .D(sig00000c15),
    .Q(sig00000b4f)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000094c (
    .C(aclk),
    .D(sig00000c14),
    .Q(sig00000b4e)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000094d (
    .C(aclk),
    .D(sig00000c13),
    .Q(sig00000b4d)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000094e (
    .C(aclk),
    .D(sig00000c12),
    .Q(sig00000b4c)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000094f (
    .C(aclk),
    .D(sig00000c11),
    .Q(sig00000b4b)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000950 (
    .C(aclk),
    .D(sig00000c10),
    .Q(sig00000b4a)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000951 (
    .C(aclk),
    .D(sig00000c0f),
    .Q(sig00000b49)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000952 (
    .C(aclk),
    .D(sig00000c0e),
    .Q(sig00000b48)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000953 (
    .C(aclk),
    .D(sig00000c0d),
    .Q(sig00000b47)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000954 (
    .C(aclk),
    .D(sig00000c0c),
    .Q(sig00000b46)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000955 (
    .C(aclk),
    .D(sig00000c0b),
    .Q(sig00000b45)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000956 (
    .C(aclk),
    .D(sig00000c0a),
    .Q(sig00000b68)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000957 (
    .C(aclk),
    .D(sig00000c09),
    .Q(sig00000b67)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000958 (
    .C(aclk),
    .D(sig00000c08),
    .Q(sig00000b66)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000959 (
    .C(aclk),
    .D(sig00000c07),
    .Q(sig00000b65)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000095a (
    .C(aclk),
    .D(sig00000c06),
    .Q(sig00000b64)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000095b (
    .C(aclk),
    .D(sig00000c05),
    .Q(sig00000b63)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000095c (
    .C(aclk),
    .D(sig00000c04),
    .Q(sig00000b62)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000095d (
    .C(aclk),
    .D(sig00000c03),
    .Q(sig00000b61)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000095e (
    .C(aclk),
    .D(sig00000c02),
    .Q(sig00000b60)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000095f (
    .C(aclk),
    .D(sig00000c01),
    .Q(sig00000b5f)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000960 (
    .C(aclk),
    .D(sig00000c00),
    .Q(sig00000b5e)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000961 (
    .C(aclk),
    .D(sig00000bff),
    .Q(sig00000b5d)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000962 (
    .C(aclk),
    .D(sig00000bfe),
    .Q(sig00000b5c)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000963 (
    .C(aclk),
    .D(sig00000bfd),
    .Q(sig00000b5b)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000964 (
    .C(aclk),
    .D(sig00000bfc),
    .Q(sig00000b5a)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000965 (
    .C(aclk),
    .D(sig00000bfb),
    .Q(sig00000b59)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000966 (
    .C(aclk),
    .D(sig00000bfa),
    .Q(sig00000b58)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000967 (
    .C(aclk),
    .D(sig00000bf9),
    .Q(sig00000b57)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000968 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000b7a),
    .Q(sig0000088b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000969 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000b79),
    .Q(sig0000088a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000096a (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000b78),
    .Q(sig00000889)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000096b (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000b77),
    .Q(sig00000888)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000096c (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000b76),
    .Q(sig00000887)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000096d (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000b75),
    .Q(sig00000886)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000096e (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000b74),
    .Q(sig00000885)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000096f (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000b73),
    .Q(sig00000884)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000970 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000b72),
    .Q(sig00000883)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000971 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000b71),
    .Q(sig00000882)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000972 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000b70),
    .Q(sig00000881)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000973 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000b6f),
    .Q(sig00000880)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000974 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000b6e),
    .Q(sig0000087f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000975 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000b6d),
    .Q(sig0000087e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000976 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000b6c),
    .Q(sig0000087d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000977 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000b6b),
    .Q(sig0000087c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000978 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000b6a),
    .Q(sig0000087b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000979 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000b69),
    .Q(sig0000087a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000097a (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000b9e),
    .Q(sig00000b8c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000097b (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000b9d),
    .Q(sig00000b8b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000097c (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000b9c),
    .Q(sig00000b8a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000097d (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000b9b),
    .Q(sig00000b89)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000097e (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000b9a),
    .Q(sig00000b88)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000097f (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000b99),
    .Q(sig00000b87)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000980 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000b98),
    .Q(sig00000b86)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000981 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000b97),
    .Q(sig00000b85)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000982 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000b96),
    .Q(sig00000b84)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000983 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000b95),
    .Q(sig00000b83)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000984 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000b94),
    .Q(sig00000b82)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000985 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000b93),
    .Q(sig00000b81)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000986 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000b92),
    .Q(sig00000b80)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000987 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000b91),
    .Q(sig00000b7f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000988 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000b90),
    .Q(sig00000b7e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000989 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000b8f),
    .Q(sig00000b7d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000098a (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000b8e),
    .Q(sig00000b7c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000098b (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000b8d),
    .Q(sig00000b7b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000098c (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000b68),
    .Q(sig00000be6)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000098d (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000b67),
    .Q(sig00000be5)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000098e (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000b66),
    .Q(sig00000be4)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000098f (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000b65),
    .Q(sig00000be3)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000990 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000b64),
    .Q(sig00000be2)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000991 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000b63),
    .Q(sig00000be1)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000992 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000b62),
    .Q(sig00000be0)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000993 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000b61),
    .Q(sig00000bdf)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000994 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000b60),
    .Q(sig00000bde)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000995 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000b5f),
    .Q(sig00000bdd)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000996 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000b5e),
    .Q(sig00000bdc)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000997 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000b5d),
    .Q(sig00000bdb)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000998 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000b5c),
    .Q(sig00000bda)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000999 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000b5b),
    .Q(sig00000bd9)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000099a (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000b5a),
    .Q(sig00000bd8)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000099b (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000b59),
    .Q(sig00000bd7)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000099c (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000b58),
    .Q(sig00000bd6)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000099d (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000b57),
    .Q(sig00000bd5)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000099e (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000bd4),
    .Q(sig00000bf8)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000099f (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000bd3),
    .Q(sig00000bf7)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000009a0 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000bd2),
    .Q(sig00000bf6)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000009a1 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000bd1),
    .Q(sig00000bf5)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000009a2 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000bd0),
    .Q(sig00000bf4)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000009a3 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000bcf),
    .Q(sig00000bf3)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000009a4 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000bce),
    .Q(sig00000bf2)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000009a5 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000bcd),
    .Q(sig00000bf1)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000009a6 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000bcc),
    .Q(sig00000bf0)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000009a7 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000bcb),
    .Q(sig00000bef)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000009a8 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000bca),
    .Q(sig00000bee)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000009a9 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000bc9),
    .Q(sig00000bed)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000009aa (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000bc8),
    .Q(sig00000bec)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000009ab (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000bc7),
    .Q(sig00000beb)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000009ac (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000bc6),
    .Q(sig00000bea)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000009ad (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000bc5),
    .Q(sig00000be9)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000009ae (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000bc4),
    .Q(sig00000be8)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000009af (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000bc3),
    .Q(sig00000be7)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000009b0 (
    .I0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .I1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .I2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .I3(sig0000087a),
    .I4(sig0000088c),
    .I5(sig0000088d),
    .O(sig00000c23)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000009b1 (
    .I0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .I1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .I2(sig0000087a),
    .I3(sig0000087b),
    .I4(sig0000088c),
    .I5(sig0000088d),
    .O(sig00000c24)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000009b2 (
    .I0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .I1(sig0000087a),
    .I2(sig0000087b),
    .I3(sig0000087c),
    .I4(sig0000088c),
    .I5(sig0000088d),
    .O(sig00000c25)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000009b3 (
    .I0(sig0000087a),
    .I1(sig0000087b),
    .I2(sig0000087c),
    .I3(sig0000087d),
    .I4(sig0000088c),
    .I5(sig0000088d),
    .O(sig00000c26)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000009b4 (
    .I0(sig0000087b),
    .I1(sig0000087c),
    .I2(sig0000087d),
    .I3(sig0000087e),
    .I4(sig0000088c),
    .I5(sig0000088d),
    .O(sig00000c27)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000009b5 (
    .I0(sig0000087c),
    .I1(sig0000087d),
    .I2(sig0000087e),
    .I3(sig0000087f),
    .I4(sig0000088c),
    .I5(sig0000088d),
    .O(sig00000c28)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000009b6 (
    .I0(sig0000087d),
    .I1(sig0000087e),
    .I2(sig0000087f),
    .I3(sig00000880),
    .I4(sig0000088c),
    .I5(sig0000088d),
    .O(sig00000c29)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000009b7 (
    .I0(sig0000087e),
    .I1(sig0000087f),
    .I2(sig00000880),
    .I3(sig00000881),
    .I4(sig0000088c),
    .I5(sig0000088d),
    .O(sig00000c2a)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000009b8 (
    .I0(sig0000087f),
    .I1(sig00000880),
    .I2(sig00000881),
    .I3(sig00000882),
    .I4(sig0000088c),
    .I5(sig0000088d),
    .O(sig00000c2b)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000009b9 (
    .I0(sig00000880),
    .I1(sig00000881),
    .I2(sig00000882),
    .I3(sig00000883),
    .I4(sig0000088c),
    .I5(sig0000088d),
    .O(sig00000c2c)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000009ba (
    .I0(sig00000881),
    .I1(sig00000882),
    .I2(sig00000883),
    .I3(sig00000884),
    .I4(sig0000088c),
    .I5(sig0000088d),
    .O(sig00000c2d)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000009bb (
    .I0(sig00000882),
    .I1(sig00000883),
    .I2(sig00000884),
    .I3(sig00000885),
    .I4(sig0000088c),
    .I5(sig0000088d),
    .O(sig00000c2e)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000009bc (
    .I0(sig00000883),
    .I1(sig00000884),
    .I2(sig00000885),
    .I3(sig00000886),
    .I4(sig0000088c),
    .I5(sig0000088d),
    .O(sig00000c2f)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000009bd (
    .I0(sig00000884),
    .I1(sig00000885),
    .I2(sig00000886),
    .I3(sig00000887),
    .I4(sig0000088c),
    .I5(sig0000088d),
    .O(sig00000c30)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000009be (
    .I0(sig00000885),
    .I1(sig00000886),
    .I2(sig00000887),
    .I3(sig00000888),
    .I4(sig0000088c),
    .I5(sig0000088d),
    .O(sig00000c31)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000009bf (
    .I0(sig00000886),
    .I1(sig00000887),
    .I2(sig00000888),
    .I3(sig00000889),
    .I4(sig0000088c),
    .I5(sig0000088d),
    .O(sig00000c32)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000009c0 (
    .I0(sig00000887),
    .I1(sig00000888),
    .I2(sig00000889),
    .I3(sig0000088a),
    .I4(sig0000088c),
    .I5(sig0000088d),
    .O(sig00000c33)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000009c1 (
    .I0(sig00000888),
    .I1(sig00000889),
    .I2(sig0000088a),
    .I3(sig0000088b),
    .I4(sig0000088c),
    .I5(sig0000088d),
    .O(sig00000c34)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000009c2 (
    .I0(sig00000889),
    .I1(sig0000088a),
    .I2(sig0000088b),
    .I3(sig0000088b),
    .I4(sig0000088c),
    .I5(sig0000088d),
    .O(sig00000c35)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000009c3 (
    .I0(sig0000088a),
    .I1(sig0000088b),
    .I2(sig0000088b),
    .I3(sig0000088b),
    .I4(sig0000088c),
    .I5(sig0000088d),
    .O(sig00000c36)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000009c4 (
    .I0(sig0000088b),
    .I1(sig0000088b),
    .I2(sig0000088b),
    .I3(sig0000088b),
    .I4(sig0000088c),
    .I5(sig0000088d),
    .O(sig00000c37)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000009c5 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000c23),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(NLW_blk000009c5_Q_UNCONNECTED)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000009c6 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000c24),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(NLW_blk000009c6_Q_UNCONNECTED)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000009c7 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000c25),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(NLW_blk000009c7_Q_UNCONNECTED)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000009c8 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000c26),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig0000008c)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000009c9 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000c27),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig0000008d)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000009ca (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000c28),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig0000008e)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000009cb (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000c29),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig0000008f)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000009cc (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000c2a),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000090)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000009cd (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000c2b),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000091)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000009ce (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000c2c),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000092)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000009cf (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000c2d),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000093)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000009d0 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000c2e),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000094)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000009d1 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000c2f),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000095)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000009d2 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000c30),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000096)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000009d3 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000c31),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000097)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000009d4 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000c32),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000098)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000009d5 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000c33),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000099)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000009d6 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000c34),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig0000009a)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000009d7 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000c35),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig0000009b)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000009d8 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000c36),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(NLW_blk000009d8_Q_UNCONNECTED)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000009d9 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000c37),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(NLW_blk000009d9_Q_UNCONNECTED)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000009da (
    .I0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .I1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .I2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .I3(sig00000868),
    .I4(sig0000088c),
    .I5(sig0000088d),
    .O(sig00000c38)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000009db (
    .I0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .I1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .I2(sig00000868),
    .I3(sig00000869),
    .I4(sig0000088c),
    .I5(sig0000088d),
    .O(sig00000c39)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000009dc (
    .I0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .I1(sig00000868),
    .I2(sig00000869),
    .I3(sig0000086a),
    .I4(sig0000088c),
    .I5(sig0000088d),
    .O(sig00000c3a)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000009dd (
    .I0(sig00000868),
    .I1(sig00000869),
    .I2(sig0000086a),
    .I3(sig0000086b),
    .I4(sig0000088c),
    .I5(sig0000088d),
    .O(sig00000c3b)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000009de (
    .I0(sig00000869),
    .I1(sig0000086a),
    .I2(sig0000086b),
    .I3(sig0000086c),
    .I4(sig0000088c),
    .I5(sig0000088d),
    .O(sig00000c3c)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000009df (
    .I0(sig0000086a),
    .I1(sig0000086b),
    .I2(sig0000086c),
    .I3(sig0000086d),
    .I4(sig0000088c),
    .I5(sig0000088d),
    .O(sig00000c3d)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000009e0 (
    .I0(sig0000086b),
    .I1(sig0000086c),
    .I2(sig0000086d),
    .I3(sig0000086e),
    .I4(sig0000088c),
    .I5(sig0000088d),
    .O(sig00000c3e)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000009e1 (
    .I0(sig0000086c),
    .I1(sig0000086d),
    .I2(sig0000086e),
    .I3(sig0000086f),
    .I4(sig0000088c),
    .I5(sig0000088d),
    .O(sig00000c3f)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000009e2 (
    .I0(sig0000086d),
    .I1(sig0000086e),
    .I2(sig0000086f),
    .I3(sig00000870),
    .I4(sig0000088c),
    .I5(sig0000088d),
    .O(sig00000c40)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000009e3 (
    .I0(sig0000086e),
    .I1(sig0000086f),
    .I2(sig00000870),
    .I3(sig00000871),
    .I4(sig0000088c),
    .I5(sig0000088d),
    .O(sig00000c41)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000009e4 (
    .I0(sig0000086f),
    .I1(sig00000870),
    .I2(sig00000871),
    .I3(sig00000872),
    .I4(sig0000088c),
    .I5(sig0000088d),
    .O(sig00000c42)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000009e5 (
    .I0(sig00000870),
    .I1(sig00000871),
    .I2(sig00000872),
    .I3(sig00000873),
    .I4(sig0000088c),
    .I5(sig0000088d),
    .O(sig00000c43)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000009e6 (
    .I0(sig00000871),
    .I1(sig00000872),
    .I2(sig00000873),
    .I3(sig00000874),
    .I4(sig0000088c),
    .I5(sig0000088d),
    .O(sig00000c44)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000009e7 (
    .I0(sig00000872),
    .I1(sig00000873),
    .I2(sig00000874),
    .I3(sig00000875),
    .I4(sig0000088c),
    .I5(sig0000088d),
    .O(sig00000c45)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000009e8 (
    .I0(sig00000873),
    .I1(sig00000874),
    .I2(sig00000875),
    .I3(sig00000876),
    .I4(sig0000088c),
    .I5(sig0000088d),
    .O(sig00000c46)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000009e9 (
    .I0(sig00000874),
    .I1(sig00000875),
    .I2(sig00000876),
    .I3(sig00000877),
    .I4(sig0000088c),
    .I5(sig0000088d),
    .O(sig00000c47)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000009ea (
    .I0(sig00000875),
    .I1(sig00000876),
    .I2(sig00000877),
    .I3(sig00000878),
    .I4(sig0000088c),
    .I5(sig0000088d),
    .O(sig00000c48)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000009eb (
    .I0(sig00000876),
    .I1(sig00000877),
    .I2(sig00000878),
    .I3(sig00000879),
    .I4(sig0000088c),
    .I5(sig0000088d),
    .O(sig00000c49)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000009ec (
    .I0(sig00000877),
    .I1(sig00000878),
    .I2(sig00000879),
    .I3(sig00000879),
    .I4(sig0000088c),
    .I5(sig0000088d),
    .O(sig00000c4a)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000009ed (
    .I0(sig00000878),
    .I1(sig00000879),
    .I2(sig00000879),
    .I3(sig00000879),
    .I4(sig0000088c),
    .I5(sig0000088d),
    .O(sig00000c4b)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000009ee (
    .I0(sig00000879),
    .I1(sig00000879),
    .I2(sig00000879),
    .I3(sig00000879),
    .I4(sig0000088c),
    .I5(sig0000088d),
    .O(sig00000c4c)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000009ef (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000c38),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(NLW_blk000009ef_Q_UNCONNECTED)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000009f0 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000c39),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(NLW_blk000009f0_Q_UNCONNECTED)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000009f1 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000c3a),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(NLW_blk000009f1_Q_UNCONNECTED)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000009f2 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000c3b),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig0000007c)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000009f3 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000c3c),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig0000007d)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000009f4 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000c3d),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig0000007e)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000009f5 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000c3e),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig0000007f)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000009f6 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000c3f),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000080)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000009f7 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000c40),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000081)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000009f8 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000c41),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000082)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000009f9 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000c42),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000083)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000009fa (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000c43),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000084)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000009fb (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000c44),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000085)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000009fc (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000c45),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000086)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000009fd (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000c46),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000087)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000009fe (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000c47),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000088)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000009ff (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000c48),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig00000089)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000a00 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000c49),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig0000008a)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000a01 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000c4a),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(sig0000008b)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000a02 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000c4b),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(NLW_blk00000a02_Q_UNCONNECTED)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000a03 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000c4c),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(NLW_blk00000a03_Q_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000a04 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000008b),
    .Q(sig00000012)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000a05 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000008a),
    .Q(sig00000011)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000a06 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000089),
    .Q(sig00000010)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000a07 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000088),
    .Q(sig0000000f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000a08 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000087),
    .Q(sig0000000e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000a09 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000086),
    .Q(sig0000000d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000a0a (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000085),
    .Q(sig0000000c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000a0b (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000084),
    .Q(sig0000000b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000a0c (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000083),
    .Q(sig0000000a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000a0d (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000082),
    .Q(sig00000009)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000a0e (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000081),
    .Q(sig00000008)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000a0f (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000080),
    .Q(sig00000007)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000a10 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000007f),
    .Q(sig00000006)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000a11 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000007e),
    .Q(sig00000005)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000a12 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000007d),
    .Q(sig00000004)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000a13 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000007c),
    .Q(sig00000003)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000a14 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000009b),
    .Q(sig00000022)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000a15 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000009a),
    .Q(sig00000021)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000a16 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000099),
    .Q(sig00000020)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000a17 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000098),
    .Q(sig0000001f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000a18 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000097),
    .Q(sig0000001e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000a19 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000096),
    .Q(sig0000001d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000a1a (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000095),
    .Q(sig0000001c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000a1b (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000094),
    .Q(sig0000001b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000a1c (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000093),
    .Q(sig0000001a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000a1d (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000092),
    .Q(sig00000019)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000a1e (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000091),
    .Q(sig00000018)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000a1f (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000090),
    .Q(sig00000017)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000a20 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000008f),
    .Q(sig00000016)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000a21 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000008e),
    .Q(sig00000015)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000a22 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000008d),
    .Q(sig00000014)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000a23 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig0000008c),
    .Q(sig00000013)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000a24 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000000ca),
    .Q(sig00000c4d)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000a25 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000c4d),
    .R(NLW_blk00000a25_R_UNCONNECTED),
    .Q(sig00000c4e)
  );
  FDR #(
    .INIT ( 1'b0 ))
  blk00000a26 (
    .C(aclk),
    .D(sig00000c4e),
    .R(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .Q(NLW_blk00000a26_Q_UNCONNECTED)
  );
  LUT4 #(
    .INIT ( 16'hAAA9 ))
  blk00000a27 (
    .I0(sig00000064),
    .I1(sig00000053),
    .I2(sig00000062),
    .I3(sig00000063),
    .O(sig00000055)
  );
  LUT6 #(
    .INIT ( 64'h5555555700000003 ))
  blk00000a28 (
    .I0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/dv_resolved_prev ),
    .I1(sig00000064),
    .I2(sig00000063),
    .I3(sig00000062),
    .I4(sig00000053),
    .I5(sig00000001),
    .O(sig0000005c)
  );
  LUT5 #(
    .INIT ( 32'h88888000 ))
  blk00000a29 (
    .I0(sig00000067),
    .I1(sig0000006a),
    .I2(sig00000066),
    .I3(sig00000052),
    .I4(sig00000002),
    .O(sig0000005f)
  );
  LUT4 #(
    .INIT ( 16'hAA80 ))
  blk00000a2a (
    .I0(sig00000067),
    .I1(sig00000066),
    .I2(sig00000052),
    .I3(sig00000002),
    .O(sig00000059)
  );
  LUT3 #(
    .INIT ( 8'hA9 ))
  blk00000a2b (
    .I0(sig00000063),
    .I1(sig00000053),
    .I2(sig00000062),
    .O(sig00000056)
  );
  LUT5 #(
    .INIT ( 32'h00000008 ))
  blk00000a2c (
    .I0(sig00000001),
    .I1(sig00000053),
    .I2(sig00000062),
    .I3(sig00000063),
    .I4(sig00000064),
    .O(sig00000060)
  );
  LUT4 #(
    .INIT ( 16'hF888 ))
  blk00000a2d (
    .I0(sig00000067),
    .I1(sig00000002),
    .I2(sig00000066),
    .I3(sig00000052),
    .O(sig0000005d)
  );
  LUT4 #(
    .INIT ( 16'h7FFF ))
  blk00000a2e (
    .I0(sig00000029),
    .I1(sig0000002a),
    .I2(sig00000027),
    .I3(sig00000028),
    .O(sig00000052)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000a2f (
    .I0(sig00000062),
    .I1(sig00000053),
    .O(sig00000057)
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  blk00000a30 (
    .I0(sig00000069),
    .I1(sig0000002c),
    .O(sig0000005e)
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  blk00000a31 (
    .I0(sig00000002),
    .I1(sig0000006f),
    .O(sig00000061)
  );
  LUT2 #(
    .INIT ( 4'hB ))
  blk00000a32 (
    .I0(sig00000065),
    .I1(sig0000006d),
    .O(s_axis_config_tready)
  );
  LUT2 #(
    .INIT ( 4'hB ))
  blk00000a33 (
    .I0(sig00000002),
    .I1(sig0000006f),
    .O(s_axis_data_tready)
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  blk00000a34 (
    .I0(sig000000c8),
    .I1(sig00000072),
    .O(sig00000137)
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  blk00000a35 (
    .I0(sig000000c7),
    .I1(sig00000072),
    .O(sig00000135)
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  blk00000a36 (
    .I0(sig000000c6),
    .I1(sig00000072),
    .O(sig00000134)
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  blk00000a37 (
    .I0(sig000000c5),
    .I1(sig00000072),
    .O(sig00000136)
  );
  LUT3 #(
    .INIT ( 8'hB0 ))
  blk00000a38 (
    .I0(sig00000121),
    .I1(sig00000002),
    .I2(sig0000002d),
    .O(sig0000011d)
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  blk00000a39 (
    .I0(sig00000027),
    .I1(sig00000121),
    .O(sig0000012c)
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  blk00000a3a (
    .I0(sig00000028),
    .I1(sig00000121),
    .O(sig0000012a)
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  blk00000a3b (
    .I0(sig00000029),
    .I1(sig00000121),
    .O(sig00000129)
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  blk00000a3c (
    .I0(sig0000002a),
    .I1(sig00000121),
    .O(sig0000012b)
  );
  LUT3 #(
    .INIT ( 8'hF2 ))
  blk00000a3d (
    .I0(sig00000002),
    .I1(sig00000121),
    .I2(sig0000002d),
    .O(sig0000011c)
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  blk00000a3e (
    .I0(sig00000205),
    .I1(sig00000150),
    .O(sig00000144)
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  blk00000a3f (
    .I0(sig00000206),
    .I1(sig00000150),
    .O(sig00000146)
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  blk00000a40 (
    .I0(sig00000207),
    .I1(sig00000150),
    .O(sig00000147)
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  blk00000a41 (
    .I0(sig00000208),
    .I1(sig00000150),
    .O(sig00000145)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk00000a42 (
    .I0(sig000000c2),
    .I1(sig000000c9),
    .I2(sig000001e1),
    .O(sig00000161)
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  blk00000a43 (
    .I0(sig0000020a),
    .I1(sig00000229),
    .O(sig00000212)
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  blk00000a44 (
    .I0(sig0000020b),
    .I1(sig00000229),
    .O(sig00000214)
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  blk00000a45 (
    .I0(sig0000020c),
    .I1(sig00000229),
    .O(sig00000215)
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  blk00000a46 (
    .I0(sig0000020d),
    .I1(sig00000229),
    .O(sig00000213)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000a47 (
    .I0(sig000002b0),
    .I1(sig000002d3),
    .O(sig00000333)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000a48 (
    .I0(sig000002ba),
    .I1(sig000002dd),
    .O(sig00000329)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000a49 (
    .I0(sig000002bb),
    .I1(sig000002de),
    .O(sig00000328)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000a4a (
    .I0(sig000002bc),
    .I1(sig000002df),
    .O(sig00000327)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000a4b (
    .I0(sig000002bd),
    .I1(sig000002e0),
    .O(sig00000326)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000a4c (
    .I0(sig000002be),
    .I1(sig000002e1),
    .O(sig00000325)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000a4d (
    .I0(sig000002bf),
    .I1(sig000002e2),
    .O(sig00000324)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000a4e (
    .I0(sig000002b1),
    .I1(sig000002d4),
    .O(sig00000332)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000a4f (
    .I0(sig000002b2),
    .I1(sig000002d5),
    .O(sig00000331)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000a50 (
    .I0(sig000002b3),
    .I1(sig000002d6),
    .O(sig00000330)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000a51 (
    .I0(sig000002b4),
    .I1(sig000002d7),
    .O(sig0000032f)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000a52 (
    .I0(sig000002b5),
    .I1(sig000002d8),
    .O(sig0000032e)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000a53 (
    .I0(sig000002b6),
    .I1(sig000002d9),
    .O(sig0000032d)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000a54 (
    .I0(sig000002b7),
    .I1(sig000002da),
    .O(sig0000032c)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000a55 (
    .I0(sig000002b8),
    .I1(sig000002db),
    .O(sig0000032b)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000a56 (
    .I0(sig000002b9),
    .I1(sig000002dc),
    .O(sig0000032a)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000a57 (
    .I0(sig000002b0),
    .I1(sig000002d3),
    .O(sig00000365)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000a58 (
    .I0(sig000002ba),
    .I1(sig000002dd),
    .O(sig0000035b)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000a59 (
    .I0(sig000002bb),
    .I1(sig000002de),
    .O(sig0000035a)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000a5a (
    .I0(sig000002bc),
    .I1(sig000002df),
    .O(sig00000359)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000a5b (
    .I0(sig000002bd),
    .I1(sig000002e0),
    .O(sig00000358)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000a5c (
    .I0(sig000002be),
    .I1(sig000002e1),
    .O(sig00000357)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000a5d (
    .I0(sig000002bf),
    .I1(sig000002e2),
    .O(sig00000356)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000a5e (
    .I0(sig000002b1),
    .I1(sig000002d4),
    .O(sig00000364)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000a5f (
    .I0(sig000002b2),
    .I1(sig000002d5),
    .O(sig00000363)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000a60 (
    .I0(sig000002b3),
    .I1(sig000002d6),
    .O(sig00000362)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000a61 (
    .I0(sig000002b4),
    .I1(sig000002d7),
    .O(sig00000361)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000a62 (
    .I0(sig000002b5),
    .I1(sig000002d8),
    .O(sig00000360)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000a63 (
    .I0(sig000002b6),
    .I1(sig000002d9),
    .O(sig0000035f)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000a64 (
    .I0(sig000002b7),
    .I1(sig000002da),
    .O(sig0000035e)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000a65 (
    .I0(sig000002b8),
    .I1(sig000002db),
    .O(sig0000035d)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000a66 (
    .I0(sig000002b9),
    .I1(sig000002dc),
    .O(sig0000035c)
  );
  LUT4 #(
    .INIT ( 16'h3CAA ))
  blk00000a67 (
    .I0(sig000001e2),
    .I1(sig000001f3),
    .I2(sig00000532),
    .I3(sig0000052d),
    .O(sig000003e8)
  );
  LUT4 #(
    .INIT ( 16'h3CAA ))
  blk00000a68 (
    .I0(sig000001e3),
    .I1(sig000001f4),
    .I2(sig00000532),
    .I3(sig0000052d),
    .O(sig000003e9)
  );
  LUT4 #(
    .INIT ( 16'h3CAA ))
  blk00000a69 (
    .I0(sig000001e4),
    .I1(sig000001f5),
    .I2(sig00000532),
    .I3(sig0000052d),
    .O(sig000003ea)
  );
  LUT4 #(
    .INIT ( 16'h3CAA ))
  blk00000a6a (
    .I0(sig000001e6),
    .I1(sig000001f7),
    .I2(sig00000532),
    .I3(sig0000052d),
    .O(sig000003ec)
  );
  LUT4 #(
    .INIT ( 16'h3CAA ))
  blk00000a6b (
    .I0(sig000001e7),
    .I1(sig000001f8),
    .I2(sig00000532),
    .I3(sig0000052d),
    .O(sig000003ed)
  );
  LUT4 #(
    .INIT ( 16'h3CAA ))
  blk00000a6c (
    .I0(sig000001e5),
    .I1(sig000001f6),
    .I2(sig00000532),
    .I3(sig0000052d),
    .O(sig000003eb)
  );
  LUT4 #(
    .INIT ( 16'h3CAA ))
  blk00000a6d (
    .I0(sig000001e8),
    .I1(sig000001f9),
    .I2(sig00000532),
    .I3(sig0000052d),
    .O(sig000003ee)
  );
  LUT4 #(
    .INIT ( 16'h3CAA ))
  blk00000a6e (
    .I0(sig000001e9),
    .I1(sig000001fa),
    .I2(sig00000532),
    .I3(sig0000052d),
    .O(sig000003ef)
  );
  LUT4 #(
    .INIT ( 16'h3CAA ))
  blk00000a6f (
    .I0(sig000001ea),
    .I1(sig000001fb),
    .I2(sig00000532),
    .I3(sig0000052d),
    .O(sig000003f0)
  );
  LUT4 #(
    .INIT ( 16'h3CAA ))
  blk00000a70 (
    .I0(sig000001eb),
    .I1(sig000001fc),
    .I2(sig00000532),
    .I3(sig0000052d),
    .O(sig000003f1)
  );
  LUT4 #(
    .INIT ( 16'h3CAA ))
  blk00000a71 (
    .I0(sig000001ed),
    .I1(sig000001fe),
    .I2(sig00000532),
    .I3(sig0000052d),
    .O(sig000003f3)
  );
  LUT4 #(
    .INIT ( 16'h3CAA ))
  blk00000a72 (
    .I0(sig000001ee),
    .I1(sig000001ff),
    .I2(sig00000532),
    .I3(sig0000052d),
    .O(sig000003f4)
  );
  LUT4 #(
    .INIT ( 16'h3CAA ))
  blk00000a73 (
    .I0(sig000001ec),
    .I1(sig000001fd),
    .I2(sig00000532),
    .I3(sig0000052d),
    .O(sig000003f2)
  );
  LUT4 #(
    .INIT ( 16'h3CAA ))
  blk00000a74 (
    .I0(sig000001ef),
    .I1(sig00000200),
    .I2(sig00000532),
    .I3(sig0000052d),
    .O(sig000003f5)
  );
  LUT4 #(
    .INIT ( 16'h3CAA ))
  blk00000a75 (
    .I0(sig000001f0),
    .I1(sig00000201),
    .I2(sig00000532),
    .I3(sig0000052d),
    .O(sig000003f6)
  );
  LUT4 #(
    .INIT ( 16'h3CAA ))
  blk00000a76 (
    .I0(sig000001f1),
    .I1(sig00000202),
    .I2(sig00000532),
    .I3(sig0000052d),
    .O(sig000003f7)
  );
  LUT4 #(
    .INIT ( 16'h7D28 ))
  blk00000a77 (
    .I0(sig0000052d),
    .I1(sig00000203),
    .I2(sig00000532),
    .I3(sig000001f2),
    .O(sig000003f8)
  );
  LUT4 #(
    .INIT ( 16'hC3AA ))
  blk00000a78 (
    .I0(sig000001f3),
    .I1(sig000001e2),
    .I2(sig00000532),
    .I3(sig0000052d),
    .O(sig0000041e)
  );
  LUT4 #(
    .INIT ( 16'hC3AA ))
  blk00000a79 (
    .I0(sig000001f4),
    .I1(sig000001e3),
    .I2(sig00000532),
    .I3(sig0000052d),
    .O(sig0000041f)
  );
  LUT4 #(
    .INIT ( 16'hC3AA ))
  blk00000a7a (
    .I0(sig000001f5),
    .I1(sig000001e4),
    .I2(sig00000532),
    .I3(sig0000052d),
    .O(sig00000420)
  );
  LUT4 #(
    .INIT ( 16'hC3AA ))
  blk00000a7b (
    .I0(sig000001f6),
    .I1(sig000001e5),
    .I2(sig00000532),
    .I3(sig0000052d),
    .O(sig00000421)
  );
  LUT4 #(
    .INIT ( 16'hC3AA ))
  blk00000a7c (
    .I0(sig000001f7),
    .I1(sig000001e6),
    .I2(sig00000532),
    .I3(sig0000052d),
    .O(sig00000422)
  );
  LUT4 #(
    .INIT ( 16'hC3AA ))
  blk00000a7d (
    .I0(sig000001f9),
    .I1(sig000001e8),
    .I2(sig00000532),
    .I3(sig0000052d),
    .O(sig00000424)
  );
  LUT4 #(
    .INIT ( 16'hC3AA ))
  blk00000a7e (
    .I0(sig000001fa),
    .I1(sig000001e9),
    .I2(sig00000532),
    .I3(sig0000052d),
    .O(sig00000425)
  );
  LUT4 #(
    .INIT ( 16'hC3AA ))
  blk00000a7f (
    .I0(sig000001f8),
    .I1(sig000001e7),
    .I2(sig00000532),
    .I3(sig0000052d),
    .O(sig00000423)
  );
  LUT4 #(
    .INIT ( 16'hC3AA ))
  blk00000a80 (
    .I0(sig000001fb),
    .I1(sig000001ea),
    .I2(sig00000532),
    .I3(sig0000052d),
    .O(sig00000426)
  );
  LUT4 #(
    .INIT ( 16'hC3AA ))
  blk00000a81 (
    .I0(sig000001fc),
    .I1(sig000001eb),
    .I2(sig00000532),
    .I3(sig0000052d),
    .O(sig00000427)
  );
  LUT4 #(
    .INIT ( 16'hC3AA ))
  blk00000a82 (
    .I0(sig000001fd),
    .I1(sig000001ec),
    .I2(sig00000532),
    .I3(sig0000052d),
    .O(sig00000428)
  );
  LUT4 #(
    .INIT ( 16'hC3AA ))
  blk00000a83 (
    .I0(sig000001fe),
    .I1(sig000001ed),
    .I2(sig00000532),
    .I3(sig0000052d),
    .O(sig00000429)
  );
  LUT4 #(
    .INIT ( 16'hC3AA ))
  blk00000a84 (
    .I0(sig00000200),
    .I1(sig000001ef),
    .I2(sig00000532),
    .I3(sig0000052d),
    .O(sig0000042b)
  );
  LUT4 #(
    .INIT ( 16'hC3AA ))
  blk00000a85 (
    .I0(sig00000201),
    .I1(sig000001f0),
    .I2(sig00000532),
    .I3(sig0000052d),
    .O(sig0000042c)
  );
  LUT4 #(
    .INIT ( 16'hC3AA ))
  blk00000a86 (
    .I0(sig000001ff),
    .I1(sig000001ee),
    .I2(sig00000532),
    .I3(sig0000052d),
    .O(sig0000042a)
  );
  LUT4 #(
    .INIT ( 16'hC3AA ))
  blk00000a87 (
    .I0(sig00000202),
    .I1(sig000001f1),
    .I2(sig00000532),
    .I3(sig0000052d),
    .O(sig0000042d)
  );
  LUT4 #(
    .INIT ( 16'hD782 ))
  blk00000a88 (
    .I0(sig0000052d),
    .I1(sig000001f2),
    .I2(sig00000532),
    .I3(sig00000203),
    .O(sig0000042e)
  );
  LUT2 #(
    .INIT ( 4'h8 ))
  blk00000a89 (
    .I0(sig0000052d),
    .I1(sig00000532),
    .O(sig000003f9)
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  blk00000a8a (
    .I0(sig0000052d),
    .I1(sig00000532),
    .O(sig0000042f)
  );
  LUT2 #(
    .INIT ( 4'h8 ))
  blk00000a8b (
    .I0(sig000001d9),
    .I1(sig000001d8),
    .O(sig00000454)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000a8c (
    .I0(sig000004f7),
    .I1(sig000004c1),
    .O(sig0000059e)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000a8d (
    .I0(sig00000501),
    .I1(sig000004cb),
    .O(sig00000593)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000a8e (
    .I0(sig00000502),
    .I1(sig000004cc),
    .O(sig00000592)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000a8f (
    .I0(sig00000503),
    .I1(sig000004cd),
    .O(sig00000591)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000a90 (
    .I0(sig00000504),
    .I1(sig000004ce),
    .O(sig00000590)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000a91 (
    .I0(sig00000505),
    .I1(sig000004cf),
    .O(sig0000058f)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000a92 (
    .I0(sig00000506),
    .I1(sig000004d0),
    .O(sig0000058e)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000a93 (
    .I0(sig00000507),
    .I1(sig000004d1),
    .O(sig0000058d)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000a94 (
    .I0(sig00000508),
    .I1(sig000004d2),
    .O(sig0000059d)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000a95 (
    .I0(sig000004f8),
    .I1(sig000004c2),
    .O(sig0000059c)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000a96 (
    .I0(sig000004f9),
    .I1(sig000004c3),
    .O(sig0000059b)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000a97 (
    .I0(sig000004fa),
    .I1(sig000004c4),
    .O(sig0000059a)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000a98 (
    .I0(sig000004fb),
    .I1(sig000004c5),
    .O(sig00000599)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000a99 (
    .I0(sig000004fc),
    .I1(sig000004c6),
    .O(sig00000598)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000a9a (
    .I0(sig000004fd),
    .I1(sig000004c7),
    .O(sig00000597)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000a9b (
    .I0(sig000004fe),
    .I1(sig000004c8),
    .O(sig00000596)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000a9c (
    .I0(sig000004ff),
    .I1(sig000004c9),
    .O(sig00000595)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000a9d (
    .I0(sig00000500),
    .I1(sig000004ca),
    .O(sig00000594)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000a9e (
    .I0(sig000004f7),
    .I1(sig000004c1),
    .O(sig000005d3)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000a9f (
    .I0(sig00000501),
    .I1(sig000004cb),
    .O(sig000005c8)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000aa0 (
    .I0(sig00000502),
    .I1(sig000004cc),
    .O(sig000005c7)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000aa1 (
    .I0(sig00000503),
    .I1(sig000004cd),
    .O(sig000005c6)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000aa2 (
    .I0(sig00000504),
    .I1(sig000004ce),
    .O(sig000005c5)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000aa3 (
    .I0(sig00000505),
    .I1(sig000004cf),
    .O(sig000005c4)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000aa4 (
    .I0(sig00000506),
    .I1(sig000004d0),
    .O(sig000005c3)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000aa5 (
    .I0(sig00000507),
    .I1(sig000004d1),
    .O(sig000005c2)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000aa6 (
    .I0(sig00000508),
    .I1(sig000004d2),
    .O(sig000005d2)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000aa7 (
    .I0(sig000004f8),
    .I1(sig000004c2),
    .O(sig000005d1)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000aa8 (
    .I0(sig000004f9),
    .I1(sig000004c3),
    .O(sig000005d0)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000aa9 (
    .I0(sig000004fa),
    .I1(sig000004c4),
    .O(sig000005cf)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000aaa (
    .I0(sig000004fb),
    .I1(sig000004c5),
    .O(sig000005ce)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000aab (
    .I0(sig000004fc),
    .I1(sig000004c6),
    .O(sig000005cd)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000aac (
    .I0(sig000004fd),
    .I1(sig000004c7),
    .O(sig000005cc)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000aad (
    .I0(sig000004fe),
    .I1(sig000004c8),
    .O(sig000005cb)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000aae (
    .I0(sig000004ff),
    .I1(sig000004c9),
    .O(sig000005ca)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000aaf (
    .I0(sig00000500),
    .I1(sig000004ca),
    .O(sig000005c9)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000ab0 (
    .I0(sig000001b2),
    .I1(sig000001b3),
    .O(sig000005f7)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk00000ab1 (
    .I0(sig0000009d),
    .I1(sig0000009c),
    .I2(sig0000088f),
    .O(sig00000867)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000ab2 (
    .I0(sig000009aa),
    .I1(sig000009cd),
    .O(sig000008d1)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000ab3 (
    .I0(sig000009a9),
    .I1(sig000009cc),
    .O(sig000008d0)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000ab4 (
    .I0(sig000009a8),
    .I1(sig000009cb),
    .O(sig000008cf)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000ab5 (
    .I0(sig000009a7),
    .I1(sig000009ca),
    .O(sig000008ce)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000ab6 (
    .I0(sig000009a6),
    .I1(sig000009c9),
    .O(sig000008cd)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000ab7 (
    .I0(sig000009a5),
    .I1(sig000009c8),
    .O(sig000008cc)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000ab8 (
    .I0(sig000009a4),
    .I1(sig000009c7),
    .O(sig000008cb)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000ab9 (
    .I0(sig000009a3),
    .I1(sig000009c6),
    .O(sig000008ca)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000aba (
    .I0(sig000009a2),
    .I1(sig000009c5),
    .O(sig000008c9)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000abb (
    .I0(sig000009b0),
    .I1(sig000009d3),
    .O(sig000008c8)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000abc (
    .I0(sig000009b0),
    .I1(sig000009d3),
    .O(sig000008d7)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000abd (
    .I0(sig000009af),
    .I1(sig000009d2),
    .O(sig000008d6)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000abe (
    .I0(sig000009ae),
    .I1(sig000009d1),
    .O(sig000008d5)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000abf (
    .I0(sig000009ad),
    .I1(sig000009d0),
    .O(sig000008d4)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000ac0 (
    .I0(sig000009ac),
    .I1(sig000009cf),
    .O(sig000008d3)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000ac1 (
    .I0(sig000009ab),
    .I1(sig000009ce),
    .O(sig000008d2)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000ac2 (
    .I0(sig000009a1),
    .I1(sig000009c4),
    .O(sig000008c7)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000ac3 (
    .I0(sig000009aa),
    .I1(sig000009cd),
    .O(sig00000903)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000ac4 (
    .I0(sig000009a9),
    .I1(sig000009cc),
    .O(sig00000902)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000ac5 (
    .I0(sig000009a8),
    .I1(sig000009cb),
    .O(sig00000901)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000ac6 (
    .I0(sig000009a7),
    .I1(sig000009ca),
    .O(sig00000900)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000ac7 (
    .I0(sig000009a6),
    .I1(sig000009c9),
    .O(sig000008ff)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000ac8 (
    .I0(sig000009a5),
    .I1(sig000009c8),
    .O(sig000008fe)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000ac9 (
    .I0(sig000009a4),
    .I1(sig000009c7),
    .O(sig000008fd)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000aca (
    .I0(sig000009a3),
    .I1(sig000009c6),
    .O(sig000008fc)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000acb (
    .I0(sig000009a2),
    .I1(sig000009c5),
    .O(sig000008fb)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000acc (
    .I0(sig000009b0),
    .I1(sig000009d3),
    .O(sig000008fa)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000acd (
    .I0(sig000009b0),
    .I1(sig000009d3),
    .O(sig00000909)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000ace (
    .I0(sig000009af),
    .I1(sig000009d2),
    .O(sig00000908)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000acf (
    .I0(sig000009ae),
    .I1(sig000009d1),
    .O(sig00000907)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000ad0 (
    .I0(sig000009ad),
    .I1(sig000009d0),
    .O(sig00000906)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000ad1 (
    .I0(sig000009ac),
    .I1(sig000009cf),
    .O(sig00000905)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000ad2 (
    .I0(sig000009ab),
    .I1(sig000009ce),
    .O(sig00000904)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000ad3 (
    .I0(sig000009a1),
    .I1(sig000009c4),
    .O(sig000008f9)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000ad4 (
    .I0(sig00000bf0),
    .I1(sig00000bba),
    .O(sig00000a41)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000ad5 (
    .I0(sig00000bef),
    .I1(sig00000bb9),
    .O(sig00000a40)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000ad6 (
    .I0(sig00000bee),
    .I1(sig00000bb8),
    .O(sig00000a3f)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000ad7 (
    .I0(sig00000bed),
    .I1(sig00000bb7),
    .O(sig00000a3e)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000ad8 (
    .I0(sig00000bec),
    .I1(sig00000bb6),
    .O(sig00000a3d)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000ad9 (
    .I0(sig00000beb),
    .I1(sig00000bb5),
    .O(sig00000a3c)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000ada (
    .I0(sig00000bea),
    .I1(sig00000bb4),
    .O(sig00000a3b)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000adb (
    .I0(sig00000be9),
    .I1(sig00000bb3),
    .O(sig00000a3a)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000adc (
    .I0(sig00000be8),
    .I1(sig00000bb2),
    .O(sig00000a39)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000add (
    .I0(sig00000bf8),
    .I1(sig00000bc2),
    .O(sig00000a38)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000ade (
    .I0(sig00000bf7),
    .I1(sig00000bc1),
    .O(sig00000a48)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000adf (
    .I0(sig00000bf6),
    .I1(sig00000bc0),
    .O(sig00000a47)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000ae0 (
    .I0(sig00000bf5),
    .I1(sig00000bbf),
    .O(sig00000a46)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000ae1 (
    .I0(sig00000bf4),
    .I1(sig00000bbe),
    .O(sig00000a45)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000ae2 (
    .I0(sig00000bf3),
    .I1(sig00000bbd),
    .O(sig00000a44)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000ae3 (
    .I0(sig00000bf2),
    .I1(sig00000bbc),
    .O(sig00000a43)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000ae4 (
    .I0(sig00000bf1),
    .I1(sig00000bbb),
    .O(sig00000a42)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000ae5 (
    .I0(sig00000be7),
    .I1(sig00000bb1),
    .O(sig00000a37)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000ae6 (
    .I0(sig00000bf0),
    .I1(sig00000bba),
    .O(sig00000a76)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000ae7 (
    .I0(sig00000bef),
    .I1(sig00000bb9),
    .O(sig00000a75)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000ae8 (
    .I0(sig00000bee),
    .I1(sig00000bb8),
    .O(sig00000a74)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000ae9 (
    .I0(sig00000bed),
    .I1(sig00000bb7),
    .O(sig00000a73)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000aea (
    .I0(sig00000bec),
    .I1(sig00000bb6),
    .O(sig00000a72)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000aeb (
    .I0(sig00000beb),
    .I1(sig00000bb5),
    .O(sig00000a71)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000aec (
    .I0(sig00000bea),
    .I1(sig00000bb4),
    .O(sig00000a70)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000aed (
    .I0(sig00000be9),
    .I1(sig00000bb3),
    .O(sig00000a6f)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000aee (
    .I0(sig00000be8),
    .I1(sig00000bb2),
    .O(sig00000a6e)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000aef (
    .I0(sig00000bf8),
    .I1(sig00000bc2),
    .O(sig00000a6d)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000af0 (
    .I0(sig00000bf7),
    .I1(sig00000bc1),
    .O(sig00000a7d)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000af1 (
    .I0(sig00000bf6),
    .I1(sig00000bc0),
    .O(sig00000a7c)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000af2 (
    .I0(sig00000bf5),
    .I1(sig00000bbf),
    .O(sig00000a7b)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000af3 (
    .I0(sig00000bf4),
    .I1(sig00000bbe),
    .O(sig00000a7a)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000af4 (
    .I0(sig00000bf3),
    .I1(sig00000bbd),
    .O(sig00000a79)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000af5 (
    .I0(sig00000bf2),
    .I1(sig00000bbc),
    .O(sig00000a78)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000af6 (
    .I0(sig00000bf1),
    .I1(sig00000bbb),
    .O(sig00000a77)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000af7 (
    .I0(sig00000be7),
    .I1(sig00000bb1),
    .O(sig00000a6c)
  );
  LUT4 #(
    .INIT ( 16'h3CAA ))
  blk00000af8 (
    .I0(sig00000895),
    .I1(sig000008a6),
    .I2(sig00000c22),
    .I3(sig00000c1d),
    .O(sig00000ad8)
  );
  LUT4 #(
    .INIT ( 16'h3CAA ))
  blk00000af9 (
    .I0(sig00000896),
    .I1(sig000008a7),
    .I2(sig00000c22),
    .I3(sig00000c1d),
    .O(sig00000ad9)
  );
  LUT4 #(
    .INIT ( 16'h3CAA ))
  blk00000afa (
    .I0(sig00000897),
    .I1(sig000008a8),
    .I2(sig00000c22),
    .I3(sig00000c1d),
    .O(sig00000ada)
  );
  LUT4 #(
    .INIT ( 16'h3CAA ))
  blk00000afb (
    .I0(sig00000899),
    .I1(sig000008aa),
    .I2(sig00000c22),
    .I3(sig00000c1d),
    .O(sig00000adc)
  );
  LUT4 #(
    .INIT ( 16'h3CAA ))
  blk00000afc (
    .I0(sig0000089a),
    .I1(sig000008ab),
    .I2(sig00000c22),
    .I3(sig00000c1d),
    .O(sig00000add)
  );
  LUT4 #(
    .INIT ( 16'h3CAA ))
  blk00000afd (
    .I0(sig00000898),
    .I1(sig000008a9),
    .I2(sig00000c22),
    .I3(sig00000c1d),
    .O(sig00000adb)
  );
  LUT4 #(
    .INIT ( 16'h3CAA ))
  blk00000afe (
    .I0(sig0000089b),
    .I1(sig000008ac),
    .I2(sig00000c22),
    .I3(sig00000c1d),
    .O(sig00000ade)
  );
  LUT4 #(
    .INIT ( 16'h3CAA ))
  blk00000aff (
    .I0(sig0000089c),
    .I1(sig000008ad),
    .I2(sig00000c22),
    .I3(sig00000c1d),
    .O(sig00000adf)
  );
  LUT4 #(
    .INIT ( 16'h3CAA ))
  blk00000b00 (
    .I0(sig0000089d),
    .I1(sig000008ae),
    .I2(sig00000c22),
    .I3(sig00000c1d),
    .O(sig00000ae0)
  );
  LUT4 #(
    .INIT ( 16'h3CAA ))
  blk00000b01 (
    .I0(sig0000089e),
    .I1(sig000008af),
    .I2(sig00000c22),
    .I3(sig00000c1d),
    .O(sig00000ae1)
  );
  LUT4 #(
    .INIT ( 16'h3CAA ))
  blk00000b02 (
    .I0(sig000008a0),
    .I1(sig000008b1),
    .I2(sig00000c22),
    .I3(sig00000c1d),
    .O(sig00000ae3)
  );
  LUT4 #(
    .INIT ( 16'h3CAA ))
  blk00000b03 (
    .I0(sig000008a1),
    .I1(sig000008b2),
    .I2(sig00000c22),
    .I3(sig00000c1d),
    .O(sig00000ae4)
  );
  LUT4 #(
    .INIT ( 16'h3CAA ))
  blk00000b04 (
    .I0(sig0000089f),
    .I1(sig000008b0),
    .I2(sig00000c22),
    .I3(sig00000c1d),
    .O(sig00000ae2)
  );
  LUT4 #(
    .INIT ( 16'h3CAA ))
  blk00000b05 (
    .I0(sig000008a2),
    .I1(sig000008b3),
    .I2(sig00000c22),
    .I3(sig00000c1d),
    .O(sig00000ae5)
  );
  LUT4 #(
    .INIT ( 16'h3CAA ))
  blk00000b06 (
    .I0(sig000008a3),
    .I1(sig000008b4),
    .I2(sig00000c22),
    .I3(sig00000c1d),
    .O(sig00000ae6)
  );
  LUT4 #(
    .INIT ( 16'h3CAA ))
  blk00000b07 (
    .I0(sig000008a4),
    .I1(sig000008b5),
    .I2(sig00000c22),
    .I3(sig00000c1d),
    .O(sig00000ae7)
  );
  LUT4 #(
    .INIT ( 16'h7D28 ))
  blk00000b08 (
    .I0(sig00000c1d),
    .I1(sig000008b6),
    .I2(sig00000c22),
    .I3(sig000008a5),
    .O(sig00000ae8)
  );
  LUT4 #(
    .INIT ( 16'hC3AA ))
  blk00000b09 (
    .I0(sig000008a6),
    .I1(sig00000895),
    .I2(sig00000c22),
    .I3(sig00000c1d),
    .O(sig00000b0e)
  );
  LUT4 #(
    .INIT ( 16'hC3AA ))
  blk00000b0a (
    .I0(sig000008a7),
    .I1(sig00000896),
    .I2(sig00000c22),
    .I3(sig00000c1d),
    .O(sig00000b0f)
  );
  LUT4 #(
    .INIT ( 16'hC3AA ))
  blk00000b0b (
    .I0(sig000008a8),
    .I1(sig00000897),
    .I2(sig00000c22),
    .I3(sig00000c1d),
    .O(sig00000b10)
  );
  LUT4 #(
    .INIT ( 16'hC3AA ))
  blk00000b0c (
    .I0(sig000008a9),
    .I1(sig00000898),
    .I2(sig00000c22),
    .I3(sig00000c1d),
    .O(sig00000b11)
  );
  LUT4 #(
    .INIT ( 16'hC3AA ))
  blk00000b0d (
    .I0(sig000008ab),
    .I1(sig0000089a),
    .I2(sig00000c22),
    .I3(sig00000c1d),
    .O(sig00000b13)
  );
  LUT4 #(
    .INIT ( 16'hC3AA ))
  blk00000b0e (
    .I0(sig000008ac),
    .I1(sig0000089b),
    .I2(sig00000c22),
    .I3(sig00000c1d),
    .O(sig00000b14)
  );
  LUT4 #(
    .INIT ( 16'hC3AA ))
  blk00000b0f (
    .I0(sig000008aa),
    .I1(sig00000899),
    .I2(sig00000c22),
    .I3(sig00000c1d),
    .O(sig00000b12)
  );
  LUT4 #(
    .INIT ( 16'hC3AA ))
  blk00000b10 (
    .I0(sig000008ad),
    .I1(sig0000089c),
    .I2(sig00000c22),
    .I3(sig00000c1d),
    .O(sig00000b15)
  );
  LUT4 #(
    .INIT ( 16'hC3AA ))
  blk00000b11 (
    .I0(sig000008ae),
    .I1(sig0000089d),
    .I2(sig00000c22),
    .I3(sig00000c1d),
    .O(sig00000b16)
  );
  LUT4 #(
    .INIT ( 16'hC3AA ))
  blk00000b12 (
    .I0(sig000008af),
    .I1(sig0000089e),
    .I2(sig00000c22),
    .I3(sig00000c1d),
    .O(sig00000b17)
  );
  LUT4 #(
    .INIT ( 16'hC3AA ))
  blk00000b13 (
    .I0(sig000008b0),
    .I1(sig0000089f),
    .I2(sig00000c22),
    .I3(sig00000c1d),
    .O(sig00000b18)
  );
  LUT4 #(
    .INIT ( 16'hC3AA ))
  blk00000b14 (
    .I0(sig000008b2),
    .I1(sig000008a1),
    .I2(sig00000c22),
    .I3(sig00000c1d),
    .O(sig00000b1a)
  );
  LUT4 #(
    .INIT ( 16'hC3AA ))
  blk00000b15 (
    .I0(sig000008b3),
    .I1(sig000008a2),
    .I2(sig00000c22),
    .I3(sig00000c1d),
    .O(sig00000b1b)
  );
  LUT4 #(
    .INIT ( 16'hC3AA ))
  blk00000b16 (
    .I0(sig000008b1),
    .I1(sig000008a0),
    .I2(sig00000c22),
    .I3(sig00000c1d),
    .O(sig00000b19)
  );
  LUT4 #(
    .INIT ( 16'hC3AA ))
  blk00000b17 (
    .I0(sig000008b4),
    .I1(sig000008a3),
    .I2(sig00000c22),
    .I3(sig00000c1d),
    .O(sig00000b1c)
  );
  LUT4 #(
    .INIT ( 16'hC3AA ))
  blk00000b18 (
    .I0(sig000008b5),
    .I1(sig000008a4),
    .I2(sig00000c22),
    .I3(sig00000c1d),
    .O(sig00000b1d)
  );
  LUT4 #(
    .INIT ( 16'hD782 ))
  blk00000b19 (
    .I0(sig00000c1d),
    .I1(sig000008a5),
    .I2(sig00000c22),
    .I3(sig000008b6),
    .O(sig00000b1e)
  );
  LUT2 #(
    .INIT ( 4'h8 ))
  blk00000b1a (
    .I0(sig00000c1d),
    .I1(sig00000c22),
    .O(sig00000ae9)
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  blk00000b1b (
    .I0(sig00000c1d),
    .I1(sig00000c22),
    .O(sig00000b1f)
  );
  LUT2 #(
    .INIT ( 4'h8 ))
  blk00000b1c (
    .I0(sig00000894),
    .I1(sig00000893),
    .O(sig00000b44)
  );
  FDSE #(
    .INIT ( 1'b0 ))
  blk00000b1d (
    .C(aclk),
    .CE(sig00000001),
    .D(sig00000055),
    .S(sig0000005c),
    .Q(sig00000064)
  );
  FDSE #(
    .INIT ( 1'b0 ))
  blk00000b1e (
    .C(aclk),
    .CE(sig00000001),
    .D(sig00000056),
    .S(sig0000005c),
    .Q(sig00000063)
  );
  FDSE #(
    .INIT ( 1'b0 ))
  blk00000b1f (
    .C(aclk),
    .CE(sig00000001),
    .D(sig00000057),
    .S(sig0000005c),
    .Q(sig00000062)
  );
  FDSE #(
    .INIT ( 1'b0 ))
  blk00000b20 (
    .C(aclk),
    .CE(sig00000001),
    .D(sig00000058),
    .S(sig0000005c),
    .Q(sig00000053)
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  blk00000b21 (
    .I0(sig00000029),
    .I1(sig00000121),
    .O(sig00000c4f)
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  blk00000b22 (
    .I0(sig00000028),
    .I1(sig00000121),
    .O(sig00000c50)
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  blk00000b23 (
    .I0(sig00000027),
    .I1(sig00000121),
    .O(sig00000c51)
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  blk00000b24 (
    .I0(sig000000c6),
    .I1(sig00000072),
    .O(sig00000c52)
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  blk00000b25 (
    .I0(sig000000c7),
    .I1(sig00000072),
    .O(sig00000c53)
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  blk00000b26 (
    .I0(sig000000c8),
    .I1(sig00000072),
    .O(sig00000c54)
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  blk00000b27 (
    .I0(sig00000205),
    .I1(sig00000150),
    .O(sig00000c55)
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  blk00000b28 (
    .I0(sig00000206),
    .I1(sig00000150),
    .O(sig00000c56)
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  blk00000b29 (
    .I0(sig00000207),
    .I1(sig00000150),
    .O(sig00000c57)
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  blk00000b2a (
    .I0(sig00000151),
    .O(sig00000c58)
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  blk00000b2b (
    .I0(sig0000020a),
    .I1(sig00000229),
    .O(sig00000c59)
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  blk00000b2c (
    .I0(sig0000020b),
    .I1(sig00000229),
    .O(sig00000c5a)
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  blk00000b2d (
    .I0(sig0000020c),
    .I1(sig00000229),
    .O(sig00000c5b)
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  blk00000b2e (
    .I0(sig00000228),
    .O(sig00000c5c)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000b2f (
    .I0(sig000002bf),
    .I1(sig000002e2),
    .O(sig00000c5d)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000b30 (
    .I0(sig000002bf),
    .I1(sig000002e2),
    .O(sig00000c5e)
  );
  LUT4 #(
    .INIT ( 16'h3CAA ))
  blk00000b31 (
    .I0(sig000001f2),
    .I1(sig00000203),
    .I2(sig00000532),
    .I3(sig0000052d),
    .O(sig00000c5f)
  );
  LUT4 #(
    .INIT ( 16'hC3AA ))
  blk00000b32 (
    .I0(sig00000203),
    .I1(sig000001f2),
    .I2(sig00000532),
    .I3(sig0000052d),
    .O(sig00000c60)
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  blk00000b33 (
    .I0(sig000001b3),
    .O(sig00000c61)
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  blk00000b34 (
    .I0(sig000001b2),
    .O(sig00000c62)
  );
  LUT4 #(
    .INIT ( 16'h3CAA ))
  blk00000b35 (
    .I0(sig000008a5),
    .I1(sig000008b6),
    .I2(sig00000c22),
    .I3(sig00000c1d),
    .O(sig00000c63)
  );
  LUT4 #(
    .INIT ( 16'hC3AA ))
  blk00000b36 (
    .I0(sig000008b6),
    .I1(sig000008a5),
    .I2(sig00000c22),
    .I3(sig00000c1d),
    .O(sig00000c64)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000b37 (
    .C(aclk),
    .D(sig00000c65),
    .Q(sig0000006d)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000b38 (
    .C(aclk),
    .D(sig00000c66),
    .Q(sig0000006f)
  );
  LUT3 #(
    .INIT ( 8'hA2 ))
  blk00000b39 (
    .I0(s_axis_config_tvalid),
    .I1(sig0000006d),
    .I2(sig00000065),
    .O(sig0000006c)
  );
  LUT3 #(
    .INIT ( 8'hA2 ))
  blk00000b3a (
    .I0(s_axis_data_tvalid),
    .I1(sig0000006f),
    .I2(sig00000002),
    .O(sig0000006e)
  );
  LUT3 #(
    .INIT ( 8'h60 ))
  blk00000b3b (
    .I0(sig000005e7),
    .I1(sig000005e8),
    .I2(sig00000806),
    .O(sig000007f6)
  );
  LUT3 #(
    .INIT ( 8'h60 ))
  blk00000b3c (
    .I0(sig000005e6),
    .I1(sig000005e8),
    .I2(sig00000826),
    .O(sig00000816)
  );
  LUT4 #(
    .INIT ( 16'hF690 ))
  blk00000b3d (
    .I0(sig000005e8),
    .I1(sig000005e7),
    .I2(sig000001a0),
    .I3(sig00000805),
    .O(sig000007f5)
  );
  LUT4 #(
    .INIT ( 16'hF690 ))
  blk00000b3e (
    .I0(sig000005e8),
    .I1(sig000005e6),
    .I2(sig000001ae),
    .I3(sig00000825),
    .O(sig00000815)
  );
  LUT4 #(
    .INIT ( 16'hF690 ))
  blk00000b3f (
    .I0(sig000005e8),
    .I1(sig000005e7),
    .I2(sig00000193),
    .I3(sig00000804),
    .O(sig000007f4)
  );
  LUT4 #(
    .INIT ( 16'hF690 ))
  blk00000b40 (
    .I0(sig000005e8),
    .I1(sig000005e6),
    .I2(sig00000199),
    .I3(sig00000824),
    .O(sig00000814)
  );
  LUT4 #(
    .INIT ( 16'hF690 ))
  blk00000b41 (
    .I0(sig000005e8),
    .I1(sig000005e7),
    .I2(sig00000198),
    .I3(sig00000803),
    .O(sig000007f3)
  );
  LUT4 #(
    .INIT ( 16'hF690 ))
  blk00000b42 (
    .I0(sig000005e8),
    .I1(sig000005e6),
    .I2(sig00000198),
    .I3(sig00000823),
    .O(sig00000813)
  );
  LUT4 #(
    .INIT ( 16'hF690 ))
  blk00000b43 (
    .I0(sig000005e8),
    .I1(sig000005e7),
    .I2(sig0000019d),
    .I3(sig00000802),
    .O(sig000007f2)
  );
  LUT4 #(
    .INIT ( 16'hF690 ))
  blk00000b44 (
    .I0(sig000005e8),
    .I1(sig000005e6),
    .I2(sig0000019d),
    .I3(sig00000822),
    .O(sig00000812)
  );
  LUT4 #(
    .INIT ( 16'hF690 ))
  blk00000b45 (
    .I0(sig000005e8),
    .I1(sig000005e7),
    .I2(sig0000019c),
    .I3(sig00000801),
    .O(sig000007f1)
  );
  LUT4 #(
    .INIT ( 16'hF690 ))
  blk00000b46 (
    .I0(sig000005e8),
    .I1(sig000005e6),
    .I2(sig0000019c),
    .I3(sig00000821),
    .O(sig00000811)
  );
  LUT4 #(
    .INIT ( 16'hF690 ))
  blk00000b47 (
    .I0(sig000005e8),
    .I1(sig000005e7),
    .I2(sig0000019b),
    .I3(sig00000800),
    .O(sig000007f0)
  );
  LUT4 #(
    .INIT ( 16'hF690 ))
  blk00000b48 (
    .I0(sig000005e8),
    .I1(sig000005e6),
    .I2(sig00000194),
    .I3(sig00000820),
    .O(sig00000810)
  );
  LUT4 #(
    .INIT ( 16'hF690 ))
  blk00000b49 (
    .I0(sig000005e8),
    .I1(sig000005e7),
    .I2(sig00000193),
    .I3(sig000007ff),
    .O(sig000007ef)
  );
  LUT4 #(
    .INIT ( 16'hF690 ))
  blk00000b4a (
    .I0(sig000005e8),
    .I1(sig000005e6),
    .I2(sig00000199),
    .I3(sig0000081f),
    .O(sig0000080f)
  );
  LUT3 #(
    .INIT ( 8'h60 ))
  blk00000b4b (
    .I0(sig000005e7),
    .I1(sig000005e8),
    .I2(sig000007fe),
    .O(sig000007ee)
  );
  LUT3 #(
    .INIT ( 8'h60 ))
  blk00000b4c (
    .I0(sig000005e6),
    .I1(sig000005e8),
    .I2(sig0000081e),
    .O(sig0000080e)
  );
  LUT4 #(
    .INIT ( 16'hF690 ))
  blk00000b4d (
    .I0(sig000005e8),
    .I1(sig000005e7),
    .I2(sig00000199),
    .I3(sig000007fd),
    .O(sig000007ed)
  );
  LUT4 #(
    .INIT ( 16'hF690 ))
  blk00000b4e (
    .I0(sig000005e8),
    .I1(sig000005e6),
    .I2(sig00000193),
    .I3(sig0000081d),
    .O(sig0000080d)
  );
  LUT4 #(
    .INIT ( 16'hF690 ))
  blk00000b4f (
    .I0(sig000005e8),
    .I1(sig000005e7),
    .I2(sig00000198),
    .I3(sig000007fc),
    .O(sig000007ec)
  );
  LUT4 #(
    .INIT ( 16'hF690 ))
  blk00000b50 (
    .I0(sig000005e8),
    .I1(sig000005e6),
    .I2(sig00000198),
    .I3(sig0000081c),
    .O(sig0000080c)
  );
  LUT4 #(
    .INIT ( 16'hF690 ))
  blk00000b51 (
    .I0(sig000005e8),
    .I1(sig000005e7),
    .I2(sig00000194),
    .I3(sig000007fb),
    .O(sig000007eb)
  );
  LUT4 #(
    .INIT ( 16'hF690 ))
  blk00000b52 (
    .I0(sig000005e8),
    .I1(sig000005e6),
    .I2(sig0000019b),
    .I3(sig0000081b),
    .O(sig0000080b)
  );
  LUT4 #(
    .INIT ( 16'hF690 ))
  blk00000b53 (
    .I0(sig000005e8),
    .I1(sig000005e7),
    .I2(sig00000194),
    .I3(sig000007fa),
    .O(sig000007ea)
  );
  LUT4 #(
    .INIT ( 16'hF690 ))
  blk00000b54 (
    .I0(sig000005e8),
    .I1(sig000005e6),
    .I2(sig0000019b),
    .I3(sig0000081a),
    .O(sig0000080a)
  );
  LUT4 #(
    .INIT ( 16'hF690 ))
  blk00000b55 (
    .I0(sig000005e8),
    .I1(sig000005e7),
    .I2(sig00000194),
    .I3(sig000007f9),
    .O(sig000007e9)
  );
  LUT4 #(
    .INIT ( 16'hF690 ))
  blk00000b56 (
    .I0(sig000005e8),
    .I1(sig000005e6),
    .I2(sig0000019b),
    .I3(sig00000819),
    .O(sig00000809)
  );
  LUT4 #(
    .INIT ( 16'hF690 ))
  blk00000b57 (
    .I0(sig000005e8),
    .I1(sig000005e7),
    .I2(sig00000194),
    .I3(sig000007f8),
    .O(sig000007e8)
  );
  LUT4 #(
    .INIT ( 16'hF690 ))
  blk00000b58 (
    .I0(sig000005e8),
    .I1(sig000005e6),
    .I2(sig0000019b),
    .I3(sig00000818),
    .O(sig00000808)
  );
  LUT3 #(
    .INIT ( 8'hF2 ))
  blk00000b59 (
    .I0(sig0000006d),
    .I1(sig00000065),
    .I2(s_axis_config_tvalid),
    .O(sig00000c65)
  );
  LUT4 #(
    .INIT ( 16'hF690 ))
  blk00000b5a (
    .I0(sig000005e8),
    .I1(sig000005e7),
    .I2(sig00000193),
    .I3(sig000007f7),
    .O(sig000007e7)
  );
  LUT4 #(
    .INIT ( 16'hF690 ))
  blk00000b5b (
    .I0(sig000005e8),
    .I1(sig000005e6),
    .I2(sig00000199),
    .I3(sig00000817),
    .O(sig00000807)
  );
  LUT3 #(
    .INIT ( 8'hF2 ))
  blk00000b5c (
    .I0(sig0000006f),
    .I1(sig00000002),
    .I2(s_axis_data_tvalid),
    .O(sig00000c66)
  );
  LUT5 #(
    .INIT ( 32'h00800000 ))
  blk00000b5d (
    .I0(sig00000027),
    .I1(sig00000029),
    .I2(sig0000002a),
    .I3(sig0000006b),
    .I4(sig00000028),
    .O(sig0000005b)
  );
  LUT6 #(
    .INIT ( 64'h0888888888888888 ))
  blk00000b5e (
    .I0(sig00000002),
    .I1(sig0000006b),
    .I2(sig00000029),
    .I3(sig0000002a),
    .I4(sig00000027),
    .I5(sig00000028),
    .O(sig00000054)
  );
  LUT6 #(
    .INIT ( 64'h2222222222F22222 ))
  blk00000b5f (
    .I0(sig00000068),
    .I1(sig0000006f),
    .I2(sig00000066),
    .I3(sig00000052),
    .I4(sig00000002),
    .I5(s_axis_data_tvalid),
    .O(sig0000005a)
  );
  MUXF7   blk00000b60 (
    .I0(sig00000c67),
    .I1(sig00000c68),
    .S(sig00000052),
    .O(sig0000002d)
  );
  LUT6 #(
    .INIT ( 64'hFFFFDC54DC54DC54 ))
  blk00000b61 (
    .I0(sig00000002),
    .I1(sig00000066),
    .I2(sig00000067),
    .I3(s_axis_data_tvalid),
    .I4(sig0000006f),
    .I5(sig00000068),
    .O(sig00000c67)
  );
  LUT4 #(
    .INIT ( 16'h8F88 ))
  blk00000b62 (
    .I0(sig00000068),
    .I1(sig0000006f),
    .I2(sig00000002),
    .I3(sig00000067),
    .O(sig00000c68)
  );
  INV   blk00000b63 (
    .I(sig000001a0),
    .O(sig000007ae)
  );
  INV   blk00000b64 (
    .I(sig00000193),
    .O(sig000007b0)
  );
  INV   blk00000b65 (
    .I(sig00000198),
    .O(sig000007b2)
  );
  INV   blk00000b66 (
    .I(sig0000019d),
    .O(sig000007b4)
  );
  INV   blk00000b67 (
    .I(sig0000019c),
    .O(sig000007b6)
  );
  INV   blk00000b68 (
    .I(sig0000019b),
    .O(sig000007b8)
  );
  INV   blk00000b69 (
    .I(sig00000193),
    .O(sig000007ba)
  );
  INV   blk00000b6a (
    .I(sig00000199),
    .O(sig000007bd)
  );
  INV   blk00000b6b (
    .I(sig00000198),
    .O(sig000007bf)
  );
  INV   blk00000b6c (
    .I(sig00000194),
    .O(sig000007c1)
  );
  INV   blk00000b6d (
    .I(sig00000194),
    .O(sig000007c3)
  );
  INV   blk00000b6e (
    .I(sig00000194),
    .O(sig000007c5)
  );
  INV   blk00000b6f (
    .I(sig00000194),
    .O(sig000007c7)
  );
  INV   blk00000b70 (
    .I(sig00000193),
    .O(sig000007c9)
  );
  INV   blk00000b71 (
    .I(sig000001ae),
    .O(sig000007cb)
  );
  INV   blk00000b72 (
    .I(sig00000199),
    .O(sig000007cd)
  );
  INV   blk00000b73 (
    .I(sig00000198),
    .O(sig000007cf)
  );
  INV   blk00000b74 (
    .I(sig0000019d),
    .O(sig000007d1)
  );
  INV   blk00000b75 (
    .I(sig0000019c),
    .O(sig000007d3)
  );
  INV   blk00000b76 (
    .I(sig00000194),
    .O(sig000007d5)
  );
  INV   blk00000b77 (
    .I(sig00000199),
    .O(sig000007d7)
  );
  INV   blk00000b78 (
    .I(sig00000193),
    .O(sig000007da)
  );
  INV   blk00000b79 (
    .I(sig00000198),
    .O(sig000007dc)
  );
  INV   blk00000b7a (
    .I(sig0000019b),
    .O(sig000007de)
  );
  INV   blk00000b7b (
    .I(sig0000019b),
    .O(sig000007e0)
  );
  INV   blk00000b7c (
    .I(sig0000019b),
    .O(sig000007e2)
  );
  INV   blk00000b7d (
    .I(sig0000019b),
    .O(sig000007e4)
  );
  INV   blk00000b7e (
    .I(sig00000199),
    .O(sig000007e6)
  );
  INV   blk00000b7f (
    .I(sig00000053),
    .O(sig00000058)
  );
  INV   blk00000b80 (
    .I(sig00000072),
    .O(sig00000075)
  );
  INV   blk00000b81 (
    .I(sig00000121),
    .O(sig00000119)
  );
  INV   blk00000b82 (
    .I(sig00000150),
    .O(sig00000157)
  );
  INV   blk00000b83 (
    .I(sig00000229),
    .O(sig00000222)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000b84 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig0000076a),
    .Q(sig00000c69),
    .Q15(NLW_blk00000b84_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000b85 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000c69),
    .Q(sig0000074a)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000b86 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000001af),
    .Q(sig00000c6a),
    .Q15(NLW_blk00000b86_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000b87 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000c6a),
    .Q(sig000005e5)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000b88 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000769),
    .Q(sig00000c6b),
    .Q15(NLW_blk00000b88_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000b89 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000c6b),
    .Q(sig00000749)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000b8a (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig0000076b),
    .Q(sig00000c6c),
    .Q15(NLW_blk00000b8a_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000b8b (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000c6c),
    .Q(sig0000074b)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000b8c (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig0000076c),
    .Q(sig00000c6d),
    .Q15(NLW_blk00000b8c_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000b8d (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000c6d),
    .Q(sig0000074c)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000b8e (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig0000076d),
    .Q(sig00000c6e),
    .Q15(NLW_blk00000b8e_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000b8f (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000c6e),
    .Q(sig0000074d)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000b90 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig0000076e),
    .Q(sig00000c6f),
    .Q15(NLW_blk00000b90_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000b91 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000c6f),
    .Q(sig0000074e)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000b92 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig0000076f),
    .Q(sig00000c70),
    .Q15(NLW_blk00000b92_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000b93 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000c70),
    .Q(sig0000074f)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000b94 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000770),
    .Q(sig00000c71),
    .Q15(NLW_blk00000b94_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000b95 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000c71),
    .Q(sig00000750)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000b96 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000773),
    .Q(sig00000c72),
    .Q15(NLW_blk00000b96_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000b97 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000c72),
    .Q(sig00000753)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000b98 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000771),
    .Q(sig00000c73),
    .Q15(NLW_blk00000b98_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000b99 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000c73),
    .Q(sig00000751)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000b9a (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000772),
    .Q(sig00000c74),
    .Q15(NLW_blk00000b9a_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000b9b (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000c74),
    .Q(sig00000752)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000b9c (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000774),
    .Q(sig00000c75),
    .Q15(NLW_blk00000b9c_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000b9d (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000c75),
    .Q(sig00000754)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000b9e (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000775),
    .Q(sig00000c76),
    .Q15(NLW_blk00000b9e_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000b9f (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000c76),
    .Q(sig00000755)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000ba0 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000776),
    .Q(sig00000c77),
    .Q15(NLW_blk00000ba0_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000ba1 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000c77),
    .Q(sig00000756)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000ba2 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000777),
    .Q(sig00000c78),
    .Q15(NLW_blk00000ba2_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000ba3 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000c78),
    .Q(sig00000757)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000ba4 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000778),
    .Q(sig00000c79),
    .Q15(NLW_blk00000ba4_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000ba5 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000c79),
    .Q(sig00000758)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000ba6 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000680),
    .Q(sig00000c7a),
    .Q15(NLW_blk00000ba6_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000ba7 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000c7a),
    .Q(sig00000643)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000ba8 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig0000068a),
    .Q(sig00000c7b),
    .Q15(NLW_blk00000ba8_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000ba9 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000c7b),
    .Q(sig00000646)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000baa (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000688),
    .Q(sig00000c7c),
    .Q15(NLW_blk00000baa_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000bab (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000c7c),
    .Q(sig00000644)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000bac (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000689),
    .Q(sig00000c7d),
    .Q15(NLW_blk00000bac_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000bad (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000c7d),
    .Q(sig00000645)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000bae (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig0000068b),
    .Q(sig00000c7e),
    .Q15(NLW_blk00000bae_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000baf (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000c7e),
    .Q(sig00000647)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000bb0 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig0000068c),
    .Q(sig00000c7f),
    .Q15(NLW_blk00000bb0_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000bb1 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000c7f),
    .Q(sig00000648)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000bb2 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig0000068d),
    .Q(sig00000c80),
    .Q15(NLW_blk00000bb2_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000bb3 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000c80),
    .Q(sig00000649)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000bb4 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig0000068e),
    .Q(sig00000c81),
    .Q15(NLW_blk00000bb4_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000bb5 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000c81),
    .Q(sig0000064a)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000bb6 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig0000068f),
    .Q(sig00000c82),
    .Q15(NLW_blk00000bb6_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000bb7 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000c82),
    .Q(sig0000064b)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000bb8 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000690),
    .Q(sig00000c83),
    .Q15(NLW_blk00000bb8_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000bb9 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000c83),
    .Q(sig0000064c)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000bba (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000691),
    .Q(sig00000c84),
    .Q15(NLW_blk00000bba_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000bbb (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000c84),
    .Q(sig0000064d)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000bbc (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000692),
    .Q(sig00000c85),
    .Q15(NLW_blk00000bbc_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000bbd (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000c85),
    .Q(sig0000064e)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000bbe (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000693),
    .Q(sig00000c86),
    .Q15(NLW_blk00000bbe_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000bbf (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000c86),
    .Q(sig0000064f)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000bc0 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000694),
    .Q(sig00000c87),
    .Q15(NLW_blk00000bc0_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000bc1 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000c87),
    .Q(sig00000650)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000bc2 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000695),
    .Q(sig00000c88),
    .Q15(NLW_blk00000bc2_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000bc3 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000c88),
    .Q(sig00000651)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000bc4 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000696),
    .Q(sig00000c89),
    .Q15(NLW_blk00000bc4_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000bc5 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000c89),
    .Q(sig00000652)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000bc6 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000697),
    .Q(sig00000c8a),
    .Q15(NLW_blk00000bc6_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000bc7 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000c8a),
    .Q(sig00000653)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000bc8 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000698),
    .Q(sig00000c8b),
    .Q15(NLW_blk00000bc8_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000bc9 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000c8b),
    .Q(sig00000654)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000bca (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig0000069c),
    .Q(sig00000c8c),
    .Q15(NLW_blk00000bca_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000bcb (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000c8c),
    .Q(sig00000634)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000bcc (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000699),
    .Q(sig00000c8d),
    .Q15(NLW_blk00000bcc_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000bcd (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000c8d),
    .Q(sig0000062a)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000bce (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig0000069b),
    .Q(sig00000c8e),
    .Q15(NLW_blk00000bce_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000bcf (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000c8e),
    .Q(sig00000633)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000bd0 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig0000069d),
    .Q(sig00000c8f),
    .Q15(NLW_blk00000bd0_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000bd1 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000c8f),
    .Q(sig00000635)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000bd2 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig0000069e),
    .Q(sig00000c90),
    .Q15(NLW_blk00000bd2_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000bd3 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000c90),
    .Q(sig00000636)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000bd4 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig0000069f),
    .Q(sig00000c91),
    .Q15(NLW_blk00000bd4_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000bd5 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000c91),
    .Q(sig00000637)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000bd6 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000006a0),
    .Q(sig00000c92),
    .Q15(NLW_blk00000bd6_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000bd7 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000c92),
    .Q(sig00000638)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000bd8 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000006a1),
    .Q(sig00000c93),
    .Q15(NLW_blk00000bd8_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000bd9 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000c93),
    .Q(sig00000639)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000bda (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000006a2),
    .Q(sig00000c94),
    .Q15(NLW_blk00000bda_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000bdb (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000c94),
    .Q(sig0000063a)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000bdc (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000006a3),
    .Q(sig00000c95),
    .Q15(NLW_blk00000bdc_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000bdd (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000c95),
    .Q(sig0000063b)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000bde (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000006a4),
    .Q(sig00000c96),
    .Q15(NLW_blk00000bde_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000bdf (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000c96),
    .Q(sig0000063c)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000be0 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000006a5),
    .Q(sig00000c97),
    .Q15(NLW_blk00000be0_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000be1 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000c97),
    .Q(sig0000063d)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000be2 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000006a6),
    .Q(sig00000c98),
    .Q15(NLW_blk00000be2_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000be3 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000c98),
    .Q(sig0000063e)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000be4 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000006a7),
    .Q(sig00000c99),
    .Q15(NLW_blk00000be4_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000be5 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000c99),
    .Q(sig0000063f)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000be6 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000006a8),
    .Q(sig00000c9a),
    .Q15(NLW_blk00000be6_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000be7 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000c9a),
    .Q(sig00000640)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000be8 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000006a9),
    .Q(sig00000c9b),
    .Q15(NLW_blk00000be8_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000be9 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000c9b),
    .Q(sig00000641)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000bea (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig0000079a),
    .Q(sig00000c9c),
    .Q15(NLW_blk00000bea_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000beb (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000c9c),
    .Q(sig000006ef)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000bec (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000797),
    .Q(sig00000c9d),
    .Q15(NLW_blk00000bec_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000bed (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000c9d),
    .Q(sig000006f2)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000bee (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000799),
    .Q(sig00000c9e),
    .Q15(NLW_blk00000bee_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000bef (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000c9e),
    .Q(sig000006f0)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000bf0 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000798),
    .Q(sig00000c9f),
    .Q15(NLW_blk00000bf0_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000bf1 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000c9f),
    .Q(sig000006f1)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000bf2 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000796),
    .Q(sig00000ca0),
    .Q15(NLW_blk00000bf2_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000bf3 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000ca0),
    .Q(sig000006f3)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000bf4 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000795),
    .Q(sig00000ca1),
    .Q15(NLW_blk00000bf4_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000bf5 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000ca1),
    .Q(sig000006f4)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000bf6 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000794),
    .Q(sig00000ca2),
    .Q15(NLW_blk00000bf6_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000bf7 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000ca2),
    .Q(sig000006f5)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000bf8 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000793),
    .Q(sig00000ca3),
    .Q15(NLW_blk00000bf8_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000bf9 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000ca3),
    .Q(sig000006f6)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000bfa (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000792),
    .Q(sig00000ca4),
    .Q15(NLW_blk00000bfa_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000bfb (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000ca4),
    .Q(sig000006f7)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000bfc (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000791),
    .Q(sig00000ca5),
    .Q15(NLW_blk00000bfc_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000bfd (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000ca5),
    .Q(sig000006f8)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000bfe (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000790),
    .Q(sig00000ca6),
    .Q15(NLW_blk00000bfe_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000bff (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000ca6),
    .Q(sig000006f9)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000c00 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig0000078f),
    .Q(sig00000ca7),
    .Q15(NLW_blk00000c00_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000c01 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000ca7),
    .Q(sig000006fa)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000c02 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig0000078e),
    .Q(sig00000ca8),
    .Q15(NLW_blk00000c02_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000c03 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000ca8),
    .Q(sig000006fb)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000c04 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig0000078d),
    .Q(sig00000ca9),
    .Q15(NLW_blk00000c04_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000c05 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000ca9),
    .Q(sig000006fc)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000c06 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig0000078c),
    .Q(sig00000caa),
    .Q15(NLW_blk00000c06_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000c07 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000caa),
    .Q(sig000006fd)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000c08 (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig0000078b),
    .Q(sig00000cab),
    .Q15(NLW_blk00000c08_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000c09 (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000cab),
    .Q(sig000006fe)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000c0a (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig0000078a),
    .Q(sig00000cac),
    .Q15(NLW_blk00000c0a_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000c0b (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000cac),
    .Q(sig000006ff)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000c0c (
    .A0(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A1(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A2(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .A3(\NlwRenamedSig_OI_U0/i_synth/axi_wrapper/blk_event_tlast_unexpected.events_to_transfer [1]),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000789),
    .Q(sig00000cad),
    .Q15(NLW_blk00000c0c_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000c0d (
    .C(aclk),
    .CE(sig00000344),
    .D(sig00000cad),
    .Q(sig00000700)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000000dc/blk000000e0  (
    .C(aclk),
    .CE(sig00000344),
    .D(\blk000000dc/sig00000cb4 ),
    .Q(sig00000120)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk000000dc/blk000000df  (
    .A0(\blk000000dc/sig00000cb3 ),
    .A1(\blk000000dc/sig00000cb2 ),
    .A2(\blk000000dc/sig00000cb2 ),
    .A3(\blk000000dc/sig00000cb2 ),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig0000011f),
    .Q(\blk000000dc/sig00000cb4 ),
    .Q15(\NLW_blk000000dc/blk000000df_Q15_UNCONNECTED )
  );
  VCC   \blk000000dc/blk000000de  (
    .P(\blk000000dc/sig00000cb3 )
  );
  GND   \blk000000dc/blk000000dd  (
    .G(\blk000000dc/sig00000cb2 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000001f6/blk000001fa  (
    .C(aclk),
    .CE(\blk000001f6/sig00000cb9 ),
    .D(\blk000001f6/sig00000cba ),
    .Q(sig000002c0)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk000001f6/blk000001f9  (
    .A0(\blk000001f6/sig00000cb8 ),
    .A1(\blk000001f6/sig00000cb9 ),
    .A2(\blk000001f6/sig00000cb9 ),
    .A3(\blk000001f6/sig00000cb8 ),
    .CE(\blk000001f6/sig00000cb9 ),
    .CLK(aclk),
    .D(sig000002c1),
    .Q(\blk000001f6/sig00000cba ),
    .Q15(\NLW_blk000001f6/blk000001f9_Q15_UNCONNECTED )
  );
  VCC   \blk000001f6/blk000001f8  (
    .P(\blk000001f6/sig00000cb9 )
  );
  GND   \blk000001f6/blk000001f7  (
    .G(\blk000001f6/sig00000cb8 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000002a3/blk000002a9  (
    .C(aclk),
    .CE(\blk000002a3/sig00000cc1 ),
    .D(\blk000002a3/sig00000cc3 ),
    .Q(sig000000c1)
  );
  SRLC32E #(
    .INIT ( 32'h00000000 ))
  \blk000002a3/blk000002a8  (
    .CLK(aclk),
    .D(sig00000206),
    .CE(\blk000002a3/sig00000cc1 ),
    .Q(\blk000002a3/sig00000cc3 ),
    .Q31(\NLW_blk000002a3/blk000002a8_Q31_UNCONNECTED ),
    .A({\blk000002a3/sig00000cc1 , \blk000002a3/sig00000cc1 , \blk000002a3/sig00000cc0 , \blk000002a3/sig00000cc1 , \blk000002a3/sig00000cc0 })
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000002a3/blk000002a7  (
    .C(aclk),
    .CE(\blk000002a3/sig00000cc1 ),
    .D(\blk000002a3/sig00000cc2 ),
    .Q(sig000000c0)
  );
  SRLC32E #(
    .INIT ( 32'h00000000 ))
  \blk000002a3/blk000002a6  (
    .CLK(aclk),
    .D(sig00000205),
    .CE(\blk000002a3/sig00000cc1 ),
    .Q(\blk000002a3/sig00000cc2 ),
    .Q31(\NLW_blk000002a3/blk000002a6_Q31_UNCONNECTED ),
    .A({\blk000002a3/sig00000cc1 , \blk000002a3/sig00000cc1 , \blk000002a3/sig00000cc0 , \blk000002a3/sig00000cc1 , \blk000002a3/sig00000cc0 })
  );
  VCC   \blk000002a3/blk000002a5  (
    .P(\blk000002a3/sig00000cc1 )
  );
  GND   \blk000002a3/blk000002a4  (
    .G(\blk000002a3/sig00000cc0 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000002aa/blk000002ae  (
    .C(aclk),
    .CE(\blk000002aa/sig00000cc8 ),
    .D(\blk000002aa/sig00000cc9 ),
    .Q(sig0000014f)
  );
  SRLC32E #(
    .INIT ( 32'h00000000 ))
  \blk000002aa/blk000002ad  (
    .CLK(aclk),
    .D(sig00000204),
    .CE(\blk000002aa/sig00000cc8 ),
    .Q(\blk000002aa/sig00000cc9 ),
    .Q31(\NLW_blk000002aa/blk000002ad_Q31_UNCONNECTED ),
    .A({\blk000002aa/sig00000cc8 , \blk000002aa/sig00000cc8 , \blk000002aa/sig00000cc7 , \blk000002aa/sig00000cc7 , \blk000002aa/sig00000cc8 })
  );
  VCC   \blk000002aa/blk000002ac  (
    .P(\blk000002aa/sig00000cc8 )
  );
  GND   \blk000002aa/blk000002ab  (
    .G(\blk000002aa/sig00000cc7 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000002af/blk000002b3  (
    .C(aclk),
    .CE(\blk000002af/sig00000cce ),
    .D(\blk000002af/sig00000ccf ),
    .Q(sig000001e0)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk000002af/blk000002b2  (
    .A0(\blk000002af/sig00000cce ),
    .A1(\blk000002af/sig00000ccd ),
    .A2(\blk000002af/sig00000ccd ),
    .A3(\blk000002af/sig00000cce ),
    .CE(\blk000002af/sig00000cce ),
    .CLK(aclk),
    .D(sig000001e1),
    .Q(\blk000002af/sig00000ccf ),
    .Q15(\NLW_blk000002af/blk000002b2_Q15_UNCONNECTED )
  );
  VCC   \blk000002af/blk000002b1  (
    .P(\blk000002af/sig00000cce )
  );
  GND   \blk000002af/blk000002b0  (
    .G(\blk000002af/sig00000ccd )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000002b4/blk000002b8  (
    .C(aclk),
    .CE(\blk000002b4/sig00000cd4 ),
    .D(\blk000002b4/sig00000cd5 ),
    .Q(sig0000009c)
  );
  SRLC32E #(
    .INIT ( 32'h00000000 ))
  \blk000002b4/blk000002b7  (
    .CLK(aclk),
    .D(sig00000162),
    .CE(\blk000002b4/sig00000cd4 ),
    .Q(\blk000002b4/sig00000cd5 ),
    .Q31(\NLW_blk000002b4/blk000002b7_Q31_UNCONNECTED ),
    .A({\blk000002b4/sig00000cd4 , \blk000002b4/sig00000cd4 , \blk000002b4/sig00000cd3 , \blk000002b4/sig00000cd4 , \blk000002b4/sig00000cd3 })
  );
  VCC   \blk000002b4/blk000002b6  (
    .P(\blk000002b4/sig00000cd4 )
  );
  GND   \blk000002b4/blk000002b5  (
    .G(\blk000002b4/sig00000cd3 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000002b9/blk000002bf  (
    .C(aclk),
    .CE(\blk000002b9/sig00000cdc ),
    .D(\blk000002b9/sig00000cde ),
    .Q(sig000001db)
  );
  SRLC32E #(
    .INIT ( 32'h00000000 ))
  \blk000002b9/blk000002be  (
    .CLK(aclk),
    .D(sig000001dd),
    .CE(\blk000002b9/sig00000cdc ),
    .Q(\blk000002b9/sig00000cde ),
    .Q31(\NLW_blk000002b9/blk000002be_Q31_UNCONNECTED ),
    .A({\blk000002b9/sig00000cdc , \blk000002b9/sig00000cdc , \blk000002b9/sig00000cdb , \blk000002b9/sig00000cdb , \blk000002b9/sig00000cdc })
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000002b9/blk000002bd  (
    .C(aclk),
    .CE(\blk000002b9/sig00000cdc ),
    .D(\blk000002b9/sig00000cdd ),
    .Q(sig000001da)
  );
  SRLC32E #(
    .INIT ( 32'h00000000 ))
  \blk000002b9/blk000002bc  (
    .CLK(aclk),
    .D(sig000001dc),
    .CE(\blk000002b9/sig00000cdc ),
    .Q(\blk000002b9/sig00000cdd ),
    .Q31(\NLW_blk000002b9/blk000002bc_Q31_UNCONNECTED ),
    .A({\blk000002b9/sig00000cdc , \blk000002b9/sig00000cdc , \blk000002b9/sig00000cdb , \blk000002b9/sig00000cdb , \blk000002b9/sig00000cdc })
  );
  VCC   \blk000002b9/blk000002bb  (
    .P(\blk000002b9/sig00000cdc )
  );
  GND   \blk000002b9/blk000002ba  (
    .G(\blk000002b9/sig00000cdb )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000002c0/blk000002c6  (
    .C(aclk),
    .CE(\blk000002c0/sig00000ce5 ),
    .D(\blk000002c0/sig00000ce7 ),
    .Q(sig000000bf)
  );
  SRLC32E #(
    .INIT ( 32'h00000000 ))
  \blk000002c0/blk000002c5  (
    .CLK(aclk),
    .D(sig000001df),
    .CE(\blk000002c0/sig00000ce5 ),
    .Q(\blk000002c0/sig00000ce7 ),
    .Q31(\NLW_blk000002c0/blk000002c5_Q31_UNCONNECTED ),
    .A({\blk000002c0/sig00000ce5 , \blk000002c0/sig00000ce5 , \blk000002c0/sig00000ce4 , \blk000002c0/sig00000ce5 , \blk000002c0/sig00000ce4 })
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000002c0/blk000002c4  (
    .C(aclk),
    .CE(\blk000002c0/sig00000ce5 ),
    .D(\blk000002c0/sig00000ce6 ),
    .Q(sig000000be)
  );
  SRLC32E #(
    .INIT ( 32'h00000000 ))
  \blk000002c0/blk000002c3  (
    .CLK(aclk),
    .D(sig000001de),
    .CE(\blk000002c0/sig00000ce5 ),
    .Q(\blk000002c0/sig00000ce6 ),
    .Q31(\NLW_blk000002c0/blk000002c3_Q31_UNCONNECTED ),
    .A({\blk000002c0/sig00000ce5 , \blk000002c0/sig00000ce5 , \blk000002c0/sig00000ce4 , \blk000002c0/sig00000ce5 , \blk000002c0/sig00000ce4 })
  );
  VCC   \blk000002c0/blk000002c2  (
    .P(\blk000002c0/sig00000ce5 )
  );
  GND   \blk000002c0/blk000002c1  (
    .G(\blk000002c0/sig00000ce4 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000003fc/blk000003ff  (
    .C(aclk),
    .CE(sig00000344),
    .D(\blk000003fc/sig00000ced ),
    .Q(sig0000052f)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk000003fc/blk000003fe  (
    .A0(\blk000003fc/sig00000cec ),
    .A1(\blk000003fc/sig00000cec ),
    .A2(\blk000003fc/sig00000cec ),
    .A3(\blk000003fc/sig00000cec ),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000530),
    .Q(\blk000003fc/sig00000ced ),
    .Q15(\NLW_blk000003fc/blk000003fe_Q15_UNCONNECTED )
  );
  GND   \blk000003fc/blk000003fd  (
    .G(\blk000003fc/sig00000cec )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000400/blk00000403  (
    .C(aclk),
    .CE(sig00000344),
    .D(\blk00000400/sig00000cf3 ),
    .Q(sig00000530)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000400/blk00000402  (
    .A0(\blk00000400/sig00000cf2 ),
    .A1(\blk00000400/sig00000cf2 ),
    .A2(\blk00000400/sig00000cf2 ),
    .A3(\blk00000400/sig00000cf2 ),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000531),
    .Q(\blk00000400/sig00000cf3 ),
    .Q15(\NLW_blk00000400/blk00000402_Q15_UNCONNECTED )
  );
  GND   \blk00000400/blk00000401  (
    .G(\blk00000400/sig00000cf2 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000404/blk00000408  (
    .C(aclk),
    .CE(\blk00000404/sig00000cf8 ),
    .D(\blk00000404/sig00000cf9 ),
    .Q(sig0000052e)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000404/blk00000407  (
    .A0(\blk00000404/sig00000cf7 ),
    .A1(\blk00000404/sig00000cf8 ),
    .A2(\blk00000404/sig00000cf7 ),
    .A3(\blk00000404/sig00000cf7 ),
    .CE(\blk00000404/sig00000cf8 ),
    .CLK(aclk),
    .D(sig0000052f),
    .Q(\blk00000404/sig00000cf9 ),
    .Q15(\NLW_blk00000404/blk00000407_Q15_UNCONNECTED )
  );
  VCC   \blk00000404/blk00000406  (
    .P(\blk00000404/sig00000cf8 )
  );
  GND   \blk00000404/blk00000405  (
    .G(\blk00000404/sig00000cf7 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000503/blk00000507  (
    .C(aclk),
    .CE(\blk00000503/sig00000cfe ),
    .D(\blk00000503/sig00000cff ),
    .Q(sig000001af)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000503/blk00000506  (
    .A0(\blk00000503/sig00000cfd ),
    .A1(\blk00000503/sig00000cfe ),
    .A2(\blk00000503/sig00000cfe ),
    .A3(\blk00000503/sig00000cfe ),
    .CE(\blk00000503/sig00000cfe ),
    .CLK(aclk),
    .D(sig00000162),
    .Q(\blk00000503/sig00000cff ),
    .Q15(\NLW_blk00000503/blk00000506_Q15_UNCONNECTED )
  );
  VCC   \blk00000503/blk00000505  (
    .P(\blk00000503/sig00000cfe )
  );
  GND   \blk00000503/blk00000504  (
    .G(\blk00000503/sig00000cfd )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000508/blk0000050b  (
    .C(aclk),
    .CE(sig00000344),
    .D(\blk00000508/sig00000d05 ),
    .Q(sig000005e8)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000508/blk0000050a  (
    .A0(\blk00000508/sig00000d04 ),
    .A1(\blk00000508/sig00000d04 ),
    .A2(\blk00000508/sig00000d04 ),
    .A3(\blk00000508/sig00000d04 ),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000005e9),
    .Q(\blk00000508/sig00000d05 ),
    .Q15(\NLW_blk00000508/blk0000050a_Q15_UNCONNECTED )
  );
  GND   \blk00000508/blk00000509  (
    .G(\blk00000508/sig00000d04 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000522/blk00000545  (
    .C(aclk),
    .CE(\blk00000522/sig00000d2b ),
    .D(\blk00000522/sig00000d2d ),
    .Q(sig00000198)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000522/blk00000544  (
    .A0(\blk00000522/sig00000d2a ),
    .A1(\blk00000522/sig00000d2a ),
    .A2(\blk00000522/sig00000d2a ),
    .A3(\blk00000522/sig00000d2a ),
    .CE(\blk00000522/sig00000d2b ),
    .CLK(aclk),
    .D(sig000005ea),
    .Q(\blk00000522/sig00000d2d ),
    .Q15(\NLW_blk00000522/blk00000544_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000522/blk00000543  (
    .C(aclk),
    .CE(\blk00000522/sig00000d2b ),
    .D(\blk00000522/sig00000d2c ),
    .Q(sig000005e7)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000522/blk00000542  (
    .A0(\blk00000522/sig00000d2a ),
    .A1(\blk00000522/sig00000d2a ),
    .A2(\blk00000522/sig00000d2a ),
    .A3(\blk00000522/sig00000d2a ),
    .CE(\blk00000522/sig00000d2b ),
    .CLK(aclk),
    .D(sig000005e5),
    .Q(\blk00000522/sig00000d2c ),
    .Q15(\NLW_blk00000522/blk00000542_Q15_UNCONNECTED )
  );
  VCC   \blk00000522/blk00000541  (
    .P(\blk00000522/sig00000d2b )
  );
  GND   \blk00000522/blk00000540  (
    .G(\blk00000522/sig00000d2a )
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  \blk00000522/blk0000053f  (
    .I0(\blk00000522/sig00000d0a ),
    .I1(\blk00000522/sig00000d19 ),
    .I2(\blk00000522/sig00000d1b ),
    .O(\blk00000522/sig00000d1e )
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  \blk00000522/blk0000053e  (
    .I0(\blk00000522/sig00000d09 ),
    .I1(\blk00000522/sig00000d0a ),
    .O(\blk00000522/sig00000d1d )
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  \blk00000522/blk0000053d  (
    .I0(\blk00000522/sig00000d0a ),
    .I1(\blk00000522/sig00000d1b ),
    .I2(\blk00000522/sig00000d19 ),
    .O(\blk00000522/sig00000d21 )
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  \blk00000522/blk0000053c  (
    .I0(\blk00000522/sig00000d0a ),
    .I1(\blk00000522/sig00000d1a ),
    .I2(\blk00000522/sig00000d16 ),
    .O(\blk00000522/sig00000d20 )
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  \blk00000522/blk0000053b  (
    .I0(\blk00000522/sig00000d0a ),
    .I1(\blk00000522/sig00000d16 ),
    .I2(\blk00000522/sig00000d1a ),
    .O(\blk00000522/sig00000d1f )
  );
  LUT2 #(
    .INIT ( 4'h8 ))
  \blk00000522/blk0000053a  (
    .I0(\blk00000522/sig00000d0a ),
    .I1(\blk00000522/sig00000d09 ),
    .O(\blk00000522/sig00000d1c )
  );
  LUT2 #(
    .INIT ( 4'h1 ))
  \blk00000522/blk00000539  (
    .I0(sig000005ea),
    .I1(sig000005eb),
    .O(\blk00000522/sig00000d29 )
  );
  LUT2 #(
    .INIT ( 4'hE ))
  \blk00000522/blk00000538  (
    .I0(sig000005eb),
    .I1(sig000005ea),
    .O(\blk00000522/sig00000d27 )
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  \blk00000522/blk00000537  (
    .I0(sig000005eb),
    .I1(sig000005ea),
    .O(\blk00000522/sig00000d26 )
  );
  LUT2 #(
    .INIT ( 4'h8 ))
  \blk00000522/blk00000536  (
    .I0(sig000005ea),
    .I1(sig000005eb),
    .O(\blk00000522/sig00000d25 )
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  \blk00000522/blk00000535  (
    .I0(sig000005ea),
    .I1(sig000005eb),
    .O(\blk00000522/sig00000d24 )
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  \blk00000522/blk00000534  (
    .I0(sig000005ea),
    .I1(sig000005eb),
    .O(\blk00000522/sig00000d23 )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000522/blk00000533  (
    .C(aclk),
    .D(\blk00000522/sig00000d1d ),
    .Q(sig000001ae)
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000522/blk00000532  (
    .C(aclk),
    .D(\blk00000522/sig00000d1c ),
    .Q(sig000001a0)
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000522/blk00000531  (
    .C(aclk),
    .D(\blk00000522/sig00000d17 ),
    .Q(sig0000019d)
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000522/blk00000530  (
    .C(aclk),
    .D(\blk00000522/sig00000d18 ),
    .Q(sig0000019c)
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000522/blk0000052f  (
    .C(aclk),
    .D(\blk00000522/sig00000d21 ),
    .Q(sig0000019b)
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000522/blk0000052e  (
    .C(aclk),
    .D(\blk00000522/sig00000d1f ),
    .Q(sig00000199)
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000522/blk0000052d  (
    .C(aclk),
    .D(\blk00000522/sig00000d1e ),
    .Q(sig00000194)
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000522/blk0000052c  (
    .C(aclk),
    .D(\blk00000522/sig00000d20 ),
    .Q(sig00000193)
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000522/blk0000052b  (
    .C(aclk),
    .D(\blk00000522/sig00000d0a ),
    .Q(sig000005e6)
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000522/blk0000052a  (
    .C(aclk),
    .D(\blk00000522/sig00000d29 ),
    .Q(\blk00000522/sig00000d09 )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000522/blk00000529  (
    .C(aclk),
    .D(\blk00000522/sig00000d27 ),
    .Q(\blk00000522/sig00000d17 )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000522/blk00000528  (
    .C(aclk),
    .D(\blk00000522/sig00000d26 ),
    .Q(\blk00000522/sig00000d18 )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000522/blk00000527  (
    .C(aclk),
    .D(\blk00000522/sig00000d23 ),
    .Q(\blk00000522/sig00000d1b )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000522/blk00000526  (
    .C(aclk),
    .D(sig000005eb),
    .Q(\blk00000522/sig00000d16 )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000522/blk00000525  (
    .C(aclk),
    .D(\blk00000522/sig00000d25 ),
    .Q(\blk00000522/sig00000d19 )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000522/blk00000524  (
    .C(aclk),
    .D(\blk00000522/sig00000d24 ),
    .Q(\blk00000522/sig00000d1a )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000522/blk00000523  (
    .C(aclk),
    .D(sig000005ec),
    .Q(\blk00000522/sig00000d0a )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000640/blk00000644  (
    .C(aclk),
    .CE(sig00000344),
    .D(\blk00000640/sig00000e36 ),
    .Q(sig00000890)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000640/blk00000643  (
    .A0(\blk00000640/sig00000e35 ),
    .A1(\blk00000640/sig00000e34 ),
    .A2(\blk00000640/sig00000e34 ),
    .A3(\blk00000640/sig00000e34 ),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig0000009d),
    .Q(\blk00000640/sig00000e36 ),
    .Q15(\NLW_blk00000640/blk00000643_Q15_UNCONNECTED )
  );
  VCC   \blk00000640/blk00000642  (
    .P(\blk00000640/sig00000e35 )
  );
  GND   \blk00000640/blk00000641  (
    .G(\blk00000640/sig00000e34 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000659/blk0000065c  (
    .C(aclk),
    .CE(sig00000344),
    .D(\blk00000659/sig00000e3c ),
    .Q(sig000009b1)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000659/blk0000065b  (
    .A0(\blk00000659/sig00000e3b ),
    .A1(\blk00000659/sig00000e3b ),
    .A2(\blk00000659/sig00000e3b ),
    .A3(\blk00000659/sig00000e3b ),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig000009b2),
    .Q(\blk00000659/sig00000e3c ),
    .Q15(\NLW_blk00000659/blk0000065b_Q15_UNCONNECTED )
  );
  GND   \blk00000659/blk0000065a  (
    .G(\blk00000659/sig00000e3b )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000007cb/blk000007cf  (
    .C(aclk),
    .CE(\blk000007cb/sig00000e41 ),
    .D(\blk000007cb/sig00000e42 ),
    .Q(sig0000088e)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk000007cb/blk000007ce  (
    .A0(\blk000007cb/sig00000e41 ),
    .A1(\blk000007cb/sig00000e41 ),
    .A2(\blk000007cb/sig00000e40 ),
    .A3(\blk000007cb/sig00000e40 ),
    .CE(\blk000007cb/sig00000e41 ),
    .CLK(aclk),
    .D(sig0000088f),
    .Q(\blk000007cb/sig00000e42 ),
    .Q15(\NLW_blk000007cb/blk000007ce_Q15_UNCONNECTED )
  );
  VCC   \blk000007cb/blk000007cd  (
    .P(\blk000007cb/sig00000e41 )
  );
  GND   \blk000007cb/blk000007cc  (
    .G(\blk000007cb/sig00000e40 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk0000083a/blk0000083d  (
    .C(aclk),
    .CE(sig00000344),
    .D(\blk0000083a/sig00000e48 ),
    .Q(sig00000c20)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk0000083a/blk0000083c  (
    .A0(\blk0000083a/sig00000e47 ),
    .A1(\blk0000083a/sig00000e47 ),
    .A2(\blk0000083a/sig00000e47 ),
    .A3(\blk0000083a/sig00000e47 ),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000c21),
    .Q(\blk0000083a/sig00000e48 ),
    .Q15(\NLW_blk0000083a/blk0000083c_Q15_UNCONNECTED )
  );
  GND   \blk0000083a/blk0000083b  (
    .G(\blk0000083a/sig00000e47 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk0000083e/blk00000841  (
    .C(aclk),
    .CE(sig00000344),
    .D(\blk0000083e/sig00000e4e ),
    .Q(sig00000c1f)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk0000083e/blk00000840  (
    .A0(\blk0000083e/sig00000e4d ),
    .A1(\blk0000083e/sig00000e4d ),
    .A2(\blk0000083e/sig00000e4d ),
    .A3(\blk0000083e/sig00000e4d ),
    .CE(sig00000344),
    .CLK(aclk),
    .D(sig00000c20),
    .Q(\blk0000083e/sig00000e4e ),
    .Q15(\NLW_blk0000083e/blk00000840_Q15_UNCONNECTED )
  );
  GND   \blk0000083e/blk0000083f  (
    .G(\blk0000083e/sig00000e4d )
  );
// synthesis translate_on
endmodule