module outputs
  reg [15 : 0] dma_respSt_first;
  wire [640 : 0] to_mem_toM_first;
  wire [584 : 0] to_child_toC_first;
  wire [527 : 0] dma_respLd_first;
  wire [102 : 0] cRqStuck_get;
  wire [67 : 0] perf_resp;
  wire RDY_cRqStuck_get,
       RDY_dma_memReq_enq,
       RDY_dma_memReq_notFull,
       RDY_dma_respLd_deq,
       RDY_dma_respLd_first,
       RDY_dma_respLd_notEmpty,
       RDY_dma_respSt_deq,
       RDY_dma_respSt_first,
       RDY_dma_respSt_notEmpty,
       RDY_perf_req,
       RDY_perf_resp,
       RDY_perf_respValid,
       RDY_perf_setStatus,
       RDY_to_child_rqFromC_enq,
       RDY_to_child_rqFromC_notFull,
       RDY_to_child_rsFromC_enq,
       RDY_to_child_rsFromC_notFull,
       RDY_to_child_toC_deq,
       RDY_to_child_toC_first,
       RDY_to_child_toC_notEmpty,
       RDY_to_mem_rsFromM_enq,
       RDY_to_mem_rsFromM_notFull,
       RDY_to_mem_toM_deq,
       RDY_to_mem_toM_first,
       RDY_to_mem_toM_notEmpty,
       dma_memReq_notFull,
       dma_respLd_notEmpty,
       dma_respSt_notEmpty,
       perf_respValid,
       to_child_rqFromC_notFull,
       to_child_rsFromC_notFull,
       to_child_toC_notEmpty,
       to_mem_rsFromM_notFull,
       to_mem_toM_notEmpty;
  // inlined wires
  reg [641 : 0] cache_toMQ_enqReq_lat_0$wget;
  reg [6 : 0] cache_rsToCIndexQ_enqReq_lat_0$wget;
  wire [656 : 0] cache_rqFromDmaQ_enqReq_lat_0$wget;
  wire [585 : 0] cache_toCQ_enqReq_lat_0$wget;
  wire [581 : 0] cache_rsFromCQ_enqReq_lat_0$wget;
  wire [528 : 0] cache_rsLdToDmaQ_enqReq_lat_0$wget;
  wire [517 : 0] cache_rsFromMQ_enqReq_lat_0$wget;
  wire [74 : 0] cache_rqFromCQ_enqReq_lat_0$wget;
  wire [16 : 0] cache_rsStToDmaQ_enqReq_lat_0$wget;
  wire [4 : 0] cache_cRqRetryIndexQ_enqReq_lat_0$wget,
	       perfReqQ_enqReq_lat_0$wget;
  wire cache_cRqRetryIndexQ_enqReq_lat_0$whas,
       cache_rsFromMQ_deqReq_lat_0$whas,
       cache_rsToCIndexQ_enqReq_lat_0$whas,
       cache_toCQ_enqReq_lat_0$whas,
       cache_toMQ_enqReq_lat_0$whas;
  // register cache_cRqRetryIndexQ_clearReq_rl
  reg cache_cRqRetryIndexQ_clearReq_rl;
  wire cache_cRqRetryIndexQ_clearReq_rl$D_IN,
       cache_cRqRetryIndexQ_clearReq_rl$EN;
  // register cache_cRqRetryIndexQ_data_0
  reg [3 : 0] cache_cRqRetryIndexQ_data_0;
  wire [3 : 0] cache_cRqRetryIndexQ_data_0$D_IN;
  wire cache_cRqRetryIndexQ_data_0$EN;
  // register cache_cRqRetryIndexQ_data_1
  reg [3 : 0] cache_cRqRetryIndexQ_data_1;
  wire [3 : 0] cache_cRqRetryIndexQ_data_1$D_IN;
  wire cache_cRqRetryIndexQ_data_1$EN;
  // register cache_cRqRetryIndexQ_data_10
  reg [3 : 0] cache_cRqRetryIndexQ_data_10;
  wire [3 : 0] cache_cRqRetryIndexQ_data_10$D_IN;
  wire cache_cRqRetryIndexQ_data_10$EN;
  // register cache_cRqRetryIndexQ_data_11
  reg [3 : 0] cache_cRqRetryIndexQ_data_11;
  wire [3 : 0] cache_cRqRetryIndexQ_data_11$D_IN;
  wire cache_cRqRetryIndexQ_data_11$EN;
  // register cache_cRqRetryIndexQ_data_12
  reg [3 : 0] cache_cRqRetryIndexQ_data_12;
  wire [3 : 0] cache_cRqRetryIndexQ_data_12$D_IN;
  wire cache_cRqRetryIndexQ_data_12$EN;
  // register cache_cRqRetryIndexQ_data_13
  reg [3 : 0] cache_cRqRetryIndexQ_data_13;
  wire [3 : 0] cache_cRqRetryIndexQ_data_13$D_IN;
  wire cache_cRqRetryIndexQ_data_13$EN;
  // register cache_cRqRetryIndexQ_data_14
  reg [3 : 0] cache_cRqRetryIndexQ_data_14;
  wire [3 : 0] cache_cRqRetryIndexQ_data_14$D_IN;
  wire cache_cRqRetryIndexQ_data_14$EN;
  // register cache_cRqRetryIndexQ_data_15
  reg [3 : 0] cache_cRqRetryIndexQ_data_15;
  wire [3 : 0] cache_cRqRetryIndexQ_data_15$D_IN;
  wire cache_cRqRetryIndexQ_data_15$EN;
  // register cache_cRqRetryIndexQ_data_2
  reg [3 : 0] cache_cRqRetryIndexQ_data_2;
  wire [3 : 0] cache_cRqRetryIndexQ_data_2$D_IN;
  wire cache_cRqRetryIndexQ_data_2$EN;
  // register cache_cRqRetryIndexQ_data_3
  reg [3 : 0] cache_cRqRetryIndexQ_data_3;
  wire [3 : 0] cache_cRqRetryIndexQ_data_3$D_IN;
  wire cache_cRqRetryIndexQ_data_3$EN;
  // register cache_cRqRetryIndexQ_data_4
  reg [3 : 0] cache_cRqRetryIndexQ_data_4;
  wire [3 : 0] cache_cRqRetryIndexQ_data_4$D_IN;
  wire cache_cRqRetryIndexQ_data_4$EN;
  // register cache_cRqRetryIndexQ_data_5
  reg [3 : 0] cache_cRqRetryIndexQ_data_5;
  wire [3 : 0] cache_cRqRetryIndexQ_data_5$D_IN;
  wire cache_cRqRetryIndexQ_data_5$EN;
  // register cache_cRqRetryIndexQ_data_6
  reg [3 : 0] cache_cRqRetryIndexQ_data_6;
  wire [3 : 0] cache_cRqRetryIndexQ_data_6$D_IN;
  wire cache_cRqRetryIndexQ_data_6$EN;
  // register cache_cRqRetryIndexQ_data_7
  reg [3 : 0] cache_cRqRetryIndexQ_data_7;
  wire [3 : 0] cache_cRqRetryIndexQ_data_7$D_IN;
  wire cache_cRqRetryIndexQ_data_7$EN;
  // register cache_cRqRetryIndexQ_data_8
  reg [3 : 0] cache_cRqRetryIndexQ_data_8;
  wire [3 : 0] cache_cRqRetryIndexQ_data_8$D_IN;
  wire cache_cRqRetryIndexQ_data_8$EN;
  // register cache_cRqRetryIndexQ_data_9
  reg [3 : 0] cache_cRqRetryIndexQ_data_9;
  wire [3 : 0] cache_cRqRetryIndexQ_data_9$D_IN;
  wire cache_cRqRetryIndexQ_data_9$EN;
  // register cache_cRqRetryIndexQ_deqP
  reg [3 : 0] cache_cRqRetryIndexQ_deqP;
  wire [3 : 0] cache_cRqRetryIndexQ_deqP$D_IN;
  wire cache_cRqRetryIndexQ_deqP$EN;
  // register cache_cRqRetryIndexQ_deqReq_rl
  reg cache_cRqRetryIndexQ_deqReq_rl;
  wire cache_cRqRetryIndexQ_deqReq_rl$D_IN, cache_cRqRetryIndexQ_deqReq_rl$EN;
  // register cache_cRqRetryIndexQ_empty
  reg cache_cRqRetryIndexQ_empty;
  wire cache_cRqRetryIndexQ_empty$D_IN, cache_cRqRetryIndexQ_empty$EN;
  // register cache_cRqRetryIndexQ_enqP
  reg [3 : 0] cache_cRqRetryIndexQ_enqP;
  wire [3 : 0] cache_cRqRetryIndexQ_enqP$D_IN;
  wire cache_cRqRetryIndexQ_enqP$EN;
  // register cache_cRqRetryIndexQ_enqReq_rl
  reg [4 : 0] cache_cRqRetryIndexQ_enqReq_rl;
  wire [4 : 0] cache_cRqRetryIndexQ_enqReq_rl$D_IN;
  wire cache_cRqRetryIndexQ_enqReq_rl$EN;
  // register cache_cRqRetryIndexQ_full
  reg cache_cRqRetryIndexQ_full;
  wire cache_cRqRetryIndexQ_full$D_IN, cache_cRqRetryIndexQ_full$EN;
  // register cache_doLdAfterReplace
  reg cache_doLdAfterReplace;
  wire cache_doLdAfterReplace$D_IN, cache_doLdAfterReplace$EN;
  // register cache_priorNewCRqSrc
  reg cache_priorNewCRqSrc;
  wire cache_priorNewCRqSrc$D_IN, cache_priorNewCRqSrc$EN;
  // register cache_rqFromCQ_clearReq_rl
  reg cache_rqFromCQ_clearReq_rl;
  wire cache_rqFromCQ_clearReq_rl$D_IN, cache_rqFromCQ_clearReq_rl$EN;
  // register cache_rqFromCQ_data_0
  reg [73 : 0] cache_rqFromCQ_data_0;
  wire [73 : 0] cache_rqFromCQ_data_0$D_IN;
  wire cache_rqFromCQ_data_0$EN;
  // register cache_rqFromCQ_data_1
  reg [73 : 0] cache_rqFromCQ_data_1;
  wire [73 : 0] cache_rqFromCQ_data_1$D_IN;
  wire cache_rqFromCQ_data_1$EN;
  // register cache_rqFromCQ_deqP
  reg cache_rqFromCQ_deqP;
  wire cache_rqFromCQ_deqP$D_IN, cache_rqFromCQ_deqP$EN;
  // register cache_rqFromCQ_deqReq_rl
  reg cache_rqFromCQ_deqReq_rl;
  wire cache_rqFromCQ_deqReq_rl$D_IN, cache_rqFromCQ_deqReq_rl$EN;
  // register cache_rqFromCQ_empty
  reg cache_rqFromCQ_empty;
  wire cache_rqFromCQ_empty$D_IN, cache_rqFromCQ_empty$EN;
  // register cache_rqFromCQ_enqP
  reg cache_rqFromCQ_enqP;
  wire cache_rqFromCQ_enqP$D_IN, cache_rqFromCQ_enqP$EN;
  // register cache_rqFromCQ_enqReq_rl
  reg [74 : 0] cache_rqFromCQ_enqReq_rl;
  wire [74 : 0] cache_rqFromCQ_enqReq_rl$D_IN;
  wire cache_rqFromCQ_enqReq_rl$EN;
  // register cache_rqFromCQ_full
  reg cache_rqFromCQ_full;
  wire cache_rqFromCQ_full$D_IN, cache_rqFromCQ_full$EN;
  // register cache_rqFromDmaQ_clearReq_rl
  reg cache_rqFromDmaQ_clearReq_rl;
  wire cache_rqFromDmaQ_clearReq_rl$D_IN, cache_rqFromDmaQ_clearReq_rl$EN;
  // register cache_rqFromDmaQ_data_0
  reg [655 : 0] cache_rqFromDmaQ_data_0;
  wire [655 : 0] cache_rqFromDmaQ_data_0$D_IN;
  wire cache_rqFromDmaQ_data_0$EN;
  // register cache_rqFromDmaQ_data_1
  reg [655 : 0] cache_rqFromDmaQ_data_1;
  wire [655 : 0] cache_rqFromDmaQ_data_1$D_IN;
  wire cache_rqFromDmaQ_data_1$EN;
  // register cache_rqFromDmaQ_deqP
  reg cache_rqFromDmaQ_deqP;
  wire cache_rqFromDmaQ_deqP$D_IN, cache_rqFromDmaQ_deqP$EN;
  // register cache_rqFromDmaQ_deqReq_rl
  reg cache_rqFromDmaQ_deqReq_rl;
  wire cache_rqFromDmaQ_deqReq_rl$D_IN, cache_rqFromDmaQ_deqReq_rl$EN;
  // register cache_rqFromDmaQ_empty
  reg cache_rqFromDmaQ_empty;
  wire cache_rqFromDmaQ_empty$D_IN, cache_rqFromDmaQ_empty$EN;
  // register cache_rqFromDmaQ_enqP
  reg cache_rqFromDmaQ_enqP;
  wire cache_rqFromDmaQ_enqP$D_IN, cache_rqFromDmaQ_enqP$EN;
  // register cache_rqFromDmaQ_enqReq_rl
  reg [656 : 0] cache_rqFromDmaQ_enqReq_rl;
  wire [656 : 0] cache_rqFromDmaQ_enqReq_rl$D_IN;
  wire cache_rqFromDmaQ_enqReq_rl$EN;
  // register cache_rqFromDmaQ_full
  reg cache_rqFromDmaQ_full;
  wire cache_rqFromDmaQ_full$D_IN, cache_rqFromDmaQ_full$EN;
  // register cache_rsFromCQ_clearReq_rl
  reg cache_rsFromCQ_clearReq_rl;
  wire cache_rsFromCQ_clearReq_rl$D_IN, cache_rsFromCQ_clearReq_rl$EN;
  // register cache_rsFromCQ_data_0
  reg [580 : 0] cache_rsFromCQ_data_0;
  wire [580 : 0] cache_rsFromCQ_data_0$D_IN;
  wire cache_rsFromCQ_data_0$EN;
  // register cache_rsFromCQ_data_1
  reg [580 : 0] cache_rsFromCQ_data_1;
  wire [580 : 0] cache_rsFromCQ_data_1$D_IN;
  wire cache_rsFromCQ_data_1$EN;
  // register cache_rsFromCQ_deqP
  reg cache_rsFromCQ_deqP;
  wire cache_rsFromCQ_deqP$D_IN, cache_rsFromCQ_deqP$EN;
  // register cache_rsFromCQ_deqReq_rl
  reg cache_rsFromCQ_deqReq_rl;
  wire cache_rsFromCQ_deqReq_rl$D_IN, cache_rsFromCQ_deqReq_rl$EN;
  // register cache_rsFromCQ_empty
  reg cache_rsFromCQ_empty;
  wire cache_rsFromCQ_empty$D_IN, cache_rsFromCQ_empty$EN;
  // register cache_rsFromCQ_enqP
  reg cache_rsFromCQ_enqP;
  wire cache_rsFromCQ_enqP$D_IN, cache_rsFromCQ_enqP$EN;
  // register cache_rsFromCQ_enqReq_rl
  reg [581 : 0] cache_rsFromCQ_enqReq_rl;
  wire [581 : 0] cache_rsFromCQ_enqReq_rl$D_IN;
  wire cache_rsFromCQ_enqReq_rl$EN;
  // register cache_rsFromCQ_full
  reg cache_rsFromCQ_full;
  wire cache_rsFromCQ_full$D_IN, cache_rsFromCQ_full$EN;
  // register cache_rsFromMQ_clearReq_rl
  reg cache_rsFromMQ_clearReq_rl;
  wire cache_rsFromMQ_clearReq_rl$D_IN, cache_rsFromMQ_clearReq_rl$EN;
  // register cache_rsFromMQ_data_0
  reg [516 : 0] cache_rsFromMQ_data_0;
  wire [516 : 0] cache_rsFromMQ_data_0$D_IN;
  wire cache_rsFromMQ_data_0$EN;
  // register cache_rsFromMQ_data_1
  reg [516 : 0] cache_rsFromMQ_data_1;
  wire [516 : 0] cache_rsFromMQ_data_1$D_IN;
  wire cache_rsFromMQ_data_1$EN;
  // register cache_rsFromMQ_deqP
  reg cache_rsFromMQ_deqP;
  wire cache_rsFromMQ_deqP$D_IN, cache_rsFromMQ_deqP$EN;
  // register cache_rsFromMQ_deqReq_rl
  reg cache_rsFromMQ_deqReq_rl;
  wire cache_rsFromMQ_deqReq_rl$D_IN, cache_rsFromMQ_deqReq_rl$EN;
  // register cache_rsFromMQ_empty
  reg cache_rsFromMQ_empty;
  wire cache_rsFromMQ_empty$D_IN, cache_rsFromMQ_empty$EN;
  // register cache_rsFromMQ_enqP
  reg cache_rsFromMQ_enqP;
  wire cache_rsFromMQ_enqP$D_IN, cache_rsFromMQ_enqP$EN;
  // register cache_rsFromMQ_enqReq_rl
  reg [517 : 0] cache_rsFromMQ_enqReq_rl;
  wire [517 : 0] cache_rsFromMQ_enqReq_rl$D_IN;
  wire cache_rsFromMQ_enqReq_rl$EN;
  // register cache_rsFromMQ_full
  reg cache_rsFromMQ_full;
  wire cache_rsFromMQ_full$D_IN, cache_rsFromMQ_full$EN;
  // register cache_rsLdToDmaQ_clearReq_rl
  reg cache_rsLdToDmaQ_clearReq_rl;
  wire cache_rsLdToDmaQ_clearReq_rl$D_IN, cache_rsLdToDmaQ_clearReq_rl$EN;
  // register cache_rsLdToDmaQ_data_0
  reg [527 : 0] cache_rsLdToDmaQ_data_0;
  wire [527 : 0] cache_rsLdToDmaQ_data_0$D_IN;
  wire cache_rsLdToDmaQ_data_0$EN;
  // register cache_rsLdToDmaQ_data_1
  reg [527 : 0] cache_rsLdToDmaQ_data_1;
  wire [527 : 0] cache_rsLdToDmaQ_data_1$D_IN;
  wire cache_rsLdToDmaQ_data_1$EN;
  // register cache_rsLdToDmaQ_deqP
  reg cache_rsLdToDmaQ_deqP;
  wire cache_rsLdToDmaQ_deqP$D_IN, cache_rsLdToDmaQ_deqP$EN;
  // register cache_rsLdToDmaQ_deqReq_rl
  reg cache_rsLdToDmaQ_deqReq_rl;
  wire cache_rsLdToDmaQ_deqReq_rl$D_IN, cache_rsLdToDmaQ_deqReq_rl$EN;
  // register cache_rsLdToDmaQ_empty
  reg cache_rsLdToDmaQ_empty;
  wire cache_rsLdToDmaQ_empty$D_IN, cache_rsLdToDmaQ_empty$EN;
  // register cache_rsLdToDmaQ_enqP
  reg cache_rsLdToDmaQ_enqP;
  wire cache_rsLdToDmaQ_enqP$D_IN, cache_rsLdToDmaQ_enqP$EN;
  // register cache_rsLdToDmaQ_enqReq_rl
  reg [528 : 0] cache_rsLdToDmaQ_enqReq_rl;
  wire [528 : 0] cache_rsLdToDmaQ_enqReq_rl$D_IN;
  wire cache_rsLdToDmaQ_enqReq_rl$EN;
  // register cache_rsLdToDmaQ_full
  reg cache_rsLdToDmaQ_full;
  wire cache_rsLdToDmaQ_full$D_IN, cache_rsLdToDmaQ_full$EN;
  // register cache_rsStToDmaQ_clearReq_rl
  reg cache_rsStToDmaQ_clearReq_rl;
  wire cache_rsStToDmaQ_clearReq_rl$D_IN, cache_rsStToDmaQ_clearReq_rl$EN;
  // register cache_rsStToDmaQ_data_0
  reg [15 : 0] cache_rsStToDmaQ_data_0;
  wire [15 : 0] cache_rsStToDmaQ_data_0$D_IN;
  wire cache_rsStToDmaQ_data_0$EN;
  // register cache_rsStToDmaQ_data_1
  reg [15 : 0] cache_rsStToDmaQ_data_1;
  wire [15 : 0] cache_rsStToDmaQ_data_1$D_IN;
  wire cache_rsStToDmaQ_data_1$EN;
  // register cache_rsStToDmaQ_deqP
  reg cache_rsStToDmaQ_deqP;
  wire cache_rsStToDmaQ_deqP$D_IN, cache_rsStToDmaQ_deqP$EN;
  // register cache_rsStToDmaQ_deqReq_rl
  reg cache_rsStToDmaQ_deqReq_rl;
  wire cache_rsStToDmaQ_deqReq_rl$D_IN, cache_rsStToDmaQ_deqReq_rl$EN;
  // register cache_rsStToDmaQ_empty
  reg cache_rsStToDmaQ_empty;
  wire cache_rsStToDmaQ_empty$D_IN, cache_rsStToDmaQ_empty$EN;
  // register cache_rsStToDmaQ_enqP
  reg cache_rsStToDmaQ_enqP;
  wire cache_rsStToDmaQ_enqP$D_IN, cache_rsStToDmaQ_enqP$EN;
  // register cache_rsStToDmaQ_enqReq_rl
  reg [16 : 0] cache_rsStToDmaQ_enqReq_rl;
  wire [16 : 0] cache_rsStToDmaQ_enqReq_rl$D_IN;
  wire cache_rsStToDmaQ_enqReq_rl$EN;
  // register cache_rsStToDmaQ_full
  reg cache_rsStToDmaQ_full;
  wire cache_rsStToDmaQ_full$D_IN, cache_rsStToDmaQ_full$EN;
  // register cache_rsToCIndexQ_clearReq_rl
  reg cache_rsToCIndexQ_clearReq_rl;
  wire cache_rsToCIndexQ_clearReq_rl$D_IN, cache_rsToCIndexQ_clearReq_rl$EN;
  // register cache_rsToCIndexQ_data_0
  reg [5 : 0] cache_rsToCIndexQ_data_0;
  wire [5 : 0] cache_rsToCIndexQ_data_0$D_IN;
  wire cache_rsToCIndexQ_data_0$EN;
  // register cache_rsToCIndexQ_data_1
  reg [5 : 0] cache_rsToCIndexQ_data_1;
  wire [5 : 0] cache_rsToCIndexQ_data_1$D_IN;
  wire cache_rsToCIndexQ_data_1$EN;
  // register cache_rsToCIndexQ_data_10
  reg [5 : 0] cache_rsToCIndexQ_data_10;
  wire [5 : 0] cache_rsToCIndexQ_data_10$D_IN;
  wire cache_rsToCIndexQ_data_10$EN;
  // register cache_rsToCIndexQ_data_11
  reg [5 : 0] cache_rsToCIndexQ_data_11;
  wire [5 : 0] cache_rsToCIndexQ_data_11$D_IN;
  wire cache_rsToCIndexQ_data_11$EN;
  // register cache_rsToCIndexQ_data_12
  reg [5 : 0] cache_rsToCIndexQ_data_12;
  wire [5 : 0] cache_rsToCIndexQ_data_12$D_IN;
  wire cache_rsToCIndexQ_data_12$EN;
  // register cache_rsToCIndexQ_data_13
  reg [5 : 0] cache_rsToCIndexQ_data_13;
  wire [5 : 0] cache_rsToCIndexQ_data_13$D_IN;
  wire cache_rsToCIndexQ_data_13$EN;
  // register cache_rsToCIndexQ_data_14
  reg [5 : 0] cache_rsToCIndexQ_data_14;
  wire [5 : 0] cache_rsToCIndexQ_data_14$D_IN;
  wire cache_rsToCIndexQ_data_14$EN;
  // register cache_rsToCIndexQ_data_15
  reg [5 : 0] cache_rsToCIndexQ_data_15;
  wire [5 : 0] cache_rsToCIndexQ_data_15$D_IN;
  wire cache_rsToCIndexQ_data_15$EN;
  // register cache_rsToCIndexQ_data_2
  reg [5 : 0] cache_rsToCIndexQ_data_2;
  wire [5 : 0] cache_rsToCIndexQ_data_2$D_IN;
  wire cache_rsToCIndexQ_data_2$EN;
  // register cache_rsToCIndexQ_data_3
  reg [5 : 0] cache_rsToCIndexQ_data_3;
  wire [5 : 0] cache_rsToCIndexQ_data_3$D_IN;
  wire cache_rsToCIndexQ_data_3$EN;
  // register cache_rsToCIndexQ_data_4
  reg [5 : 0] cache_rsToCIndexQ_data_4;
  wire [5 : 0] cache_rsToCIndexQ_data_4$D_IN;
  wire cache_rsToCIndexQ_data_4$EN;
  // register cache_rsToCIndexQ_data_5
  reg [5 : 0] cache_rsToCIndexQ_data_5;
  wire [5 : 0] cache_rsToCIndexQ_data_5$D_IN;
  wire cache_rsToCIndexQ_data_5$EN;
  // register cache_rsToCIndexQ_data_6
  reg [5 : 0] cache_rsToCIndexQ_data_6;
  wire [5 : 0] cache_rsToCIndexQ_data_6$D_IN;
  wire cache_rsToCIndexQ_data_6$EN;
  // register cache_rsToCIndexQ_data_7
  reg [5 : 0] cache_rsToCIndexQ_data_7;
  wire [5 : 0] cache_rsToCIndexQ_data_7$D_IN;
  wire cache_rsToCIndexQ_data_7$EN;
  // register cache_rsToCIndexQ_data_8
  reg [5 : 0] cache_rsToCIndexQ_data_8;
  wire [5 : 0] cache_rsToCIndexQ_data_8$D_IN;
  wire cache_rsToCIndexQ_data_8$EN;
  // register cache_rsToCIndexQ_data_9
  reg [5 : 0] cache_rsToCIndexQ_data_9;
  wire [5 : 0] cache_rsToCIndexQ_data_9$D_IN;
  wire cache_rsToCIndexQ_data_9$EN;
  // register cache_rsToCIndexQ_deqP
  reg [3 : 0] cache_rsToCIndexQ_deqP;
  wire [3 : 0] cache_rsToCIndexQ_deqP$D_IN;
  wire cache_rsToCIndexQ_deqP$EN;
  // register cache_rsToCIndexQ_deqReq_rl
  reg cache_rsToCIndexQ_deqReq_rl;
  wire cache_rsToCIndexQ_deqReq_rl$D_IN, cache_rsToCIndexQ_deqReq_rl$EN;
  // register cache_rsToCIndexQ_empty
  reg cache_rsToCIndexQ_empty;
  wire cache_rsToCIndexQ_empty$D_IN, cache_rsToCIndexQ_empty$EN;
  // register cache_rsToCIndexQ_enqP
  reg [3 : 0] cache_rsToCIndexQ_enqP;
  wire [3 : 0] cache_rsToCIndexQ_enqP$D_IN;
  wire cache_rsToCIndexQ_enqP$EN;
  // register cache_rsToCIndexQ_enqReq_rl
  reg [6 : 0] cache_rsToCIndexQ_enqReq_rl;
  wire [6 : 0] cache_rsToCIndexQ_enqReq_rl$D_IN;
  wire cache_rsToCIndexQ_enqReq_rl$EN;
  // register cache_rsToCIndexQ_full
  reg cache_rsToCIndexQ_full;
  wire cache_rsToCIndexQ_full$D_IN, cache_rsToCIndexQ_full$EN;
  // register cache_toCQ_clearReq_rl
  reg cache_toCQ_clearReq_rl;
  wire cache_toCQ_clearReq_rl$D_IN, cache_toCQ_clearReq_rl$EN;
  // register cache_toCQ_data_0
  reg [584 : 0] cache_toCQ_data_0;
  wire [584 : 0] cache_toCQ_data_0$D_IN;
  wire cache_toCQ_data_0$EN;
  // register cache_toCQ_data_1
  reg [584 : 0] cache_toCQ_data_1;
  wire [584 : 0] cache_toCQ_data_1$D_IN;
  wire cache_toCQ_data_1$EN;
  // register cache_toCQ_deqP
  reg cache_toCQ_deqP;
  wire cache_toCQ_deqP$D_IN, cache_toCQ_deqP$EN;
  // register cache_toCQ_deqReq_rl
  reg cache_toCQ_deqReq_rl;
  wire cache_toCQ_deqReq_rl$D_IN, cache_toCQ_deqReq_rl$EN;
  // register cache_toCQ_empty
  reg cache_toCQ_empty;
  wire cache_toCQ_empty$D_IN, cache_toCQ_empty$EN;
  // register cache_toCQ_enqP
  reg cache_toCQ_enqP;
  wire cache_toCQ_enqP$D_IN, cache_toCQ_enqP$EN;
  // register cache_toCQ_enqReq_rl
  reg [585 : 0] cache_toCQ_enqReq_rl;
  wire [585 : 0] cache_toCQ_enqReq_rl$D_IN;
  wire cache_toCQ_enqReq_rl$EN;
  // register cache_toCQ_full
  reg cache_toCQ_full;
  wire cache_toCQ_full$D_IN, cache_toCQ_full$EN;
  // register cache_toMQ_clearReq_rl
  reg cache_toMQ_clearReq_rl;
  wire cache_toMQ_clearReq_rl$D_IN, cache_toMQ_clearReq_rl$EN;
  // register cache_toMQ_data_0
  reg [640 : 0] cache_toMQ_data_0;
  wire [640 : 0] cache_toMQ_data_0$D_IN;
  wire cache_toMQ_data_0$EN;
  // register cache_toMQ_data_1
  reg [640 : 0] cache_toMQ_data_1;
  wire [640 : 0] cache_toMQ_data_1$D_IN;
  wire cache_toMQ_data_1$EN;
  // register cache_toMQ_deqP
  reg cache_toMQ_deqP;
  wire cache_toMQ_deqP$D_IN, cache_toMQ_deqP$EN;
  // register cache_toMQ_deqReq_rl
  reg cache_toMQ_deqReq_rl;
  wire cache_toMQ_deqReq_rl$D_IN, cache_toMQ_deqReq_rl$EN;
  // register cache_toMQ_empty
  reg cache_toMQ_empty;
  wire cache_toMQ_empty$D_IN, cache_toMQ_empty$EN;
  // register cache_toMQ_enqP
  reg cache_toMQ_enqP;
  wire cache_toMQ_enqP$D_IN, cache_toMQ_enqP$EN;
  // register cache_toMQ_enqReq_rl
  reg [641 : 0] cache_toMQ_enqReq_rl;
  wire [641 : 0] cache_toMQ_enqReq_rl$D_IN;
  wire cache_toMQ_enqReq_rl$EN;
  // register cache_toMQ_full
  reg cache_toMQ_full;
  wire cache_toMQ_full$D_IN, cache_toMQ_full$EN;
  // register cache_whichCRq
  reg [3 : 0] cache_whichCRq;
  wire [3 : 0] cache_whichCRq$D_IN;
  wire cache_whichCRq$EN;
  // register perfReqQ_clearReq_rl
  reg perfReqQ_clearReq_rl;
  wire perfReqQ_clearReq_rl$D_IN, perfReqQ_clearReq_rl$EN;
  // register perfReqQ_data_0
  reg [3 : 0] perfReqQ_data_0;
  wire [3 : 0] perfReqQ_data_0$D_IN;
  wire perfReqQ_data_0$EN;
  // register perfReqQ_deqReq_rl
  reg perfReqQ_deqReq_rl;
  wire perfReqQ_deqReq_rl$D_IN, perfReqQ_deqReq_rl$EN;
  // register perfReqQ_empty
  reg perfReqQ_empty;
  wire perfReqQ_empty$D_IN, perfReqQ_empty$EN;
  // register perfReqQ_enqReq_rl
  reg [4 : 0] perfReqQ_enqReq_rl;
  wire [4 : 0] perfReqQ_enqReq_rl$D_IN;
  wire perfReqQ_enqReq_rl$EN;
  // register perfReqQ_full
  reg perfReqQ_full;
  wire perfReqQ_full$D_IN, perfReqQ_full$EN;
  // ports of submodule cache_cRqMshr
  reg [512 : 0] cache_cRqMshr$pipelineResp_setData_d;
  reg [64 : 0] cache_cRqMshr$pipelineResp_setStateSlot_slot;
  reg [3 : 0] cache_cRqMshr$sendRsToDmaC_getRq_n,
	      cache_cRqMshr$sendRsToDmaC_releaseEntry_n;
  reg [2 : 0] cache_cRqMshr$pipelineResp_setStateSlot_state;
  wire [512 : 0] cache_cRqMshr$mRsDeq_setData_d,
		 cache_cRqMshr$pipelineResp_getData,
		 cache_cRqMshr$sendRsToDmaC_getData,
		 cache_cRqMshr$sendToM_getData,
		 cache_cRqMshr$transfer_getEmptyEntryInit_d;
  wire [167 : 0] cache_cRqMshr$stuck_get;
  wire [151 : 0] cache_cRqMshr$pipelineResp_getRq,
		 cache_cRqMshr$sendRqToC_getRq,
		 cache_cRqMshr$sendRsToDmaC_getRq,
		 cache_cRqMshr$sendToM_getRq,
		 cache_cRqMshr$transfer_getEmptyEntryInit_r,
		 cache_cRqMshr$transfer_getRq,
		 cache_cRqMshr$transfer_hasEmptyEntry_r;
  wire [64 : 0] cache_cRqMshr$pipelineResp_getSlot,
		cache_cRqMshr$sendRqToC_getSlot,
		cache_cRqMshr$sendRqToC_setSlot_s,
		cache_cRqMshr$sendToM_getSlot,
		cache_cRqMshr$transfer_getSlot;
  wire [63 : 0] cache_cRqMshr$pipelineResp_searchEndOfChain_addr;
  wire [4 : 0] cache_cRqMshr$pipelineResp_getAddrSucc,
	       cache_cRqMshr$pipelineResp_getRepSucc,
	       cache_cRqMshr$pipelineResp_searchEndOfChain,
	       cache_cRqMshr$pipelineResp_setAddrSucc_succ,
	       cache_cRqMshr$pipelineResp_setRepSucc_succ,
	       cache_cRqMshr$sendRqToC_searchNeedRqChild,
	       cache_cRqMshr$sendRqToC_searchNeedRqChild_suggestIdx;
  wire [3 : 0] cache_cRqMshr$mRsDeq_setData_n,
	       cache_cRqMshr$pipelineResp_getAddrSucc_n,
	       cache_cRqMshr$pipelineResp_getData_n,
	       cache_cRqMshr$pipelineResp_getRepSucc_n,
	       cache_cRqMshr$pipelineResp_getRq_n,
	       cache_cRqMshr$pipelineResp_getSlot_n,
	       cache_cRqMshr$pipelineResp_getState_n,
	       cache_cRqMshr$pipelineResp_setAddrSucc_n,
	       cache_cRqMshr$pipelineResp_setData_n,
	       cache_cRqMshr$pipelineResp_setRepSucc_n,
	       cache_cRqMshr$pipelineResp_setStateSlot_n,
	       cache_cRqMshr$sendRqToC_getRq_n,
	       cache_cRqMshr$sendRqToC_getSlot_n,
	       cache_cRqMshr$sendRqToC_getState_n,
	       cache_cRqMshr$sendRqToC_setSlot_n,
	       cache_cRqMshr$sendRsToDmaC_getData_n,
	       cache_cRqMshr$sendToM_getData_n,
	       cache_cRqMshr$sendToM_getRq_n,
	       cache_cRqMshr$sendToM_getSlot_n,
	       cache_cRqMshr$transfer_getEmptyEntryInit,
	       cache_cRqMshr$transfer_getRq_n,
	       cache_cRqMshr$transfer_getSlot_n;
  wire [2 : 0] cache_cRqMshr$pipelineResp_getState,
	       cache_cRqMshr$sendRqToC_getState;
  wire cache_cRqMshr$EN_mRsDeq_setData,
       cache_cRqMshr$EN_pipelineResp_setAddrSucc,
       cache_cRqMshr$EN_pipelineResp_setData,
       cache_cRqMshr$EN_pipelineResp_setRepSucc,
       cache_cRqMshr$EN_pipelineResp_setStateSlot,
       cache_cRqMshr$EN_sendRqToC_setSlot,
       cache_cRqMshr$EN_sendRsToDmaC_releaseEntry,
       cache_cRqMshr$EN_stuck_get,
       cache_cRqMshr$EN_transfer_getEmptyEntryInit,
       cache_cRqMshr$RDY_sendRsToDmaC_releaseEntry,
       cache_cRqMshr$RDY_stuck_get,
       cache_cRqMshr$RDY_transfer_getEmptyEntryInit;
  // ports of submodule cache_cRqRetryIndexQ_clearReq_dummy2_0
  wire cache_cRqRetryIndexQ_clearReq_dummy2_0$D_IN,
       cache_cRqRetryIndexQ_clearReq_dummy2_0$EN;
  // ports of submodule cache_cRqRetryIndexQ_clearReq_dummy2_1
  wire cache_cRqRetryIndexQ_clearReq_dummy2_1$D_IN,
       cache_cRqRetryIndexQ_clearReq_dummy2_1$EN,
       cache_cRqRetryIndexQ_clearReq_dummy2_1$Q_OUT;
  // ports of submodule cache_cRqRetryIndexQ_deqReq_dummy2_0
  wire cache_cRqRetryIndexQ_deqReq_dummy2_0$D_IN,
       cache_cRqRetryIndexQ_deqReq_dummy2_0$EN;
  // ports of submodule cache_cRqRetryIndexQ_deqReq_dummy2_1
  wire cache_cRqRetryIndexQ_deqReq_dummy2_1$D_IN,
       cache_cRqRetryIndexQ_deqReq_dummy2_1$EN;
  // ports of submodule cache_cRqRetryIndexQ_deqReq_dummy2_2
  wire cache_cRqRetryIndexQ_deqReq_dummy2_2$D_IN,
       cache_cRqRetryIndexQ_deqReq_dummy2_2$EN,
       cache_cRqRetryIndexQ_deqReq_dummy2_2$Q_OUT;
  // ports of submodule cache_cRqRetryIndexQ_enqReq_dummy2_0
  wire cache_cRqRetryIndexQ_enqReq_dummy2_0$D_IN,
       cache_cRqRetryIndexQ_enqReq_dummy2_0$EN;
  // ports of submodule cache_cRqRetryIndexQ_enqReq_dummy2_1
  wire cache_cRqRetryIndexQ_enqReq_dummy2_1$D_IN,
       cache_cRqRetryIndexQ_enqReq_dummy2_1$EN;
  // ports of submodule cache_cRqRetryIndexQ_enqReq_dummy2_2
  wire cache_cRqRetryIndexQ_enqReq_dummy2_2$D_IN,
       cache_cRqRetryIndexQ_enqReq_dummy2_2$EN,
       cache_cRqRetryIndexQ_enqReq_dummy2_2$Q_OUT;
  // ports of submodule cache_pipeline
  reg [583 : 0] cache_pipeline$send_r;
  reg [573 : 0] cache_pipeline$deqWrite_wrRam;
  reg [4 : 0] cache_pipeline$deqWrite_swapRq;
  reg cache_pipeline$deqWrite_updateRep;
  wire [584 : 0] cache_pipeline$first, cache_pipeline$unguard_first;
  wire cache_pipeline$EN_deqWrite,
       cache_pipeline$EN_send,
       cache_pipeline$RDY_deqWrite,
       cache_pipeline$RDY_first,
       cache_pipeline$RDY_send,
       cache_pipeline$RDY_unguard_first,
       cache_pipeline$notEmpty;
  // ports of submodule cache_rqFromCQ_clearReq_dummy2_0
  wire cache_rqFromCQ_clearReq_dummy2_0$D_IN,
       cache_rqFromCQ_clearReq_dummy2_0$EN;
  // ports of submodule cache_rqFromCQ_clearReq_dummy2_1
  wire cache_rqFromCQ_clearReq_dummy2_1$D_IN,
       cache_rqFromCQ_clearReq_dummy2_1$EN,
       cache_rqFromCQ_clearReq_dummy2_1$Q_OUT;
  // ports of submodule cache_rqFromCQ_deqReq_dummy2_0
  wire cache_rqFromCQ_deqReq_dummy2_0$D_IN, cache_rqFromCQ_deqReq_dummy2_0$EN;
  // ports of submodule cache_rqFromCQ_deqReq_dummy2_1
  wire cache_rqFromCQ_deqReq_dummy2_1$D_IN, cache_rqFromCQ_deqReq_dummy2_1$EN;
  // ports of submodule cache_rqFromCQ_deqReq_dummy2_2
  wire cache_rqFromCQ_deqReq_dummy2_2$D_IN,
       cache_rqFromCQ_deqReq_dummy2_2$EN,
       cache_rqFromCQ_deqReq_dummy2_2$Q_OUT;
  // ports of submodule cache_rqFromCQ_enqReq_dummy2_0
  wire cache_rqFromCQ_enqReq_dummy2_0$D_IN, cache_rqFromCQ_enqReq_dummy2_0$EN;
  // ports of submodule cache_rqFromCQ_enqReq_dummy2_1
  wire cache_rqFromCQ_enqReq_dummy2_1$D_IN, cache_rqFromCQ_enqReq_dummy2_1$EN;
  // ports of submodule cache_rqFromCQ_enqReq_dummy2_2
  wire cache_rqFromCQ_enqReq_dummy2_2$D_IN,
       cache_rqFromCQ_enqReq_dummy2_2$EN,
       cache_rqFromCQ_enqReq_dummy2_2$Q_OUT;
  // ports of submodule cache_rqFromDmaQ_clearReq_dummy2_0
  wire cache_rqFromDmaQ_clearReq_dummy2_0$D_IN,
       cache_rqFromDmaQ_clearReq_dummy2_0$EN;
  // ports of submodule cache_rqFromDmaQ_clearReq_dummy2_1
  wire cache_rqFromDmaQ_clearReq_dummy2_1$D_IN,
       cache_rqFromDmaQ_clearReq_dummy2_1$EN,
       cache_rqFromDmaQ_clearReq_dummy2_1$Q_OUT;
  // ports of submodule cache_rqFromDmaQ_deqReq_dummy2_0
  wire cache_rqFromDmaQ_deqReq_dummy2_0$D_IN,
       cache_rqFromDmaQ_deqReq_dummy2_0$EN;
  // ports of submodule cache_rqFromDmaQ_deqReq_dummy2_1
  wire cache_rqFromDmaQ_deqReq_dummy2_1$D_IN,
       cache_rqFromDmaQ_deqReq_dummy2_1$EN;
  // ports of submodule cache_rqFromDmaQ_deqReq_dummy2_2
  wire cache_rqFromDmaQ_deqReq_dummy2_2$D_IN,
       cache_rqFromDmaQ_deqReq_dummy2_2$EN,
       cache_rqFromDmaQ_deqReq_dummy2_2$Q_OUT;
  // ports of submodule cache_rqFromDmaQ_enqReq_dummy2_0
  wire cache_rqFromDmaQ_enqReq_dummy2_0$D_IN,
       cache_rqFromDmaQ_enqReq_dummy2_0$EN;
  // ports of submodule cache_rqFromDmaQ_enqReq_dummy2_1
  wire cache_rqFromDmaQ_enqReq_dummy2_1$D_IN,
       cache_rqFromDmaQ_enqReq_dummy2_1$EN;
  // ports of submodule cache_rqFromDmaQ_enqReq_dummy2_2
  wire cache_rqFromDmaQ_enqReq_dummy2_2$D_IN,
       cache_rqFromDmaQ_enqReq_dummy2_2$EN,
       cache_rqFromDmaQ_enqReq_dummy2_2$Q_OUT;
  // ports of submodule cache_rsFromCQ_clearReq_dummy2_0
  wire cache_rsFromCQ_clearReq_dummy2_0$D_IN,
       cache_rsFromCQ_clearReq_dummy2_0$EN;
  // ports of submodule cache_rsFromCQ_clearReq_dummy2_1
  wire cache_rsFromCQ_clearReq_dummy2_1$D_IN,
       cache_rsFromCQ_clearReq_dummy2_1$EN,
       cache_rsFromCQ_clearReq_dummy2_1$Q_OUT;
  // ports of submodule cache_rsFromCQ_deqReq_dummy2_0
  wire cache_rsFromCQ_deqReq_dummy2_0$D_IN, cache_rsFromCQ_deqReq_dummy2_0$EN;
  // ports of submodule cache_rsFromCQ_deqReq_dummy2_1
  wire cache_rsFromCQ_deqReq_dummy2_1$D_IN, cache_rsFromCQ_deqReq_dummy2_1$EN;
  // ports of submodule cache_rsFromCQ_deqReq_dummy2_2
  wire cache_rsFromCQ_deqReq_dummy2_2$D_IN,
       cache_rsFromCQ_deqReq_dummy2_2$EN,
       cache_rsFromCQ_deqReq_dummy2_2$Q_OUT;
  // ports of submodule cache_rsFromCQ_enqReq_dummy2_0
  wire cache_rsFromCQ_enqReq_dummy2_0$D_IN, cache_rsFromCQ_enqReq_dummy2_0$EN;
  // ports of submodule cache_rsFromCQ_enqReq_dummy2_1
  wire cache_rsFromCQ_enqReq_dummy2_1$D_IN, cache_rsFromCQ_enqReq_dummy2_1$EN;
  // ports of submodule cache_rsFromCQ_enqReq_dummy2_2
  wire cache_rsFromCQ_enqReq_dummy2_2$D_IN,
       cache_rsFromCQ_enqReq_dummy2_2$EN,
       cache_rsFromCQ_enqReq_dummy2_2$Q_OUT;
  // ports of submodule cache_rsFromMQ_clearReq_dummy2_0
  wire cache_rsFromMQ_clearReq_dummy2_0$D_IN,
       cache_rsFromMQ_clearReq_dummy2_0$EN;
  // ports of submodule cache_rsFromMQ_clearReq_dummy2_1
  wire cache_rsFromMQ_clearReq_dummy2_1$D_IN,
       cache_rsFromMQ_clearReq_dummy2_1$EN,
       cache_rsFromMQ_clearReq_dummy2_1$Q_OUT;
  // ports of submodule cache_rsFromMQ_deqReq_dummy2_0
  wire cache_rsFromMQ_deqReq_dummy2_0$D_IN, cache_rsFromMQ_deqReq_dummy2_0$EN;
  // ports of submodule cache_rsFromMQ_deqReq_dummy2_1
  wire cache_rsFromMQ_deqReq_dummy2_1$D_IN, cache_rsFromMQ_deqReq_dummy2_1$EN;
  // ports of submodule cache_rsFromMQ_deqReq_dummy2_2
  wire cache_rsFromMQ_deqReq_dummy2_2$D_IN,
       cache_rsFromMQ_deqReq_dummy2_2$EN,
       cache_rsFromMQ_deqReq_dummy2_2$Q_OUT;
  // ports of submodule cache_rsFromMQ_enqReq_dummy2_0
  wire cache_rsFromMQ_enqReq_dummy2_0$D_IN, cache_rsFromMQ_enqReq_dummy2_0$EN;
  // ports of submodule cache_rsFromMQ_enqReq_dummy2_1
  wire cache_rsFromMQ_enqReq_dummy2_1$D_IN, cache_rsFromMQ_enqReq_dummy2_1$EN;
  // ports of submodule cache_rsFromMQ_enqReq_dummy2_2
  wire cache_rsFromMQ_enqReq_dummy2_2$D_IN,
       cache_rsFromMQ_enqReq_dummy2_2$EN,
       cache_rsFromMQ_enqReq_dummy2_2$Q_OUT;
  // ports of submodule cache_rsLdToDmaIndexQ
  wire [3 : 0] cache_rsLdToDmaIndexQ$D_IN, cache_rsLdToDmaIndexQ$D_OUT;
  wire cache_rsLdToDmaIndexQ$CLR,
       cache_rsLdToDmaIndexQ$DEQ,
       cache_rsLdToDmaIndexQ$EMPTY_N,
       cache_rsLdToDmaIndexQ$ENQ,
       cache_rsLdToDmaIndexQ$FULL_N;
  // ports of submodule cache_rsLdToDmaIndexQ_mRsDeq
  wire [3 : 0] cache_rsLdToDmaIndexQ_mRsDeq$D_IN,
	       cache_rsLdToDmaIndexQ_mRsDeq$D_OUT;
  wire cache_rsLdToDmaIndexQ_mRsDeq$CLR,
       cache_rsLdToDmaIndexQ_mRsDeq$DEQ,
       cache_rsLdToDmaIndexQ_mRsDeq$EMPTY_N,
       cache_rsLdToDmaIndexQ_mRsDeq$ENQ,
       cache_rsLdToDmaIndexQ_mRsDeq$FULL_N;
  // ports of submodule cache_rsLdToDmaIndexQ_pipelineResp
  wire [3 : 0] cache_rsLdToDmaIndexQ_pipelineResp$D_IN,
	       cache_rsLdToDmaIndexQ_pipelineResp$D_OUT;
  wire cache_rsLdToDmaIndexQ_pipelineResp$CLR,
       cache_rsLdToDmaIndexQ_pipelineResp$DEQ,
       cache_rsLdToDmaIndexQ_pipelineResp$EMPTY_N,
       cache_rsLdToDmaIndexQ_pipelineResp$ENQ,
       cache_rsLdToDmaIndexQ_pipelineResp$FULL_N;
  // ports of submodule cache_rsLdToDmaQ_clearReq_dummy2_0
  wire cache_rsLdToDmaQ_clearReq_dummy2_0$D_IN,
       cache_rsLdToDmaQ_clearReq_dummy2_0$EN;
  // ports of submodule cache_rsLdToDmaQ_clearReq_dummy2_1
  wire cache_rsLdToDmaQ_clearReq_dummy2_1$D_IN,
       cache_rsLdToDmaQ_clearReq_dummy2_1$EN,
       cache_rsLdToDmaQ_clearReq_dummy2_1$Q_OUT;
  // ports of submodule cache_rsLdToDmaQ_deqReq_dummy2_0
  wire cache_rsLdToDmaQ_deqReq_dummy2_0$D_IN,
       cache_rsLdToDmaQ_deqReq_dummy2_0$EN;
  // ports of submodule cache_rsLdToDmaQ_deqReq_dummy2_1
  wire cache_rsLdToDmaQ_deqReq_dummy2_1$D_IN,
       cache_rsLdToDmaQ_deqReq_dummy2_1$EN;
  // ports of submodule cache_rsLdToDmaQ_deqReq_dummy2_2
  wire cache_rsLdToDmaQ_deqReq_dummy2_2$D_IN,
       cache_rsLdToDmaQ_deqReq_dummy2_2$EN,
       cache_rsLdToDmaQ_deqReq_dummy2_2$Q_OUT;
  // ports of submodule cache_rsLdToDmaQ_enqReq_dummy2_0
  wire cache_rsLdToDmaQ_enqReq_dummy2_0$D_IN,
       cache_rsLdToDmaQ_enqReq_dummy2_0$EN;
  // ports of submodule cache_rsLdToDmaQ_enqReq_dummy2_1
  wire cache_rsLdToDmaQ_enqReq_dummy2_1$D_IN,
       cache_rsLdToDmaQ_enqReq_dummy2_1$EN;
  // ports of submodule cache_rsLdToDmaQ_enqReq_dummy2_2
  wire cache_rsLdToDmaQ_enqReq_dummy2_2$D_IN,
       cache_rsLdToDmaQ_enqReq_dummy2_2$EN,
       cache_rsLdToDmaQ_enqReq_dummy2_2$Q_OUT;
  // ports of submodule cache_rsStToDmaIndexQ
  wire [3 : 0] cache_rsStToDmaIndexQ$D_IN, cache_rsStToDmaIndexQ$D_OUT;
  wire cache_rsStToDmaIndexQ$CLR,
       cache_rsStToDmaIndexQ$DEQ,
       cache_rsStToDmaIndexQ$EMPTY_N,
       cache_rsStToDmaIndexQ$ENQ,
       cache_rsStToDmaIndexQ$FULL_N;
  // ports of submodule cache_rsStToDmaIndexQ_pipelineResp
  wire [3 : 0] cache_rsStToDmaIndexQ_pipelineResp$D_IN,
	       cache_rsStToDmaIndexQ_pipelineResp$D_OUT;
  wire cache_rsStToDmaIndexQ_pipelineResp$CLR,
       cache_rsStToDmaIndexQ_pipelineResp$DEQ,
       cache_rsStToDmaIndexQ_pipelineResp$EMPTY_N,
       cache_rsStToDmaIndexQ_pipelineResp$ENQ,
       cache_rsStToDmaIndexQ_pipelineResp$FULL_N;
  // ports of submodule cache_rsStToDmaIndexQ_sendToM
  wire [3 : 0] cache_rsStToDmaIndexQ_sendToM$D_IN,
	       cache_rsStToDmaIndexQ_sendToM$D_OUT;
  wire cache_rsStToDmaIndexQ_sendToM$CLR,
       cache_rsStToDmaIndexQ_sendToM$DEQ,
       cache_rsStToDmaIndexQ_sendToM$EMPTY_N,
       cache_rsStToDmaIndexQ_sendToM$ENQ,
       cache_rsStToDmaIndexQ_sendToM$FULL_N;
  // ports of submodule cache_rsStToDmaQ_clearReq_dummy2_0
  wire cache_rsStToDmaQ_clearReq_dummy2_0$D_IN,
       cache_rsStToDmaQ_clearReq_dummy2_0$EN;
  // ports of submodule cache_rsStToDmaQ_clearReq_dummy2_1
  wire cache_rsStToDmaQ_clearReq_dummy2_1$D_IN,
       cache_rsStToDmaQ_clearReq_dummy2_1$EN,
       cache_rsStToDmaQ_clearReq_dummy2_1$Q_OUT;
  // ports of submodule cache_rsStToDmaQ_deqReq_dummy2_0
  wire cache_rsStToDmaQ_deqReq_dummy2_0$D_IN,
       cache_rsStToDmaQ_deqReq_dummy2_0$EN;
  // ports of submodule cache_rsStToDmaQ_deqReq_dummy2_1
  wire cache_rsStToDmaQ_deqReq_dummy2_1$D_IN,
       cache_rsStToDmaQ_deqReq_dummy2_1$EN;
  // ports of submodule cache_rsStToDmaQ_deqReq_dummy2_2
  wire cache_rsStToDmaQ_deqReq_dummy2_2$D_IN,
       cache_rsStToDmaQ_deqReq_dummy2_2$EN,
       cache_rsStToDmaQ_deqReq_dummy2_2$Q_OUT;
  // ports of submodule cache_rsStToDmaQ_enqReq_dummy2_0
  wire cache_rsStToDmaQ_enqReq_dummy2_0$D_IN,
       cache_rsStToDmaQ_enqReq_dummy2_0$EN;
  // ports of submodule cache_rsStToDmaQ_enqReq_dummy2_1
  wire cache_rsStToDmaQ_enqReq_dummy2_1$D_IN,
       cache_rsStToDmaQ_enqReq_dummy2_1$EN;
  // ports of submodule cache_rsStToDmaQ_enqReq_dummy2_2
  wire cache_rsStToDmaQ_enqReq_dummy2_2$D_IN,
       cache_rsStToDmaQ_enqReq_dummy2_2$EN,
       cache_rsStToDmaQ_enqReq_dummy2_2$Q_OUT;
  // ports of submodule cache_rsToCIndexQ_clearReq_dummy2_0
  wire cache_rsToCIndexQ_clearReq_dummy2_0$D_IN,
       cache_rsToCIndexQ_clearReq_dummy2_0$EN;
  // ports of submodule cache_rsToCIndexQ_clearReq_dummy2_1
  wire cache_rsToCIndexQ_clearReq_dummy2_1$D_IN,
       cache_rsToCIndexQ_clearReq_dummy2_1$EN,
       cache_rsToCIndexQ_clearReq_dummy2_1$Q_OUT;
  // ports of submodule cache_rsToCIndexQ_deqReq_dummy2_0
  wire cache_rsToCIndexQ_deqReq_dummy2_0$D_IN,
       cache_rsToCIndexQ_deqReq_dummy2_0$EN;
  // ports of submodule cache_rsToCIndexQ_deqReq_dummy2_1
  wire cache_rsToCIndexQ_deqReq_dummy2_1$D_IN,
       cache_rsToCIndexQ_deqReq_dummy2_1$EN;
  // ports of submodule cache_rsToCIndexQ_deqReq_dummy2_2
  wire cache_rsToCIndexQ_deqReq_dummy2_2$D_IN,
       cache_rsToCIndexQ_deqReq_dummy2_2$EN,
       cache_rsToCIndexQ_deqReq_dummy2_2$Q_OUT;
  // ports of submodule cache_rsToCIndexQ_enqReq_dummy2_0
  wire cache_rsToCIndexQ_enqReq_dummy2_0$D_IN,
       cache_rsToCIndexQ_enqReq_dummy2_0$EN;
  // ports of submodule cache_rsToCIndexQ_enqReq_dummy2_1
  wire cache_rsToCIndexQ_enqReq_dummy2_1$D_IN,
       cache_rsToCIndexQ_enqReq_dummy2_1$EN;
  // ports of submodule cache_rsToCIndexQ_enqReq_dummy2_2
  wire cache_rsToCIndexQ_enqReq_dummy2_2$D_IN,
       cache_rsToCIndexQ_enqReq_dummy2_2$EN,
       cache_rsToCIndexQ_enqReq_dummy2_2$Q_OUT;
  // ports of submodule cache_toCQ_clearReq_dummy2_0
  wire cache_toCQ_clearReq_dummy2_0$D_IN, cache_toCQ_clearReq_dummy2_0$EN;
  // ports of submodule cache_toCQ_clearReq_dummy2_1
  wire cache_toCQ_clearReq_dummy2_1$D_IN,
       cache_toCQ_clearReq_dummy2_1$EN,
       cache_toCQ_clearReq_dummy2_1$Q_OUT;
  // ports of submodule cache_toCQ_deqReq_dummy2_0
  wire cache_toCQ_deqReq_dummy2_0$D_IN, cache_toCQ_deqReq_dummy2_0$EN;
  // ports of submodule cache_toCQ_deqReq_dummy2_1
  wire cache_toCQ_deqReq_dummy2_1$D_IN, cache_toCQ_deqReq_dummy2_1$EN;
  // ports of submodule cache_toCQ_deqReq_dummy2_2
  wire cache_toCQ_deqReq_dummy2_2$D_IN,
       cache_toCQ_deqReq_dummy2_2$EN,
       cache_toCQ_deqReq_dummy2_2$Q_OUT;
  // ports of submodule cache_toCQ_enqReq_dummy2_0
  wire cache_toCQ_enqReq_dummy2_0$D_IN, cache_toCQ_enqReq_dummy2_0$EN;
  // ports of submodule cache_toCQ_enqReq_dummy2_1
  wire cache_toCQ_enqReq_dummy2_1$D_IN, cache_toCQ_enqReq_dummy2_1$EN;
  // ports of submodule cache_toCQ_enqReq_dummy2_2
  wire cache_toCQ_enqReq_dummy2_2$D_IN,
       cache_toCQ_enqReq_dummy2_2$EN,
       cache_toCQ_enqReq_dummy2_2$Q_OUT;
  // ports of submodule cache_toMInfoQ
  wire [5 : 0] cache_toMInfoQ$D_IN, cache_toMInfoQ$D_OUT;
  wire cache_toMInfoQ$CLR,
       cache_toMInfoQ$DEQ,
       cache_toMInfoQ$EMPTY_N,
       cache_toMInfoQ$ENQ,
       cache_toMInfoQ$FULL_N;
  // ports of submodule cache_toMQ_clearReq_dummy2_0
  wire cache_toMQ_clearReq_dummy2_0$D_IN, cache_toMQ_clearReq_dummy2_0$EN;
  // ports of submodule cache_toMQ_clearReq_dummy2_1
  wire cache_toMQ_clearReq_dummy2_1$D_IN,
       cache_toMQ_clearReq_dummy2_1$EN,
       cache_toMQ_clearReq_dummy2_1$Q_OUT;
  // ports of submodule cache_toMQ_deqReq_dummy2_0
  wire cache_toMQ_deqReq_dummy2_0$D_IN, cache_toMQ_deqReq_dummy2_0$EN;
  // ports of submodule cache_toMQ_deqReq_dummy2_1
  wire cache_toMQ_deqReq_dummy2_1$D_IN, cache_toMQ_deqReq_dummy2_1$EN;
  // ports of submodule cache_toMQ_deqReq_dummy2_2
  wire cache_toMQ_deqReq_dummy2_2$D_IN,
       cache_toMQ_deqReq_dummy2_2$EN,
       cache_toMQ_deqReq_dummy2_2$Q_OUT;
  // ports of submodule cache_toMQ_enqReq_dummy2_0
  wire cache_toMQ_enqReq_dummy2_0$D_IN, cache_toMQ_enqReq_dummy2_0$EN;
  // ports of submodule cache_toMQ_enqReq_dummy2_1
  wire cache_toMQ_enqReq_dummy2_1$D_IN, cache_toMQ_enqReq_dummy2_1$EN;
  // ports of submodule cache_toMQ_enqReq_dummy2_2
  wire cache_toMQ_enqReq_dummy2_2$D_IN,
       cache_toMQ_enqReq_dummy2_2$EN,
       cache_toMQ_enqReq_dummy2_2$Q_OUT;
  // ports of submodule perfReqQ_clearReq_dummy2_0
  wire perfReqQ_clearReq_dummy2_0$D_IN, perfReqQ_clearReq_dummy2_0$EN;
  // ports of submodule perfReqQ_clearReq_dummy2_1
  wire perfReqQ_clearReq_dummy2_1$D_IN,
       perfReqQ_clearReq_dummy2_1$EN,
       perfReqQ_clearReq_dummy2_1$Q_OUT;
  // ports of submodule perfReqQ_deqReq_dummy2_0
  wire perfReqQ_deqReq_dummy2_0$D_IN, perfReqQ_deqReq_dummy2_0$EN;
  // ports of submodule perfReqQ_deqReq_dummy2_1
  wire perfReqQ_deqReq_dummy2_1$D_IN, perfReqQ_deqReq_dummy2_1$EN;
  // ports of submodule perfReqQ_deqReq_dummy2_2
  wire perfReqQ_deqReq_dummy2_2$D_IN,
       perfReqQ_deqReq_dummy2_2$EN,
       perfReqQ_deqReq_dummy2_2$Q_OUT;
  // ports of submodule perfReqQ_enqReq_dummy2_0
  wire perfReqQ_enqReq_dummy2_0$D_IN, perfReqQ_enqReq_dummy2_0$EN;
  // ports of submodule perfReqQ_enqReq_dummy2_1
  wire perfReqQ_enqReq_dummy2_1$D_IN, perfReqQ_enqReq_dummy2_1$EN;
  // ports of submodule perfReqQ_enqReq_dummy2_2
  wire perfReqQ_enqReq_dummy2_2$D_IN,
       perfReqQ_enqReq_dummy2_2$EN,
       perfReqQ_enqReq_dummy2_2$Q_OUT;
  // rule scheduling signals
  wire CAN_FIRE_RL_cache_cRqRetryIndexQ_canonicalize,
       CAN_FIRE_RL_cache_cRqRetryIndexQ_clearReq_canon,
       CAN_FIRE_RL_cache_cRqRetryIndexQ_deqReq_canon,
       CAN_FIRE_RL_cache_cRqRetryIndexQ_enqReq_canon,
       CAN_FIRE_RL_cache_cRqTransfer_new_child,
       CAN_FIRE_RL_cache_cRqTransfer_new_dma,
       CAN_FIRE_RL_cache_cRqTransfer_retry,
       CAN_FIRE_RL_cache_cRsTransfer,
       CAN_FIRE_RL_cache_mRsDeq_nonRefill,
       CAN_FIRE_RL_cache_mRsTransfer,
       CAN_FIRE_RL_cache_mergeRsLdToDmaIndexQ_mRsDeq,
       CAN_FIRE_RL_cache_mergeRsLdToDmaIndexQ_pipelineResp,
       CAN_FIRE_RL_cache_mergeRsStToDmaIndexQ_pipelineResp,
       CAN_FIRE_RL_cache_mergeRsStToDmaIndexQ_sendToM,
       CAN_FIRE_RL_cache_pipelineResp_cRq,
       CAN_FIRE_RL_cache_pipelineResp_cRs,
       CAN_FIRE_RL_cache_pipelineResp_mRs,
       CAN_FIRE_RL_cache_rqFromCQ_canonicalize,
       CAN_FIRE_RL_cache_rqFromCQ_clearReq_canon,
       CAN_FIRE_RL_cache_rqFromCQ_deqReq_canon,
       CAN_FIRE_RL_cache_rqFromCQ_enqReq_canon,
       CAN_FIRE_RL_cache_rqFromDmaQ_canonicalize,
       CAN_FIRE_RL_cache_rqFromDmaQ_clearReq_canon,
       CAN_FIRE_RL_cache_rqFromDmaQ_deqReq_canon,
       CAN_FIRE_RL_cache_rqFromDmaQ_enqReq_canon,
       CAN_FIRE_RL_cache_rsFromCQ_canonicalize,
       CAN_FIRE_RL_cache_rsFromCQ_clearReq_canon,
       CAN_FIRE_RL_cache_rsFromCQ_deqReq_canon,
       CAN_FIRE_RL_cache_rsFromCQ_enqReq_canon,
       CAN_FIRE_RL_cache_rsFromMQ_canonicalize,
       CAN_FIRE_RL_cache_rsFromMQ_clearReq_canon,
       CAN_FIRE_RL_cache_rsFromMQ_deqReq_canon,
       CAN_FIRE_RL_cache_rsFromMQ_enqReq_canon,
       CAN_FIRE_RL_cache_rsLdToDmaQ_canonicalize,
       CAN_FIRE_RL_cache_rsLdToDmaQ_clearReq_canon,
       CAN_FIRE_RL_cache_rsLdToDmaQ_deqReq_canon,
       CAN_FIRE_RL_cache_rsLdToDmaQ_enqReq_canon,
       CAN_FIRE_RL_cache_rsStToDmaQ_canonicalize,
       CAN_FIRE_RL_cache_rsStToDmaQ_clearReq_canon,
       CAN_FIRE_RL_cache_rsStToDmaQ_deqReq_canon,
       CAN_FIRE_RL_cache_rsStToDmaQ_enqReq_canon,
       CAN_FIRE_RL_cache_rsToCIndexQ_canonicalize,
       CAN_FIRE_RL_cache_rsToCIndexQ_clearReq_canon,
       CAN_FIRE_RL_cache_rsToCIndexQ_deqReq_canon,
       CAN_FIRE_RL_cache_rsToCIndexQ_enqReq_canon,
       CAN_FIRE_RL_cache_sendRqToC,
       CAN_FIRE_RL_cache_sendRsLdToDma,
       CAN_FIRE_RL_cache_sendRsStToDma,
       CAN_FIRE_RL_cache_sendRsToC,
       CAN_FIRE_RL_cache_sendToM,
       CAN_FIRE_RL_cache_toCQ_canonicalize,
       CAN_FIRE_RL_cache_toCQ_clearReq_canon,
       CAN_FIRE_RL_cache_toCQ_deqReq_canon,
       CAN_FIRE_RL_cache_toCQ_enqReq_canon,
       CAN_FIRE_RL_cache_toMQ_canonicalize,
       CAN_FIRE_RL_cache_toMQ_clearReq_canon,
       CAN_FIRE_RL_cache_toMQ_deqReq_canon,
       CAN_FIRE_RL_cache_toMQ_enqReq_canon,
       CAN_FIRE_RL_perfReqQ_canonicalize,
       CAN_FIRE_RL_perfReqQ_clearReq_canon,
       CAN_FIRE_RL_perfReqQ_deqReq_canon,
       CAN_FIRE_RL_perfReqQ_enqReq_canon,
       CAN_FIRE_cRqStuck_get,
       CAN_FIRE_dma_memReq_enq,
       CAN_FIRE_dma_respLd_deq,
       CAN_FIRE_dma_respSt_deq,
       CAN_FIRE_perf_req,
       CAN_FIRE_perf_resp,
       CAN_FIRE_perf_setStatus,
       CAN_FIRE_to_child_rqFromC_enq,
       CAN_FIRE_to_child_rsFromC_enq,
       CAN_FIRE_to_child_toC_deq,
       CAN_FIRE_to_mem_rsFromM_enq,
       CAN_FIRE_to_mem_toM_deq,
       WILL_FIRE_RL_cache_cRqRetryIndexQ_canonicalize,
       WILL_FIRE_RL_cache_cRqRetryIndexQ_clearReq_canon,
       WILL_FIRE_RL_cache_cRqRetryIndexQ_deqReq_canon,
       WILL_FIRE_RL_cache_cRqRetryIndexQ_enqReq_canon,
       WILL_FIRE_RL_cache_cRqTransfer_new_child,
       WILL_FIRE_RL_cache_cRqTransfer_new_dma,
       WILL_FIRE_RL_cache_cRqTransfer_retry,
       WILL_FIRE_RL_cache_cRsTransfer,
       WILL_FIRE_RL_cache_mRsDeq_nonRefill,
       WILL_FIRE_RL_cache_mRsTransfer,
       WILL_FIRE_RL_cache_mergeRsLdToDmaIndexQ_mRsDeq,
       WILL_FIRE_RL_cache_mergeRsLdToDmaIndexQ_pipelineResp,
       WILL_FIRE_RL_cache_mergeRsStToDmaIndexQ_pipelineResp,
       WILL_FIRE_RL_cache_mergeRsStToDmaIndexQ_sendToM,
       WILL_FIRE_RL_cache_pipelineResp_cRq,
       WILL_FIRE_RL_cache_pipelineResp_cRs,
       WILL_FIRE_RL_cache_pipelineResp_mRs,
       WILL_FIRE_RL_cache_rqFromCQ_canonicalize,
       WILL_FIRE_RL_cache_rqFromCQ_clearReq_canon,
       WILL_FIRE_RL_cache_rqFromCQ_deqReq_canon,
       WILL_FIRE_RL_cache_rqFromCQ_enqReq_canon,
       WILL_FIRE_RL_cache_rqFromDmaQ_canonicalize,
       WILL_FIRE_RL_cache_rqFromDmaQ_clearReq_canon,
       WILL_FIRE_RL_cache_rqFromDmaQ_deqReq_canon,
       WILL_FIRE_RL_cache_rqFromDmaQ_enqReq_canon,
       WILL_FIRE_RL_cache_rsFromCQ_canonicalize,
       WILL_FIRE_RL_cache_rsFromCQ_clearReq_canon,
       WILL_FIRE_RL_cache_rsFromCQ_deqReq_canon,
       WILL_FIRE_RL_cache_rsFromCQ_enqReq_canon,
       WILL_FIRE_RL_cache_rsFromMQ_canonicalize,
       WILL_FIRE_RL_cache_rsFromMQ_clearReq_canon,
       WILL_FIRE_RL_cache_rsFromMQ_deqReq_canon,
       WILL_FIRE_RL_cache_rsFromMQ_enqReq_canon,
       WILL_FIRE_RL_cache_rsLdToDmaQ_canonicalize,
       WILL_FIRE_RL_cache_rsLdToDmaQ_clearReq_canon,
       WILL_FIRE_RL_cache_rsLdToDmaQ_deqReq_canon,
       WILL_FIRE_RL_cache_rsLdToDmaQ_enqReq_canon,
       WILL_FIRE_RL_cache_rsStToDmaQ_canonicalize,
       WILL_FIRE_RL_cache_rsStToDmaQ_clearReq_canon,
       WILL_FIRE_RL_cache_rsStToDmaQ_deqReq_canon,
       WILL_FIRE_RL_cache_rsStToDmaQ_enqReq_canon,
       WILL_FIRE_RL_cache_rsToCIndexQ_canonicalize,
       WILL_FIRE_RL_cache_rsToCIndexQ_clearReq_canon,
       WILL_FIRE_RL_cache_rsToCIndexQ_deqReq_canon,
       WILL_FIRE_RL_cache_rsToCIndexQ_enqReq_canon,
       WILL_FIRE_RL_cache_sendRqToC,
       WILL_FIRE_RL_cache_sendRsLdToDma,
       WILL_FIRE_RL_cache_sendRsStToDma,
       WILL_FIRE_RL_cache_sendRsToC,
       WILL_FIRE_RL_cache_sendToM,
       WILL_FIRE_RL_cache_toCQ_canonicalize,
       WILL_FIRE_RL_cache_toCQ_clearReq_canon,
       WILL_FIRE_RL_cache_toCQ_deqReq_canon,
       WILL_FIRE_RL_cache_toCQ_enqReq_canon,
       WILL_FIRE_RL_cache_toMQ_canonicalize,
       WILL_FIRE_RL_cache_toMQ_clearReq_canon,
       WILL_FIRE_RL_cache_toMQ_deqReq_canon,
       WILL_FIRE_RL_cache_toMQ_enqReq_canon,
       WILL_FIRE_RL_perfReqQ_canonicalize,
       WILL_FIRE_RL_perfReqQ_clearReq_canon,
       WILL_FIRE_RL_perfReqQ_deqReq_canon,
       WILL_FIRE_RL_perfReqQ_enqReq_canon,
       WILL_FIRE_cRqStuck_get,
       WILL_FIRE_dma_memReq_enq,
       WILL_FIRE_dma_respLd_deq,
       WILL_FIRE_dma_respSt_deq,
       WILL_FIRE_perf_req,
       WILL_FIRE_perf_resp,
       WILL_FIRE_perf_setStatus,
       WILL_FIRE_to_child_rqFromC_enq,
       WILL_FIRE_to_child_rsFromC_enq,
       WILL_FIRE_to_child_toC_deq,
       WILL_FIRE_to_mem_rsFromM_enq,
       WILL_FIRE_to_mem_toM_deq;
  // inputs to muxes for submodule ports
  reg [3 : 0] MUX_cache_cRqMshr$sendRsToDmaC_getData_1__VAL_2,
	      MUX_cache_cRqMshr$transfer_getRq_1__VAL_2;
  wire [585 : 0] MUX_cache_toCQ_enqReq_lat_0$wset_1__VAL_1,
		 MUX_cache_toCQ_enqReq_lat_0$wset_1__VAL_2;
  wire [583 : 0] MUX_cache_pipeline$send_1__VAL_1,
		 MUX_cache_pipeline$send_1__VAL_2,
		 MUX_cache_pipeline$send_1__VAL_3,
		 MUX_cache_pipeline$send_1__VAL_4,
		 MUX_cache_pipeline$send_1__VAL_5;
  wire [573 : 0] MUX_cache_pipeline$deqWrite_2__VAL_1,
		 MUX_cache_pipeline$deqWrite_2__VAL_2,
		 MUX_cache_pipeline$deqWrite_2__VAL_3;
  wire [512 : 0] MUX_cache_cRqMshr$pipelineResp_setData_2__VAL_1,
		 MUX_cache_cRqMshr$pipelineResp_setData_2__VAL_2,
		 MUX_cache_cRqMshr$pipelineResp_setData_2__VAL_3,
		 MUX_cache_cRqMshr$transfer_getEmptyEntryInit_2__VAL_2;
  wire [151 : 0] MUX_cache_cRqMshr$transfer_getEmptyEntryInit_1__VAL_1,
		 MUX_cache_cRqMshr$transfer_getEmptyEntryInit_1__VAL_2;
  wire [64 : 0] MUX_cache_cRqMshr$pipelineResp_setStateSlot_3__VAL_1,
		MUX_cache_cRqMshr$pipelineResp_setStateSlot_3__VAL_2;
  wire [6 : 0] MUX_cache_rsToCIndexQ_enqReq_lat_0$wset_1__VAL_1,
	       MUX_cache_rsToCIndexQ_enqReq_lat_0$wset_1__VAL_2,
	       MUX_cache_rsToCIndexQ_enqReq_lat_0$wset_1__VAL_3;
  wire [5 : 0] MUX_cache_toMInfoQ$enq_1__VAL_1,
	       MUX_cache_toMInfoQ$enq_1__VAL_2;
  wire [4 : 0] MUX_cache_cRqRetryIndexQ_enqReq_lat_0$wset_1__VAL_1,
	       MUX_cache_cRqRetryIndexQ_enqReq_lat_0$wset_1__VAL_2,
	       MUX_cache_pipeline$deqWrite_1__VAL_2,
	       MUX_cache_pipeline$deqWrite_1__VAL_3;
  wire [2 : 0] MUX_cache_cRqMshr$pipelineResp_setStateSlot_2__VAL_1,
	       MUX_cache_cRqMshr$pipelineResp_setStateSlot_2__VAL_2;
  wire MUX_cache_cRqMshr$pipelineResp_setData_1__SEL_1,
       MUX_cache_cRqMshr$pipelineResp_setData_1__SEL_2,
       MUX_cache_cRqMshr$pipelineResp_setStateSlot_1__SEL_1,
       MUX_cache_cRqRetryIndexQ_enqReq_dummy2_0$write_1__SEL_1,
       MUX_cache_cRqRetryIndexQ_enqReq_dummy2_0$write_1__SEL_2,
       MUX_cache_pipeline$deqWrite_3__VAL_2,
       MUX_cache_pipeline$deqWrite_3__VAL_3,
       MUX_cache_rsLdToDmaIndexQ_pipelineResp$enq_1__SEL_1,
       MUX_cache_rsStToDmaIndexQ_pipelineResp$enq_1__SEL_1,
       MUX_cache_rsToCIndexQ_enqReq_dummy2_0$write_1__SEL_1,
       MUX_cache_rsToCIndexQ_enqReq_dummy2_0$write_1__SEL_2,
       MUX_cache_toMInfoQ$enq_1__SEL_1;
  // remaining internal signals
  reg [63 : 0] CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q232,
	       CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q233,
	       CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q267,
	       CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q91,
	       CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q92,
	       CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q93,
	       CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q98,
	       CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q99,
	       CASE_cache_rsFromCQ_deqP_0_cache_rsFromCQ_data_ETC__q236,
	       CASE_cache_rsFromCQ_deqP_0_cache_rsFromCQ_data_ETC__q237,
	       CASE_cache_rsFromCQ_deqP_0_cache_rsFromCQ_data_ETC__q243,
	       CASE_cache_rsFromCQ_deqP_0_cache_rsFromCQ_data_ETC__q69,
	       CASE_cache_rsFromCQ_deqP_0_cache_rsFromCQ_data_ETC__q70,
	       CASE_cache_rsFromCQ_deqP_0_cache_rsFromCQ_data_ETC__q71,
	       CASE_cache_rsFromCQ_deqP_0_cache_rsFromCQ_data_ETC__q72,
	       CASE_cache_rsFromCQ_deqP_0_cache_rsFromCQ_data_ETC__q75,
	       CASE_cache_rsFromCQ_deqP_0_cache_rsFromCQ_data_ETC__q76,
	       CASE_cache_rsFromMQ_deqP_0_cache_rsFromMQ_data_ETC__q1,
	       CASE_cache_rsFromMQ_deqP_0_cache_rsFromMQ_data_ETC__q2,
	       CASE_cache_rsFromMQ_deqP_0_cache_rsFromMQ_data_ETC__q226,
	       CASE_cache_rsFromMQ_deqP_0_cache_rsFromMQ_data_ETC__q227,
	       CASE_cache_rsFromMQ_deqP_0_cache_rsFromMQ_data_ETC__q3,
	       CASE_cache_rsFromMQ_deqP_0_cache_rsFromMQ_data_ETC__q4,
	       CASE_cache_rsFromMQ_deqP_0_cache_rsFromMQ_data_ETC__q73,
	       CASE_cache_rsFromMQ_deqP_0_cache_rsFromMQ_data_ETC__q74,
	       CASE_cache_rsLdToDmaQ_deqP_0_cache_rsLdToDmaQ__ETC__q257,
	       CASE_cache_rsLdToDmaQ_deqP_0_cache_rsLdToDmaQ__ETC__q258,
	       CASE_cache_rsLdToDmaQ_deqP_0_cache_rsLdToDmaQ__ETC__q259,
	       CASE_cache_rsLdToDmaQ_deqP_0_cache_rsLdToDmaQ__ETC__q85,
	       CASE_cache_rsLdToDmaQ_deqP_0_cache_rsLdToDmaQ__ETC__q86,
	       CASE_cache_rsLdToDmaQ_deqP_0_cache_rsLdToDmaQ__ETC__q87,
	       CASE_cache_rsLdToDmaQ_deqP_0_cache_rsLdToDmaQ__ETC__q96,
	       CASE_cache_rsLdToDmaQ_deqP_0_cache_rsLdToDmaQ__ETC__q97,
	       CASE_cache_toCQ_deqP_0_cache_toCQ_data_0_BITS__ETC__q234,
	       CASE_cache_toCQ_deqP_0_cache_toCQ_data_0_BITS__ETC__q235,
	       CASE_cache_toCQ_deqP_0_cache_toCQ_data_0_BITS__ETC__q239,
	       CASE_cache_toCQ_deqP_0_cache_toCQ_data_0_BITS__ETC__q247,
	       CASE_cache_toCQ_deqP_0_cache_toCQ_data_0_BITS__ETC__q249,
	       CASE_cache_toCQ_deqP_0_cache_toCQ_data_0_BITS__ETC__q88,
	       CASE_cache_toCQ_deqP_0_cache_toCQ_data_0_BITS__ETC__q89,
	       CASE_cache_toCQ_deqP_0_cache_toCQ_data_0_BITS__ETC__q90,
	       CASE_cache_toCQ_deqP_0_cache_toCQ_data_0_BITS__ETC__q94,
	       CASE_cache_toCQ_deqP_0_cache_toCQ_data_0_BITS__ETC__q95,
	       CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BITS__ETC__q220,
	       CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BITS__ETC__q221,
	       CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BITS__ETC__q222,
	       CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BITS__ETC__q223,
	       CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BITS__ETC__q224,
	       CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BITS__ETC__q225,
	       CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BITS__ETC__q245,
	       CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BITS__ETC__q246,
	       CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BITS__ETC__q251,
	       CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BITS__ETC__q252,
	       addr__h257616,
	       addr__h273361;
  reg [15 : 0] CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q266,
	       x__h456399;
  reg [3 : 0] x__h248737, x__h456804;
  reg [2 : 0] x__h257564, x__h445950;
  reg [1 : 0] CASE_cache_cRqMshrpipelineResp_getRq_BITS_82__ETC__q79,
	      CASE_cache_pipelinefirst_BITS_580_TO_579_0_ca_ETC__q84,
	      CASE_cache_rqFromCQ_deqP_0_cache_rqFromCQ_data_ETC__q230,
	      CASE_cache_rqFromCQ_deqP_0_cache_rqFromCQ_data_ETC__q265,
	      CASE_cache_rsFromCQ_deqP_0_cache_rsFromCQ_data_ETC__q244,
	      CASE_cache_toCQ_deqP_0_cache_toCQ_data_0_BITS__ETC__q248,
	      CASE_cache_toCQ_deqP_0_cache_toCQ_data_0_BITS__ETC__q250,
	      SEL_ARR_IF_cache_cRqMshr_sendRqToC_getSlot_IF__ETC___d2522,
	      SEL_ARR_cache_pipeline_first__581_BITS_519_TO__ETC___d3403,
	      SEL_ARR_cache_rsToCIndexQ_data_0_391_BITS_1_TO_ETC___d2445,
	      x__h249082,
	      x__h275130,
	      x__h444361,
	      x__h444405;
  reg CASE_cache_pipelineunguard_first_BITS_584_TO__ETC__q77,
      CASE_cache_rqFromCQ_deqP_0_cache_rqFromCQ_data_ETC__q231,
      CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q10,
      CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q11,
      CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q12,
      CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q13,
      CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q14,
      CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q15,
      CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q16,
      CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q17,
      CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q18,
      CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q19,
      CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q20,
      CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q21,
      CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q22,
      CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q23,
      CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q24,
      CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q25,
      CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q26,
      CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q27,
      CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q28,
      CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q29,
      CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q30,
      CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q31,
      CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q32,
      CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q33,
      CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q34,
      CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q35,
      CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q36,
      CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q37,
      CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q38,
      CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q39,
      CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q40,
      CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q41,
      CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q42,
      CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q43,
      CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q44,
      CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q45,
      CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q46,
      CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q47,
      CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q48,
      CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q49,
      CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q5,
      CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q50,
      CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q51,
      CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q52,
      CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q53,
      CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q54,
      CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q55,
      CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q56,
      CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q57,
      CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q58,
      CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q59,
      CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q6,
      CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q60,
      CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q61,
      CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q62,
      CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q63,
      CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q64,
      CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q65,
      CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q66,
      CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q67,
      CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q68,
      CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q7,
      CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q8,
      CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q9,
      CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q106,
      CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q107,
      CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q110,
      CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q111,
      CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q114,
      CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q115,
      CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q118,
      CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q119,
      CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q122,
      CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q123,
      CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q126,
      CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q127,
      CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q130,
      CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q131,
      CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q134,
      CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q135,
      CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q138,
      CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q139,
      CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q142,
      CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q143,
      CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q146,
      CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q147,
      CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q150,
      CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q151,
      CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q154,
      CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q155,
      CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q158,
      CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q159,
      CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q162,
      CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q163,
      CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q166,
      CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q167,
      CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q170,
      CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q171,
      CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q174,
      CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q175,
      CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q178,
      CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q179,
      CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q182,
      CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q183,
      CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q186,
      CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q187,
      CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q190,
      CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q191,
      CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q194,
      CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q195,
      CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q198,
      CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q199,
      CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q202,
      CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q203,
      CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q206,
      CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q207,
      CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q210,
      CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q211,
      CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q214,
      CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q215,
      CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q218,
      CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q219,
      CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q228,
      CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q229,
      CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q80,
      CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q81,
      CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q82,
      CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q83,
      CASE_cache_rsFromCQ_deqP_0_cache_rsFromCQ_data_ETC__q242,
      CASE_cache_rsFromMQ_deqP_0_NOT_cache_rsFromMQ__ETC__q263,
      CASE_cache_rsFromMQ_deqP_0_cache_rsFromMQ_data_ETC__q262,
      CASE_cache_toCQ_deqP_0_NOT_cache_toCQ_data_0_B_ETC__q255,
      CASE_cache_toCQ_deqP_0_cache_toCQ_data_0_BIT_5_ETC__q238,
      CASE_cache_toCQ_deqP_0_cache_toCQ_data_0_BIT_5_ETC__q256,
      CASE_cache_toMInfoQD_OUT_BITS_1_TO_0_0_NOT_ca_ETC__q264,
      CASE_cache_toMQ_deqP_0_NOT_cache_toMQ_data_0_B_ETC__q260,
      CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_4_ETC__q253,
      CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q100,
      CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q101,
      CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q102,
      CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q103,
      CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q104,
      CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q105,
      CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q108,
      CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q109,
      CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q112,
      CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q113,
      CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q116,
      CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q117,
      CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q120,
      CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q121,
      CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q124,
      CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q125,
      CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q128,
      CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q129,
      CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q132,
      CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q133,
      CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q136,
      CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q137,
      CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q140,
      CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q141,
      CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q144,
      CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q145,
      CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q148,
      CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q149,
      CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q152,
      CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q153,
      CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q156,
      CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q157,
      CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q160,
      CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q161,
      CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q164,
      CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q165,
      CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q168,
      CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q169,
      CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q172,
      CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q173,
      CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q176,
      CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q177,
      CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q180,
      CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q181,
      CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q184,
      CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q185,
      CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q188,
      CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q189,
      CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q192,
      CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q193,
      CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q196,
      CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q197,
      CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q200,
      CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q201,
      CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q204,
      CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q205,
      CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q208,
      CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q209,
      CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q212,
      CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q213,
      CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q216,
      CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q217,
      CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q240,
      CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q241,
      CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_6_ETC__q261,
      CASE_child13067_0_cache_cRqMshrsendRqToC_getS_ETC__q254,
      SEL_ARR_cache_cRqMshr_pipelineResp_getSlot_IF__ETC___d3431,
      SEL_ARR_cache_cRqMshr_pipelineResp_getSlot_IF__ETC___d3446;
  wire [641 : 0] IF_cache_doLdAfterReplace_007_THEN_2_CONCAT_DO_ETC___d2016;
  wire [639 : 0] DONTCARE_CONCAT_SEL_ARR_cache_toMQ_data_0_050__ETC___d4073,
		 IF_SEL_ARR_NOT_cache_toMQ_data_0_050_BIT_640_0_ETC___d4404,
		 IF_cache_toMQ_enqReq_dummy2_2_read__54_AND_IF__ETC___d703,
		 SEL_ARR_cache_toMQ_data_0_050_BITS_639_TO_576__ETC___d4402;
  wire [583 : 0] DONTCARE_CONCAT_SEL_ARR_cache_toCQ_data_0_917__ETC___d3940,
		 IF_SEL_ARR_NOT_cache_toCQ_data_0_917_BIT_584_9_ETC___d4000,
		 IF_cache_toCQ_enqReq_dummy2_2_read__53_AND_IF__ETC___d302,
		 SEL_ARR_cache_toCQ_data_0_917_BITS_583_TO_520__ETC___d3998;
  wire [580 : 0] SEL_ARR_cache_rsFromCQ_data_0_855_BITS_580_TO__ETC___d1910;
  wire [573 : 0] IF_NOT_cache_pipeline_first__581_BITS_525_TO_5_ETC___d2999,
		 IF_cache_cRqMshr_pipelineResp_searchEndOfChain_ETC___d3012,
		 IF_cache_pipeline_first__581_BITS_525_TO_524_6_ETC___d3010,
		 IF_cache_pipeline_first__581_BIT_512_308_THEN__ETC___d3660,
		 cache_cRqMshr_pipelineResp_getRq_IF_cache_pipe_ETC___d2995,
		 cache_cRqMshr_pipelineResp_getRq_IF_cache_pipe_ETC___d3658;
  wire [514 : 0] SEL_ARR_cache_rsFromCQ_data_0_855_BIT_514_865__ETC___d1909;
  wire [512 : 0] SEL_ARR_cache_toCQ_data_0_917_BIT_515_953_cach_ETC___d3992;
  wire [511 : 0] IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2991,
		 IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3656,
		 IF_cache_pipeline_first__581_BITS_519_TO_518_5_ETC___d2993,
		 SEL_ARR_cache_rsFromCQ_data_0_855_BITS_513_TO__ETC___d1904,
		 SEL_ARR_cache_rsFromMQ_data_0_914_BITS_516_TO__ETC___d1966,
		 SEL_ARR_cache_toMQ_data_0_050_BITS_511_TO_448__ETC___d4401;
  wire [447 : 0] SEL_ARR_cache_rqFromDmaQ_data_0_129_BITS_527_T_ETC___d1845,
		 SEL_ARR_cache_rsLdToDmaQ_data_0_004_BITS_527_T_ETC___d4036,
		 SEL_ARR_cache_toCQ_data_0_917_BITS_514_TO_451__ETC___d3987;
  wire [383 : 0] IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2916,
		 IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3613,
		 SEL_ARR_cache_rsFromCQ_data_0_855_BITS_513_TO__ETC___d1895,
		 SEL_ARR_cache_rsFromMQ_data_0_914_BITS_516_TO__ETC___d1957,
		 SEL_ARR_cache_toMQ_data_0_050_BITS_511_TO_448__ETC___d4392;
  wire [319 : 0] SEL_ARR_cache_rqFromDmaQ_data_0_129_BITS_527_T_ETC___d1836,
		 SEL_ARR_cache_rsLdToDmaQ_data_0_004_BITS_527_T_ETC___d4027,
		 SEL_ARR_cache_toCQ_data_0_917_BITS_514_TO_451__ETC___d3978;
  wire [255 : 0] IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2844,
		 IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3573,
		 SEL_ARR_cache_rsFromCQ_data_0_855_BITS_513_TO__ETC___d1886,
		 SEL_ARR_cache_rsFromMQ_data_0_914_BITS_516_TO__ETC___d1948,
		 SEL_ARR_cache_toMQ_data_0_050_BITS_511_TO_448__ETC___d4383;
  wire [191 : 0] SEL_ARR_cache_rqFromDmaQ_data_0_129_BITS_527_T_ETC___d1827,
		 SEL_ARR_cache_rsLdToDmaQ_data_0_004_BITS_527_T_ETC___d4018,
		 SEL_ARR_cache_toCQ_data_0_917_BITS_514_TO_451__ETC___d3969;
  wire [127 : 0] IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2772,
		 IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3533;
  wire [85 : 0] SEL_ARR_cache_rqFromCQ_data_0_090_BITS_7_TO_6__ETC___d1118;
  wire [64 : 0] IF_IF_SEL_ARR_cache_pipeline_first__581_BITS_5_ETC___d3709,
		IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3078,
		IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3096,
		IF_cache_pipeline_first__581_BITS_525_TO_524_6_ETC___d3095,
		cache_cRqMshr_pipelineResp_getSlot_IF_cache_pi_ETC___d3754;
  wire [63 : 0] IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2808,
		IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2880,
		IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2952,
		IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3553,
		IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3593,
		IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3633,
		SEL_ARR_cache_rqFromDmaQ_data_0_129_BIT_591_57_ETC___d1806,
		SEL_ARR_cache_toMQ_data_0_050_BIT_575_078_cach_ETC___d4365,
		addr__h288271,
		cache_cRqMshrpipelineResp_getData_BITS_63_TO_0__q78,
		rqAddr__h313360;
  wire [61 : 0] SEL_ARR_cache_rqFromDmaQ_data_0_129_BIT_591_57_ETC___d1801,
		SEL_ARR_cache_toMQ_data_0_050_BIT_575_078_cach_ETC___d4356;
  wire [59 : 0] SEL_ARR_cache_rqFromDmaQ_data_0_129_BIT_591_57_ETC___d1796,
		SEL_ARR_cache_toMQ_data_0_050_BIT_575_078_cach_ETC___d4347;
  wire [57 : 0] SEL_ARR_cache_rqFromDmaQ_data_0_129_BIT_591_57_ETC___d1791,
		SEL_ARR_cache_toMQ_data_0_050_BIT_575_078_cach_ETC___d4338;
  wire [55 : 0] IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2732,
		IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2767,
		IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2839,
		IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2911,
		IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2986,
		IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3511,
		IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3530,
		IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3570,
		IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3610,
		IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3653,
		SEL_ARR_cache_rqFromDmaQ_data_0_129_BIT_591_57_ETC___d1786,
		SEL_ARR_cache_toMQ_data_0_050_BIT_575_078_cach_ETC___d4329;
  wire [53 : 0] SEL_ARR_cache_rqFromDmaQ_data_0_129_BIT_591_57_ETC___d1781,
		SEL_ARR_cache_toMQ_data_0_050_BIT_575_078_cach_ETC___d4320;
  wire [51 : 0] SEL_ARR_cache_rqFromDmaQ_data_0_129_BIT_591_57_ETC___d1776,
		SEL_ARR_cache_toMQ_data_0_050_BIT_575_078_cach_ETC___d4311;
  wire [49 : 0] SEL_ARR_cache_rqFromDmaQ_data_0_129_BIT_591_57_ETC___d1771,
		SEL_ARR_cache_toMQ_data_0_050_BIT_575_078_cach_ETC___d4302;
  wire [47 : 0] IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2799,
		IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2871,
		IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2943,
		IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3548,
		IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3588,
		IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3628,
		SEL_ARR_cache_rqFromDmaQ_data_0_129_BIT_591_57_ETC___d1766,
		SEL_ARR_cache_toMQ_data_0_050_BIT_575_078_cach_ETC___d4293;
  wire [45 : 0] SEL_ARR_cache_rqFromDmaQ_data_0_129_BIT_591_57_ETC___d1761,
		SEL_ARR_cache_toMQ_data_0_050_BIT_575_078_cach_ETC___d4284;
  wire [43 : 0] SEL_ARR_cache_rqFromDmaQ_data_0_129_BIT_591_57_ETC___d1756,
		SEL_ARR_cache_toMQ_data_0_050_BIT_575_078_cach_ETC___d4275;
  wire [41 : 0] SEL_ARR_cache_rqFromDmaQ_data_0_129_BIT_591_57_ETC___d1751,
		SEL_ARR_cache_toMQ_data_0_050_BIT_575_078_cach_ETC___d4266;
  wire [39 : 0] IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2723,
		IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2758,
		IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2830,
		IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2902,
		IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2977,
		IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3506,
		IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3525,
		IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3565,
		IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3605,
		IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3648,
		SEL_ARR_cache_rqFromDmaQ_data_0_129_BIT_591_57_ETC___d1746,
		SEL_ARR_cache_toMQ_data_0_050_BIT_575_078_cach_ETC___d4257;
  wire [37 : 0] SEL_ARR_cache_rqFromDmaQ_data_0_129_BIT_591_57_ETC___d1741,
		SEL_ARR_cache_toMQ_data_0_050_BIT_575_078_cach_ETC___d4248;
  wire [35 : 0] SEL_ARR_cache_rqFromDmaQ_data_0_129_BIT_591_57_ETC___d1736,
		SEL_ARR_cache_toMQ_data_0_050_BIT_575_078_cach_ETC___d4239;
  wire [33 : 0] SEL_ARR_cache_rqFromDmaQ_data_0_129_BIT_591_57_ETC___d1731,
		SEL_ARR_cache_toMQ_data_0_050_BIT_575_078_cach_ETC___d4230;
  wire [31 : 0] IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2790,
		IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2862,
		IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2934,
		SEL_ARR_cache_rqFromDmaQ_data_0_129_BIT_591_57_ETC___d1726,
		SEL_ARR_cache_toMQ_data_0_050_BIT_575_078_cach_ETC___d4221;
  wire [29 : 0] SEL_ARR_cache_rqFromDmaQ_data_0_129_BIT_591_57_ETC___d1721,
		SEL_ARR_cache_toMQ_data_0_050_BIT_575_078_cach_ETC___d4212;
  wire [27 : 0] SEL_ARR_cache_rqFromDmaQ_data_0_129_BIT_591_57_ETC___d1716,
		SEL_ARR_cache_toMQ_data_0_050_BIT_575_078_cach_ETC___d4203;
  wire [25 : 0] SEL_ARR_cache_rqFromDmaQ_data_0_129_BIT_591_57_ETC___d1711,
		SEL_ARR_cache_toMQ_data_0_050_BIT_575_078_cach_ETC___d4194;
  wire [23 : 0] IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2714,
		IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2749,
		IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2821,
		IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2893,
		IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2968,
		SEL_ARR_cache_rqFromDmaQ_data_0_129_BIT_591_57_ETC___d1706,
		SEL_ARR_cache_toMQ_data_0_050_BIT_575_078_cach_ETC___d4185;
  wire [21 : 0] SEL_ARR_cache_rqFromDmaQ_data_0_129_BIT_591_57_ETC___d1701,
		SEL_ARR_cache_toMQ_data_0_050_BIT_575_078_cach_ETC___d4176;
  wire [19 : 0] SEL_ARR_cache_rqFromDmaQ_data_0_129_BIT_591_57_ETC___d1696,
		SEL_ARR_cache_toMQ_data_0_050_BIT_575_078_cach_ETC___d4167;
  wire [17 : 0] SEL_ARR_cache_rqFromDmaQ_data_0_129_BIT_591_57_ETC___d1691,
		SEL_ARR_cache_toMQ_data_0_050_BIT_575_078_cach_ETC___d4158;
  wire [15 : 0] SEL_ARR_cache_rqFromDmaQ_data_0_129_BIT_591_57_ETC___d1686,
		SEL_ARR_cache_toMQ_data_0_050_BIT_575_078_cach_ETC___d4149;
  wire [13 : 0] IF_IF_cache_cRqMshr_pipelineResp_getRq_IF_cach_ETC___d2699,
		IF_IF_cache_cRqMshr_pipelineResp_getRq_IF_cach_ETC___d3397,
		IF_NOT_cache_pipeline_first__581_BITS_525_TO_5_ETC___d3000,
		IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3493,
		IF_cache_pipeline_first__581_BITS_519_TO_518_5_ETC___d2693,
		SEL_ARR_cache_rqFromDmaQ_data_0_129_BIT_591_57_ETC___d1681,
		SEL_ARR_cache_toMQ_data_0_050_BIT_575_078_cach_ETC___d4140;
  wire [12 : 0] _0_CONCAT_IF_cache_pipeline_first__581_BITS_523_ETC___d3043;
  wire [11 : 0] SEL_ARR_cache_rqFromDmaQ_data_0_129_BIT_591_57_ETC___d1676,
		SEL_ARR_cache_toMQ_data_0_050_BIT_575_078_cach_ETC___d4131;
  wire [9 : 0] SEL_ARR_cache_rqFromDmaQ_data_0_129_BIT_591_57_ETC___d1671,
	       SEL_ARR_cache_toMQ_data_0_050_BIT_575_078_cach_ETC___d4122;
  wire [7 : 0] IF_SEL_ARR_cache_pipeline_first__581_BITS_519__ETC___d3694,
	       IF_cache_pipeline_first__581_BITS_523_TO_522_6_ETC___d3041,
	       SEL_ARR_cache_rqFromDmaQ_data_0_129_BIT_591_57_ETC___d1666,
	       SEL_ARR_cache_toMQ_data_0_050_BIT_575_078_cach_ETC___d4113;
  wire [5 : 0] IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2697,
	       IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3396,
	       SEL_ARR_cache_rqFromDmaQ_data_0_129_BIT_591_57_ETC___d1661,
	       SEL_ARR_cache_toMQ_data_0_050_BIT_575_078_cach_ETC___d4104;
  wire [4 : 0] IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2678,
	       IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2683,
	       IF_cache_pipeline_first__581_BITS_519_TO_518_5_ETC___d2676,
	       IF_cache_pipeline_first__581_BITS_525_TO_524_6_ETC___d2682,
	       IF_cache_pipeline_first__581_BIT_512_308_THEN__ETC___d3486;
  wire [3 : 0] SEL_ARR_cache_rqFromDmaQ_data_0_129_BIT_591_57_ETC___d1656,
	       SEL_ARR_cache_toMQ_data_0_050_BIT_575_078_cach_ETC___d4095,
	       _theResult_____2__h234513,
	       _theResult_____2__h245988,
	       next_deqP___1__h234850,
	       next_deqP___1__h246325,
	       pipeOutCRqIdx__h314276,
	       v__h232953,
	       v__h233236,
	       v__h242396,
	       v__h242679;
  wire [2 : 0] IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3027,
	       IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3033,
	       IF_cache_pipeline_first__581_BITS_519_TO_518_5_ETC___d3025,
	       IF_cache_pipeline_first__581_BITS_525_TO_524_6_ETC___d3032;
  wire [1 : 0] IF_IF_cache_pipeline_first__581_BITS_584_TO_58_ETC___d3672,
	       IF_IF_cache_pipeline_first__581_BITS_584_TO_58_ETC___d3684,
	       IF_IF_cache_pipeline_first__581_BITS_584_TO_58_ETC___d3697,
	       IF_NOT_SEL_ARR_NOT_cache_rqFromDmaQ_data_0_129_ETC___d1646,
	       IF_NOT_cache_cRqMshr_pipelineResp_getRq_IF_cac_ETC___d3054,
	       IF_NOT_cache_cRqMshr_pipelineResp_getRq_IF_cac_ETC___d3063,
	       IF_NOT_cache_cRqMshr_pipelineResp_getRq_IF_cac_ETC___d3073,
	       IF_SEL_ARR_cache_cRqMshr_pipelineResp_getSlot__ETC___d3712,
	       IF_SEL_ARR_cache_cRqMshr_pipelineResp_getSlot__ETC___d3713,
	       IF_SEL_ARR_cache_cRqMshr_pipelineResp_getSlot__ETC___d3726,
	       IF_SEL_ARR_cache_cRqMshr_pipelineResp_getSlot__ETC___d3727,
	       IF_SEL_ARR_cache_cRqMshr_pipelineResp_getSlot__ETC___d3741,
	       IF_SEL_ARR_cache_cRqMshr_pipelineResp_getSlot__ETC___d3742,
	       IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2597,
	       IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2686,
	       IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3048,
	       IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3057,
	       IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3067,
	       IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3173,
	       IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3388,
	       IF_cache_pipeline_first__581_BITS_525_TO_524_6_ETC___d3171,
	       child__h313067;
  wire IF_IF_cache_cRqMshr_pipelineResp_getRq_IF_cach_ETC___d2635,
       IF_NOT_cache_pipeline_first__581_BITS_525_TO_5_ETC___d2654,
       IF_NOT_cache_pipeline_first__581_BITS_525_TO_5_ETC___d2657,
       IF_SEL_ARR_IF_cache_cRqMshr_pipelineResp_getSl_ETC___d3481,
       IF_SEL_ARR_IF_cache_cRqMshr_pipelineResp_getSl_ETC___d3482,
       IF_SEL_ARR_cache_cRqMshr_pipelineResp_getSlot__ETC___d3454,
       IF_SEL_ARR_cache_cRqMshr_pipelineResp_getSlot__ETC___d3455,
       IF_SEL_ARR_cache_cRqMshr_pipelineResp_getSlot__ETC___d3458,
       IF_SEL_ARR_cache_cRqMshr_pipelineResp_getSlot__ETC___d3459,
       IF_SEL_ARR_cache_cRqMshr_pipelineResp_getSlot__ETC___d3462,
       IF_SEL_ARR_cache_cRqMshr_pipelineResp_getSlot__ETC___d3463,
       IF_SEL_ARR_cache_cRqMshr_pipelineResp_getSlot__ETC___d3484,
       IF_SEL_ARR_cache_cRqMshr_pipelineResp_getSlot__ETC___d3804,
       IF_SEL_ARR_cache_cRqMshr_pipelineResp_getSlot__ETC___d3814,
       IF_SEL_ARR_cache_cRqMshr_pipelineResp_getSlot__ETC___d3830,
       IF_SEL_ARR_cache_pipeline_first__581_BITS_519__ETC___d3417,
       IF_SEL_ARR_cache_pipeline_first__581_BITS_519__ETC___d3418,
       IF_SEL_ARR_cache_pipeline_first__581_BITS_519__ETC___d3488,
       IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2626,
       IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2627,
       IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3014,
       IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3022,
       IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3155,
       IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3156,
       IF_cache_cRqRetryIndexQ_deqReq_dummy2_2_read___ETC___d854,
       IF_cache_cRqRetryIndexQ_deqReq_lat_1_whas__11__ETC___d817,
       IF_cache_cRqRetryIndexQ_enqReq_lat_1_whas__01__ETC___d833,
       IF_cache_pipeline_RDY_first__579_AND_cache_cRq_ETC___d2613,
       IF_cache_pipeline_first__581_BITS_525_TO_524_6_ETC___d2667,
       IF_cache_pipeline_first__581_BIT_517_582_THEN__ETC___d3124,
       IF_cache_rqFromCQ_deqReq_dummy2_2_read__7_AND__ETC___d55,
       IF_cache_rqFromCQ_deqReq_lat_1_whas__3_THEN_ca_ETC___d19,
       IF_cache_rqFromCQ_enqReq_lat_1_whas_THEN_cache_ETC___d39,
       IF_cache_rqFromDmaQ_deqReq_dummy2_2_read__53_A_ETC___d361,
       IF_cache_rqFromDmaQ_deqReq_lat_1_whas__19_THEN_ETC___d325,
       IF_cache_rqFromDmaQ_enqReq_lat_1_whas__09_THEN_ETC___d345,
       IF_cache_rsFromCQ_deqReq_dummy2_2_read__39_AND_ETC___d147,
       IF_cache_rsFromCQ_deqReq_lat_1_whas__05_THEN_c_ETC___d111,
       IF_cache_rsFromCQ_enqReq_lat_1_whas__5_THEN_ca_ETC___d131,
       IF_cache_rsFromMQ_deqReq_dummy2_2_read__54_AND_ETC___d762,
       IF_cache_rsFromMQ_deqReq_lat_1_whas__20_THEN_c_ETC___d726,
       IF_cache_rsFromMQ_enqReq_lat_1_whas__10_THEN_c_ETC___d746,
       IF_cache_rsLdToDmaQ_deqReq_dummy2_2_read__44_A_ETC___d452,
       IF_cache_rsLdToDmaQ_deqReq_lat_1_whas__10_THEN_ETC___d416,
       IF_cache_rsLdToDmaQ_enqReq_lat_1_whas__00_THEN_ETC___d436,
       IF_cache_rsStToDmaQ_deqReq_dummy2_2_read__35_A_ETC___d543,
       IF_cache_rsStToDmaQ_deqReq_lat_1_whas__01_THEN_ETC___d507,
       IF_cache_rsStToDmaQ_enqReq_lat_1_whas__91_THEN_ETC___d527,
       IF_cache_rsToCIndexQ_deqReq_dummy2_2_read__64__ETC___d977,
       IF_cache_rsToCIndexQ_deqReq_lat_1_whas__34_THE_ETC___d940,
       IF_cache_rsToCIndexQ_enqReq_lat_1_whas__24_THE_ETC___d956,
       IF_cache_toCQ_deqReq_dummy2_2_read__61_AND_IF__ETC___d269,
       IF_cache_toCQ_deqReq_lat_1_whas__32_THEN_cache_ETC___d238,
       IF_cache_toCQ_enqReq_lat_1_whas__87_THEN_cache_ETC___d196,
       IF_cache_toMQ_deqReq_dummy2_2_read__62_AND_IF__ETC___d670,
       IF_cache_toMQ_deqReq_lat_1_whas__33_THEN_cache_ETC___d639,
       IF_cache_toMQ_enqReq_lat_1_whas__88_THEN_cache_ETC___d597,
       IF_perfReqQ_enqReq_lat_1_whas__839_THEN_perfRe_ETC___d3875,
       NOT_IF_cache_pipeline_first__581_BITS_584_TO_5_ETC___d3191,
       NOT_SEL_ARR_NOT_cache_rqFromDmaQ_data_0_129_BI_ETC___d1584,
       NOT_SEL_ARR_NOT_cache_rqFromDmaQ_data_0_129_BI_ETC___d1586,
       NOT_SEL_ARR_NOT_cache_rqFromDmaQ_data_0_129_BI_ETC___d1588,
       NOT_SEL_ARR_NOT_cache_rqFromDmaQ_data_0_129_BI_ETC___d1590,
       NOT_SEL_ARR_NOT_cache_rqFromDmaQ_data_0_129_BI_ETC___d1592,
       NOT_SEL_ARR_NOT_cache_rqFromDmaQ_data_0_129_BI_ETC___d1594,
       NOT_SEL_ARR_NOT_cache_rqFromDmaQ_data_0_129_BI_ETC___d1596,
       NOT_SEL_ARR_NOT_cache_rqFromDmaQ_data_0_129_BI_ETC___d1598,
       NOT_SEL_ARR_NOT_cache_rqFromDmaQ_data_0_129_BI_ETC___d1600,
       NOT_SEL_ARR_NOT_cache_rqFromDmaQ_data_0_129_BI_ETC___d1602,
       NOT_SEL_ARR_NOT_cache_rqFromDmaQ_data_0_129_BI_ETC___d1604,
       NOT_SEL_ARR_NOT_cache_rqFromDmaQ_data_0_129_BI_ETC___d1606,
       NOT_SEL_ARR_NOT_cache_rqFromDmaQ_data_0_129_BI_ETC___d1608,
       NOT_SEL_ARR_NOT_cache_rqFromDmaQ_data_0_129_BI_ETC___d1610,
       NOT_SEL_ARR_NOT_cache_rqFromDmaQ_data_0_129_BI_ETC___d1612,
       NOT_SEL_ARR_NOT_cache_rqFromDmaQ_data_0_129_BI_ETC___d1614,
       NOT_SEL_ARR_NOT_cache_rqFromDmaQ_data_0_129_BI_ETC___d1616,
       NOT_SEL_ARR_NOT_cache_rqFromDmaQ_data_0_129_BI_ETC___d1618,
       NOT_SEL_ARR_NOT_cache_rqFromDmaQ_data_0_129_BI_ETC___d1620,
       NOT_SEL_ARR_NOT_cache_rqFromDmaQ_data_0_129_BI_ETC___d1622,
       NOT_SEL_ARR_NOT_cache_rqFromDmaQ_data_0_129_BI_ETC___d1624,
       NOT_SEL_ARR_NOT_cache_rqFromDmaQ_data_0_129_BI_ETC___d1626,
       NOT_SEL_ARR_NOT_cache_rqFromDmaQ_data_0_129_BI_ETC___d1628,
       NOT_SEL_ARR_NOT_cache_rqFromDmaQ_data_0_129_BI_ETC___d1630,
       NOT_SEL_ARR_NOT_cache_rqFromDmaQ_data_0_129_BI_ETC___d1632,
       NOT_SEL_ARR_NOT_cache_rqFromDmaQ_data_0_129_BI_ETC___d1634,
       NOT_SEL_ARR_NOT_cache_rqFromDmaQ_data_0_129_BI_ETC___d1636,
       NOT_SEL_ARR_NOT_cache_rqFromDmaQ_data_0_129_BI_ETC___d1638,
       NOT_SEL_ARR_NOT_cache_rqFromDmaQ_data_0_129_BI_ETC___d1640,
       NOT_SEL_ARR_NOT_cache_rqFromDmaQ_data_0_129_BI_ETC___d1642,
       NOT_SEL_ARR_NOT_cache_rqFromDmaQ_data_0_129_BI_ETC___d1644,
       NOT_SEL_ARR_cache_cRqMshr_sendRqToC_getSlot_IF_ETC___d2508,
       NOT_cache_cRqMshr_pipelineResp_getRq_IF_cache__ETC___d3264,
       NOT_cache_cRqMshr_pipelineResp_getRq_IF_cache__ETC___d3290,
       NOT_cache_cRqMshr_pipelineResp_getRq_IF_cache__ETC___d3299,
       NOT_cache_cRqMshr_pipelineResp_getSlot_IF_cach_ETC___d3369,
       NOT_cache_cRqMshr_pipelineResp_searchEndOfChai_ETC___d3114,
       NOT_cache_cRqMshr_pipelineResp_searchEndOfChai_ETC___d3353,
       NOT_cache_cRqRetryIndexQ_clearReq_dummy2_1_rea_ETC___d853,
       NOT_cache_cRqRetryIndexQ_enqReq_dummy2_2_read__ETC___d876,
       NOT_cache_pipeline_first__581_BITS_516_TO_513__ETC___d2637,
       NOT_cache_pipeline_first__581_BITS_516_TO_513__ETC___d3798,
       NOT_cache_pipeline_first__581_BITS_519_TO_518__ETC___d3275,
       NOT_cache_pipeline_first__581_BITS_519_TO_518__ETC___d3281,
       NOT_cache_pipeline_first__581_BITS_525_TO_524__ETC___d3019,
       NOT_cache_pipeline_first__581_BIT_512_308_309__ETC___d3801,
       NOT_cache_pipeline_first__581_BIT_512_308_309__ETC___d3809,
       NOT_cache_pipeline_first__581_BIT_512_308_309__ETC___d3827,
       NOT_cache_pipeline_first__581_BIT_517_582_105__ETC___d3133,
       NOT_cache_pipeline_first__581_BIT_517_582_105__ETC___d3143,
       NOT_cache_pipeline_first__581_BIT_517_582_105__ETC___d3149,
       NOT_cache_pipeline_first__581_BIT_517_582_105__ETC___d3316,
       NOT_cache_pipeline_first__581_BIT_517_582_105__ETC___d3320,
       NOT_cache_pipeline_first__581_BIT_517_582_105__ETC___d3324,
       NOT_cache_pipeline_first__581_BIT_517_582_105__ETC___d3328,
       NOT_cache_pipeline_first__581_BIT_517_582_105__ETC___d3332,
       NOT_cache_pipeline_first__581_BIT_517_582_105__ETC___d3340,
       NOT_cache_pipeline_first__581_BIT_517_582_105__ETC___d3345,
       NOT_cache_pipeline_first__581_BIT_517_582_105__ETC___d3351,
       NOT_cache_pipeline_first__581_BIT_517_582_105__ETC___d3359,
       NOT_cache_rqFromCQ_clearReq_dummy2_1_read__8_9_ETC___d33,
       NOT_cache_rqFromCQ_enqReq_dummy2_2_read__4_9_O_ETC___d78,
       NOT_cache_rqFromDmaQ_clearReq_dummy2_1_read__3_ETC___d339,
       NOT_cache_rqFromDmaQ_enqReq_dummy2_2_read__40__ETC___d384,
       NOT_cache_rsFromCQ_clearReq_dummy2_1_read__20__ETC___d125,
       NOT_cache_rsFromCQ_enqReq_dummy2_2_read__26_61_ETC___d170,
       NOT_cache_rsFromMQ_clearReq_dummy2_1_read__35__ETC___d740,
       NOT_cache_rsFromMQ_enqReq_dummy2_2_read__41_76_ETC___d785,
       NOT_cache_rsLdToDmaQ_clearReq_dummy2_1_read__2_ETC___d430,
       NOT_cache_rsLdToDmaQ_enqReq_dummy2_2_read__31__ETC___d475,
       NOT_cache_rsStToDmaQ_clearReq_dummy2_1_read__1_ETC___d521,
       NOT_cache_rsStToDmaQ_enqReq_dummy2_2_read__22__ETC___d566,
       NOT_cache_rsToCIndexQ_clearReq_dummy2_1_read___ETC___d976,
       NOT_cache_rsToCIndexQ_enqReq_dummy2_2_read__51_ETC___d999,
       NOT_cache_toCQ_clearReq_dummy2_1_read__47_48_O_ETC___d252,
       NOT_cache_toCQ_enqReq_dummy2_2_read__53_83_OR__ETC___d292,
       NOT_cache_toMQ_clearReq_dummy2_1_read__48_49_O_ETC___d653,
       NOT_cache_toMQ_enqReq_dummy2_2_read__54_84_OR__ETC___d693,
       NOT_perfReqQ_clearReq_dummy2_1_read__864_865_O_ETC___d3869,
       NOT_perfReqQ_enqReq_dummy2_2_read__870_890_OR__ETC___d3900,
       SEL_ARR_IF_cache_cRqMshr_pipelineResp_getSlot__ETC___d3440,
       _0_OR_IF_SEL_ARR_cache_pipeline_first__581_BITS_ETC___d3423,
       _0_OR_NOT_CASE_IF_cache_pipeline_first__581_BIT_ETC___d3468,
       _0_OR_NOT_cache_pipeline_first__581_BITS_519_TO_ETC___d2614,
       _theResult_____2__h119142,
       _theResult_____2__h135235,
       _theResult_____2__h142737,
       _theResult_____2__h208521,
       _theResult_____2__h22297,
       _theResult_____2__h225016,
       _theResult_____2__h37990,
       _theResult_____2__h7215,
       cache_cRqMshr_pipelineResp_getRq_IF_cache_pipe_ETC___d3123,
       cache_cRqMshr_pipelineResp_getRq_IF_cache_pipe_ETC___d3166,
       cache_cRqMshr_pipelineResp_searchEndOfChain_ca_ETC___d2669,
       cache_cRqMshr_sendRqToC_searchNeedRqChild_1_CO_ETC___d2482,
       cache_cRqRetryIndexQ_enqReq_dummy2_2_read__28__ETC___d864,
       cache_pipeline_RDY_deqWrite__580_AND_IF_cache__ETC___d2671,
       cache_pipeline_RDY_deqWrite__580_AND_NOT_cache_ETC___d3471,
       cache_pipeline_first__581_BITS_516_TO_513_583__ETC___d2588,
       cache_pipeline_first__581_BITS_516_TO_513_583__ETC___d3103,
       cache_pipeline_first__581_BITS_516_TO_513_583__ETC___d3287,
       cache_pipeline_first__581_BITS_516_TO_513_583__ETC___d3295,
       cache_pipeline_first__581_BITS_519_TO_518_594__ETC___d2598,
       cache_pipeline_first__581_BITS_519_TO_518_594__ETC___d2618,
       cache_pipeline_first__581_BITS_519_TO_518_594__ETC___d3126,
       cache_pipeline_first__581_BITS_519_TO_518_594__ETC___d3136,
       cache_pipeline_first__581_BITS_519_TO_518_594__ETC___d3192,
       cache_pipeline_first__581_BITS_519_TO_518_594__ETC___d3196,
       cache_pipeline_first__581_BITS_519_TO_518_594__ETC___d3265,
       cache_pipeline_first__581_BITS_519_TO_518_594__ETC___d3271,
       cache_pipeline_first__581_BITS_521_TO_520_600__ETC___d2601,
       cache_pipeline_first__581_BITS_521_TO_520_600__ETC___d2621,
       cache_pipeline_first__581_BITS_523_TO_522_603__ETC___d2604,
       cache_pipeline_first__581_BITS_523_TO_522_603__ETC___d2624,
       cache_pipeline_first__581_BITS_573_TO_526_644__ETC___d2646,
       cache_pipeline_first__581_BIT_517_582_AND_NOT__ETC___d3820,
       cache_pipeline_first__581_BIT_517_582_AND_NOT__ETC___d3824,
       cache_pipeline_first__581_BIT_517_582_AND_cach_ETC___d3129,
       cache_pipeline_first__581_BIT_517_582_AND_cach_ETC___d3139,
       cache_pipeline_first__581_BIT_517_582_AND_cach_ETC___d3146,
       cache_pipeline_first__581_BIT_517_582_AND_cach_ETC___d3195,
       cache_pipeline_first__581_BIT_517_582_AND_cach_ETC___d3199,
       cache_pipeline_first__581_BIT_517_582_AND_cach_ETC___d3268,
       cache_pipeline_first__581_BIT_517_582_AND_cach_ETC___d3274,
       cache_pipeline_first__581_BIT_517_582_AND_cach_ETC___d3278,
       cache_pipeline_first__581_BIT_517_582_AND_cach_ETC___d3284,
       cache_rqFromCQ_enqReq_dummy2_2_read__4_AND_IF__ETC___d65,
       cache_rqFromDmaQ_enqReq_dummy2_2_read__40_AND__ETC___d371,
       cache_rsFromCQ_enqReq_dummy2_2_read__26_AND_IF_ETC___d157,
       cache_rsFromMQ_enqReq_dummy2_2_read__41_AND_IF_ETC___d772,
       cache_rsLdToDmaQ_enqReq_dummy2_2_read__31_AND__ETC___d462,
       cache_rsStToDmaQ_enqReq_dummy2_2_read__22_AND__ETC___d553,
       cache_rsToCIndexQ_enqReq_dummy2_2_read__51_AND_ETC___d987,
       cache_toCQ_enqReq_dummy2_2_read__53_AND_IF_cac_ETC___d279,
       cache_toMQ_enqReq_dummy2_2_read__54_AND_IF_cac_ETC___d680,
       next_deqP___1__h119479,
       next_deqP___1__h135572,
       next_deqP___1__h143074,
       next_deqP___1__h208858,
       next_deqP___1__h225353,
       next_deqP___1__h22634,
       next_deqP___1__h38327,
       next_deqP___1__h7552,
       perfReqQ_enqReq_dummy2_2_read__870_AND_IF_perf_ETC___d3887,
       v__h129259,
       v__h129542,
       v__h142239,
       v__h142522,
       v__h16641,
       v__h168573,
       v__h168856,
       v__h16924,
       v__h218716,
       v__h218999,
       v__h31944,
       v__h32227,
       v__h6037,
       v__h6320,
       v__h72082,
       v__h72365;
  // value method to_child_rsFromC_notFull
  assign to_child_rsFromC_notFull = !cache_rsFromCQ_full ;
  assign RDY_to_child_rsFromC_notFull = 1'd1 ;
  // action method to_child_rsFromC_enq
  assign RDY_to_child_rsFromC_enq = !cache_rsFromCQ_full ;
  assign CAN_FIRE_to_child_rsFromC_enq = !cache_rsFromCQ_full ;
  assign WILL_FIRE_to_child_rsFromC_enq = EN_to_child_rsFromC_enq ;
  // value method to_child_rqFromC_notFull
  assign to_child_rqFromC_notFull = !cache_rqFromCQ_full ;
  assign RDY_to_child_rqFromC_notFull = 1'd1 ;
  // action method to_child_rqFromC_enq
  assign RDY_to_child_rqFromC_enq = !cache_rqFromCQ_full ;
  assign CAN_FIRE_to_child_rqFromC_enq = !cache_rqFromCQ_full ;
  assign WILL_FIRE_to_child_rqFromC_enq = EN_to_child_rqFromC_enq ;
  // value method to_child_toC_notEmpty
  assign to_child_toC_notEmpty = !cache_toCQ_empty ;
  assign RDY_to_child_toC_notEmpty = 1'd1 ;
  // action method to_child_toC_deq
  assign RDY_to_child_toC_deq = !cache_toCQ_empty ;
  assign CAN_FIRE_to_child_toC_deq = !cache_toCQ_empty ;
  assign WILL_FIRE_to_child_toC_deq = EN_to_child_toC_deq ;
  // value method to_child_toC_first
  assign to_child_toC_first =
	     { CASE_cache_toCQ_deqP_0_cache_toCQ_data_0_BIT_5_ETC__q256,
	       IF_SEL_ARR_NOT_cache_toCQ_data_0_917_BIT_584_9_ETC___d4000 } ;
  assign RDY_to_child_toC_first = !cache_toCQ_empty ;
  // value method dma_memReq_notFull
  assign dma_memReq_notFull = !cache_rqFromDmaQ_full ;
  assign RDY_dma_memReq_notFull = 1'd1 ;
  // action method dma_memReq_enq
  assign RDY_dma_memReq_enq = !cache_rqFromDmaQ_full ;
  assign CAN_FIRE_dma_memReq_enq = !cache_rqFromDmaQ_full ;
  assign WILL_FIRE_dma_memReq_enq = EN_dma_memReq_enq ;
  // value method dma_respLd_notEmpty
  assign dma_respLd_notEmpty = !cache_rsLdToDmaQ_empty ;
  assign RDY_dma_respLd_notEmpty = 1'd1 ;
  // action method dma_respLd_deq
  assign RDY_dma_respLd_deq = !cache_rsLdToDmaQ_empty ;
  assign CAN_FIRE_dma_respLd_deq = !cache_rsLdToDmaQ_empty ;
  assign WILL_FIRE_dma_respLd_deq = EN_dma_respLd_deq ;
  // value method dma_respLd_first
  assign dma_respLd_first =
	     { SEL_ARR_cache_rsLdToDmaQ_data_0_004_BITS_527_T_ETC___d4036,
	       CASE_cache_rsLdToDmaQ_deqP_0_cache_rsLdToDmaQ__ETC__q259,
	       x__h456399 } ;
  assign RDY_dma_respLd_first = !cache_rsLdToDmaQ_empty ;
  // value method dma_respSt_notEmpty
  assign dma_respSt_notEmpty = !cache_rsStToDmaQ_empty ;
  assign RDY_dma_respSt_notEmpty = 1'd1 ;
  // action method dma_respSt_deq
  assign RDY_dma_respSt_deq = !cache_rsStToDmaQ_empty ;
  assign CAN_FIRE_dma_respSt_deq = !cache_rsStToDmaQ_empty ;
  assign WILL_FIRE_dma_respSt_deq = EN_dma_respSt_deq ;
  // value method dma_respSt_first
  always@(cache_rsStToDmaQ_deqP or
	  cache_rsStToDmaQ_data_0 or cache_rsStToDmaQ_data_1)
  begin
    case (cache_rsStToDmaQ_deqP)
      1'd0: dma_respSt_first = cache_rsStToDmaQ_data_0;
      1'd1: dma_respSt_first = cache_rsStToDmaQ_data_1;
    endcase
  end
  assign RDY_dma_respSt_first = !cache_rsStToDmaQ_empty ;
  // value method to_mem_toM_notEmpty
  assign to_mem_toM_notEmpty = !cache_toMQ_empty ;
  assign RDY_to_mem_toM_notEmpty = 1'd1 ;
  // action method to_mem_toM_deq
  assign RDY_to_mem_toM_deq = !cache_toMQ_empty ;
  assign CAN_FIRE_to_mem_toM_deq = !cache_toMQ_empty ;
  assign WILL_FIRE_to_mem_toM_deq = EN_to_mem_toM_deq ;
  // value method to_mem_toM_first
  assign to_mem_toM_first =
	     { CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_6_ETC__q261,
	       IF_SEL_ARR_NOT_cache_toMQ_data_0_050_BIT_640_0_ETC___d4404 } ;
  assign RDY_to_mem_toM_first = !cache_toMQ_empty ;
  // value method to_mem_rsFromM_notFull
  assign to_mem_rsFromM_notFull = !cache_rsFromMQ_full ;
  assign RDY_to_mem_rsFromM_notFull = 1'd1 ;
  // action method to_mem_rsFromM_enq
  assign RDY_to_mem_rsFromM_enq = !cache_rsFromMQ_full ;
  assign CAN_FIRE_to_mem_rsFromM_enq = !cache_rsFromMQ_full ;
  assign WILL_FIRE_to_mem_rsFromM_enq = EN_to_mem_rsFromM_enq ;
  // actionvalue method cRqStuck_get
  assign cRqStuck_get =
	     { cache_cRqMshr$stuck_get[32:16],
	       cache_cRqMshr$stuck_get[167:100],
	       cache_cRqMshr$stuck_get[98:97],
	       cache_cRqMshr$stuck_get[15:0] } ;
  assign RDY_cRqStuck_get = cache_cRqMshr$RDY_stuck_get ;
  assign CAN_FIRE_cRqStuck_get = cache_cRqMshr$RDY_stuck_get ;
  assign WILL_FIRE_cRqStuck_get = EN_cRqStuck_get ;
  // action method perf_setStatus
  assign RDY_perf_setStatus = 1'd1 ;
  assign CAN_FIRE_perf_setStatus = 1'd1 ;
  assign WILL_FIRE_perf_setStatus = EN_perf_setStatus ;
  // action method perf_req
  assign RDY_perf_req = !perfReqQ_full ;
  assign CAN_FIRE_perf_req = !perfReqQ_full ;
  assign WILL_FIRE_perf_req = EN_perf_req ;
  // actionvalue method perf_resp
  assign perf_resp = { perfReqQ_data_0, 64'd0 } ;
  assign RDY_perf_resp = !perfReqQ_empty ;
  assign CAN_FIRE_perf_resp = !perfReqQ_empty ;
  assign WILL_FIRE_perf_resp = EN_perf_resp ;
  // value method perf_respValid
  assign perf_respValid = !perfReqQ_empty ;
  assign RDY_perf_respValid = 1'd1 ;
  // submodule cache_cRqMshr
  mkLastLvCRqMshr cache_cRqMshr(.CLK(CLK),
				.RST_N(RST_N),
				.mRsDeq_setData_d(cache_cRqMshr$mRsDeq_setData_d),
				.mRsDeq_setData_n(cache_cRqMshr$mRsDeq_setData_n),
				.pipelineResp_getAddrSucc_n(cache_cRqMshr$pipelineResp_getAddrSucc_n),
				.pipelineResp_getData_n(cache_cRqMshr$pipelineResp_getData_n),
				.pipelineResp_getRepSucc_n(cache_cRqMshr$pipelineResp_getRepSucc_n),
				.pipelineResp_getRq_n(cache_cRqMshr$pipelineResp_getRq_n),
				.pipelineResp_getSlot_n(cache_cRqMshr$pipelineResp_getSlot_n),
				.pipelineResp_getState_n(cache_cRqMshr$pipelineResp_getState_n),
				.pipelineResp_searchEndOfChain_addr(cache_cRqMshr$pipelineResp_searchEndOfChain_addr),
				.pipelineResp_setAddrSucc_n(cache_cRqMshr$pipelineResp_setAddrSucc_n),
				.pipelineResp_setAddrSucc_succ(cache_cRqMshr$pipelineResp_setAddrSucc_succ),
				.pipelineResp_setData_d(cache_cRqMshr$pipelineResp_setData_d),
				.pipelineResp_setData_n(cache_cRqMshr$pipelineResp_setData_n),
				.pipelineResp_setRepSucc_n(cache_cRqMshr$pipelineResp_setRepSucc_n),
				.pipelineResp_setRepSucc_succ(cache_cRqMshr$pipelineResp_setRepSucc_succ),
				.pipelineResp_setStateSlot_n(cache_cRqMshr$pipelineResp_setStateSlot_n),
				.pipelineResp_setStateSlot_slot(cache_cRqMshr$pipelineResp_setStateSlot_slot),
				.pipelineResp_setStateSlot_state(cache_cRqMshr$pipelineResp_setStateSlot_state),
				.sendRqToC_getRq_n(cache_cRqMshr$sendRqToC_getRq_n),
				.sendRqToC_getSlot_n(cache_cRqMshr$sendRqToC_getSlot_n),
				.sendRqToC_getState_n(cache_cRqMshr$sendRqToC_getState_n),
				.sendRqToC_searchNeedRqChild_suggestIdx(cache_cRqMshr$sendRqToC_searchNeedRqChild_suggestIdx),
				.sendRqToC_setSlot_n(cache_cRqMshr$sendRqToC_setSlot_n),
				.sendRqToC_setSlot_s(cache_cRqMshr$sendRqToC_setSlot_s),
				.sendRsToDmaC_getData_n(cache_cRqMshr$sendRsToDmaC_getData_n),
				.sendRsToDmaC_getRq_n(cache_cRqMshr$sendRsToDmaC_getRq_n),
				.sendRsToDmaC_releaseEntry_n(cache_cRqMshr$sendRsToDmaC_releaseEntry_n),
				.sendToM_getData_n(cache_cRqMshr$sendToM_getData_n),
				.sendToM_getRq_n(cache_cRqMshr$sendToM_getRq_n),
				.sendToM_getSlot_n(cache_cRqMshr$sendToM_getSlot_n),
				.transfer_getEmptyEntryInit_d(cache_cRqMshr$transfer_getEmptyEntryInit_d),
				.transfer_getEmptyEntryInit_r(cache_cRqMshr$transfer_getEmptyEntryInit_r),
				.transfer_getRq_n(cache_cRqMshr$transfer_getRq_n),
				.transfer_getSlot_n(cache_cRqMshr$transfer_getSlot_n),
				.transfer_hasEmptyEntry_r(cache_cRqMshr$transfer_hasEmptyEntry_r),
				.EN_transfer_getEmptyEntryInit(cache_cRqMshr$EN_transfer_getEmptyEntryInit),
				.EN_mRsDeq_setData(cache_cRqMshr$EN_mRsDeq_setData),
				.EN_sendRsToDmaC_releaseEntry(cache_cRqMshr$EN_sendRsToDmaC_releaseEntry),
				.EN_sendRqToC_setSlot(cache_cRqMshr$EN_sendRqToC_setSlot),
				.EN_pipelineResp_setData(cache_cRqMshr$EN_pipelineResp_setData),
				.EN_pipelineResp_setStateSlot(cache_cRqMshr$EN_pipelineResp_setStateSlot),
				.EN_pipelineResp_setAddrSucc(cache_cRqMshr$EN_pipelineResp_setAddrSucc),
				.EN_pipelineResp_setRepSucc(cache_cRqMshr$EN_pipelineResp_setRepSucc),
				.EN_stuck_get(cache_cRqMshr$EN_stuck_get),
				.transfer_getRq(cache_cRqMshr$transfer_getRq),
				.RDY_transfer_getRq(),
				.transfer_getSlot(cache_cRqMshr$transfer_getSlot),
				.RDY_transfer_getSlot(),
				.transfer_getEmptyEntryInit(cache_cRqMshr$transfer_getEmptyEntryInit),
				.RDY_transfer_getEmptyEntryInit(cache_cRqMshr$RDY_transfer_getEmptyEntryInit),
				.transfer_hasEmptyEntry(),
				.RDY_transfer_hasEmptyEntry(),
				.RDY_mRsDeq_setData(),
				.sendToM_getRq(cache_cRqMshr$sendToM_getRq),
				.RDY_sendToM_getRq(),
				.sendToM_getSlot(cache_cRqMshr$sendToM_getSlot),
				.RDY_sendToM_getSlot(),
				.sendToM_getData(cache_cRqMshr$sendToM_getData),
				.RDY_sendToM_getData(),
				.sendRsToDmaC_getRq(cache_cRqMshr$sendRsToDmaC_getRq),
				.RDY_sendRsToDmaC_getRq(),
				.sendRsToDmaC_getData(cache_cRqMshr$sendRsToDmaC_getData),
				.RDY_sendRsToDmaC_getData(),
				.RDY_sendRsToDmaC_releaseEntry(cache_cRqMshr$RDY_sendRsToDmaC_releaseEntry),
				.sendRqToC_getRq(cache_cRqMshr$sendRqToC_getRq),
				.RDY_sendRqToC_getRq(),
				.sendRqToC_getState(cache_cRqMshr$sendRqToC_getState),
				.RDY_sendRqToC_getState(),
				.sendRqToC_getSlot(cache_cRqMshr$sendRqToC_getSlot),
				.RDY_sendRqToC_getSlot(),
				.RDY_sendRqToC_setSlot(),
				.sendRqToC_searchNeedRqChild(cache_cRqMshr$sendRqToC_searchNeedRqChild),
				.RDY_sendRqToC_searchNeedRqChild(),
				.pipelineResp_getRq(cache_cRqMshr$pipelineResp_getRq),
				.RDY_pipelineResp_getRq(),
				.pipelineResp_getState(cache_cRqMshr$pipelineResp_getState),
				.RDY_pipelineResp_getState(),
				.pipelineResp_getSlot(cache_cRqMshr$pipelineResp_getSlot),
				.RDY_pipelineResp_getSlot(),
				.pipelineResp_getData(cache_cRqMshr$pipelineResp_getData),
				.RDY_pipelineResp_getData(),
				.pipelineResp_getAddrSucc(cache_cRqMshr$pipelineResp_getAddrSucc),
				.RDY_pipelineResp_getAddrSucc(),
				.pipelineResp_getRepSucc(cache_cRqMshr$pipelineResp_getRepSucc),
				.RDY_pipelineResp_getRepSucc(),
				.RDY_pipelineResp_setData(),
				.RDY_pipelineResp_setStateSlot(),
				.RDY_pipelineResp_setAddrSucc(),
				.RDY_pipelineResp_setRepSucc(),
				.pipelineResp_searchEndOfChain(cache_cRqMshr$pipelineResp_searchEndOfChain),
				.RDY_pipelineResp_searchEndOfChain(),
				.stuck_get(cache_cRqMshr$stuck_get),
				.RDY_stuck_get(cache_cRqMshr$RDY_stuck_get));
  // submodule cache_cRqRetryIndexQ_clearReq_dummy2_0
  RevertReg #(.width(32'd1),
	      .init(1'd1)) cache_cRqRetryIndexQ_clearReq_dummy2_0(.CLK(CLK),
								  .D_IN(cache_cRqRetryIndexQ_clearReq_dummy2_0$D_IN),
								  .EN(cache_cRqRetryIndexQ_clearReq_dummy2_0$EN),
								  .Q_OUT());
  // submodule cache_cRqRetryIndexQ_clearReq_dummy2_1
  RevertReg #(.width(32'd1),
	      .init(1'd1)) cache_cRqRetryIndexQ_clearReq_dummy2_1(.CLK(CLK),
								  .D_IN(cache_cRqRetryIndexQ_clearReq_dummy2_1$D_IN),
								  .EN(cache_cRqRetryIndexQ_clearReq_dummy2_1$EN),
								  .Q_OUT(cache_cRqRetryIndexQ_clearReq_dummy2_1$Q_OUT));
  // submodule cache_cRqRetryIndexQ_deqReq_dummy2_0
  RevertReg #(.width(32'd1),
	      .init(1'd1)) cache_cRqRetryIndexQ_deqReq_dummy2_0(.CLK(CLK),
								.D_IN(cache_cRqRetryIndexQ_deqReq_dummy2_0$D_IN),
								.EN(cache_cRqRetryIndexQ_deqReq_dummy2_0$EN),
								.Q_OUT());
  // submodule cache_cRqRetryIndexQ_deqReq_dummy2_1
  RevertReg #(.width(32'd1),
	      .init(1'd1)) cache_cRqRetryIndexQ_deqReq_dummy2_1(.CLK(CLK),
								.D_IN(cache_cRqRetryIndexQ_deqReq_dummy2_1$D_IN),
								.EN(cache_cRqRetryIndexQ_deqReq_dummy2_1$EN),
								.Q_OUT());
  // submodule cache_cRqRetryIndexQ_deqReq_dummy2_2
  RevertReg #(.width(32'd1),
	      .init(1'd1)) cache_cRqRetryIndexQ_deqReq_dummy2_2(.CLK(CLK),
								.D_IN(cache_cRqRetryIndexQ_deqReq_dummy2_2$D_IN),
								.EN(cache_cRqRetryIndexQ_deqReq_dummy2_2$EN),
								.Q_OUT(cache_cRqRetryIndexQ_deqReq_dummy2_2$Q_OUT));
  // submodule cache_cRqRetryIndexQ_enqReq_dummy2_0
  RevertReg #(.width(32'd1),
	      .init(1'd1)) cache_cRqRetryIndexQ_enqReq_dummy2_0(.CLK(CLK),
								.D_IN(cache_cRqRetryIndexQ_enqReq_dummy2_0$D_IN),
								.EN(cache_cRqRetryIndexQ_enqReq_dummy2_0$EN),
								.Q_OUT());
  // submodule cache_cRqRetryIndexQ_enqReq_dummy2_1
  RevertReg #(.width(32'd1),
	      .init(1'd1)) cache_cRqRetryIndexQ_enqReq_dummy2_1(.CLK(CLK),
								.D_IN(cache_cRqRetryIndexQ_enqReq_dummy2_1$D_IN),
								.EN(cache_cRqRetryIndexQ_enqReq_dummy2_1$EN),
								.Q_OUT());
  // submodule cache_cRqRetryIndexQ_enqReq_dummy2_2
  RevertReg #(.width(32'd1),
	      .init(1'd1)) cache_cRqRetryIndexQ_enqReq_dummy2_2(.CLK(CLK),
								.D_IN(cache_cRqRetryIndexQ_enqReq_dummy2_2$D_IN),
								.EN(cache_cRqRetryIndexQ_enqReq_dummy2_2$EN),
								.Q_OUT(cache_cRqRetryIndexQ_enqReq_dummy2_2$Q_OUT));
  // submodule cache_pipeline
  mkLLPipeline cache_pipeline(.CLK(CLK),
			      .RST_N(RST_N),
			      .deqWrite_swapRq(cache_pipeline$deqWrite_swapRq),
			      .deqWrite_updateRep(cache_pipeline$deqWrite_updateRep),
			      .deqWrite_wrRam(cache_pipeline$deqWrite_wrRam),
			      .send_r(cache_pipeline$send_r),
			      .EN_send(cache_pipeline$EN_send),
			      .EN_deqWrite(cache_pipeline$EN_deqWrite),
			      .RDY_send(cache_pipeline$RDY_send),
			      .notEmpty(cache_pipeline$notEmpty),
			      .RDY_notEmpty(),
			      .first(cache_pipeline$first),
			      .RDY_first(cache_pipeline$RDY_first),
			      .unguard_first(cache_pipeline$unguard_first),
			      .RDY_unguard_first(cache_pipeline$RDY_unguard_first),
			      .RDY_deqWrite(cache_pipeline$RDY_deqWrite));
  // submodule cache_rqFromCQ_clearReq_dummy2_0
  RevertReg #(.width(32'd1),
	      .init(1'd1)) cache_rqFromCQ_clearReq_dummy2_0(.CLK(CLK),
							    .D_IN(cache_rqFromCQ_clearReq_dummy2_0$D_IN),
							    .EN(cache_rqFromCQ_clearReq_dummy2_0$EN),
							    .Q_OUT());
  // submodule cache_rqFromCQ_clearReq_dummy2_1
  RevertReg #(.width(32'd1),
	      .init(1'd1)) cache_rqFromCQ_clearReq_dummy2_1(.CLK(CLK),
							    .D_IN(cache_rqFromCQ_clearReq_dummy2_1$D_IN),
							    .EN(cache_rqFromCQ_clearReq_dummy2_1$EN),
							    .Q_OUT(cache_rqFromCQ_clearReq_dummy2_1$Q_OUT));
  // submodule cache_rqFromCQ_deqReq_dummy2_0
  RevertReg #(.width(32'd1),
	      .init(1'd1)) cache_rqFromCQ_deqReq_dummy2_0(.CLK(CLK),
							  .D_IN(cache_rqFromCQ_deqReq_dummy2_0$D_IN),
							  .EN(cache_rqFromCQ_deqReq_dummy2_0$EN),
							  .Q_OUT());
  // submodule cache_rqFromCQ_deqReq_dummy2_1
  RevertReg #(.width(32'd1),
	      .init(1'd1)) cache_rqFromCQ_deqReq_dummy2_1(.CLK(CLK),
							  .D_IN(cache_rqFromCQ_deqReq_dummy2_1$D_IN),
							  .EN(cache_rqFromCQ_deqReq_dummy2_1$EN),
							  .Q_OUT());
  // submodule cache_rqFromCQ_deqReq_dummy2_2
  RevertReg #(.width(32'd1),
	      .init(1'd1)) cache_rqFromCQ_deqReq_dummy2_2(.CLK(CLK),
							  .D_IN(cache_rqFromCQ_deqReq_dummy2_2$D_IN),
							  .EN(cache_rqFromCQ_deqReq_dummy2_2$EN),
							  .Q_OUT(cache_rqFromCQ_deqReq_dummy2_2$Q_OUT));
  // submodule cache_rqFromCQ_enqReq_dummy2_0
  RevertReg #(.width(32'd1),
	      .init(1'd1)) cache_rqFromCQ_enqReq_dummy2_0(.CLK(CLK),
							  .D_IN(cache_rqFromCQ_enqReq_dummy2_0$D_IN),
							  .EN(cache_rqFromCQ_enqReq_dummy2_0$EN),
							  .Q_OUT());
  // submodule cache_rqFromCQ_enqReq_dummy2_1
  RevertReg #(.width(32'd1),
	      .init(1'd1)) cache_rqFromCQ_enqReq_dummy2_1(.CLK(CLK),
							  .D_IN(cache_rqFromCQ_enqReq_dummy2_1$D_IN),
							  .EN(cache_rqFromCQ_enqReq_dummy2_1$EN),
							  .Q_OUT());
  // submodule cache_rqFromCQ_enqReq_dummy2_2
  RevertReg #(.width(32'd1),
	      .init(1'd1)) cache_rqFromCQ_enqReq_dummy2_2(.CLK(CLK),
							  .D_IN(cache_rqFromCQ_enqReq_dummy2_2$D_IN),
							  .EN(cache_rqFromCQ_enqReq_dummy2_2$EN),
							  .Q_OUT(cache_rqFromCQ_enqReq_dummy2_2$Q_OUT));
  // submodule cache_rqFromDmaQ_clearReq_dummy2_0
  RevertReg #(.width(32'd1),
	      .init(1'd1)) cache_rqFromDmaQ_clearReq_dummy2_0(.CLK(CLK),
							      .D_IN(cache_rqFromDmaQ_clearReq_dummy2_0$D_IN),
							      .EN(cache_rqFromDmaQ_clearReq_dummy2_0$EN),
							      .Q_OUT());
  // submodule cache_rqFromDmaQ_clearReq_dummy2_1
  RevertReg #(.width(32'd1),
	      .init(1'd1)) cache_rqFromDmaQ_clearReq_dummy2_1(.CLK(CLK),
							      .D_IN(cache_rqFromDmaQ_clearReq_dummy2_1$D_IN),
							      .EN(cache_rqFromDmaQ_clearReq_dummy2_1$EN),
							      .Q_OUT(cache_rqFromDmaQ_clearReq_dummy2_1$Q_OUT));
  // submodule cache_rqFromDmaQ_deqReq_dummy2_0
  RevertReg #(.width(32'd1),
	      .init(1'd1)) cache_rqFromDmaQ_deqReq_dummy2_0(.CLK(CLK),
							    .D_IN(cache_rqFromDmaQ_deqReq_dummy2_0$D_IN),
							    .EN(cache_rqFromDmaQ_deqReq_dummy2_0$EN),
							    .Q_OUT());
  // submodule cache_rqFromDmaQ_deqReq_dummy2_1
  RevertReg #(.width(32'd1),
	      .init(1'd1)) cache_rqFromDmaQ_deqReq_dummy2_1(.CLK(CLK),
							    .D_IN(cache_rqFromDmaQ_deqReq_dummy2_1$D_IN),
							    .EN(cache_rqFromDmaQ_deqReq_dummy2_1$EN),
							    .Q_OUT());
  // submodule cache_rqFromDmaQ_deqReq_dummy2_2
  RevertReg #(.width(32'd1),
	      .init(1'd1)) cache_rqFromDmaQ_deqReq_dummy2_2(.CLK(CLK),
							    .D_IN(cache_rqFromDmaQ_deqReq_dummy2_2$D_IN),
							    .EN(cache_rqFromDmaQ_deqReq_dummy2_2$EN),
							    .Q_OUT(cache_rqFromDmaQ_deqReq_dummy2_2$Q_OUT));
  // submodule cache_rqFromDmaQ_enqReq_dummy2_0
  RevertReg #(.width(32'd1),
	      .init(1'd1)) cache_rqFromDmaQ_enqReq_dummy2_0(.CLK(CLK),
							    .D_IN(cache_rqFromDmaQ_enqReq_dummy2_0$D_IN),
							    .EN(cache_rqFromDmaQ_enqReq_dummy2_0$EN),
							    .Q_OUT());
  // submodule cache_rqFromDmaQ_enqReq_dummy2_1
  RevertReg #(.width(32'd1),
	      .init(1'd1)) cache_rqFromDmaQ_enqReq_dummy2_1(.CLK(CLK),
							    .D_IN(cache_rqFromDmaQ_enqReq_dummy2_1$D_IN),
							    .EN(cache_rqFromDmaQ_enqReq_dummy2_1$EN),
							    .Q_OUT());
  // submodule cache_rqFromDmaQ_enqReq_dummy2_2
  RevertReg #(.width(32'd1),
	      .init(1'd1)) cache_rqFromDmaQ_enqReq_dummy2_2(.CLK(CLK),
							    .D_IN(cache_rqFromDmaQ_enqReq_dummy2_2$D_IN),
							    .EN(cache_rqFromDmaQ_enqReq_dummy2_2$EN),
							    .Q_OUT(cache_rqFromDmaQ_enqReq_dummy2_2$Q_OUT));
  // submodule cache_rsFromCQ_clearReq_dummy2_0
  RevertReg #(.width(32'd1),
	      .init(1'd1)) cache_rsFromCQ_clearReq_dummy2_0(.CLK(CLK),
							    .D_IN(cache_rsFromCQ_clearReq_dummy2_0$D_IN),
							    .EN(cache_rsFromCQ_clearReq_dummy2_0$EN),
							    .Q_OUT());
  // submodule cache_rsFromCQ_clearReq_dummy2_1
  RevertReg #(.width(32'd1),
	      .init(1'd1)) cache_rsFromCQ_clearReq_dummy2_1(.CLK(CLK),
							    .D_IN(cache_rsFromCQ_clearReq_dummy2_1$D_IN),
							    .EN(cache_rsFromCQ_clearReq_dummy2_1$EN),
							    .Q_OUT(cache_rsFromCQ_clearReq_dummy2_1$Q_OUT));
  // submodule cache_rsFromCQ_deqReq_dummy2_0
  RevertReg #(.width(32'd1),
	      .init(1'd1)) cache_rsFromCQ_deqReq_dummy2_0(.CLK(CLK),
							  .D_IN(cache_rsFromCQ_deqReq_dummy2_0$D_IN),
							  .EN(cache_rsFromCQ_deqReq_dummy2_0$EN),
							  .Q_OUT());
  // submodule cache_rsFromCQ_deqReq_dummy2_1
  RevertReg #(.width(32'd1),
	      .init(1'd1)) cache_rsFromCQ_deqReq_dummy2_1(.CLK(CLK),
							  .D_IN(cache_rsFromCQ_deqReq_dummy2_1$D_IN),
							  .EN(cache_rsFromCQ_deqReq_dummy2_1$EN),
							  .Q_OUT());
  // submodule cache_rsFromCQ_deqReq_dummy2_2
  RevertReg #(.width(32'd1),
	      .init(1'd1)) cache_rsFromCQ_deqReq_dummy2_2(.CLK(CLK),
							  .D_IN(cache_rsFromCQ_deqReq_dummy2_2$D_IN),
							  .EN(cache_rsFromCQ_deqReq_dummy2_2$EN),
							  .Q_OUT(cache_rsFromCQ_deqReq_dummy2_2$Q_OUT));
  // submodule cache_rsFromCQ_enqReq_dummy2_0
  RevertReg #(.width(32'd1),
	      .init(1'd1)) cache_rsFromCQ_enqReq_dummy2_0(.CLK(CLK),
							  .D_IN(cache_rsFromCQ_enqReq_dummy2_0$D_IN),
							  .EN(cache_rsFromCQ_enqReq_dummy2_0$EN),
							  .Q_OUT());
  // submodule cache_rsFromCQ_enqReq_dummy2_1
  RevertReg #(.width(32'd1),
	      .init(1'd1)) cache_rsFromCQ_enqReq_dummy2_1(.CLK(CLK),
							  .D_IN(cache_rsFromCQ_enqReq_dummy2_1$D_IN),
							  .EN(cache_rsFromCQ_enqReq_dummy2_1$EN),
							  .Q_OUT());
  // submodule cache_rsFromCQ_enqReq_dummy2_2
  RevertReg #(.width(32'd1),
	      .init(1'd1)) cache_rsFromCQ_enqReq_dummy2_2(.CLK(CLK),
							  .D_IN(cache_rsFromCQ_enqReq_dummy2_2$D_IN),
							  .EN(cache_rsFromCQ_enqReq_dummy2_2$EN),
							  .Q_OUT(cache_rsFromCQ_enqReq_dummy2_2$Q_OUT));
  // submodule cache_rsFromMQ_clearReq_dummy2_0
  RevertReg #(.width(32'd1),
	      .init(1'd1)) cache_rsFromMQ_clearReq_dummy2_0(.CLK(CLK),
							    .D_IN(cache_rsFromMQ_clearReq_dummy2_0$D_IN),
							    .EN(cache_rsFromMQ_clearReq_dummy2_0$EN),
							    .Q_OUT());
  // submodule cache_rsFromMQ_clearReq_dummy2_1
  RevertReg #(.width(32'd1),
	      .init(1'd1)) cache_rsFromMQ_clearReq_dummy2_1(.CLK(CLK),
							    .D_IN(cache_rsFromMQ_clearReq_dummy2_1$D_IN),
							    .EN(cache_rsFromMQ_clearReq_dummy2_1$EN),
							    .Q_OUT(cache_rsFromMQ_clearReq_dummy2_1$Q_OUT));
  // submodule cache_rsFromMQ_deqReq_dummy2_0
  RevertReg #(.width(32'd1),
	      .init(1'd1)) cache_rsFromMQ_deqReq_dummy2_0(.CLK(CLK),
							  .D_IN(cache_rsFromMQ_deqReq_dummy2_0$D_IN),
							  .EN(cache_rsFromMQ_deqReq_dummy2_0$EN),
							  .Q_OUT());
  // submodule cache_rsFromMQ_deqReq_dummy2_1
  RevertReg #(.width(32'd1),
	      .init(1'd1)) cache_rsFromMQ_deqReq_dummy2_1(.CLK(CLK),
							  .D_IN(cache_rsFromMQ_deqReq_dummy2_1$D_IN),
							  .EN(cache_rsFromMQ_deqReq_dummy2_1$EN),
							  .Q_OUT());
  // submodule cache_rsFromMQ_deqReq_dummy2_2
  RevertReg #(.width(32'd1),
	      .init(1'd1)) cache_rsFromMQ_deqReq_dummy2_2(.CLK(CLK),
							  .D_IN(cache_rsFromMQ_deqReq_dummy2_2$D_IN),
							  .EN(cache_rsFromMQ_deqReq_dummy2_2$EN),
							  .Q_OUT(cache_rsFromMQ_deqReq_dummy2_2$Q_OUT));
  // submodule cache_rsFromMQ_enqReq_dummy2_0
  RevertReg #(.width(32'd1),
	      .init(1'd1)) cache_rsFromMQ_enqReq_dummy2_0(.CLK(CLK),
							  .D_IN(cache_rsFromMQ_enqReq_dummy2_0$D_IN),
							  .EN(cache_rsFromMQ_enqReq_dummy2_0$EN),
							  .Q_OUT());
  // submodule cache_rsFromMQ_enqReq_dummy2_1
  RevertReg #(.width(32'd1),
	      .init(1'd1)) cache_rsFromMQ_enqReq_dummy2_1(.CLK(CLK),
							  .D_IN(cache_rsFromMQ_enqReq_dummy2_1$D_IN),
							  .EN(cache_rsFromMQ_enqReq_dummy2_1$EN),
							  .Q_OUT());
  // submodule cache_rsFromMQ_enqReq_dummy2_2
  RevertReg #(.width(32'd1),
	      .init(1'd1)) cache_rsFromMQ_enqReq_dummy2_2(.CLK(CLK),
							  .D_IN(cache_rsFromMQ_enqReq_dummy2_2$D_IN),
							  .EN(cache_rsFromMQ_enqReq_dummy2_2$EN),
							  .Q_OUT(cache_rsFromMQ_enqReq_dummy2_2$Q_OUT));
  // submodule cache_rsLdToDmaIndexQ
  SizedFIFO #(.p1width(32'd4),
	      .p2depth(32'd16),
	      .p3cntr_width(32'd4),
	      .guarded(1'd1)) cache_rsLdToDmaIndexQ(.RST(RST_N),
						    .CLK(CLK),
						    .D_IN(cache_rsLdToDmaIndexQ$D_IN),
						    .ENQ(cache_rsLdToDmaIndexQ$ENQ),
						    .DEQ(cache_rsLdToDmaIndexQ$DEQ),
						    .CLR(cache_rsLdToDmaIndexQ$CLR),
						    .D_OUT(cache_rsLdToDmaIndexQ$D_OUT),
						    .FULL_N(cache_rsLdToDmaIndexQ$FULL_N),
						    .EMPTY_N(cache_rsLdToDmaIndexQ$EMPTY_N));
  // submodule cache_rsLdToDmaIndexQ_mRsDeq
  FIFO2 #(.width(32'd4),
	  .guarded(1'd1)) cache_rsLdToDmaIndexQ_mRsDeq(.RST(RST_N),
						       .CLK(CLK),
						       .D_IN(cache_rsLdToDmaIndexQ_mRsDeq$D_IN),
						       .ENQ(cache_rsLdToDmaIndexQ_mRsDeq$ENQ),
						       .DEQ(cache_rsLdToDmaIndexQ_mRsDeq$DEQ),
						       .CLR(cache_rsLdToDmaIndexQ_mRsDeq$CLR),
						       .D_OUT(cache_rsLdToDmaIndexQ_mRsDeq$D_OUT),
						       .FULL_N(cache_rsLdToDmaIndexQ_mRsDeq$FULL_N),
						       .EMPTY_N(cache_rsLdToDmaIndexQ_mRsDeq$EMPTY_N));
  // submodule cache_rsLdToDmaIndexQ_pipelineResp
  FIFO2 #(.width(32'd4),
	  .guarded(1'd1)) cache_rsLdToDmaIndexQ_pipelineResp(.RST(RST_N),
							     .CLK(CLK),
							     .D_IN(cache_rsLdToDmaIndexQ_pipelineResp$D_IN),
							     .ENQ(cache_rsLdToDmaIndexQ_pipelineResp$ENQ),
							     .DEQ(cache_rsLdToDmaIndexQ_pipelineResp$DEQ),
							     .CLR(cache_rsLdToDmaIndexQ_pipelineResp$CLR),
							     .D_OUT(cache_rsLdToDmaIndexQ_pipelineResp$D_OUT),
							     .FULL_N(cache_rsLdToDmaIndexQ_pipelineResp$FULL_N),
							     .EMPTY_N(cache_rsLdToDmaIndexQ_pipelineResp$EMPTY_N));
  // submodule cache_rsLdToDmaQ_clearReq_dummy2_0
  RevertReg #(.width(32'd1),
	      .init(1'd1)) cache_rsLdToDmaQ_clearReq_dummy2_0(.CLK(CLK),
							      .D_IN(cache_rsLdToDmaQ_clearReq_dummy2_0$D_IN),
							      .EN(cache_rsLdToDmaQ_clearReq_dummy2_0$EN),
							      .Q_OUT());
  // submodule cache_rsLdToDmaQ_clearReq_dummy2_1
  RevertReg #(.width(32'd1),
	      .init(1'd1)) cache_rsLdToDmaQ_clearReq_dummy2_1(.CLK(CLK),
							      .D_IN(cache_rsLdToDmaQ_clearReq_dummy2_1$D_IN),
							      .EN(cache_rsLdToDmaQ_clearReq_dummy2_1$EN),
							      .Q_OUT(cache_rsLdToDmaQ_clearReq_dummy2_1$Q_OUT));
  // submodule cache_rsLdToDmaQ_deqReq_dummy2_0
  RevertReg #(.width(32'd1),
	      .init(1'd1)) cache_rsLdToDmaQ_deqReq_dummy2_0(.CLK(CLK),
							    .D_IN(cache_rsLdToDmaQ_deqReq_dummy2_0$D_IN),
							    .EN(cache_rsLdToDmaQ_deqReq_dummy2_0$EN),
							    .Q_OUT());
  // submodule cache_rsLdToDmaQ_deqReq_dummy2_1
  RevertReg #(.width(32'd1),
	      .init(1'd1)) cache_rsLdToDmaQ_deqReq_dummy2_1(.CLK(CLK),
							    .D_IN(cache_rsLdToDmaQ_deqReq_dummy2_1$D_IN),
							    .EN(cache_rsLdToDmaQ_deqReq_dummy2_1$EN),
							    .Q_OUT());
  // submodule cache_rsLdToDmaQ_deqReq_dummy2_2
  RevertReg #(.width(32'd1),
	      .init(1'd1)) cache_rsLdToDmaQ_deqReq_dummy2_2(.CLK(CLK),
							    .D_IN(cache_rsLdToDmaQ_deqReq_dummy2_2$D_IN),
							    .EN(cache_rsLdToDmaQ_deqReq_dummy2_2$EN),
							    .Q_OUT(cache_rsLdToDmaQ_deqReq_dummy2_2$Q_OUT));
  // submodule cache_rsLdToDmaQ_enqReq_dummy2_0
  RevertReg #(.width(32'd1),
	      .init(1'd1)) cache_rsLdToDmaQ_enqReq_dummy2_0(.CLK(CLK),
							    .D_IN(cache_rsLdToDmaQ_enqReq_dummy2_0$D_IN),
							    .EN(cache_rsLdToDmaQ_enqReq_dummy2_0$EN),
							    .Q_OUT());
  // submodule cache_rsLdToDmaQ_enqReq_dummy2_1
  RevertReg #(.width(32'd1),
	      .init(1'd1)) cache_rsLdToDmaQ_enqReq_dummy2_1(.CLK(CLK),
							    .D_IN(cache_rsLdToDmaQ_enqReq_dummy2_1$D_IN),
							    .EN(cache_rsLdToDmaQ_enqReq_dummy2_1$EN),
							    .Q_OUT());
  // submodule cache_rsLdToDmaQ_enqReq_dummy2_2
  RevertReg #(.width(32'd1),
	      .init(1'd1)) cache_rsLdToDmaQ_enqReq_dummy2_2(.CLK(CLK),
							    .D_IN(cache_rsLdToDmaQ_enqReq_dummy2_2$D_IN),
							    .EN(cache_rsLdToDmaQ_enqReq_dummy2_2$EN),
							    .Q_OUT(cache_rsLdToDmaQ_enqReq_dummy2_2$Q_OUT));
  // submodule cache_rsStToDmaIndexQ
  SizedFIFO #(.p1width(32'd4),
	      .p2depth(32'd16),
	      .p3cntr_width(32'd4),
	      .guarded(1'd1)) cache_rsStToDmaIndexQ(.RST(RST_N),
						    .CLK(CLK),
						    .D_IN(cache_rsStToDmaIndexQ$D_IN),
						    .ENQ(cache_rsStToDmaIndexQ$ENQ),
						    .DEQ(cache_rsStToDmaIndexQ$DEQ),
						    .CLR(cache_rsStToDmaIndexQ$CLR),
						    .D_OUT(cache_rsStToDmaIndexQ$D_OUT),
						    .FULL_N(cache_rsStToDmaIndexQ$FULL_N),
						    .EMPTY_N(cache_rsStToDmaIndexQ$EMPTY_N));
  // submodule cache_rsStToDmaIndexQ_pipelineResp
  FIFO2 #(.width(32'd4),
	  .guarded(1'd1)) cache_rsStToDmaIndexQ_pipelineResp(.RST(RST_N),
							     .CLK(CLK),
							     .D_IN(cache_rsStToDmaIndexQ_pipelineResp$D_IN),
							     .ENQ(cache_rsStToDmaIndexQ_pipelineResp$ENQ),
							     .DEQ(cache_rsStToDmaIndexQ_pipelineResp$DEQ),
							     .CLR(cache_rsStToDmaIndexQ_pipelineResp$CLR),
							     .D_OUT(cache_rsStToDmaIndexQ_pipelineResp$D_OUT),
							     .FULL_N(cache_rsStToDmaIndexQ_pipelineResp$FULL_N),
							     .EMPTY_N(cache_rsStToDmaIndexQ_pipelineResp$EMPTY_N));
  // submodule cache_rsStToDmaIndexQ_sendToM
  FIFO2 #(.width(32'd4),
	  .guarded(1'd1)) cache_rsStToDmaIndexQ_sendToM(.RST(RST_N),
							.CLK(CLK),
							.D_IN(cache_rsStToDmaIndexQ_sendToM$D_IN),
							.ENQ(cache_rsStToDmaIndexQ_sendToM$ENQ),
							.DEQ(cache_rsStToDmaIndexQ_sendToM$DEQ),
							.CLR(cache_rsStToDmaIndexQ_sendToM$CLR),
							.D_OUT(cache_rsStToDmaIndexQ_sendToM$D_OUT),
							.FULL_N(cache_rsStToDmaIndexQ_sendToM$FULL_N),
							.EMPTY_N(cache_rsStToDmaIndexQ_sendToM$EMPTY_N));
  // submodule cache_rsStToDmaQ_clearReq_dummy2_0
  RevertReg #(.width(32'd1),
	      .init(1'd1)) cache_rsStToDmaQ_clearReq_dummy2_0(.CLK(CLK),
							      .D_IN(cache_rsStToDmaQ_clearReq_dummy2_0$D_IN),
							      .EN(cache_rsStToDmaQ_clearReq_dummy2_0$EN),
							      .Q_OUT());
  // submodule cache_rsStToDmaQ_clearReq_dummy2_1
  RevertReg #(.width(32'd1),
	      .init(1'd1)) cache_rsStToDmaQ_clearReq_dummy2_1(.CLK(CLK),
							      .D_IN(cache_rsStToDmaQ_clearReq_dummy2_1$D_IN),
							      .EN(cache_rsStToDmaQ_clearReq_dummy2_1$EN),
							      .Q_OUT(cache_rsStToDmaQ_clearReq_dummy2_1$Q_OUT));
  // submodule cache_rsStToDmaQ_deqReq_dummy2_0
  RevertReg #(.width(32'd1),
	      .init(1'd1)) cache_rsStToDmaQ_deqReq_dummy2_0(.CLK(CLK),
							    .D_IN(cache_rsStToDmaQ_deqReq_dummy2_0$D_IN),
							    .EN(cache_rsStToDmaQ_deqReq_dummy2_0$EN),
							    .Q_OUT());
  // submodule cache_rsStToDmaQ_deqReq_dummy2_1
  RevertReg #(.width(32'd1),
	      .init(1'd1)) cache_rsStToDmaQ_deqReq_dummy2_1(.CLK(CLK),
							    .D_IN(cache_rsStToDmaQ_deqReq_dummy2_1$D_IN),
							    .EN(cache_rsStToDmaQ_deqReq_dummy2_1$EN),
							    .Q_OUT());
  // submodule cache_rsStToDmaQ_deqReq_dummy2_2
  RevertReg #(.width(32'd1),
	      .init(1'd1)) cache_rsStToDmaQ_deqReq_dummy2_2(.CLK(CLK),
							    .D_IN(cache_rsStToDmaQ_deqReq_dummy2_2$D_IN),
							    .EN(cache_rsStToDmaQ_deqReq_dummy2_2$EN),
							    .Q_OUT(cache_rsStToDmaQ_deqReq_dummy2_2$Q_OUT));
  // submodule cache_rsStToDmaQ_enqReq_dummy2_0
  RevertReg #(.width(32'd1),
	      .init(1'd1)) cache_rsStToDmaQ_enqReq_dummy2_0(.CLK(CLK),
							    .D_IN(cache_rsStToDmaQ_enqReq_dummy2_0$D_IN),
							    .EN(cache_rsStToDmaQ_enqReq_dummy2_0$EN),
							    .Q_OUT());
  // submodule cache_rsStToDmaQ_enqReq_dummy2_1
  RevertReg #(.width(32'd1),
	      .init(1'd1)) cache_rsStToDmaQ_enqReq_dummy2_1(.CLK(CLK),
							    .D_IN(cache_rsStToDmaQ_enqReq_dummy2_1$D_IN),
							    .EN(cache_rsStToDmaQ_enqReq_dummy2_1$EN),
							    .Q_OUT());
  // submodule cache_rsStToDmaQ_enqReq_dummy2_2
  RevertReg #(.width(32'd1),
	      .init(1'd1)) cache_rsStToDmaQ_enqReq_dummy2_2(.CLK(CLK),
							    .D_IN(cache_rsStToDmaQ_enqReq_dummy2_2$D_IN),
							    .EN(cache_rsStToDmaQ_enqReq_dummy2_2$EN),
							    .Q_OUT(cache_rsStToDmaQ_enqReq_dummy2_2$Q_OUT));
  // submodule cache_rsToCIndexQ_clearReq_dummy2_0
  RevertReg #(.width(32'd1),
	      .init(1'd1)) cache_rsToCIndexQ_clearReq_dummy2_0(.CLK(CLK),
							       .D_IN(cache_rsToCIndexQ_clearReq_dummy2_0$D_IN),
							       .EN(cache_rsToCIndexQ_clearReq_dummy2_0$EN),
							       .Q_OUT());
  // submodule cache_rsToCIndexQ_clearReq_dummy2_1
  RevertReg #(.width(32'd1),
	      .init(1'd1)) cache_rsToCIndexQ_clearReq_dummy2_1(.CLK(CLK),
							       .D_IN(cache_rsToCIndexQ_clearReq_dummy2_1$D_IN),
							       .EN(cache_rsToCIndexQ_clearReq_dummy2_1$EN),
							       .Q_OUT(cache_rsToCIndexQ_clearReq_dummy2_1$Q_OUT));
  // submodule cache_rsToCIndexQ_deqReq_dummy2_0
  RevertReg #(.width(32'd1),
	      .init(1'd1)) cache_rsToCIndexQ_deqReq_dummy2_0(.CLK(CLK),
							     .D_IN(cache_rsToCIndexQ_deqReq_dummy2_0$D_IN),
							     .EN(cache_rsToCIndexQ_deqReq_dummy2_0$EN),
							     .Q_OUT());
  // submodule cache_rsToCIndexQ_deqReq_dummy2_1
  RevertReg #(.width(32'd1),
	      .init(1'd1)) cache_rsToCIndexQ_deqReq_dummy2_1(.CLK(CLK),
							     .D_IN(cache_rsToCIndexQ_deqReq_dummy2_1$D_IN),
							     .EN(cache_rsToCIndexQ_deqReq_dummy2_1$EN),
							     .Q_OUT());
  // submodule cache_rsToCIndexQ_deqReq_dummy2_2
  RevertReg #(.width(32'd1),
	      .init(1'd1)) cache_rsToCIndexQ_deqReq_dummy2_2(.CLK(CLK),
							     .D_IN(cache_rsToCIndexQ_deqReq_dummy2_2$D_IN),
							     .EN(cache_rsToCIndexQ_deqReq_dummy2_2$EN),
							     .Q_OUT(cache_rsToCIndexQ_deqReq_dummy2_2$Q_OUT));
  // submodule cache_rsToCIndexQ_enqReq_dummy2_0
  RevertReg #(.width(32'd1),
	      .init(1'd1)) cache_rsToCIndexQ_enqReq_dummy2_0(.CLK(CLK),
							     .D_IN(cache_rsToCIndexQ_enqReq_dummy2_0$D_IN),
							     .EN(cache_rsToCIndexQ_enqReq_dummy2_0$EN),
							     .Q_OUT());
  // submodule cache_rsToCIndexQ_enqReq_dummy2_1
  RevertReg #(.width(32'd1),
	      .init(1'd1)) cache_rsToCIndexQ_enqReq_dummy2_1(.CLK(CLK),
							     .D_IN(cache_rsToCIndexQ_enqReq_dummy2_1$D_IN),
							     .EN(cache_rsToCIndexQ_enqReq_dummy2_1$EN),
							     .Q_OUT());
  // submodule cache_rsToCIndexQ_enqReq_dummy2_2
  RevertReg #(.width(32'd1),
	      .init(1'd1)) cache_rsToCIndexQ_enqReq_dummy2_2(.CLK(CLK),
							     .D_IN(cache_rsToCIndexQ_enqReq_dummy2_2$D_IN),
							     .EN(cache_rsToCIndexQ_enqReq_dummy2_2$EN),
							     .Q_OUT(cache_rsToCIndexQ_enqReq_dummy2_2$Q_OUT));
  // submodule cache_toCQ_clearReq_dummy2_0
  RevertReg #(.width(32'd1),
	      .init(1'd1)) cache_toCQ_clearReq_dummy2_0(.CLK(CLK),
							.D_IN(cache_toCQ_clearReq_dummy2_0$D_IN),
							.EN(cache_toCQ_clearReq_dummy2_0$EN),
							.Q_OUT());
  // submodule cache_toCQ_clearReq_dummy2_1
  RevertReg #(.width(32'd1),
	      .init(1'd1)) cache_toCQ_clearReq_dummy2_1(.CLK(CLK),
							.D_IN(cache_toCQ_clearReq_dummy2_1$D_IN),
							.EN(cache_toCQ_clearReq_dummy2_1$EN),
							.Q_OUT(cache_toCQ_clearReq_dummy2_1$Q_OUT));
  // submodule cache_toCQ_deqReq_dummy2_0
  RevertReg #(.width(32'd1),
	      .init(1'd1)) cache_toCQ_deqReq_dummy2_0(.CLK(CLK),
						      .D_IN(cache_toCQ_deqReq_dummy2_0$D_IN),
						      .EN(cache_toCQ_deqReq_dummy2_0$EN),
						      .Q_OUT());
  // submodule cache_toCQ_deqReq_dummy2_1
  RevertReg #(.width(32'd1),
	      .init(1'd1)) cache_toCQ_deqReq_dummy2_1(.CLK(CLK),
						      .D_IN(cache_toCQ_deqReq_dummy2_1$D_IN),
						      .EN(cache_toCQ_deqReq_dummy2_1$EN),
						      .Q_OUT());
  // submodule cache_toCQ_deqReq_dummy2_2
  RevertReg #(.width(32'd1),
	      .init(1'd1)) cache_toCQ_deqReq_dummy2_2(.CLK(CLK),
						      .D_IN(cache_toCQ_deqReq_dummy2_2$D_IN),
						      .EN(cache_toCQ_deqReq_dummy2_2$EN),
						      .Q_OUT(cache_toCQ_deqReq_dummy2_2$Q_OUT));
  // submodule cache_toCQ_enqReq_dummy2_0
  RevertReg #(.width(32'd1),
	      .init(1'd1)) cache_toCQ_enqReq_dummy2_0(.CLK(CLK),
						      .D_IN(cache_toCQ_enqReq_dummy2_0$D_IN),
						      .EN(cache_toCQ_enqReq_dummy2_0$EN),
						      .Q_OUT());
  // submodule cache_toCQ_enqReq_dummy2_1
  RevertReg #(.width(32'd1),
	      .init(1'd1)) cache_toCQ_enqReq_dummy2_1(.CLK(CLK),
						      .D_IN(cache_toCQ_enqReq_dummy2_1$D_IN),
						      .EN(cache_toCQ_enqReq_dummy2_1$EN),
						      .Q_OUT());
  // submodule cache_toCQ_enqReq_dummy2_2
  RevertReg #(.width(32'd1),
	      .init(1'd1)) cache_toCQ_enqReq_dummy2_2(.CLK(CLK),
						      .D_IN(cache_toCQ_enqReq_dummy2_2$D_IN),
						      .EN(cache_toCQ_enqReq_dummy2_2$EN),
						      .Q_OUT(cache_toCQ_enqReq_dummy2_2$Q_OUT));
  // submodule cache_toMInfoQ
  SizedFIFO #(.p1width(32'd6),
	      .p2depth(32'd16),
	      .p3cntr_width(32'd4),
	      .guarded(1'd1)) cache_toMInfoQ(.RST(RST_N),
					     .CLK(CLK),
					     .D_IN(cache_toMInfoQ$D_IN),
					     .ENQ(cache_toMInfoQ$ENQ),
					     .DEQ(cache_toMInfoQ$DEQ),
					     .CLR(cache_toMInfoQ$CLR),
					     .D_OUT(cache_toMInfoQ$D_OUT),
					     .FULL_N(cache_toMInfoQ$FULL_N),
					     .EMPTY_N(cache_toMInfoQ$EMPTY_N));
  // submodule cache_toMQ_clearReq_dummy2_0
  RevertReg #(.width(32'd1),
	      .init(1'd1)) cache_toMQ_clearReq_dummy2_0(.CLK(CLK),
							.D_IN(cache_toMQ_clearReq_dummy2_0$D_IN),
							.EN(cache_toMQ_clearReq_dummy2_0$EN),
							.Q_OUT());
  // submodule cache_toMQ_clearReq_dummy2_1
  RevertReg #(.width(32'd1),
	      .init(1'd1)) cache_toMQ_clearReq_dummy2_1(.CLK(CLK),
							.D_IN(cache_toMQ_clearReq_dummy2_1$D_IN),
							.EN(cache_toMQ_clearReq_dummy2_1$EN),
							.Q_OUT(cache_toMQ_clearReq_dummy2_1$Q_OUT));
  // submodule cache_toMQ_deqReq_dummy2_0
  RevertReg #(.width(32'd1),
	      .init(1'd1)) cache_toMQ_deqReq_dummy2_0(.CLK(CLK),
						      .D_IN(cache_toMQ_deqReq_dummy2_0$D_IN),
						      .EN(cache_toMQ_deqReq_dummy2_0$EN),
						      .Q_OUT());
  // submodule cache_toMQ_deqReq_dummy2_1
  RevertReg #(.width(32'd1),
	      .init(1'd1)) cache_toMQ_deqReq_dummy2_1(.CLK(CLK),
						      .D_IN(cache_toMQ_deqReq_dummy2_1$D_IN),
						      .EN(cache_toMQ_deqReq_dummy2_1$EN),
						      .Q_OUT());
  // submodule cache_toMQ_deqReq_dummy2_2
  RevertReg #(.width(32'd1),
	      .init(1'd1)) cache_toMQ_deqReq_dummy2_2(.CLK(CLK),
						      .D_IN(cache_toMQ_deqReq_dummy2_2$D_IN),
						      .EN(cache_toMQ_deqReq_dummy2_2$EN),
						      .Q_OUT(cache_toMQ_deqReq_dummy2_2$Q_OUT));
  // submodule cache_toMQ_enqReq_dummy2_0
  RevertReg #(.width(32'd1),
	      .init(1'd1)) cache_toMQ_enqReq_dummy2_0(.CLK(CLK),
						      .D_IN(cache_toMQ_enqReq_dummy2_0$D_IN),
						      .EN(cache_toMQ_enqReq_dummy2_0$EN),
						      .Q_OUT());
  // submodule cache_toMQ_enqReq_dummy2_1
  RevertReg #(.width(32'd1),
	      .init(1'd1)) cache_toMQ_enqReq_dummy2_1(.CLK(CLK),
						      .D_IN(cache_toMQ_enqReq_dummy2_1$D_IN),
						      .EN(cache_toMQ_enqReq_dummy2_1$EN),
						      .Q_OUT());
  // submodule cache_toMQ_enqReq_dummy2_2
  RevertReg #(.width(32'd1),
	      .init(1'd1)) cache_toMQ_enqReq_dummy2_2(.CLK(CLK),
						      .D_IN(cache_toMQ_enqReq_dummy2_2$D_IN),
						      .EN(cache_toMQ_enqReq_dummy2_2$EN),
						      .Q_OUT(cache_toMQ_enqReq_dummy2_2$Q_OUT));
  // submodule perfReqQ_clearReq_dummy2_0
  RevertReg #(.width(32'd1),
	      .init(1'd1)) perfReqQ_clearReq_dummy2_0(.CLK(CLK),
						      .D_IN(perfReqQ_clearReq_dummy2_0$D_IN),
						      .EN(perfReqQ_clearReq_dummy2_0$EN),
						      .Q_OUT());
  // submodule perfReqQ_clearReq_dummy2_1
  RevertReg #(.width(32'd1),
	      .init(1'd1)) perfReqQ_clearReq_dummy2_1(.CLK(CLK),
						      .D_IN(perfReqQ_clearReq_dummy2_1$D_IN),
						      .EN(perfReqQ_clearReq_dummy2_1$EN),
						      .Q_OUT(perfReqQ_clearReq_dummy2_1$Q_OUT));
  // submodule perfReqQ_deqReq_dummy2_0
  RevertReg #(.width(32'd1), .init(1'd1)) perfReqQ_deqReq_dummy2_0(.CLK(CLK),
								   .D_IN(perfReqQ_deqReq_dummy2_0$D_IN),
								   .EN(perfReqQ_deqReq_dummy2_0$EN),
								   .Q_OUT());
  // submodule perfReqQ_deqReq_dummy2_1
  RevertReg #(.width(32'd1), .init(1'd1)) perfReqQ_deqReq_dummy2_1(.CLK(CLK),
								   .D_IN(perfReqQ_deqReq_dummy2_1$D_IN),
								   .EN(perfReqQ_deqReq_dummy2_1$EN),
								   .Q_OUT());
  // submodule perfReqQ_deqReq_dummy2_2
  RevertReg #(.width(32'd1), .init(1'd1)) perfReqQ_deqReq_dummy2_2(.CLK(CLK),
								   .D_IN(perfReqQ_deqReq_dummy2_2$D_IN),
								   .EN(perfReqQ_deqReq_dummy2_2$EN),
								   .Q_OUT(perfReqQ_deqReq_dummy2_2$Q_OUT));
  // submodule perfReqQ_enqReq_dummy2_0
  RevertReg #(.width(32'd1), .init(1'd1)) perfReqQ_enqReq_dummy2_0(.CLK(CLK),
								   .D_IN(perfReqQ_enqReq_dummy2_0$D_IN),
								   .EN(perfReqQ_enqReq_dummy2_0$EN),
								   .Q_OUT());
  // submodule perfReqQ_enqReq_dummy2_1
  RevertReg #(.width(32'd1), .init(1'd1)) perfReqQ_enqReq_dummy2_1(.CLK(CLK),
								   .D_IN(perfReqQ_enqReq_dummy2_1$D_IN),
								   .EN(perfReqQ_enqReq_dummy2_1$EN),
								   .Q_OUT());
  // submodule perfReqQ_enqReq_dummy2_2
  RevertReg #(.width(32'd1), .init(1'd1)) perfReqQ_enqReq_dummy2_2(.CLK(CLK),
								   .D_IN(perfReqQ_enqReq_dummy2_2$D_IN),
								   .EN(perfReqQ_enqReq_dummy2_2$EN),
								   .Q_OUT(perfReqQ_enqReq_dummy2_2$Q_OUT));
  // rule RL_cache_mergeRsLdToDmaIndexQ_mRsDeq
  assign CAN_FIRE_RL_cache_mergeRsLdToDmaIndexQ_mRsDeq =
	     cache_rsLdToDmaIndexQ_mRsDeq$EMPTY_N &&
	     cache_rsLdToDmaIndexQ$FULL_N ;
  assign WILL_FIRE_RL_cache_mergeRsLdToDmaIndexQ_mRsDeq =
	     CAN_FIRE_RL_cache_mergeRsLdToDmaIndexQ_mRsDeq &&
	     !WILL_FIRE_RL_cache_mergeRsLdToDmaIndexQ_pipelineResp ;
  // rule RL_cache_mergeRsLdToDmaIndexQ_pipelineResp
  assign CAN_FIRE_RL_cache_mergeRsLdToDmaIndexQ_pipelineResp =
	     cache_rsLdToDmaIndexQ$FULL_N &&
	     cache_rsLdToDmaIndexQ_pipelineResp$EMPTY_N ;
  assign WILL_FIRE_RL_cache_mergeRsLdToDmaIndexQ_pipelineResp =
	     CAN_FIRE_RL_cache_mergeRsLdToDmaIndexQ_pipelineResp ;
  // rule RL_cache_mergeRsStToDmaIndexQ_sendToM
  assign CAN_FIRE_RL_cache_mergeRsStToDmaIndexQ_sendToM =
	     cache_rsStToDmaIndexQ_sendToM$EMPTY_N &&
	     cache_rsStToDmaIndexQ$FULL_N ;
  assign WILL_FIRE_RL_cache_mergeRsStToDmaIndexQ_sendToM =
	     CAN_FIRE_RL_cache_mergeRsStToDmaIndexQ_sendToM &&
	     !WILL_FIRE_RL_cache_mergeRsStToDmaIndexQ_pipelineResp ;
  // rule RL_cache_mergeRsStToDmaIndexQ_pipelineResp
  assign CAN_FIRE_RL_cache_mergeRsStToDmaIndexQ_pipelineResp =
	     cache_rsStToDmaIndexQ$FULL_N &&
	     cache_rsStToDmaIndexQ_pipelineResp$EMPTY_N ;
  assign WILL_FIRE_RL_cache_mergeRsStToDmaIndexQ_pipelineResp =
	     CAN_FIRE_RL_cache_mergeRsStToDmaIndexQ_pipelineResp ;
  // rule RL_cache_sendToM
  assign CAN_FIRE_RL_cache_sendToM =
	     cache_toMInfoQ$EMPTY_N &&
	     CASE_cache_toMInfoQD_OUT_BITS_1_TO_0_0_NOT_ca_ETC__q264 ;
  assign WILL_FIRE_RL_cache_sendToM = CAN_FIRE_RL_cache_sendToM ;
  // rule RL_cache_sendRsToC
  assign CAN_FIRE_RL_cache_sendRsToC =
	     !cache_toCQ_full && !cache_rsToCIndexQ_empty &&
	     cache_cRqMshr$RDY_sendRsToDmaC_releaseEntry ;
  assign WILL_FIRE_RL_cache_sendRsToC =
	     CAN_FIRE_RL_cache_sendRsToC &&
	     !WILL_FIRE_RL_cache_sendRsStToDma &&
	     !WILL_FIRE_RL_cache_sendRsLdToDma ;
  // rule RL_cache_sendRqToC
  assign CAN_FIRE_RL_cache_sendRqToC =
	     !cache_toCQ_full &&
	     cache_cRqMshr_sendRqToC_searchNeedRqChild_1_CO_ETC___d2482 &&
	     cache_rsToCIndexQ_empty ;
  assign WILL_FIRE_RL_cache_sendRqToC = CAN_FIRE_RL_cache_sendRqToC ;
  // rule RL_cache_sendRsLdToDma
  assign CAN_FIRE_RL_cache_sendRsLdToDma =
	     !cache_rsLdToDmaQ_full &&
	     cache_cRqMshr$RDY_sendRsToDmaC_releaseEntry &&
	     cache_rsLdToDmaIndexQ$EMPTY_N ;
  assign WILL_FIRE_RL_cache_sendRsLdToDma = CAN_FIRE_RL_cache_sendRsLdToDma ;
  // rule RL_cache_mRsDeq_nonRefill
  assign CAN_FIRE_RL_cache_mRsDeq_nonRefill =
	     !cache_rsFromMQ_empty && cache_rsLdToDmaIndexQ_mRsDeq$FULL_N &&
	     CASE_cache_rsFromMQ_deqP_0_NOT_cache_rsFromMQ__ETC__q263 ;
  assign WILL_FIRE_RL_cache_mRsDeq_nonRefill =
	     CAN_FIRE_RL_cache_mRsDeq_nonRefill ;
  // rule RL_cache_sendRsStToDma
  assign CAN_FIRE_RL_cache_sendRsStToDma =
	     !cache_rsStToDmaQ_full &&
	     cache_cRqMshr$RDY_sendRsToDmaC_releaseEntry &&
	     cache_rsStToDmaIndexQ$EMPTY_N ;
  assign WILL_FIRE_RL_cache_sendRsStToDma =
	     CAN_FIRE_RL_cache_sendRsStToDma &&
	     !WILL_FIRE_RL_cache_sendRsLdToDma ;
  // rule RL_cache_pipelineResp_cRq
  assign CAN_FIRE_RL_cache_pipelineResp_cRq =
	     cache_pipeline$RDY_first &&
	     cache_pipeline_RDY_deqWrite__580_AND_IF_cache__ETC___d2671 &&
	     cache_pipeline$first[584:583] == 2'd0 ;
  assign WILL_FIRE_RL_cache_pipelineResp_cRq =
	     CAN_FIRE_RL_cache_pipelineResp_cRq ;
  // rule RL_cache_pipelineResp_mRs
  assign CAN_FIRE_RL_cache_pipelineResp_mRs =
	     !cache_rsToCIndexQ_full && cache_pipeline$RDY_first &&
	     cache_pipeline$RDY_deqWrite &&
	     cache_pipeline$first[584:583] == 2'd2 ;
  assign WILL_FIRE_RL_cache_pipelineResp_mRs =
	     CAN_FIRE_RL_cache_pipelineResp_mRs ;
  // rule RL_cache_pipelineResp_cRs
  assign CAN_FIRE_RL_cache_pipelineResp_cRs =
	     cache_pipeline$RDY_first &&
	     cache_pipeline_RDY_deqWrite__580_AND_NOT_cache_ETC___d3471 &&
	     cache_pipeline$first[584:583] == 2'd1 ;
  assign WILL_FIRE_RL_cache_pipelineResp_cRs =
	     CAN_FIRE_RL_cache_pipelineResp_cRs ;
  // rule RL_cache_cRqTransfer_retry
  assign CAN_FIRE_RL_cache_cRqTransfer_retry =
	     !cache_cRqRetryIndexQ_empty && cache_pipeline$RDY_send ;
  assign WILL_FIRE_RL_cache_cRqTransfer_retry =
	     CAN_FIRE_RL_cache_cRqTransfer_retry &&
	     !WILL_FIRE_RL_cache_cRsTransfer &&
	     !WILL_FIRE_RL_cache_mRsTransfer ;
  // rule RL_cache_cRqTransfer_new_child
  assign CAN_FIRE_RL_cache_cRqTransfer_new_child =
	     !cache_rqFromCQ_empty && cache_pipeline$RDY_send &&
	     cache_cRqMshr$RDY_transfer_getEmptyEntryInit &&
	     cache_cRqRetryIndexQ_empty &&
	     (!cache_priorNewCRqSrc || cache_rqFromDmaQ_empty) ;
  assign WILL_FIRE_RL_cache_cRqTransfer_new_child =
	     CAN_FIRE_RL_cache_cRqTransfer_new_child &&
	     !WILL_FIRE_RL_cache_cRsTransfer &&
	     !WILL_FIRE_RL_cache_mRsTransfer ;
  // rule RL_cache_cRqTransfer_new_dma
  assign CAN_FIRE_RL_cache_cRqTransfer_new_dma =
	     !cache_rqFromDmaQ_empty && cache_pipeline$RDY_send &&
	     cache_cRqMshr$RDY_transfer_getEmptyEntryInit &&
	     cache_cRqRetryIndexQ_empty &&
	     (cache_priorNewCRqSrc || cache_rqFromCQ_empty) ;
  assign WILL_FIRE_RL_cache_cRqTransfer_new_dma =
	     CAN_FIRE_RL_cache_cRqTransfer_new_dma &&
	     !WILL_FIRE_RL_cache_cRsTransfer &&
	     !WILL_FIRE_RL_cache_mRsTransfer ;
  // rule RL_cache_cRsTransfer
  assign CAN_FIRE_RL_cache_cRsTransfer =
	     !cache_rsFromCQ_empty && cache_pipeline$RDY_send ;
  assign WILL_FIRE_RL_cache_cRsTransfer =
	     CAN_FIRE_RL_cache_cRsTransfer &&
	     !WILL_FIRE_RL_cache_mRsTransfer ;
  // rule RL_cache_mRsTransfer
  assign CAN_FIRE_RL_cache_mRsTransfer =
	     !cache_rsFromMQ_empty && cache_pipeline$RDY_send &&
	     CASE_cache_rsFromMQ_deqP_0_cache_rsFromMQ_data_ETC__q262 ;
  assign WILL_FIRE_RL_cache_mRsTransfer = CAN_FIRE_RL_cache_mRsTransfer ;
  // rule RL_cache_rqFromCQ_canonicalize
  assign CAN_FIRE_RL_cache_rqFromCQ_canonicalize = 1'd1 ;
  assign WILL_FIRE_RL_cache_rqFromCQ_canonicalize = 1'd1 ;
  // rule RL_cache_rqFromCQ_enqReq_canon
  assign CAN_FIRE_RL_cache_rqFromCQ_enqReq_canon = 1'd1 ;
  assign WILL_FIRE_RL_cache_rqFromCQ_enqReq_canon = 1'd1 ;
  // rule RL_cache_rqFromCQ_deqReq_canon
  assign CAN_FIRE_RL_cache_rqFromCQ_deqReq_canon = 1'd1 ;
  assign WILL_FIRE_RL_cache_rqFromCQ_deqReq_canon = 1'd1 ;
  // rule RL_cache_rqFromCQ_clearReq_canon
  assign CAN_FIRE_RL_cache_rqFromCQ_clearReq_canon = 1'd1 ;
  assign WILL_FIRE_RL_cache_rqFromCQ_clearReq_canon = 1'd1 ;
  // rule RL_cache_rsFromCQ_canonicalize
  assign CAN_FIRE_RL_cache_rsFromCQ_canonicalize = 1'd1 ;
  assign WILL_FIRE_RL_cache_rsFromCQ_canonicalize = 1'd1 ;
  // rule RL_cache_rsFromCQ_enqReq_canon
  assign CAN_FIRE_RL_cache_rsFromCQ_enqReq_canon = 1'd1 ;
  assign WILL_FIRE_RL_cache_rsFromCQ_enqReq_canon = 1'd1 ;
  // rule RL_cache_rsFromCQ_deqReq_canon
  assign CAN_FIRE_RL_cache_rsFromCQ_deqReq_canon = 1'd1 ;
  assign WILL_FIRE_RL_cache_rsFromCQ_deqReq_canon = 1'd1 ;
  // rule RL_cache_rsFromCQ_clearReq_canon
  assign CAN_FIRE_RL_cache_rsFromCQ_clearReq_canon = 1'd1 ;
  assign WILL_FIRE_RL_cache_rsFromCQ_clearReq_canon = 1'd1 ;
  // rule RL_cache_toCQ_canonicalize
  assign CAN_FIRE_RL_cache_toCQ_canonicalize = 1'd1 ;
  assign WILL_FIRE_RL_cache_toCQ_canonicalize = 1'd1 ;
  // rule RL_cache_toCQ_enqReq_canon
  assign CAN_FIRE_RL_cache_toCQ_enqReq_canon = 1'd1 ;
  assign WILL_FIRE_RL_cache_toCQ_enqReq_canon = 1'd1 ;
  // rule RL_cache_toCQ_deqReq_canon
  assign CAN_FIRE_RL_cache_toCQ_deqReq_canon = 1'd1 ;
  assign WILL_FIRE_RL_cache_toCQ_deqReq_canon = 1'd1 ;
  // rule RL_cache_toCQ_clearReq_canon
  assign CAN_FIRE_RL_cache_toCQ_clearReq_canon = 1'd1 ;
  assign WILL_FIRE_RL_cache_toCQ_clearReq_canon = 1'd1 ;
  // rule RL_cache_rqFromDmaQ_canonicalize
  assign CAN_FIRE_RL_cache_rqFromDmaQ_canonicalize = 1'd1 ;
  assign WILL_FIRE_RL_cache_rqFromDmaQ_canonicalize = 1'd1 ;
  // rule RL_cache_rqFromDmaQ_enqReq_canon
  assign CAN_FIRE_RL_cache_rqFromDmaQ_enqReq_canon = 1'd1 ;
  assign WILL_FIRE_RL_cache_rqFromDmaQ_enqReq_canon = 1'd1 ;
  // rule RL_cache_rqFromDmaQ_deqReq_canon
  assign CAN_FIRE_RL_cache_rqFromDmaQ_deqReq_canon = 1'd1 ;
  assign WILL_FIRE_RL_cache_rqFromDmaQ_deqReq_canon = 1'd1 ;
  // rule RL_cache_rqFromDmaQ_clearReq_canon
  assign CAN_FIRE_RL_cache_rqFromDmaQ_clearReq_canon = 1'd1 ;
  assign WILL_FIRE_RL_cache_rqFromDmaQ_clearReq_canon = 1'd1 ;
  // rule RL_cache_rsLdToDmaQ_canonicalize
  assign CAN_FIRE_RL_cache_rsLdToDmaQ_canonicalize = 1'd1 ;
  assign WILL_FIRE_RL_cache_rsLdToDmaQ_canonicalize = 1'd1 ;
  // rule RL_cache_rsLdToDmaQ_enqReq_canon
  assign CAN_FIRE_RL_cache_rsLdToDmaQ_enqReq_canon = 1'd1 ;
  assign WILL_FIRE_RL_cache_rsLdToDmaQ_enqReq_canon = 1'd1 ;
  // rule RL_cache_rsLdToDmaQ_deqReq_canon
  assign CAN_FIRE_RL_cache_rsLdToDmaQ_deqReq_canon = 1'd1 ;
  assign WILL_FIRE_RL_cache_rsLdToDmaQ_deqReq_canon = 1'd1 ;
  // rule RL_cache_rsLdToDmaQ_clearReq_canon
  assign CAN_FIRE_RL_cache_rsLdToDmaQ_clearReq_canon = 1'd1 ;
  assign WILL_FIRE_RL_cache_rsLdToDmaQ_clearReq_canon = 1'd1 ;
  // rule RL_cache_rsStToDmaQ_canonicalize
  assign CAN_FIRE_RL_cache_rsStToDmaQ_canonicalize = 1'd1 ;
  assign WILL_FIRE_RL_cache_rsStToDmaQ_canonicalize = 1'd1 ;
  // rule RL_cache_rsStToDmaQ_enqReq_canon
  assign CAN_FIRE_RL_cache_rsStToDmaQ_enqReq_canon = 1'd1 ;
  assign WILL_FIRE_RL_cache_rsStToDmaQ_enqReq_canon = 1'd1 ;
  // rule RL_cache_rsStToDmaQ_deqReq_canon
  assign CAN_FIRE_RL_cache_rsStToDmaQ_deqReq_canon = 1'd1 ;
  assign WILL_FIRE_RL_cache_rsStToDmaQ_deqReq_canon = 1'd1 ;
  // rule RL_cache_rsStToDmaQ_clearReq_canon
  assign CAN_FIRE_RL_cache_rsStToDmaQ_clearReq_canon = 1'd1 ;
  assign WILL_FIRE_RL_cache_rsStToDmaQ_clearReq_canon = 1'd1 ;
  // rule RL_cache_toMQ_canonicalize
  assign CAN_FIRE_RL_cache_toMQ_canonicalize = 1'd1 ;
  assign WILL_FIRE_RL_cache_toMQ_canonicalize = 1'd1 ;
  // rule RL_cache_toMQ_enqReq_canon
  assign CAN_FIRE_RL_cache_toMQ_enqReq_canon = 1'd1 ;
  assign WILL_FIRE_RL_cache_toMQ_enqReq_canon = 1'd1 ;
  // rule RL_cache_toMQ_deqReq_canon
  assign CAN_FIRE_RL_cache_toMQ_deqReq_canon = 1'd1 ;
  assign WILL_FIRE_RL_cache_toMQ_deqReq_canon = 1'd1 ;
  // rule RL_cache_toMQ_clearReq_canon
  assign CAN_FIRE_RL_cache_toMQ_clearReq_canon = 1'd1 ;
  assign WILL_FIRE_RL_cache_toMQ_clearReq_canon = 1'd1 ;
  // rule RL_cache_rsFromMQ_canonicalize
  assign CAN_FIRE_RL_cache_rsFromMQ_canonicalize = 1'd1 ;
  assign WILL_FIRE_RL_cache_rsFromMQ_canonicalize = 1'd1 ;
  // rule RL_cache_rsFromMQ_enqReq_canon
  assign CAN_FIRE_RL_cache_rsFromMQ_enqReq_canon = 1'd1 ;
  assign WILL_FIRE_RL_cache_rsFromMQ_enqReq_canon = 1'd1 ;
  // rule RL_cache_rsFromMQ_deqReq_canon
  assign CAN_FIRE_RL_cache_rsFromMQ_deqReq_canon = 1'd1 ;
  assign WILL_FIRE_RL_cache_rsFromMQ_deqReq_canon = 1'd1 ;
  // rule RL_cache_rsFromMQ_clearReq_canon
  assign CAN_FIRE_RL_cache_rsFromMQ_clearReq_canon = 1'd1 ;
  assign WILL_FIRE_RL_cache_rsFromMQ_clearReq_canon = 1'd1 ;
  // rule RL_cache_cRqRetryIndexQ_canonicalize
  assign CAN_FIRE_RL_cache_cRqRetryIndexQ_canonicalize = 1'd1 ;
  assign WILL_FIRE_RL_cache_cRqRetryIndexQ_canonicalize = 1'd1 ;
  // rule RL_cache_cRqRetryIndexQ_enqReq_canon
  assign CAN_FIRE_RL_cache_cRqRetryIndexQ_enqReq_canon = 1'd1 ;
  assign WILL_FIRE_RL_cache_cRqRetryIndexQ_enqReq_canon = 1'd1 ;
  // rule RL_cache_cRqRetryIndexQ_deqReq_canon
  assign CAN_FIRE_RL_cache_cRqRetryIndexQ_deqReq_canon = 1'd1 ;
  assign WILL_FIRE_RL_cache_cRqRetryIndexQ_deqReq_canon = 1'd1 ;
  // rule RL_cache_cRqRetryIndexQ_clearReq_canon
  assign CAN_FIRE_RL_cache_cRqRetryIndexQ_clearReq_canon = 1'd1 ;
  assign WILL_FIRE_RL_cache_cRqRetryIndexQ_clearReq_canon = 1'd1 ;
  // rule RL_cache_rsToCIndexQ_canonicalize
  assign CAN_FIRE_RL_cache_rsToCIndexQ_canonicalize = 1'd1 ;
  assign WILL_FIRE_RL_cache_rsToCIndexQ_canonicalize = 1'd1 ;
  // rule RL_cache_rsToCIndexQ_enqReq_canon
  assign CAN_FIRE_RL_cache_rsToCIndexQ_enqReq_canon = 1'd1 ;
  assign WILL_FIRE_RL_cache_rsToCIndexQ_enqReq_canon = 1'd1 ;
  // rule RL_cache_rsToCIndexQ_deqReq_canon
  assign CAN_FIRE_RL_cache_rsToCIndexQ_deqReq_canon = 1'd1 ;
  assign WILL_FIRE_RL_cache_rsToCIndexQ_deqReq_canon = 1'd1 ;
  // rule RL_cache_rsToCIndexQ_clearReq_canon
  assign CAN_FIRE_RL_cache_rsToCIndexQ_clearReq_canon = 1'd1 ;
  assign WILL_FIRE_RL_cache_rsToCIndexQ_clearReq_canon = 1'd1 ;
  // rule RL_perfReqQ_canonicalize
  assign CAN_FIRE_RL_perfReqQ_canonicalize = 1'd1 ;
  assign WILL_FIRE_RL_perfReqQ_canonicalize = 1'd1 ;
  // rule RL_perfReqQ_enqReq_canon
  assign CAN_FIRE_RL_perfReqQ_enqReq_canon = 1'd1 ;
  assign WILL_FIRE_RL_perfReqQ_enqReq_canon = 1'd1 ;
  // rule RL_perfReqQ_deqReq_canon
  assign CAN_FIRE_RL_perfReqQ_deqReq_canon = 1'd1 ;
  assign WILL_FIRE_RL_perfReqQ_deqReq_canon = 1'd1 ;
  // rule RL_perfReqQ_clearReq_canon
  assign CAN_FIRE_RL_perfReqQ_clearReq_canon = 1'd1 ;
  assign WILL_FIRE_RL_perfReqQ_clearReq_canon = 1'd1 ;
  // inputs to muxes for submodule ports
  assign MUX_cache_cRqMshr$pipelineResp_setData_1__SEL_1 =
	     WILL_FIRE_RL_cache_pipelineResp_cRq &&
	     (cache_pipeline$first[517] &&
	      cache_pipeline_first__581_BITS_516_TO_513_583__ETC___d3103 ||
	      !cache_pipeline$first[517] &&
	      NOT_cache_cRqMshr_pipelineResp_searchEndOfChai_ETC___d3114) ;
  assign MUX_cache_cRqMshr$pipelineResp_setData_1__SEL_2 =
	     WILL_FIRE_RL_cache_pipelineResp_cRs &&
	     cache_pipeline$first[517] &&
	     (cache_pipeline$first[512] &&
	      IF_SEL_ARR_cache_pipeline_first__581_BITS_519__ETC___d3488 ||
	      !cache_pipeline$first[512] &&
	      IF_SEL_ARR_cache_cRqMshr_pipelineResp_getSlot__ETC___d3484) ;
  assign MUX_cache_cRqMshr$pipelineResp_setStateSlot_1__SEL_1 =
	     WILL_FIRE_RL_cache_pipelineResp_cRs &&
	     cache_pipeline$first[517] ;
  assign MUX_cache_cRqRetryIndexQ_enqReq_dummy2_0$write_1__SEL_1 =
	     WILL_FIRE_RL_cache_pipelineResp_cRq &&
	     NOT_cache_pipeline_first__581_BIT_517_582_105__ETC___d3332 ;
  assign MUX_cache_cRqRetryIndexQ_enqReq_dummy2_0$write_1__SEL_2 =
	     WILL_FIRE_RL_cache_pipelineResp_cRs &&
	     cache_pipeline$first[517] &&
	     cache_pipeline$first[512] &&
	     IF_SEL_ARR_cache_pipeline_first__581_BITS_519__ETC___d3488 &&
	     cache_cRqMshr$pipelineResp_getRepSucc[4] ;
  assign MUX_cache_rsLdToDmaIndexQ_pipelineResp$enq_1__SEL_1 =
	     WILL_FIRE_RL_cache_pipelineResp_cRq &&
	     (cache_pipeline_first__581_BIT_517_582_AND_cach_ETC___d3139 ||
	      NOT_cache_pipeline_first__581_BIT_517_582_105__ETC___d3143) ;
  assign MUX_cache_rsStToDmaIndexQ_pipelineResp$enq_1__SEL_1 =
	     WILL_FIRE_RL_cache_pipelineResp_cRq &&
	     (cache_pipeline_first__581_BIT_517_582_AND_cach_ETC___d3129 ||
	      NOT_cache_pipeline_first__581_BIT_517_582_105__ETC___d3133) ;
  assign MUX_cache_rsToCIndexQ_enqReq_dummy2_0$write_1__SEL_1 =
	     WILL_FIRE_RL_cache_pipelineResp_cRq &&
	     (cache_pipeline_first__581_BIT_517_582_AND_cach_ETC___d3146 ||
	      NOT_cache_pipeline_first__581_BIT_517_582_105__ETC___d3149) ;
  assign MUX_cache_rsToCIndexQ_enqReq_dummy2_0$write_1__SEL_2 =
	     WILL_FIRE_RL_cache_pipelineResp_cRs &&
	     cache_pipeline$first[517] &&
	     !cache_pipeline$first[512] &&
	     IF_SEL_ARR_cache_cRqMshr_pipelineResp_getSlot__ETC___d3484 &&
	     !cache_cRqMshr$pipelineResp_getRq[16] ;
  assign MUX_cache_toMInfoQ$enq_1__SEL_1 =
	     WILL_FIRE_RL_cache_pipelineResp_cRq &&
	     (cache_pipeline$first[517] &&
	      cache_pipeline_first__581_BITS_516_TO_513_583__ETC___d2588 &&
	      !cache_cRqMshr$pipelineResp_getRq[16] &&
	      IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3156 &&
	      cache_pipeline$first[525:524] == 2'd0 ||
	      !cache_pipeline$first[517] &&
	      (!cache_cRqMshr$pipelineResp_searchEndOfChain[4] ||
	       cache_cRqMshr$pipelineResp_getState != 3'd1) &&
	      cache_cRqMshr_pipelineResp_getRq_IF_cache_pipe_ETC___d3166) ;
  always@(cache_rsToCIndexQ_deqP or
	  cache_rsToCIndexQ_data_0 or
	  cache_rsToCIndexQ_data_1 or
	  cache_rsToCIndexQ_data_2 or
	  cache_rsToCIndexQ_data_3 or
	  cache_rsToCIndexQ_data_4 or
	  cache_rsToCIndexQ_data_5 or
	  cache_rsToCIndexQ_data_6 or
	  cache_rsToCIndexQ_data_7 or
	  cache_rsToCIndexQ_data_8 or
	  cache_rsToCIndexQ_data_9 or
	  cache_rsToCIndexQ_data_10 or
	  cache_rsToCIndexQ_data_11 or
	  cache_rsToCIndexQ_data_12 or
	  cache_rsToCIndexQ_data_13 or
	  cache_rsToCIndexQ_data_14 or cache_rsToCIndexQ_data_15)
  begin
    case (cache_rsToCIndexQ_deqP)
      4'd0:
	  MUX_cache_cRqMshr$sendRsToDmaC_getData_1__VAL_2 =
	      cache_rsToCIndexQ_data_0[5:2];
      4'd1:
	  MUX_cache_cRqMshr$sendRsToDmaC_getData_1__VAL_2 =
	      cache_rsToCIndexQ_data_1[5:2];
      4'd2:
	  MUX_cache_cRqMshr$sendRsToDmaC_getData_1__VAL_2 =
	      cache_rsToCIndexQ_data_2[5:2];
      4'd3:
	  MUX_cache_cRqMshr$sendRsToDmaC_getData_1__VAL_2 =
	      cache_rsToCIndexQ_data_3[5:2];
      4'd4:
	  MUX_cache_cRqMshr$sendRsToDmaC_getData_1__VAL_2 =
	      cache_rsToCIndexQ_data_4[5:2];
      4'd5:
	  MUX_cache_cRqMshr$sendRsToDmaC_getData_1__VAL_2 =
	      cache_rsToCIndexQ_data_5[5:2];
      4'd6:
	  MUX_cache_cRqMshr$sendRsToDmaC_getData_1__VAL_2 =
	      cache_rsToCIndexQ_data_6[5:2];
      4'd7:
	  MUX_cache_cRqMshr$sendRsToDmaC_getData_1__VAL_2 =
	      cache_rsToCIndexQ_data_7[5:2];
      4'd8:
	  MUX_cache_cRqMshr$sendRsToDmaC_getData_1__VAL_2 =
	      cache_rsToCIndexQ_data_8[5:2];
      4'd9:
	  MUX_cache_cRqMshr$sendRsToDmaC_getData_1__VAL_2 =
	      cache_rsToCIndexQ_data_9[5:2];
      4'd10:
	  MUX_cache_cRqMshr$sendRsToDmaC_getData_1__VAL_2 =
	      cache_rsToCIndexQ_data_10[5:2];
      4'd11:
	  MUX_cache_cRqMshr$sendRsToDmaC_getData_1__VAL_2 =
	      cache_rsToCIndexQ_data_11[5:2];
      4'd12:
	  MUX_cache_cRqMshr$sendRsToDmaC_getData_1__VAL_2 =
	      cache_rsToCIndexQ_data_12[5:2];
      4'd13:
	  MUX_cache_cRqMshr$sendRsToDmaC_getData_1__VAL_2 =
	      cache_rsToCIndexQ_data_13[5:2];
      4'd14:
	  MUX_cache_cRqMshr$sendRsToDmaC_getData_1__VAL_2 =
	      cache_rsToCIndexQ_data_14[5:2];
      4'd15:
	  MUX_cache_cRqMshr$sendRsToDmaC_getData_1__VAL_2 =
	      cache_rsToCIndexQ_data_15[5:2];
    endcase
  end
  always@(cache_rsFromMQ_deqP or
	  cache_rsFromMQ_data_0 or cache_rsFromMQ_data_1)
  begin
    case (cache_rsFromMQ_deqP)
      1'd0:
	  MUX_cache_cRqMshr$transfer_getRq_1__VAL_2 =
	      cache_rsFromMQ_data_0[3:0];
      1'd1:
	  MUX_cache_cRqMshr$transfer_getRq_1__VAL_2 =
	      cache_rsFromMQ_data_1[3:0];
    endcase
  end
  assign MUX_cache_cRqMshr$pipelineResp_setData_2__VAL_1 =
	     { IF_cache_pipeline_first__581_BIT_517_582_THEN__ETC___d3124,
	       cache_pipeline$first[511:0] } ;
  assign MUX_cache_cRqMshr$pipelineResp_setData_2__VAL_2 =
	     { cache_pipeline$first[512] ?
		 cache_pipeline$first[525:524] == 2'd3 :
		 cache_cRqMshr$pipelineResp_getRq[16] ||
		 CASE_cache_cRqMshrpipelineResp_getRq_BITS_82__ETC__q79 ==
		 2'd0,
	       cache_pipeline$first[511:0] } ;
  assign MUX_cache_cRqMshr$pipelineResp_setData_2__VAL_3 =
	     { CASE_cache_cRqMshrpipelineResp_getRq_BITS_82__ETC__q79 == 2'd0,
	       cache_pipeline$first[511:0] } ;
  assign MUX_cache_cRqMshr$pipelineResp_setStateSlot_2__VAL_1 =
	     cache_pipeline$first[512] ?
	       (IF_SEL_ARR_cache_pipeline_first__581_BITS_519__ETC___d3488 ?
		  3'd3 :
		  3'd2) :
	       (IF_SEL_ARR_cache_cRqMshr_pipelineResp_getSlot__ETC___d3484 ?
		  3'd4 :
		  3'd3) ;
  assign MUX_cache_cRqMshr$pipelineResp_setStateSlot_2__VAL_2 =
	     cache_pipeline$first[517] ?
	       (cache_pipeline_first__581_BITS_516_TO_513_583__ETC___d2588 ?
		  IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3027 :
		  3'd5) :
	       ((cache_cRqMshr$pipelineResp_searchEndOfChain[4] &&
		 cache_cRqMshr$pipelineResp_getState == 3'd1) ?
		  3'd5 :
		  IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3033) ;
  assign MUX_cache_cRqMshr$pipelineResp_setStateSlot_3__VAL_1 =
	     cache_pipeline$first[512] ?
	       IF_IF_SEL_ARR_cache_pipeline_first__581_BITS_5_ETC___d3709 :
	       cache_cRqMshr_pipelineResp_getSlot_IF_cache_pi_ETC___d3754 ;
  assign MUX_cache_cRqMshr$pipelineResp_setStateSlot_3__VAL_2 =
	     cache_pipeline$first[517] ?
	       (cache_pipeline_first__581_BITS_516_TO_513_583__ETC___d2588 ?
		  IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3078 :
		  65'h15555555555554222) :
	       ((cache_cRqMshr$pipelineResp_searchEndOfChain[4] &&
		 cache_cRqMshr$pipelineResp_getState == 3'd1) ?
		  65'h15555555555554222 :
		  IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3096) ;
  assign MUX_cache_cRqMshr$transfer_getEmptyEntryInit_1__VAL_1 =
	     { addr__h257616,
	       CASE_cache_rqFromCQ_deqP_0_cache_rqFromCQ_data_ETC__q265,
	       SEL_ARR_cache_rqFromCQ_data_0_090_BITS_7_TO_6__ETC___d1118 } ;
  assign MUX_cache_cRqMshr$transfer_getEmptyEntryInit_1__VAL_2 =
	     { addr__h273361,
	       2'd0,
	       IF_NOT_SEL_ARR_NOT_cache_rqFromDmaQ_data_0_129_ETC___d1646,
	       3'd2,
	       SEL_ARR_cache_rqFromDmaQ_data_0_129_BIT_591_57_ETC___d1806,
	       1'd1,
	       CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q266 } ;
  assign MUX_cache_cRqMshr$transfer_getEmptyEntryInit_2__VAL_2 =
	     { !CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q68 ||
	       NOT_SEL_ARR_NOT_cache_rqFromDmaQ_data_0_129_BI_ETC___d1644,
	       SEL_ARR_cache_rqFromDmaQ_data_0_129_BITS_527_T_ETC___d1845,
	       CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q267 } ;
  assign MUX_cache_cRqRetryIndexQ_enqReq_lat_0$wset_1__VAL_1 =
	     { 1'd1, cache_cRqMshr$pipelineResp_getAddrSucc[3:0] } ;
  assign MUX_cache_cRqRetryIndexQ_enqReq_lat_0$wset_1__VAL_2 =
	     { 1'd1, cache_cRqMshr$pipelineResp_getRepSucc[3:0] } ;
  assign MUX_cache_pipeline$deqWrite_1__VAL_2 =
	     cache_pipeline$first[517] ?
	       (cache_pipeline_first__581_BITS_516_TO_513_583__ETC___d2588 ?
		  IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2678 :
		  5'd10) :
	       ((cache_cRqMshr$pipelineResp_searchEndOfChain[4] &&
		 cache_cRqMshr$pipelineResp_getState == 3'd1) ?
		  5'd10 :
		  IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2683) ;
  assign MUX_cache_pipeline$deqWrite_1__VAL_3 =
	     cache_pipeline$first[517] ?
	       IF_cache_pipeline_first__581_BIT_512_308_THEN__ETC___d3486 :
	       5'd10 ;
  assign MUX_cache_pipeline$deqWrite_2__VAL_1 =
	     { cache_cRqMshr$pipelineResp_getRq[151:104],
	       IF_IF_cache_cRqMshr_pipelineResp_getRq_IF_cach_ETC___d3397,
	       cache_pipeline$first[511:0] } ;
  assign MUX_cache_pipeline$deqWrite_2__VAL_2 =
	     cache_pipeline$first[517] ?
	       (cache_pipeline_first__581_BITS_516_TO_513_583__ETC___d2588 ?
		  cache_cRqMshr_pipelineResp_getRq_IF_cache_pipe_ETC___d2995 :
		  cache_pipeline$first[573:0]) :
	       IF_cache_cRqMshr_pipelineResp_searchEndOfChain_ETC___d3012 ;
  assign MUX_cache_pipeline$deqWrite_2__VAL_3 =
	     cache_pipeline$first[517] ?
	       IF_cache_pipeline_first__581_BIT_512_308_THEN__ETC___d3660 :
	       cache_pipeline$first[573:0] ;
  assign MUX_cache_pipeline$deqWrite_3__VAL_2 =
	     cache_pipeline$first[517] ?
	       cache_pipeline_first__581_BITS_516_TO_513_583__ETC___d2588 &&
	       IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3014 :
	       (!cache_cRqMshr$pipelineResp_searchEndOfChain[4] ||
		cache_cRqMshr$pipelineResp_getState != 3'd1) &&
	       IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3022 ;
  assign MUX_cache_pipeline$deqWrite_3__VAL_3 =
	     cache_pipeline$first[517] && !cache_pipeline$first[512] &&
	     IF_SEL_ARR_cache_cRqMshr_pipelineResp_getSlot__ETC___d3484 ;
  assign MUX_cache_pipeline$send_1__VAL_1 =
	     { 516'h2AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA,
	       cache_cRqMshr$transfer_getRq[151:88],
	       x__h248737 } ;
  assign MUX_cache_pipeline$send_1__VAL_2 =
	     { 516'h2AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA,
	       addr__h257616,
	       cache_cRqMshr$transfer_getEmptyEntryInit } ;
  assign MUX_cache_pipeline$send_1__VAL_3 =
	     { 516'h2AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA,
	       addr__h273361,
	       cache_cRqMshr$transfer_getEmptyEntryInit } ;
  assign MUX_cache_pipeline$send_1__VAL_4 =
	     { 3'd2,
	       SEL_ARR_cache_rsFromCQ_data_0_855_BITS_580_TO__ETC___d1910 } ;
  assign MUX_cache_pipeline$send_1__VAL_5 =
	     { 2'd2,
	       cache_cRqMshr$transfer_getRq[151:88],
	       (cache_cRqMshr$transfer_getRq[85:84] == 2'd3) ?
		 cache_cRqMshr$transfer_getRq[85:84] :
		 2'd2,
	       SEL_ARR_cache_rsFromMQ_data_0_914_BITS_516_TO__ETC___d1966,
	       cache_cRqMshr$transfer_getSlot[64:61] } ;
  assign MUX_cache_rsToCIndexQ_enqReq_lat_0$wset_1__VAL_1 =
	     { 1'd1,
	       cache_pipeline$first[582:579],
	       cache_cRqMshr$pipelineResp_getRq[85:84] } ;
  assign MUX_cache_rsToCIndexQ_enqReq_lat_0$wset_1__VAL_2 =
	     { 1'd1,
	       cache_pipeline$first[516:513],
	       cache_cRqMshr$pipelineResp_getRq[85:84] } ;
  assign MUX_cache_rsToCIndexQ_enqReq_lat_0$wset_1__VAL_3 =
	     { 1'd1,
	       cache_pipeline$first[516:513],
	       IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3388 } ;
  assign MUX_cache_toCQ_enqReq_lat_0$wset_1__VAL_1 =
	     { 2'd3,
	       cache_cRqMshr$sendRsToDmaC_getRq[151:88],
	       SEL_ARR_cache_rsToCIndexQ_data_0_391_BITS_1_TO_ETC___d2445,
	       cache_cRqMshr$sendRsToDmaC_getRq[82:81],
	       cache_cRqMshr$sendRsToDmaC_getData,
	       cache_cRqMshr$sendRsToDmaC_getRq[2:0] } ;
  assign MUX_cache_toCQ_enqReq_lat_0$wset_1__VAL_2 =
	     { 518'h2AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA,
	       rqAddr__h313360,
	       SEL_ARR_IF_cache_cRqMshr_sendRqToC_getSlot_IF__ETC___d2522,
	       (cache_cRqMshr$sendRqToC_getSlot[3:2] != 2'd1 &&
		cache_cRqMshr$sendRqToC_getSlot[7:6] != 2'd1) ?
		 2'd2 :
		 ((cache_cRqMshr$sendRqToC_getSlot[3:2] == 2'd1) ?
		    2'd0 :
		    2'd1) } ;
  assign MUX_cache_toMInfoQ$enq_1__VAL_1 =
	     { cache_pipeline$first[582:579],
	       cache_pipeline$first[517] ?
		 2'd0 :
		 IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3173 } ;
  assign MUX_cache_toMInfoQ$enq_1__VAL_2 =
	     { cache_pipeline$first[516:513],
	       IF_cache_pipeline_first__581_BITS_525_TO_524_6_ETC___d3171 } ;
  // inlined wires
  assign cache_rqFromCQ_enqReq_lat_0$wget = { 1'd1, to_child_rqFromC_enq_x } ;
  assign cache_rsFromCQ_enqReq_lat_0$wget = { 1'd1, to_child_rsFromC_enq_x } ;
  assign cache_toCQ_enqReq_lat_0$wget =
	     WILL_FIRE_RL_cache_sendRsToC ?
	       MUX_cache_toCQ_enqReq_lat_0$wset_1__VAL_1 :
	       MUX_cache_toCQ_enqReq_lat_0$wset_1__VAL_2 ;
  assign cache_toCQ_enqReq_lat_0$whas =
	     WILL_FIRE_RL_cache_sendRsToC || WILL_FIRE_RL_cache_sendRqToC ;
  assign cache_rqFromDmaQ_enqReq_lat_0$wget = { 1'd1, dma_memReq_enq_x } ;
  assign cache_rsLdToDmaQ_enqReq_lat_0$wget =
	     { 1'd1,
	       cache_cRqMshr$sendRsToDmaC_getData[511:0],
	       cache_cRqMshr$sendRsToDmaC_getRq[15:0] } ;
  assign cache_rsStToDmaQ_enqReq_lat_0$wget =
	     { 1'd1, cache_cRqMshr$sendRsToDmaC_getRq[15:0] } ;
  always@(cache_toMInfoQ$D_OUT or
	  IF_cache_doLdAfterReplace_007_THEN_2_CONCAT_DO_ETC___d2016 or
	  cache_cRqMshr$sendToM_getRq or cache_cRqMshr$sendToM_getData)
  begin
    case (cache_toMInfoQ$D_OUT[1:0])
      2'd0:
	  cache_toMQ_enqReq_lat_0$wget =
	      { 573'h12AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA,
		cache_cRqMshr$sendToM_getRq[151:88],
		!cache_cRqMshr$sendToM_getRq[16],
		cache_toMInfoQ$D_OUT[5:2] };
      2'd1:
	  cache_toMQ_enqReq_lat_0$wget =
	      { 2'd3,
		cache_cRqMshr$sendToM_getRq[151:88],
		cache_cRqMshr$sendToM_getRq[80:17],
		cache_cRqMshr$sendToM_getData[511:0] };
      default: cache_toMQ_enqReq_lat_0$wget =
		   IF_cache_doLdAfterReplace_007_THEN_2_CONCAT_DO_ETC___d2016;
    endcase
  end
  assign cache_toMQ_enqReq_lat_0$whas =
	     WILL_FIRE_RL_cache_sendToM &&
	     (cache_toMInfoQ$D_OUT[1:0] == 2'd0 ||
	      cache_toMInfoQ$D_OUT[1:0] == 2'd1 ||
	      cache_toMInfoQ$D_OUT[1:0] == 2'd2) ;
  assign cache_rsFromMQ_enqReq_lat_0$wget = { 1'd1, to_mem_rsFromM_enq_x } ;
  assign cache_rsFromMQ_deqReq_lat_0$whas =
	     WILL_FIRE_RL_cache_mRsDeq_nonRefill ||
	     WILL_FIRE_RL_cache_mRsTransfer ;
  assign cache_cRqRetryIndexQ_enqReq_lat_0$wget =
	     MUX_cache_cRqRetryIndexQ_enqReq_dummy2_0$write_1__SEL_1 ?
	       MUX_cache_cRqRetryIndexQ_enqReq_lat_0$wset_1__VAL_1 :
	       MUX_cache_cRqRetryIndexQ_enqReq_lat_0$wset_1__VAL_2 ;
  assign cache_cRqRetryIndexQ_enqReq_lat_0$whas =
	     MUX_cache_cRqRetryIndexQ_enqReq_dummy2_0$write_1__SEL_1 ||
	     MUX_cache_cRqRetryIndexQ_enqReq_dummy2_0$write_1__SEL_2 ;
  always@(MUX_cache_rsToCIndexQ_enqReq_dummy2_0$write_1__SEL_1 or
	  MUX_cache_rsToCIndexQ_enqReq_lat_0$wset_1__VAL_1 or
	  MUX_cache_rsToCIndexQ_enqReq_dummy2_0$write_1__SEL_2 or
	  MUX_cache_rsToCIndexQ_enqReq_lat_0$wset_1__VAL_2 or
	  WILL_FIRE_RL_cache_pipelineResp_mRs or
	  MUX_cache_rsToCIndexQ_enqReq_lat_0$wset_1__VAL_3)
  begin
    case (1'b1) // synopsys parallel_case
      MUX_cache_rsToCIndexQ_enqReq_dummy2_0$write_1__SEL_1:
	  cache_rsToCIndexQ_enqReq_lat_0$wget =
	      MUX_cache_rsToCIndexQ_enqReq_lat_0$wset_1__VAL_1;
      MUX_cache_rsToCIndexQ_enqReq_dummy2_0$write_1__SEL_2:
	  cache_rsToCIndexQ_enqReq_lat_0$wget =
	      MUX_cache_rsToCIndexQ_enqReq_lat_0$wset_1__VAL_2;
      WILL_FIRE_RL_cache_pipelineResp_mRs:
	  cache_rsToCIndexQ_enqReq_lat_0$wget =
	      MUX_cache_rsToCIndexQ_enqReq_lat_0$wset_1__VAL_3;
      default: cache_rsToCIndexQ_enqReq_lat_0$wget =
		   7'b0101010 /* unspecified value */ ;
    endcase
  end
  assign cache_rsToCIndexQ_enqReq_lat_0$whas =
	     MUX_cache_rsToCIndexQ_enqReq_dummy2_0$write_1__SEL_1 ||
	     MUX_cache_rsToCIndexQ_enqReq_dummy2_0$write_1__SEL_2 ||
	     WILL_FIRE_RL_cache_pipelineResp_mRs ;
  assign perfReqQ_enqReq_lat_0$wget = { 1'd1, perf_req_r } ;
  // register cache_cRqRetryIndexQ_clearReq_rl
  assign cache_cRqRetryIndexQ_clearReq_rl$D_IN = 1'd0 ;
  assign cache_cRqRetryIndexQ_clearReq_rl$EN = 1'd1 ;
  // register cache_cRqRetryIndexQ_data_0
  assign cache_cRqRetryIndexQ_data_0$D_IN =
	     cache_cRqRetryIndexQ_enqReq_lat_0$whas ?
	       cache_cRqRetryIndexQ_enqReq_lat_0$wget[3:0] :
	       cache_cRqRetryIndexQ_enqReq_rl[3:0] ;
  assign cache_cRqRetryIndexQ_data_0$EN =
	     cache_cRqRetryIndexQ_enqP == 4'd0 &&
	     NOT_cache_cRqRetryIndexQ_clearReq_dummy2_1_rea_ETC___d853 &&
	     cache_cRqRetryIndexQ_enqReq_dummy2_2$Q_OUT &&
	     IF_cache_cRqRetryIndexQ_enqReq_lat_1_whas__01__ETC___d833 ;
  // register cache_cRqRetryIndexQ_data_1
  assign cache_cRqRetryIndexQ_data_1$D_IN = cache_cRqRetryIndexQ_data_0$D_IN ;
  assign cache_cRqRetryIndexQ_data_1$EN =
	     cache_cRqRetryIndexQ_enqP == 4'd1 &&
	     NOT_cache_cRqRetryIndexQ_clearReq_dummy2_1_rea_ETC___d853 &&
	     cache_cRqRetryIndexQ_enqReq_dummy2_2$Q_OUT &&
	     IF_cache_cRqRetryIndexQ_enqReq_lat_1_whas__01__ETC___d833 ;
  // register cache_cRqRetryIndexQ_data_10
  assign cache_cRqRetryIndexQ_data_10$D_IN =
	     cache_cRqRetryIndexQ_data_0$D_IN ;
  assign cache_cRqRetryIndexQ_data_10$EN =
	     cache_cRqRetryIndexQ_enqP == 4'd10 &&
	     NOT_cache_cRqRetryIndexQ_clearReq_dummy2_1_rea_ETC___d853 &&
	     cache_cRqRetryIndexQ_enqReq_dummy2_2$Q_OUT &&
	     IF_cache_cRqRetryIndexQ_enqReq_lat_1_whas__01__ETC___d833 ;
  // register cache_cRqRetryIndexQ_data_11
  assign cache_cRqRetryIndexQ_data_11$D_IN =
	     cache_cRqRetryIndexQ_data_0$D_IN ;
  assign cache_cRqRetryIndexQ_data_11$EN =
	     cache_cRqRetryIndexQ_enqP == 4'd11 &&
	     NOT_cache_cRqRetryIndexQ_clearReq_dummy2_1_rea_ETC___d853 &&
	     cache_cRqRetryIndexQ_enqReq_dummy2_2$Q_OUT &&
	     IF_cache_cRqRetryIndexQ_enqReq_lat_1_whas__01__ETC___d833 ;
  // register cache_cRqRetryIndexQ_data_12
  assign cache_cRqRetryIndexQ_data_12$D_IN =
	     cache_cRqRetryIndexQ_data_0$D_IN ;
  assign cache_cRqRetryIndexQ_data_12$EN =
	     cache_cRqRetryIndexQ_enqP == 4'd12 &&
	     NOT_cache_cRqRetryIndexQ_clearReq_dummy2_1_rea_ETC___d853 &&
	     cache_cRqRetryIndexQ_enqReq_dummy2_2$Q_OUT &&
	     IF_cache_cRqRetryIndexQ_enqReq_lat_1_whas__01__ETC___d833 ;
  // register cache_cRqRetryIndexQ_data_13
  assign cache_cRqRetryIndexQ_data_13$D_IN =
	     cache_cRqRetryIndexQ_data_0$D_IN ;
  assign cache_cRqRetryIndexQ_data_13$EN =
	     cache_cRqRetryIndexQ_enqP == 4'd13 &&
	     NOT_cache_cRqRetryIndexQ_clearReq_dummy2_1_rea_ETC___d853 &&
	     cache_cRqRetryIndexQ_enqReq_dummy2_2$Q_OUT &&
	     IF_cache_cRqRetryIndexQ_enqReq_lat_1_whas__01__ETC___d833 ;
  // register cache_cRqRetryIndexQ_data_14
  assign cache_cRqRetryIndexQ_data_14$D_IN =
	     cache_cRqRetryIndexQ_data_0$D_IN ;
  assign cache_cRqRetryIndexQ_data_14$EN =
	     cache_cRqRetryIndexQ_enqP == 4'd14 &&
	     NOT_cache_cRqRetryIndexQ_clearReq_dummy2_1_rea_ETC___d853 &&
	     cache_cRqRetryIndexQ_enqReq_dummy2_2$Q_OUT &&
	     IF_cache_cRqRetryIndexQ_enqReq_lat_1_whas__01__ETC___d833 ;
  // register cache_cRqRetryIndexQ_data_15
  assign cache_cRqRetryIndexQ_data_15$D_IN =
	     cache_cRqRetryIndexQ_data_0$D_IN ;
  assign cache_cRqRetryIndexQ_data_15$EN =
	     cache_cRqRetryIndexQ_enqP == 4'd15 &&
	     NOT_cache_cRqRetryIndexQ_clearReq_dummy2_1_rea_ETC___d853 &&
	     cache_cRqRetryIndexQ_enqReq_dummy2_2$Q_OUT &&
	     IF_cache_cRqRetryIndexQ_enqReq_lat_1_whas__01__ETC___d833 ;
  // register cache_cRqRetryIndexQ_data_2
  assign cache_cRqRetryIndexQ_data_2$D_IN = cache_cRqRetryIndexQ_data_0$D_IN ;
  assign cache_cRqRetryIndexQ_data_2$EN =
	     cache_cRqRetryIndexQ_enqP == 4'd2 &&
	     NOT_cache_cRqRetryIndexQ_clearReq_dummy2_1_rea_ETC___d853 &&
	     cache_cRqRetryIndexQ_enqReq_dummy2_2$Q_OUT &&
	     IF_cache_cRqRetryIndexQ_enqReq_lat_1_whas__01__ETC___d833 ;
  // register cache_cRqRetryIndexQ_data_3
  assign cache_cRqRetryIndexQ_data_3$D_IN = cache_cRqRetryIndexQ_data_0$D_IN ;
  assign cache_cRqRetryIndexQ_data_3$EN =
	     cache_cRqRetryIndexQ_enqP == 4'd3 &&
	     NOT_cache_cRqRetryIndexQ_clearReq_dummy2_1_rea_ETC___d853 &&
	     cache_cRqRetryIndexQ_enqReq_dummy2_2$Q_OUT &&
	     IF_cache_cRqRetryIndexQ_enqReq_lat_1_whas__01__ETC___d833 ;
  // register cache_cRqRetryIndexQ_data_4
  assign cache_cRqRetryIndexQ_data_4$D_IN = cache_cRqRetryIndexQ_data_0$D_IN ;
  assign cache_cRqRetryIndexQ_data_4$EN =
	     cache_cRqRetryIndexQ_enqP == 4'd4 &&
	     NOT_cache_cRqRetryIndexQ_clearReq_dummy2_1_rea_ETC___d853 &&
	     cache_cRqRetryIndexQ_enqReq_dummy2_2$Q_OUT &&
	     IF_cache_cRqRetryIndexQ_enqReq_lat_1_whas__01__ETC___d833 ;
  // register cache_cRqRetryIndexQ_data_5
  assign cache_cRqRetryIndexQ_data_5$D_IN = cache_cRqRetryIndexQ_data_0$D_IN ;
  assign cache_cRqRetryIndexQ_data_5$EN =
	     cache_cRqRetryIndexQ_enqP == 4'd5 &&
	     NOT_cache_cRqRetryIndexQ_clearReq_dummy2_1_rea_ETC___d853 &&
	     cache_cRqRetryIndexQ_enqReq_dummy2_2$Q_OUT &&
	     IF_cache_cRqRetryIndexQ_enqReq_lat_1_whas__01__ETC___d833 ;
  // register cache_cRqRetryIndexQ_data_6
  assign cache_cRqRetryIndexQ_data_6$D_IN = cache_cRqRetryIndexQ_data_0$D_IN ;
  assign cache_cRqRetryIndexQ_data_6$EN =
	     cache_cRqRetryIndexQ_enqP == 4'd6 &&
	     NOT_cache_cRqRetryIndexQ_clearReq_dummy2_1_rea_ETC___d853 &&
	     cache_cRqRetryIndexQ_enqReq_dummy2_2$Q_OUT &&
	     IF_cache_cRqRetryIndexQ_enqReq_lat_1_whas__01__ETC___d833 ;
  // register cache_cRqRetryIndexQ_data_7
  assign cache_cRqRetryIndexQ_data_7$D_IN = cache_cRqRetryIndexQ_data_0$D_IN ;
  assign cache_cRqRetryIndexQ_data_7$EN =
	     cache_cRqRetryIndexQ_enqP == 4'd7 &&
	     NOT_cache_cRqRetryIndexQ_clearReq_dummy2_1_rea_ETC___d853 &&
	     cache_cRqRetryIndexQ_enqReq_dummy2_2$Q_OUT &&
	     IF_cache_cRqRetryIndexQ_enqReq_lat_1_whas__01__ETC___d833 ;
  // register cache_cRqRetryIndexQ_data_8
  assign cache_cRqRetryIndexQ_data_8$D_IN = cache_cRqRetryIndexQ_data_0$D_IN ;
  assign cache_cRqRetryIndexQ_data_8$EN =
	     cache_cRqRetryIndexQ_enqP == 4'd8 &&
	     NOT_cache_cRqRetryIndexQ_clearReq_dummy2_1_rea_ETC___d853 &&
	     cache_cRqRetryIndexQ_enqReq_dummy2_2$Q_OUT &&
	     IF_cache_cRqRetryIndexQ_enqReq_lat_1_whas__01__ETC___d833 ;
  // register cache_cRqRetryIndexQ_data_9
  assign cache_cRqRetryIndexQ_data_9$D_IN = cache_cRqRetryIndexQ_data_0$D_IN ;
  assign cache_cRqRetryIndexQ_data_9$EN =
	     cache_cRqRetryIndexQ_enqP == 4'd9 &&
	     NOT_cache_cRqRetryIndexQ_clearReq_dummy2_1_rea_ETC___d853 &&
	     cache_cRqRetryIndexQ_enqReq_dummy2_2$Q_OUT &&
	     IF_cache_cRqRetryIndexQ_enqReq_lat_1_whas__01__ETC___d833 ;
  // register cache_cRqRetryIndexQ_deqP
  assign cache_cRqRetryIndexQ_deqP$D_IN =
	     (cache_cRqRetryIndexQ_clearReq_dummy2_1$Q_OUT &&
	      cache_cRqRetryIndexQ_clearReq_rl) ?
	       4'd0 :
	       _theResult_____2__h234513 ;
  assign cache_cRqRetryIndexQ_deqP$EN = 1'd1 ;
  // register cache_cRqRetryIndexQ_deqReq_rl
  assign cache_cRqRetryIndexQ_deqReq_rl$D_IN = 1'd0 ;
  assign cache_cRqRetryIndexQ_deqReq_rl$EN = 1'd1 ;
  // register cache_cRqRetryIndexQ_empty
  assign cache_cRqRetryIndexQ_empty$D_IN =
	     cache_cRqRetryIndexQ_clearReq_dummy2_1$Q_OUT &&
	     cache_cRqRetryIndexQ_clearReq_rl ||
	     IF_cache_cRqRetryIndexQ_deqReq_dummy2_2_read___ETC___d854 &&
	     NOT_cache_cRqRetryIndexQ_enqReq_dummy2_2_read__ETC___d876 ;
  assign cache_cRqRetryIndexQ_empty$EN = 1'd1 ;
  // register cache_cRqRetryIndexQ_enqP
  assign cache_cRqRetryIndexQ_enqP$D_IN =
	     (cache_cRqRetryIndexQ_clearReq_dummy2_1$Q_OUT &&
	      cache_cRqRetryIndexQ_clearReq_rl) ?
	       4'd0 :
	       v__h232953 ;
  assign cache_cRqRetryIndexQ_enqP$EN = 1'd1 ;
  // register cache_cRqRetryIndexQ_enqReq_rl
  assign cache_cRqRetryIndexQ_enqReq_rl$D_IN = 5'd10 ;
  assign cache_cRqRetryIndexQ_enqReq_rl$EN = 1'd1 ;
  // register cache_cRqRetryIndexQ_full
  assign cache_cRqRetryIndexQ_full$D_IN =
	     NOT_cache_cRqRetryIndexQ_clearReq_dummy2_1_rea_ETC___d853 &&
	     IF_cache_cRqRetryIndexQ_deqReq_dummy2_2_read___ETC___d854 &&
	     cache_cRqRetryIndexQ_enqReq_dummy2_2_read__28__ETC___d864 ;
  assign cache_cRqRetryIndexQ_full$EN = 1'd1 ;
  // register cache_doLdAfterReplace
  assign cache_doLdAfterReplace$D_IN = !cache_doLdAfterReplace ;
  assign cache_doLdAfterReplace$EN =
	     WILL_FIRE_RL_cache_sendToM && cache_toMInfoQ$D_OUT[1:0] == 2'd2 ;
  // register cache_priorNewCRqSrc
  assign cache_priorNewCRqSrc$D_IN = !cache_priorNewCRqSrc ;
  assign cache_priorNewCRqSrc$EN =
	     WILL_FIRE_RL_cache_cRqTransfer_new_dma ||
	     WILL_FIRE_RL_cache_cRqTransfer_new_child ;
  // register cache_rqFromCQ_clearReq_rl
  assign cache_rqFromCQ_clearReq_rl$D_IN = 1'd0 ;
  assign cache_rqFromCQ_clearReq_rl$EN = 1'd1 ;
  // register cache_rqFromCQ_data_0
  assign cache_rqFromCQ_data_0$D_IN =
	     EN_to_child_rqFromC_enq ?
	       cache_rqFromCQ_enqReq_lat_0$wget[73:0] :
	       cache_rqFromCQ_enqReq_rl[73:0] ;
  assign cache_rqFromCQ_data_0$EN =
	     cache_rqFromCQ_enqP == 1'd0 &&
	     NOT_cache_rqFromCQ_clearReq_dummy2_1_read__8_9_ETC___d33 &&
	     cache_rqFromCQ_enqReq_dummy2_2$Q_OUT &&
	     IF_cache_rqFromCQ_enqReq_lat_1_whas_THEN_cache_ETC___d39 ;
  // register cache_rqFromCQ_data_1
  assign cache_rqFromCQ_data_1$D_IN =
	     EN_to_child_rqFromC_enq ?
	       cache_rqFromCQ_enqReq_lat_0$wget[73:0] :
	       cache_rqFromCQ_enqReq_rl[73:0] ;
  assign cache_rqFromCQ_data_1$EN =
	     cache_rqFromCQ_enqP == 1'd1 &&
	     NOT_cache_rqFromCQ_clearReq_dummy2_1_read__8_9_ETC___d33 &&
	     cache_rqFromCQ_enqReq_dummy2_2$Q_OUT &&
	     IF_cache_rqFromCQ_enqReq_lat_1_whas_THEN_cache_ETC___d39 ;
  // register cache_rqFromCQ_deqP
  assign cache_rqFromCQ_deqP$D_IN =
	     NOT_cache_rqFromCQ_clearReq_dummy2_1_read__8_9_ETC___d33 &&
	     _theResult_____2__h7215 ;
  assign cache_rqFromCQ_deqP$EN = 1'd1 ;
  // register cache_rqFromCQ_deqReq_rl
  assign cache_rqFromCQ_deqReq_rl$D_IN = 1'd0 ;
  assign cache_rqFromCQ_deqReq_rl$EN = 1'd1 ;
  // register cache_rqFromCQ_empty
  assign cache_rqFromCQ_empty$D_IN =
	     cache_rqFromCQ_clearReq_dummy2_1$Q_OUT &&
	     cache_rqFromCQ_clearReq_rl ||
	     IF_cache_rqFromCQ_deqReq_dummy2_2_read__7_AND__ETC___d55 &&
	     NOT_cache_rqFromCQ_enqReq_dummy2_2_read__4_9_O_ETC___d78 ;
  assign cache_rqFromCQ_empty$EN = 1'd1 ;
  // register cache_rqFromCQ_enqP
  assign cache_rqFromCQ_enqP$D_IN =
	     NOT_cache_rqFromCQ_clearReq_dummy2_1_read__8_9_ETC___d33 &&
	     v__h6037 ;
  assign cache_rqFromCQ_enqP$EN = 1'd1 ;
  // register cache_rqFromCQ_enqReq_rl
  assign cache_rqFromCQ_enqReq_rl$D_IN = 75'h2AAAAAAAAAAAAAAAAAA ;
  assign cache_rqFromCQ_enqReq_rl$EN = 1'd1 ;
  // register cache_rqFromCQ_full
  assign cache_rqFromCQ_full$D_IN =
	     NOT_cache_rqFromCQ_clearReq_dummy2_1_read__8_9_ETC___d33 &&
	     IF_cache_rqFromCQ_deqReq_dummy2_2_read__7_AND__ETC___d55 &&
	     cache_rqFromCQ_enqReq_dummy2_2_read__4_AND_IF__ETC___d65 ;
  assign cache_rqFromCQ_full$EN = 1'd1 ;
  // register cache_rqFromDmaQ_clearReq_rl
  assign cache_rqFromDmaQ_clearReq_rl$D_IN = 1'd0 ;
  assign cache_rqFromDmaQ_clearReq_rl$EN = 1'd1 ;
  // register cache_rqFromDmaQ_data_0
  assign cache_rqFromDmaQ_data_0$D_IN =
	     EN_dma_memReq_enq ?
	       cache_rqFromDmaQ_enqReq_lat_0$wget[655:0] :
	       cache_rqFromDmaQ_enqReq_rl[655:0] ;
  assign cache_rqFromDmaQ_data_0$EN =
	     cache_rqFromDmaQ_enqP == 1'd0 &&
	     NOT_cache_rqFromDmaQ_clearReq_dummy2_1_read__3_ETC___d339 &&
	     cache_rqFromDmaQ_enqReq_dummy2_2$Q_OUT &&
	     IF_cache_rqFromDmaQ_enqReq_lat_1_whas__09_THEN_ETC___d345 ;
  // register cache_rqFromDmaQ_data_1
  assign cache_rqFromDmaQ_data_1$D_IN =
	     EN_dma_memReq_enq ?
	       cache_rqFromDmaQ_enqReq_lat_0$wget[655:0] :
	       cache_rqFromDmaQ_enqReq_rl[655:0] ;
  assign cache_rqFromDmaQ_data_1$EN =
	     cache_rqFromDmaQ_enqP == 1'd1 &&
	     NOT_cache_rqFromDmaQ_clearReq_dummy2_1_read__3_ETC___d339 &&
	     cache_rqFromDmaQ_enqReq_dummy2_2$Q_OUT &&
	     IF_cache_rqFromDmaQ_enqReq_lat_1_whas__09_THEN_ETC___d345 ;
  // register cache_rqFromDmaQ_deqP
  assign cache_rqFromDmaQ_deqP$D_IN =
	     NOT_cache_rqFromDmaQ_clearReq_dummy2_1_read__3_ETC___d339 &&
	     _theResult_____2__h119142 ;
  assign cache_rqFromDmaQ_deqP$EN = 1'd1 ;
  // register cache_rqFromDmaQ_deqReq_rl
  assign cache_rqFromDmaQ_deqReq_rl$D_IN = 1'd0 ;
  assign cache_rqFromDmaQ_deqReq_rl$EN = 1'd1 ;
  // register cache_rqFromDmaQ_empty
  assign cache_rqFromDmaQ_empty$D_IN =
	     cache_rqFromDmaQ_clearReq_dummy2_1$Q_OUT &&
	     cache_rqFromDmaQ_clearReq_rl ||
	     IF_cache_rqFromDmaQ_deqReq_dummy2_2_read__53_A_ETC___d361 &&
	     NOT_cache_rqFromDmaQ_enqReq_dummy2_2_read__40__ETC___d384 ;
  assign cache_rqFromDmaQ_empty$EN = 1'd1 ;
  // register cache_rqFromDmaQ_enqP
  assign cache_rqFromDmaQ_enqP$D_IN =
	     NOT_cache_rqFromDmaQ_clearReq_dummy2_1_read__3_ETC___d339 &&
	     v__h72082 ;
  assign cache_rqFromDmaQ_enqP$EN = 1'd1 ;
  // register cache_rqFromDmaQ_enqReq_rl
  assign cache_rqFromDmaQ_enqReq_rl$D_IN =
	     657'h0AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA ;
  assign cache_rqFromDmaQ_enqReq_rl$EN = 1'd1 ;
  // register cache_rqFromDmaQ_full
  assign cache_rqFromDmaQ_full$D_IN =
	     NOT_cache_rqFromDmaQ_clearReq_dummy2_1_read__3_ETC___d339 &&
	     IF_cache_rqFromDmaQ_deqReq_dummy2_2_read__53_A_ETC___d361 &&
	     cache_rqFromDmaQ_enqReq_dummy2_2_read__40_AND__ETC___d371 ;
  assign cache_rqFromDmaQ_full$EN = 1'd1 ;
  // register cache_rsFromCQ_clearReq_rl
  assign cache_rsFromCQ_clearReq_rl$D_IN = 1'd0 ;
  assign cache_rsFromCQ_clearReq_rl$EN = 1'd1 ;
  // register cache_rsFromCQ_data_0
  assign cache_rsFromCQ_data_0$D_IN =
	     EN_to_child_rsFromC_enq ?
	       cache_rsFromCQ_enqReq_lat_0$wget[580:0] :
	       cache_rsFromCQ_enqReq_rl[580:0] ;
  assign cache_rsFromCQ_data_0$EN =
	     cache_rsFromCQ_enqP == 1'd0 &&
	     NOT_cache_rsFromCQ_clearReq_dummy2_1_read__20__ETC___d125 &&
	     cache_rsFromCQ_enqReq_dummy2_2$Q_OUT &&
	     IF_cache_rsFromCQ_enqReq_lat_1_whas__5_THEN_ca_ETC___d131 ;
  // register cache_rsFromCQ_data_1
  assign cache_rsFromCQ_data_1$D_IN =
	     EN_to_child_rsFromC_enq ?
	       cache_rsFromCQ_enqReq_lat_0$wget[580:0] :
	       cache_rsFromCQ_enqReq_rl[580:0] ;
  assign cache_rsFromCQ_data_1$EN =
	     cache_rsFromCQ_enqP == 1'd1 &&
	     NOT_cache_rsFromCQ_clearReq_dummy2_1_read__20__ETC___d125 &&
	     cache_rsFromCQ_enqReq_dummy2_2$Q_OUT &&
	     IF_cache_rsFromCQ_enqReq_lat_1_whas__5_THEN_ca_ETC___d131 ;
  // register cache_rsFromCQ_deqP
  assign cache_rsFromCQ_deqP$D_IN =
	     NOT_cache_rsFromCQ_clearReq_dummy2_1_read__20__ETC___d125 &&
	     _theResult_____2__h22297 ;
  assign cache_rsFromCQ_deqP$EN = 1'd1 ;
  // register cache_rsFromCQ_deqReq_rl
  assign cache_rsFromCQ_deqReq_rl$D_IN = 1'd0 ;
  assign cache_rsFromCQ_deqReq_rl$EN = 1'd1 ;
  // register cache_rsFromCQ_empty
  assign cache_rsFromCQ_empty$D_IN =
	     cache_rsFromCQ_clearReq_dummy2_1$Q_OUT &&
	     cache_rsFromCQ_clearReq_rl ||
	     IF_cache_rsFromCQ_deqReq_dummy2_2_read__39_AND_ETC___d147 &&
	     NOT_cache_rsFromCQ_enqReq_dummy2_2_read__26_61_ETC___d170 ;
  assign cache_rsFromCQ_empty$EN = 1'd1 ;
  // register cache_rsFromCQ_enqP
  assign cache_rsFromCQ_enqP$D_IN =
	     NOT_cache_rsFromCQ_clearReq_dummy2_1_read__20__ETC___d125 &&
	     v__h16641 ;
  assign cache_rsFromCQ_enqP$EN = 1'd1 ;
  // register cache_rsFromCQ_enqReq_rl
  assign cache_rsFromCQ_enqReq_rl$D_IN =
	     582'h0AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA ;
  assign cache_rsFromCQ_enqReq_rl$EN = 1'd1 ;
  // register cache_rsFromCQ_full
  assign cache_rsFromCQ_full$D_IN =
	     NOT_cache_rsFromCQ_clearReq_dummy2_1_read__20__ETC___d125 &&
	     IF_cache_rsFromCQ_deqReq_dummy2_2_read__39_AND_ETC___d147 &&
	     cache_rsFromCQ_enqReq_dummy2_2_read__26_AND_IF_ETC___d157 ;
  assign cache_rsFromCQ_full$EN = 1'd1 ;
  // register cache_rsFromMQ_clearReq_rl
  assign cache_rsFromMQ_clearReq_rl$D_IN = 1'd0 ;
  assign cache_rsFromMQ_clearReq_rl$EN = 1'd1 ;
  // register cache_rsFromMQ_data_0
  assign cache_rsFromMQ_data_0$D_IN =
	     EN_to_mem_rsFromM_enq ?
	       cache_rsFromMQ_enqReq_lat_0$wget[516:0] :
	       cache_rsFromMQ_enqReq_rl[516:0] ;
  assign cache_rsFromMQ_data_0$EN =
	     cache_rsFromMQ_enqP == 1'd0 &&
	     NOT_cache_rsFromMQ_clearReq_dummy2_1_read__35__ETC___d740 &&
	     cache_rsFromMQ_enqReq_dummy2_2$Q_OUT &&
	     IF_cache_rsFromMQ_enqReq_lat_1_whas__10_THEN_c_ETC___d746 ;
  // register cache_rsFromMQ_data_1
  assign cache_rsFromMQ_data_1$D_IN =
	     EN_to_mem_rsFromM_enq ?
	       cache_rsFromMQ_enqReq_lat_0$wget[516:0] :
	       cache_rsFromMQ_enqReq_rl[516:0] ;
  assign cache_rsFromMQ_data_1$EN =
	     cache_rsFromMQ_enqP == 1'd1 &&
	     NOT_cache_rsFromMQ_clearReq_dummy2_1_read__35__ETC___d740 &&
	     cache_rsFromMQ_enqReq_dummy2_2$Q_OUT &&
	     IF_cache_rsFromMQ_enqReq_lat_1_whas__10_THEN_c_ETC___d746 ;
  // register cache_rsFromMQ_deqP
  assign cache_rsFromMQ_deqP$D_IN =
	     NOT_cache_rsFromMQ_clearReq_dummy2_1_read__35__ETC___d740 &&
	     _theResult_____2__h225016 ;
  assign cache_rsFromMQ_deqP$EN = 1'd1 ;
  // register cache_rsFromMQ_deqReq_rl
  assign cache_rsFromMQ_deqReq_rl$D_IN = 1'd0 ;
  assign cache_rsFromMQ_deqReq_rl$EN = 1'd1 ;
  // register cache_rsFromMQ_empty
  assign cache_rsFromMQ_empty$D_IN =
	     cache_rsFromMQ_clearReq_dummy2_1$Q_OUT &&
	     cache_rsFromMQ_clearReq_rl ||
	     IF_cache_rsFromMQ_deqReq_dummy2_2_read__54_AND_ETC___d762 &&
	     NOT_cache_rsFromMQ_enqReq_dummy2_2_read__41_76_ETC___d785 ;
  assign cache_rsFromMQ_empty$EN = 1'd1 ;
  // register cache_rsFromMQ_enqP
  assign cache_rsFromMQ_enqP$D_IN =
	     NOT_cache_rsFromMQ_clearReq_dummy2_1_read__35__ETC___d740 &&
	     v__h218716 ;
  assign cache_rsFromMQ_enqP$EN = 1'd1 ;
  // register cache_rsFromMQ_enqReq_rl
  assign cache_rsFromMQ_enqReq_rl$D_IN =
	     518'h0AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA ;
  assign cache_rsFromMQ_enqReq_rl$EN = 1'd1 ;
  // register cache_rsFromMQ_full
  assign cache_rsFromMQ_full$D_IN =
	     NOT_cache_rsFromMQ_clearReq_dummy2_1_read__35__ETC___d740 &&
	     IF_cache_rsFromMQ_deqReq_dummy2_2_read__54_AND_ETC___d762 &&
	     cache_rsFromMQ_enqReq_dummy2_2_read__41_AND_IF_ETC___d772 ;
  assign cache_rsFromMQ_full$EN = 1'd1 ;
  // register cache_rsLdToDmaQ_clearReq_rl
  assign cache_rsLdToDmaQ_clearReq_rl$D_IN = 1'd0 ;
  assign cache_rsLdToDmaQ_clearReq_rl$EN = 1'd1 ;
  // register cache_rsLdToDmaQ_data_0
  assign cache_rsLdToDmaQ_data_0$D_IN =
	     CAN_FIRE_RL_cache_sendRsLdToDma ?
	       cache_rsLdToDmaQ_enqReq_lat_0$wget[527:0] :
	       cache_rsLdToDmaQ_enqReq_rl[527:0] ;
  assign cache_rsLdToDmaQ_data_0$EN =
	     cache_rsLdToDmaQ_enqP == 1'd0 &&
	     NOT_cache_rsLdToDmaQ_clearReq_dummy2_1_read__2_ETC___d430 &&
	     cache_rsLdToDmaQ_enqReq_dummy2_2$Q_OUT &&
	     IF_cache_rsLdToDmaQ_enqReq_lat_1_whas__00_THEN_ETC___d436 ;
  // register cache_rsLdToDmaQ_data_1
  assign cache_rsLdToDmaQ_data_1$D_IN =
	     CAN_FIRE_RL_cache_sendRsLdToDma ?
	       cache_rsLdToDmaQ_enqReq_lat_0$wget[527:0] :
	       cache_rsLdToDmaQ_enqReq_rl[527:0] ;
  assign cache_rsLdToDmaQ_data_1$EN =
	     cache_rsLdToDmaQ_enqP == 1'd1 &&
	     NOT_cache_rsLdToDmaQ_clearReq_dummy2_1_read__2_ETC___d430 &&
	     cache_rsLdToDmaQ_enqReq_dummy2_2$Q_OUT &&
	     IF_cache_rsLdToDmaQ_enqReq_lat_1_whas__00_THEN_ETC___d436 ;
  // register cache_rsLdToDmaQ_deqP
  assign cache_rsLdToDmaQ_deqP$D_IN =
	     NOT_cache_rsLdToDmaQ_clearReq_dummy2_1_read__2_ETC___d430 &&
	     _theResult_____2__h135235 ;
  assign cache_rsLdToDmaQ_deqP$EN = 1'd1 ;
  // register cache_rsLdToDmaQ_deqReq_rl
  assign cache_rsLdToDmaQ_deqReq_rl$D_IN = 1'd0 ;
  assign cache_rsLdToDmaQ_deqReq_rl$EN = 1'd1 ;
  // register cache_rsLdToDmaQ_empty
  assign cache_rsLdToDmaQ_empty$D_IN =
	     cache_rsLdToDmaQ_clearReq_dummy2_1$Q_OUT &&
	     cache_rsLdToDmaQ_clearReq_rl ||
	     IF_cache_rsLdToDmaQ_deqReq_dummy2_2_read__44_A_ETC___d452 &&
	     NOT_cache_rsLdToDmaQ_enqReq_dummy2_2_read__31__ETC___d475 ;
  assign cache_rsLdToDmaQ_empty$EN = 1'd1 ;
  // register cache_rsLdToDmaQ_enqP
  assign cache_rsLdToDmaQ_enqP$D_IN =
	     NOT_cache_rsLdToDmaQ_clearReq_dummy2_1_read__2_ETC___d430 &&
	     v__h129259 ;
  assign cache_rsLdToDmaQ_enqP$EN = 1'd1 ;
  // register cache_rsLdToDmaQ_enqReq_rl
  assign cache_rsLdToDmaQ_enqReq_rl$D_IN =
	     529'h0AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA ;
  assign cache_rsLdToDmaQ_enqReq_rl$EN = 1'd1 ;
  // register cache_rsLdToDmaQ_full
  assign cache_rsLdToDmaQ_full$D_IN =
	     NOT_cache_rsLdToDmaQ_clearReq_dummy2_1_read__2_ETC___d430 &&
	     IF_cache_rsLdToDmaQ_deqReq_dummy2_2_read__44_A_ETC___d452 &&
	     cache_rsLdToDmaQ_enqReq_dummy2_2_read__31_AND__ETC___d462 ;
  assign cache_rsLdToDmaQ_full$EN = 1'd1 ;
  // register cache_rsStToDmaQ_clearReq_rl
  assign cache_rsStToDmaQ_clearReq_rl$D_IN = 1'd0 ;
  assign cache_rsStToDmaQ_clearReq_rl$EN = 1'd1 ;
  // register cache_rsStToDmaQ_data_0
  assign cache_rsStToDmaQ_data_0$D_IN =
	     WILL_FIRE_RL_cache_sendRsStToDma ?
	       cache_rsStToDmaQ_enqReq_lat_0$wget[15:0] :
	       cache_rsStToDmaQ_enqReq_rl[15:0] ;
  assign cache_rsStToDmaQ_data_0$EN =
	     cache_rsStToDmaQ_enqP == 1'd0 &&
	     NOT_cache_rsStToDmaQ_clearReq_dummy2_1_read__1_ETC___d521 &&
	     cache_rsStToDmaQ_enqReq_dummy2_2$Q_OUT &&
	     IF_cache_rsStToDmaQ_enqReq_lat_1_whas__91_THEN_ETC___d527 ;
  // register cache_rsStToDmaQ_data_1
  assign cache_rsStToDmaQ_data_1$D_IN =
	     WILL_FIRE_RL_cache_sendRsStToDma ?
	       cache_rsStToDmaQ_enqReq_lat_0$wget[15:0] :
	       cache_rsStToDmaQ_enqReq_rl[15:0] ;
  assign cache_rsStToDmaQ_data_1$EN =
	     cache_rsStToDmaQ_enqP == 1'd1 &&
	     NOT_cache_rsStToDmaQ_clearReq_dummy2_1_read__1_ETC___d521 &&
	     cache_rsStToDmaQ_enqReq_dummy2_2$Q_OUT &&
	     IF_cache_rsStToDmaQ_enqReq_lat_1_whas__91_THEN_ETC___d527 ;
  // register cache_rsStToDmaQ_deqP
  assign cache_rsStToDmaQ_deqP$D_IN =
	     NOT_cache_rsStToDmaQ_clearReq_dummy2_1_read__1_ETC___d521 &&
	     _theResult_____2__h142737 ;
  assign cache_rsStToDmaQ_deqP$EN = 1'd1 ;
  // register cache_rsStToDmaQ_deqReq_rl
  assign cache_rsStToDmaQ_deqReq_rl$D_IN = 1'd0 ;
  assign cache_rsStToDmaQ_deqReq_rl$EN = 1'd1 ;
  // register cache_rsStToDmaQ_empty
  assign cache_rsStToDmaQ_empty$D_IN =
	     cache_rsStToDmaQ_clearReq_dummy2_1$Q_OUT &&
	     cache_rsStToDmaQ_clearReq_rl ||
	     IF_cache_rsStToDmaQ_deqReq_dummy2_2_read__35_A_ETC___d543 &&
	     NOT_cache_rsStToDmaQ_enqReq_dummy2_2_read__22__ETC___d566 ;
  assign cache_rsStToDmaQ_empty$EN = 1'd1 ;
  // register cache_rsStToDmaQ_enqP
  assign cache_rsStToDmaQ_enqP$D_IN =
	     NOT_cache_rsStToDmaQ_clearReq_dummy2_1_read__1_ETC___d521 &&
	     v__h142239 ;
  assign cache_rsStToDmaQ_enqP$EN = 1'd1 ;
  // register cache_rsStToDmaQ_enqReq_rl
  assign cache_rsStToDmaQ_enqReq_rl$D_IN = 17'd43690 ;
  assign cache_rsStToDmaQ_enqReq_rl$EN = 1'd1 ;
  // register cache_rsStToDmaQ_full
  assign cache_rsStToDmaQ_full$D_IN =
	     NOT_cache_rsStToDmaQ_clearReq_dummy2_1_read__1_ETC___d521 &&
	     IF_cache_rsStToDmaQ_deqReq_dummy2_2_read__35_A_ETC___d543 &&
	     cache_rsStToDmaQ_enqReq_dummy2_2_read__22_AND__ETC___d553 ;
  assign cache_rsStToDmaQ_full$EN = 1'd1 ;
  // register cache_rsToCIndexQ_clearReq_rl
  assign cache_rsToCIndexQ_clearReq_rl$D_IN = 1'd0 ;
  assign cache_rsToCIndexQ_clearReq_rl$EN = 1'd1 ;
  // register cache_rsToCIndexQ_data_0
  assign cache_rsToCIndexQ_data_0$D_IN =
	     cache_rsToCIndexQ_enqReq_lat_0$whas ?
	       cache_rsToCIndexQ_enqReq_lat_0$wget[5:0] :
	       cache_rsToCIndexQ_enqReq_rl[5:0] ;
  assign cache_rsToCIndexQ_data_0$EN =
	     cache_rsToCIndexQ_enqP == 4'd0 &&
	     NOT_cache_rsToCIndexQ_clearReq_dummy2_1_read___ETC___d976 &&
	     cache_rsToCIndexQ_enqReq_dummy2_2$Q_OUT &&
	     IF_cache_rsToCIndexQ_enqReq_lat_1_whas__24_THE_ETC___d956 ;
  // register cache_rsToCIndexQ_data_1
  assign cache_rsToCIndexQ_data_1$D_IN = cache_rsToCIndexQ_data_0$D_IN ;
  assign cache_rsToCIndexQ_data_1$EN =
	     cache_rsToCIndexQ_enqP == 4'd1 &&
	     NOT_cache_rsToCIndexQ_clearReq_dummy2_1_read___ETC___d976 &&
	     cache_rsToCIndexQ_enqReq_dummy2_2$Q_OUT &&
	     IF_cache_rsToCIndexQ_enqReq_lat_1_whas__24_THE_ETC___d956 ;
  // register cache_rsToCIndexQ_data_10
  assign cache_rsToCIndexQ_data_10$D_IN = cache_rsToCIndexQ_data_0$D_IN ;
  assign cache_rsToCIndexQ_data_10$EN =
	     cache_rsToCIndexQ_enqP == 4'd10 &&
	     NOT_cache_rsToCIndexQ_clearReq_dummy2_1_read___ETC___d976 &&
	     cache_rsToCIndexQ_enqReq_dummy2_2$Q_OUT &&
	     IF_cache_rsToCIndexQ_enqReq_lat_1_whas__24_THE_ETC___d956 ;
  // register cache_rsToCIndexQ_data_11
  assign cache_rsToCIndexQ_data_11$D_IN = cache_rsToCIndexQ_data_0$D_IN ;
  assign cache_rsToCIndexQ_data_11$EN =
	     cache_rsToCIndexQ_enqP == 4'd11 &&
	     NOT_cache_rsToCIndexQ_clearReq_dummy2_1_read___ETC___d976 &&
	     cache_rsToCIndexQ_enqReq_dummy2_2$Q_OUT &&
	     IF_cache_rsToCIndexQ_enqReq_lat_1_whas__24_THE_ETC___d956 ;
  // register cache_rsToCIndexQ_data_12
  assign cache_rsToCIndexQ_data_12$D_IN = cache_rsToCIndexQ_data_0$D_IN ;
  assign cache_rsToCIndexQ_data_12$EN =
	     cache_rsToCIndexQ_enqP == 4'd12 &&
	     NOT_cache_rsToCIndexQ_clearReq_dummy2_1_read___ETC___d976 &&
	     cache_rsToCIndexQ_enqReq_dummy2_2$Q_OUT &&
	     IF_cache_rsToCIndexQ_enqReq_lat_1_whas__24_THE_ETC___d956 ;
  // register cache_rsToCIndexQ_data_13
  assign cache_rsToCIndexQ_data_13$D_IN = cache_rsToCIndexQ_data_0$D_IN ;
  assign cache_rsToCIndexQ_data_13$EN =
	     cache_rsToCIndexQ_enqP == 4'd13 &&
	     NOT_cache_rsToCIndexQ_clearReq_dummy2_1_read___ETC___d976 &&
	     cache_rsToCIndexQ_enqReq_dummy2_2$Q_OUT &&
	     IF_cache_rsToCIndexQ_enqReq_lat_1_whas__24_THE_ETC___d956 ;
  // register cache_rsToCIndexQ_data_14
  assign cache_rsToCIndexQ_data_14$D_IN = cache_rsToCIndexQ_data_0$D_IN ;
  assign cache_rsToCIndexQ_data_14$EN =
	     cache_rsToCIndexQ_enqP == 4'd14 &&
	     NOT_cache_rsToCIndexQ_clearReq_dummy2_1_read___ETC___d976 &&
	     cache_rsToCIndexQ_enqReq_dummy2_2$Q_OUT &&
	     IF_cache_rsToCIndexQ_enqReq_lat_1_whas__24_THE_ETC___d956 ;
  // register cache_rsToCIndexQ_data_15
  assign cache_rsToCIndexQ_data_15$D_IN = cache_rsToCIndexQ_data_0$D_IN ;
  assign cache_rsToCIndexQ_data_15$EN =
	     cache_rsToCIndexQ_enqP == 4'd15 &&
	     NOT_cache_rsToCIndexQ_clearReq_dummy2_1_read___ETC___d976 &&
	     cache_rsToCIndexQ_enqReq_dummy2_2$Q_OUT &&
	     IF_cache_rsToCIndexQ_enqReq_lat_1_whas__24_THE_ETC___d956 ;
  // register cache_rsToCIndexQ_data_2
  assign cache_rsToCIndexQ_data_2$D_IN = cache_rsToCIndexQ_data_0$D_IN ;
  assign cache_rsToCIndexQ_data_2$EN =
	     cache_rsToCIndexQ_enqP == 4'd2 &&
	     NOT_cache_rsToCIndexQ_clearReq_dummy2_1_read___ETC___d976 &&
	     cache_rsToCIndexQ_enqReq_dummy2_2$Q_OUT &&
	     IF_cache_rsToCIndexQ_enqReq_lat_1_whas__24_THE_ETC___d956 ;
  // register cache_rsToCIndexQ_data_3
  assign cache_rsToCIndexQ_data_3$D_IN = cache_rsToCIndexQ_data_0$D_IN ;
  assign cache_rsToCIndexQ_data_3$EN =
	     cache_rsToCIndexQ_enqP == 4'd3 &&
	     NOT_cache_rsToCIndexQ_clearReq_dummy2_1_read___ETC___d976 &&
	     cache_rsToCIndexQ_enqReq_dummy2_2$Q_OUT &&
	     IF_cache_rsToCIndexQ_enqReq_lat_1_whas__24_THE_ETC___d956 ;
  // register cache_rsToCIndexQ_data_4
  assign cache_rsToCIndexQ_data_4$D_IN = cache_rsToCIndexQ_data_0$D_IN ;
  assign cache_rsToCIndexQ_data_4$EN =
	     cache_rsToCIndexQ_enqP == 4'd4 &&
	     NOT_cache_rsToCIndexQ_clearReq_dummy2_1_read___ETC___d976 &&
	     cache_rsToCIndexQ_enqReq_dummy2_2$Q_OUT &&
	     IF_cache_rsToCIndexQ_enqReq_lat_1_whas__24_THE_ETC___d956 ;
  // register cache_rsToCIndexQ_data_5
  assign cache_rsToCIndexQ_data_5$D_IN = cache_rsToCIndexQ_data_0$D_IN ;
  assign cache_rsToCIndexQ_data_5$EN =
	     cache_rsToCIndexQ_enqP == 4'd5 &&
	     NOT_cache_rsToCIndexQ_clearReq_dummy2_1_read___ETC___d976 &&
	     cache_rsToCIndexQ_enqReq_dummy2_2$Q_OUT &&
	     IF_cache_rsToCIndexQ_enqReq_lat_1_whas__24_THE_ETC___d956 ;
  // register cache_rsToCIndexQ_data_6
  assign cache_rsToCIndexQ_data_6$D_IN = cache_rsToCIndexQ_data_0$D_IN ;
  assign cache_rsToCIndexQ_data_6$EN =
	     cache_rsToCIndexQ_enqP == 4'd6 &&
	     NOT_cache_rsToCIndexQ_clearReq_dummy2_1_read___ETC___d976 &&
	     cache_rsToCIndexQ_enqReq_dummy2_2$Q_OUT &&
	     IF_cache_rsToCIndexQ_enqReq_lat_1_whas__24_THE_ETC___d956 ;
  // register cache_rsToCIndexQ_data_7
  assign cache_rsToCIndexQ_data_7$D_IN = cache_rsToCIndexQ_data_0$D_IN ;
  assign cache_rsToCIndexQ_data_7$EN =
	     cache_rsToCIndexQ_enqP == 4'd7 &&
	     NOT_cache_rsToCIndexQ_clearReq_dummy2_1_read___ETC___d976 &&
	     cache_rsToCIndexQ_enqReq_dummy2_2$Q_OUT &&
	     IF_cache_rsToCIndexQ_enqReq_lat_1_whas__24_THE_ETC___d956 ;
  // register cache_rsToCIndexQ_data_8
  assign cache_rsToCIndexQ_data_8$D_IN = cache_rsToCIndexQ_data_0$D_IN ;
  assign cache_rsToCIndexQ_data_8$EN =
	     cache_rsToCIndexQ_enqP == 4'd8 &&
	     NOT_cache_rsToCIndexQ_clearReq_dummy2_1_read___ETC___d976 &&
	     cache_rsToCIndexQ_enqReq_dummy2_2$Q_OUT &&
	     IF_cache_rsToCIndexQ_enqReq_lat_1_whas__24_THE_ETC___d956 ;
  // register cache_rsToCIndexQ_data_9
  assign cache_rsToCIndexQ_data_9$D_IN = cache_rsToCIndexQ_data_0$D_IN ;
  assign cache_rsToCIndexQ_data_9$EN =
	     cache_rsToCIndexQ_enqP == 4'd9 &&
	     NOT_cache_rsToCIndexQ_clearReq_dummy2_1_read___ETC___d976 &&
	     cache_rsToCIndexQ_enqReq_dummy2_2$Q_OUT &&
	     IF_cache_rsToCIndexQ_enqReq_lat_1_whas__24_THE_ETC___d956 ;
  // register cache_rsToCIndexQ_deqP
  assign cache_rsToCIndexQ_deqP$D_IN =
	     (cache_rsToCIndexQ_clearReq_dummy2_1$Q_OUT &&
	      cache_rsToCIndexQ_clearReq_rl) ?
	       4'd0 :
	       _theResult_____2__h245988 ;
  assign cache_rsToCIndexQ_deqP$EN = 1'd1 ;
  // register cache_rsToCIndexQ_deqReq_rl
  assign cache_rsToCIndexQ_deqReq_rl$D_IN = 1'd0 ;
  assign cache_rsToCIndexQ_deqReq_rl$EN = 1'd1 ;
  // register cache_rsToCIndexQ_empty
  assign cache_rsToCIndexQ_empty$D_IN =
	     cache_rsToCIndexQ_clearReq_dummy2_1$Q_OUT &&
	     cache_rsToCIndexQ_clearReq_rl ||
	     IF_cache_rsToCIndexQ_deqReq_dummy2_2_read__64__ETC___d977 &&
	     NOT_cache_rsToCIndexQ_enqReq_dummy2_2_read__51_ETC___d999 ;
  assign cache_rsToCIndexQ_empty$EN = 1'd1 ;
  // register cache_rsToCIndexQ_enqP
  assign cache_rsToCIndexQ_enqP$D_IN =
	     (cache_rsToCIndexQ_clearReq_dummy2_1$Q_OUT &&
	      cache_rsToCIndexQ_clearReq_rl) ?
	       4'd0 :
	       v__h242396 ;
  assign cache_rsToCIndexQ_enqP$EN = 1'd1 ;
  // register cache_rsToCIndexQ_enqReq_rl
  assign cache_rsToCIndexQ_enqReq_rl$D_IN = 7'd42 ;
  assign cache_rsToCIndexQ_enqReq_rl$EN = 1'd1 ;
  // register cache_rsToCIndexQ_full
  assign cache_rsToCIndexQ_full$D_IN =
	     NOT_cache_rsToCIndexQ_clearReq_dummy2_1_read___ETC___d976 &&
	     IF_cache_rsToCIndexQ_deqReq_dummy2_2_read__64__ETC___d977 &&
	     cache_rsToCIndexQ_enqReq_dummy2_2_read__51_AND_ETC___d987 ;
  assign cache_rsToCIndexQ_full$EN = 1'd1 ;
  // register cache_toCQ_clearReq_rl
  assign cache_toCQ_clearReq_rl$D_IN = 1'd0 ;
  assign cache_toCQ_clearReq_rl$EN = 1'd1 ;
  // register cache_toCQ_data_0
  assign cache_toCQ_data_0$D_IN =
	     { cache_toCQ_enqReq_lat_0$whas ?
		 cache_toCQ_enqReq_lat_0$wget[584] :
		 cache_toCQ_enqReq_rl[584],
	       IF_cache_toCQ_enqReq_dummy2_2_read__53_AND_IF__ETC___d302 } ;
  assign cache_toCQ_data_0$EN =
	     cache_toCQ_enqP == 1'd0 &&
	     NOT_cache_toCQ_clearReq_dummy2_1_read__47_48_O_ETC___d252 &&
	     cache_toCQ_enqReq_dummy2_2$Q_OUT &&
	     IF_cache_toCQ_enqReq_lat_1_whas__87_THEN_cache_ETC___d196 ;
  // register cache_toCQ_data_1
  assign cache_toCQ_data_1$D_IN = cache_toCQ_data_0$D_IN ;
  assign cache_toCQ_data_1$EN =
	     cache_toCQ_enqP == 1'd1 &&
	     NOT_cache_toCQ_clearReq_dummy2_1_read__47_48_O_ETC___d252 &&
	     cache_toCQ_enqReq_dummy2_2$Q_OUT &&
	     IF_cache_toCQ_enqReq_lat_1_whas__87_THEN_cache_ETC___d196 ;
  // register cache_toCQ_deqP
  assign cache_toCQ_deqP$D_IN =
	     NOT_cache_toCQ_clearReq_dummy2_1_read__47_48_O_ETC___d252 &&
	     _theResult_____2__h37990 ;
  assign cache_toCQ_deqP$EN = 1'd1 ;
  // register cache_toCQ_deqReq_rl
  assign cache_toCQ_deqReq_rl$D_IN = 1'd0 ;
  assign cache_toCQ_deqReq_rl$EN = 1'd1 ;
  // register cache_toCQ_empty
  assign cache_toCQ_empty$D_IN =
	     cache_toCQ_clearReq_dummy2_1$Q_OUT && cache_toCQ_clearReq_rl ||
	     IF_cache_toCQ_deqReq_dummy2_2_read__61_AND_IF__ETC___d269 &&
	     NOT_cache_toCQ_enqReq_dummy2_2_read__53_83_OR__ETC___d292 ;
  assign cache_toCQ_empty$EN = 1'd1 ;
  // register cache_toCQ_enqP
  assign cache_toCQ_enqP$D_IN =
	     NOT_cache_toCQ_clearReq_dummy2_1_read__47_48_O_ETC___d252 &&
	     v__h31944 ;
  assign cache_toCQ_enqP$EN = 1'd1 ;
  // register cache_toCQ_enqReq_rl
  assign cache_toCQ_enqReq_rl$D_IN =
	     586'h0AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA ;
  assign cache_toCQ_enqReq_rl$EN = 1'd1 ;
  // register cache_toCQ_full
  assign cache_toCQ_full$D_IN =
	     NOT_cache_toCQ_clearReq_dummy2_1_read__47_48_O_ETC___d252 &&
	     IF_cache_toCQ_deqReq_dummy2_2_read__61_AND_IF__ETC___d269 &&
	     cache_toCQ_enqReq_dummy2_2_read__53_AND_IF_cac_ETC___d279 ;
  assign cache_toCQ_full$EN = 1'd1 ;
  // register cache_toMQ_clearReq_rl
  assign cache_toMQ_clearReq_rl$D_IN = 1'd0 ;
  assign cache_toMQ_clearReq_rl$EN = 1'd1 ;
  // register cache_toMQ_data_0
  assign cache_toMQ_data_0$D_IN =
	     { cache_toMQ_enqReq_lat_0$whas ?
		 cache_toMQ_enqReq_lat_0$wget[640] :
		 cache_toMQ_enqReq_rl[640],
	       IF_cache_toMQ_enqReq_dummy2_2_read__54_AND_IF__ETC___d703 } ;
  assign cache_toMQ_data_0$EN =
	     cache_toMQ_enqP == 1'd0 &&
	     NOT_cache_toMQ_clearReq_dummy2_1_read__48_49_O_ETC___d653 &&
	     cache_toMQ_enqReq_dummy2_2$Q_OUT &&
	     IF_cache_toMQ_enqReq_lat_1_whas__88_THEN_cache_ETC___d597 ;
  // register cache_toMQ_data_1
  assign cache_toMQ_data_1$D_IN = cache_toMQ_data_0$D_IN ;
  assign cache_toMQ_data_1$EN =
	     cache_toMQ_enqP == 1'd1 &&
	     NOT_cache_toMQ_clearReq_dummy2_1_read__48_49_O_ETC___d653 &&
	     cache_toMQ_enqReq_dummy2_2$Q_OUT &&
	     IF_cache_toMQ_enqReq_lat_1_whas__88_THEN_cache_ETC___d597 ;
  // register cache_toMQ_deqP
  assign cache_toMQ_deqP$D_IN =
	     NOT_cache_toMQ_clearReq_dummy2_1_read__48_49_O_ETC___d653 &&
	     _theResult_____2__h208521 ;
  assign cache_toMQ_deqP$EN = 1'd1 ;
  // register cache_toMQ_deqReq_rl
  assign cache_toMQ_deqReq_rl$D_IN = 1'd0 ;
  assign cache_toMQ_deqReq_rl$EN = 1'd1 ;
  // register cache_toMQ_empty
  assign cache_toMQ_empty$D_IN =
	     cache_toMQ_clearReq_dummy2_1$Q_OUT && cache_toMQ_clearReq_rl ||
	     IF_cache_toMQ_deqReq_dummy2_2_read__62_AND_IF__ETC___d670 &&
	     NOT_cache_toMQ_enqReq_dummy2_2_read__54_84_OR__ETC___d693 ;
  assign cache_toMQ_empty$EN = 1'd1 ;
  // register cache_toMQ_enqP
  assign cache_toMQ_enqP$D_IN =
	     NOT_cache_toMQ_clearReq_dummy2_1_read__48_49_O_ETC___d653 &&
	     v__h168573 ;
  assign cache_toMQ_enqP$EN = 1'd1 ;
  // register cache_toMQ_enqReq_rl
  assign cache_toMQ_enqReq_rl$D_IN =
	     642'h055555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555554AAAAAAAAAAAAAAAAA ;
  assign cache_toMQ_enqReq_rl$EN = 1'd1 ;
  // register cache_toMQ_full
  assign cache_toMQ_full$D_IN =
	     NOT_cache_toMQ_clearReq_dummy2_1_read__48_49_O_ETC___d653 &&
	     IF_cache_toMQ_deqReq_dummy2_2_read__62_AND_IF__ETC___d670 &&
	     cache_toMQ_enqReq_dummy2_2_read__54_AND_IF_cac_ETC___d680 ;
  assign cache_toMQ_full$EN = 1'd1 ;
  // register cache_whichCRq
  assign cache_whichCRq$D_IN =
	     (cache_whichCRq == 4'd15) ? 4'd0 : cache_whichCRq + 4'd1 ;
  assign cache_whichCRq$EN = CAN_FIRE_RL_cache_sendRqToC ;
  // register perfReqQ_clearReq_rl
  assign perfReqQ_clearReq_rl$D_IN = 1'd0 ;
  assign perfReqQ_clearReq_rl$EN = 1'd1 ;
  // register perfReqQ_data_0
  assign perfReqQ_data_0$D_IN =
	     EN_perf_req ?
	       perfReqQ_enqReq_lat_0$wget[3:0] :
	       perfReqQ_enqReq_rl[3:0] ;
  assign perfReqQ_data_0$EN =
	     NOT_perfReqQ_clearReq_dummy2_1_read__864_865_O_ETC___d3869 &&
	     perfReqQ_enqReq_dummy2_2$Q_OUT &&
	     IF_perfReqQ_enqReq_lat_1_whas__839_THEN_perfRe_ETC___d3875 ;
  // register perfReqQ_deqReq_rl
  assign perfReqQ_deqReq_rl$D_IN = 1'd0 ;
  assign perfReqQ_deqReq_rl$EN = 1'd1 ;
  // register perfReqQ_empty
  assign perfReqQ_empty$D_IN =
	     perfReqQ_clearReq_dummy2_1$Q_OUT && perfReqQ_clearReq_rl ||
	     NOT_perfReqQ_enqReq_dummy2_2_read__870_890_OR__ETC___d3900 ;
  assign perfReqQ_empty$EN = 1'd1 ;
  // register perfReqQ_enqReq_rl
  assign perfReqQ_enqReq_rl$D_IN = 5'd10 ;
  assign perfReqQ_enqReq_rl$EN = 1'd1 ;
  // register perfReqQ_full
  assign perfReqQ_full$D_IN =
	     NOT_perfReqQ_clearReq_dummy2_1_read__864_865_O_ETC___d3869 &&
	     perfReqQ_enqReq_dummy2_2_read__870_AND_IF_perf_ETC___d3887 ;
  assign perfReqQ_full$EN = 1'd1 ;
  // submodule cache_cRqMshr
  assign cache_cRqMshr$mRsDeq_setData_d =
	     { 1'd1,
	       SEL_ARR_cache_rsFromMQ_data_0_914_BITS_516_TO__ETC___d1966 } ;
  assign cache_cRqMshr$mRsDeq_setData_n =
	     MUX_cache_cRqMshr$transfer_getRq_1__VAL_2 ;
  assign cache_cRqMshr$pipelineResp_getAddrSucc_n = pipeOutCRqIdx__h314276 ;
  assign cache_cRqMshr$pipelineResp_getData_n =
	     WILL_FIRE_RL_cache_pipelineResp_cRq ?
	       cache_pipeline$first[582:579] :
	       cache_pipeline$first[516:513] ;
  assign cache_cRqMshr$pipelineResp_getRepSucc_n = pipeOutCRqIdx__h314276 ;
  assign cache_cRqMshr$pipelineResp_getRq_n = pipeOutCRqIdx__h314276 ;
  assign cache_cRqMshr$pipelineResp_getSlot_n = pipeOutCRqIdx__h314276 ;
  assign cache_cRqMshr$pipelineResp_getState_n = pipeOutCRqIdx__h314276 ;
  assign cache_cRqMshr$pipelineResp_searchEndOfChain_addr =
	     cache_cRqMshr$pipelineResp_getRq[151:88] ;
  assign cache_cRqMshr$pipelineResp_setAddrSucc_n =
	     cache_cRqMshr$pipelineResp_searchEndOfChain[3:0] ;
  assign cache_cRqMshr$pipelineResp_setAddrSucc_succ =
	     { 1'd1, cache_pipeline$first[582:579] } ;
  always@(MUX_cache_cRqMshr$pipelineResp_setData_1__SEL_1 or
	  MUX_cache_cRqMshr$pipelineResp_setData_2__VAL_1 or
	  MUX_cache_cRqMshr$pipelineResp_setData_1__SEL_2 or
	  MUX_cache_cRqMshr$pipelineResp_setData_2__VAL_2 or
	  WILL_FIRE_RL_cache_pipelineResp_mRs or
	  MUX_cache_cRqMshr$pipelineResp_setData_2__VAL_3)
  begin
    case (1'b1) // synopsys parallel_case
      MUX_cache_cRqMshr$pipelineResp_setData_1__SEL_1:
	  cache_cRqMshr$pipelineResp_setData_d =
	      MUX_cache_cRqMshr$pipelineResp_setData_2__VAL_1;
      MUX_cache_cRqMshr$pipelineResp_setData_1__SEL_2:
	  cache_cRqMshr$pipelineResp_setData_d =
	      MUX_cache_cRqMshr$pipelineResp_setData_2__VAL_2;
      WILL_FIRE_RL_cache_pipelineResp_mRs:
	  cache_cRqMshr$pipelineResp_setData_d =
	      MUX_cache_cRqMshr$pipelineResp_setData_2__VAL_3;
      default: cache_cRqMshr$pipelineResp_setData_d =
		   513'h0AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA /* unspecified value */ ;
    endcase
  end
  assign cache_cRqMshr$pipelineResp_setData_n =
	     (MUX_cache_cRqMshr$pipelineResp_setData_1__SEL_2 ||
	      WILL_FIRE_RL_cache_pipelineResp_mRs) ?
	       cache_pipeline$first[516:513] :
	       cache_pipeline$first[582:579] ;
  assign cache_cRqMshr$pipelineResp_setRepSucc_n =
	     cache_pipeline$first[516:513] ;
  assign cache_cRqMshr$pipelineResp_setRepSucc_succ =
	     { 1'd1, cache_pipeline$first[582:579] } ;
  assign cache_cRqMshr$pipelineResp_setStateSlot_n =
	     (MUX_cache_cRqMshr$pipelineResp_setStateSlot_1__SEL_1 ||
	      WILL_FIRE_RL_cache_pipelineResp_mRs) ?
	       cache_pipeline$first[516:513] :
	       cache_pipeline$first[582:579] ;
  always@(MUX_cache_cRqMshr$pipelineResp_setStateSlot_1__SEL_1 or
	  MUX_cache_cRqMshr$pipelineResp_setStateSlot_3__VAL_1 or
	  WILL_FIRE_RL_cache_pipelineResp_cRq or
	  MUX_cache_cRqMshr$pipelineResp_setStateSlot_3__VAL_2 or
	  WILL_FIRE_RL_cache_pipelineResp_mRs)
  begin
    case (1'b1) // synopsys parallel_case
      MUX_cache_cRqMshr$pipelineResp_setStateSlot_1__SEL_1:
	  cache_cRqMshr$pipelineResp_setStateSlot_slot =
	      MUX_cache_cRqMshr$pipelineResp_setStateSlot_3__VAL_1;
      WILL_FIRE_RL_cache_pipelineResp_cRq:
	  cache_cRqMshr$pipelineResp_setStateSlot_slot =
	      MUX_cache_cRqMshr$pipelineResp_setStateSlot_3__VAL_2;
      WILL_FIRE_RL_cache_pipelineResp_mRs:
	  cache_cRqMshr$pipelineResp_setStateSlot_slot =
	      65'h0AAAAAAAAAAAAAAAA /* unspecified value */ ;
      default: cache_cRqMshr$pipelineResp_setStateSlot_slot =
		   65'h0AAAAAAAAAAAAAAAA /* unspecified value */ ;
    endcase
  end
  always@(MUX_cache_cRqMshr$pipelineResp_setStateSlot_1__SEL_1 or
	  MUX_cache_cRqMshr$pipelineResp_setStateSlot_2__VAL_1 or
	  WILL_FIRE_RL_cache_pipelineResp_cRq or
	  MUX_cache_cRqMshr$pipelineResp_setStateSlot_2__VAL_2 or
	  WILL_FIRE_RL_cache_pipelineResp_mRs)
  begin
    case (1'b1) // synopsys parallel_case
      MUX_cache_cRqMshr$pipelineResp_setStateSlot_1__SEL_1:
	  cache_cRqMshr$pipelineResp_setStateSlot_state =
	      MUX_cache_cRqMshr$pipelineResp_setStateSlot_2__VAL_1;
      WILL_FIRE_RL_cache_pipelineResp_cRq:
	  cache_cRqMshr$pipelineResp_setStateSlot_state =
	      MUX_cache_cRqMshr$pipelineResp_setStateSlot_2__VAL_2;
      WILL_FIRE_RL_cache_pipelineResp_mRs:
	  cache_cRqMshr$pipelineResp_setStateSlot_state = 3'd4;
      default: cache_cRqMshr$pipelineResp_setStateSlot_state =
		   3'b010 /* unspecified value */ ;
    endcase
  end
  assign cache_cRqMshr$sendRqToC_getRq_n =
	     cache_cRqMshr$sendRqToC_searchNeedRqChild[3:0] ;
  assign cache_cRqMshr$sendRqToC_getSlot_n =
	     cache_cRqMshr$sendRqToC_searchNeedRqChild[3:0] ;
  assign cache_cRqMshr$sendRqToC_getState_n =
	     cache_cRqMshr$sendRqToC_searchNeedRqChild[3:0] ;
  assign cache_cRqMshr$sendRqToC_searchNeedRqChild_suggestIdx =
	     { 1'd1, cache_whichCRq } ;
  assign cache_cRqMshr$sendRqToC_setSlot_n =
	     cache_cRqMshr$sendRqToC_searchNeedRqChild[3:0] ;
  assign cache_cRqMshr$sendRqToC_setSlot_s =
	     { cache_cRqMshr$sendRqToC_getSlot[64:12],
	       (cache_cRqMshr$sendRqToC_getSlot[3:2] != 2'd1 &&
		cache_cRqMshr$sendRqToC_getSlot[7:6] != 2'd1) ?
		 2'd2 :
		 cache_cRqMshr$sendRqToC_getSlot[11:10],
	       ((cache_cRqMshr$sendRqToC_getSlot[3:2] == 2'd1 ||
		 cache_cRqMshr$sendRqToC_getSlot[7:6] == 2'd1) &&
		cache_cRqMshr$sendRqToC_getSlot[11:10] == 2'd1) ?
		 cache_cRqMshr$sendRqToC_getSlot[9:8] :
		 ((cache_cRqMshr$sendRqToC_getSlot[3:2] != 2'd1 &&
		   cache_cRqMshr$sendRqToC_getSlot[7:6] != 2'd1) ?
		    SEL_ARR_IF_cache_cRqMshr_sendRqToC_getSlot_IF__ETC___d2522 :
		    cache_cRqMshr$sendRqToC_getSlot[9:8]),
	       (cache_cRqMshr$sendRqToC_getSlot[7:6] == 2'd1 &&
		cache_cRqMshr$sendRqToC_getSlot[3:2] != 2'd1) ?
		 2'd2 :
		 cache_cRqMshr$sendRqToC_getSlot[7:6],
	       (cache_cRqMshr$sendRqToC_getSlot[3:2] == 2'd1 &&
		cache_cRqMshr$sendRqToC_getSlot[7:6] == 2'd1) ?
		 cache_cRqMshr$sendRqToC_getSlot[5:4] :
		 ((cache_cRqMshr$sendRqToC_getSlot[7:6] == 2'd1 &&
		   cache_cRqMshr$sendRqToC_getSlot[3:2] != 2'd1) ?
		    SEL_ARR_IF_cache_cRqMshr_sendRqToC_getSlot_IF__ETC___d2522 :
		    cache_cRqMshr$sendRqToC_getSlot[5:4]),
	       (cache_cRqMshr$sendRqToC_getSlot[3:2] == 2'd1) ?
		 2'd2 :
		 cache_cRqMshr$sendRqToC_getSlot[3:2],
	       (cache_cRqMshr$sendRqToC_getSlot[3:2] == 2'd1) ?
		 SEL_ARR_IF_cache_cRqMshr_sendRqToC_getSlot_IF__ETC___d2522 :
		 cache_cRqMshr$sendRqToC_getSlot[1:0] } ;
  assign cache_cRqMshr$sendRsToDmaC_getData_n =
	     WILL_FIRE_RL_cache_sendRsLdToDma ?
	       cache_rsLdToDmaIndexQ$D_OUT :
	       MUX_cache_cRqMshr$sendRsToDmaC_getData_1__VAL_2 ;
  always@(WILL_FIRE_RL_cache_sendRsLdToDma or
	  cache_rsLdToDmaIndexQ$D_OUT or
	  WILL_FIRE_RL_cache_sendRsToC or
	  MUX_cache_cRqMshr$sendRsToDmaC_getData_1__VAL_2 or
	  WILL_FIRE_RL_cache_sendRsStToDma or cache_rsStToDmaIndexQ$D_OUT)
  begin
    case (1'b1) // synopsys parallel_case
      WILL_FIRE_RL_cache_sendRsLdToDma:
	  cache_cRqMshr$sendRsToDmaC_getRq_n = cache_rsLdToDmaIndexQ$D_OUT;
      WILL_FIRE_RL_cache_sendRsToC:
	  cache_cRqMshr$sendRsToDmaC_getRq_n =
	      MUX_cache_cRqMshr$sendRsToDmaC_getData_1__VAL_2;
      WILL_FIRE_RL_cache_sendRsStToDma:
	  cache_cRqMshr$sendRsToDmaC_getRq_n = cache_rsStToDmaIndexQ$D_OUT;
      default: cache_cRqMshr$sendRsToDmaC_getRq_n =
		   4'b1010 /* unspecified value */ ;
    endcase
  end
  always@(WILL_FIRE_RL_cache_sendRsLdToDma or
	  cache_rsLdToDmaIndexQ$D_OUT or
	  WILL_FIRE_RL_cache_sendRsToC or
	  MUX_cache_cRqMshr$sendRsToDmaC_getData_1__VAL_2 or
	  WILL_FIRE_RL_cache_sendRsStToDma or cache_rsStToDmaIndexQ$D_OUT)
  begin
    case (1'b1) // synopsys parallel_case
      WILL_FIRE_RL_cache_sendRsLdToDma:
	  cache_cRqMshr$sendRsToDmaC_releaseEntry_n =
	      cache_rsLdToDmaIndexQ$D_OUT;
      WILL_FIRE_RL_cache_sendRsToC:
	  cache_cRqMshr$sendRsToDmaC_releaseEntry_n =
	      MUX_cache_cRqMshr$sendRsToDmaC_getData_1__VAL_2;
      WILL_FIRE_RL_cache_sendRsStToDma:
	  cache_cRqMshr$sendRsToDmaC_releaseEntry_n =
	      cache_rsStToDmaIndexQ$D_OUT;
      default: cache_cRqMshr$sendRsToDmaC_releaseEntry_n =
		   4'b1010 /* unspecified value */ ;
    endcase
  end
  assign cache_cRqMshr$sendToM_getData_n = cache_toMInfoQ$D_OUT[5:2] ;
  assign cache_cRqMshr$sendToM_getRq_n = cache_toMInfoQ$D_OUT[5:2] ;
  assign cache_cRqMshr$sendToM_getSlot_n = cache_toMInfoQ$D_OUT[5:2] ;
  assign cache_cRqMshr$transfer_getEmptyEntryInit_d =
	     WILL_FIRE_RL_cache_cRqTransfer_new_child ?
	       513'h0AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA :
	       MUX_cache_cRqMshr$transfer_getEmptyEntryInit_2__VAL_2 ;
  assign cache_cRqMshr$transfer_getEmptyEntryInit_r =
	     WILL_FIRE_RL_cache_cRqTransfer_new_child ?
	       MUX_cache_cRqMshr$transfer_getEmptyEntryInit_1__VAL_1 :
	       MUX_cache_cRqMshr$transfer_getEmptyEntryInit_1__VAL_2 ;
  assign cache_cRqMshr$transfer_getRq_n =
	     WILL_FIRE_RL_cache_cRqTransfer_retry ?
	       x__h248737 :
	       MUX_cache_cRqMshr$transfer_getRq_1__VAL_2 ;
  assign cache_cRqMshr$transfer_getSlot_n =
	     MUX_cache_cRqMshr$transfer_getRq_1__VAL_2 ;
  assign cache_cRqMshr$transfer_hasEmptyEntry_r = 152'h0 ;
  assign cache_cRqMshr$EN_transfer_getEmptyEntryInit =
	     WILL_FIRE_RL_cache_cRqTransfer_new_child ||
	     WILL_FIRE_RL_cache_cRqTransfer_new_dma ;
  assign cache_cRqMshr$EN_mRsDeq_setData =
	     CAN_FIRE_RL_cache_mRsDeq_nonRefill ;
  assign cache_cRqMshr$EN_sendRsToDmaC_releaseEntry =
	     WILL_FIRE_RL_cache_sendRsLdToDma ||
	     WILL_FIRE_RL_cache_sendRsToC ||
	     WILL_FIRE_RL_cache_sendRsStToDma ;
  assign cache_cRqMshr$EN_sendRqToC_setSlot = CAN_FIRE_RL_cache_sendRqToC ;
  assign cache_cRqMshr$EN_pipelineResp_setData =
	     MUX_cache_cRqMshr$pipelineResp_setData_1__SEL_1 ||
	     MUX_cache_cRqMshr$pipelineResp_setData_1__SEL_2 ||
	     WILL_FIRE_RL_cache_pipelineResp_mRs ;
  assign cache_cRqMshr$EN_pipelineResp_setStateSlot =
	     WILL_FIRE_RL_cache_pipelineResp_cRs &&
	     cache_pipeline$first[517] ||
	     WILL_FIRE_RL_cache_pipelineResp_cRq ||
	     WILL_FIRE_RL_cache_pipelineResp_mRs ;
  assign cache_cRqMshr$EN_pipelineResp_setAddrSucc =
	     WILL_FIRE_RL_cache_pipelineResp_cRq &&
	     (cache_pipeline$first[517] &&
	      !cache_pipeline_first__581_BITS_516_TO_513_583__ETC___d2588 &&
	      cache_cRqMshr$pipelineResp_searchEndOfChain[4] ||
	      !cache_pipeline$first[517] &&
	      cache_cRqMshr$pipelineResp_searchEndOfChain[4] &&
	      cache_cRqMshr$pipelineResp_getState == 3'd1) ;
  assign cache_cRqMshr$EN_pipelineResp_setRepSucc =
	     WILL_FIRE_RL_cache_pipelineResp_cRq &&
	     cache_pipeline$first[517] &&
	     !cache_pipeline_first__581_BITS_516_TO_513_583__ETC___d2588 &&
	     !cache_cRqMshr$pipelineResp_searchEndOfChain[4] ;
  assign cache_cRqMshr$EN_stuck_get = EN_cRqStuck_get ;
  // submodule cache_cRqRetryIndexQ_clearReq_dummy2_0
  assign cache_cRqRetryIndexQ_clearReq_dummy2_0$D_IN = 1'b0 ;
  assign cache_cRqRetryIndexQ_clearReq_dummy2_0$EN = 1'b0 ;
  // submodule cache_cRqRetryIndexQ_clearReq_dummy2_1
  assign cache_cRqRetryIndexQ_clearReq_dummy2_1$D_IN = 1'd1 ;
  assign cache_cRqRetryIndexQ_clearReq_dummy2_1$EN = 1'd1 ;
  // submodule cache_cRqRetryIndexQ_deqReq_dummy2_0
  assign cache_cRqRetryIndexQ_deqReq_dummy2_0$D_IN = 1'd1 ;
  assign cache_cRqRetryIndexQ_deqReq_dummy2_0$EN =
	     WILL_FIRE_RL_cache_cRqTransfer_retry ;
  // submodule cache_cRqRetryIndexQ_deqReq_dummy2_1
  assign cache_cRqRetryIndexQ_deqReq_dummy2_1$D_IN = 1'b0 ;
  assign cache_cRqRetryIndexQ_deqReq_dummy2_1$EN = 1'b0 ;
  // submodule cache_cRqRetryIndexQ_deqReq_dummy2_2
  assign cache_cRqRetryIndexQ_deqReq_dummy2_2$D_IN = 1'd1 ;
  assign cache_cRqRetryIndexQ_deqReq_dummy2_2$EN = 1'd1 ;
  // submodule cache_cRqRetryIndexQ_enqReq_dummy2_0
  assign cache_cRqRetryIndexQ_enqReq_dummy2_0$D_IN = 1'd1 ;
  assign cache_cRqRetryIndexQ_enqReq_dummy2_0$EN =
	     WILL_FIRE_RL_cache_pipelineResp_cRq &&
	     NOT_cache_pipeline_first__581_BIT_517_582_105__ETC___d3332 ||
	     WILL_FIRE_RL_cache_pipelineResp_cRs &&
	     cache_pipeline$first[517] &&
	     cache_pipeline$first[512] &&
	     IF_SEL_ARR_cache_pipeline_first__581_BITS_519__ETC___d3488 &&
	     cache_cRqMshr$pipelineResp_getRepSucc[4] ;
  // submodule cache_cRqRetryIndexQ_enqReq_dummy2_1
  assign cache_cRqRetryIndexQ_enqReq_dummy2_1$D_IN = 1'b0 ;
  assign cache_cRqRetryIndexQ_enqReq_dummy2_1$EN = 1'b0 ;
  // submodule cache_cRqRetryIndexQ_enqReq_dummy2_2
  assign cache_cRqRetryIndexQ_enqReq_dummy2_2$D_IN = 1'd1 ;
  assign cache_cRqRetryIndexQ_enqReq_dummy2_2$EN = 1'd1 ;
  // submodule cache_pipeline
  always@(WILL_FIRE_RL_cache_pipelineResp_mRs or
	  cache_cRqMshr$pipelineResp_getAddrSucc or
	  WILL_FIRE_RL_cache_pipelineResp_cRq or
	  MUX_cache_pipeline$deqWrite_1__VAL_2 or
	  WILL_FIRE_RL_cache_pipelineResp_cRs or
	  MUX_cache_pipeline$deqWrite_1__VAL_3)
  begin
    case (1'b1) // synopsys parallel_case
      WILL_FIRE_RL_cache_pipelineResp_mRs:
	  cache_pipeline$deqWrite_swapRq =
	      cache_cRqMshr$pipelineResp_getAddrSucc;
      WILL_FIRE_RL_cache_pipelineResp_cRq:
	  cache_pipeline$deqWrite_swapRq =
	      MUX_cache_pipeline$deqWrite_1__VAL_2;
      WILL_FIRE_RL_cache_pipelineResp_cRs:
	  cache_pipeline$deqWrite_swapRq =
	      MUX_cache_pipeline$deqWrite_1__VAL_3;
      default: cache_pipeline$deqWrite_swapRq =
		   5'b01010 /* unspecified value */ ;
    endcase
  end
  always@(WILL_FIRE_RL_cache_pipelineResp_mRs or
	  WILL_FIRE_RL_cache_pipelineResp_cRq or
	  MUX_cache_pipeline$deqWrite_3__VAL_2 or
	  WILL_FIRE_RL_cache_pipelineResp_cRs or
	  MUX_cache_pipeline$deqWrite_3__VAL_3)
  begin
    case (1'b1) // synopsys parallel_case
      WILL_FIRE_RL_cache_pipelineResp_mRs:
	  cache_pipeline$deqWrite_updateRep = 1'd1;
      WILL_FIRE_RL_cache_pipelineResp_cRq:
	  cache_pipeline$deqWrite_updateRep =
	      MUX_cache_pipeline$deqWrite_3__VAL_2;
      WILL_FIRE_RL_cache_pipelineResp_cRs:
	  cache_pipeline$deqWrite_updateRep =
	      MUX_cache_pipeline$deqWrite_3__VAL_3;
      default: cache_pipeline$deqWrite_updateRep =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(WILL_FIRE_RL_cache_pipelineResp_mRs or
	  MUX_cache_pipeline$deqWrite_2__VAL_1 or
	  WILL_FIRE_RL_cache_pipelineResp_cRq or
	  MUX_cache_pipeline$deqWrite_2__VAL_2 or
	  WILL_FIRE_RL_cache_pipelineResp_cRs or
	  MUX_cache_pipeline$deqWrite_2__VAL_3)
  begin
    case (1'b1) // synopsys parallel_case
      WILL_FIRE_RL_cache_pipelineResp_mRs:
	  cache_pipeline$deqWrite_wrRam =
	      MUX_cache_pipeline$deqWrite_2__VAL_1;
      WILL_FIRE_RL_cache_pipelineResp_cRq:
	  cache_pipeline$deqWrite_wrRam =
	      MUX_cache_pipeline$deqWrite_2__VAL_2;
      WILL_FIRE_RL_cache_pipelineResp_cRs:
	  cache_pipeline$deqWrite_wrRam =
	      MUX_cache_pipeline$deqWrite_2__VAL_3;
      default: cache_pipeline$deqWrite_wrRam =
		   574'h2AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA /* unspecified value */ ;
    endcase
  end
  always@(WILL_FIRE_RL_cache_cRqTransfer_retry or
	  MUX_cache_pipeline$send_1__VAL_1 or
	  WILL_FIRE_RL_cache_cRqTransfer_new_child or
	  MUX_cache_pipeline$send_1__VAL_2 or
	  WILL_FIRE_RL_cache_cRqTransfer_new_dma or
	  MUX_cache_pipeline$send_1__VAL_3 or
	  WILL_FIRE_RL_cache_cRsTransfer or
	  MUX_cache_pipeline$send_1__VAL_4 or
	  WILL_FIRE_RL_cache_mRsTransfer or MUX_cache_pipeline$send_1__VAL_5)
  begin
    case (1'b1) // synopsys parallel_case
      WILL_FIRE_RL_cache_cRqTransfer_retry:
	  cache_pipeline$send_r = MUX_cache_pipeline$send_1__VAL_1;
      WILL_FIRE_RL_cache_cRqTransfer_new_child:
	  cache_pipeline$send_r = MUX_cache_pipeline$send_1__VAL_2;
      WILL_FIRE_RL_cache_cRqTransfer_new_dma:
	  cache_pipeline$send_r = MUX_cache_pipeline$send_1__VAL_3;
      WILL_FIRE_RL_cache_cRsTransfer:
	  cache_pipeline$send_r = MUX_cache_pipeline$send_1__VAL_4;
      WILL_FIRE_RL_cache_mRsTransfer:
	  cache_pipeline$send_r = MUX_cache_pipeline$send_1__VAL_5;
      default: cache_pipeline$send_r =
		   584'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA /* unspecified value */ ;
    endcase
  end
  assign cache_pipeline$EN_send =
	     WILL_FIRE_RL_cache_cRqTransfer_retry ||
	     WILL_FIRE_RL_cache_cRqTransfer_new_child ||
	     WILL_FIRE_RL_cache_cRqTransfer_new_dma ||
	     WILL_FIRE_RL_cache_cRsTransfer ||
	     WILL_FIRE_RL_cache_mRsTransfer ;
  assign cache_pipeline$EN_deqWrite =
	     WILL_FIRE_RL_cache_pipelineResp_mRs ||
	     WILL_FIRE_RL_cache_pipelineResp_cRq ||
	     WILL_FIRE_RL_cache_pipelineResp_cRs ;
  // submodule cache_rqFromCQ_clearReq_dummy2_0
  assign cache_rqFromCQ_clearReq_dummy2_0$D_IN = 1'b0 ;
  assign cache_rqFromCQ_clearReq_dummy2_0$EN = 1'b0 ;
  // submodule cache_rqFromCQ_clearReq_dummy2_1
  assign cache_rqFromCQ_clearReq_dummy2_1$D_IN = 1'd1 ;
  assign cache_rqFromCQ_clearReq_dummy2_1$EN = 1'd1 ;
  // submodule cache_rqFromCQ_deqReq_dummy2_0
  assign cache_rqFromCQ_deqReq_dummy2_0$D_IN = 1'd1 ;
  assign cache_rqFromCQ_deqReq_dummy2_0$EN =
	     WILL_FIRE_RL_cache_cRqTransfer_new_child ;
  // submodule cache_rqFromCQ_deqReq_dummy2_1
  assign cache_rqFromCQ_deqReq_dummy2_1$D_IN = 1'b0 ;
  assign cache_rqFromCQ_deqReq_dummy2_1$EN = 1'b0 ;
  // submodule cache_rqFromCQ_deqReq_dummy2_2
  assign cache_rqFromCQ_deqReq_dummy2_2$D_IN = 1'd1 ;
  assign cache_rqFromCQ_deqReq_dummy2_2$EN = 1'd1 ;
  // submodule cache_rqFromCQ_enqReq_dummy2_0
  assign cache_rqFromCQ_enqReq_dummy2_0$D_IN = 1'd1 ;
  assign cache_rqFromCQ_enqReq_dummy2_0$EN = EN_to_child_rqFromC_enq ;
  // submodule cache_rqFromCQ_enqReq_dummy2_1
  assign cache_rqFromCQ_enqReq_dummy2_1$D_IN = 1'b0 ;
  assign cache_rqFromCQ_enqReq_dummy2_1$EN = 1'b0 ;
  // submodule cache_rqFromCQ_enqReq_dummy2_2
  assign cache_rqFromCQ_enqReq_dummy2_2$D_IN = 1'd1 ;
  assign cache_rqFromCQ_enqReq_dummy2_2$EN = 1'd1 ;
  // submodule cache_rqFromDmaQ_clearReq_dummy2_0
  assign cache_rqFromDmaQ_clearReq_dummy2_0$D_IN = 1'b0 ;
  assign cache_rqFromDmaQ_clearReq_dummy2_0$EN = 1'b0 ;
  // submodule cache_rqFromDmaQ_clearReq_dummy2_1
  assign cache_rqFromDmaQ_clearReq_dummy2_1$D_IN = 1'd1 ;
  assign cache_rqFromDmaQ_clearReq_dummy2_1$EN = 1'd1 ;
  // submodule cache_rqFromDmaQ_deqReq_dummy2_0
  assign cache_rqFromDmaQ_deqReq_dummy2_0$D_IN = 1'd1 ;
  assign cache_rqFromDmaQ_deqReq_dummy2_0$EN =
	     WILL_FIRE_RL_cache_cRqTransfer_new_dma ;
  // submodule cache_rqFromDmaQ_deqReq_dummy2_1
  assign cache_rqFromDmaQ_deqReq_dummy2_1$D_IN = 1'b0 ;
  assign cache_rqFromDmaQ_deqReq_dummy2_1$EN = 1'b0 ;
  // submodule cache_rqFromDmaQ_deqReq_dummy2_2
  assign cache_rqFromDmaQ_deqReq_dummy2_2$D_IN = 1'd1 ;
  assign cache_rqFromDmaQ_deqReq_dummy2_2$EN = 1'd1 ;
  // submodule cache_rqFromDmaQ_enqReq_dummy2_0
  assign cache_rqFromDmaQ_enqReq_dummy2_0$D_IN = 1'd1 ;
  assign cache_rqFromDmaQ_enqReq_dummy2_0$EN = EN_dma_memReq_enq ;
  // submodule cache_rqFromDmaQ_enqReq_dummy2_1
  assign cache_rqFromDmaQ_enqReq_dummy2_1$D_IN = 1'b0 ;
  assign cache_rqFromDmaQ_enqReq_dummy2_1$EN = 1'b0 ;
  // submodule cache_rqFromDmaQ_enqReq_dummy2_2
  assign cache_rqFromDmaQ_enqReq_dummy2_2$D_IN = 1'd1 ;
  assign cache_rqFromDmaQ_enqReq_dummy2_2$EN = 1'd1 ;
  // submodule cache_rsFromCQ_clearReq_dummy2_0
  assign cache_rsFromCQ_clearReq_dummy2_0$D_IN = 1'b0 ;
  assign cache_rsFromCQ_clearReq_dummy2_0$EN = 1'b0 ;
  // submodule cache_rsFromCQ_clearReq_dummy2_1
  assign cache_rsFromCQ_clearReq_dummy2_1$D_IN = 1'd1 ;
  assign cache_rsFromCQ_clearReq_dummy2_1$EN = 1'd1 ;
  // submodule cache_rsFromCQ_deqReq_dummy2_0
  assign cache_rsFromCQ_deqReq_dummy2_0$D_IN = 1'd1 ;
  assign cache_rsFromCQ_deqReq_dummy2_0$EN = WILL_FIRE_RL_cache_cRsTransfer ;
  // submodule cache_rsFromCQ_deqReq_dummy2_1
  assign cache_rsFromCQ_deqReq_dummy2_1$D_IN = 1'b0 ;
  assign cache_rsFromCQ_deqReq_dummy2_1$EN = 1'b0 ;
  // submodule cache_rsFromCQ_deqReq_dummy2_2
  assign cache_rsFromCQ_deqReq_dummy2_2$D_IN = 1'd1 ;
  assign cache_rsFromCQ_deqReq_dummy2_2$EN = 1'd1 ;
  // submodule cache_rsFromCQ_enqReq_dummy2_0
  assign cache_rsFromCQ_enqReq_dummy2_0$D_IN = 1'd1 ;
  assign cache_rsFromCQ_enqReq_dummy2_0$EN = EN_to_child_rsFromC_enq ;
  // submodule cache_rsFromCQ_enqReq_dummy2_1
  assign cache_rsFromCQ_enqReq_dummy2_1$D_IN = 1'b0 ;
  assign cache_rsFromCQ_enqReq_dummy2_1$EN = 1'b0 ;
  // submodule cache_rsFromCQ_enqReq_dummy2_2
  assign cache_rsFromCQ_enqReq_dummy2_2$D_IN = 1'd1 ;
  assign cache_rsFromCQ_enqReq_dummy2_2$EN = 1'd1 ;
  // submodule cache_rsFromMQ_clearReq_dummy2_0
  assign cache_rsFromMQ_clearReq_dummy2_0$D_IN = 1'b0 ;
  assign cache_rsFromMQ_clearReq_dummy2_0$EN = 1'b0 ;
  // submodule cache_rsFromMQ_clearReq_dummy2_1
  assign cache_rsFromMQ_clearReq_dummy2_1$D_IN = 1'd1 ;
  assign cache_rsFromMQ_clearReq_dummy2_1$EN = 1'd1 ;
  // submodule cache_rsFromMQ_deqReq_dummy2_0
  assign cache_rsFromMQ_deqReq_dummy2_0$D_IN = 1'd1 ;
  assign cache_rsFromMQ_deqReq_dummy2_0$EN =
	     cache_rsFromMQ_deqReq_lat_0$whas ;
  // submodule cache_rsFromMQ_deqReq_dummy2_1
  assign cache_rsFromMQ_deqReq_dummy2_1$D_IN = 1'b0 ;
  assign cache_rsFromMQ_deqReq_dummy2_1$EN = 1'b0 ;
  // submodule cache_rsFromMQ_deqReq_dummy2_2
  assign cache_rsFromMQ_deqReq_dummy2_2$D_IN = 1'd1 ;
  assign cache_rsFromMQ_deqReq_dummy2_2$EN = 1'd1 ;
  // submodule cache_rsFromMQ_enqReq_dummy2_0
  assign cache_rsFromMQ_enqReq_dummy2_0$D_IN = 1'd1 ;
  assign cache_rsFromMQ_enqReq_dummy2_0$EN = EN_to_mem_rsFromM_enq ;
  // submodule cache_rsFromMQ_enqReq_dummy2_1
  assign cache_rsFromMQ_enqReq_dummy2_1$D_IN = 1'b0 ;
  assign cache_rsFromMQ_enqReq_dummy2_1$EN = 1'b0 ;
  // submodule cache_rsFromMQ_enqReq_dummy2_2
  assign cache_rsFromMQ_enqReq_dummy2_2$D_IN = 1'd1 ;
  assign cache_rsFromMQ_enqReq_dummy2_2$EN = 1'd1 ;
  // submodule cache_rsLdToDmaIndexQ
  assign cache_rsLdToDmaIndexQ$D_IN =
	     WILL_FIRE_RL_cache_mergeRsLdToDmaIndexQ_mRsDeq ?
	       cache_rsLdToDmaIndexQ_mRsDeq$D_OUT :
	       cache_rsLdToDmaIndexQ_pipelineResp$D_OUT ;
  assign cache_rsLdToDmaIndexQ$ENQ =
	     WILL_FIRE_RL_cache_mergeRsLdToDmaIndexQ_mRsDeq ||
	     WILL_FIRE_RL_cache_mergeRsLdToDmaIndexQ_pipelineResp ;
  assign cache_rsLdToDmaIndexQ$DEQ = CAN_FIRE_RL_cache_sendRsLdToDma ;
  assign cache_rsLdToDmaIndexQ$CLR = 1'b0 ;
  // submodule cache_rsLdToDmaIndexQ_mRsDeq
  assign cache_rsLdToDmaIndexQ_mRsDeq$D_IN =
	     MUX_cache_cRqMshr$transfer_getRq_1__VAL_2 ;
  assign cache_rsLdToDmaIndexQ_mRsDeq$ENQ =
	     CAN_FIRE_RL_cache_mRsDeq_nonRefill ;
  assign cache_rsLdToDmaIndexQ_mRsDeq$DEQ =
	     WILL_FIRE_RL_cache_mergeRsLdToDmaIndexQ_mRsDeq ;
  assign cache_rsLdToDmaIndexQ_mRsDeq$CLR = 1'b0 ;
  // submodule cache_rsLdToDmaIndexQ_pipelineResp
  assign cache_rsLdToDmaIndexQ_pipelineResp$D_IN =
	     MUX_cache_rsLdToDmaIndexQ_pipelineResp$enq_1__SEL_1 ?
	       cache_pipeline$first[582:579] :
	       cache_pipeline$first[516:513] ;
  assign cache_rsLdToDmaIndexQ_pipelineResp$ENQ =
	     WILL_FIRE_RL_cache_pipelineResp_cRq &&
	     (cache_pipeline_first__581_BIT_517_582_AND_cach_ETC___d3139 ||
	      NOT_cache_pipeline_first__581_BIT_517_582_105__ETC___d3143) ||
	     WILL_FIRE_RL_cache_pipelineResp_cRs &&
	     cache_pipeline_first__581_BIT_517_582_AND_NOT__ETC___d3824 ;
  assign cache_rsLdToDmaIndexQ_pipelineResp$DEQ =
	     CAN_FIRE_RL_cache_mergeRsLdToDmaIndexQ_pipelineResp ;
  assign cache_rsLdToDmaIndexQ_pipelineResp$CLR = 1'b0 ;
  // submodule cache_rsLdToDmaQ_clearReq_dummy2_0
  assign cache_rsLdToDmaQ_clearReq_dummy2_0$D_IN = 1'b0 ;
  assign cache_rsLdToDmaQ_clearReq_dummy2_0$EN = 1'b0 ;
  // submodule cache_rsLdToDmaQ_clearReq_dummy2_1
  assign cache_rsLdToDmaQ_clearReq_dummy2_1$D_IN = 1'd1 ;
  assign cache_rsLdToDmaQ_clearReq_dummy2_1$EN = 1'd1 ;
  // submodule cache_rsLdToDmaQ_deqReq_dummy2_0
  assign cache_rsLdToDmaQ_deqReq_dummy2_0$D_IN = 1'd1 ;
  assign cache_rsLdToDmaQ_deqReq_dummy2_0$EN = EN_dma_respLd_deq ;
  // submodule cache_rsLdToDmaQ_deqReq_dummy2_1
  assign cache_rsLdToDmaQ_deqReq_dummy2_1$D_IN = 1'b0 ;
  assign cache_rsLdToDmaQ_deqReq_dummy2_1$EN = 1'b0 ;
  // submodule cache_rsLdToDmaQ_deqReq_dummy2_2
  assign cache_rsLdToDmaQ_deqReq_dummy2_2$D_IN = 1'd1 ;
  assign cache_rsLdToDmaQ_deqReq_dummy2_2$EN = 1'd1 ;
  // submodule cache_rsLdToDmaQ_enqReq_dummy2_0
  assign cache_rsLdToDmaQ_enqReq_dummy2_0$D_IN = 1'd1 ;
  assign cache_rsLdToDmaQ_enqReq_dummy2_0$EN =
	     CAN_FIRE_RL_cache_sendRsLdToDma ;
  // submodule cache_rsLdToDmaQ_enqReq_dummy2_1
  assign cache_rsLdToDmaQ_enqReq_dummy2_1$D_IN = 1'b0 ;
  assign cache_rsLdToDmaQ_enqReq_dummy2_1$EN = 1'b0 ;
  // submodule cache_rsLdToDmaQ_enqReq_dummy2_2
  assign cache_rsLdToDmaQ_enqReq_dummy2_2$D_IN = 1'd1 ;
  assign cache_rsLdToDmaQ_enqReq_dummy2_2$EN = 1'd1 ;
  // submodule cache_rsStToDmaIndexQ
  assign cache_rsStToDmaIndexQ$D_IN =
	     WILL_FIRE_RL_cache_mergeRsStToDmaIndexQ_sendToM ?
	       cache_rsStToDmaIndexQ_sendToM$D_OUT :
	       cache_rsStToDmaIndexQ_pipelineResp$D_OUT ;
  assign cache_rsStToDmaIndexQ$ENQ =
	     WILL_FIRE_RL_cache_mergeRsStToDmaIndexQ_sendToM ||
	     WILL_FIRE_RL_cache_mergeRsStToDmaIndexQ_pipelineResp ;
  assign cache_rsStToDmaIndexQ$DEQ = WILL_FIRE_RL_cache_sendRsStToDma ;
  assign cache_rsStToDmaIndexQ$CLR = 1'b0 ;
  // submodule cache_rsStToDmaIndexQ_pipelineResp
  assign cache_rsStToDmaIndexQ_pipelineResp$D_IN =
	     MUX_cache_rsStToDmaIndexQ_pipelineResp$enq_1__SEL_1 ?
	       cache_pipeline$first[582:579] :
	       cache_pipeline$first[516:513] ;
  assign cache_rsStToDmaIndexQ_pipelineResp$ENQ =
	     WILL_FIRE_RL_cache_pipelineResp_cRq &&
	     (cache_pipeline_first__581_BIT_517_582_AND_cach_ETC___d3129 ||
	      NOT_cache_pipeline_first__581_BIT_517_582_105__ETC___d3133) ||
	     WILL_FIRE_RL_cache_pipelineResp_cRs &&
	     cache_pipeline_first__581_BIT_517_582_AND_NOT__ETC___d3820 ;
  assign cache_rsStToDmaIndexQ_pipelineResp$DEQ =
	     CAN_FIRE_RL_cache_mergeRsStToDmaIndexQ_pipelineResp ;
  assign cache_rsStToDmaIndexQ_pipelineResp$CLR = 1'b0 ;
  // submodule cache_rsStToDmaIndexQ_sendToM
  assign cache_rsStToDmaIndexQ_sendToM$D_IN = cache_toMInfoQ$D_OUT[5:2] ;
  assign cache_rsStToDmaIndexQ_sendToM$ENQ =
	     WILL_FIRE_RL_cache_sendToM && cache_toMInfoQ$D_OUT[1:0] == 2'd1 ;
  assign cache_rsStToDmaIndexQ_sendToM$DEQ =
	     WILL_FIRE_RL_cache_mergeRsStToDmaIndexQ_sendToM ;
  assign cache_rsStToDmaIndexQ_sendToM$CLR = 1'b0 ;
  // submodule cache_rsStToDmaQ_clearReq_dummy2_0
  assign cache_rsStToDmaQ_clearReq_dummy2_0$D_IN = 1'b0 ;
  assign cache_rsStToDmaQ_clearReq_dummy2_0$EN = 1'b0 ;
  // submodule cache_rsStToDmaQ_clearReq_dummy2_1
  assign cache_rsStToDmaQ_clearReq_dummy2_1$D_IN = 1'd1 ;
  assign cache_rsStToDmaQ_clearReq_dummy2_1$EN = 1'd1 ;
  // submodule cache_rsStToDmaQ_deqReq_dummy2_0
  assign cache_rsStToDmaQ_deqReq_dummy2_0$D_IN = 1'd1 ;
  assign cache_rsStToDmaQ_deqReq_dummy2_0$EN = EN_dma_respSt_deq ;
  // submodule cache_rsStToDmaQ_deqReq_dummy2_1
  assign cache_rsStToDmaQ_deqReq_dummy2_1$D_IN = 1'b0 ;
  assign cache_rsStToDmaQ_deqReq_dummy2_1$EN = 1'b0 ;
  // submodule cache_rsStToDmaQ_deqReq_dummy2_2
  assign cache_rsStToDmaQ_deqReq_dummy2_2$D_IN = 1'd1 ;
  assign cache_rsStToDmaQ_deqReq_dummy2_2$EN = 1'd1 ;
  // submodule cache_rsStToDmaQ_enqReq_dummy2_0
  assign cache_rsStToDmaQ_enqReq_dummy2_0$D_IN = 1'd1 ;
  assign cache_rsStToDmaQ_enqReq_dummy2_0$EN =
	     WILL_FIRE_RL_cache_sendRsStToDma ;
  // submodule cache_rsStToDmaQ_enqReq_dummy2_1
  assign cache_rsStToDmaQ_enqReq_dummy2_1$D_IN = 1'b0 ;
  assign cache_rsStToDmaQ_enqReq_dummy2_1$EN = 1'b0 ;
  // submodule cache_rsStToDmaQ_enqReq_dummy2_2
  assign cache_rsStToDmaQ_enqReq_dummy2_2$D_IN = 1'd1 ;
  assign cache_rsStToDmaQ_enqReq_dummy2_2$EN = 1'd1 ;
  // submodule cache_rsToCIndexQ_clearReq_dummy2_0
  assign cache_rsToCIndexQ_clearReq_dummy2_0$D_IN = 1'b0 ;
  assign cache_rsToCIndexQ_clearReq_dummy2_0$EN = 1'b0 ;
  // submodule cache_rsToCIndexQ_clearReq_dummy2_1
  assign cache_rsToCIndexQ_clearReq_dummy2_1$D_IN = 1'd1 ;
  assign cache_rsToCIndexQ_clearReq_dummy2_1$EN = 1'd1 ;
  // submodule cache_rsToCIndexQ_deqReq_dummy2_0
  assign cache_rsToCIndexQ_deqReq_dummy2_0$D_IN = 1'd1 ;
  assign cache_rsToCIndexQ_deqReq_dummy2_0$EN = WILL_FIRE_RL_cache_sendRsToC ;
  // submodule cache_rsToCIndexQ_deqReq_dummy2_1
  assign cache_rsToCIndexQ_deqReq_dummy2_1$D_IN = 1'b0 ;
  assign cache_rsToCIndexQ_deqReq_dummy2_1$EN = 1'b0 ;
  // submodule cache_rsToCIndexQ_deqReq_dummy2_2
  assign cache_rsToCIndexQ_deqReq_dummy2_2$D_IN = 1'd1 ;
  assign cache_rsToCIndexQ_deqReq_dummy2_2$EN = 1'd1 ;
  // submodule cache_rsToCIndexQ_enqReq_dummy2_0
  assign cache_rsToCIndexQ_enqReq_dummy2_0$D_IN = 1'd1 ;
  assign cache_rsToCIndexQ_enqReq_dummy2_0$EN =
	     WILL_FIRE_RL_cache_pipelineResp_cRq &&
	     (cache_pipeline_first__581_BIT_517_582_AND_cach_ETC___d3146 ||
	      NOT_cache_pipeline_first__581_BIT_517_582_105__ETC___d3149) ||
	     WILL_FIRE_RL_cache_pipelineResp_cRs &&
	     cache_pipeline$first[517] &&
	     !cache_pipeline$first[512] &&
	     IF_SEL_ARR_cache_cRqMshr_pipelineResp_getSlot__ETC___d3484 &&
	     !cache_cRqMshr$pipelineResp_getRq[16] ||
	     WILL_FIRE_RL_cache_pipelineResp_mRs ;
  // submodule cache_rsToCIndexQ_enqReq_dummy2_1
  assign cache_rsToCIndexQ_enqReq_dummy2_1$D_IN = 1'b0 ;
  assign cache_rsToCIndexQ_enqReq_dummy2_1$EN = 1'b0 ;
  // submodule cache_rsToCIndexQ_enqReq_dummy2_2
  assign cache_rsToCIndexQ_enqReq_dummy2_2$D_IN = 1'd1 ;
  assign cache_rsToCIndexQ_enqReq_dummy2_2$EN = 1'd1 ;
  // submodule cache_toCQ_clearReq_dummy2_0
  assign cache_toCQ_clearReq_dummy2_0$D_IN = 1'b0 ;
  assign cache_toCQ_clearReq_dummy2_0$EN = 1'b0 ;
  // submodule cache_toCQ_clearReq_dummy2_1
  assign cache_toCQ_clearReq_dummy2_1$D_IN = 1'd1 ;
  assign cache_toCQ_clearReq_dummy2_1$EN = 1'd1 ;
  // submodule cache_toCQ_deqReq_dummy2_0
  assign cache_toCQ_deqReq_dummy2_0$D_IN = 1'd1 ;
  assign cache_toCQ_deqReq_dummy2_0$EN = EN_to_child_toC_deq ;
  // submodule cache_toCQ_deqReq_dummy2_1
  assign cache_toCQ_deqReq_dummy2_1$D_IN = 1'b0 ;
  assign cache_toCQ_deqReq_dummy2_1$EN = 1'b0 ;
  // submodule cache_toCQ_deqReq_dummy2_2
  assign cache_toCQ_deqReq_dummy2_2$D_IN = 1'd1 ;
  assign cache_toCQ_deqReq_dummy2_2$EN = 1'd1 ;
  // submodule cache_toCQ_enqReq_dummy2_0
  assign cache_toCQ_enqReq_dummy2_0$D_IN = 1'd1 ;
  assign cache_toCQ_enqReq_dummy2_0$EN =
	     WILL_FIRE_RL_cache_sendRqToC || WILL_FIRE_RL_cache_sendRsToC ;
  // submodule cache_toCQ_enqReq_dummy2_1
  assign cache_toCQ_enqReq_dummy2_1$D_IN = 1'b0 ;
  assign cache_toCQ_enqReq_dummy2_1$EN = 1'b0 ;
  // submodule cache_toCQ_enqReq_dummy2_2
  assign cache_toCQ_enqReq_dummy2_2$D_IN = 1'd1 ;
  assign cache_toCQ_enqReq_dummy2_2$EN = 1'd1 ;
  // submodule cache_toMInfoQ
  assign cache_toMInfoQ$D_IN =
	     MUX_cache_toMInfoQ$enq_1__SEL_1 ?
	       MUX_cache_toMInfoQ$enq_1__VAL_1 :
	       MUX_cache_toMInfoQ$enq_1__VAL_2 ;
  assign cache_toMInfoQ$ENQ =
	     MUX_cache_toMInfoQ$enq_1__SEL_1 ||
	     WILL_FIRE_RL_cache_pipelineResp_cRs &&
	     cache_pipeline$first[517] &&
	     cache_pipeline$first[512] &&
	     IF_SEL_ARR_cache_pipeline_first__581_BITS_519__ETC___d3488 ;
  assign cache_toMInfoQ$DEQ =
	     WILL_FIRE_RL_cache_sendToM &&
	     (cache_toMInfoQ$D_OUT[1:0] == 2'd0 ||
	      cache_toMInfoQ$D_OUT[1:0] == 2'd1 ||
	      cache_toMInfoQ$D_OUT[1:0] == 2'd2 && cache_doLdAfterReplace) ;
  assign cache_toMInfoQ$CLR = 1'b0 ;
  // submodule cache_toMQ_clearReq_dummy2_0
  assign cache_toMQ_clearReq_dummy2_0$D_IN = 1'b0 ;
  assign cache_toMQ_clearReq_dummy2_0$EN = 1'b0 ;
  // submodule cache_toMQ_clearReq_dummy2_1
  assign cache_toMQ_clearReq_dummy2_1$D_IN = 1'd1 ;
  assign cache_toMQ_clearReq_dummy2_1$EN = 1'd1 ;
  // submodule cache_toMQ_deqReq_dummy2_0
  assign cache_toMQ_deqReq_dummy2_0$D_IN = 1'd1 ;
  assign cache_toMQ_deqReq_dummy2_0$EN = EN_to_mem_toM_deq ;
  // submodule cache_toMQ_deqReq_dummy2_1
  assign cache_toMQ_deqReq_dummy2_1$D_IN = 1'b0 ;
  assign cache_toMQ_deqReq_dummy2_1$EN = 1'b0 ;
  // submodule cache_toMQ_deqReq_dummy2_2
  assign cache_toMQ_deqReq_dummy2_2$D_IN = 1'd1 ;
  assign cache_toMQ_deqReq_dummy2_2$EN = 1'd1 ;
  // submodule cache_toMQ_enqReq_dummy2_0
  assign cache_toMQ_enqReq_dummy2_0$D_IN = 1'd1 ;
  assign cache_toMQ_enqReq_dummy2_0$EN = cache_toMQ_enqReq_lat_0$whas ;
  // submodule cache_toMQ_enqReq_dummy2_1
  assign cache_toMQ_enqReq_dummy2_1$D_IN = 1'b0 ;
  assign cache_toMQ_enqReq_dummy2_1$EN = 1'b0 ;
  // submodule cache_toMQ_enqReq_dummy2_2
  assign cache_toMQ_enqReq_dummy2_2$D_IN = 1'd1 ;
  assign cache_toMQ_enqReq_dummy2_2$EN = 1'd1 ;
  // submodule perfReqQ_clearReq_dummy2_0
  assign perfReqQ_clearReq_dummy2_0$D_IN = 1'b0 ;
  assign perfReqQ_clearReq_dummy2_0$EN = 1'b0 ;
  // submodule perfReqQ_clearReq_dummy2_1
  assign perfReqQ_clearReq_dummy2_1$D_IN = 1'd1 ;
  assign perfReqQ_clearReq_dummy2_1$EN = 1'd1 ;
  // submodule perfReqQ_deqReq_dummy2_0
  assign perfReqQ_deqReq_dummy2_0$D_IN = 1'd1 ;
  assign perfReqQ_deqReq_dummy2_0$EN = EN_perf_resp ;
  // submodule perfReqQ_deqReq_dummy2_1
  assign perfReqQ_deqReq_dummy2_1$D_IN = 1'b0 ;
  assign perfReqQ_deqReq_dummy2_1$EN = 1'b0 ;
  // submodule perfReqQ_deqReq_dummy2_2
  assign perfReqQ_deqReq_dummy2_2$D_IN = 1'd1 ;
  assign perfReqQ_deqReq_dummy2_2$EN = 1'd1 ;
  // submodule perfReqQ_enqReq_dummy2_0
  assign perfReqQ_enqReq_dummy2_0$D_IN = 1'd1 ;
  assign perfReqQ_enqReq_dummy2_0$EN = EN_perf_req ;
  // submodule perfReqQ_enqReq_dummy2_1
  assign perfReqQ_enqReq_dummy2_1$D_IN = 1'b0 ;
  assign perfReqQ_enqReq_dummy2_1$EN = 1'b0 ;
  // submodule perfReqQ_enqReq_dummy2_2
  assign perfReqQ_enqReq_dummy2_2$D_IN = 1'd1 ;
  assign perfReqQ_enqReq_dummy2_2$EN = 1'd1 ;
  // remaining internal signals
  assign DONTCARE_CONCAT_SEL_ARR_cache_toCQ_data_0_917__ETC___d3940 =
	     { 516'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA,
	       CASE_cache_toCQ_deqP_0_cache_toCQ_data_0_BITS__ETC__q249,
	       CASE_cache_toCQ_deqP_0_cache_toCQ_data_0_BITS__ETC__q250,
	       x__h444361 } ;
  assign DONTCARE_CONCAT_SEL_ARR_cache_toMQ_data_0_050__ETC___d4073 =
	     { 571'h2AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA,
	       CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BITS__ETC__q252,
	       CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_4_ETC__q253,
	       x__h456804 } ;
  assign IF_IF_SEL_ARR_cache_pipeline_first__581_BITS_5_ETC___d3709 =
	     IF_SEL_ARR_cache_pipeline_first__581_BITS_519__ETC___d3488 ?
	       { cache_pipeline$first[578:575],
		 cache_pipeline$first[573:526],
		 13'd4642 } :
	       { cache_cRqMshr$pipelineResp_getSlot[64:12],
		 IF_SEL_ARR_cache_pipeline_first__581_BITS_519__ETC___d3694,
		 (SEL_ARR_cache_pipeline_first__581_BITS_519_TO__ETC___d3403 ==
		  2'd0) ?
		   IF_IF_cache_pipeline_first__581_BITS_584_TO_58_ETC___d3697 :
		   cache_cRqMshr$pipelineResp_getSlot[3:2],
		 cache_cRqMshr$pipelineResp_getSlot[1:0] } ;
  assign IF_IF_cache_cRqMshr_pipelineResp_getRq_IF_cach_ETC___d2635 =
	     IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2627 ?
	       !cache_rsToCIndexQ_full :
	       cache_pipeline$first[525:524] != 2'd0 ||
	       cache_toMInfoQ$FULL_N ;
  assign IF_IF_cache_cRqMshr_pipelineResp_getRq_IF_cach_ETC___d2699 =
	     IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2627 ?
	       { IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2686,
		 IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2697,
		 cache_cRqMshr$pipelineResp_getAddrSucc,
		 1'd0 } :
	       { cache_pipeline$first[525:518],
		 1'd1,
		 cache_pipeline$first[582:579],
		 1'd0 } ;
  assign IF_IF_cache_cRqMshr_pipelineResp_getRq_IF_cach_ETC___d3397 =
	     { (IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3388 ==
		2'd3) ?
		 IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3388 :
		 cache_pipeline$first[525:524],
	       IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3396,
	       cache_cRqMshr$pipelineResp_getAddrSucc,
	       1'd0 } ;
  assign IF_IF_cache_pipeline_first__581_BITS_584_TO_58_ETC___d3672 =
	     (cache_pipeline$first[580:579] == 2'd2 ||
	      cache_cRqMshr$pipelineResp_getSlot[11:10] == 2'd0) ?
	       2'd0 :
	       cache_cRqMshr$pipelineResp_getSlot[11:10] ;
  assign IF_IF_cache_pipeline_first__581_BITS_584_TO_58_ETC___d3684 =
	     (cache_pipeline$first[580:579] == 2'd1 ||
	      cache_cRqMshr$pipelineResp_getSlot[7:6] == 2'd0) ?
	       2'd0 :
	       cache_cRqMshr$pipelineResp_getSlot[7:6] ;
  assign IF_IF_cache_pipeline_first__581_BITS_584_TO_58_ETC___d3697 =
	     (cache_pipeline$first[580:579] == 2'd0 ||
	      cache_cRqMshr$pipelineResp_getSlot[3:2] == 2'd0) ?
	       2'd0 :
	       cache_cRqMshr$pipelineResp_getSlot[3:2] ;
  assign IF_NOT_SEL_ARR_NOT_cache_rqFromDmaQ_data_0_129_ETC___d1646 =
	     (!CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q68 ||
	      NOT_SEL_ARR_NOT_cache_rqFromDmaQ_data_0_129_BI_ETC___d1644) ?
	       2'd3 :
	       2'd1 ;
  assign IF_NOT_cache_cRqMshr_pipelineResp_getRq_IF_cac_ETC___d3054 =
	     (cache_cRqMshr$pipelineResp_getRq[82:81] != 2'd2 &&
	      !cache_pipeline_first__581_BITS_523_TO_522_603__ETC___d2604) ?
	       IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2597 :
	       cache_cRqMshr$pipelineResp_getRq[87:86] ;
  assign IF_NOT_cache_cRqMshr_pipelineResp_getRq_IF_cac_ETC___d3063 =
	     (cache_cRqMshr$pipelineResp_getRq[82:81] != 2'd1 &&
	      !cache_pipeline_first__581_BITS_521_TO_520_600__ETC___d2601) ?
	       IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2597 :
	       cache_cRqMshr$pipelineResp_getRq[87:86] ;
  assign IF_NOT_cache_cRqMshr_pipelineResp_getRq_IF_cac_ETC___d3073 =
	     (cache_cRqMshr$pipelineResp_getRq[82:81] != 2'd0 &&
	      !cache_pipeline_first__581_BITS_519_TO_518_594__ETC___d2598) ?
	       IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2597 :
	       cache_cRqMshr$pipelineResp_getRq[87:86] ;
  assign IF_NOT_cache_pipeline_first__581_BITS_525_TO_5_ETC___d2654 =
	     (cache_pipeline$first[525:524] != 2'd0 &&
	      cache_pipeline_first__581_BITS_573_TO_526_644__ETC___d2646) ?
	       _0_OR_NOT_cache_pipeline_first__581_BITS_519_TO_ETC___d2614 :
	       cache_toMInfoQ$FULL_N &&
	       (!cache_cRqMshr$pipelineResp_getAddrSucc[4] ||
		!cache_cRqRetryIndexQ_full) ;
  assign IF_NOT_cache_pipeline_first__581_BITS_525_TO_5_ETC___d2657 =
	     (cache_pipeline$first[525:524] != 2'd0 &&
	      IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2627) ?
	       !cache_rsToCIndexQ_full :
	       cache_pipeline$first[525:524] != 2'd0 ||
	       cache_toMInfoQ$FULL_N ;
  assign IF_NOT_cache_pipeline_first__581_BITS_525_TO_5_ETC___d2999 =
	     (cache_pipeline$first[525:524] != 2'd0 &&
	      cache_pipeline_first__581_BITS_573_TO_526_644__ETC___d2646) ?
	       { cache_cRqMshr$pipelineResp_getRq[151:104],
		 IF_cache_pipeline_first__581_BITS_519_TO_518_5_ETC___d2693,
		 IF_cache_pipeline_first__581_BITS_519_TO_518_5_ETC___d2993 } :
	       cache_pipeline$first[573:0] ;
  assign IF_NOT_cache_pipeline_first__581_BITS_525_TO_5_ETC___d3000 =
	     (cache_pipeline$first[525:524] != 2'd0 &&
	      IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2627) ?
	       { IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2686,
		 IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2697,
		 cache_cRqMshr$pipelineResp_getAddrSucc,
		 1'd0 } :
	       { cache_pipeline$first[525:518],
		 1'd1,
		 cache_pipeline$first[582:579],
		 1'd0 } ;
  assign IF_SEL_ARR_IF_cache_cRqMshr_pipelineResp_getSl_ETC___d3481 =
	     SEL_ARR_IF_cache_cRqMshr_pipelineResp_getSlot__ETC___d3440 ?
	       cache_cRqMshr$pipelineResp_getSlot[3:2] == 2'd0 &&
	       cache_cRqMshr$pipelineResp_getSlot[7:6] == 2'd0 &&
	       cache_cRqMshr$pipelineResp_getSlot[11:10] == 2'd0 :
	       (cache_pipeline$first[580:579] == 2'd0 ||
		cache_cRqMshr$pipelineResp_getSlot[3:2] == 2'd0) &&
	       (cache_pipeline$first[580:579] == 2'd1 ||
		cache_cRqMshr$pipelineResp_getSlot[7:6] == 2'd0) &&
	       (cache_pipeline$first[580:579] == 2'd2 ||
		cache_cRqMshr$pipelineResp_getSlot[11:10] == 2'd0) ;
  assign IF_SEL_ARR_IF_cache_cRqMshr_pipelineResp_getSl_ETC___d3482 =
	     SEL_ARR_IF_cache_cRqMshr_pipelineResp_getSlot__ETC___d3440 ?
	       cache_cRqMshr$pipelineResp_getSlot[3:2] == 2'd0 &&
	       cache_cRqMshr$pipelineResp_getSlot[7:6] == 2'd0 &&
	       cache_cRqMshr$pipelineResp_getSlot[11:10] == 2'd0 :
	       (cache_pipeline$first[580:579] == 2'd0 ||
		cache_cRqMshr$pipelineResp_getSlot[3:2] == 2'd0) &&
	       (cache_pipeline$first[580:579] == 2'd1 ||
		cache_cRqMshr$pipelineResp_getSlot[7:6] == 2'd0) &&
	       (cache_pipeline$first[580:579] == 2'd2 ||
		cache_cRqMshr$pipelineResp_getSlot[11:10] == 2'd0) ;
  assign IF_SEL_ARR_NOT_cache_toCQ_data_0_917_BIT_584_9_ETC___d4000 =
	     CASE_cache_toCQ_deqP_0_NOT_cache_toCQ_data_0_B_ETC__q255 ?
	       DONTCARE_CONCAT_SEL_ARR_cache_toCQ_data_0_917__ETC___d3940 :
	       SEL_ARR_cache_toCQ_data_0_917_BITS_583_TO_520__ETC___d3998 ;
  assign IF_SEL_ARR_NOT_cache_toMQ_data_0_050_BIT_640_0_ETC___d4404 =
	     CASE_cache_toMQ_deqP_0_NOT_cache_toMQ_data_0_B_ETC__q260 ?
	       DONTCARE_CONCAT_SEL_ARR_cache_toMQ_data_0_050__ETC___d4073 :
	       SEL_ARR_cache_toMQ_data_0_050_BITS_639_TO_576__ETC___d4402 ;
  assign IF_SEL_ARR_cache_cRqMshr_pipelineResp_getSlot__ETC___d3454 =
	     SEL_ARR_cache_cRqMshr_pipelineResp_getSlot_IF__ETC___d3446 ?
	       (SEL_ARR_IF_cache_cRqMshr_pipelineResp_getSlot__ETC___d3440 ?
		  cache_cRqMshr$pipelineResp_getSlot[3:2] != 2'd0 :
		  cache_pipeline$first[580:579] != 2'd0 &&
		  cache_cRqMshr$pipelineResp_getSlot[3:2] != 2'd0) :
	       cache_cRqMshr$pipelineResp_getSlot[3:2] != 2'd0 ;
  assign IF_SEL_ARR_cache_cRqMshr_pipelineResp_getSlot__ETC___d3455 =
	     SEL_ARR_cache_cRqMshr_pipelineResp_getSlot_IF__ETC___d3431 ?
	       (SEL_ARR_IF_cache_cRqMshr_pipelineResp_getSlot__ETC___d3440 ?
		  cache_cRqMshr$pipelineResp_getSlot[3:2] != 2'd0 :
		  cache_pipeline$first[580:579] != 2'd0 &&
		  cache_cRqMshr$pipelineResp_getSlot[3:2] != 2'd0) :
	       IF_SEL_ARR_cache_cRqMshr_pipelineResp_getSlot__ETC___d3454 ;
  assign IF_SEL_ARR_cache_cRqMshr_pipelineResp_getSlot__ETC___d3458 =
	     SEL_ARR_cache_cRqMshr_pipelineResp_getSlot_IF__ETC___d3446 ?
	       (SEL_ARR_IF_cache_cRqMshr_pipelineResp_getSlot__ETC___d3440 ?
		  cache_cRqMshr$pipelineResp_getSlot[7:6] != 2'd0 :
		  cache_pipeline$first[580:579] != 2'd1 &&
		  cache_cRqMshr$pipelineResp_getSlot[7:6] != 2'd0) :
	       cache_cRqMshr$pipelineResp_getSlot[7:6] != 2'd0 ;
  assign IF_SEL_ARR_cache_cRqMshr_pipelineResp_getSlot__ETC___d3459 =
	     SEL_ARR_cache_cRqMshr_pipelineResp_getSlot_IF__ETC___d3431 ?
	       (SEL_ARR_IF_cache_cRqMshr_pipelineResp_getSlot__ETC___d3440 ?
		  cache_cRqMshr$pipelineResp_getSlot[7:6] != 2'd0 :
		  cache_pipeline$first[580:579] != 2'd1 &&
		  cache_cRqMshr$pipelineResp_getSlot[7:6] != 2'd0) :
	       IF_SEL_ARR_cache_cRqMshr_pipelineResp_getSlot__ETC___d3458 ;
  assign IF_SEL_ARR_cache_cRqMshr_pipelineResp_getSlot__ETC___d3462 =
	     SEL_ARR_cache_cRqMshr_pipelineResp_getSlot_IF__ETC___d3446 ?
	       (SEL_ARR_IF_cache_cRqMshr_pipelineResp_getSlot__ETC___d3440 ?
		  cache_cRqMshr$pipelineResp_getSlot[11:10] != 2'd0 :
		  cache_pipeline$first[580:579] != 2'd2 &&
		  cache_cRqMshr$pipelineResp_getSlot[11:10] != 2'd0) :
	       cache_cRqMshr$pipelineResp_getSlot[11:10] != 2'd0 ;
  assign IF_SEL_ARR_cache_cRqMshr_pipelineResp_getSlot__ETC___d3463 =
	     SEL_ARR_cache_cRqMshr_pipelineResp_getSlot_IF__ETC___d3431 ?
	       (SEL_ARR_IF_cache_cRqMshr_pipelineResp_getSlot__ETC___d3440 ?
		  cache_cRqMshr$pipelineResp_getSlot[11:10] != 2'd0 :
		  cache_pipeline$first[580:579] != 2'd2 &&
		  cache_cRqMshr$pipelineResp_getSlot[11:10] != 2'd0) :
	       IF_SEL_ARR_cache_cRqMshr_pipelineResp_getSlot__ETC___d3462 ;
  assign IF_SEL_ARR_cache_cRqMshr_pipelineResp_getSlot__ETC___d3484 =
	     SEL_ARR_cache_cRqMshr_pipelineResp_getSlot_IF__ETC___d3431 ?
	       IF_SEL_ARR_IF_cache_cRqMshr_pipelineResp_getSl_ETC___d3481 :
	       (SEL_ARR_cache_cRqMshr_pipelineResp_getSlot_IF__ETC___d3446 ?
		  IF_SEL_ARR_IF_cache_cRqMshr_pipelineResp_getSl_ETC___d3482 :
		  cache_cRqMshr$pipelineResp_getSlot[3:2] == 2'd0 &&
		  cache_cRqMshr$pipelineResp_getSlot[7:6] == 2'd0 &&
		  cache_cRqMshr$pipelineResp_getSlot[11:10] == 2'd0) ;
  assign IF_SEL_ARR_cache_cRqMshr_pipelineResp_getSlot__ETC___d3712 =
	     SEL_ARR_cache_cRqMshr_pipelineResp_getSlot_IF__ETC___d3446 ?
	       (SEL_ARR_IF_cache_cRqMshr_pipelineResp_getSlot__ETC___d3440 ?
		  cache_cRqMshr$pipelineResp_getSlot[11:10] :
		  IF_IF_cache_pipeline_first__581_BITS_584_TO_58_ETC___d3672) :
	       cache_cRqMshr$pipelineResp_getSlot[11:10] ;
  assign IF_SEL_ARR_cache_cRqMshr_pipelineResp_getSlot__ETC___d3713 =
	     SEL_ARR_cache_cRqMshr_pipelineResp_getSlot_IF__ETC___d3431 ?
	       (SEL_ARR_IF_cache_cRqMshr_pipelineResp_getSlot__ETC___d3440 ?
		  cache_cRqMshr$pipelineResp_getSlot[11:10] :
		  IF_IF_cache_pipeline_first__581_BITS_584_TO_58_ETC___d3672) :
	       IF_SEL_ARR_cache_cRqMshr_pipelineResp_getSlot__ETC___d3712 ;
  assign IF_SEL_ARR_cache_cRqMshr_pipelineResp_getSlot__ETC___d3726 =
	     SEL_ARR_cache_cRqMshr_pipelineResp_getSlot_IF__ETC___d3446 ?
	       (SEL_ARR_IF_cache_cRqMshr_pipelineResp_getSlot__ETC___d3440 ?
		  cache_cRqMshr$pipelineResp_getSlot[7:6] :
		  IF_IF_cache_pipeline_first__581_BITS_584_TO_58_ETC___d3684) :
	       cache_cRqMshr$pipelineResp_getSlot[7:6] ;
  assign IF_SEL_ARR_cache_cRqMshr_pipelineResp_getSlot__ETC___d3727 =
	     SEL_ARR_cache_cRqMshr_pipelineResp_getSlot_IF__ETC___d3431 ?
	       (SEL_ARR_IF_cache_cRqMshr_pipelineResp_getSlot__ETC___d3440 ?
		  cache_cRqMshr$pipelineResp_getSlot[7:6] :
		  IF_IF_cache_pipeline_first__581_BITS_584_TO_58_ETC___d3684) :
	       IF_SEL_ARR_cache_cRqMshr_pipelineResp_getSlot__ETC___d3726 ;
  assign IF_SEL_ARR_cache_cRqMshr_pipelineResp_getSlot__ETC___d3741 =
	     SEL_ARR_cache_cRqMshr_pipelineResp_getSlot_IF__ETC___d3446 ?
	       (SEL_ARR_IF_cache_cRqMshr_pipelineResp_getSlot__ETC___d3440 ?
		  cache_cRqMshr$pipelineResp_getSlot[3:2] :
		  IF_IF_cache_pipeline_first__581_BITS_584_TO_58_ETC___d3697) :
	       cache_cRqMshr$pipelineResp_getSlot[3:2] ;
  assign IF_SEL_ARR_cache_cRqMshr_pipelineResp_getSlot__ETC___d3742 =
	     SEL_ARR_cache_cRqMshr_pipelineResp_getSlot_IF__ETC___d3431 ?
	       (SEL_ARR_IF_cache_cRqMshr_pipelineResp_getSlot__ETC___d3440 ?
		  cache_cRqMshr$pipelineResp_getSlot[3:2] :
		  IF_IF_cache_pipeline_first__581_BITS_584_TO_58_ETC___d3697) :
	       IF_SEL_ARR_cache_cRqMshr_pipelineResp_getSlot__ETC___d3741 ;
  assign IF_SEL_ARR_cache_cRqMshr_pipelineResp_getSlot__ETC___d3804 =
	     IF_SEL_ARR_cache_cRqMshr_pipelineResp_getSlot__ETC___d3484 &&
	     cache_cRqMshr$pipelineResp_getRq[16] &&
	     (!cache_pipeline_first__581_BITS_573_TO_526_644__ETC___d2646 ||
	      cache_pipeline$first[525:524] == 2'd0) ;
  assign IF_SEL_ARR_cache_cRqMshr_pipelineResp_getSlot__ETC___d3814 =
	     IF_SEL_ARR_cache_cRqMshr_pipelineResp_getSlot__ETC___d3484 &&
	     cache_cRqMshr$pipelineResp_getRq[16] &&
	     cache_cRqMshr$pipelineResp_getData[512] !=
	     (cache_cRqMshr$pipelineResp_getRq[17] ||
	      cache_cRqMshr$pipelineResp_getRq[18] ||
	      cache_cRqMshr$pipelineResp_getRq[19] ||
	      cache_cRqMshr$pipelineResp_getRq[20] ||
	      cache_cRqMshr$pipelineResp_getRq[21] ||
	      cache_cRqMshr$pipelineResp_getRq[22] ||
	      cache_cRqMshr$pipelineResp_getRq[23] ||
	      cache_cRqMshr$pipelineResp_getRq[24] ||
	      cache_cRqMshr$pipelineResp_getRq[25] ||
	      cache_cRqMshr$pipelineResp_getRq[26] ||
	      cache_cRqMshr$pipelineResp_getRq[27] ||
	      cache_cRqMshr$pipelineResp_getRq[28] ||
	      cache_cRqMshr$pipelineResp_getRq[29] ||
	      cache_cRqMshr$pipelineResp_getRq[30] ||
	      cache_cRqMshr$pipelineResp_getRq[31] ||
	      cache_cRqMshr$pipelineResp_getRq[32] ||
	      cache_cRqMshr$pipelineResp_getRq[33] ||
	      cache_cRqMshr$pipelineResp_getRq[34] ||
	      cache_cRqMshr$pipelineResp_getRq[35] ||
	      cache_cRqMshr$pipelineResp_getRq[36] ||
	      cache_cRqMshr$pipelineResp_getRq[37] ||
	      cache_cRqMshr$pipelineResp_getRq[38] ||
	      cache_cRqMshr$pipelineResp_getRq[39] ||
	      cache_cRqMshr$pipelineResp_getRq[40] ||
	      cache_cRqMshr$pipelineResp_getRq[41] ||
	      cache_cRqMshr$pipelineResp_getRq[42] ||
	      cache_cRqMshr$pipelineResp_getRq[43] ||
	      cache_cRqMshr$pipelineResp_getRq[44] ||
	      cache_cRqMshr$pipelineResp_getRq[45] ||
	      cache_cRqMshr$pipelineResp_getRq[46] ||
	      cache_cRqMshr$pipelineResp_getRq[47] ||
	      cache_cRqMshr$pipelineResp_getRq[48] ||
	      cache_cRqMshr$pipelineResp_getRq[49] ||
	      cache_cRqMshr$pipelineResp_getRq[50] ||
	      cache_cRqMshr$pipelineResp_getRq[51] ||
	      cache_cRqMshr$pipelineResp_getRq[52] ||
	      cache_cRqMshr$pipelineResp_getRq[53] ||
	      cache_cRqMshr$pipelineResp_getRq[54] ||
	      cache_cRqMshr$pipelineResp_getRq[55] ||
	      cache_cRqMshr$pipelineResp_getRq[56] ||
	      cache_cRqMshr$pipelineResp_getRq[57] ||
	      cache_cRqMshr$pipelineResp_getRq[58] ||
	      cache_cRqMshr$pipelineResp_getRq[59] ||
	      cache_cRqMshr$pipelineResp_getRq[60] ||
	      cache_cRqMshr$pipelineResp_getRq[61] ||
	      cache_cRqMshr$pipelineResp_getRq[62] ||
	      cache_cRqMshr$pipelineResp_getRq[63] ||
	      cache_cRqMshr$pipelineResp_getRq[64] ||
	      cache_cRqMshr$pipelineResp_getRq[65] ||
	      cache_cRqMshr$pipelineResp_getRq[66] ||
	      cache_cRqMshr$pipelineResp_getRq[67] ||
	      cache_cRqMshr$pipelineResp_getRq[68] ||
	      cache_cRqMshr$pipelineResp_getRq[69] ||
	      cache_cRqMshr$pipelineResp_getRq[70] ||
	      cache_cRqMshr$pipelineResp_getRq[71] ||
	      cache_cRqMshr$pipelineResp_getRq[72] ||
	      cache_cRqMshr$pipelineResp_getRq[73] ||
	      cache_cRqMshr$pipelineResp_getRq[74] ||
	      cache_cRqMshr$pipelineResp_getRq[75] ||
	      cache_cRqMshr$pipelineResp_getRq[76] ||
	      cache_cRqMshr$pipelineResp_getRq[77] ||
	      cache_cRqMshr$pipelineResp_getRq[78] ||
	      cache_cRqMshr$pipelineResp_getRq[79] ||
	      cache_cRqMshr$pipelineResp_getRq[80]) ;
  assign IF_SEL_ARR_cache_cRqMshr_pipelineResp_getSlot__ETC___d3830 =
	     IF_SEL_ARR_cache_cRqMshr_pipelineResp_getSlot__ETC___d3484 &&
	     !cache_cRqMshr$pipelineResp_getRq[16] &&
	     (!cache_pipeline_first__581_BITS_573_TO_526_644__ETC___d2646 ||
	      cache_pipeline$first[525:524] == 2'd0) ;
  assign IF_SEL_ARR_cache_pipeline_first__581_BITS_519__ETC___d3417 =
	     (SEL_ARR_cache_pipeline_first__581_BITS_519_TO__ETC___d3403 ==
	      2'd0) ?
	       cache_pipeline$first[580:579] != 2'd1 &&
	       cache_cRqMshr$pipelineResp_getSlot[7:6] != 2'd0 ||
	       cache_pipeline$first[580:579] != 2'd2 &&
	       cache_cRqMshr$pipelineResp_getSlot[11:10] != 2'd0 :
	       cache_cRqMshr$pipelineResp_getSlot[7:6] != 2'd0 ||
	       cache_cRqMshr$pipelineResp_getSlot[11:10] != 2'd0 ;
  assign IF_SEL_ARR_cache_pipeline_first__581_BITS_519__ETC___d3418 =
	     ((SEL_ARR_cache_pipeline_first__581_BITS_519_TO__ETC___d3403 ==
	       2'd0) ?
		cache_pipeline$first[580:579] != 2'd0 &&
		cache_cRqMshr$pipelineResp_getSlot[3:2] != 2'd0 :
		cache_cRqMshr$pipelineResp_getSlot[3:2] != 2'd0) ||
	     IF_SEL_ARR_cache_pipeline_first__581_BITS_519__ETC___d3417 ;
  assign IF_SEL_ARR_cache_pipeline_first__581_BITS_519__ETC___d3488 =
	     (SEL_ARR_cache_pipeline_first__581_BITS_519_TO__ETC___d3403 ==
	      2'd0) ?
	       (cache_pipeline$first[580:579] == 2'd0 ||
		cache_cRqMshr$pipelineResp_getSlot[3:2] == 2'd0) &&
	       (cache_pipeline$first[580:579] == 2'd1 ||
		cache_cRqMshr$pipelineResp_getSlot[7:6] == 2'd0) &&
	       (cache_pipeline$first[580:579] == 2'd2 ||
		cache_cRqMshr$pipelineResp_getSlot[11:10] == 2'd0) :
	       cache_cRqMshr$pipelineResp_getSlot[3:2] == 2'd0 &&
	       cache_cRqMshr$pipelineResp_getSlot[7:6] == 2'd0 &&
	       cache_cRqMshr$pipelineResp_getSlot[11:10] == 2'd0 ;
  assign IF_SEL_ARR_cache_pipeline_first__581_BITS_519__ETC___d3694 =
	     { (SEL_ARR_cache_pipeline_first__581_BITS_519_TO__ETC___d3403 ==
		2'd0) ?
		 IF_IF_cache_pipeline_first__581_BITS_584_TO_58_ETC___d3672 :
		 cache_cRqMshr$pipelineResp_getSlot[11:10],
	       cache_cRqMshr$pipelineResp_getSlot[9:8],
	       (SEL_ARR_cache_pipeline_first__581_BITS_519_TO__ETC___d3403 ==
		2'd0) ?
		 IF_IF_cache_pipeline_first__581_BITS_584_TO_58_ETC___d3684 :
		 cache_cRqMshr$pipelineResp_getSlot[7:6],
	       cache_cRqMshr$pipelineResp_getSlot[5:4] } ;
  assign IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2597 =
	     (cache_cRqMshr$pipelineResp_getRq[85:84] == 2'd1) ?
	       cache_cRqMshr$pipelineResp_getRq[85:84] :
	       2'd0 ;
  assign IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2626 =
	     ((cache_cRqMshr$pipelineResp_getRq[82:81] == 2'd1) ?
		cache_pipeline_first__581_BITS_521_TO_520_600__ETC___d2621 :
		cache_pipeline_first__581_BITS_521_TO_520_600__ETC___d2601) &&
	     ((cache_cRqMshr$pipelineResp_getRq[82:81] == 2'd2) ?
		cache_pipeline_first__581_BITS_523_TO_522_603__ETC___d2624 :
		cache_pipeline_first__581_BITS_523_TO_522_603__ETC___d2604) ;
  assign IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2627 =
	     ((cache_cRqMshr$pipelineResp_getRq[82:81] == 2'd0) ?
		cache_pipeline_first__581_BITS_519_TO_518_594__ETC___d2618 :
		cache_pipeline_first__581_BITS_519_TO_518_594__ETC___d2598) &&
	     IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2626 ;
  assign IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2678 =
	     cache_cRqMshr$pipelineResp_getRq[16] ?
	       IF_cache_pipeline_first__581_BITS_519_TO_518_5_ETC___d2676 :
	       (IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2627 ?
		  cache_cRqMshr$pipelineResp_getAddrSucc :
		  5'd10) ;
  assign IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2683 =
	     cache_cRqMshr$pipelineResp_getRq[16] ?
	       ((cache_pipeline$first[525:524] != 2'd0 &&
		 cache_pipeline_first__581_BITS_573_TO_526_644__ETC___d2646) ?
		  IF_cache_pipeline_first__581_BITS_519_TO_518_5_ETC___d2676 :
		  5'd10) :
	       IF_cache_pipeline_first__581_BITS_525_TO_524_6_ETC___d2682 ;
  assign IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2686 =
	     (cache_cRqMshr$pipelineResp_getRq[85:84] == 2'd3) ?
	       cache_cRqMshr$pipelineResp_getRq[85:84] :
	       cache_pipeline$first[525:524] ;
  assign IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2697 =
	     { (cache_cRqMshr$pipelineResp_getRq[82:81] == 2'd2) ?
		 cache_cRqMshr$pipelineResp_getRq[85:84] :
		 cache_pipeline$first[523:522],
	       (cache_cRqMshr$pipelineResp_getRq[82:81] == 2'd1) ?
		 cache_cRqMshr$pipelineResp_getRq[85:84] :
		 cache_pipeline$first[521:520],
	       (cache_cRqMshr$pipelineResp_getRq[82:81] == 2'd0) ?
		 cache_cRqMshr$pipelineResp_getRq[85:84] :
		 cache_pipeline$first[519:518] } ;
  assign IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2714 =
	     { cache_cRqMshr$pipelineResp_getRq[80] ?
		 cache_cRqMshr$pipelineResp_getData[511:504] :
		 cache_pipeline$first[511:504],
	       cache_cRqMshr$pipelineResp_getRq[79] ?
		 cache_cRqMshr$pipelineResp_getData[503:496] :
		 cache_pipeline$first[503:496],
	       cache_cRqMshr$pipelineResp_getRq[78] ?
		 cache_cRqMshr$pipelineResp_getData[495:488] :
		 cache_pipeline$first[495:488] } ;
  assign IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2723 =
	     { IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2714,
	       cache_cRqMshr$pipelineResp_getRq[77] ?
		 cache_cRqMshr$pipelineResp_getData[487:480] :
		 cache_pipeline$first[487:480],
	       cache_cRqMshr$pipelineResp_getRq[76] ?
		 cache_cRqMshr$pipelineResp_getData[479:472] :
		 cache_pipeline$first[479:472] } ;
  assign IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2732 =
	     { IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2723,
	       cache_cRqMshr$pipelineResp_getRq[75] ?
		 cache_cRqMshr$pipelineResp_getData[471:464] :
		 cache_pipeline$first[471:464],
	       cache_cRqMshr$pipelineResp_getRq[74] ?
		 cache_cRqMshr$pipelineResp_getData[463:456] :
		 cache_pipeline$first[463:456] } ;
  assign IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2749 =
	     { cache_cRqMshr$pipelineResp_getRq[72] ?
		 cache_cRqMshr$pipelineResp_getData[447:440] :
		 cache_pipeline$first[447:440],
	       cache_cRqMshr$pipelineResp_getRq[71] ?
		 cache_cRqMshr$pipelineResp_getData[439:432] :
		 cache_pipeline$first[439:432],
	       cache_cRqMshr$pipelineResp_getRq[70] ?
		 cache_cRqMshr$pipelineResp_getData[431:424] :
		 cache_pipeline$first[431:424] } ;
  assign IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2758 =
	     { IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2749,
	       cache_cRqMshr$pipelineResp_getRq[69] ?
		 cache_cRqMshr$pipelineResp_getData[423:416] :
		 cache_pipeline$first[423:416],
	       cache_cRqMshr$pipelineResp_getRq[68] ?
		 cache_cRqMshr$pipelineResp_getData[415:408] :
		 cache_pipeline$first[415:408] } ;
  assign IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2767 =
	     { IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2758,
	       cache_cRqMshr$pipelineResp_getRq[67] ?
		 cache_cRqMshr$pipelineResp_getData[407:400] :
		 cache_pipeline$first[407:400],
	       cache_cRqMshr$pipelineResp_getRq[66] ?
		 cache_cRqMshr$pipelineResp_getData[399:392] :
		 cache_pipeline$first[399:392] } ;
  assign IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2772 =
	     { IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2732,
	       cache_cRqMshr$pipelineResp_getRq[73] ?
		 cache_cRqMshr$pipelineResp_getData[455:448] :
		 cache_pipeline$first[455:448],
	       IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2767,
	       cache_cRqMshr$pipelineResp_getRq[65] ?
		 cache_cRqMshr$pipelineResp_getData[391:384] :
		 cache_pipeline$first[391:384] } ;
  assign IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2790 =
	     { cache_cRqMshr$pipelineResp_getRq[64] ?
		 cache_cRqMshr$pipelineResp_getData[383:376] :
		 cache_pipeline$first[383:376],
	       cache_cRqMshr$pipelineResp_getRq[63] ?
		 cache_cRqMshr$pipelineResp_getData[375:368] :
		 cache_pipeline$first[375:368],
	       cache_cRqMshr$pipelineResp_getRq[62] ?
		 cache_cRqMshr$pipelineResp_getData[367:360] :
		 cache_pipeline$first[367:360],
	       cache_cRqMshr$pipelineResp_getRq[61] ?
		 cache_cRqMshr$pipelineResp_getData[359:352] :
		 cache_pipeline$first[359:352] } ;
  assign IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2799 =
	     { IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2790,
	       cache_cRqMshr$pipelineResp_getRq[60] ?
		 cache_cRqMshr$pipelineResp_getData[351:344] :
		 cache_pipeline$first[351:344],
	       cache_cRqMshr$pipelineResp_getRq[59] ?
		 cache_cRqMshr$pipelineResp_getData[343:336] :
		 cache_pipeline$first[343:336] } ;
  assign IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2808 =
	     { IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2799,
	       cache_cRqMshr$pipelineResp_getRq[58] ?
		 cache_cRqMshr$pipelineResp_getData[335:328] :
		 cache_pipeline$first[335:328],
	       cache_cRqMshr$pipelineResp_getRq[57] ?
		 cache_cRqMshr$pipelineResp_getData[327:320] :
		 cache_pipeline$first[327:320] } ;
  assign IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2821 =
	     { cache_cRqMshr$pipelineResp_getRq[56] ?
		 cache_cRqMshr$pipelineResp_getData[319:312] :
		 cache_pipeline$first[319:312],
	       cache_cRqMshr$pipelineResp_getRq[55] ?
		 cache_cRqMshr$pipelineResp_getData[311:304] :
		 cache_pipeline$first[311:304],
	       cache_cRqMshr$pipelineResp_getRq[54] ?
		 cache_cRqMshr$pipelineResp_getData[303:296] :
		 cache_pipeline$first[303:296] } ;
  assign IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2830 =
	     { IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2821,
	       cache_cRqMshr$pipelineResp_getRq[53] ?
		 cache_cRqMshr$pipelineResp_getData[295:288] :
		 cache_pipeline$first[295:288],
	       cache_cRqMshr$pipelineResp_getRq[52] ?
		 cache_cRqMshr$pipelineResp_getData[287:280] :
		 cache_pipeline$first[287:280] } ;
  assign IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2839 =
	     { IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2830,
	       cache_cRqMshr$pipelineResp_getRq[51] ?
		 cache_cRqMshr$pipelineResp_getData[279:272] :
		 cache_pipeline$first[279:272],
	       cache_cRqMshr$pipelineResp_getRq[50] ?
		 cache_cRqMshr$pipelineResp_getData[271:264] :
		 cache_pipeline$first[271:264] } ;
  assign IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2844 =
	     { IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2772,
	       IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2808,
	       IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2839,
	       cache_cRqMshr$pipelineResp_getRq[49] ?
		 cache_cRqMshr$pipelineResp_getData[263:256] :
		 cache_pipeline$first[263:256] } ;
  assign IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2862 =
	     { cache_cRqMshr$pipelineResp_getRq[48] ?
		 cache_cRqMshr$pipelineResp_getData[255:248] :
		 cache_pipeline$first[255:248],
	       cache_cRqMshr$pipelineResp_getRq[47] ?
		 cache_cRqMshr$pipelineResp_getData[247:240] :
		 cache_pipeline$first[247:240],
	       cache_cRqMshr$pipelineResp_getRq[46] ?
		 cache_cRqMshr$pipelineResp_getData[239:232] :
		 cache_pipeline$first[239:232],
	       cache_cRqMshr$pipelineResp_getRq[45] ?
		 cache_cRqMshr$pipelineResp_getData[231:224] :
		 cache_pipeline$first[231:224] } ;
  assign IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2871 =
	     { IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2862,
	       cache_cRqMshr$pipelineResp_getRq[44] ?
		 cache_cRqMshr$pipelineResp_getData[223:216] :
		 cache_pipeline$first[223:216],
	       cache_cRqMshr$pipelineResp_getRq[43] ?
		 cache_cRqMshr$pipelineResp_getData[215:208] :
		 cache_pipeline$first[215:208] } ;
  assign IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2880 =
	     { IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2871,
	       cache_cRqMshr$pipelineResp_getRq[42] ?
		 cache_cRqMshr$pipelineResp_getData[207:200] :
		 cache_pipeline$first[207:200],
	       cache_cRqMshr$pipelineResp_getRq[41] ?
		 cache_cRqMshr$pipelineResp_getData[199:192] :
		 cache_pipeline$first[199:192] } ;
  assign IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2893 =
	     { cache_cRqMshr$pipelineResp_getRq[40] ?
		 cache_cRqMshr$pipelineResp_getData[191:184] :
		 cache_pipeline$first[191:184],
	       cache_cRqMshr$pipelineResp_getRq[39] ?
		 cache_cRqMshr$pipelineResp_getData[183:176] :
		 cache_pipeline$first[183:176],
	       cache_cRqMshr$pipelineResp_getRq[38] ?
		 cache_cRqMshr$pipelineResp_getData[175:168] :
		 cache_pipeline$first[175:168] } ;
  assign IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2902 =
	     { IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2893,
	       cache_cRqMshr$pipelineResp_getRq[37] ?
		 cache_cRqMshr$pipelineResp_getData[167:160] :
		 cache_pipeline$first[167:160],
	       cache_cRqMshr$pipelineResp_getRq[36] ?
		 cache_cRqMshr$pipelineResp_getData[159:152] :
		 cache_pipeline$first[159:152] } ;
  assign IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2911 =
	     { IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2902,
	       cache_cRqMshr$pipelineResp_getRq[35] ?
		 cache_cRqMshr$pipelineResp_getData[151:144] :
		 cache_pipeline$first[151:144],
	       cache_cRqMshr$pipelineResp_getRq[34] ?
		 cache_cRqMshr$pipelineResp_getData[143:136] :
		 cache_pipeline$first[143:136] } ;
  assign IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2916 =
	     { IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2844,
	       IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2880,
	       IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2911,
	       cache_cRqMshr$pipelineResp_getRq[33] ?
		 cache_cRqMshr$pipelineResp_getData[135:128] :
		 cache_pipeline$first[135:128] } ;
  assign IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2934 =
	     { cache_cRqMshr$pipelineResp_getRq[32] ?
		 cache_cRqMshr$pipelineResp_getData[127:120] :
		 cache_pipeline$first[127:120],
	       cache_cRqMshr$pipelineResp_getRq[31] ?
		 cache_cRqMshr$pipelineResp_getData[119:112] :
		 cache_pipeline$first[119:112],
	       cache_cRqMshr$pipelineResp_getRq[30] ?
		 cache_cRqMshr$pipelineResp_getData[111:104] :
		 cache_pipeline$first[111:104],
	       cache_cRqMshr$pipelineResp_getRq[29] ?
		 cache_cRqMshr$pipelineResp_getData[103:96] :
		 cache_pipeline$first[103:96] } ;
  assign IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2943 =
	     { IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2934,
	       cache_cRqMshr$pipelineResp_getRq[28] ?
		 cache_cRqMshr$pipelineResp_getData[95:88] :
		 cache_pipeline$first[95:88],
	       cache_cRqMshr$pipelineResp_getRq[27] ?
		 cache_cRqMshr$pipelineResp_getData[87:80] :
		 cache_pipeline$first[87:80] } ;
  assign IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2952 =
	     { IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2943,
	       cache_cRqMshr$pipelineResp_getRq[26] ?
		 cache_cRqMshr$pipelineResp_getData[79:72] :
		 cache_pipeline$first[79:72],
	       cache_cRqMshr$pipelineResp_getRq[25] ?
		 cache_cRqMshr$pipelineResp_getData[71:64] :
		 cache_pipeline$first[71:64] } ;
  assign IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2968 =
	     { cache_cRqMshr$pipelineResp_getRq[24] ?
		 cache_cRqMshrpipelineResp_getData_BITS_63_TO_0__q78[63:56] :
		 cache_pipeline$first[63:56],
	       cache_cRqMshr$pipelineResp_getRq[23] ?
		 cache_cRqMshrpipelineResp_getData_BITS_63_TO_0__q78[55:48] :
		 cache_pipeline$first[55:48],
	       cache_cRqMshr$pipelineResp_getRq[22] ?
		 cache_cRqMshrpipelineResp_getData_BITS_63_TO_0__q78[47:40] :
		 cache_pipeline$first[47:40] } ;
  assign IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2977 =
	     { IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2968,
	       cache_cRqMshr$pipelineResp_getRq[21] ?
		 cache_cRqMshrpipelineResp_getData_BITS_63_TO_0__q78[39:32] :
		 cache_pipeline$first[39:32],
	       cache_cRqMshr$pipelineResp_getRq[20] ?
		 cache_cRqMshrpipelineResp_getData_BITS_63_TO_0__q78[31:24] :
		 cache_pipeline$first[31:24] } ;
  assign IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2986 =
	     { IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2977,
	       cache_cRqMshr$pipelineResp_getRq[19] ?
		 cache_cRqMshrpipelineResp_getData_BITS_63_TO_0__q78[23:16] :
		 cache_pipeline$first[23:16],
	       cache_cRqMshr$pipelineResp_getRq[18] ?
		 cache_cRqMshrpipelineResp_getData_BITS_63_TO_0__q78[15:8] :
		 cache_pipeline$first[15:8] } ;
  assign IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2991 =
	     { IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2916,
	       IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2952,
	       IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2986,
	       cache_cRqMshr$pipelineResp_getRq[17] ?
		 cache_cRqMshrpipelineResp_getData_BITS_63_TO_0__q78[7:0] :
		 cache_pipeline$first[7:0] } ;
  assign IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3014 =
	     cache_cRqMshr$pipelineResp_getRq[16] ?
	       cache_pipeline_first__581_BITS_519_TO_518_594__ETC___d2598 &&
	       cache_pipeline_first__581_BITS_521_TO_520_600__ETC___d2601 &&
	       cache_pipeline_first__581_BITS_523_TO_522_603__ETC___d2604 :
	       IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2627 ;
  assign IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3022 =
	     cache_cRqMshr$pipelineResp_getRq[16] ?
	       NOT_cache_pipeline_first__581_BITS_525_TO_524__ETC___d3019 :
	       cache_pipeline_first__581_BITS_573_TO_526_644__ETC___d2646 &&
	       cache_pipeline$first[525:524] != 2'd0 &&
	       IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2627 ;
  assign IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3027 =
	     cache_cRqMshr$pipelineResp_getRq[16] ?
	       IF_cache_pipeline_first__581_BITS_519_TO_518_5_ETC___d3025 :
	       (IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2627 ?
		  3'd4 :
		  3'd3) ;
  assign IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3033 =
	     cache_cRqMshr$pipelineResp_getRq[16] ?
	       ((cache_pipeline$first[525:524] != 2'd0 &&
		 cache_pipeline_first__581_BITS_573_TO_526_644__ETC___d2646) ?
		  IF_cache_pipeline_first__581_BITS_519_TO_518_5_ETC___d3025 :
		  3'd4) :
	       IF_cache_pipeline_first__581_BITS_525_TO_524_6_ETC___d3032 ;
  assign IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3048 =
	     (cache_cRqMshr$pipelineResp_getRq[82:81] == 2'd2) ?
	       (cache_pipeline_first__581_BITS_523_TO_522_603__ETC___d2624 ?
		  2'd0 :
		  2'd2) :
	       (cache_pipeline_first__581_BITS_523_TO_522_603__ETC___d2604 ?
		  2'd0 :
		  2'd1) ;
  assign IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3057 =
	     (cache_cRqMshr$pipelineResp_getRq[82:81] == 2'd1) ?
	       (cache_pipeline_first__581_BITS_521_TO_520_600__ETC___d2621 ?
		  2'd0 :
		  2'd2) :
	       (cache_pipeline_first__581_BITS_521_TO_520_600__ETC___d2601 ?
		  2'd0 :
		  2'd1) ;
  assign IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3067 =
	     (cache_cRqMshr$pipelineResp_getRq[82:81] == 2'd0) ?
	       (cache_pipeline_first__581_BITS_519_TO_518_594__ETC___d2618 ?
		  2'd0 :
		  2'd2) :
	       (cache_pipeline_first__581_BITS_519_TO_518_594__ETC___d2598 ?
		  2'd0 :
		  2'd1) ;
  assign IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3078 =
	     cache_cRqMshr$pipelineResp_getRq[16] ?
	       { cache_pipeline$first[578:575],
		 48'hAAAAAAAAAAAA,
		 _0_CONCAT_IF_cache_pipeline_first__581_BITS_523_ETC___d3043 } :
	       { cache_pipeline$first[578:575],
		 48'hAAAAAAAAAAAA,
		 cache_pipeline$first[525:524] == 2'd0,
		 IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3048,
		 IF_NOT_cache_cRqMshr_pipelineResp_getRq_IF_cac_ETC___d3054,
		 IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3057,
		 IF_NOT_cache_cRqMshr_pipelineResp_getRq_IF_cac_ETC___d3063,
		 IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3067,
		 IF_NOT_cache_cRqMshr_pipelineResp_getRq_IF_cac_ETC___d3073 } ;
  assign IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3096 =
	     cache_cRqMshr$pipelineResp_getRq[16] ?
	       { cache_pipeline$first[578:575],
		 48'hAAAAAAAAAAAA,
		 _0_CONCAT_IF_cache_pipeline_first__581_BITS_523_ETC___d3043 } :
	       IF_cache_pipeline_first__581_BITS_525_TO_524_6_ETC___d3095 ;
  assign IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3155 =
	     ((cache_cRqMshr$pipelineResp_getRq[82:81] == 2'd1) ?
		!cache_pipeline_first__581_BITS_521_TO_520_600__ETC___d2621 :
		!cache_pipeline_first__581_BITS_521_TO_520_600__ETC___d2601) ||
	     ((cache_cRqMshr$pipelineResp_getRq[82:81] == 2'd2) ?
		!cache_pipeline_first__581_BITS_523_TO_522_603__ETC___d2624 :
		!cache_pipeline_first__581_BITS_523_TO_522_603__ETC___d2604) ;
  assign IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3156 =
	     ((cache_cRqMshr$pipelineResp_getRq[82:81] == 2'd0) ?
		!cache_pipeline_first__581_BITS_519_TO_518_594__ETC___d2618 :
		!cache_pipeline_first__581_BITS_519_TO_518_594__ETC___d2598) ||
	     IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3155 ;
  assign IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3173 =
	     cache_cRqMshr$pipelineResp_getRq[16] ?
	       ((cache_cRqMshr$pipelineResp_getRq[85:84] == 2'd3) ?
		  2'd1 :
		  2'd0) :
	       ((cache_pipeline$first[525:524] == 2'd0 ||
		 cache_pipeline_first__581_BITS_573_TO_526_644__ETC___d2646) ?
		  2'd0 :
		  IF_cache_pipeline_first__581_BITS_525_TO_524_6_ETC___d3171) ;
  assign IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3388 =
	     (cache_cRqMshr$pipelineResp_getRq[85:84] == 2'd1 &&
	      cache_cRqMshr$pipelineResp_getRq[83] &&
	      cache_pipeline$first[519:518] == 2'd0 &&
	      cache_pipeline$first[521:520] == 2'd0 &&
	      cache_pipeline$first[523:522] == 2'd0) ?
	       2'd2 :
	       cache_cRqMshr$pipelineResp_getRq[85:84] ;
  assign IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3396 =
	     { (cache_cRqMshr$pipelineResp_getRq[82:81] == 2'd2) ?
		 IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3388 :
		 cache_pipeline$first[523:522],
	       (cache_cRqMshr$pipelineResp_getRq[82:81] == 2'd1) ?
		 IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3388 :
		 cache_pipeline$first[521:520],
	       (cache_cRqMshr$pipelineResp_getRq[82:81] == 2'd0) ?
		 IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3388 :
		 cache_pipeline$first[519:518] } ;
  assign IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3493 =
	     { IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2686,
	       cache_cRqMshr$pipelineResp_getRq[16] ?
		 cache_pipeline$first[523:518] :
		 IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2697,
	       cache_cRqMshr$pipelineResp_getAddrSucc,
	       1'd0 } ;
  assign IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3506 =
	     { IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2714,
	       cache_cRqMshr$pipelineResp_getRq[77] ?
		 cache_cRqMshr$pipelineResp_getData[487:480] :
		 cache_pipeline$first[487:480],
	       cache_cRqMshr$pipelineResp_getRq[76] ?
		 cache_cRqMshr$pipelineResp_getData[479:472] :
		 cache_pipeline$first[479:472] } ;
  assign IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3511 =
	     { IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3506,
	       cache_cRqMshr$pipelineResp_getRq[75] ?
		 cache_cRqMshr$pipelineResp_getData[471:464] :
		 cache_pipeline$first[471:464],
	       cache_cRqMshr$pipelineResp_getRq[74] ?
		 cache_cRqMshr$pipelineResp_getData[463:456] :
		 cache_pipeline$first[463:456] } ;
  assign IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3525 =
	     { IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2749,
	       cache_cRqMshr$pipelineResp_getRq[69] ?
		 cache_cRqMshr$pipelineResp_getData[423:416] :
		 cache_pipeline$first[423:416],
	       cache_cRqMshr$pipelineResp_getRq[68] ?
		 cache_cRqMshr$pipelineResp_getData[415:408] :
		 cache_pipeline$first[415:408] } ;
  assign IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3530 =
	     { IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3525,
	       cache_cRqMshr$pipelineResp_getRq[67] ?
		 cache_cRqMshr$pipelineResp_getData[407:400] :
		 cache_pipeline$first[407:400],
	       cache_cRqMshr$pipelineResp_getRq[66] ?
		 cache_cRqMshr$pipelineResp_getData[399:392] :
		 cache_pipeline$first[399:392] } ;
  assign IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3533 =
	     { IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3511,
	       cache_cRqMshr$pipelineResp_getRq[73] ?
		 cache_cRqMshr$pipelineResp_getData[455:448] :
		 cache_pipeline$first[455:448],
	       IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3530,
	       cache_cRqMshr$pipelineResp_getRq[65] ?
		 cache_cRqMshr$pipelineResp_getData[391:384] :
		 cache_pipeline$first[391:384] } ;
  assign IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3548 =
	     { IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2790,
	       cache_cRqMshr$pipelineResp_getRq[60] ?
		 cache_cRqMshr$pipelineResp_getData[351:344] :
		 cache_pipeline$first[351:344],
	       cache_cRqMshr$pipelineResp_getRq[59] ?
		 cache_cRqMshr$pipelineResp_getData[343:336] :
		 cache_pipeline$first[343:336] } ;
  assign IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3553 =
	     { IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3548,
	       cache_cRqMshr$pipelineResp_getRq[58] ?
		 cache_cRqMshr$pipelineResp_getData[335:328] :
		 cache_pipeline$first[335:328],
	       cache_cRqMshr$pipelineResp_getRq[57] ?
		 cache_cRqMshr$pipelineResp_getData[327:320] :
		 cache_pipeline$first[327:320] } ;
  assign IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3565 =
	     { IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2821,
	       cache_cRqMshr$pipelineResp_getRq[53] ?
		 cache_cRqMshr$pipelineResp_getData[295:288] :
		 cache_pipeline$first[295:288],
	       cache_cRqMshr$pipelineResp_getRq[52] ?
		 cache_cRqMshr$pipelineResp_getData[287:280] :
		 cache_pipeline$first[287:280] } ;
  assign IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3570 =
	     { IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3565,
	       cache_cRqMshr$pipelineResp_getRq[51] ?
		 cache_cRqMshr$pipelineResp_getData[279:272] :
		 cache_pipeline$first[279:272],
	       cache_cRqMshr$pipelineResp_getRq[50] ?
		 cache_cRqMshr$pipelineResp_getData[271:264] :
		 cache_pipeline$first[271:264] } ;
  assign IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3573 =
	     { IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3533,
	       IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3553,
	       IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3570,
	       cache_cRqMshr$pipelineResp_getRq[49] ?
		 cache_cRqMshr$pipelineResp_getData[263:256] :
		 cache_pipeline$first[263:256] } ;
  assign IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3588 =
	     { IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2862,
	       cache_cRqMshr$pipelineResp_getRq[44] ?
		 cache_cRqMshr$pipelineResp_getData[223:216] :
		 cache_pipeline$first[223:216],
	       cache_cRqMshr$pipelineResp_getRq[43] ?
		 cache_cRqMshr$pipelineResp_getData[215:208] :
		 cache_pipeline$first[215:208] } ;
  assign IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3593 =
	     { IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3588,
	       cache_cRqMshr$pipelineResp_getRq[42] ?
		 cache_cRqMshr$pipelineResp_getData[207:200] :
		 cache_pipeline$first[207:200],
	       cache_cRqMshr$pipelineResp_getRq[41] ?
		 cache_cRqMshr$pipelineResp_getData[199:192] :
		 cache_pipeline$first[199:192] } ;
  assign IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3605 =
	     { IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2893,
	       cache_cRqMshr$pipelineResp_getRq[37] ?
		 cache_cRqMshr$pipelineResp_getData[167:160] :
		 cache_pipeline$first[167:160],
	       cache_cRqMshr$pipelineResp_getRq[36] ?
		 cache_cRqMshr$pipelineResp_getData[159:152] :
		 cache_pipeline$first[159:152] } ;
  assign IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3610 =
	     { IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3605,
	       cache_cRqMshr$pipelineResp_getRq[35] ?
		 cache_cRqMshr$pipelineResp_getData[151:144] :
		 cache_pipeline$first[151:144],
	       cache_cRqMshr$pipelineResp_getRq[34] ?
		 cache_cRqMshr$pipelineResp_getData[143:136] :
		 cache_pipeline$first[143:136] } ;
  assign IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3613 =
	     { IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3573,
	       IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3593,
	       IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3610,
	       cache_cRqMshr$pipelineResp_getRq[33] ?
		 cache_cRqMshr$pipelineResp_getData[135:128] :
		 cache_pipeline$first[135:128] } ;
  assign IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3628 =
	     { IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2934,
	       cache_cRqMshr$pipelineResp_getRq[28] ?
		 cache_cRqMshr$pipelineResp_getData[95:88] :
		 cache_pipeline$first[95:88],
	       cache_cRqMshr$pipelineResp_getRq[27] ?
		 cache_cRqMshr$pipelineResp_getData[87:80] :
		 cache_pipeline$first[87:80] } ;
  assign IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3633 =
	     { IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3628,
	       cache_cRqMshr$pipelineResp_getRq[26] ?
		 cache_cRqMshr$pipelineResp_getData[79:72] :
		 cache_pipeline$first[79:72],
	       cache_cRqMshr$pipelineResp_getRq[25] ?
		 cache_cRqMshr$pipelineResp_getData[71:64] :
		 cache_pipeline$first[71:64] } ;
  assign IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3648 =
	     { IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2968,
	       cache_cRqMshr$pipelineResp_getRq[21] ?
		 cache_cRqMshrpipelineResp_getData_BITS_63_TO_0__q78[39:32] :
		 cache_pipeline$first[39:32],
	       cache_cRqMshr$pipelineResp_getRq[20] ?
		 cache_cRqMshrpipelineResp_getData_BITS_63_TO_0__q78[31:24] :
		 cache_pipeline$first[31:24] } ;
  assign IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3653 =
	     { IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3648,
	       cache_cRqMshr$pipelineResp_getRq[19] ?
		 cache_cRqMshrpipelineResp_getData_BITS_63_TO_0__q78[23:16] :
		 cache_pipeline$first[23:16],
	       cache_cRqMshr$pipelineResp_getRq[18] ?
		 cache_cRqMshrpipelineResp_getData_BITS_63_TO_0__q78[15:8] :
		 cache_pipeline$first[15:8] } ;
  assign IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3656 =
	     { IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3613,
	       IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3633,
	       IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3653,
	       cache_cRqMshr$pipelineResp_getRq[17] ?
		 cache_cRqMshrpipelineResp_getData_BITS_63_TO_0__q78[7:0] :
		 cache_pipeline$first[7:0] } ;
  assign IF_cache_cRqMshr_pipelineResp_searchEndOfChain_ETC___d3012 =
	     (cache_cRqMshr$pipelineResp_searchEndOfChain[4] &&
	      cache_cRqMshr$pipelineResp_getState == 3'd1) ?
	       cache_pipeline$first[573:0] :
	       (cache_cRqMshr$pipelineResp_getRq[16] ?
		  IF_NOT_cache_pipeline_first__581_BITS_525_TO_5_ETC___d2999 :
		  IF_cache_pipeline_first__581_BITS_525_TO_524_6_ETC___d3010) ;
  assign IF_cache_cRqRetryIndexQ_deqReq_dummy2_2_read___ETC___d854 =
	     _theResult_____2__h234513 == v__h232953 ;
  assign IF_cache_cRqRetryIndexQ_deqReq_lat_1_whas__11__ETC___d817 =
	     WILL_FIRE_RL_cache_cRqTransfer_retry ||
	     cache_cRqRetryIndexQ_deqReq_rl ;
  assign IF_cache_cRqRetryIndexQ_enqReq_lat_1_whas__01__ETC___d833 =
	     cache_cRqRetryIndexQ_enqReq_lat_0$whas ?
	       cache_cRqRetryIndexQ_enqReq_lat_0$wget[4] :
	       cache_cRqRetryIndexQ_enqReq_rl[4] ;
  assign IF_cache_doLdAfterReplace_007_THEN_2_CONCAT_DO_ETC___d2016 =
	     cache_doLdAfterReplace ?
	       { 573'h12AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA,
		 cache_cRqMshr$sendToM_getRq[151:88],
		 1'd1,
		 cache_toMInfoQ$D_OUT[5:2] } :
	       { 2'd3,
		 addr__h288271,
		 64'hFFFFFFFFFFFFFFFF,
		 cache_cRqMshr$sendToM_getData[511:0] } ;
  assign IF_cache_pipeline_RDY_first__579_AND_cache_cRq_ETC___d2613 =
	     (cache_pipeline$RDY_first &&
	      cache_cRqMshr$pipelineResp_getRq[85:84] == 2'd3) ?
	       cache_rsStToDmaIndexQ_pipelineResp$FULL_N :
	       cache_rsLdToDmaIndexQ_pipelineResp$FULL_N ;
  assign IF_cache_pipeline_first__581_BITS_519_TO_518_5_ETC___d2676 =
	     (cache_pipeline_first__581_BITS_519_TO_518_594__ETC___d2598 &&
	      cache_pipeline_first__581_BITS_521_TO_520_600__ETC___d2601 &&
	      cache_pipeline_first__581_BITS_523_TO_522_603__ETC___d2604) ?
	       cache_cRqMshr$pipelineResp_getAddrSucc :
	       5'd10 ;
  assign IF_cache_pipeline_first__581_BITS_519_TO_518_5_ETC___d2693 =
	     (cache_pipeline_first__581_BITS_519_TO_518_594__ETC___d2598 &&
	      cache_pipeline_first__581_BITS_521_TO_520_600__ETC___d2601 &&
	      cache_pipeline_first__581_BITS_523_TO_522_603__ETC___d2604) ?
	       { IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2686,
		 cache_pipeline$first[523:518],
		 cache_cRqMshr$pipelineResp_getAddrSucc,
		 1'd0 } :
	       { cache_pipeline$first[525:518],
		 1'd1,
		 cache_pipeline$first[582:579],
		 1'd0 } ;
  assign IF_cache_pipeline_first__581_BITS_519_TO_518_5_ETC___d2993 =
	     (cache_pipeline_first__581_BITS_519_TO_518_594__ETC___d2598 &&
	      cache_pipeline_first__581_BITS_521_TO_520_600__ETC___d2601 &&
	      cache_pipeline_first__581_BITS_523_TO_522_603__ETC___d2604) ?
	       IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2991 :
	       cache_pipeline$first[511:0] ;
  assign IF_cache_pipeline_first__581_BITS_519_TO_518_5_ETC___d3025 =
	     (cache_pipeline_first__581_BITS_519_TO_518_594__ETC___d2598 &&
	      cache_pipeline_first__581_BITS_521_TO_520_600__ETC___d2601 &&
	      cache_pipeline_first__581_BITS_523_TO_522_603__ETC___d2604) ?
	       3'd4 :
	       3'd3 ;
  assign IF_cache_pipeline_first__581_BITS_523_TO_522_6_ETC___d3041 =
	     { cache_pipeline_first__581_BITS_523_TO_522_603__ETC___d2604 ?
		 4'd2 :
		 { 2'd1,
		   IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2597 },
	       cache_pipeline_first__581_BITS_521_TO_520_600__ETC___d2601 ?
		 4'd2 :
		 { 2'd1,
		   IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2597 } } ;
  assign IF_cache_pipeline_first__581_BITS_525_TO_524_6_ETC___d2667 =
	     (cache_pipeline$first[525:524] == 2'd0 ||
	      cache_pipeline_first__581_BITS_573_TO_526_644__ETC___d2646) ?
	       IF_NOT_cache_pipeline_first__581_BITS_525_TO_5_ETC___d2657 :
	       cache_pipeline$first[519:518] != 2'd0 ||
	       cache_pipeline$first[521:520] != 2'd0 ||
	       cache_pipeline$first[523:522] != 2'd0 ||
	       cache_toMInfoQ$FULL_N ;
  assign IF_cache_pipeline_first__581_BITS_525_TO_524_6_ETC___d2682 =
	     (cache_pipeline$first[525:524] == 2'd0 ||
	      cache_pipeline_first__581_BITS_573_TO_526_644__ETC___d2646) ?
	       ((cache_pipeline$first[525:524] != 2'd0 &&
		 IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2627) ?
		  cache_cRqMshr$pipelineResp_getAddrSucc :
		  5'd10) :
	       5'd10 ;
  assign IF_cache_pipeline_first__581_BITS_525_TO_524_6_ETC___d3010 =
	     (cache_pipeline$first[525:524] == 2'd0 ||
	      cache_pipeline_first__581_BITS_573_TO_526_644__ETC___d2646) ?
	       { cache_cRqMshr$pipelineResp_getRq[151:104],
		 IF_NOT_cache_pipeline_first__581_BITS_525_TO_5_ETC___d3000,
		 cache_pipeline$first[511:0] } :
	       ((cache_pipeline$first[519:518] == 2'd0 &&
		 cache_pipeline$first[521:520] == 2'd0 &&
		 cache_pipeline$first[523:522] == 2'd0) ?
		  { cache_cRqMshr$pipelineResp_getRq[151:104],
		    9'd1,
		    cache_pipeline$first[582:579],
		    513'h0AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA } :
		  { cache_pipeline$first[573:518],
		    1'd1,
		    cache_pipeline$first[582:579],
		    1'd1,
		    cache_pipeline$first[511:0] }) ;
  assign IF_cache_pipeline_first__581_BITS_525_TO_524_6_ETC___d3032 =
	     (cache_pipeline$first[525:524] == 2'd0 ||
	      cache_pipeline_first__581_BITS_573_TO_526_644__ETC___d2646) ?
	       ((cache_pipeline$first[525:524] != 2'd0 &&
		 IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2627) ?
		  3'd4 :
		  3'd3) :
	       ((cache_pipeline$first[519:518] == 2'd0 &&
		 cache_pipeline$first[521:520] == 2'd0 &&
		 cache_pipeline$first[523:522] == 2'd0) ?
		  3'd3 :
		  3'd2) ;
  assign IF_cache_pipeline_first__581_BITS_525_TO_524_6_ETC___d3095 =
	     (cache_pipeline$first[525:524] == 2'd0 ||
	      cache_pipeline_first__581_BITS_573_TO_526_644__ETC___d2646) ?
	       { cache_pipeline$first[578:575],
		 48'hAAAAAAAAAAAA,
		 cache_pipeline$first[525:524] == 2'd0,
		 IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3048,
		 IF_NOT_cache_cRqMshr_pipelineResp_getRq_IF_cac_ETC___d3054,
		 IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3057,
		 IF_NOT_cache_cRqMshr_pipelineResp_getRq_IF_cac_ETC___d3063,
		 IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3067,
		 IF_NOT_cache_cRqMshr_pipelineResp_getRq_IF_cac_ETC___d3073 } :
	       { cache_pipeline$first[578:575],
		 cache_pipeline$first[573:526],
		 cache_pipeline$first[519:518] == 2'd0 &&
		 cache_pipeline$first[521:520] == 2'd0 &&
		 cache_pipeline$first[523:522] == 2'd0,
		 (cache_pipeline$first[519:518] == 2'd0 &&
		  cache_pipeline$first[521:520] == 2'd0 &&
		  cache_pipeline$first[523:522] == 2'd0) ?
		   12'd546 :
		   { (cache_pipeline$first[523:522] == 2'd0) ?
		       cache_pipeline$first[523:520] :
		       4'd4,
		     (cache_pipeline$first[521:520] == 2'd0) ?
		       cache_pipeline$first[521:518] :
		       4'd4,
		     (cache_pipeline$first[519:518] == 2'd0) ?
		       cache_pipeline$first[519:516] :
		       4'd4 } } ;
  assign IF_cache_pipeline_first__581_BITS_525_TO_524_6_ETC___d3171 =
	     (cache_pipeline$first[525:524] == 2'd3) ? 2'd2 : 2'd0 ;
  assign IF_cache_pipeline_first__581_BIT_512_308_THEN__ETC___d3486 =
	     cache_pipeline$first[512] ?
	       5'd10 :
	       (IF_SEL_ARR_cache_cRqMshr_pipelineResp_getSlot__ETC___d3484 ?
		  cache_cRqMshr$pipelineResp_getAddrSucc :
		  5'd10) ;
  assign IF_cache_pipeline_first__581_BIT_512_308_THEN__ETC___d3660 =
	     cache_pipeline$first[512] ?
	       (IF_SEL_ARR_cache_pipeline_first__581_BITS_519__ETC___d3488 ?
		  { cache_cRqMshr$pipelineResp_getRq[151:104],
		    9'd1,
		    cache_pipeline$first[516:513],
		    513'h0AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA } :
		  cache_pipeline$first[573:0]) :
	       (IF_SEL_ARR_cache_cRqMshr_pipelineResp_getSlot__ETC___d3484 ?
		  cache_cRqMshr_pipelineResp_getRq_IF_cache_pipe_ETC___d3658 :
		  cache_pipeline$first[573:0]) ;
  assign IF_cache_pipeline_first__581_BIT_517_582_THEN__ETC___d3124 =
	     cache_pipeline$first[517] ?
	       cache_cRqMshr$pipelineResp_getRq[16] ||
	       CASE_cache_cRqMshrpipelineResp_getRq_BITS_82__ETC__q79 ==
	       2'd0 :
	       cache_cRqMshr_pipelineResp_getRq_IF_cache_pipe_ETC___d3123 ;
  assign IF_cache_rqFromCQ_deqReq_dummy2_2_read__7_AND__ETC___d55 =
	     _theResult_____2__h7215 == v__h6037 ;
  assign IF_cache_rqFromCQ_deqReq_lat_1_whas__3_THEN_ca_ETC___d19 =
	     WILL_FIRE_RL_cache_cRqTransfer_new_child ||
	     cache_rqFromCQ_deqReq_rl ;
  assign IF_cache_rqFromCQ_enqReq_lat_1_whas_THEN_cache_ETC___d39 =
	     EN_to_child_rqFromC_enq ?
	       cache_rqFromCQ_enqReq_lat_0$wget[74] :
	       cache_rqFromCQ_enqReq_rl[74] ;
  assign IF_cache_rqFromDmaQ_deqReq_dummy2_2_read__53_A_ETC___d361 =
	     _theResult_____2__h119142 == v__h72082 ;
  assign IF_cache_rqFromDmaQ_deqReq_lat_1_whas__19_THEN_ETC___d325 =
	     WILL_FIRE_RL_cache_cRqTransfer_new_dma ||
	     cache_rqFromDmaQ_deqReq_rl ;
  assign IF_cache_rqFromDmaQ_enqReq_lat_1_whas__09_THEN_ETC___d345 =
	     EN_dma_memReq_enq ?
	       cache_rqFromDmaQ_enqReq_lat_0$wget[656] :
	       cache_rqFromDmaQ_enqReq_rl[656] ;
  assign IF_cache_rsFromCQ_deqReq_dummy2_2_read__39_AND_ETC___d147 =
	     _theResult_____2__h22297 == v__h16641 ;
  assign IF_cache_rsFromCQ_deqReq_lat_1_whas__05_THEN_c_ETC___d111 =
	     WILL_FIRE_RL_cache_cRsTransfer || cache_rsFromCQ_deqReq_rl ;
  assign IF_cache_rsFromCQ_enqReq_lat_1_whas__5_THEN_ca_ETC___d131 =
	     EN_to_child_rsFromC_enq ?
	       cache_rsFromCQ_enqReq_lat_0$wget[581] :
	       cache_rsFromCQ_enqReq_rl[581] ;
  assign IF_cache_rsFromMQ_deqReq_dummy2_2_read__54_AND_ETC___d762 =
	     _theResult_____2__h225016 == v__h218716 ;
  assign IF_cache_rsFromMQ_deqReq_lat_1_whas__20_THEN_c_ETC___d726 =
	     cache_rsFromMQ_deqReq_lat_0$whas || cache_rsFromMQ_deqReq_rl ;
  assign IF_cache_rsFromMQ_enqReq_lat_1_whas__10_THEN_c_ETC___d746 =
	     EN_to_mem_rsFromM_enq ?
	       cache_rsFromMQ_enqReq_lat_0$wget[517] :
	       cache_rsFromMQ_enqReq_rl[517] ;
  assign IF_cache_rsLdToDmaQ_deqReq_dummy2_2_read__44_A_ETC___d452 =
	     _theResult_____2__h135235 == v__h129259 ;
  assign IF_cache_rsLdToDmaQ_deqReq_lat_1_whas__10_THEN_ETC___d416 =
	     EN_dma_respLd_deq || cache_rsLdToDmaQ_deqReq_rl ;
  assign IF_cache_rsLdToDmaQ_enqReq_lat_1_whas__00_THEN_ETC___d436 =
	     CAN_FIRE_RL_cache_sendRsLdToDma ?
	       cache_rsLdToDmaQ_enqReq_lat_0$wget[528] :
	       cache_rsLdToDmaQ_enqReq_rl[528] ;
  assign IF_cache_rsStToDmaQ_deqReq_dummy2_2_read__35_A_ETC___d543 =
	     _theResult_____2__h142737 == v__h142239 ;
  assign IF_cache_rsStToDmaQ_deqReq_lat_1_whas__01_THEN_ETC___d507 =
	     EN_dma_respSt_deq || cache_rsStToDmaQ_deqReq_rl ;
  assign IF_cache_rsStToDmaQ_enqReq_lat_1_whas__91_THEN_ETC___d527 =
	     WILL_FIRE_RL_cache_sendRsStToDma ?
	       cache_rsStToDmaQ_enqReq_lat_0$wget[16] :
	       cache_rsStToDmaQ_enqReq_rl[16] ;
  assign IF_cache_rsToCIndexQ_deqReq_dummy2_2_read__64__ETC___d977 =
	     _theResult_____2__h245988 == v__h242396 ;
  assign IF_cache_rsToCIndexQ_deqReq_lat_1_whas__34_THE_ETC___d940 =
	     WILL_FIRE_RL_cache_sendRsToC || cache_rsToCIndexQ_deqReq_rl ;
  assign IF_cache_rsToCIndexQ_enqReq_lat_1_whas__24_THE_ETC___d956 =
	     cache_rsToCIndexQ_enqReq_lat_0$whas ?
	       cache_rsToCIndexQ_enqReq_lat_0$wget[6] :
	       cache_rsToCIndexQ_enqReq_rl[6] ;
  assign IF_cache_toCQ_deqReq_dummy2_2_read__61_AND_IF__ETC___d269 =
	     _theResult_____2__h37990 == v__h31944 ;
  assign IF_cache_toCQ_deqReq_lat_1_whas__32_THEN_cache_ETC___d238 =
	     EN_to_child_toC_deq || cache_toCQ_deqReq_rl ;
  assign IF_cache_toCQ_enqReq_dummy2_2_read__53_AND_IF__ETC___d302 =
	     (cache_toCQ_enqReq_dummy2_2$Q_OUT &&
	      IF_cache_toCQ_enqReq_lat_1_whas__87_THEN_cache_ETC___d196 &&
	      (cache_toCQ_enqReq_lat_0$whas ?
		 !cache_toCQ_enqReq_lat_0$wget[584] :
		 !cache_toCQ_enqReq_rl[584])) ?
	       { 516'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA,
		 cache_toCQ_enqReq_lat_0$whas ?
		   cache_toCQ_enqReq_lat_0$wget[67:0] :
		   cache_toCQ_enqReq_rl[67:0] } :
	       (cache_toCQ_enqReq_lat_0$whas ?
		  cache_toCQ_enqReq_lat_0$wget[583:0] :
		  cache_toCQ_enqReq_rl[583:0]) ;
  assign IF_cache_toCQ_enqReq_lat_1_whas__87_THEN_cache_ETC___d196 =
	     cache_toCQ_enqReq_lat_0$whas ?
	       cache_toCQ_enqReq_lat_0$wget[585] :
	       cache_toCQ_enqReq_rl[585] ;
  assign IF_cache_toMQ_deqReq_dummy2_2_read__62_AND_IF__ETC___d670 =
	     _theResult_____2__h208521 == v__h168573 ;
  assign IF_cache_toMQ_deqReq_lat_1_whas__33_THEN_cache_ETC___d639 =
	     EN_to_mem_toM_deq || cache_toMQ_deqReq_rl ;
  assign IF_cache_toMQ_enqReq_dummy2_2_read__54_AND_IF__ETC___d703 =
	     (cache_toMQ_enqReq_dummy2_2$Q_OUT &&
	      IF_cache_toMQ_enqReq_lat_1_whas__88_THEN_cache_ETC___d597 &&
	      (cache_toMQ_enqReq_lat_0$whas ?
		 !cache_toMQ_enqReq_lat_0$wget[640] :
		 !cache_toMQ_enqReq_rl[640])) ?
	       { 571'h2AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA,
		 cache_toMQ_enqReq_lat_0$whas ?
		   cache_toMQ_enqReq_lat_0$wget[68:0] :
		   cache_toMQ_enqReq_rl[68:0] } :
	       (cache_toMQ_enqReq_lat_0$whas ?
		  cache_toMQ_enqReq_lat_0$wget[639:0] :
		  cache_toMQ_enqReq_rl[639:0]) ;
  assign IF_cache_toMQ_enqReq_lat_1_whas__88_THEN_cache_ETC___d597 =
	     cache_toMQ_enqReq_lat_0$whas ?
	       cache_toMQ_enqReq_lat_0$wget[641] :
	       cache_toMQ_enqReq_rl[641] ;
  assign IF_perfReqQ_enqReq_lat_1_whas__839_THEN_perfRe_ETC___d3875 =
	     EN_perf_req ?
	       perfReqQ_enqReq_lat_0$wget[4] :
	       perfReqQ_enqReq_rl[4] ;
  assign NOT_IF_cache_pipeline_first__581_BITS_584_TO_5_ETC___d3191 =
	     cache_pipeline$first[582:579] != pipeOutCRqIdx__h314276 ;
  assign NOT_SEL_ARR_NOT_cache_rqFromDmaQ_data_0_129_BI_ETC___d1584 =
	     !CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q5 ||
	     !CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q6 ||
	     !CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q7 ;
  assign NOT_SEL_ARR_NOT_cache_rqFromDmaQ_data_0_129_BI_ETC___d1586 =
	     !CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q8 ||
	     !CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q9 ||
	     NOT_SEL_ARR_NOT_cache_rqFromDmaQ_data_0_129_BI_ETC___d1584 ;
  assign NOT_SEL_ARR_NOT_cache_rqFromDmaQ_data_0_129_BI_ETC___d1588 =
	     !CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q10 ||
	     !CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q11 ||
	     NOT_SEL_ARR_NOT_cache_rqFromDmaQ_data_0_129_BI_ETC___d1586 ;
  assign NOT_SEL_ARR_NOT_cache_rqFromDmaQ_data_0_129_BI_ETC___d1590 =
	     !CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q12 ||
	     !CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q13 ||
	     NOT_SEL_ARR_NOT_cache_rqFromDmaQ_data_0_129_BI_ETC___d1588 ;
  assign NOT_SEL_ARR_NOT_cache_rqFromDmaQ_data_0_129_BI_ETC___d1592 =
	     !CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q14 ||
	     !CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q15 ||
	     NOT_SEL_ARR_NOT_cache_rqFromDmaQ_data_0_129_BI_ETC___d1590 ;
  assign NOT_SEL_ARR_NOT_cache_rqFromDmaQ_data_0_129_BI_ETC___d1594 =
	     !CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q16 ||
	     !CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q17 ||
	     NOT_SEL_ARR_NOT_cache_rqFromDmaQ_data_0_129_BI_ETC___d1592 ;
  assign NOT_SEL_ARR_NOT_cache_rqFromDmaQ_data_0_129_BI_ETC___d1596 =
	     !CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q18 ||
	     !CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q19 ||
	     NOT_SEL_ARR_NOT_cache_rqFromDmaQ_data_0_129_BI_ETC___d1594 ;
  assign NOT_SEL_ARR_NOT_cache_rqFromDmaQ_data_0_129_BI_ETC___d1598 =
	     !CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q20 ||
	     !CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q21 ||
	     NOT_SEL_ARR_NOT_cache_rqFromDmaQ_data_0_129_BI_ETC___d1596 ;
  assign NOT_SEL_ARR_NOT_cache_rqFromDmaQ_data_0_129_BI_ETC___d1600 =
	     !CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q22 ||
	     !CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q23 ||
	     NOT_SEL_ARR_NOT_cache_rqFromDmaQ_data_0_129_BI_ETC___d1598 ;
  assign NOT_SEL_ARR_NOT_cache_rqFromDmaQ_data_0_129_BI_ETC___d1602 =
	     !CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q24 ||
	     !CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q25 ||
	     NOT_SEL_ARR_NOT_cache_rqFromDmaQ_data_0_129_BI_ETC___d1600 ;
  assign NOT_SEL_ARR_NOT_cache_rqFromDmaQ_data_0_129_BI_ETC___d1604 =
	     !CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q26 ||
	     !CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q27 ||
	     NOT_SEL_ARR_NOT_cache_rqFromDmaQ_data_0_129_BI_ETC___d1602 ;
  assign NOT_SEL_ARR_NOT_cache_rqFromDmaQ_data_0_129_BI_ETC___d1606 =
	     !CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q28 ||
	     !CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q29 ||
	     NOT_SEL_ARR_NOT_cache_rqFromDmaQ_data_0_129_BI_ETC___d1604 ;
  assign NOT_SEL_ARR_NOT_cache_rqFromDmaQ_data_0_129_BI_ETC___d1608 =
	     !CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q30 ||
	     !CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q31 ||
	     NOT_SEL_ARR_NOT_cache_rqFromDmaQ_data_0_129_BI_ETC___d1606 ;
  assign NOT_SEL_ARR_NOT_cache_rqFromDmaQ_data_0_129_BI_ETC___d1610 =
	     !CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q32 ||
	     !CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q33 ||
	     NOT_SEL_ARR_NOT_cache_rqFromDmaQ_data_0_129_BI_ETC___d1608 ;
  assign NOT_SEL_ARR_NOT_cache_rqFromDmaQ_data_0_129_BI_ETC___d1612 =
	     !CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q34 ||
	     !CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q35 ||
	     NOT_SEL_ARR_NOT_cache_rqFromDmaQ_data_0_129_BI_ETC___d1610 ;
  assign NOT_SEL_ARR_NOT_cache_rqFromDmaQ_data_0_129_BI_ETC___d1614 =
	     !CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q36 ||
	     !CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q37 ||
	     NOT_SEL_ARR_NOT_cache_rqFromDmaQ_data_0_129_BI_ETC___d1612 ;
  assign NOT_SEL_ARR_NOT_cache_rqFromDmaQ_data_0_129_BI_ETC___d1616 =
	     !CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q38 ||
	     !CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q39 ||
	     NOT_SEL_ARR_NOT_cache_rqFromDmaQ_data_0_129_BI_ETC___d1614 ;
  assign NOT_SEL_ARR_NOT_cache_rqFromDmaQ_data_0_129_BI_ETC___d1618 =
	     !CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q40 ||
	     !CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q41 ||
	     NOT_SEL_ARR_NOT_cache_rqFromDmaQ_data_0_129_BI_ETC___d1616 ;
  assign NOT_SEL_ARR_NOT_cache_rqFromDmaQ_data_0_129_BI_ETC___d1620 =
	     !CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q42 ||
	     !CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q43 ||
	     NOT_SEL_ARR_NOT_cache_rqFromDmaQ_data_0_129_BI_ETC___d1618 ;
  assign NOT_SEL_ARR_NOT_cache_rqFromDmaQ_data_0_129_BI_ETC___d1622 =
	     !CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q44 ||
	     !CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q45 ||
	     NOT_SEL_ARR_NOT_cache_rqFromDmaQ_data_0_129_BI_ETC___d1620 ;
  assign NOT_SEL_ARR_NOT_cache_rqFromDmaQ_data_0_129_BI_ETC___d1624 =
	     !CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q46 ||
	     !CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q47 ||
	     NOT_SEL_ARR_NOT_cache_rqFromDmaQ_data_0_129_BI_ETC___d1622 ;
  assign NOT_SEL_ARR_NOT_cache_rqFromDmaQ_data_0_129_BI_ETC___d1626 =
	     !CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q48 ||
	     !CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q49 ||
	     NOT_SEL_ARR_NOT_cache_rqFromDmaQ_data_0_129_BI_ETC___d1624 ;
  assign NOT_SEL_ARR_NOT_cache_rqFromDmaQ_data_0_129_BI_ETC___d1628 =
	     !CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q50 ||
	     !CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q51 ||
	     NOT_SEL_ARR_NOT_cache_rqFromDmaQ_data_0_129_BI_ETC___d1626 ;
  assign NOT_SEL_ARR_NOT_cache_rqFromDmaQ_data_0_129_BI_ETC___d1630 =
	     !CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q52 ||
	     !CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q53 ||
	     NOT_SEL_ARR_NOT_cache_rqFromDmaQ_data_0_129_BI_ETC___d1628 ;
  assign NOT_SEL_ARR_NOT_cache_rqFromDmaQ_data_0_129_BI_ETC___d1632 =
	     !CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q54 ||
	     !CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q55 ||
	     NOT_SEL_ARR_NOT_cache_rqFromDmaQ_data_0_129_BI_ETC___d1630 ;
  assign NOT_SEL_ARR_NOT_cache_rqFromDmaQ_data_0_129_BI_ETC___d1634 =
	     !CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q56 ||
	     !CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q57 ||
	     NOT_SEL_ARR_NOT_cache_rqFromDmaQ_data_0_129_BI_ETC___d1632 ;
  assign NOT_SEL_ARR_NOT_cache_rqFromDmaQ_data_0_129_BI_ETC___d1636 =
	     !CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q58 ||
	     !CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q59 ||
	     NOT_SEL_ARR_NOT_cache_rqFromDmaQ_data_0_129_BI_ETC___d1634 ;
  assign NOT_SEL_ARR_NOT_cache_rqFromDmaQ_data_0_129_BI_ETC___d1638 =
	     !CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q60 ||
	     !CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q61 ||
	     NOT_SEL_ARR_NOT_cache_rqFromDmaQ_data_0_129_BI_ETC___d1636 ;
  assign NOT_SEL_ARR_NOT_cache_rqFromDmaQ_data_0_129_BI_ETC___d1640 =
	     !CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q62 ||
	     !CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q63 ||
	     NOT_SEL_ARR_NOT_cache_rqFromDmaQ_data_0_129_BI_ETC___d1638 ;
  assign NOT_SEL_ARR_NOT_cache_rqFromDmaQ_data_0_129_BI_ETC___d1642 =
	     !CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q64 ||
	     !CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q65 ||
	     NOT_SEL_ARR_NOT_cache_rqFromDmaQ_data_0_129_BI_ETC___d1640 ;
  assign NOT_SEL_ARR_NOT_cache_rqFromDmaQ_data_0_129_BI_ETC___d1644 =
	     !CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q66 ||
	     !CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q67 ||
	     NOT_SEL_ARR_NOT_cache_rqFromDmaQ_data_0_129_BI_ETC___d1642 ;
  assign NOT_SEL_ARR_cache_cRqMshr_sendRqToC_getSlot_IF_ETC___d2508 =
	     !CASE_child13067_0_cache_cRqMshrsendRqToC_getS_ETC__q254 ;
  assign NOT_cache_cRqMshr_pipelineResp_getRq_IF_cache__ETC___d3264 =
	     (cache_cRqMshr$pipelineResp_getRq[17] ||
	      cache_cRqMshr$pipelineResp_getRq[18] ||
	      cache_cRqMshr$pipelineResp_getRq[19] ||
	      cache_cRqMshr$pipelineResp_getRq[20] ||
	      cache_cRqMshr$pipelineResp_getRq[21] ||
	      cache_cRqMshr$pipelineResp_getRq[22] ||
	      cache_cRqMshr$pipelineResp_getRq[23] ||
	      cache_cRqMshr$pipelineResp_getRq[24] ||
	      cache_cRqMshr$pipelineResp_getRq[25] ||
	      cache_cRqMshr$pipelineResp_getRq[26] ||
	      cache_cRqMshr$pipelineResp_getRq[27] ||
	      cache_cRqMshr$pipelineResp_getRq[28] ||
	      cache_cRqMshr$pipelineResp_getRq[29] ||
	      cache_cRqMshr$pipelineResp_getRq[30] ||
	      cache_cRqMshr$pipelineResp_getRq[31] ||
	      cache_cRqMshr$pipelineResp_getRq[32] ||
	      cache_cRqMshr$pipelineResp_getRq[33] ||
	      cache_cRqMshr$pipelineResp_getRq[34] ||
	      cache_cRqMshr$pipelineResp_getRq[35] ||
	      cache_cRqMshr$pipelineResp_getRq[36] ||
	      cache_cRqMshr$pipelineResp_getRq[37] ||
	      cache_cRqMshr$pipelineResp_getRq[38] ||
	      cache_cRqMshr$pipelineResp_getRq[39] ||
	      cache_cRqMshr$pipelineResp_getRq[40] ||
	      cache_cRqMshr$pipelineResp_getRq[41] ||
	      cache_cRqMshr$pipelineResp_getRq[42] ||
	      cache_cRqMshr$pipelineResp_getRq[43] ||
	      cache_cRqMshr$pipelineResp_getRq[44] ||
	      cache_cRqMshr$pipelineResp_getRq[45] ||
	      cache_cRqMshr$pipelineResp_getRq[46] ||
	      cache_cRqMshr$pipelineResp_getRq[47] ||
	      cache_cRqMshr$pipelineResp_getRq[48] ||
	      cache_cRqMshr$pipelineResp_getRq[49] ||
	      cache_cRqMshr$pipelineResp_getRq[50] ||
	      cache_cRqMshr$pipelineResp_getRq[51] ||
	      cache_cRqMshr$pipelineResp_getRq[52] ||
	      cache_cRqMshr$pipelineResp_getRq[53] ||
	      cache_cRqMshr$pipelineResp_getRq[54] ||
	      cache_cRqMshr$pipelineResp_getRq[55] ||
	      cache_cRqMshr$pipelineResp_getRq[56] ||
	      cache_cRqMshr$pipelineResp_getRq[57] ||
	      cache_cRqMshr$pipelineResp_getRq[58] ||
	      cache_cRqMshr$pipelineResp_getRq[59] ||
	      cache_cRqMshr$pipelineResp_getRq[60] ||
	      cache_cRqMshr$pipelineResp_getRq[61] ||
	      cache_cRqMshr$pipelineResp_getRq[62] ||
	      cache_cRqMshr$pipelineResp_getRq[63] ||
	      cache_cRqMshr$pipelineResp_getRq[64] ||
	      cache_cRqMshr$pipelineResp_getRq[65] ||
	      cache_cRqMshr$pipelineResp_getRq[66] ||
	      cache_cRqMshr$pipelineResp_getRq[67] ||
	      cache_cRqMshr$pipelineResp_getRq[68] ||
	      cache_cRqMshr$pipelineResp_getRq[69] ||
	      cache_cRqMshr$pipelineResp_getRq[70] ||
	      cache_cRqMshr$pipelineResp_getRq[71] ||
	      cache_cRqMshr$pipelineResp_getRq[72] ||
	      cache_cRqMshr$pipelineResp_getRq[73] ||
	      cache_cRqMshr$pipelineResp_getRq[74] ||
	      cache_cRqMshr$pipelineResp_getRq[75] ||
	      cache_cRqMshr$pipelineResp_getRq[76] ||
	      cache_cRqMshr$pipelineResp_getRq[77] ||
	      cache_cRqMshr$pipelineResp_getRq[78] ||
	      cache_cRqMshr$pipelineResp_getRq[79] ||
	      cache_cRqMshr$pipelineResp_getRq[80]) !=
	     (cache_cRqMshr$pipelineResp_getRq[85:84] == 2'd3) ;
  assign NOT_cache_cRqMshr_pipelineResp_getRq_IF_cache__ETC___d3290 =
	     !cache_cRqMshr$pipelineResp_getRq[16] &&
	     IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2627 &&
	     (!cache_pipeline_first__581_BITS_573_TO_526_644__ETC___d2646 ||
	      cache_pipeline$first[525:524] == 2'd0) ;
  assign NOT_cache_cRqMshr_pipelineResp_getRq_IF_cache__ETC___d3299 =
	     !cache_cRqMshr$pipelineResp_getRq[16] &&
	     IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3156 &&
	     cache_pipeline$first[525:524] == 2'd0 &&
	     (cache_pipeline$first[519:518] != 2'd0 ||
	      cache_pipeline$first[521:520] != 2'd0 ||
	      cache_pipeline$first[523:522] != 2'd0) ;
  assign NOT_cache_cRqMshr_pipelineResp_getSlot_IF_cach_ETC___d3369 =
	     cache_cRqMshr$pipelineResp_getSlot[64:61] !=
	     cache_pipeline$first[578:575] ;
  assign NOT_cache_cRqMshr_pipelineResp_searchEndOfChai_ETC___d3114 =
	     (!cache_cRqMshr$pipelineResp_searchEndOfChain[4] ||
	      cache_cRqMshr$pipelineResp_getState != 3'd1) &&
	     (cache_cRqMshr$pipelineResp_getRq[16] &&
	      NOT_cache_pipeline_first__581_BITS_525_TO_524__ETC___d3019 ||
	      !cache_cRqMshr$pipelineResp_getRq[16] &&
	      (cache_pipeline_first__581_BITS_573_TO_526_644__ETC___d2646 &&
	       cache_pipeline$first[525:524] != 2'd0 &&
	       IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2627 ||
	       cache_pipeline$first[525:524] != 2'd0 &&
	       !cache_pipeline_first__581_BITS_573_TO_526_644__ETC___d2646 &&
	       cache_pipeline$first[519:518] == 2'd0 &&
	       cache_pipeline$first[521:520] == 2'd0 &&
	       cache_pipeline$first[523:522] == 2'd0)) ;
  assign NOT_cache_cRqMshr_pipelineResp_searchEndOfChai_ETC___d3353 =
	     (!cache_cRqMshr$pipelineResp_searchEndOfChain[4] ||
	      cache_cRqMshr$pipelineResp_getState != 3'd1) &&
	     !cache_cRqMshr$pipelineResp_getRq[16] &&
	     cache_pipeline$first[525:524] == 2'd0 &&
	     (cache_pipeline$first[519:518] != 2'd0 ||
	      cache_pipeline$first[521:520] != 2'd0 ||
	      cache_pipeline$first[523:522] != 2'd0) ;
  assign NOT_cache_cRqRetryIndexQ_clearReq_dummy2_1_rea_ETC___d853 =
	     !cache_cRqRetryIndexQ_clearReq_dummy2_1$Q_OUT ||
	     !cache_cRqRetryIndexQ_clearReq_rl ;
  assign NOT_cache_cRqRetryIndexQ_enqReq_dummy2_2_read__ETC___d876 =
	     (!cache_cRqRetryIndexQ_enqReq_dummy2_2$Q_OUT ||
	      (cache_cRqRetryIndexQ_enqReq_lat_0$whas ?
		 !cache_cRqRetryIndexQ_enqReq_lat_0$wget[4] :
		 !cache_cRqRetryIndexQ_enqReq_rl[4])) &&
	     (cache_cRqRetryIndexQ_deqReq_dummy2_2$Q_OUT &&
	      IF_cache_cRqRetryIndexQ_deqReq_lat_1_whas__11__ETC___d817 ||
	      cache_cRqRetryIndexQ_empty) ;
  assign NOT_cache_pipeline_first__581_BITS_516_TO_513__ETC___d2637 =
	     !cache_pipeline_first__581_BITS_516_TO_513_583__ETC___d2588 ||
	     (cache_cRqMshr$pipelineResp_getRq[16] ?
		_0_OR_NOT_cache_pipeline_first__581_BITS_519_TO_ETC___d2614 :
		IF_IF_cache_cRqMshr_pipelineResp_getRq_IF_cach_ETC___d2635) ;
  assign NOT_cache_pipeline_first__581_BITS_516_TO_513__ETC___d3798 =
	     cache_pipeline$first[516:513] != pipeOutCRqIdx__h314276 ;
  assign NOT_cache_pipeline_first__581_BITS_519_TO_518__ETC___d3275 =
	     (!cache_pipeline_first__581_BITS_519_TO_518_594__ETC___d2598 ||
	      !cache_pipeline_first__581_BITS_521_TO_520_600__ETC___d2601 ||
	      !cache_pipeline_first__581_BITS_523_TO_522_603__ETC___d2604) &&
	     (!cache_pipeline_first__581_BITS_573_TO_526_644__ETC___d2646 ||
	      cache_pipeline$first[525:524] == 2'd0) ;
  assign NOT_cache_pipeline_first__581_BITS_519_TO_518__ETC___d3281 =
	     (!cache_pipeline_first__581_BITS_519_TO_518_594__ETC___d2598 ||
	      !cache_pipeline_first__581_BITS_521_TO_520_600__ETC___d2601 ||
	      !cache_pipeline_first__581_BITS_523_TO_522_603__ETC___d2604) &&
	     cache_cRqMshr$pipelineResp_getSlot[12] ;
  assign NOT_cache_pipeline_first__581_BITS_525_TO_524__ETC___d3019 =
	     cache_pipeline$first[525:524] != 2'd0 &&
	     cache_pipeline_first__581_BITS_573_TO_526_644__ETC___d2646 &&
	     cache_pipeline_first__581_BITS_519_TO_518_594__ETC___d2598 &&
	     cache_pipeline_first__581_BITS_521_TO_520_600__ETC___d2601 &&
	     cache_pipeline_first__581_BITS_523_TO_522_603__ETC___d2604 ;
  assign NOT_cache_pipeline_first__581_BIT_512_308_309__ETC___d3801 =
	     !cache_pipeline$first[512] &&
	     IF_SEL_ARR_cache_cRqMshr_pipelineResp_getSlot__ETC___d3484 &&
	     cache_cRqMshr$pipelineResp_getRq[16] &&
	     NOT_cache_pipeline_first__581_BITS_516_TO_513__ETC___d3798 ;
  assign NOT_cache_pipeline_first__581_BIT_512_308_309__ETC___d3809 =
	     !cache_pipeline$first[512] &&
	     IF_SEL_ARR_cache_cRqMshr_pipelineResp_getSlot__ETC___d3484 &&
	     cache_cRqMshr$pipelineResp_getRq[16] &&
	     NOT_cache_cRqMshr_pipelineResp_getRq_IF_cache__ETC___d3264 ;
  assign NOT_cache_pipeline_first__581_BIT_512_308_309__ETC___d3827 =
	     !cache_pipeline$first[512] &&
	     IF_SEL_ARR_cache_cRqMshr_pipelineResp_getSlot__ETC___d3484 &&
	     !cache_cRqMshr$pipelineResp_getRq[16] &&
	     NOT_cache_pipeline_first__581_BITS_516_TO_513__ETC___d3798 ;
  assign NOT_cache_pipeline_first__581_BIT_517_582_105__ETC___d3133 =
	     !cache_pipeline$first[517] &&
	     (!cache_cRqMshr$pipelineResp_searchEndOfChain[4] ||
	      cache_cRqMshr$pipelineResp_getState != 3'd1) &&
	     cache_cRqMshr$pipelineResp_getRq[16] &&
	     cache_pipeline$first[525:524] != 2'd0 &&
	     cache_pipeline_first__581_BITS_573_TO_526_644__ETC___d2646 &&
	     cache_pipeline_first__581_BITS_519_TO_518_594__ETC___d3126 ;
  assign NOT_cache_pipeline_first__581_BIT_517_582_105__ETC___d3143 =
	     !cache_pipeline$first[517] &&
	     (!cache_cRqMshr$pipelineResp_searchEndOfChain[4] ||
	      cache_cRqMshr$pipelineResp_getState != 3'd1) &&
	     cache_cRqMshr$pipelineResp_getRq[16] &&
	     cache_pipeline$first[525:524] != 2'd0 &&
	     cache_pipeline_first__581_BITS_573_TO_526_644__ETC___d2646 &&
	     cache_pipeline_first__581_BITS_519_TO_518_594__ETC___d3136 ;
  assign NOT_cache_pipeline_first__581_BIT_517_582_105__ETC___d3149 =
	     !cache_pipeline$first[517] &&
	     (!cache_cRqMshr$pipelineResp_searchEndOfChain[4] ||
	      cache_cRqMshr$pipelineResp_getState != 3'd1) &&
	     !cache_cRqMshr$pipelineResp_getRq[16] &&
	     cache_pipeline_first__581_BITS_573_TO_526_644__ETC___d2646 &&
	     cache_pipeline$first[525:524] != 2'd0 &&
	     IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2627 ;
  assign NOT_cache_pipeline_first__581_BIT_517_582_105__ETC___d3316 =
	     !cache_pipeline$first[517] &&
	     (!cache_cRqMshr$pipelineResp_searchEndOfChain[4] ||
	      cache_cRqMshr$pipelineResp_getState != 3'd1) &&
	     cache_cRqMshr$pipelineResp_getRq[16] &&
	     cache_pipeline$first[525:524] != 2'd0 &&
	     cache_pipeline_first__581_BITS_573_TO_526_644__ETC___d2646 &&
	     cache_pipeline_first__581_BITS_519_TO_518_594__ETC___d3192 ;
  assign NOT_cache_pipeline_first__581_BIT_517_582_105__ETC___d3320 =
	     !cache_pipeline$first[517] &&
	     (!cache_cRqMshr$pipelineResp_searchEndOfChain[4] ||
	      cache_cRqMshr$pipelineResp_getState != 3'd1) &&
	     cache_cRqMshr$pipelineResp_getRq[16] &&
	     cache_pipeline$first[525:524] != 2'd0 &&
	     cache_pipeline_first__581_BITS_573_TO_526_644__ETC___d2646 &&
	     cache_pipeline_first__581_BITS_519_TO_518_594__ETC___d3265 ;
  assign NOT_cache_pipeline_first__581_BIT_517_582_105__ETC___d3324 =
	     !cache_pipeline$first[517] &&
	     (!cache_cRqMshr$pipelineResp_searchEndOfChain[4] ||
	      cache_cRqMshr$pipelineResp_getState != 3'd1) &&
	     cache_cRqMshr$pipelineResp_getRq[16] &&
	     cache_pipeline$first[525:524] != 2'd0 &&
	     cache_pipeline_first__581_BITS_573_TO_526_644__ETC___d2646 &&
	     cache_pipeline_first__581_BITS_519_TO_518_594__ETC___d3271 ;
  assign NOT_cache_pipeline_first__581_BIT_517_582_105__ETC___d3328 =
	     !cache_pipeline$first[517] &&
	     (!cache_cRqMshr$pipelineResp_searchEndOfChain[4] ||
	      cache_cRqMshr$pipelineResp_getState != 3'd1) &&
	     cache_cRqMshr$pipelineResp_getRq[16] &&
	     cache_pipeline$first[525:524] != 2'd0 &&
	     cache_pipeline_first__581_BITS_573_TO_526_644__ETC___d2646 &&
	     NOT_cache_pipeline_first__581_BITS_519_TO_518__ETC___d3281 ;
  assign NOT_cache_pipeline_first__581_BIT_517_582_105__ETC___d3332 =
	     !cache_pipeline$first[517] &&
	     (!cache_cRqMshr$pipelineResp_searchEndOfChain[4] ||
	      cache_cRqMshr$pipelineResp_getState != 3'd1) &&
	     cache_cRqMshr$pipelineResp_getRq[16] &&
	     (cache_pipeline$first[525:524] == 2'd0 ||
	      !cache_pipeline_first__581_BITS_573_TO_526_644__ETC___d2646) &&
	     cache_cRqMshr$pipelineResp_getAddrSucc[4] ;
  assign NOT_cache_pipeline_first__581_BIT_517_582_105__ETC___d3340 =
	     !cache_pipeline$first[517] &&
	     (!cache_cRqMshr$pipelineResp_searchEndOfChain[4] ||
	      cache_cRqMshr$pipelineResp_getState != 3'd1) &&
	     cache_cRqMshr$pipelineResp_getRq[16] &&
	     (cache_pipeline$first[525:524] == 2'd0 ||
	      !cache_pipeline_first__581_BITS_573_TO_526_644__ETC___d2646) &&
	     cache_cRqMshr$pipelineResp_getRepSucc[4] ;
  assign NOT_cache_pipeline_first__581_BIT_517_582_105__ETC___d3345 =
	     !cache_pipeline$first[517] &&
	     (!cache_cRqMshr$pipelineResp_searchEndOfChain[4] ||
	      cache_cRqMshr$pipelineResp_getState != 3'd1) &&
	     !cache_cRqMshr$pipelineResp_getRq[16] &&
	     cache_pipeline_first__581_BITS_573_TO_526_644__ETC___d2646 &&
	     cache_pipeline$first[525:524] != 2'd0 &&
	     IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2627 &&
	     NOT_IF_cache_pipeline_first__581_BITS_584_TO_5_ETC___d3191 ;
  assign NOT_cache_pipeline_first__581_BIT_517_582_105__ETC___d3351 =
	     !cache_pipeline$first[517] &&
	     (!cache_cRqMshr$pipelineResp_searchEndOfChain[4] ||
	      cache_cRqMshr$pipelineResp_getState != 3'd1) &&
	     !cache_cRqMshr$pipelineResp_getRq[16] &&
	     (cache_pipeline$first[525:524] == 2'd0 ||
	      cache_pipeline_first__581_BITS_573_TO_526_644__ETC___d2646) &&
	     (cache_pipeline$first[525:524] == 2'd0 ||
	      IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3156) &&
	     cache_cRqMshr$pipelineResp_getSlot[12] ;
  assign NOT_cache_pipeline_first__581_BIT_517_582_105__ETC___d3359 =
	     !cache_pipeline$first[517] &&
	     (!cache_cRqMshr$pipelineResp_searchEndOfChain[4] ||
	      cache_cRqMshr$pipelineResp_getState != 3'd1) &&
	     !cache_cRqMshr$pipelineResp_getRq[16] &&
	     cache_pipeline$first[525:524] != 2'd0 &&
	     !cache_pipeline_first__581_BITS_573_TO_526_644__ETC___d2646 &&
	     cache_pipeline$first[519:518] == 2'd0 &&
	     cache_pipeline$first[521:520] == 2'd0 &&
	     cache_pipeline$first[523:522] == 2'd0 &&
	     cache_cRqMshr$pipelineResp_getRepSucc[4] ;
  assign NOT_cache_rqFromCQ_clearReq_dummy2_1_read__8_9_ETC___d33 =
	     !cache_rqFromCQ_clearReq_dummy2_1$Q_OUT ||
	     !cache_rqFromCQ_clearReq_rl ;
  assign NOT_cache_rqFromCQ_enqReq_dummy2_2_read__4_9_O_ETC___d78 =
	     (!cache_rqFromCQ_enqReq_dummy2_2$Q_OUT ||
	      (EN_to_child_rqFromC_enq ?
		 !cache_rqFromCQ_enqReq_lat_0$wget[74] :
		 !cache_rqFromCQ_enqReq_rl[74])) &&
	     (cache_rqFromCQ_deqReq_dummy2_2$Q_OUT &&
	      IF_cache_rqFromCQ_deqReq_lat_1_whas__3_THEN_ca_ETC___d19 ||
	      cache_rqFromCQ_empty) ;
  assign NOT_cache_rqFromDmaQ_clearReq_dummy2_1_read__3_ETC___d339 =
	     !cache_rqFromDmaQ_clearReq_dummy2_1$Q_OUT ||
	     !cache_rqFromDmaQ_clearReq_rl ;
  assign NOT_cache_rqFromDmaQ_enqReq_dummy2_2_read__40__ETC___d384 =
	     (!cache_rqFromDmaQ_enqReq_dummy2_2$Q_OUT ||
	      (EN_dma_memReq_enq ?
		 !cache_rqFromDmaQ_enqReq_lat_0$wget[656] :
		 !cache_rqFromDmaQ_enqReq_rl[656])) &&
	     (cache_rqFromDmaQ_deqReq_dummy2_2$Q_OUT &&
	      IF_cache_rqFromDmaQ_deqReq_lat_1_whas__19_THEN_ETC___d325 ||
	      cache_rqFromDmaQ_empty) ;
  assign NOT_cache_rsFromCQ_clearReq_dummy2_1_read__20__ETC___d125 =
	     !cache_rsFromCQ_clearReq_dummy2_1$Q_OUT ||
	     !cache_rsFromCQ_clearReq_rl ;
  assign NOT_cache_rsFromCQ_enqReq_dummy2_2_read__26_61_ETC___d170 =
	     (!cache_rsFromCQ_enqReq_dummy2_2$Q_OUT ||
	      (EN_to_child_rsFromC_enq ?
		 !cache_rsFromCQ_enqReq_lat_0$wget[581] :
		 !cache_rsFromCQ_enqReq_rl[581])) &&
	     (cache_rsFromCQ_deqReq_dummy2_2$Q_OUT &&
	      IF_cache_rsFromCQ_deqReq_lat_1_whas__05_THEN_c_ETC___d111 ||
	      cache_rsFromCQ_empty) ;
  assign NOT_cache_rsFromMQ_clearReq_dummy2_1_read__35__ETC___d740 =
	     !cache_rsFromMQ_clearReq_dummy2_1$Q_OUT ||
	     !cache_rsFromMQ_clearReq_rl ;
  assign NOT_cache_rsFromMQ_enqReq_dummy2_2_read__41_76_ETC___d785 =
	     (!cache_rsFromMQ_enqReq_dummy2_2$Q_OUT ||
	      (EN_to_mem_rsFromM_enq ?
		 !cache_rsFromMQ_enqReq_lat_0$wget[517] :
		 !cache_rsFromMQ_enqReq_rl[517])) &&
	     (cache_rsFromMQ_deqReq_dummy2_2$Q_OUT &&
	      IF_cache_rsFromMQ_deqReq_lat_1_whas__20_THEN_c_ETC___d726 ||
	      cache_rsFromMQ_empty) ;
  assign NOT_cache_rsLdToDmaQ_clearReq_dummy2_1_read__2_ETC___d430 =
	     !cache_rsLdToDmaQ_clearReq_dummy2_1$Q_OUT ||
	     !cache_rsLdToDmaQ_clearReq_rl ;
  assign NOT_cache_rsLdToDmaQ_enqReq_dummy2_2_read__31__ETC___d475 =
	     (!cache_rsLdToDmaQ_enqReq_dummy2_2$Q_OUT ||
	      (CAN_FIRE_RL_cache_sendRsLdToDma ?
		 !cache_rsLdToDmaQ_enqReq_lat_0$wget[528] :
		 !cache_rsLdToDmaQ_enqReq_rl[528])) &&
	     (cache_rsLdToDmaQ_deqReq_dummy2_2$Q_OUT &&
	      IF_cache_rsLdToDmaQ_deqReq_lat_1_whas__10_THEN_ETC___d416 ||
	      cache_rsLdToDmaQ_empty) ;
  assign NOT_cache_rsStToDmaQ_clearReq_dummy2_1_read__1_ETC___d521 =
	     !cache_rsStToDmaQ_clearReq_dummy2_1$Q_OUT ||
	     !cache_rsStToDmaQ_clearReq_rl ;
  assign NOT_cache_rsStToDmaQ_enqReq_dummy2_2_read__22__ETC___d566 =
	     (!cache_rsStToDmaQ_enqReq_dummy2_2$Q_OUT ||
	      (WILL_FIRE_RL_cache_sendRsStToDma ?
		 !cache_rsStToDmaQ_enqReq_lat_0$wget[16] :
		 !cache_rsStToDmaQ_enqReq_rl[16])) &&
	     (cache_rsStToDmaQ_deqReq_dummy2_2$Q_OUT &&
	      IF_cache_rsStToDmaQ_deqReq_lat_1_whas__01_THEN_ETC___d507 ||
	      cache_rsStToDmaQ_empty) ;
  assign NOT_cache_rsToCIndexQ_clearReq_dummy2_1_read___ETC___d976 =
	     !cache_rsToCIndexQ_clearReq_dummy2_1$Q_OUT ||
	     !cache_rsToCIndexQ_clearReq_rl ;
  assign NOT_cache_rsToCIndexQ_enqReq_dummy2_2_read__51_ETC___d999 =
	     (!cache_rsToCIndexQ_enqReq_dummy2_2$Q_OUT ||
	      (cache_rsToCIndexQ_enqReq_lat_0$whas ?
		 !cache_rsToCIndexQ_enqReq_lat_0$wget[6] :
		 !cache_rsToCIndexQ_enqReq_rl[6])) &&
	     (cache_rsToCIndexQ_deqReq_dummy2_2$Q_OUT &&
	      IF_cache_rsToCIndexQ_deqReq_lat_1_whas__34_THE_ETC___d940 ||
	      cache_rsToCIndexQ_empty) ;
  assign NOT_cache_toCQ_clearReq_dummy2_1_read__47_48_O_ETC___d252 =
	     !cache_toCQ_clearReq_dummy2_1$Q_OUT || !cache_toCQ_clearReq_rl ;
  assign NOT_cache_toCQ_enqReq_dummy2_2_read__53_83_OR__ETC___d292 =
	     (!cache_toCQ_enqReq_dummy2_2$Q_OUT ||
	      (cache_toCQ_enqReq_lat_0$whas ?
		 !cache_toCQ_enqReq_lat_0$wget[585] :
		 !cache_toCQ_enqReq_rl[585])) &&
	     (cache_toCQ_deqReq_dummy2_2$Q_OUT &&
	      IF_cache_toCQ_deqReq_lat_1_whas__32_THEN_cache_ETC___d238 ||
	      cache_toCQ_empty) ;
  assign NOT_cache_toMQ_clearReq_dummy2_1_read__48_49_O_ETC___d653 =
	     !cache_toMQ_clearReq_dummy2_1$Q_OUT || !cache_toMQ_clearReq_rl ;
  assign NOT_cache_toMQ_enqReq_dummy2_2_read__54_84_OR__ETC___d693 =
	     (!cache_toMQ_enqReq_dummy2_2$Q_OUT ||
	      (cache_toMQ_enqReq_lat_0$whas ?
		 !cache_toMQ_enqReq_lat_0$wget[641] :
		 !cache_toMQ_enqReq_rl[641])) &&
	     (cache_toMQ_deqReq_dummy2_2$Q_OUT &&
	      IF_cache_toMQ_deqReq_lat_1_whas__33_THEN_cache_ETC___d639 ||
	      cache_toMQ_empty) ;
  assign NOT_perfReqQ_clearReq_dummy2_1_read__864_865_O_ETC___d3869 =
	     !perfReqQ_clearReq_dummy2_1$Q_OUT || !perfReqQ_clearReq_rl ;
  assign NOT_perfReqQ_enqReq_dummy2_2_read__870_890_OR__ETC___d3900 =
	     (!perfReqQ_enqReq_dummy2_2$Q_OUT ||
	      (EN_perf_req ?
		 !perfReqQ_enqReq_lat_0$wget[4] :
		 !perfReqQ_enqReq_rl[4])) &&
	     (perfReqQ_deqReq_dummy2_2$Q_OUT &&
	      (EN_perf_resp || perfReqQ_deqReq_rl) ||
	      perfReqQ_empty) ;
  assign SEL_ARR_IF_cache_cRqMshr_pipelineResp_getSlot__ETC___d3440 =
	     CASE_cache_pipelinefirst_BITS_580_TO_579_0_ca_ETC__q84 <
	     SEL_ARR_cache_pipeline_first__581_BITS_519_TO__ETC___d3403 ;
  assign SEL_ARR_cache_rqFromCQ_data_0_090_BITS_7_TO_6__ETC___d1118 =
	     { CASE_cache_rqFromCQ_deqP_0_cache_rqFromCQ_data_ETC__q230,
	       CASE_cache_rqFromCQ_deqP_0_cache_rqFromCQ_data_ETC__q231,
	       x__h249082,
	       78'h2AAAAAAAAAAAAAAA8AAA,
	       x__h257564 } ;
  assign SEL_ARR_cache_rqFromDmaQ_data_0_129_BITS_527_T_ETC___d1827 =
	     { CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q91,
	       CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q92,
	       CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q93 } ;
  assign SEL_ARR_cache_rqFromDmaQ_data_0_129_BITS_527_T_ETC___d1836 =
	     { SEL_ARR_cache_rqFromDmaQ_data_0_129_BITS_527_T_ETC___d1827,
	       CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q98,
	       CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q99 } ;
  assign SEL_ARR_cache_rqFromDmaQ_data_0_129_BITS_527_T_ETC___d1845 =
	     { SEL_ARR_cache_rqFromDmaQ_data_0_129_BITS_527_T_ETC___d1836,
	       CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q232,
	       CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q233 } ;
  assign SEL_ARR_cache_rqFromDmaQ_data_0_129_BIT_591_57_ETC___d1656 =
	     { CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q80,
	       CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q81,
	       CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q82,
	       CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q83 } ;
  assign SEL_ARR_cache_rqFromDmaQ_data_0_129_BIT_591_57_ETC___d1661 =
	     { SEL_ARR_cache_rqFromDmaQ_data_0_129_BIT_591_57_ETC___d1656,
	       CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q106,
	       CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q107 } ;
  assign SEL_ARR_cache_rqFromDmaQ_data_0_129_BIT_591_57_ETC___d1666 =
	     { SEL_ARR_cache_rqFromDmaQ_data_0_129_BIT_591_57_ETC___d1661,
	       CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q110,
	       CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q111 } ;
  assign SEL_ARR_cache_rqFromDmaQ_data_0_129_BIT_591_57_ETC___d1671 =
	     { SEL_ARR_cache_rqFromDmaQ_data_0_129_BIT_591_57_ETC___d1666,
	       CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q114,
	       CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q115 } ;
  assign SEL_ARR_cache_rqFromDmaQ_data_0_129_BIT_591_57_ETC___d1676 =
	     { SEL_ARR_cache_rqFromDmaQ_data_0_129_BIT_591_57_ETC___d1671,
	       CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q118,
	       CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q119 } ;
  assign SEL_ARR_cache_rqFromDmaQ_data_0_129_BIT_591_57_ETC___d1681 =
	     { SEL_ARR_cache_rqFromDmaQ_data_0_129_BIT_591_57_ETC___d1676,
	       CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q122,
	       CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q123 } ;
  assign SEL_ARR_cache_rqFromDmaQ_data_0_129_BIT_591_57_ETC___d1686 =
	     { SEL_ARR_cache_rqFromDmaQ_data_0_129_BIT_591_57_ETC___d1681,
	       CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q126,
	       CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q127 } ;
  assign SEL_ARR_cache_rqFromDmaQ_data_0_129_BIT_591_57_ETC___d1691 =
	     { SEL_ARR_cache_rqFromDmaQ_data_0_129_BIT_591_57_ETC___d1686,
	       CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q130,
	       CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q131 } ;
  assign SEL_ARR_cache_rqFromDmaQ_data_0_129_BIT_591_57_ETC___d1696 =
	     { SEL_ARR_cache_rqFromDmaQ_data_0_129_BIT_591_57_ETC___d1691,
	       CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q134,
	       CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q135 } ;
  assign SEL_ARR_cache_rqFromDmaQ_data_0_129_BIT_591_57_ETC___d1701 =
	     { SEL_ARR_cache_rqFromDmaQ_data_0_129_BIT_591_57_ETC___d1696,
	       CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q138,
	       CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q139 } ;
  assign SEL_ARR_cache_rqFromDmaQ_data_0_129_BIT_591_57_ETC___d1706 =
	     { SEL_ARR_cache_rqFromDmaQ_data_0_129_BIT_591_57_ETC___d1701,
	       CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q142,
	       CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q143 } ;
  assign SEL_ARR_cache_rqFromDmaQ_data_0_129_BIT_591_57_ETC___d1711 =
	     { SEL_ARR_cache_rqFromDmaQ_data_0_129_BIT_591_57_ETC___d1706,
	       CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q146,
	       CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q147 } ;
  assign SEL_ARR_cache_rqFromDmaQ_data_0_129_BIT_591_57_ETC___d1716 =
	     { SEL_ARR_cache_rqFromDmaQ_data_0_129_BIT_591_57_ETC___d1711,
	       CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q150,
	       CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q151 } ;
  assign SEL_ARR_cache_rqFromDmaQ_data_0_129_BIT_591_57_ETC___d1721 =
	     { SEL_ARR_cache_rqFromDmaQ_data_0_129_BIT_591_57_ETC___d1716,
	       CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q154,
	       CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q155 } ;
  assign SEL_ARR_cache_rqFromDmaQ_data_0_129_BIT_591_57_ETC___d1726 =
	     { SEL_ARR_cache_rqFromDmaQ_data_0_129_BIT_591_57_ETC___d1721,
	       CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q158,
	       CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q159 } ;
  assign SEL_ARR_cache_rqFromDmaQ_data_0_129_BIT_591_57_ETC___d1731 =
	     { SEL_ARR_cache_rqFromDmaQ_data_0_129_BIT_591_57_ETC___d1726,
	       CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q162,
	       CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q163 } ;
  assign SEL_ARR_cache_rqFromDmaQ_data_0_129_BIT_591_57_ETC___d1736 =
	     { SEL_ARR_cache_rqFromDmaQ_data_0_129_BIT_591_57_ETC___d1731,
	       CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q166,
	       CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q167 } ;
  assign SEL_ARR_cache_rqFromDmaQ_data_0_129_BIT_591_57_ETC___d1741 =
	     { SEL_ARR_cache_rqFromDmaQ_data_0_129_BIT_591_57_ETC___d1736,
	       CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q170,
	       CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q171 } ;
  assign SEL_ARR_cache_rqFromDmaQ_data_0_129_BIT_591_57_ETC___d1746 =
	     { SEL_ARR_cache_rqFromDmaQ_data_0_129_BIT_591_57_ETC___d1741,
	       CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q174,
	       CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q175 } ;
  assign SEL_ARR_cache_rqFromDmaQ_data_0_129_BIT_591_57_ETC___d1751 =
	     { SEL_ARR_cache_rqFromDmaQ_data_0_129_BIT_591_57_ETC___d1746,
	       CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q178,
	       CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q179 } ;
  assign SEL_ARR_cache_rqFromDmaQ_data_0_129_BIT_591_57_ETC___d1756 =
	     { SEL_ARR_cache_rqFromDmaQ_data_0_129_BIT_591_57_ETC___d1751,
	       CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q182,
	       CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q183 } ;
  assign SEL_ARR_cache_rqFromDmaQ_data_0_129_BIT_591_57_ETC___d1761 =
	     { SEL_ARR_cache_rqFromDmaQ_data_0_129_BIT_591_57_ETC___d1756,
	       CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q186,
	       CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q187 } ;
  assign SEL_ARR_cache_rqFromDmaQ_data_0_129_BIT_591_57_ETC___d1766 =
	     { SEL_ARR_cache_rqFromDmaQ_data_0_129_BIT_591_57_ETC___d1761,
	       CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q190,
	       CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q191 } ;
  assign SEL_ARR_cache_rqFromDmaQ_data_0_129_BIT_591_57_ETC___d1771 =
	     { SEL_ARR_cache_rqFromDmaQ_data_0_129_BIT_591_57_ETC___d1766,
	       CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q194,
	       CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q195 } ;
  assign SEL_ARR_cache_rqFromDmaQ_data_0_129_BIT_591_57_ETC___d1776 =
	     { SEL_ARR_cache_rqFromDmaQ_data_0_129_BIT_591_57_ETC___d1771,
	       CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q198,
	       CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q199 } ;
  assign SEL_ARR_cache_rqFromDmaQ_data_0_129_BIT_591_57_ETC___d1781 =
	     { SEL_ARR_cache_rqFromDmaQ_data_0_129_BIT_591_57_ETC___d1776,
	       CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q202,
	       CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q203 } ;
  assign SEL_ARR_cache_rqFromDmaQ_data_0_129_BIT_591_57_ETC___d1786 =
	     { SEL_ARR_cache_rqFromDmaQ_data_0_129_BIT_591_57_ETC___d1781,
	       CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q206,
	       CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q207 } ;
  assign SEL_ARR_cache_rqFromDmaQ_data_0_129_BIT_591_57_ETC___d1791 =
	     { SEL_ARR_cache_rqFromDmaQ_data_0_129_BIT_591_57_ETC___d1786,
	       CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q210,
	       CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q211 } ;
  assign SEL_ARR_cache_rqFromDmaQ_data_0_129_BIT_591_57_ETC___d1796 =
	     { SEL_ARR_cache_rqFromDmaQ_data_0_129_BIT_591_57_ETC___d1791,
	       CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q214,
	       CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q215 } ;
  assign SEL_ARR_cache_rqFromDmaQ_data_0_129_BIT_591_57_ETC___d1801 =
	     { SEL_ARR_cache_rqFromDmaQ_data_0_129_BIT_591_57_ETC___d1796,
	       CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q218,
	       CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q219 } ;
  assign SEL_ARR_cache_rqFromDmaQ_data_0_129_BIT_591_57_ETC___d1806 =
	     { SEL_ARR_cache_rqFromDmaQ_data_0_129_BIT_591_57_ETC___d1801,
	       CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q228,
	       CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q229 } ;
  assign SEL_ARR_cache_rsFromCQ_data_0_855_BITS_513_TO__ETC___d1886 =
	     { CASE_cache_rsFromCQ_deqP_0_cache_rsFromCQ_data_ETC__q69,
	       CASE_cache_rsFromCQ_deqP_0_cache_rsFromCQ_data_ETC__q70,
	       CASE_cache_rsFromCQ_deqP_0_cache_rsFromCQ_data_ETC__q71,
	       CASE_cache_rsFromCQ_deqP_0_cache_rsFromCQ_data_ETC__q72 } ;
  assign SEL_ARR_cache_rsFromCQ_data_0_855_BITS_513_TO__ETC___d1895 =
	     { SEL_ARR_cache_rsFromCQ_data_0_855_BITS_513_TO__ETC___d1886,
	       CASE_cache_rsFromCQ_deqP_0_cache_rsFromCQ_data_ETC__q75,
	       CASE_cache_rsFromCQ_deqP_0_cache_rsFromCQ_data_ETC__q76 } ;
  assign SEL_ARR_cache_rsFromCQ_data_0_855_BITS_513_TO__ETC___d1904 =
	     { SEL_ARR_cache_rsFromCQ_data_0_855_BITS_513_TO__ETC___d1895,
	       CASE_cache_rsFromCQ_deqP_0_cache_rsFromCQ_data_ETC__q236,
	       CASE_cache_rsFromCQ_deqP_0_cache_rsFromCQ_data_ETC__q237 } ;
  assign SEL_ARR_cache_rsFromCQ_data_0_855_BITS_580_TO__ETC___d1910 =
	     { CASE_cache_rsFromCQ_deqP_0_cache_rsFromCQ_data_ETC__q243,
	       CASE_cache_rsFromCQ_deqP_0_cache_rsFromCQ_data_ETC__q244,
	       SEL_ARR_cache_rsFromCQ_data_0_855_BIT_514_865__ETC___d1909 } ;
  assign SEL_ARR_cache_rsFromCQ_data_0_855_BIT_514_865__ETC___d1909 =
	     { CASE_cache_rsFromCQ_deqP_0_cache_rsFromCQ_data_ETC__q242,
	       SEL_ARR_cache_rsFromCQ_data_0_855_BITS_513_TO__ETC___d1904,
	       x__h275130 } ;
  assign SEL_ARR_cache_rsFromMQ_data_0_914_BITS_516_TO__ETC___d1948 =
	     { CASE_cache_rsFromMQ_deqP_0_cache_rsFromMQ_data_ETC__q1,
	       CASE_cache_rsFromMQ_deqP_0_cache_rsFromMQ_data_ETC__q2,
	       CASE_cache_rsFromMQ_deqP_0_cache_rsFromMQ_data_ETC__q3,
	       CASE_cache_rsFromMQ_deqP_0_cache_rsFromMQ_data_ETC__q4 } ;
  assign SEL_ARR_cache_rsFromMQ_data_0_914_BITS_516_TO__ETC___d1957 =
	     { SEL_ARR_cache_rsFromMQ_data_0_914_BITS_516_TO__ETC___d1948,
	       CASE_cache_rsFromMQ_deqP_0_cache_rsFromMQ_data_ETC__q73,
	       CASE_cache_rsFromMQ_deqP_0_cache_rsFromMQ_data_ETC__q74 } ;
  assign SEL_ARR_cache_rsFromMQ_data_0_914_BITS_516_TO__ETC___d1966 =
	     { SEL_ARR_cache_rsFromMQ_data_0_914_BITS_516_TO__ETC___d1957,
	       CASE_cache_rsFromMQ_deqP_0_cache_rsFromMQ_data_ETC__q226,
	       CASE_cache_rsFromMQ_deqP_0_cache_rsFromMQ_data_ETC__q227 } ;
  assign SEL_ARR_cache_rsLdToDmaQ_data_0_004_BITS_527_T_ETC___d4018 =
	     { CASE_cache_rsLdToDmaQ_deqP_0_cache_rsLdToDmaQ__ETC__q85,
	       CASE_cache_rsLdToDmaQ_deqP_0_cache_rsLdToDmaQ__ETC__q86,
	       CASE_cache_rsLdToDmaQ_deqP_0_cache_rsLdToDmaQ__ETC__q87 } ;
  assign SEL_ARR_cache_rsLdToDmaQ_data_0_004_BITS_527_T_ETC___d4027 =
	     { SEL_ARR_cache_rsLdToDmaQ_data_0_004_BITS_527_T_ETC___d4018,
	       CASE_cache_rsLdToDmaQ_deqP_0_cache_rsLdToDmaQ__ETC__q96,
	       CASE_cache_rsLdToDmaQ_deqP_0_cache_rsLdToDmaQ__ETC__q97 } ;
  assign SEL_ARR_cache_rsLdToDmaQ_data_0_004_BITS_527_T_ETC___d4036 =
	     { SEL_ARR_cache_rsLdToDmaQ_data_0_004_BITS_527_T_ETC___d4027,
	       CASE_cache_rsLdToDmaQ_deqP_0_cache_rsLdToDmaQ__ETC__q257,
	       CASE_cache_rsLdToDmaQ_deqP_0_cache_rsLdToDmaQ__ETC__q258 } ;
  assign SEL_ARR_cache_toCQ_data_0_917_BITS_514_TO_451__ETC___d3969 =
	     { CASE_cache_toCQ_deqP_0_cache_toCQ_data_0_BITS__ETC__q88,
	       CASE_cache_toCQ_deqP_0_cache_toCQ_data_0_BITS__ETC__q89,
	       CASE_cache_toCQ_deqP_0_cache_toCQ_data_0_BITS__ETC__q90 } ;
  assign SEL_ARR_cache_toCQ_data_0_917_BITS_514_TO_451__ETC___d3978 =
	     { SEL_ARR_cache_toCQ_data_0_917_BITS_514_TO_451__ETC___d3969,
	       CASE_cache_toCQ_deqP_0_cache_toCQ_data_0_BITS__ETC__q94,
	       CASE_cache_toCQ_deqP_0_cache_toCQ_data_0_BITS__ETC__q95 } ;
  assign SEL_ARR_cache_toCQ_data_0_917_BITS_514_TO_451__ETC___d3987 =
	     { SEL_ARR_cache_toCQ_data_0_917_BITS_514_TO_451__ETC___d3978,
	       CASE_cache_toCQ_deqP_0_cache_toCQ_data_0_BITS__ETC__q234,
	       CASE_cache_toCQ_deqP_0_cache_toCQ_data_0_BITS__ETC__q235 } ;
  assign SEL_ARR_cache_toCQ_data_0_917_BITS_583_TO_520__ETC___d3998 =
	     { CASE_cache_toCQ_deqP_0_cache_toCQ_data_0_BITS__ETC__q247,
	       CASE_cache_toCQ_deqP_0_cache_toCQ_data_0_BITS__ETC__q248,
	       x__h444405,
	       SEL_ARR_cache_toCQ_data_0_917_BIT_515_953_cach_ETC___d3992,
	       x__h445950 } ;
  assign SEL_ARR_cache_toCQ_data_0_917_BIT_515_953_cach_ETC___d3992 =
	     { CASE_cache_toCQ_deqP_0_cache_toCQ_data_0_BIT_5_ETC__q238,
	       SEL_ARR_cache_toCQ_data_0_917_BITS_514_TO_451__ETC___d3987,
	       CASE_cache_toCQ_deqP_0_cache_toCQ_data_0_BITS__ETC__q239 } ;
  assign SEL_ARR_cache_toMQ_data_0_050_BITS_511_TO_448__ETC___d4383 =
	     { CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BITS__ETC__q220,
	       CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BITS__ETC__q221,
	       CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BITS__ETC__q222,
	       CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BITS__ETC__q223 } ;
  assign SEL_ARR_cache_toMQ_data_0_050_BITS_511_TO_448__ETC___d4392 =
	     { SEL_ARR_cache_toMQ_data_0_050_BITS_511_TO_448__ETC___d4383,
	       CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BITS__ETC__q224,
	       CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BITS__ETC__q225 } ;
  assign SEL_ARR_cache_toMQ_data_0_050_BITS_511_TO_448__ETC___d4401 =
	     { SEL_ARR_cache_toMQ_data_0_050_BITS_511_TO_448__ETC___d4392,
	       CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BITS__ETC__q245,
	       CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BITS__ETC__q246 } ;
  assign SEL_ARR_cache_toMQ_data_0_050_BITS_639_TO_576__ETC___d4402 =
	     { CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BITS__ETC__q251,
	       SEL_ARR_cache_toMQ_data_0_050_BIT_575_078_cach_ETC___d4365,
	       SEL_ARR_cache_toMQ_data_0_050_BITS_511_TO_448__ETC___d4401 } ;
  assign SEL_ARR_cache_toMQ_data_0_050_BIT_575_078_cach_ETC___d4095 =
	     { CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q100,
	       CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q101,
	       CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q102,
	       CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q103 } ;
  assign SEL_ARR_cache_toMQ_data_0_050_BIT_575_078_cach_ETC___d4104 =
	     { SEL_ARR_cache_toMQ_data_0_050_BIT_575_078_cach_ETC___d4095,
	       CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q104,
	       CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q105 } ;
  assign SEL_ARR_cache_toMQ_data_0_050_BIT_575_078_cach_ETC___d4113 =
	     { SEL_ARR_cache_toMQ_data_0_050_BIT_575_078_cach_ETC___d4104,
	       CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q108,
	       CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q109 } ;
  assign SEL_ARR_cache_toMQ_data_0_050_BIT_575_078_cach_ETC___d4122 =
	     { SEL_ARR_cache_toMQ_data_0_050_BIT_575_078_cach_ETC___d4113,
	       CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q112,
	       CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q113 } ;
  assign SEL_ARR_cache_toMQ_data_0_050_BIT_575_078_cach_ETC___d4131 =
	     { SEL_ARR_cache_toMQ_data_0_050_BIT_575_078_cach_ETC___d4122,
	       CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q116,
	       CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q117 } ;
  assign SEL_ARR_cache_toMQ_data_0_050_BIT_575_078_cach_ETC___d4140 =
	     { SEL_ARR_cache_toMQ_data_0_050_BIT_575_078_cach_ETC___d4131,
	       CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q120,
	       CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q121 } ;
  assign SEL_ARR_cache_toMQ_data_0_050_BIT_575_078_cach_ETC___d4149 =
	     { SEL_ARR_cache_toMQ_data_0_050_BIT_575_078_cach_ETC___d4140,
	       CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q124,
	       CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q125 } ;
  assign SEL_ARR_cache_toMQ_data_0_050_BIT_575_078_cach_ETC___d4158 =
	     { SEL_ARR_cache_toMQ_data_0_050_BIT_575_078_cach_ETC___d4149,
	       CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q128,
	       CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q129 } ;
  assign SEL_ARR_cache_toMQ_data_0_050_BIT_575_078_cach_ETC___d4167 =
	     { SEL_ARR_cache_toMQ_data_0_050_BIT_575_078_cach_ETC___d4158,
	       CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q132,
	       CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q133 } ;
  assign SEL_ARR_cache_toMQ_data_0_050_BIT_575_078_cach_ETC___d4176 =
	     { SEL_ARR_cache_toMQ_data_0_050_BIT_575_078_cach_ETC___d4167,
	       CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q136,
	       CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q137 } ;
  assign SEL_ARR_cache_toMQ_data_0_050_BIT_575_078_cach_ETC___d4185 =
	     { SEL_ARR_cache_toMQ_data_0_050_BIT_575_078_cach_ETC___d4176,
	       CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q140,
	       CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q141 } ;
  assign SEL_ARR_cache_toMQ_data_0_050_BIT_575_078_cach_ETC___d4194 =
	     { SEL_ARR_cache_toMQ_data_0_050_BIT_575_078_cach_ETC___d4185,
	       CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q144,
	       CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q145 } ;
  assign SEL_ARR_cache_toMQ_data_0_050_BIT_575_078_cach_ETC___d4203 =
	     { SEL_ARR_cache_toMQ_data_0_050_BIT_575_078_cach_ETC___d4194,
	       CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q148,
	       CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q149 } ;
  assign SEL_ARR_cache_toMQ_data_0_050_BIT_575_078_cach_ETC___d4212 =
	     { SEL_ARR_cache_toMQ_data_0_050_BIT_575_078_cach_ETC___d4203,
	       CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q152,
	       CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q153 } ;
  assign SEL_ARR_cache_toMQ_data_0_050_BIT_575_078_cach_ETC___d4221 =
	     { SEL_ARR_cache_toMQ_data_0_050_BIT_575_078_cach_ETC___d4212,
	       CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q156,
	       CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q157 } ;
  assign SEL_ARR_cache_toMQ_data_0_050_BIT_575_078_cach_ETC___d4230 =
	     { SEL_ARR_cache_toMQ_data_0_050_BIT_575_078_cach_ETC___d4221,
	       CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q160,
	       CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q161 } ;
  assign SEL_ARR_cache_toMQ_data_0_050_BIT_575_078_cach_ETC___d4239 =
	     { SEL_ARR_cache_toMQ_data_0_050_BIT_575_078_cach_ETC___d4230,
	       CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q164,
	       CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q165 } ;
  assign SEL_ARR_cache_toMQ_data_0_050_BIT_575_078_cach_ETC___d4248 =
	     { SEL_ARR_cache_toMQ_data_0_050_BIT_575_078_cach_ETC___d4239,
	       CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q168,
	       CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q169 } ;
  assign SEL_ARR_cache_toMQ_data_0_050_BIT_575_078_cach_ETC___d4257 =
	     { SEL_ARR_cache_toMQ_data_0_050_BIT_575_078_cach_ETC___d4248,
	       CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q172,
	       CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q173 } ;
  assign SEL_ARR_cache_toMQ_data_0_050_BIT_575_078_cach_ETC___d4266 =
	     { SEL_ARR_cache_toMQ_data_0_050_BIT_575_078_cach_ETC___d4257,
	       CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q176,
	       CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q177 } ;
  assign SEL_ARR_cache_toMQ_data_0_050_BIT_575_078_cach_ETC___d4275 =
	     { SEL_ARR_cache_toMQ_data_0_050_BIT_575_078_cach_ETC___d4266,
	       CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q180,
	       CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q181 } ;
  assign SEL_ARR_cache_toMQ_data_0_050_BIT_575_078_cach_ETC___d4284 =
	     { SEL_ARR_cache_toMQ_data_0_050_BIT_575_078_cach_ETC___d4275,
	       CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q184,
	       CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q185 } ;
  assign SEL_ARR_cache_toMQ_data_0_050_BIT_575_078_cach_ETC___d4293 =
	     { SEL_ARR_cache_toMQ_data_0_050_BIT_575_078_cach_ETC___d4284,
	       CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q188,
	       CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q189 } ;
  assign SEL_ARR_cache_toMQ_data_0_050_BIT_575_078_cach_ETC___d4302 =
	     { SEL_ARR_cache_toMQ_data_0_050_BIT_575_078_cach_ETC___d4293,
	       CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q192,
	       CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q193 } ;
  assign SEL_ARR_cache_toMQ_data_0_050_BIT_575_078_cach_ETC___d4311 =
	     { SEL_ARR_cache_toMQ_data_0_050_BIT_575_078_cach_ETC___d4302,
	       CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q196,
	       CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q197 } ;
  assign SEL_ARR_cache_toMQ_data_0_050_BIT_575_078_cach_ETC___d4320 =
	     { SEL_ARR_cache_toMQ_data_0_050_BIT_575_078_cach_ETC___d4311,
	       CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q200,
	       CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q201 } ;
  assign SEL_ARR_cache_toMQ_data_0_050_BIT_575_078_cach_ETC___d4329 =
	     { SEL_ARR_cache_toMQ_data_0_050_BIT_575_078_cach_ETC___d4320,
	       CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q204,
	       CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q205 } ;
  assign SEL_ARR_cache_toMQ_data_0_050_BIT_575_078_cach_ETC___d4338 =
	     { SEL_ARR_cache_toMQ_data_0_050_BIT_575_078_cach_ETC___d4329,
	       CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q208,
	       CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q209 } ;
  assign SEL_ARR_cache_toMQ_data_0_050_BIT_575_078_cach_ETC___d4347 =
	     { SEL_ARR_cache_toMQ_data_0_050_BIT_575_078_cach_ETC___d4338,
	       CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q212,
	       CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q213 } ;
  assign SEL_ARR_cache_toMQ_data_0_050_BIT_575_078_cach_ETC___d4356 =
	     { SEL_ARR_cache_toMQ_data_0_050_BIT_575_078_cach_ETC___d4347,
	       CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q216,
	       CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q217 } ;
  assign SEL_ARR_cache_toMQ_data_0_050_BIT_575_078_cach_ETC___d4365 =
	     { SEL_ARR_cache_toMQ_data_0_050_BIT_575_078_cach_ETC___d4356,
	       CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q240,
	       CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q241 } ;
  assign _0_CONCAT_IF_cache_pipeline_first__581_BITS_523_ETC___d3043 =
	     { 1'd0,
	       IF_cache_pipeline_first__581_BITS_523_TO_522_6_ETC___d3041,
	       cache_pipeline_first__581_BITS_519_TO_518_594__ETC___d2598 ?
		 4'd2 :
		 { 2'd1,
		   IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2597 } } ;
  assign _0_OR_IF_SEL_ARR_cache_pipeline_first__581_BITS_ETC___d3423 =
	     IF_SEL_ARR_cache_pipeline_first__581_BITS_519__ETC___d3418 ||
	     cache_toMInfoQ$FULL_N &&
	     (!cache_cRqMshr$pipelineResp_getRepSucc[4] ||
	      !cache_cRqRetryIndexQ_full) ;
  assign _0_OR_NOT_CASE_IF_cache_pipeline_first__581_BIT_ETC___d3468 =
	     IF_SEL_ARR_cache_cRqMshr_pipelineResp_getSlot__ETC___d3455 ||
	     IF_SEL_ARR_cache_cRqMshr_pipelineResp_getSlot__ETC___d3459 ||
	     IF_SEL_ARR_cache_cRqMshr_pipelineResp_getSlot__ETC___d3463 ||
	     (cache_cRqMshr$pipelineResp_getRq[16] ?
		IF_cache_pipeline_RDY_first__579_AND_cache_cRq_ETC___d2613 :
		!cache_rsToCIndexQ_full) ;
  assign _0_OR_NOT_cache_pipeline_first__581_BITS_519_TO_ETC___d2614 =
	     !cache_pipeline_first__581_BITS_519_TO_518_594__ETC___d2598 ||
	     !cache_pipeline_first__581_BITS_521_TO_520_600__ETC___d2601 ||
	     !cache_pipeline_first__581_BITS_523_TO_522_603__ETC___d2604 ||
	     IF_cache_pipeline_RDY_first__579_AND_cache_cRq_ETC___d2613 ;
  assign _theResult_____2__h119142 =
	     (cache_rqFromDmaQ_deqReq_dummy2_2$Q_OUT &&
	      IF_cache_rqFromDmaQ_deqReq_lat_1_whas__19_THEN_ETC___d325) ?
	       next_deqP___1__h119479 :
	       cache_rqFromDmaQ_deqP ;
  assign _theResult_____2__h135235 =
	     (cache_rsLdToDmaQ_deqReq_dummy2_2$Q_OUT &&
	      IF_cache_rsLdToDmaQ_deqReq_lat_1_whas__10_THEN_ETC___d416) ?
	       next_deqP___1__h135572 :
	       cache_rsLdToDmaQ_deqP ;
  assign _theResult_____2__h142737 =
	     (cache_rsStToDmaQ_deqReq_dummy2_2$Q_OUT &&
	      IF_cache_rsStToDmaQ_deqReq_lat_1_whas__01_THEN_ETC___d507) ?
	       next_deqP___1__h143074 :
	       cache_rsStToDmaQ_deqP ;
  assign _theResult_____2__h208521 =
	     (cache_toMQ_deqReq_dummy2_2$Q_OUT &&
	      IF_cache_toMQ_deqReq_lat_1_whas__33_THEN_cache_ETC___d639) ?
	       next_deqP___1__h208858 :
	       cache_toMQ_deqP ;
  assign _theResult_____2__h22297 =
	     (cache_rsFromCQ_deqReq_dummy2_2$Q_OUT &&
	      IF_cache_rsFromCQ_deqReq_lat_1_whas__05_THEN_c_ETC___d111) ?
	       next_deqP___1__h22634 :
	       cache_rsFromCQ_deqP ;
  assign _theResult_____2__h225016 =
	     (cache_rsFromMQ_deqReq_dummy2_2$Q_OUT &&
	      IF_cache_rsFromMQ_deqReq_lat_1_whas__20_THEN_c_ETC___d726) ?
	       next_deqP___1__h225353 :
	       cache_rsFromMQ_deqP ;
  assign _theResult_____2__h234513 =
	     (cache_cRqRetryIndexQ_deqReq_dummy2_2$Q_OUT &&
	      IF_cache_cRqRetryIndexQ_deqReq_lat_1_whas__11__ETC___d817) ?
	       next_deqP___1__h234850 :
	       cache_cRqRetryIndexQ_deqP ;
  assign _theResult_____2__h245988 =
	     (cache_rsToCIndexQ_deqReq_dummy2_2$Q_OUT &&
	      IF_cache_rsToCIndexQ_deqReq_lat_1_whas__34_THE_ETC___d940) ?
	       next_deqP___1__h246325 :
	       cache_rsToCIndexQ_deqP ;
  assign _theResult_____2__h37990 =
	     (cache_toCQ_deqReq_dummy2_2$Q_OUT &&
	      IF_cache_toCQ_deqReq_lat_1_whas__32_THEN_cache_ETC___d238) ?
	       next_deqP___1__h38327 :
	       cache_toCQ_deqP ;
  assign _theResult_____2__h7215 =
	     (cache_rqFromCQ_deqReq_dummy2_2$Q_OUT &&
	      IF_cache_rqFromCQ_deqReq_lat_1_whas__3_THEN_ca_ETC___d19) ?
	       next_deqP___1__h7552 :
	       cache_rqFromCQ_deqP ;
  assign addr__h288271 =
	     { cache_cRqMshr$sendToM_getSlot[60:13],
	       cache_cRqMshr$sendToM_getRq[103:88] } ;
  assign cache_cRqMshr_pipelineResp_getRq_IF_cache_pipe_ETC___d2995 =
	     { cache_cRqMshr$pipelineResp_getRq[151:104],
	       cache_cRqMshr$pipelineResp_getRq[16] ?
		 IF_cache_pipeline_first__581_BITS_519_TO_518_5_ETC___d2693 :
		 IF_IF_cache_cRqMshr_pipelineResp_getRq_IF_cach_ETC___d2699,
	       cache_cRqMshr$pipelineResp_getRq[16] ?
		 IF_cache_pipeline_first__581_BITS_519_TO_518_5_ETC___d2993 :
		 cache_pipeline$first[511:0] } ;
  assign cache_cRqMshr_pipelineResp_getRq_IF_cache_pipe_ETC___d3123 =
	     cache_cRqMshr$pipelineResp_getRq[16] ||
	     ((cache_pipeline$first[525:524] == 2'd0 ||
	       cache_pipeline_first__581_BITS_573_TO_526_644__ETC___d2646) ?
		CASE_cache_cRqMshrpipelineResp_getRq_BITS_82__ETC__q79 ==
		2'd0 :
		cache_pipeline$first[525:524] == 2'd3) ;
  assign cache_cRqMshr_pipelineResp_getRq_IF_cache_pipe_ETC___d3166 =
	     cache_cRqMshr$pipelineResp_getRq[16] &&
	     (cache_pipeline$first[525:524] == 2'd0 ||
	      !cache_pipeline_first__581_BITS_573_TO_526_644__ETC___d2646) ||
	     !cache_cRqMshr$pipelineResp_getRq[16] &&
	     (cache_pipeline$first[525:524] == 2'd0 ||
	      !cache_pipeline_first__581_BITS_573_TO_526_644__ETC___d2646 &&
	      cache_pipeline$first[519:518] == 2'd0 &&
	      cache_pipeline$first[521:520] == 2'd0 &&
	      cache_pipeline$first[523:522] == 2'd0) ;
  assign cache_cRqMshr_pipelineResp_getRq_IF_cache_pipe_ETC___d3658 =
	     { cache_cRqMshr$pipelineResp_getRq[151:104],
	       IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3493,
	       cache_cRqMshr$pipelineResp_getRq[16] ?
		 IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3656 :
		 cache_pipeline$first[511:0] } ;
  assign cache_cRqMshr_pipelineResp_getSlot_IF_cache_pi_ETC___d3754 =
	     { cache_cRqMshr$pipelineResp_getSlot[64:12],
	       IF_SEL_ARR_cache_cRqMshr_pipelineResp_getSlot__ETC___d3713,
	       cache_cRqMshr$pipelineResp_getSlot[9:8],
	       IF_SEL_ARR_cache_cRqMshr_pipelineResp_getSlot__ETC___d3727,
	       cache_cRqMshr$pipelineResp_getSlot[5:4],
	       IF_SEL_ARR_cache_cRqMshr_pipelineResp_getSlot__ETC___d3742,
	       cache_cRqMshr$pipelineResp_getSlot[1:0] } ;
  assign cache_cRqMshr_pipelineResp_searchEndOfChain_ca_ETC___d2669 =
	     cache_cRqMshr$pipelineResp_searchEndOfChain[4] &&
	     cache_cRqMshr$pipelineResp_getState == 3'd1 ||
	     (cache_cRqMshr$pipelineResp_getRq[16] ?
		IF_NOT_cache_pipeline_first__581_BITS_525_TO_5_ETC___d2654 :
		IF_cache_pipeline_first__581_BITS_525_TO_524_6_ETC___d2667) ;
  assign cache_cRqMshr_sendRqToC_searchNeedRqChild_1_CO_ETC___d2482 =
	     cache_cRqMshr$sendRqToC_searchNeedRqChild[4] &&
	     (!cache_pipeline$notEmpty || cache_pipeline$RDY_unguard_first) &&
	     (!cache_pipeline$notEmpty ||
	      CASE_cache_pipelineunguard_first_BITS_584_TO__ETC__q77) ;
  assign cache_cRqMshrpipelineResp_getData_BITS_63_TO_0__q78 =
	     cache_cRqMshr$pipelineResp_getData[63:0] ;
  assign cache_cRqRetryIndexQ_enqReq_dummy2_2_read__28__ETC___d864 =
	     cache_cRqRetryIndexQ_enqReq_dummy2_2$Q_OUT &&
	     IF_cache_cRqRetryIndexQ_enqReq_lat_1_whas__01__ETC___d833 ||
	     (!cache_cRqRetryIndexQ_deqReq_dummy2_2$Q_OUT ||
	      !WILL_FIRE_RL_cache_cRqTransfer_retry &&
	      !cache_cRqRetryIndexQ_deqReq_rl) &&
	     cache_cRqRetryIndexQ_full ;
  assign cache_pipeline_RDY_deqWrite__580_AND_IF_cache__ETC___d2671 =
	     cache_pipeline$RDY_deqWrite &&
	     (cache_pipeline$first[517] ?
		NOT_cache_pipeline_first__581_BITS_516_TO_513__ETC___d2637 :
		cache_cRqMshr_pipelineResp_searchEndOfChain_ca_ETC___d2669) ;
  assign cache_pipeline_RDY_deqWrite__580_AND_NOT_cache_ETC___d3471 =
	     cache_pipeline$RDY_deqWrite &&
	     (!cache_pipeline$first[517] ||
	      (cache_pipeline$first[512] ?
		 _0_OR_IF_SEL_ARR_cache_pipeline_first__581_BITS_ETC___d3423 :
		 _0_OR_NOT_CASE_IF_cache_pipeline_first__581_BIT_ETC___d3468)) ;
  assign cache_pipeline_first__581_BITS_516_TO_513_583__ETC___d2588 =
	     cache_pipeline$first[516:513] == cache_pipeline$first[582:579] ;
  assign cache_pipeline_first__581_BITS_516_TO_513_583__ETC___d3103 =
	     cache_pipeline_first__581_BITS_516_TO_513_583__ETC___d2588 &&
	     (cache_cRqMshr$pipelineResp_getRq[16] &&
	      cache_pipeline_first__581_BITS_519_TO_518_594__ETC___d2598 &&
	      cache_pipeline_first__581_BITS_521_TO_520_600__ETC___d2601 &&
	      cache_pipeline_first__581_BITS_523_TO_522_603__ETC___d2604 ||
	      !cache_cRqMshr$pipelineResp_getRq[16] &&
	      IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2627) ;
  assign cache_pipeline_first__581_BITS_516_TO_513_583__ETC___d3287 =
	     cache_pipeline_first__581_BITS_516_TO_513_583__ETC___d2588 &&
	     !cache_cRqMshr$pipelineResp_getRq[16] &&
	     IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2627 &&
	     NOT_IF_cache_pipeline_first__581_BITS_584_TO_5_ETC___d3191 ;
  assign cache_pipeline_first__581_BITS_516_TO_513_583__ETC___d3295 =
	     cache_pipeline_first__581_BITS_516_TO_513_583__ETC___d2588 &&
	     !cache_cRqMshr$pipelineResp_getRq[16] &&
	     IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d3156 &&
	     cache_cRqMshr$pipelineResp_getSlot[12] ;
  assign cache_pipeline_first__581_BITS_519_TO_518_594__ETC___d2598 =
	     cache_pipeline$first[519:518] <=
	     IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2597 ;
  assign cache_pipeline_first__581_BITS_519_TO_518_594__ETC___d2618 =
	     cache_pipeline$first[519:518] <=
	     cache_cRqMshr$pipelineResp_getRq[87:86] ;
  assign cache_pipeline_first__581_BITS_519_TO_518_594__ETC___d3126 =
	     cache_pipeline_first__581_BITS_519_TO_518_594__ETC___d2598 &&
	     cache_pipeline_first__581_BITS_521_TO_520_600__ETC___d2601 &&
	     cache_pipeline_first__581_BITS_523_TO_522_603__ETC___d2604 &&
	     cache_cRqMshr$pipelineResp_getRq[85:84] == 2'd3 ;
  assign cache_pipeline_first__581_BITS_519_TO_518_594__ETC___d3136 =
	     cache_pipeline_first__581_BITS_519_TO_518_594__ETC___d2598 &&
	     cache_pipeline_first__581_BITS_521_TO_520_600__ETC___d2601 &&
	     cache_pipeline_first__581_BITS_523_TO_522_603__ETC___d2604 &&
	     cache_cRqMshr$pipelineResp_getRq[85:84] != 2'd3 ;
  assign cache_pipeline_first__581_BITS_519_TO_518_594__ETC___d3192 =
	     cache_pipeline_first__581_BITS_519_TO_518_594__ETC___d2598 &&
	     cache_pipeline_first__581_BITS_521_TO_520_600__ETC___d2601 &&
	     cache_pipeline_first__581_BITS_523_TO_522_603__ETC___d2604 &&
	     NOT_IF_cache_pipeline_first__581_BITS_584_TO_5_ETC___d3191 ;
  assign cache_pipeline_first__581_BITS_519_TO_518_594__ETC___d3196 =
	     cache_pipeline_first__581_BITS_519_TO_518_594__ETC___d2598 &&
	     cache_pipeline_first__581_BITS_521_TO_520_600__ETC___d2601 &&
	     cache_pipeline_first__581_BITS_523_TO_522_603__ETC___d2604 &&
	     (!cache_pipeline_first__581_BITS_573_TO_526_644__ETC___d2646 ||
	      cache_pipeline$first[525:524] == 2'd0) ;
  assign cache_pipeline_first__581_BITS_519_TO_518_594__ETC___d3265 =
	     cache_pipeline_first__581_BITS_519_TO_518_594__ETC___d2598 &&
	     cache_pipeline_first__581_BITS_521_TO_520_600__ETC___d2601 &&
	     cache_pipeline_first__581_BITS_523_TO_522_603__ETC___d2604 &&
	     NOT_cache_cRqMshr_pipelineResp_getRq_IF_cache__ETC___d3264 ;
  assign cache_pipeline_first__581_BITS_519_TO_518_594__ETC___d3271 =
	     cache_pipeline_first__581_BITS_519_TO_518_594__ETC___d2598 &&
	     cache_pipeline_first__581_BITS_521_TO_520_600__ETC___d2601 &&
	     cache_pipeline_first__581_BITS_523_TO_522_603__ETC___d2604 &&
	     cache_cRqMshr$pipelineResp_getData[512] !=
	     (cache_cRqMshr$pipelineResp_getRq[17] ||
	      cache_cRqMshr$pipelineResp_getRq[18] ||
	      cache_cRqMshr$pipelineResp_getRq[19] ||
	      cache_cRqMshr$pipelineResp_getRq[20] ||
	      cache_cRqMshr$pipelineResp_getRq[21] ||
	      cache_cRqMshr$pipelineResp_getRq[22] ||
	      cache_cRqMshr$pipelineResp_getRq[23] ||
	      cache_cRqMshr$pipelineResp_getRq[24] ||
	      cache_cRqMshr$pipelineResp_getRq[25] ||
	      cache_cRqMshr$pipelineResp_getRq[26] ||
	      cache_cRqMshr$pipelineResp_getRq[27] ||
	      cache_cRqMshr$pipelineResp_getRq[28] ||
	      cache_cRqMshr$pipelineResp_getRq[29] ||
	      cache_cRqMshr$pipelineResp_getRq[30] ||
	      cache_cRqMshr$pipelineResp_getRq[31] ||
	      cache_cRqMshr$pipelineResp_getRq[32] ||
	      cache_cRqMshr$pipelineResp_getRq[33] ||
	      cache_cRqMshr$pipelineResp_getRq[34] ||
	      cache_cRqMshr$pipelineResp_getRq[35] ||
	      cache_cRqMshr$pipelineResp_getRq[36] ||
	      cache_cRqMshr$pipelineResp_getRq[37] ||
	      cache_cRqMshr$pipelineResp_getRq[38] ||
	      cache_cRqMshr$pipelineResp_getRq[39] ||
	      cache_cRqMshr$pipelineResp_getRq[40] ||
	      cache_cRqMshr$pipelineResp_getRq[41] ||
	      cache_cRqMshr$pipelineResp_getRq[42] ||
	      cache_cRqMshr$pipelineResp_getRq[43] ||
	      cache_cRqMshr$pipelineResp_getRq[44] ||
	      cache_cRqMshr$pipelineResp_getRq[45] ||
	      cache_cRqMshr$pipelineResp_getRq[46] ||
	      cache_cRqMshr$pipelineResp_getRq[47] ||
	      cache_cRqMshr$pipelineResp_getRq[48] ||
	      cache_cRqMshr$pipelineResp_getRq[49] ||
	      cache_cRqMshr$pipelineResp_getRq[50] ||
	      cache_cRqMshr$pipelineResp_getRq[51] ||
	      cache_cRqMshr$pipelineResp_getRq[52] ||
	      cache_cRqMshr$pipelineResp_getRq[53] ||
	      cache_cRqMshr$pipelineResp_getRq[54] ||
	      cache_cRqMshr$pipelineResp_getRq[55] ||
	      cache_cRqMshr$pipelineResp_getRq[56] ||
	      cache_cRqMshr$pipelineResp_getRq[57] ||
	      cache_cRqMshr$pipelineResp_getRq[58] ||
	      cache_cRqMshr$pipelineResp_getRq[59] ||
	      cache_cRqMshr$pipelineResp_getRq[60] ||
	      cache_cRqMshr$pipelineResp_getRq[61] ||
	      cache_cRqMshr$pipelineResp_getRq[62] ||
	      cache_cRqMshr$pipelineResp_getRq[63] ||
	      cache_cRqMshr$pipelineResp_getRq[64] ||
	      cache_cRqMshr$pipelineResp_getRq[65] ||
	      cache_cRqMshr$pipelineResp_getRq[66] ||
	      cache_cRqMshr$pipelineResp_getRq[67] ||
	      cache_cRqMshr$pipelineResp_getRq[68] ||
	      cache_cRqMshr$pipelineResp_getRq[69] ||
	      cache_cRqMshr$pipelineResp_getRq[70] ||
	      cache_cRqMshr$pipelineResp_getRq[71] ||
	      cache_cRqMshr$pipelineResp_getRq[72] ||
	      cache_cRqMshr$pipelineResp_getRq[73] ||
	      cache_cRqMshr$pipelineResp_getRq[74] ||
	      cache_cRqMshr$pipelineResp_getRq[75] ||
	      cache_cRqMshr$pipelineResp_getRq[76] ||
	      cache_cRqMshr$pipelineResp_getRq[77] ||
	      cache_cRqMshr$pipelineResp_getRq[78] ||
	      cache_cRqMshr$pipelineResp_getRq[79] ||
	      cache_cRqMshr$pipelineResp_getRq[80]) ;
  assign cache_pipeline_first__581_BITS_521_TO_520_600__ETC___d2601 =
	     cache_pipeline$first[521:520] <=
	     IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2597 ;
  assign cache_pipeline_first__581_BITS_521_TO_520_600__ETC___d2621 =
	     cache_pipeline$first[521:520] <=
	     cache_cRqMshr$pipelineResp_getRq[87:86] ;
  assign cache_pipeline_first__581_BITS_523_TO_522_603__ETC___d2604 =
	     cache_pipeline$first[523:522] <=
	     IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2597 ;
  assign cache_pipeline_first__581_BITS_523_TO_522_603__ETC___d2624 =
	     cache_pipeline$first[523:522] <=
	     cache_cRqMshr$pipelineResp_getRq[87:86] ;
  assign cache_pipeline_first__581_BITS_573_TO_526_644__ETC___d2646 =
	     cache_pipeline$first[573:526] ==
	     cache_cRqMshr$pipelineResp_getRq[151:104] ;
  assign cache_pipeline_first__581_BIT_517_582_AND_NOT__ETC___d3820 =
	     cache_pipeline$first[517] && !cache_pipeline$first[512] &&
	     IF_SEL_ARR_cache_cRqMshr_pipelineResp_getSlot__ETC___d3484 &&
	     cache_cRqMshr$pipelineResp_getRq[16] &&
	     cache_cRqMshr$pipelineResp_getRq[85:84] == 2'd3 ;
  assign cache_pipeline_first__581_BIT_517_582_AND_NOT__ETC___d3824 =
	     cache_pipeline$first[517] && !cache_pipeline$first[512] &&
	     IF_SEL_ARR_cache_cRqMshr_pipelineResp_getSlot__ETC___d3484 &&
	     cache_cRqMshr$pipelineResp_getRq[16] &&
	     cache_cRqMshr$pipelineResp_getRq[85:84] != 2'd3 ;
  assign cache_pipeline_first__581_BIT_517_582_AND_cach_ETC___d3129 =
	     cache_pipeline$first[517] &&
	     cache_pipeline_first__581_BITS_516_TO_513_583__ETC___d2588 &&
	     cache_cRqMshr$pipelineResp_getRq[16] &&
	     cache_pipeline_first__581_BITS_519_TO_518_594__ETC___d3126 ;
  assign cache_pipeline_first__581_BIT_517_582_AND_cach_ETC___d3139 =
	     cache_pipeline$first[517] &&
	     cache_pipeline_first__581_BITS_516_TO_513_583__ETC___d2588 &&
	     cache_cRqMshr$pipelineResp_getRq[16] &&
	     cache_pipeline_first__581_BITS_519_TO_518_594__ETC___d3136 ;
  assign cache_pipeline_first__581_BIT_517_582_AND_cach_ETC___d3146 =
	     cache_pipeline$first[517] &&
	     cache_pipeline_first__581_BITS_516_TO_513_583__ETC___d2588 &&
	     !cache_cRqMshr$pipelineResp_getRq[16] &&
	     IF_cache_cRqMshr_pipelineResp_getRq_IF_cache_p_ETC___d2627 ;
  assign cache_pipeline_first__581_BIT_517_582_AND_cach_ETC___d3195 =
	     cache_pipeline$first[517] &&
	     cache_pipeline_first__581_BITS_516_TO_513_583__ETC___d2588 &&
	     cache_cRqMshr$pipelineResp_getRq[16] &&
	     cache_pipeline_first__581_BITS_519_TO_518_594__ETC___d3192 ;
  assign cache_pipeline_first__581_BIT_517_582_AND_cach_ETC___d3199 =
	     cache_pipeline$first[517] &&
	     cache_pipeline_first__581_BITS_516_TO_513_583__ETC___d2588 &&
	     cache_cRqMshr$pipelineResp_getRq[16] &&
	     cache_pipeline_first__581_BITS_519_TO_518_594__ETC___d3196 ;
  assign cache_pipeline_first__581_BIT_517_582_AND_cach_ETC___d3268 =
	     cache_pipeline$first[517] &&
	     cache_pipeline_first__581_BITS_516_TO_513_583__ETC___d2588 &&
	     cache_cRqMshr$pipelineResp_getRq[16] &&
	     cache_pipeline_first__581_BITS_519_TO_518_594__ETC___d3265 ;
  assign cache_pipeline_first__581_BIT_517_582_AND_cach_ETC___d3274 =
	     cache_pipeline$first[517] &&
	     cache_pipeline_first__581_BITS_516_TO_513_583__ETC___d2588 &&
	     cache_cRqMshr$pipelineResp_getRq[16] &&
	     cache_pipeline_first__581_BITS_519_TO_518_594__ETC___d3271 ;
  assign cache_pipeline_first__581_BIT_517_582_AND_cach_ETC___d3278 =
	     cache_pipeline$first[517] &&
	     cache_pipeline_first__581_BITS_516_TO_513_583__ETC___d2588 &&
	     cache_cRqMshr$pipelineResp_getRq[16] &&
	     NOT_cache_pipeline_first__581_BITS_519_TO_518__ETC___d3275 ;
  assign cache_pipeline_first__581_BIT_517_582_AND_cach_ETC___d3284 =
	     cache_pipeline$first[517] &&
	     cache_pipeline_first__581_BITS_516_TO_513_583__ETC___d2588 &&
	     cache_cRqMshr$pipelineResp_getRq[16] &&
	     NOT_cache_pipeline_first__581_BITS_519_TO_518__ETC___d3281 ;
  assign cache_rqFromCQ_enqReq_dummy2_2_read__4_AND_IF__ETC___d65 =
	     cache_rqFromCQ_enqReq_dummy2_2$Q_OUT &&
	     IF_cache_rqFromCQ_enqReq_lat_1_whas_THEN_cache_ETC___d39 ||
	     (!cache_rqFromCQ_deqReq_dummy2_2$Q_OUT ||
	      !WILL_FIRE_RL_cache_cRqTransfer_new_child &&
	      !cache_rqFromCQ_deqReq_rl) &&
	     cache_rqFromCQ_full ;
  assign cache_rqFromDmaQ_enqReq_dummy2_2_read__40_AND__ETC___d371 =
	     cache_rqFromDmaQ_enqReq_dummy2_2$Q_OUT &&
	     IF_cache_rqFromDmaQ_enqReq_lat_1_whas__09_THEN_ETC___d345 ||
	     (!cache_rqFromDmaQ_deqReq_dummy2_2$Q_OUT ||
	      !WILL_FIRE_RL_cache_cRqTransfer_new_dma &&
	      !cache_rqFromDmaQ_deqReq_rl) &&
	     cache_rqFromDmaQ_full ;
  assign cache_rsFromCQ_enqReq_dummy2_2_read__26_AND_IF_ETC___d157 =
	     cache_rsFromCQ_enqReq_dummy2_2$Q_OUT &&
	     IF_cache_rsFromCQ_enqReq_lat_1_whas__5_THEN_ca_ETC___d131 ||
	     (!cache_rsFromCQ_deqReq_dummy2_2$Q_OUT ||
	      !WILL_FIRE_RL_cache_cRsTransfer && !cache_rsFromCQ_deqReq_rl) &&
	     cache_rsFromCQ_full ;
  assign cache_rsFromMQ_enqReq_dummy2_2_read__41_AND_IF_ETC___d772 =
	     cache_rsFromMQ_enqReq_dummy2_2$Q_OUT &&
	     IF_cache_rsFromMQ_enqReq_lat_1_whas__10_THEN_c_ETC___d746 ||
	     (!cache_rsFromMQ_deqReq_dummy2_2$Q_OUT ||
	      !cache_rsFromMQ_deqReq_lat_0$whas &&
	      !cache_rsFromMQ_deqReq_rl) &&
	     cache_rsFromMQ_full ;
  assign cache_rsLdToDmaQ_enqReq_dummy2_2_read__31_AND__ETC___d462 =
	     cache_rsLdToDmaQ_enqReq_dummy2_2$Q_OUT &&
	     IF_cache_rsLdToDmaQ_enqReq_lat_1_whas__00_THEN_ETC___d436 ||
	     (!cache_rsLdToDmaQ_deqReq_dummy2_2$Q_OUT ||
	      !EN_dma_respLd_deq && !cache_rsLdToDmaQ_deqReq_rl) &&
	     cache_rsLdToDmaQ_full ;
  assign cache_rsStToDmaQ_enqReq_dummy2_2_read__22_AND__ETC___d553 =
	     cache_rsStToDmaQ_enqReq_dummy2_2$Q_OUT &&
	     IF_cache_rsStToDmaQ_enqReq_lat_1_whas__91_THEN_ETC___d527 ||
	     (!cache_rsStToDmaQ_deqReq_dummy2_2$Q_OUT ||
	      !EN_dma_respSt_deq && !cache_rsStToDmaQ_deqReq_rl) &&
	     cache_rsStToDmaQ_full ;
  assign cache_rsToCIndexQ_enqReq_dummy2_2_read__51_AND_ETC___d987 =
	     cache_rsToCIndexQ_enqReq_dummy2_2$Q_OUT &&
	     IF_cache_rsToCIndexQ_enqReq_lat_1_whas__24_THE_ETC___d956 ||
	     (!cache_rsToCIndexQ_deqReq_dummy2_2$Q_OUT ||
	      !WILL_FIRE_RL_cache_sendRsToC &&
	      !cache_rsToCIndexQ_deqReq_rl) &&
	     cache_rsToCIndexQ_full ;
  assign cache_toCQ_enqReq_dummy2_2_read__53_AND_IF_cac_ETC___d279 =
	     cache_toCQ_enqReq_dummy2_2$Q_OUT &&
	     IF_cache_toCQ_enqReq_lat_1_whas__87_THEN_cache_ETC___d196 ||
	     (!cache_toCQ_deqReq_dummy2_2$Q_OUT ||
	      !EN_to_child_toC_deq && !cache_toCQ_deqReq_rl) &&
	     cache_toCQ_full ;
  assign cache_toMQ_enqReq_dummy2_2_read__54_AND_IF_cac_ETC___d680 =
	     cache_toMQ_enqReq_dummy2_2$Q_OUT &&
	     IF_cache_toMQ_enqReq_lat_1_whas__88_THEN_cache_ETC___d597 ||
	     (!cache_toMQ_deqReq_dummy2_2$Q_OUT ||
	      !EN_to_mem_toM_deq && !cache_toMQ_deqReq_rl) &&
	     cache_toMQ_full ;
  assign child__h313067 =
	     (cache_cRqMshr$sendRqToC_getSlot[3:2] != 2'd1 &&
	      cache_cRqMshr$sendRqToC_getSlot[7:6] != 2'd1) ?
	       2'd2 :
	       ((cache_cRqMshr$sendRqToC_getSlot[3:2] == 2'd1) ?
		  2'd0 :
		  2'd1) ;
  assign next_deqP___1__h119479 = cache_rqFromDmaQ_deqP + 1'd1 ;
  assign next_deqP___1__h135572 = cache_rsLdToDmaQ_deqP + 1'd1 ;
  assign next_deqP___1__h143074 = cache_rsStToDmaQ_deqP + 1'd1 ;
  assign next_deqP___1__h208858 = cache_toMQ_deqP + 1'd1 ;
  assign next_deqP___1__h225353 = cache_rsFromMQ_deqP + 1'd1 ;
  assign next_deqP___1__h22634 = cache_rsFromCQ_deqP + 1'd1 ;
  assign next_deqP___1__h234850 =
	     (cache_cRqRetryIndexQ_deqP == 4'd15) ?
	       4'd0 :
	       cache_cRqRetryIndexQ_deqP + 4'd1 ;
  assign next_deqP___1__h246325 =
	     (cache_rsToCIndexQ_deqP == 4'd15) ?
	       4'd0 :
	       cache_rsToCIndexQ_deqP + 4'd1 ;
  assign next_deqP___1__h38327 = cache_toCQ_deqP + 1'd1 ;
  assign next_deqP___1__h7552 = cache_rqFromCQ_deqP + 1'd1 ;
  assign perfReqQ_enqReq_dummy2_2_read__870_AND_IF_perf_ETC___d3887 =
	     perfReqQ_enqReq_dummy2_2$Q_OUT &&
	     IF_perfReqQ_enqReq_lat_1_whas__839_THEN_perfRe_ETC___d3875 ||
	     (!perfReqQ_deqReq_dummy2_2$Q_OUT ||
	      !EN_perf_resp && !perfReqQ_deqReq_rl) &&
	     perfReqQ_full ;
  assign pipeOutCRqIdx__h314276 =
	     (cache_pipeline$first[584:583] == 2'd0) ?
	       cache_pipeline$first[582:579] :
	       (cache_pipeline$first[517] ?
		  cache_pipeline$first[516:513] :
		  4'd0) ;
  assign rqAddr__h313360 =
	     (cache_cRqMshr$sendRqToC_getState == 3'd3) ?
	       cache_cRqMshr$sendRqToC_getRq[151:88] :
	       { cache_cRqMshr$sendRqToC_getSlot[60:13],
		 cache_cRqMshr$sendRqToC_getRq[103:88] } ;
  assign v__h129259 =
	     (cache_rsLdToDmaQ_enqReq_dummy2_2$Q_OUT &&
	      IF_cache_rsLdToDmaQ_enqReq_lat_1_whas__00_THEN_ETC___d436) ?
	       v__h129542 :
	       cache_rsLdToDmaQ_enqP ;
  assign v__h129542 = cache_rsLdToDmaQ_enqP + 1'd1 ;
  assign v__h142239 =
	     (cache_rsStToDmaQ_enqReq_dummy2_2$Q_OUT &&
	      IF_cache_rsStToDmaQ_enqReq_lat_1_whas__91_THEN_ETC___d527) ?
	       v__h142522 :
	       cache_rsStToDmaQ_enqP ;
  assign v__h142522 = cache_rsStToDmaQ_enqP + 1'd1 ;
  assign v__h16641 =
	     (cache_rsFromCQ_enqReq_dummy2_2$Q_OUT &&
	      IF_cache_rsFromCQ_enqReq_lat_1_whas__5_THEN_ca_ETC___d131) ?
	       v__h16924 :
	       cache_rsFromCQ_enqP ;
  assign v__h168573 =
	     (cache_toMQ_enqReq_dummy2_2$Q_OUT &&
	      IF_cache_toMQ_enqReq_lat_1_whas__88_THEN_cache_ETC___d597) ?
	       v__h168856 :
	       cache_toMQ_enqP ;
  assign v__h168856 = cache_toMQ_enqP + 1'd1 ;
  assign v__h16924 = cache_rsFromCQ_enqP + 1'd1 ;
  assign v__h218716 =
	     (cache_rsFromMQ_enqReq_dummy2_2$Q_OUT &&
	      IF_cache_rsFromMQ_enqReq_lat_1_whas__10_THEN_c_ETC___d746) ?
	       v__h218999 :
	       cache_rsFromMQ_enqP ;
  assign v__h218999 = cache_rsFromMQ_enqP + 1'd1 ;
  assign v__h232953 =
	     (cache_cRqRetryIndexQ_enqReq_dummy2_2$Q_OUT &&
	      IF_cache_cRqRetryIndexQ_enqReq_lat_1_whas__01__ETC___d833) ?
	       v__h233236 :
	       cache_cRqRetryIndexQ_enqP ;
  assign v__h233236 =
	     (cache_cRqRetryIndexQ_enqP == 4'd15) ?
	       4'd0 :
	       cache_cRqRetryIndexQ_enqP + 4'd1 ;
  assign v__h242396 =
	     (cache_rsToCIndexQ_enqReq_dummy2_2$Q_OUT &&
	      IF_cache_rsToCIndexQ_enqReq_lat_1_whas__24_THE_ETC___d956) ?
	       v__h242679 :
	       cache_rsToCIndexQ_enqP ;
  assign v__h242679 =
	     (cache_rsToCIndexQ_enqP == 4'd15) ?
	       4'd0 :
	       cache_rsToCIndexQ_enqP + 4'd1 ;
  assign v__h31944 =
	     (cache_toCQ_enqReq_dummy2_2$Q_OUT &&
	      IF_cache_toCQ_enqReq_lat_1_whas__87_THEN_cache_ETC___d196) ?
	       v__h32227 :
	       cache_toCQ_enqP ;
  assign v__h32227 = cache_toCQ_enqP + 1'd1 ;
  assign v__h6037 =
	     (cache_rqFromCQ_enqReq_dummy2_2$Q_OUT &&
	      IF_cache_rqFromCQ_enqReq_lat_1_whas_THEN_cache_ETC___d39) ?
	       v__h6320 :
	       cache_rqFromCQ_enqP ;
  assign v__h6320 = cache_rqFromCQ_enqP + 1'd1 ;
  assign v__h72082 =
	     (cache_rqFromDmaQ_enqReq_dummy2_2$Q_OUT &&
	      IF_cache_rqFromDmaQ_enqReq_lat_1_whas__09_THEN_ETC___d345) ?
	       v__h72365 :
	       cache_rqFromDmaQ_enqP ;
  assign v__h72365 = cache_rqFromDmaQ_enqP + 1'd1 ;
  always@(cache_rqFromCQ_deqP or
	  cache_rqFromCQ_data_0 or cache_rqFromCQ_data_1)
  begin
    case (cache_rqFromCQ_deqP)
      1'd0: x__h257564 = cache_rqFromCQ_data_0[4:2];
      1'd1: x__h257564 = cache_rqFromCQ_data_1[4:2];
    endcase
  end
  always@(cache_rqFromCQ_deqP or
	  cache_rqFromCQ_data_0 or cache_rqFromCQ_data_1)
  begin
    case (cache_rqFromCQ_deqP)
      1'd0: addr__h257616 = cache_rqFromCQ_data_0[73:10];
      1'd1: addr__h257616 = cache_rqFromCQ_data_1[73:10];
    endcase
  end
  always@(cache_cRqRetryIndexQ_deqP or
	  cache_cRqRetryIndexQ_data_0 or
	  cache_cRqRetryIndexQ_data_1 or
	  cache_cRqRetryIndexQ_data_2 or
	  cache_cRqRetryIndexQ_data_3 or
	  cache_cRqRetryIndexQ_data_4 or
	  cache_cRqRetryIndexQ_data_5 or
	  cache_cRqRetryIndexQ_data_6 or
	  cache_cRqRetryIndexQ_data_7 or
	  cache_cRqRetryIndexQ_data_8 or
	  cache_cRqRetryIndexQ_data_9 or
	  cache_cRqRetryIndexQ_data_10 or
	  cache_cRqRetryIndexQ_data_11 or
	  cache_cRqRetryIndexQ_data_12 or
	  cache_cRqRetryIndexQ_data_13 or
	  cache_cRqRetryIndexQ_data_14 or cache_cRqRetryIndexQ_data_15)
  begin
    case (cache_cRqRetryIndexQ_deqP)
      4'd0: x__h248737 = cache_cRqRetryIndexQ_data_0;
      4'd1: x__h248737 = cache_cRqRetryIndexQ_data_1;
      4'd2: x__h248737 = cache_cRqRetryIndexQ_data_2;
      4'd3: x__h248737 = cache_cRqRetryIndexQ_data_3;
      4'd4: x__h248737 = cache_cRqRetryIndexQ_data_4;
      4'd5: x__h248737 = cache_cRqRetryIndexQ_data_5;
      4'd6: x__h248737 = cache_cRqRetryIndexQ_data_6;
      4'd7: x__h248737 = cache_cRqRetryIndexQ_data_7;
      4'd8: x__h248737 = cache_cRqRetryIndexQ_data_8;
      4'd9: x__h248737 = cache_cRqRetryIndexQ_data_9;
      4'd10: x__h248737 = cache_cRqRetryIndexQ_data_10;
      4'd11: x__h248737 = cache_cRqRetryIndexQ_data_11;
      4'd12: x__h248737 = cache_cRqRetryIndexQ_data_12;
      4'd13: x__h248737 = cache_cRqRetryIndexQ_data_13;
      4'd14: x__h248737 = cache_cRqRetryIndexQ_data_14;
      4'd15: x__h248737 = cache_cRqRetryIndexQ_data_15;
    endcase
  end
  always@(cache_rqFromCQ_deqP or
	  cache_rqFromCQ_data_0 or cache_rqFromCQ_data_1)
  begin
    case (cache_rqFromCQ_deqP)
      1'd0: x__h249082 = cache_rqFromCQ_data_0[1:0];
      1'd1: x__h249082 = cache_rqFromCQ_data_1[1:0];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0: addr__h273361 = cache_rqFromDmaQ_data_0[655:592];
      1'd1: addr__h273361 = cache_rqFromDmaQ_data_1[655:592];
    endcase
  end
  always@(cache_toCQ_deqP or cache_toCQ_data_0 or cache_toCQ_data_1)
  begin
    case (cache_toCQ_deqP)
      1'd0: x__h444361 = cache_toCQ_data_0[1:0];
      1'd1: x__h444361 = cache_toCQ_data_1[1:0];
    endcase
  end
  always@(cache_toCQ_deqP or cache_toCQ_data_0 or cache_toCQ_data_1)
  begin
    case (cache_toCQ_deqP)
      1'd0: x__h444405 = cache_toCQ_data_0[517:516];
      1'd1: x__h444405 = cache_toCQ_data_1[517:516];
    endcase
  end
  always@(cache_toCQ_deqP or cache_toCQ_data_0 or cache_toCQ_data_1)
  begin
    case (cache_toCQ_deqP)
      1'd0: x__h445950 = cache_toCQ_data_0[2:0];
      1'd1: x__h445950 = cache_toCQ_data_1[2:0];
    endcase
  end
  always@(cache_toMQ_deqP or cache_toMQ_data_0 or cache_toMQ_data_1)
  begin
    case (cache_toMQ_deqP)
      1'd0: x__h456804 = cache_toMQ_data_0[3:0];
      1'd1: x__h456804 = cache_toMQ_data_1[3:0];
    endcase
  end
  always@(cache_rsLdToDmaQ_deqP or
	  cache_rsLdToDmaQ_data_0 or cache_rsLdToDmaQ_data_1)
  begin
    case (cache_rsLdToDmaQ_deqP)
      1'd0: x__h456399 = cache_rsLdToDmaQ_data_0[15:0];
      1'd1: x__h456399 = cache_rsLdToDmaQ_data_1[15:0];
    endcase
  end
  always@(cache_rsFromCQ_deqP or
	  cache_rsFromCQ_data_0 or cache_rsFromCQ_data_1)
  begin
    case (cache_rsFromCQ_deqP)
      1'd0: x__h275130 = cache_rsFromCQ_data_0[1:0];
      1'd1: x__h275130 = cache_rsFromCQ_data_1[1:0];
    endcase
  end
  always@(cache_rsFromMQ_deqP or
	  cache_rsFromMQ_data_0 or cache_rsFromMQ_data_1)
  begin
    case (cache_rsFromMQ_deqP)
      1'd0:
	  CASE_cache_rsFromMQ_deqP_0_cache_rsFromMQ_data_ETC__q1 =
	      cache_rsFromMQ_data_0[516:453];
      1'd1:
	  CASE_cache_rsFromMQ_deqP_0_cache_rsFromMQ_data_ETC__q1 =
	      cache_rsFromMQ_data_1[516:453];
    endcase
  end
  always@(cache_rsFromMQ_deqP or
	  cache_rsFromMQ_data_0 or cache_rsFromMQ_data_1)
  begin
    case (cache_rsFromMQ_deqP)
      1'd0:
	  CASE_cache_rsFromMQ_deqP_0_cache_rsFromMQ_data_ETC__q2 =
	      cache_rsFromMQ_data_0[452:389];
      1'd1:
	  CASE_cache_rsFromMQ_deqP_0_cache_rsFromMQ_data_ETC__q2 =
	      cache_rsFromMQ_data_1[452:389];
    endcase
  end
  always@(cache_rsFromMQ_deqP or
	  cache_rsFromMQ_data_0 or cache_rsFromMQ_data_1)
  begin
    case (cache_rsFromMQ_deqP)
      1'd0:
	  CASE_cache_rsFromMQ_deqP_0_cache_rsFromMQ_data_ETC__q3 =
	      cache_rsFromMQ_data_0[388:325];
      1'd1:
	  CASE_cache_rsFromMQ_deqP_0_cache_rsFromMQ_data_ETC__q3 =
	      cache_rsFromMQ_data_1[388:325];
    endcase
  end
  always@(cache_rsFromMQ_deqP or
	  cache_rsFromMQ_data_0 or cache_rsFromMQ_data_1)
  begin
    case (cache_rsFromMQ_deqP)
      1'd0:
	  CASE_cache_rsFromMQ_deqP_0_cache_rsFromMQ_data_ETC__q4 =
	      cache_rsFromMQ_data_0[324:261];
      1'd1:
	  CASE_cache_rsFromMQ_deqP_0_cache_rsFromMQ_data_ETC__q4 =
	      cache_rsFromMQ_data_1[324:261];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q5 =
	      !cache_rqFromDmaQ_data_0[589];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q5 =
	      !cache_rqFromDmaQ_data_1[589];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q6 =
	      !cache_rqFromDmaQ_data_0[590];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q6 =
	      !cache_rqFromDmaQ_data_1[590];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q7 =
	      !cache_rqFromDmaQ_data_0[591];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q7 =
	      !cache_rqFromDmaQ_data_1[591];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q8 =
	      !cache_rqFromDmaQ_data_0[587];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q8 =
	      !cache_rqFromDmaQ_data_1[587];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q9 =
	      !cache_rqFromDmaQ_data_0[588];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q9 =
	      !cache_rqFromDmaQ_data_1[588];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q10 =
	      !cache_rqFromDmaQ_data_0[585];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q10 =
	      !cache_rqFromDmaQ_data_1[585];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q11 =
	      !cache_rqFromDmaQ_data_0[586];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q11 =
	      !cache_rqFromDmaQ_data_1[586];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q12 =
	      !cache_rqFromDmaQ_data_0[583];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q12 =
	      !cache_rqFromDmaQ_data_1[583];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q13 =
	      !cache_rqFromDmaQ_data_0[584];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q13 =
	      !cache_rqFromDmaQ_data_1[584];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q14 =
	      !cache_rqFromDmaQ_data_0[581];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q14 =
	      !cache_rqFromDmaQ_data_1[581];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q15 =
	      !cache_rqFromDmaQ_data_0[582];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q15 =
	      !cache_rqFromDmaQ_data_1[582];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q16 =
	      !cache_rqFromDmaQ_data_0[579];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q16 =
	      !cache_rqFromDmaQ_data_1[579];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q17 =
	      !cache_rqFromDmaQ_data_0[580];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q17 =
	      !cache_rqFromDmaQ_data_1[580];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q18 =
	      !cache_rqFromDmaQ_data_0[577];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q18 =
	      !cache_rqFromDmaQ_data_1[577];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q19 =
	      !cache_rqFromDmaQ_data_0[578];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q19 =
	      !cache_rqFromDmaQ_data_1[578];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q20 =
	      !cache_rqFromDmaQ_data_0[575];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q20 =
	      !cache_rqFromDmaQ_data_1[575];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q21 =
	      !cache_rqFromDmaQ_data_0[576];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q21 =
	      !cache_rqFromDmaQ_data_1[576];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q22 =
	      !cache_rqFromDmaQ_data_0[573];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q22 =
	      !cache_rqFromDmaQ_data_1[573];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q23 =
	      !cache_rqFromDmaQ_data_0[574];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q23 =
	      !cache_rqFromDmaQ_data_1[574];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q24 =
	      !cache_rqFromDmaQ_data_0[571];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q24 =
	      !cache_rqFromDmaQ_data_1[571];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q25 =
	      !cache_rqFromDmaQ_data_0[572];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q25 =
	      !cache_rqFromDmaQ_data_1[572];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q26 =
	      !cache_rqFromDmaQ_data_0[569];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q26 =
	      !cache_rqFromDmaQ_data_1[569];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q27 =
	      !cache_rqFromDmaQ_data_0[570];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q27 =
	      !cache_rqFromDmaQ_data_1[570];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q28 =
	      !cache_rqFromDmaQ_data_0[567];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q28 =
	      !cache_rqFromDmaQ_data_1[567];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q29 =
	      !cache_rqFromDmaQ_data_0[568];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q29 =
	      !cache_rqFromDmaQ_data_1[568];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q30 =
	      !cache_rqFromDmaQ_data_0[565];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q30 =
	      !cache_rqFromDmaQ_data_1[565];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q31 =
	      !cache_rqFromDmaQ_data_0[566];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q31 =
	      !cache_rqFromDmaQ_data_1[566];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q32 =
	      !cache_rqFromDmaQ_data_0[563];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q32 =
	      !cache_rqFromDmaQ_data_1[563];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q33 =
	      !cache_rqFromDmaQ_data_0[564];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q33 =
	      !cache_rqFromDmaQ_data_1[564];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q34 =
	      !cache_rqFromDmaQ_data_0[561];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q34 =
	      !cache_rqFromDmaQ_data_1[561];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q35 =
	      !cache_rqFromDmaQ_data_0[562];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q35 =
	      !cache_rqFromDmaQ_data_1[562];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q36 =
	      !cache_rqFromDmaQ_data_0[559];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q36 =
	      !cache_rqFromDmaQ_data_1[559];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q37 =
	      !cache_rqFromDmaQ_data_0[560];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q37 =
	      !cache_rqFromDmaQ_data_1[560];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q38 =
	      !cache_rqFromDmaQ_data_0[557];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q38 =
	      !cache_rqFromDmaQ_data_1[557];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q39 =
	      !cache_rqFromDmaQ_data_0[558];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q39 =
	      !cache_rqFromDmaQ_data_1[558];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q40 =
	      !cache_rqFromDmaQ_data_0[555];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q40 =
	      !cache_rqFromDmaQ_data_1[555];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q41 =
	      !cache_rqFromDmaQ_data_0[556];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q41 =
	      !cache_rqFromDmaQ_data_1[556];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q42 =
	      !cache_rqFromDmaQ_data_0[553];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q42 =
	      !cache_rqFromDmaQ_data_1[553];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q43 =
	      !cache_rqFromDmaQ_data_0[554];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q43 =
	      !cache_rqFromDmaQ_data_1[554];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q44 =
	      !cache_rqFromDmaQ_data_0[551];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q44 =
	      !cache_rqFromDmaQ_data_1[551];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q45 =
	      !cache_rqFromDmaQ_data_0[552];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q45 =
	      !cache_rqFromDmaQ_data_1[552];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q46 =
	      !cache_rqFromDmaQ_data_0[549];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q46 =
	      !cache_rqFromDmaQ_data_1[549];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q47 =
	      !cache_rqFromDmaQ_data_0[550];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q47 =
	      !cache_rqFromDmaQ_data_1[550];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q48 =
	      !cache_rqFromDmaQ_data_0[547];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q48 =
	      !cache_rqFromDmaQ_data_1[547];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q49 =
	      !cache_rqFromDmaQ_data_0[548];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q49 =
	      !cache_rqFromDmaQ_data_1[548];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q50 =
	      !cache_rqFromDmaQ_data_0[545];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q50 =
	      !cache_rqFromDmaQ_data_1[545];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q51 =
	      !cache_rqFromDmaQ_data_0[546];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q51 =
	      !cache_rqFromDmaQ_data_1[546];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q52 =
	      !cache_rqFromDmaQ_data_0[543];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q52 =
	      !cache_rqFromDmaQ_data_1[543];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q53 =
	      !cache_rqFromDmaQ_data_0[544];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q53 =
	      !cache_rqFromDmaQ_data_1[544];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q54 =
	      !cache_rqFromDmaQ_data_0[541];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q54 =
	      !cache_rqFromDmaQ_data_1[541];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q55 =
	      !cache_rqFromDmaQ_data_0[542];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q55 =
	      !cache_rqFromDmaQ_data_1[542];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q56 =
	      !cache_rqFromDmaQ_data_0[539];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q56 =
	      !cache_rqFromDmaQ_data_1[539];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q57 =
	      !cache_rqFromDmaQ_data_0[540];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q57 =
	      !cache_rqFromDmaQ_data_1[540];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q58 =
	      !cache_rqFromDmaQ_data_0[537];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q58 =
	      !cache_rqFromDmaQ_data_1[537];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q59 =
	      !cache_rqFromDmaQ_data_0[538];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q59 =
	      !cache_rqFromDmaQ_data_1[538];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q60 =
	      !cache_rqFromDmaQ_data_0[535];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q60 =
	      !cache_rqFromDmaQ_data_1[535];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q61 =
	      !cache_rqFromDmaQ_data_0[536];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q61 =
	      !cache_rqFromDmaQ_data_1[536];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q62 =
	      !cache_rqFromDmaQ_data_0[533];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q62 =
	      !cache_rqFromDmaQ_data_1[533];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q63 =
	      !cache_rqFromDmaQ_data_0[534];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q63 =
	      !cache_rqFromDmaQ_data_1[534];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q64 =
	      !cache_rqFromDmaQ_data_0[531];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q64 =
	      !cache_rqFromDmaQ_data_1[531];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q65 =
	      !cache_rqFromDmaQ_data_0[532];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q65 =
	      !cache_rqFromDmaQ_data_1[532];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q66 =
	      !cache_rqFromDmaQ_data_0[529];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q66 =
	      !cache_rqFromDmaQ_data_1[529];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q67 =
	      !cache_rqFromDmaQ_data_0[530];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q67 =
	      !cache_rqFromDmaQ_data_1[530];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q68 =
	      !cache_rqFromDmaQ_data_0[528];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_NOT_cache_rqFromD_ETC__q68 =
	      !cache_rqFromDmaQ_data_1[528];
    endcase
  end
  always@(cache_rsFromCQ_deqP or
	  cache_rsFromCQ_data_0 or cache_rsFromCQ_data_1)
  begin
    case (cache_rsFromCQ_deqP)
      1'd0:
	  CASE_cache_rsFromCQ_deqP_0_cache_rsFromCQ_data_ETC__q69 =
	      cache_rsFromCQ_data_0[513:450];
      1'd1:
	  CASE_cache_rsFromCQ_deqP_0_cache_rsFromCQ_data_ETC__q69 =
	      cache_rsFromCQ_data_1[513:450];
    endcase
  end
  always@(cache_rsFromCQ_deqP or
	  cache_rsFromCQ_data_0 or cache_rsFromCQ_data_1)
  begin
    case (cache_rsFromCQ_deqP)
      1'd0:
	  CASE_cache_rsFromCQ_deqP_0_cache_rsFromCQ_data_ETC__q70 =
	      cache_rsFromCQ_data_0[449:386];
      1'd1:
	  CASE_cache_rsFromCQ_deqP_0_cache_rsFromCQ_data_ETC__q70 =
	      cache_rsFromCQ_data_1[449:386];
    endcase
  end
  always@(cache_rsFromCQ_deqP or
	  cache_rsFromCQ_data_0 or cache_rsFromCQ_data_1)
  begin
    case (cache_rsFromCQ_deqP)
      1'd0:
	  CASE_cache_rsFromCQ_deqP_0_cache_rsFromCQ_data_ETC__q71 =
	      cache_rsFromCQ_data_0[385:322];
      1'd1:
	  CASE_cache_rsFromCQ_deqP_0_cache_rsFromCQ_data_ETC__q71 =
	      cache_rsFromCQ_data_1[385:322];
    endcase
  end
  always@(cache_rsFromCQ_deqP or
	  cache_rsFromCQ_data_0 or cache_rsFromCQ_data_1)
  begin
    case (cache_rsFromCQ_deqP)
      1'd0:
	  CASE_cache_rsFromCQ_deqP_0_cache_rsFromCQ_data_ETC__q72 =
	      cache_rsFromCQ_data_0[321:258];
      1'd1:
	  CASE_cache_rsFromCQ_deqP_0_cache_rsFromCQ_data_ETC__q72 =
	      cache_rsFromCQ_data_1[321:258];
    endcase
  end
  always@(cache_rsFromMQ_deqP or
	  cache_rsFromMQ_data_0 or cache_rsFromMQ_data_1)
  begin
    case (cache_rsFromMQ_deqP)
      1'd0:
	  CASE_cache_rsFromMQ_deqP_0_cache_rsFromMQ_data_ETC__q73 =
	      cache_rsFromMQ_data_0[260:197];
      1'd1:
	  CASE_cache_rsFromMQ_deqP_0_cache_rsFromMQ_data_ETC__q73 =
	      cache_rsFromMQ_data_1[260:197];
    endcase
  end
  always@(cache_rsFromMQ_deqP or
	  cache_rsFromMQ_data_0 or cache_rsFromMQ_data_1)
  begin
    case (cache_rsFromMQ_deqP)
      1'd0:
	  CASE_cache_rsFromMQ_deqP_0_cache_rsFromMQ_data_ETC__q74 =
	      cache_rsFromMQ_data_0[196:133];
      1'd1:
	  CASE_cache_rsFromMQ_deqP_0_cache_rsFromMQ_data_ETC__q74 =
	      cache_rsFromMQ_data_1[196:133];
    endcase
  end
  always@(cache_rsFromCQ_deqP or
	  cache_rsFromCQ_data_0 or cache_rsFromCQ_data_1)
  begin
    case (cache_rsFromCQ_deqP)
      1'd0:
	  CASE_cache_rsFromCQ_deqP_0_cache_rsFromCQ_data_ETC__q75 =
	      cache_rsFromCQ_data_0[257:194];
      1'd1:
	  CASE_cache_rsFromCQ_deqP_0_cache_rsFromCQ_data_ETC__q75 =
	      cache_rsFromCQ_data_1[257:194];
    endcase
  end
  always@(cache_rsFromCQ_deqP or
	  cache_rsFromCQ_data_0 or cache_rsFromCQ_data_1)
  begin
    case (cache_rsFromCQ_deqP)
      1'd0:
	  CASE_cache_rsFromCQ_deqP_0_cache_rsFromCQ_data_ETC__q76 =
	      cache_rsFromCQ_data_0[193:130];
      1'd1:
	  CASE_cache_rsFromCQ_deqP_0_cache_rsFromCQ_data_ETC__q76 =
	      cache_rsFromCQ_data_1[193:130];
    endcase
  end
  always@(cache_pipeline$unguard_first or
	  cache_cRqMshr$sendRqToC_searchNeedRqChild)
  begin
    case (cache_pipeline$unguard_first[584:583])
      2'd0:
	  CASE_cache_pipelineunguard_first_BITS_584_TO__ETC__q77 =
	      cache_pipeline$unguard_first[582:579] !=
	      cache_cRqMshr$sendRqToC_searchNeedRqChild[3:0];
      2'd2:
	  CASE_cache_pipelineunguard_first_BITS_584_TO__ETC__q77 =
	      !cache_pipeline$unguard_first[517] ||
	      cache_pipeline$unguard_first[516:513] !=
	      cache_cRqMshr$sendRqToC_searchNeedRqChild[3:0];
      default: CASE_cache_pipelineunguard_first_BITS_584_TO__ETC__q77 =
		   cache_pipeline$unguard_first[584:583] != 2'd1 ||
		   !cache_pipeline$unguard_first[517] ||
		   cache_pipeline$unguard_first[516:513] !=
		   cache_cRqMshr$sendRqToC_searchNeedRqChild[3:0];
    endcase
  end
  always@(cache_cRqMshr$pipelineResp_getRq or cache_pipeline$first)
  begin
    case (cache_cRqMshr$pipelineResp_getRq[82:81])
      2'd0:
	  CASE_cache_cRqMshrpipelineResp_getRq_BITS_82__ETC__q79 =
	      cache_pipeline$first[519:518];
      2'd1:
	  CASE_cache_cRqMshrpipelineResp_getRq_BITS_82__ETC__q79 =
	      cache_pipeline$first[521:520];
      2'd2:
	  CASE_cache_cRqMshrpipelineResp_getRq_BITS_82__ETC__q79 =
	      cache_pipeline$first[523:522];
      2'd3:
	  CASE_cache_cRqMshrpipelineResp_getRq_BITS_82__ETC__q79 =
	      2'b10 /* unspecified value */ ;
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q80 =
	      cache_rqFromDmaQ_data_0[591];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q80 =
	      cache_rqFromDmaQ_data_1[591];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q81 =
	      cache_rqFromDmaQ_data_0[590];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q81 =
	      cache_rqFromDmaQ_data_1[590];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q82 =
	      cache_rqFromDmaQ_data_0[589];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q82 =
	      cache_rqFromDmaQ_data_1[589];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q83 =
	      cache_rqFromDmaQ_data_0[588];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q83 =
	      cache_rqFromDmaQ_data_1[588];
    endcase
  end
  always@(cache_pipeline$first)
  begin
    case (cache_pipeline$first[580:579])
      2'd0:
	  SEL_ARR_cache_pipeline_first__581_BITS_519_TO__ETC___d3403 =
	      cache_pipeline$first[519:518];
      2'd1:
	  SEL_ARR_cache_pipeline_first__581_BITS_519_TO__ETC___d3403 =
	      cache_pipeline$first[521:520];
      2'd2:
	  SEL_ARR_cache_pipeline_first__581_BITS_519_TO__ETC___d3403 =
	      cache_pipeline$first[523:522];
      2'd3:
	  SEL_ARR_cache_pipeline_first__581_BITS_519_TO__ETC___d3403 =
	      2'b10 /* unspecified value */ ;
    endcase
  end
  always@(cache_pipeline$first or cache_cRqMshr$pipelineResp_getSlot)
  begin
    case (cache_pipeline$first[580:579])
      2'd0:
	  CASE_cache_pipelinefirst_BITS_580_TO_579_0_ca_ETC__q84 =
	      cache_cRqMshr$pipelineResp_getSlot[1:0];
      2'd1:
	  CASE_cache_pipelinefirst_BITS_580_TO_579_0_ca_ETC__q84 =
	      cache_cRqMshr$pipelineResp_getSlot[5:4];
      2'd2:
	  CASE_cache_pipelinefirst_BITS_580_TO_579_0_ca_ETC__q84 =
	      cache_cRqMshr$pipelineResp_getSlot[9:8];
      2'd3:
	  CASE_cache_pipelinefirst_BITS_580_TO_579_0_ca_ETC__q84 =
	      2'b10 /* unspecified value */ ;
    endcase
  end
  always@(cache_pipeline$first or cache_cRqMshr$pipelineResp_getSlot)
  begin
    case (cache_pipeline$first[580:579])
      2'd0:
	  SEL_ARR_cache_cRqMshr_pipelineResp_getSlot_IF__ETC___d3446 =
	      cache_cRqMshr$pipelineResp_getSlot[3:2] == 2'd2;
      2'd1:
	  SEL_ARR_cache_cRqMshr_pipelineResp_getSlot_IF__ETC___d3446 =
	      cache_cRqMshr$pipelineResp_getSlot[7:6] == 2'd2;
      2'd2:
	  SEL_ARR_cache_cRqMshr_pipelineResp_getSlot_IF__ETC___d3446 =
	      cache_cRqMshr$pipelineResp_getSlot[11:10] == 2'd2;
      2'd3:
	  SEL_ARR_cache_cRqMshr_pipelineResp_getSlot_IF__ETC___d3446 =
	      1'b0 /* unspecified value */ ;
    endcase
  end
  always@(cache_pipeline$first or cache_cRqMshr$pipelineResp_getSlot)
  begin
    case (cache_pipeline$first[580:579])
      2'd0:
	  SEL_ARR_cache_cRqMshr_pipelineResp_getSlot_IF__ETC___d3431 =
	      cache_cRqMshr$pipelineResp_getSlot[3:2] == 2'd1;
      2'd1:
	  SEL_ARR_cache_cRqMshr_pipelineResp_getSlot_IF__ETC___d3431 =
	      cache_cRqMshr$pipelineResp_getSlot[7:6] == 2'd1;
      2'd2:
	  SEL_ARR_cache_cRqMshr_pipelineResp_getSlot_IF__ETC___d3431 =
	      cache_cRqMshr$pipelineResp_getSlot[11:10] == 2'd1;
      2'd3:
	  SEL_ARR_cache_cRqMshr_pipelineResp_getSlot_IF__ETC___d3431 =
	      1'b0 /* unspecified value */ ;
    endcase
  end
  always@(cache_rsLdToDmaQ_deqP or
	  cache_rsLdToDmaQ_data_0 or cache_rsLdToDmaQ_data_1)
  begin
    case (cache_rsLdToDmaQ_deqP)
      1'd0:
	  CASE_cache_rsLdToDmaQ_deqP_0_cache_rsLdToDmaQ__ETC__q85 =
	      cache_rsLdToDmaQ_data_0[527:464];
      1'd1:
	  CASE_cache_rsLdToDmaQ_deqP_0_cache_rsLdToDmaQ__ETC__q85 =
	      cache_rsLdToDmaQ_data_1[527:464];
    endcase
  end
  always@(cache_rsLdToDmaQ_deqP or
	  cache_rsLdToDmaQ_data_0 or cache_rsLdToDmaQ_data_1)
  begin
    case (cache_rsLdToDmaQ_deqP)
      1'd0:
	  CASE_cache_rsLdToDmaQ_deqP_0_cache_rsLdToDmaQ__ETC__q86 =
	      cache_rsLdToDmaQ_data_0[463:400];
      1'd1:
	  CASE_cache_rsLdToDmaQ_deqP_0_cache_rsLdToDmaQ__ETC__q86 =
	      cache_rsLdToDmaQ_data_1[463:400];
    endcase
  end
  always@(cache_rsLdToDmaQ_deqP or
	  cache_rsLdToDmaQ_data_0 or cache_rsLdToDmaQ_data_1)
  begin
    case (cache_rsLdToDmaQ_deqP)
      1'd0:
	  CASE_cache_rsLdToDmaQ_deqP_0_cache_rsLdToDmaQ__ETC__q87 =
	      cache_rsLdToDmaQ_data_0[399:336];
      1'd1:
	  CASE_cache_rsLdToDmaQ_deqP_0_cache_rsLdToDmaQ__ETC__q87 =
	      cache_rsLdToDmaQ_data_1[399:336];
    endcase
  end
  always@(cache_toCQ_deqP or cache_toCQ_data_0 or cache_toCQ_data_1)
  begin
    case (cache_toCQ_deqP)
      1'd0:
	  CASE_cache_toCQ_deqP_0_cache_toCQ_data_0_BITS__ETC__q88 =
	      cache_toCQ_data_0[514:451];
      1'd1:
	  CASE_cache_toCQ_deqP_0_cache_toCQ_data_0_BITS__ETC__q88 =
	      cache_toCQ_data_1[514:451];
    endcase
  end
  always@(cache_toCQ_deqP or cache_toCQ_data_0 or cache_toCQ_data_1)
  begin
    case (cache_toCQ_deqP)
      1'd0:
	  CASE_cache_toCQ_deqP_0_cache_toCQ_data_0_BITS__ETC__q89 =
	      cache_toCQ_data_0[450:387];
      1'd1:
	  CASE_cache_toCQ_deqP_0_cache_toCQ_data_0_BITS__ETC__q89 =
	      cache_toCQ_data_1[450:387];
    endcase
  end
  always@(cache_toCQ_deqP or cache_toCQ_data_0 or cache_toCQ_data_1)
  begin
    case (cache_toCQ_deqP)
      1'd0:
	  CASE_cache_toCQ_deqP_0_cache_toCQ_data_0_BITS__ETC__q90 =
	      cache_toCQ_data_0[386:323];
      1'd1:
	  CASE_cache_toCQ_deqP_0_cache_toCQ_data_0_BITS__ETC__q90 =
	      cache_toCQ_data_1[386:323];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q91 =
	      cache_rqFromDmaQ_data_0[527:464];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q91 =
	      cache_rqFromDmaQ_data_1[527:464];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q92 =
	      cache_rqFromDmaQ_data_0[463:400];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q92 =
	      cache_rqFromDmaQ_data_1[463:400];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q93 =
	      cache_rqFromDmaQ_data_0[399:336];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q93 =
	      cache_rqFromDmaQ_data_1[399:336];
    endcase
  end
  always@(cache_toCQ_deqP or cache_toCQ_data_0 or cache_toCQ_data_1)
  begin
    case (cache_toCQ_deqP)
      1'd0:
	  CASE_cache_toCQ_deqP_0_cache_toCQ_data_0_BITS__ETC__q94 =
	      cache_toCQ_data_0[322:259];
      1'd1:
	  CASE_cache_toCQ_deqP_0_cache_toCQ_data_0_BITS__ETC__q94 =
	      cache_toCQ_data_1[322:259];
    endcase
  end
  always@(cache_toCQ_deqP or cache_toCQ_data_0 or cache_toCQ_data_1)
  begin
    case (cache_toCQ_deqP)
      1'd0:
	  CASE_cache_toCQ_deqP_0_cache_toCQ_data_0_BITS__ETC__q95 =
	      cache_toCQ_data_0[258:195];
      1'd1:
	  CASE_cache_toCQ_deqP_0_cache_toCQ_data_0_BITS__ETC__q95 =
	      cache_toCQ_data_1[258:195];
    endcase
  end
  always@(cache_rsLdToDmaQ_deqP or
	  cache_rsLdToDmaQ_data_0 or cache_rsLdToDmaQ_data_1)
  begin
    case (cache_rsLdToDmaQ_deqP)
      1'd0:
	  CASE_cache_rsLdToDmaQ_deqP_0_cache_rsLdToDmaQ__ETC__q96 =
	      cache_rsLdToDmaQ_data_0[335:272];
      1'd1:
	  CASE_cache_rsLdToDmaQ_deqP_0_cache_rsLdToDmaQ__ETC__q96 =
	      cache_rsLdToDmaQ_data_1[335:272];
    endcase
  end
  always@(cache_rsLdToDmaQ_deqP or
	  cache_rsLdToDmaQ_data_0 or cache_rsLdToDmaQ_data_1)
  begin
    case (cache_rsLdToDmaQ_deqP)
      1'd0:
	  CASE_cache_rsLdToDmaQ_deqP_0_cache_rsLdToDmaQ__ETC__q97 =
	      cache_rsLdToDmaQ_data_0[271:208];
      1'd1:
	  CASE_cache_rsLdToDmaQ_deqP_0_cache_rsLdToDmaQ__ETC__q97 =
	      cache_rsLdToDmaQ_data_1[271:208];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q98 =
	      cache_rqFromDmaQ_data_0[335:272];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q98 =
	      cache_rqFromDmaQ_data_1[335:272];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q99 =
	      cache_rqFromDmaQ_data_0[271:208];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q99 =
	      cache_rqFromDmaQ_data_1[271:208];
    endcase
  end
  always@(cache_toMQ_deqP or cache_toMQ_data_0 or cache_toMQ_data_1)
  begin
    case (cache_toMQ_deqP)
      1'd0:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q100 =
	      cache_toMQ_data_0[575];
      1'd1:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q100 =
	      cache_toMQ_data_1[575];
    endcase
  end
  always@(cache_toMQ_deqP or cache_toMQ_data_0 or cache_toMQ_data_1)
  begin
    case (cache_toMQ_deqP)
      1'd0:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q101 =
	      cache_toMQ_data_0[574];
      1'd1:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q101 =
	      cache_toMQ_data_1[574];
    endcase
  end
  always@(cache_toMQ_deqP or cache_toMQ_data_0 or cache_toMQ_data_1)
  begin
    case (cache_toMQ_deqP)
      1'd0:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q102 =
	      cache_toMQ_data_0[573];
      1'd1:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q102 =
	      cache_toMQ_data_1[573];
    endcase
  end
  always@(cache_toMQ_deqP or cache_toMQ_data_0 or cache_toMQ_data_1)
  begin
    case (cache_toMQ_deqP)
      1'd0:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q103 =
	      cache_toMQ_data_0[572];
      1'd1:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q103 =
	      cache_toMQ_data_1[572];
    endcase
  end
  always@(cache_toMQ_deqP or cache_toMQ_data_0 or cache_toMQ_data_1)
  begin
    case (cache_toMQ_deqP)
      1'd0:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q104 =
	      cache_toMQ_data_0[571];
      1'd1:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q104 =
	      cache_toMQ_data_1[571];
    endcase
  end
  always@(cache_toMQ_deqP or cache_toMQ_data_0 or cache_toMQ_data_1)
  begin
    case (cache_toMQ_deqP)
      1'd0:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q105 =
	      cache_toMQ_data_0[570];
      1'd1:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q105 =
	      cache_toMQ_data_1[570];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q106 =
	      cache_rqFromDmaQ_data_0[587];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q106 =
	      cache_rqFromDmaQ_data_1[587];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q107 =
	      cache_rqFromDmaQ_data_0[586];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q107 =
	      cache_rqFromDmaQ_data_1[586];
    endcase
  end
  always@(cache_toMQ_deqP or cache_toMQ_data_0 or cache_toMQ_data_1)
  begin
    case (cache_toMQ_deqP)
      1'd0:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q108 =
	      cache_toMQ_data_0[569];
      1'd1:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q108 =
	      cache_toMQ_data_1[569];
    endcase
  end
  always@(cache_toMQ_deqP or cache_toMQ_data_0 or cache_toMQ_data_1)
  begin
    case (cache_toMQ_deqP)
      1'd0:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q109 =
	      cache_toMQ_data_0[568];
      1'd1:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q109 =
	      cache_toMQ_data_1[568];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q110 =
	      cache_rqFromDmaQ_data_0[585];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q110 =
	      cache_rqFromDmaQ_data_1[585];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q111 =
	      cache_rqFromDmaQ_data_0[584];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q111 =
	      cache_rqFromDmaQ_data_1[584];
    endcase
  end
  always@(cache_toMQ_deqP or cache_toMQ_data_0 or cache_toMQ_data_1)
  begin
    case (cache_toMQ_deqP)
      1'd0:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q112 =
	      cache_toMQ_data_0[567];
      1'd1:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q112 =
	      cache_toMQ_data_1[567];
    endcase
  end
  always@(cache_toMQ_deqP or cache_toMQ_data_0 or cache_toMQ_data_1)
  begin
    case (cache_toMQ_deqP)
      1'd0:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q113 =
	      cache_toMQ_data_0[566];
      1'd1:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q113 =
	      cache_toMQ_data_1[566];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q114 =
	      cache_rqFromDmaQ_data_0[583];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q114 =
	      cache_rqFromDmaQ_data_1[583];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q115 =
	      cache_rqFromDmaQ_data_0[582];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q115 =
	      cache_rqFromDmaQ_data_1[582];
    endcase
  end
  always@(cache_toMQ_deqP or cache_toMQ_data_0 or cache_toMQ_data_1)
  begin
    case (cache_toMQ_deqP)
      1'd0:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q116 =
	      cache_toMQ_data_0[565];
      1'd1:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q116 =
	      cache_toMQ_data_1[565];
    endcase
  end
  always@(cache_toMQ_deqP or cache_toMQ_data_0 or cache_toMQ_data_1)
  begin
    case (cache_toMQ_deqP)
      1'd0:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q117 =
	      cache_toMQ_data_0[564];
      1'd1:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q117 =
	      cache_toMQ_data_1[564];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q118 =
	      cache_rqFromDmaQ_data_0[581];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q118 =
	      cache_rqFromDmaQ_data_1[581];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q119 =
	      cache_rqFromDmaQ_data_0[580];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q119 =
	      cache_rqFromDmaQ_data_1[580];
    endcase
  end
  always@(cache_toMQ_deqP or cache_toMQ_data_0 or cache_toMQ_data_1)
  begin
    case (cache_toMQ_deqP)
      1'd0:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q120 =
	      cache_toMQ_data_0[563];
      1'd1:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q120 =
	      cache_toMQ_data_1[563];
    endcase
  end
  always@(cache_toMQ_deqP or cache_toMQ_data_0 or cache_toMQ_data_1)
  begin
    case (cache_toMQ_deqP)
      1'd0:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q121 =
	      cache_toMQ_data_0[562];
      1'd1:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q121 =
	      cache_toMQ_data_1[562];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q122 =
	      cache_rqFromDmaQ_data_0[579];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q122 =
	      cache_rqFromDmaQ_data_1[579];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q123 =
	      cache_rqFromDmaQ_data_0[578];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q123 =
	      cache_rqFromDmaQ_data_1[578];
    endcase
  end
  always@(cache_toMQ_deqP or cache_toMQ_data_0 or cache_toMQ_data_1)
  begin
    case (cache_toMQ_deqP)
      1'd0:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q124 =
	      cache_toMQ_data_0[561];
      1'd1:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q124 =
	      cache_toMQ_data_1[561];
    endcase
  end
  always@(cache_toMQ_deqP or cache_toMQ_data_0 or cache_toMQ_data_1)
  begin
    case (cache_toMQ_deqP)
      1'd0:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q125 =
	      cache_toMQ_data_0[560];
      1'd1:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q125 =
	      cache_toMQ_data_1[560];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q126 =
	      cache_rqFromDmaQ_data_0[577];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q126 =
	      cache_rqFromDmaQ_data_1[577];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q127 =
	      cache_rqFromDmaQ_data_0[576];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q127 =
	      cache_rqFromDmaQ_data_1[576];
    endcase
  end
  always@(cache_toMQ_deqP or cache_toMQ_data_0 or cache_toMQ_data_1)
  begin
    case (cache_toMQ_deqP)
      1'd0:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q128 =
	      cache_toMQ_data_0[559];
      1'd1:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q128 =
	      cache_toMQ_data_1[559];
    endcase
  end
  always@(cache_toMQ_deqP or cache_toMQ_data_0 or cache_toMQ_data_1)
  begin
    case (cache_toMQ_deqP)
      1'd0:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q129 =
	      cache_toMQ_data_0[558];
      1'd1:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q129 =
	      cache_toMQ_data_1[558];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q130 =
	      cache_rqFromDmaQ_data_0[575];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q130 =
	      cache_rqFromDmaQ_data_1[575];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q131 =
	      cache_rqFromDmaQ_data_0[574];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q131 =
	      cache_rqFromDmaQ_data_1[574];
    endcase
  end
  always@(cache_toMQ_deqP or cache_toMQ_data_0 or cache_toMQ_data_1)
  begin
    case (cache_toMQ_deqP)
      1'd0:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q132 =
	      cache_toMQ_data_0[557];
      1'd1:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q132 =
	      cache_toMQ_data_1[557];
    endcase
  end
  always@(cache_toMQ_deqP or cache_toMQ_data_0 or cache_toMQ_data_1)
  begin
    case (cache_toMQ_deqP)
      1'd0:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q133 =
	      cache_toMQ_data_0[556];
      1'd1:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q133 =
	      cache_toMQ_data_1[556];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q134 =
	      cache_rqFromDmaQ_data_0[573];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q134 =
	      cache_rqFromDmaQ_data_1[573];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q135 =
	      cache_rqFromDmaQ_data_0[572];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q135 =
	      cache_rqFromDmaQ_data_1[572];
    endcase
  end
  always@(cache_toMQ_deqP or cache_toMQ_data_0 or cache_toMQ_data_1)
  begin
    case (cache_toMQ_deqP)
      1'd0:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q136 =
	      cache_toMQ_data_0[555];
      1'd1:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q136 =
	      cache_toMQ_data_1[555];
    endcase
  end
  always@(cache_toMQ_deqP or cache_toMQ_data_0 or cache_toMQ_data_1)
  begin
    case (cache_toMQ_deqP)
      1'd0:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q137 =
	      cache_toMQ_data_0[554];
      1'd1:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q137 =
	      cache_toMQ_data_1[554];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q138 =
	      cache_rqFromDmaQ_data_0[571];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q138 =
	      cache_rqFromDmaQ_data_1[571];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q139 =
	      cache_rqFromDmaQ_data_0[570];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q139 =
	      cache_rqFromDmaQ_data_1[570];
    endcase
  end
  always@(cache_toMQ_deqP or cache_toMQ_data_0 or cache_toMQ_data_1)
  begin
    case (cache_toMQ_deqP)
      1'd0:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q140 =
	      cache_toMQ_data_0[553];
      1'd1:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q140 =
	      cache_toMQ_data_1[553];
    endcase
  end
  always@(cache_toMQ_deqP or cache_toMQ_data_0 or cache_toMQ_data_1)
  begin
    case (cache_toMQ_deqP)
      1'd0:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q141 =
	      cache_toMQ_data_0[552];
      1'd1:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q141 =
	      cache_toMQ_data_1[552];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q142 =
	      cache_rqFromDmaQ_data_0[569];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q142 =
	      cache_rqFromDmaQ_data_1[569];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q143 =
	      cache_rqFromDmaQ_data_0[568];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q143 =
	      cache_rqFromDmaQ_data_1[568];
    endcase
  end
  always@(cache_toMQ_deqP or cache_toMQ_data_0 or cache_toMQ_data_1)
  begin
    case (cache_toMQ_deqP)
      1'd0:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q144 =
	      cache_toMQ_data_0[551];
      1'd1:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q144 =
	      cache_toMQ_data_1[551];
    endcase
  end
  always@(cache_toMQ_deqP or cache_toMQ_data_0 or cache_toMQ_data_1)
  begin
    case (cache_toMQ_deqP)
      1'd0:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q145 =
	      cache_toMQ_data_0[550];
      1'd1:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q145 =
	      cache_toMQ_data_1[550];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q146 =
	      cache_rqFromDmaQ_data_0[567];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q146 =
	      cache_rqFromDmaQ_data_1[567];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q147 =
	      cache_rqFromDmaQ_data_0[566];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q147 =
	      cache_rqFromDmaQ_data_1[566];
    endcase
  end
  always@(cache_toMQ_deqP or cache_toMQ_data_0 or cache_toMQ_data_1)
  begin
    case (cache_toMQ_deqP)
      1'd0:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q148 =
	      cache_toMQ_data_0[549];
      1'd1:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q148 =
	      cache_toMQ_data_1[549];
    endcase
  end
  always@(cache_toMQ_deqP or cache_toMQ_data_0 or cache_toMQ_data_1)
  begin
    case (cache_toMQ_deqP)
      1'd0:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q149 =
	      cache_toMQ_data_0[548];
      1'd1:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q149 =
	      cache_toMQ_data_1[548];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q150 =
	      cache_rqFromDmaQ_data_0[565];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q150 =
	      cache_rqFromDmaQ_data_1[565];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q151 =
	      cache_rqFromDmaQ_data_0[564];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q151 =
	      cache_rqFromDmaQ_data_1[564];
    endcase
  end
  always@(cache_toMQ_deqP or cache_toMQ_data_0 or cache_toMQ_data_1)
  begin
    case (cache_toMQ_deqP)
      1'd0:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q152 =
	      cache_toMQ_data_0[547];
      1'd1:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q152 =
	      cache_toMQ_data_1[547];
    endcase
  end
  always@(cache_toMQ_deqP or cache_toMQ_data_0 or cache_toMQ_data_1)
  begin
    case (cache_toMQ_deqP)
      1'd0:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q153 =
	      cache_toMQ_data_0[546];
      1'd1:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q153 =
	      cache_toMQ_data_1[546];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q154 =
	      cache_rqFromDmaQ_data_0[563];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q154 =
	      cache_rqFromDmaQ_data_1[563];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q155 =
	      cache_rqFromDmaQ_data_0[562];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q155 =
	      cache_rqFromDmaQ_data_1[562];
    endcase
  end
  always@(cache_toMQ_deqP or cache_toMQ_data_0 or cache_toMQ_data_1)
  begin
    case (cache_toMQ_deqP)
      1'd0:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q156 =
	      cache_toMQ_data_0[545];
      1'd1:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q156 =
	      cache_toMQ_data_1[545];
    endcase
  end
  always@(cache_toMQ_deqP or cache_toMQ_data_0 or cache_toMQ_data_1)
  begin
    case (cache_toMQ_deqP)
      1'd0:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q157 =
	      cache_toMQ_data_0[544];
      1'd1:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q157 =
	      cache_toMQ_data_1[544];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q158 =
	      cache_rqFromDmaQ_data_0[561];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q158 =
	      cache_rqFromDmaQ_data_1[561];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q159 =
	      cache_rqFromDmaQ_data_0[560];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q159 =
	      cache_rqFromDmaQ_data_1[560];
    endcase
  end
  always@(cache_toMQ_deqP or cache_toMQ_data_0 or cache_toMQ_data_1)
  begin
    case (cache_toMQ_deqP)
      1'd0:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q160 =
	      cache_toMQ_data_0[543];
      1'd1:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q160 =
	      cache_toMQ_data_1[543];
    endcase
  end
  always@(cache_toMQ_deqP or cache_toMQ_data_0 or cache_toMQ_data_1)
  begin
    case (cache_toMQ_deqP)
      1'd0:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q161 =
	      cache_toMQ_data_0[542];
      1'd1:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q161 =
	      cache_toMQ_data_1[542];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q162 =
	      cache_rqFromDmaQ_data_0[559];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q162 =
	      cache_rqFromDmaQ_data_1[559];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q163 =
	      cache_rqFromDmaQ_data_0[558];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q163 =
	      cache_rqFromDmaQ_data_1[558];
    endcase
  end
  always@(cache_toMQ_deqP or cache_toMQ_data_0 or cache_toMQ_data_1)
  begin
    case (cache_toMQ_deqP)
      1'd0:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q164 =
	      cache_toMQ_data_0[541];
      1'd1:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q164 =
	      cache_toMQ_data_1[541];
    endcase
  end
  always@(cache_toMQ_deqP or cache_toMQ_data_0 or cache_toMQ_data_1)
  begin
    case (cache_toMQ_deqP)
      1'd0:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q165 =
	      cache_toMQ_data_0[540];
      1'd1:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q165 =
	      cache_toMQ_data_1[540];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q166 =
	      cache_rqFromDmaQ_data_0[557];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q166 =
	      cache_rqFromDmaQ_data_1[557];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q167 =
	      cache_rqFromDmaQ_data_0[556];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q167 =
	      cache_rqFromDmaQ_data_1[556];
    endcase
  end
  always@(cache_toMQ_deqP or cache_toMQ_data_0 or cache_toMQ_data_1)
  begin
    case (cache_toMQ_deqP)
      1'd0:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q168 =
	      cache_toMQ_data_0[539];
      1'd1:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q168 =
	      cache_toMQ_data_1[539];
    endcase
  end
  always@(cache_toMQ_deqP or cache_toMQ_data_0 or cache_toMQ_data_1)
  begin
    case (cache_toMQ_deqP)
      1'd0:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q169 =
	      cache_toMQ_data_0[538];
      1'd1:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q169 =
	      cache_toMQ_data_1[538];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q170 =
	      cache_rqFromDmaQ_data_0[555];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q170 =
	      cache_rqFromDmaQ_data_1[555];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q171 =
	      cache_rqFromDmaQ_data_0[554];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q171 =
	      cache_rqFromDmaQ_data_1[554];
    endcase
  end
  always@(cache_toMQ_deqP or cache_toMQ_data_0 or cache_toMQ_data_1)
  begin
    case (cache_toMQ_deqP)
      1'd0:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q172 =
	      cache_toMQ_data_0[537];
      1'd1:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q172 =
	      cache_toMQ_data_1[537];
    endcase
  end
  always@(cache_toMQ_deqP or cache_toMQ_data_0 or cache_toMQ_data_1)
  begin
    case (cache_toMQ_deqP)
      1'd0:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q173 =
	      cache_toMQ_data_0[536];
      1'd1:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q173 =
	      cache_toMQ_data_1[536];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q174 =
	      cache_rqFromDmaQ_data_0[553];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q174 =
	      cache_rqFromDmaQ_data_1[553];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q175 =
	      cache_rqFromDmaQ_data_0[552];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q175 =
	      cache_rqFromDmaQ_data_1[552];
    endcase
  end
  always@(cache_toMQ_deqP or cache_toMQ_data_0 or cache_toMQ_data_1)
  begin
    case (cache_toMQ_deqP)
      1'd0:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q176 =
	      cache_toMQ_data_0[535];
      1'd1:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q176 =
	      cache_toMQ_data_1[535];
    endcase
  end
  always@(cache_toMQ_deqP or cache_toMQ_data_0 or cache_toMQ_data_1)
  begin
    case (cache_toMQ_deqP)
      1'd0:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q177 =
	      cache_toMQ_data_0[534];
      1'd1:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q177 =
	      cache_toMQ_data_1[534];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q178 =
	      cache_rqFromDmaQ_data_0[551];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q178 =
	      cache_rqFromDmaQ_data_1[551];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q179 =
	      cache_rqFromDmaQ_data_0[550];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q179 =
	      cache_rqFromDmaQ_data_1[550];
    endcase
  end
  always@(cache_toMQ_deqP or cache_toMQ_data_0 or cache_toMQ_data_1)
  begin
    case (cache_toMQ_deqP)
      1'd0:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q180 =
	      cache_toMQ_data_0[533];
      1'd1:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q180 =
	      cache_toMQ_data_1[533];
    endcase
  end
  always@(cache_toMQ_deqP or cache_toMQ_data_0 or cache_toMQ_data_1)
  begin
    case (cache_toMQ_deqP)
      1'd0:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q181 =
	      cache_toMQ_data_0[532];
      1'd1:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q181 =
	      cache_toMQ_data_1[532];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q182 =
	      cache_rqFromDmaQ_data_0[549];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q182 =
	      cache_rqFromDmaQ_data_1[549];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q183 =
	      cache_rqFromDmaQ_data_0[548];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q183 =
	      cache_rqFromDmaQ_data_1[548];
    endcase
  end
  always@(cache_toMQ_deqP or cache_toMQ_data_0 or cache_toMQ_data_1)
  begin
    case (cache_toMQ_deqP)
      1'd0:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q184 =
	      cache_toMQ_data_0[531];
      1'd1:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q184 =
	      cache_toMQ_data_1[531];
    endcase
  end
  always@(cache_toMQ_deqP or cache_toMQ_data_0 or cache_toMQ_data_1)
  begin
    case (cache_toMQ_deqP)
      1'd0:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q185 =
	      cache_toMQ_data_0[530];
      1'd1:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q185 =
	      cache_toMQ_data_1[530];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q186 =
	      cache_rqFromDmaQ_data_0[547];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q186 =
	      cache_rqFromDmaQ_data_1[547];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q187 =
	      cache_rqFromDmaQ_data_0[546];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q187 =
	      cache_rqFromDmaQ_data_1[546];
    endcase
  end
  always@(cache_toMQ_deqP or cache_toMQ_data_0 or cache_toMQ_data_1)
  begin
    case (cache_toMQ_deqP)
      1'd0:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q188 =
	      cache_toMQ_data_0[529];
      1'd1:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q188 =
	      cache_toMQ_data_1[529];
    endcase
  end
  always@(cache_toMQ_deqP or cache_toMQ_data_0 or cache_toMQ_data_1)
  begin
    case (cache_toMQ_deqP)
      1'd0:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q189 =
	      cache_toMQ_data_0[528];
      1'd1:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q189 =
	      cache_toMQ_data_1[528];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q190 =
	      cache_rqFromDmaQ_data_0[545];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q190 =
	      cache_rqFromDmaQ_data_1[545];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q191 =
	      cache_rqFromDmaQ_data_0[544];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q191 =
	      cache_rqFromDmaQ_data_1[544];
    endcase
  end
  always@(cache_toMQ_deqP or cache_toMQ_data_0 or cache_toMQ_data_1)
  begin
    case (cache_toMQ_deqP)
      1'd0:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q192 =
	      cache_toMQ_data_0[527];
      1'd1:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q192 =
	      cache_toMQ_data_1[527];
    endcase
  end
  always@(cache_toMQ_deqP or cache_toMQ_data_0 or cache_toMQ_data_1)
  begin
    case (cache_toMQ_deqP)
      1'd0:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q193 =
	      cache_toMQ_data_0[526];
      1'd1:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q193 =
	      cache_toMQ_data_1[526];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q194 =
	      cache_rqFromDmaQ_data_0[543];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q194 =
	      cache_rqFromDmaQ_data_1[543];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q195 =
	      cache_rqFromDmaQ_data_0[542];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q195 =
	      cache_rqFromDmaQ_data_1[542];
    endcase
  end
  always@(cache_toMQ_deqP or cache_toMQ_data_0 or cache_toMQ_data_1)
  begin
    case (cache_toMQ_deqP)
      1'd0:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q196 =
	      cache_toMQ_data_0[525];
      1'd1:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q196 =
	      cache_toMQ_data_1[525];
    endcase
  end
  always@(cache_toMQ_deqP or cache_toMQ_data_0 or cache_toMQ_data_1)
  begin
    case (cache_toMQ_deqP)
      1'd0:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q197 =
	      cache_toMQ_data_0[524];
      1'd1:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q197 =
	      cache_toMQ_data_1[524];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q198 =
	      cache_rqFromDmaQ_data_0[541];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q198 =
	      cache_rqFromDmaQ_data_1[541];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q199 =
	      cache_rqFromDmaQ_data_0[540];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q199 =
	      cache_rqFromDmaQ_data_1[540];
    endcase
  end
  always@(cache_toMQ_deqP or cache_toMQ_data_0 or cache_toMQ_data_1)
  begin
    case (cache_toMQ_deqP)
      1'd0:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q200 =
	      cache_toMQ_data_0[523];
      1'd1:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q200 =
	      cache_toMQ_data_1[523];
    endcase
  end
  always@(cache_toMQ_deqP or cache_toMQ_data_0 or cache_toMQ_data_1)
  begin
    case (cache_toMQ_deqP)
      1'd0:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q201 =
	      cache_toMQ_data_0[522];
      1'd1:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q201 =
	      cache_toMQ_data_1[522];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q202 =
	      cache_rqFromDmaQ_data_0[539];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q202 =
	      cache_rqFromDmaQ_data_1[539];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q203 =
	      cache_rqFromDmaQ_data_0[538];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q203 =
	      cache_rqFromDmaQ_data_1[538];
    endcase
  end
  always@(cache_toMQ_deqP or cache_toMQ_data_0 or cache_toMQ_data_1)
  begin
    case (cache_toMQ_deqP)
      1'd0:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q204 =
	      cache_toMQ_data_0[521];
      1'd1:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q204 =
	      cache_toMQ_data_1[521];
    endcase
  end
  always@(cache_toMQ_deqP or cache_toMQ_data_0 or cache_toMQ_data_1)
  begin
    case (cache_toMQ_deqP)
      1'd0:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q205 =
	      cache_toMQ_data_0[520];
      1'd1:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q205 =
	      cache_toMQ_data_1[520];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q206 =
	      cache_rqFromDmaQ_data_0[537];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q206 =
	      cache_rqFromDmaQ_data_1[537];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q207 =
	      cache_rqFromDmaQ_data_0[536];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q207 =
	      cache_rqFromDmaQ_data_1[536];
    endcase
  end
  always@(cache_toMQ_deqP or cache_toMQ_data_0 or cache_toMQ_data_1)
  begin
    case (cache_toMQ_deqP)
      1'd0:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q208 =
	      cache_toMQ_data_0[519];
      1'd1:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q208 =
	      cache_toMQ_data_1[519];
    endcase
  end
  always@(cache_toMQ_deqP or cache_toMQ_data_0 or cache_toMQ_data_1)
  begin
    case (cache_toMQ_deqP)
      1'd0:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q209 =
	      cache_toMQ_data_0[518];
      1'd1:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q209 =
	      cache_toMQ_data_1[518];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q210 =
	      cache_rqFromDmaQ_data_0[535];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q210 =
	      cache_rqFromDmaQ_data_1[535];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q211 =
	      cache_rqFromDmaQ_data_0[534];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q211 =
	      cache_rqFromDmaQ_data_1[534];
    endcase
  end
  always@(cache_toMQ_deqP or cache_toMQ_data_0 or cache_toMQ_data_1)
  begin
    case (cache_toMQ_deqP)
      1'd0:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q212 =
	      cache_toMQ_data_0[517];
      1'd1:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q212 =
	      cache_toMQ_data_1[517];
    endcase
  end
  always@(cache_toMQ_deqP or cache_toMQ_data_0 or cache_toMQ_data_1)
  begin
    case (cache_toMQ_deqP)
      1'd0:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q213 =
	      cache_toMQ_data_0[516];
      1'd1:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q213 =
	      cache_toMQ_data_1[516];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q214 =
	      cache_rqFromDmaQ_data_0[533];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q214 =
	      cache_rqFromDmaQ_data_1[533];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q215 =
	      cache_rqFromDmaQ_data_0[532];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q215 =
	      cache_rqFromDmaQ_data_1[532];
    endcase
  end
  always@(cache_toMQ_deqP or cache_toMQ_data_0 or cache_toMQ_data_1)
  begin
    case (cache_toMQ_deqP)
      1'd0:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q216 =
	      cache_toMQ_data_0[515];
      1'd1:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q216 =
	      cache_toMQ_data_1[515];
    endcase
  end
  always@(cache_toMQ_deqP or cache_toMQ_data_0 or cache_toMQ_data_1)
  begin
    case (cache_toMQ_deqP)
      1'd0:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q217 =
	      cache_toMQ_data_0[514];
      1'd1:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q217 =
	      cache_toMQ_data_1[514];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q218 =
	      cache_rqFromDmaQ_data_0[531];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q218 =
	      cache_rqFromDmaQ_data_1[531];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q219 =
	      cache_rqFromDmaQ_data_0[530];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q219 =
	      cache_rqFromDmaQ_data_1[530];
    endcase
  end
  always@(cache_toMQ_deqP or cache_toMQ_data_0 or cache_toMQ_data_1)
  begin
    case (cache_toMQ_deqP)
      1'd0:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BITS__ETC__q220 =
	      cache_toMQ_data_0[511:448];
      1'd1:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BITS__ETC__q220 =
	      cache_toMQ_data_1[511:448];
    endcase
  end
  always@(cache_toMQ_deqP or cache_toMQ_data_0 or cache_toMQ_data_1)
  begin
    case (cache_toMQ_deqP)
      1'd0:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BITS__ETC__q221 =
	      cache_toMQ_data_0[447:384];
      1'd1:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BITS__ETC__q221 =
	      cache_toMQ_data_1[447:384];
    endcase
  end
  always@(cache_toMQ_deqP or cache_toMQ_data_0 or cache_toMQ_data_1)
  begin
    case (cache_toMQ_deqP)
      1'd0:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BITS__ETC__q222 =
	      cache_toMQ_data_0[383:320];
      1'd1:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BITS__ETC__q222 =
	      cache_toMQ_data_1[383:320];
    endcase
  end
  always@(cache_toMQ_deqP or cache_toMQ_data_0 or cache_toMQ_data_1)
  begin
    case (cache_toMQ_deqP)
      1'd0:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BITS__ETC__q223 =
	      cache_toMQ_data_0[319:256];
      1'd1:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BITS__ETC__q223 =
	      cache_toMQ_data_1[319:256];
    endcase
  end
  always@(cache_toMQ_deqP or cache_toMQ_data_0 or cache_toMQ_data_1)
  begin
    case (cache_toMQ_deqP)
      1'd0:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BITS__ETC__q224 =
	      cache_toMQ_data_0[255:192];
      1'd1:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BITS__ETC__q224 =
	      cache_toMQ_data_1[255:192];
    endcase
  end
  always@(cache_toMQ_deqP or cache_toMQ_data_0 or cache_toMQ_data_1)
  begin
    case (cache_toMQ_deqP)
      1'd0:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BITS__ETC__q225 =
	      cache_toMQ_data_0[191:128];
      1'd1:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BITS__ETC__q225 =
	      cache_toMQ_data_1[191:128];
    endcase
  end
  always@(child__h313067 or cache_cRqMshr$sendRqToC_getSlot)
  begin
    case (child__h313067)
      2'd0:
	  SEL_ARR_IF_cache_cRqMshr_sendRqToC_getSlot_IF__ETC___d2522 =
	      cache_cRqMshr$sendRqToC_getSlot[1:0];
      2'd1:
	  SEL_ARR_IF_cache_cRqMshr_sendRqToC_getSlot_IF__ETC___d2522 =
	      cache_cRqMshr$sendRqToC_getSlot[5:4];
      2'd2:
	  SEL_ARR_IF_cache_cRqMshr_sendRqToC_getSlot_IF__ETC___d2522 =
	      cache_cRqMshr$sendRqToC_getSlot[9:8];
      2'd3:
	  SEL_ARR_IF_cache_cRqMshr_sendRqToC_getSlot_IF__ETC___d2522 =
	      2'b10 /* unspecified value */ ;
    endcase
  end
  always@(cache_rsFromMQ_deqP or
	  cache_rsFromMQ_data_0 or cache_rsFromMQ_data_1)
  begin
    case (cache_rsFromMQ_deqP)
      1'd0:
	  CASE_cache_rsFromMQ_deqP_0_cache_rsFromMQ_data_ETC__q226 =
	      cache_rsFromMQ_data_0[132:69];
      1'd1:
	  CASE_cache_rsFromMQ_deqP_0_cache_rsFromMQ_data_ETC__q226 =
	      cache_rsFromMQ_data_1[132:69];
    endcase
  end
  always@(cache_rsFromMQ_deqP or
	  cache_rsFromMQ_data_0 or cache_rsFromMQ_data_1)
  begin
    case (cache_rsFromMQ_deqP)
      1'd0:
	  CASE_cache_rsFromMQ_deqP_0_cache_rsFromMQ_data_ETC__q227 =
	      cache_rsFromMQ_data_0[68:5];
      1'd1:
	  CASE_cache_rsFromMQ_deqP_0_cache_rsFromMQ_data_ETC__q227 =
	      cache_rsFromMQ_data_1[68:5];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q228 =
	      cache_rqFromDmaQ_data_0[529];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q228 =
	      cache_rqFromDmaQ_data_1[529];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q229 =
	      cache_rqFromDmaQ_data_0[528];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q229 =
	      cache_rqFromDmaQ_data_1[528];
    endcase
  end
  always@(cache_rqFromCQ_deqP or
	  cache_rqFromCQ_data_0 or cache_rqFromCQ_data_1)
  begin
    case (cache_rqFromCQ_deqP)
      1'd0:
	  CASE_cache_rqFromCQ_deqP_0_cache_rqFromCQ_data_ETC__q230 =
	      cache_rqFromCQ_data_0[7:6];
      1'd1:
	  CASE_cache_rqFromCQ_deqP_0_cache_rqFromCQ_data_ETC__q230 =
	      cache_rqFromCQ_data_1[7:6];
    endcase
  end
  always@(cache_rqFromCQ_deqP or
	  cache_rqFromCQ_data_0 or cache_rqFromCQ_data_1)
  begin
    case (cache_rqFromCQ_deqP)
      1'd0:
	  CASE_cache_rqFromCQ_deqP_0_cache_rqFromCQ_data_ETC__q231 =
	      cache_rqFromCQ_data_0[5];
      1'd1:
	  CASE_cache_rqFromCQ_deqP_0_cache_rqFromCQ_data_ETC__q231 =
	      cache_rqFromCQ_data_1[5];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q232 =
	      cache_rqFromDmaQ_data_0[207:144];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q232 =
	      cache_rqFromDmaQ_data_1[207:144];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q233 =
	      cache_rqFromDmaQ_data_0[143:80];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q233 =
	      cache_rqFromDmaQ_data_1[143:80];
    endcase
  end
  always@(cache_toCQ_deqP or cache_toCQ_data_0 or cache_toCQ_data_1)
  begin
    case (cache_toCQ_deqP)
      1'd0:
	  CASE_cache_toCQ_deqP_0_cache_toCQ_data_0_BITS__ETC__q234 =
	      cache_toCQ_data_0[194:131];
      1'd1:
	  CASE_cache_toCQ_deqP_0_cache_toCQ_data_0_BITS__ETC__q234 =
	      cache_toCQ_data_1[194:131];
    endcase
  end
  always@(cache_toCQ_deqP or cache_toCQ_data_0 or cache_toCQ_data_1)
  begin
    case (cache_toCQ_deqP)
      1'd0:
	  CASE_cache_toCQ_deqP_0_cache_toCQ_data_0_BITS__ETC__q235 =
	      cache_toCQ_data_0[130:67];
      1'd1:
	  CASE_cache_toCQ_deqP_0_cache_toCQ_data_0_BITS__ETC__q235 =
	      cache_toCQ_data_1[130:67];
    endcase
  end
  always@(cache_rsFromCQ_deqP or
	  cache_rsFromCQ_data_0 or cache_rsFromCQ_data_1)
  begin
    case (cache_rsFromCQ_deqP)
      1'd0:
	  CASE_cache_rsFromCQ_deqP_0_cache_rsFromCQ_data_ETC__q236 =
	      cache_rsFromCQ_data_0[129:66];
      1'd1:
	  CASE_cache_rsFromCQ_deqP_0_cache_rsFromCQ_data_ETC__q236 =
	      cache_rsFromCQ_data_1[129:66];
    endcase
  end
  always@(cache_rsFromCQ_deqP or
	  cache_rsFromCQ_data_0 or cache_rsFromCQ_data_1)
  begin
    case (cache_rsFromCQ_deqP)
      1'd0:
	  CASE_cache_rsFromCQ_deqP_0_cache_rsFromCQ_data_ETC__q237 =
	      cache_rsFromCQ_data_0[65:2];
      1'd1:
	  CASE_cache_rsFromCQ_deqP_0_cache_rsFromCQ_data_ETC__q237 =
	      cache_rsFromCQ_data_1[65:2];
    endcase
  end
  always@(cache_toCQ_deqP or cache_toCQ_data_0 or cache_toCQ_data_1)
  begin
    case (cache_toCQ_deqP)
      1'd0:
	  CASE_cache_toCQ_deqP_0_cache_toCQ_data_0_BIT_5_ETC__q238 =
	      cache_toCQ_data_0[515];
      1'd1:
	  CASE_cache_toCQ_deqP_0_cache_toCQ_data_0_BIT_5_ETC__q238 =
	      cache_toCQ_data_1[515];
    endcase
  end
  always@(cache_toCQ_deqP or cache_toCQ_data_0 or cache_toCQ_data_1)
  begin
    case (cache_toCQ_deqP)
      1'd0:
	  CASE_cache_toCQ_deqP_0_cache_toCQ_data_0_BITS__ETC__q239 =
	      cache_toCQ_data_0[66:3];
      1'd1:
	  CASE_cache_toCQ_deqP_0_cache_toCQ_data_0_BITS__ETC__q239 =
	      cache_toCQ_data_1[66:3];
    endcase
  end
  always@(cache_rsToCIndexQ_deqP or
	  cache_rsToCIndexQ_data_0 or
	  cache_rsToCIndexQ_data_1 or
	  cache_rsToCIndexQ_data_2 or
	  cache_rsToCIndexQ_data_3 or
	  cache_rsToCIndexQ_data_4 or
	  cache_rsToCIndexQ_data_5 or
	  cache_rsToCIndexQ_data_6 or
	  cache_rsToCIndexQ_data_7 or
	  cache_rsToCIndexQ_data_8 or
	  cache_rsToCIndexQ_data_9 or
	  cache_rsToCIndexQ_data_10 or
	  cache_rsToCIndexQ_data_11 or
	  cache_rsToCIndexQ_data_12 or
	  cache_rsToCIndexQ_data_13 or
	  cache_rsToCIndexQ_data_14 or cache_rsToCIndexQ_data_15)
  begin
    case (cache_rsToCIndexQ_deqP)
      4'd0:
	  SEL_ARR_cache_rsToCIndexQ_data_0_391_BITS_1_TO_ETC___d2445 =
	      cache_rsToCIndexQ_data_0[1:0];
      4'd1:
	  SEL_ARR_cache_rsToCIndexQ_data_0_391_BITS_1_TO_ETC___d2445 =
	      cache_rsToCIndexQ_data_1[1:0];
      4'd2:
	  SEL_ARR_cache_rsToCIndexQ_data_0_391_BITS_1_TO_ETC___d2445 =
	      cache_rsToCIndexQ_data_2[1:0];
      4'd3:
	  SEL_ARR_cache_rsToCIndexQ_data_0_391_BITS_1_TO_ETC___d2445 =
	      cache_rsToCIndexQ_data_3[1:0];
      4'd4:
	  SEL_ARR_cache_rsToCIndexQ_data_0_391_BITS_1_TO_ETC___d2445 =
	      cache_rsToCIndexQ_data_4[1:0];
      4'd5:
	  SEL_ARR_cache_rsToCIndexQ_data_0_391_BITS_1_TO_ETC___d2445 =
	      cache_rsToCIndexQ_data_5[1:0];
      4'd6:
	  SEL_ARR_cache_rsToCIndexQ_data_0_391_BITS_1_TO_ETC___d2445 =
	      cache_rsToCIndexQ_data_6[1:0];
      4'd7:
	  SEL_ARR_cache_rsToCIndexQ_data_0_391_BITS_1_TO_ETC___d2445 =
	      cache_rsToCIndexQ_data_7[1:0];
      4'd8:
	  SEL_ARR_cache_rsToCIndexQ_data_0_391_BITS_1_TO_ETC___d2445 =
	      cache_rsToCIndexQ_data_8[1:0];
      4'd9:
	  SEL_ARR_cache_rsToCIndexQ_data_0_391_BITS_1_TO_ETC___d2445 =
	      cache_rsToCIndexQ_data_9[1:0];
      4'd10:
	  SEL_ARR_cache_rsToCIndexQ_data_0_391_BITS_1_TO_ETC___d2445 =
	      cache_rsToCIndexQ_data_10[1:0];
      4'd11:
	  SEL_ARR_cache_rsToCIndexQ_data_0_391_BITS_1_TO_ETC___d2445 =
	      cache_rsToCIndexQ_data_11[1:0];
      4'd12:
	  SEL_ARR_cache_rsToCIndexQ_data_0_391_BITS_1_TO_ETC___d2445 =
	      cache_rsToCIndexQ_data_12[1:0];
      4'd13:
	  SEL_ARR_cache_rsToCIndexQ_data_0_391_BITS_1_TO_ETC___d2445 =
	      cache_rsToCIndexQ_data_13[1:0];
      4'd14:
	  SEL_ARR_cache_rsToCIndexQ_data_0_391_BITS_1_TO_ETC___d2445 =
	      cache_rsToCIndexQ_data_14[1:0];
      4'd15:
	  SEL_ARR_cache_rsToCIndexQ_data_0_391_BITS_1_TO_ETC___d2445 =
	      cache_rsToCIndexQ_data_15[1:0];
    endcase
  end
  always@(cache_toMQ_deqP or cache_toMQ_data_0 or cache_toMQ_data_1)
  begin
    case (cache_toMQ_deqP)
      1'd0:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q240 =
	      cache_toMQ_data_0[513];
      1'd1:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q240 =
	      cache_toMQ_data_1[513];
    endcase
  end
  always@(cache_toMQ_deqP or cache_toMQ_data_0 or cache_toMQ_data_1)
  begin
    case (cache_toMQ_deqP)
      1'd0:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q241 =
	      cache_toMQ_data_0[512];
      1'd1:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_5_ETC__q241 =
	      cache_toMQ_data_1[512];
    endcase
  end
  always@(cache_rsFromCQ_deqP or
	  cache_rsFromCQ_data_0 or cache_rsFromCQ_data_1)
  begin
    case (cache_rsFromCQ_deqP)
      1'd0:
	  CASE_cache_rsFromCQ_deqP_0_cache_rsFromCQ_data_ETC__q242 =
	      cache_rsFromCQ_data_0[514];
      1'd1:
	  CASE_cache_rsFromCQ_deqP_0_cache_rsFromCQ_data_ETC__q242 =
	      cache_rsFromCQ_data_1[514];
    endcase
  end
  always@(cache_rsFromCQ_deqP or
	  cache_rsFromCQ_data_0 or cache_rsFromCQ_data_1)
  begin
    case (cache_rsFromCQ_deqP)
      1'd0:
	  CASE_cache_rsFromCQ_deqP_0_cache_rsFromCQ_data_ETC__q243 =
	      cache_rsFromCQ_data_0[580:517];
      1'd1:
	  CASE_cache_rsFromCQ_deqP_0_cache_rsFromCQ_data_ETC__q243 =
	      cache_rsFromCQ_data_1[580:517];
    endcase
  end
  always@(cache_rsFromCQ_deqP or
	  cache_rsFromCQ_data_0 or cache_rsFromCQ_data_1)
  begin
    case (cache_rsFromCQ_deqP)
      1'd0:
	  CASE_cache_rsFromCQ_deqP_0_cache_rsFromCQ_data_ETC__q244 =
	      cache_rsFromCQ_data_0[516:515];
      1'd1:
	  CASE_cache_rsFromCQ_deqP_0_cache_rsFromCQ_data_ETC__q244 =
	      cache_rsFromCQ_data_1[516:515];
    endcase
  end
  always@(cache_toMQ_deqP or cache_toMQ_data_0 or cache_toMQ_data_1)
  begin
    case (cache_toMQ_deqP)
      1'd0:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BITS__ETC__q245 =
	      cache_toMQ_data_0[127:64];
      1'd1:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BITS__ETC__q245 =
	      cache_toMQ_data_1[127:64];
    endcase
  end
  always@(cache_toMQ_deqP or cache_toMQ_data_0 or cache_toMQ_data_1)
  begin
    case (cache_toMQ_deqP)
      1'd0:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BITS__ETC__q246 =
	      cache_toMQ_data_0[63:0];
      1'd1:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BITS__ETC__q246 =
	      cache_toMQ_data_1[63:0];
    endcase
  end
  always@(cache_toCQ_deqP or cache_toCQ_data_0 or cache_toCQ_data_1)
  begin
    case (cache_toCQ_deqP)
      1'd0:
	  CASE_cache_toCQ_deqP_0_cache_toCQ_data_0_BITS__ETC__q247 =
	      cache_toCQ_data_0[583:520];
      1'd1:
	  CASE_cache_toCQ_deqP_0_cache_toCQ_data_0_BITS__ETC__q247 =
	      cache_toCQ_data_1[583:520];
    endcase
  end
  always@(cache_toCQ_deqP or cache_toCQ_data_0 or cache_toCQ_data_1)
  begin
    case (cache_toCQ_deqP)
      1'd0:
	  CASE_cache_toCQ_deqP_0_cache_toCQ_data_0_BITS__ETC__q248 =
	      cache_toCQ_data_0[519:518];
      1'd1:
	  CASE_cache_toCQ_deqP_0_cache_toCQ_data_0_BITS__ETC__q248 =
	      cache_toCQ_data_1[519:518];
    endcase
  end
  always@(cache_toCQ_deqP or cache_toCQ_data_0 or cache_toCQ_data_1)
  begin
    case (cache_toCQ_deqP)
      1'd0:
	  CASE_cache_toCQ_deqP_0_cache_toCQ_data_0_BITS__ETC__q249 =
	      cache_toCQ_data_0[67:4];
      1'd1:
	  CASE_cache_toCQ_deqP_0_cache_toCQ_data_0_BITS__ETC__q249 =
	      cache_toCQ_data_1[67:4];
    endcase
  end
  always@(cache_toCQ_deqP or cache_toCQ_data_0 or cache_toCQ_data_1)
  begin
    case (cache_toCQ_deqP)
      1'd0:
	  CASE_cache_toCQ_deqP_0_cache_toCQ_data_0_BITS__ETC__q250 =
	      cache_toCQ_data_0[3:2];
      1'd1:
	  CASE_cache_toCQ_deqP_0_cache_toCQ_data_0_BITS__ETC__q250 =
	      cache_toCQ_data_1[3:2];
    endcase
  end
  always@(cache_toMQ_deqP or cache_toMQ_data_0 or cache_toMQ_data_1)
  begin
    case (cache_toMQ_deqP)
      1'd0:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BITS__ETC__q251 =
	      cache_toMQ_data_0[639:576];
      1'd1:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BITS__ETC__q251 =
	      cache_toMQ_data_1[639:576];
    endcase
  end
  always@(cache_toMQ_deqP or cache_toMQ_data_0 or cache_toMQ_data_1)
  begin
    case (cache_toMQ_deqP)
      1'd0:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BITS__ETC__q252 =
	      cache_toMQ_data_0[68:5];
      1'd1:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BITS__ETC__q252 =
	      cache_toMQ_data_1[68:5];
    endcase
  end
  always@(cache_toMQ_deqP or cache_toMQ_data_0 or cache_toMQ_data_1)
  begin
    case (cache_toMQ_deqP)
      1'd0:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_4_ETC__q253 =
	      cache_toMQ_data_0[4];
      1'd1:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_4_ETC__q253 =
	      cache_toMQ_data_1[4];
    endcase
  end
  always@(child__h313067 or cache_cRqMshr$sendRqToC_getSlot)
  begin
    case (child__h313067)
      2'd0:
	  CASE_child13067_0_cache_cRqMshrsendRqToC_getS_ETC__q254 =
	      cache_cRqMshr$sendRqToC_getSlot[3:2] == 2'd1;
      2'd1:
	  CASE_child13067_0_cache_cRqMshrsendRqToC_getS_ETC__q254 =
	      cache_cRqMshr$sendRqToC_getSlot[7:6] == 2'd1;
      2'd2:
	  CASE_child13067_0_cache_cRqMshrsendRqToC_getS_ETC__q254 =
	      cache_cRqMshr$sendRqToC_getSlot[11:10] == 2'd1;
      2'd3:
	  CASE_child13067_0_cache_cRqMshrsendRqToC_getS_ETC__q254 =
	      1'b0 /* unspecified value */ ;
    endcase
  end
  always@(cache_toCQ_deqP or cache_toCQ_data_0 or cache_toCQ_data_1)
  begin
    case (cache_toCQ_deqP)
      1'd0:
	  CASE_cache_toCQ_deqP_0_NOT_cache_toCQ_data_0_B_ETC__q255 =
	      !cache_toCQ_data_0[584];
      1'd1:
	  CASE_cache_toCQ_deqP_0_NOT_cache_toCQ_data_0_B_ETC__q255 =
	      !cache_toCQ_data_1[584];
    endcase
  end
  always@(cache_toCQ_deqP or cache_toCQ_data_0 or cache_toCQ_data_1)
  begin
    case (cache_toCQ_deqP)
      1'd0:
	  CASE_cache_toCQ_deqP_0_cache_toCQ_data_0_BIT_5_ETC__q256 =
	      cache_toCQ_data_0[584];
      1'd1:
	  CASE_cache_toCQ_deqP_0_cache_toCQ_data_0_BIT_5_ETC__q256 =
	      cache_toCQ_data_1[584];
    endcase
  end
  always@(cache_rsLdToDmaQ_deqP or
	  cache_rsLdToDmaQ_data_0 or cache_rsLdToDmaQ_data_1)
  begin
    case (cache_rsLdToDmaQ_deqP)
      1'd0:
	  CASE_cache_rsLdToDmaQ_deqP_0_cache_rsLdToDmaQ__ETC__q257 =
	      cache_rsLdToDmaQ_data_0[207:144];
      1'd1:
	  CASE_cache_rsLdToDmaQ_deqP_0_cache_rsLdToDmaQ__ETC__q257 =
	      cache_rsLdToDmaQ_data_1[207:144];
    endcase
  end
  always@(cache_rsLdToDmaQ_deqP or
	  cache_rsLdToDmaQ_data_0 or cache_rsLdToDmaQ_data_1)
  begin
    case (cache_rsLdToDmaQ_deqP)
      1'd0:
	  CASE_cache_rsLdToDmaQ_deqP_0_cache_rsLdToDmaQ__ETC__q258 =
	      cache_rsLdToDmaQ_data_0[143:80];
      1'd1:
	  CASE_cache_rsLdToDmaQ_deqP_0_cache_rsLdToDmaQ__ETC__q258 =
	      cache_rsLdToDmaQ_data_1[143:80];
    endcase
  end
  always@(cache_rsLdToDmaQ_deqP or
	  cache_rsLdToDmaQ_data_0 or cache_rsLdToDmaQ_data_1)
  begin
    case (cache_rsLdToDmaQ_deqP)
      1'd0:
	  CASE_cache_rsLdToDmaQ_deqP_0_cache_rsLdToDmaQ__ETC__q259 =
	      cache_rsLdToDmaQ_data_0[79:16];
      1'd1:
	  CASE_cache_rsLdToDmaQ_deqP_0_cache_rsLdToDmaQ__ETC__q259 =
	      cache_rsLdToDmaQ_data_1[79:16];
    endcase
  end
  always@(cache_toMQ_deqP or cache_toMQ_data_0 or cache_toMQ_data_1)
  begin
    case (cache_toMQ_deqP)
      1'd0:
	  CASE_cache_toMQ_deqP_0_NOT_cache_toMQ_data_0_B_ETC__q260 =
	      !cache_toMQ_data_0[640];
      1'd1:
	  CASE_cache_toMQ_deqP_0_NOT_cache_toMQ_data_0_B_ETC__q260 =
	      !cache_toMQ_data_1[640];
    endcase
  end
  always@(cache_toMQ_deqP or cache_toMQ_data_0 or cache_toMQ_data_1)
  begin
    case (cache_toMQ_deqP)
      1'd0:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_6_ETC__q261 =
	      cache_toMQ_data_0[640];
      1'd1:
	  CASE_cache_toMQ_deqP_0_cache_toMQ_data_0_BIT_6_ETC__q261 =
	      cache_toMQ_data_1[640];
    endcase
  end
  always@(cache_rsFromMQ_deqP or
	  cache_rsFromMQ_data_0 or cache_rsFromMQ_data_1)
  begin
    case (cache_rsFromMQ_deqP)
      1'd0:
	  CASE_cache_rsFromMQ_deqP_0_cache_rsFromMQ_data_ETC__q262 =
	      cache_rsFromMQ_data_0[4];
      1'd1:
	  CASE_cache_rsFromMQ_deqP_0_cache_rsFromMQ_data_ETC__q262 =
	      cache_rsFromMQ_data_1[4];
    endcase
  end
  always@(cache_rsFromMQ_deqP or
	  cache_rsFromMQ_data_0 or cache_rsFromMQ_data_1)
  begin
    case (cache_rsFromMQ_deqP)
      1'd0:
	  CASE_cache_rsFromMQ_deqP_0_NOT_cache_rsFromMQ__ETC__q263 =
	      !cache_rsFromMQ_data_0[4];
      1'd1:
	  CASE_cache_rsFromMQ_deqP_0_NOT_cache_rsFromMQ__ETC__q263 =
	      !cache_rsFromMQ_data_1[4];
    endcase
  end
  always@(cache_toMInfoQ$D_OUT or
	  cache_toMQ_full or cache_rsStToDmaIndexQ_sendToM$FULL_N)
  begin
    case (cache_toMInfoQ$D_OUT[1:0])
      2'd0:
	  CASE_cache_toMInfoQD_OUT_BITS_1_TO_0_0_NOT_ca_ETC__q264 =
	      !cache_toMQ_full;
      2'd1:
	  CASE_cache_toMInfoQD_OUT_BITS_1_TO_0_0_NOT_ca_ETC__q264 =
	      !cache_toMQ_full && cache_rsStToDmaIndexQ_sendToM$FULL_N;
      default: CASE_cache_toMInfoQD_OUT_BITS_1_TO_0_0_NOT_ca_ETC__q264 =
		   cache_toMInfoQ$D_OUT[1:0] != 2'd2 || !cache_toMQ_full;
    endcase
  end
  always@(cache_rqFromCQ_deqP or
	  cache_rqFromCQ_data_0 or cache_rqFromCQ_data_1)
  begin
    case (cache_rqFromCQ_deqP)
      1'd0:
	  CASE_cache_rqFromCQ_deqP_0_cache_rqFromCQ_data_ETC__q265 =
	      cache_rqFromCQ_data_0[9:8];
      1'd1:
	  CASE_cache_rqFromCQ_deqP_0_cache_rqFromCQ_data_ETC__q265 =
	      cache_rqFromCQ_data_1[9:8];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q266 =
	      cache_rqFromDmaQ_data_0[15:0];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q266 =
	      cache_rqFromDmaQ_data_1[15:0];
    endcase
  end
  always@(cache_rqFromDmaQ_deqP or
	  cache_rqFromDmaQ_data_0 or cache_rqFromDmaQ_data_1)
  begin
    case (cache_rqFromDmaQ_deqP)
      1'd0:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q267 =
	      cache_rqFromDmaQ_data_0[79:16];
      1'd1:
	  CASE_cache_rqFromDmaQ_deqP_0_cache_rqFromDmaQ__ETC__q267 =
	      cache_rqFromDmaQ_data_1[79:16];
    endcase
  end
  // handling of inlined registers
  always@(posedge CLK)
  begin
    if (RST_N == `BSV_RESET_VALUE)
      begin
        cache_cRqRetryIndexQ_clearReq_rl <= `BSV_ASSIGNMENT_DELAY 1'd0;
	cache_cRqRetryIndexQ_data_0 <= `BSV_ASSIGNMENT_DELAY 4'd0;
	cache_cRqRetryIndexQ_data_1 <= `BSV_ASSIGNMENT_DELAY 4'd0;
	cache_cRqRetryIndexQ_data_10 <= `BSV_ASSIGNMENT_DELAY 4'd0;
	cache_cRqRetryIndexQ_data_11 <= `BSV_ASSIGNMENT_DELAY 4'd0;
	cache_cRqRetryIndexQ_data_12 <= `BSV_ASSIGNMENT_DELAY 4'd0;
	cache_cRqRetryIndexQ_data_13 <= `BSV_ASSIGNMENT_DELAY 4'd0;
	cache_cRqRetryIndexQ_data_14 <= `BSV_ASSIGNMENT_DELAY 4'd0;
	cache_cRqRetryIndexQ_data_15 <= `BSV_ASSIGNMENT_DELAY 4'd0;
	cache_cRqRetryIndexQ_data_2 <= `BSV_ASSIGNMENT_DELAY 4'd0;
	cache_cRqRetryIndexQ_data_3 <= `BSV_ASSIGNMENT_DELAY 4'd0;
	cache_cRqRetryIndexQ_data_4 <= `BSV_ASSIGNMENT_DELAY 4'd0;
	cache_cRqRetryIndexQ_data_5 <= `BSV_ASSIGNMENT_DELAY 4'd0;
	cache_cRqRetryIndexQ_data_6 <= `BSV_ASSIGNMENT_DELAY 4'd0;
	cache_cRqRetryIndexQ_data_7 <= `BSV_ASSIGNMENT_DELAY 4'd0;
	cache_cRqRetryIndexQ_data_8 <= `BSV_ASSIGNMENT_DELAY 4'd0;
	cache_cRqRetryIndexQ_data_9 <= `BSV_ASSIGNMENT_DELAY 4'd0;
	cache_cRqRetryIndexQ_deqP <= `BSV_ASSIGNMENT_DELAY 4'd0;
	cache_cRqRetryIndexQ_deqReq_rl <= `BSV_ASSIGNMENT_DELAY 1'd0;
	cache_cRqRetryIndexQ_empty <= `BSV_ASSIGNMENT_DELAY 1'd1;
	cache_cRqRetryIndexQ_enqP <= `BSV_ASSIGNMENT_DELAY 4'd0;
	cache_cRqRetryIndexQ_enqReq_rl <= `BSV_ASSIGNMENT_DELAY 5'd10;
	cache_cRqRetryIndexQ_full <= `BSV_ASSIGNMENT_DELAY 1'd0;
	cache_doLdAfterReplace <= `BSV_ASSIGNMENT_DELAY 1'd0;
	cache_priorNewCRqSrc <= `BSV_ASSIGNMENT_DELAY 1'd0;
	cache_rqFromCQ_clearReq_rl <= `BSV_ASSIGNMENT_DELAY 1'd0;
	cache_rqFromCQ_data_0 <= `BSV_ASSIGNMENT_DELAY 74'd0;
	cache_rqFromCQ_data_1 <= `BSV_ASSIGNMENT_DELAY 74'd0;
	cache_rqFromCQ_deqP <= `BSV_ASSIGNMENT_DELAY 1'd0;
	cache_rqFromCQ_deqReq_rl <= `BSV_ASSIGNMENT_DELAY 1'd0;
	cache_rqFromCQ_empty <= `BSV_ASSIGNMENT_DELAY 1'd1;
	cache_rqFromCQ_enqP <= `BSV_ASSIGNMENT_DELAY 1'd0;
	cache_rqFromCQ_enqReq_rl <= `BSV_ASSIGNMENT_DELAY
	    75'h2AAAAAAAAAAAAAAAAAA;
	cache_rqFromCQ_full <= `BSV_ASSIGNMENT_DELAY 1'd0;
	cache_rqFromDmaQ_clearReq_rl <= `BSV_ASSIGNMENT_DELAY 1'd0;
	cache_rqFromDmaQ_data_0 <= `BSV_ASSIGNMENT_DELAY 656'd0;
	cache_rqFromDmaQ_data_1 <= `BSV_ASSIGNMENT_DELAY 656'd0;
	cache_rqFromDmaQ_deqP <= `BSV_ASSIGNMENT_DELAY 1'd0;
	cache_rqFromDmaQ_deqReq_rl <= `BSV_ASSIGNMENT_DELAY 1'd0;
	cache_rqFromDmaQ_empty <= `BSV_ASSIGNMENT_DELAY 1'd1;
	cache_rqFromDmaQ_enqP <= `BSV_ASSIGNMENT_DELAY 1'd0;
	cache_rqFromDmaQ_enqReq_rl <= `BSV_ASSIGNMENT_DELAY
	    657'h0AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
	cache_rqFromDmaQ_full <= `BSV_ASSIGNMENT_DELAY 1'd0;
	cache_rsFromCQ_clearReq_rl <= `BSV_ASSIGNMENT_DELAY 1'd0;
	cache_rsFromCQ_data_0 <= `BSV_ASSIGNMENT_DELAY
	    581'h000000000000000002AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA8;
	cache_rsFromCQ_data_1 <= `BSV_ASSIGNMENT_DELAY
	    581'h000000000000000002AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA8;
	cache_rsFromCQ_deqP <= `BSV_ASSIGNMENT_DELAY 1'd0;
	cache_rsFromCQ_deqReq_rl <= `BSV_ASSIGNMENT_DELAY 1'd0;
	cache_rsFromCQ_empty <= `BSV_ASSIGNMENT_DELAY 1'd1;
	cache_rsFromCQ_enqP <= `BSV_ASSIGNMENT_DELAY 1'd0;
	cache_rsFromCQ_enqReq_rl <= `BSV_ASSIGNMENT_DELAY
	    582'h0AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
	cache_rsFromCQ_full <= `BSV_ASSIGNMENT_DELAY 1'd0;
	cache_rsFromMQ_clearReq_rl <= `BSV_ASSIGNMENT_DELAY 1'd0;
	cache_rsFromMQ_data_0 <= `BSV_ASSIGNMENT_DELAY 517'd0;
	cache_rsFromMQ_data_1 <= `BSV_ASSIGNMENT_DELAY 517'd0;
	cache_rsFromMQ_deqP <= `BSV_ASSIGNMENT_DELAY 1'd0;
	cache_rsFromMQ_deqReq_rl <= `BSV_ASSIGNMENT_DELAY 1'd0;
	cache_rsFromMQ_empty <= `BSV_ASSIGNMENT_DELAY 1'd1;
	cache_rsFromMQ_enqP <= `BSV_ASSIGNMENT_DELAY 1'd0;
	cache_rsFromMQ_enqReq_rl <= `BSV_ASSIGNMENT_DELAY
	    518'h0AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
	cache_rsFromMQ_full <= `BSV_ASSIGNMENT_DELAY 1'd0;
	cache_rsLdToDmaQ_clearReq_rl <= `BSV_ASSIGNMENT_DELAY 1'd0;
	cache_rsLdToDmaQ_data_0 <= `BSV_ASSIGNMENT_DELAY 528'd0;
	cache_rsLdToDmaQ_data_1 <= `BSV_ASSIGNMENT_DELAY 528'd0;
	cache_rsLdToDmaQ_deqP <= `BSV_ASSIGNMENT_DELAY 1'd0;
	cache_rsLdToDmaQ_deqReq_rl <= `BSV_ASSIGNMENT_DELAY 1'd0;
	cache_rsLdToDmaQ_empty <= `BSV_ASSIGNMENT_DELAY 1'd1;
	cache_rsLdToDmaQ_enqP <= `BSV_ASSIGNMENT_DELAY 1'd0;
	cache_rsLdToDmaQ_enqReq_rl <= `BSV_ASSIGNMENT_DELAY
	    529'h0AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
	cache_rsLdToDmaQ_full <= `BSV_ASSIGNMENT_DELAY 1'd0;
	cache_rsStToDmaQ_clearReq_rl <= `BSV_ASSIGNMENT_DELAY 1'd0;
	cache_rsStToDmaQ_data_0 <= `BSV_ASSIGNMENT_DELAY 16'd0;
	cache_rsStToDmaQ_data_1 <= `BSV_ASSIGNMENT_DELAY 16'd0;
	cache_rsStToDmaQ_deqP <= `BSV_ASSIGNMENT_DELAY 1'd0;
	cache_rsStToDmaQ_deqReq_rl <= `BSV_ASSIGNMENT_DELAY 1'd0;
	cache_rsStToDmaQ_empty <= `BSV_ASSIGNMENT_DELAY 1'd1;
	cache_rsStToDmaQ_enqP <= `BSV_ASSIGNMENT_DELAY 1'd0;
	cache_rsStToDmaQ_enqReq_rl <= `BSV_ASSIGNMENT_DELAY 17'd43690;
	cache_rsStToDmaQ_full <= `BSV_ASSIGNMENT_DELAY 1'd0;
	cache_rsToCIndexQ_clearReq_rl <= `BSV_ASSIGNMENT_DELAY 1'd0;
	cache_rsToCIndexQ_data_0 <= `BSV_ASSIGNMENT_DELAY 6'd0;
	cache_rsToCIndexQ_data_1 <= `BSV_ASSIGNMENT_DELAY 6'd0;
	cache_rsToCIndexQ_data_10 <= `BSV_ASSIGNMENT_DELAY 6'd0;
	cache_rsToCIndexQ_data_11 <= `BSV_ASSIGNMENT_DELAY 6'd0;
	cache_rsToCIndexQ_data_12 <= `BSV_ASSIGNMENT_DELAY 6'd0;
	cache_rsToCIndexQ_data_13 <= `BSV_ASSIGNMENT_DELAY 6'd0;
	cache_rsToCIndexQ_data_14 <= `BSV_ASSIGNMENT_DELAY 6'd0;
	cache_rsToCIndexQ_data_15 <= `BSV_ASSIGNMENT_DELAY 6'd0;
	cache_rsToCIndexQ_data_2 <= `BSV_ASSIGNMENT_DELAY 6'd0;
	cache_rsToCIndexQ_data_3 <= `BSV_ASSIGNMENT_DELAY 6'd0;
	cache_rsToCIndexQ_data_4 <= `BSV_ASSIGNMENT_DELAY 6'd0;
	cache_rsToCIndexQ_data_5 <= `BSV_ASSIGNMENT_DELAY 6'd0;
	cache_rsToCIndexQ_data_6 <= `BSV_ASSIGNMENT_DELAY 6'd0;
	cache_rsToCIndexQ_data_7 <= `BSV_ASSIGNMENT_DELAY 6'd0;
	cache_rsToCIndexQ_data_8 <= `BSV_ASSIGNMENT_DELAY 6'd0;
	cache_rsToCIndexQ_data_9 <= `BSV_ASSIGNMENT_DELAY 6'd0;
	cache_rsToCIndexQ_deqP <= `BSV_ASSIGNMENT_DELAY 4'd0;
	cache_rsToCIndexQ_deqReq_rl <= `BSV_ASSIGNMENT_DELAY 1'd0;
	cache_rsToCIndexQ_empty <= `BSV_ASSIGNMENT_DELAY 1'd1;
	cache_rsToCIndexQ_enqP <= `BSV_ASSIGNMENT_DELAY 4'd0;
	cache_rsToCIndexQ_enqReq_rl <= `BSV_ASSIGNMENT_DELAY 7'd42;
	cache_rsToCIndexQ_full <= `BSV_ASSIGNMENT_DELAY 1'd0;
	cache_toCQ_clearReq_rl <= `BSV_ASSIGNMENT_DELAY 1'd0;
	cache_toCQ_data_0 <= `BSV_ASSIGNMENT_DELAY
	    585'h0AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA00000000000000000;
	cache_toCQ_data_1 <= `BSV_ASSIGNMENT_DELAY
	    585'h0AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA00000000000000000;
	cache_toCQ_deqP <= `BSV_ASSIGNMENT_DELAY 1'd0;
	cache_toCQ_deqReq_rl <= `BSV_ASSIGNMENT_DELAY 1'd0;
	cache_toCQ_empty <= `BSV_ASSIGNMENT_DELAY 1'd1;
	cache_toCQ_enqP <= `BSV_ASSIGNMENT_DELAY 1'd0;
	cache_toCQ_enqReq_rl <= `BSV_ASSIGNMENT_DELAY
	    586'h0AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
	cache_toCQ_full <= `BSV_ASSIGNMENT_DELAY 1'd0;
	cache_toMQ_clearReq_rl <= `BSV_ASSIGNMENT_DELAY 1'd0;
	cache_toMQ_data_0 <= `BSV_ASSIGNMENT_DELAY
	    641'h05555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555400000000000000000;
	cache_toMQ_data_1 <= `BSV_ASSIGNMENT_DELAY
	    641'h05555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555555400000000000000000;
	cache_toMQ_deqP <= `BSV_ASSIGNMENT_DELAY 1'd0;
	cache_toMQ_deqReq_rl <= `BSV_ASSIGNMENT_DELAY 1'd0;
	cache_toMQ_empty <= `BSV_ASSIGNMENT_DELAY 1'd1;
	cache_toMQ_enqP <= `BSV_ASSIGNMENT_DELAY 1'd0;
	cache_toMQ_enqReq_rl <= `BSV_ASSIGNMENT_DELAY
	    642'h0AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
	cache_toMQ_full <= `BSV_ASSIGNMENT_DELAY 1'd0;
	cache_whichCRq <= `BSV_ASSIGNMENT_DELAY 4'd0;
	perfReqQ_clearReq_rl <= `BSV_ASSIGNMENT_DELAY 1'd0;
	perfReqQ_data_0 <= `BSV_ASSIGNMENT_DELAY 4'd0;
	perfReqQ_deqReq_rl <= `BSV_ASSIGNMENT_DELAY 1'd0;
	perfReqQ_empty <= `BSV_ASSIGNMENT_DELAY 1'd1;
	perfReqQ_enqReq_rl <= `BSV_ASSIGNMENT_DELAY 5'd10;
	perfReqQ_full <= `BSV_ASSIGNMENT_DELAY 1'd0;
      end
    else
      begin
        if (cache_cRqRetryIndexQ_clearReq_rl$EN)
	  cache_cRqRetryIndexQ_clearReq_rl <= `BSV_ASSIGNMENT_DELAY
	      cache_cRqRetryIndexQ_clearReq_rl$D_IN;
	if (cache_cRqRetryIndexQ_data_0$EN)
	  cache_cRqRetryIndexQ_data_0 <= `BSV_ASSIGNMENT_DELAY
	      cache_cRqRetryIndexQ_data_0$D_IN;
	if (cache_cRqRetryIndexQ_data_1$EN)
	  cache_cRqRetryIndexQ_data_1 <= `BSV_ASSIGNMENT_DELAY
	      cache_cRqRetryIndexQ_data_1$D_IN;
	if (cache_cRqRetryIndexQ_data_10$EN)
	  cache_cRqRetryIndexQ_data_10 <= `BSV_ASSIGNMENT_DELAY
	      cache_cRqRetryIndexQ_data_10$D_IN;
	if (cache_cRqRetryIndexQ_data_11$EN)
	  cache_cRqRetryIndexQ_data_11 <= `BSV_ASSIGNMENT_DELAY
	      cache_cRqRetryIndexQ_data_11$D_IN;
	if (cache_cRqRetryIndexQ_data_12$EN)
	  cache_cRqRetryIndexQ_data_12 <= `BSV_ASSIGNMENT_DELAY
	      cache_cRqRetryIndexQ_data_12$D_IN;
	if (cache_cRqRetryIndexQ_data_13$EN)
	  cache_cRqRetryIndexQ_data_13 <= `BSV_ASSIGNMENT_DELAY
	      cache_cRqRetryIndexQ_data_13$D_IN;
	if (cache_cRqRetryIndexQ_data_14$EN)
	  cache_cRqRetryIndexQ_data_14 <= `BSV_ASSIGNMENT_DELAY
	      cache_cRqRetryIndexQ_data_14$D_IN;
	if (cache_cRqRetryIndexQ_data_15$EN)
	  cache_cRqRetryIndexQ_data_15 <= `BSV_ASSIGNMENT_DELAY
	      cache_cRqRetryIndexQ_data_15$D_IN;
	if (cache_cRqRetryIndexQ_data_2$EN)
	  cache_cRqRetryIndexQ_data_2 <= `BSV_ASSIGNMENT_DELAY
	      cache_cRqRetryIndexQ_data_2$D_IN;
	if (cache_cRqRetryIndexQ_data_3$EN)
	  cache_cRqRetryIndexQ_data_3 <= `BSV_ASSIGNMENT_DELAY
	      cache_cRqRetryIndexQ_data_3$D_IN;
	if (cache_cRqRetryIndexQ_data_4$EN)
	  cache_cRqRetryIndexQ_data_4 <= `BSV_ASSIGNMENT_DELAY
	      cache_cRqRetryIndexQ_data_4$D_IN;
	if (cache_cRqRetryIndexQ_data_5$EN)
	  cache_cRqRetryIndexQ_data_5 <= `BSV_ASSIGNMENT_DELAY
	      cache_cRqRetryIndexQ_data_5$D_IN;
	if (cache_cRqRetryIndexQ_data_6$EN)
	  cache_cRqRetryIndexQ_data_6 <= `BSV_ASSIGNMENT_DELAY
	      cache_cRqRetryIndexQ_data_6$D_IN;
	if (cache_cRqRetryIndexQ_data_7$EN)
	  cache_cRqRetryIndexQ_data_7 <= `BSV_ASSIGNMENT_DELAY
	      cache_cRqRetryIndexQ_data_7$D_IN;
	if (cache_cRqRetryIndexQ_data_8$EN)
	  cache_cRqRetryIndexQ_data_8 <= `BSV_ASSIGNMENT_DELAY
	      cache_cRqRetryIndexQ_data_8$D_IN;
	if (cache_cRqRetryIndexQ_data_9$EN)
	  cache_cRqRetryIndexQ_data_9 <= `BSV_ASSIGNMENT_DELAY
	      cache_cRqRetryIndexQ_data_9$D_IN;
	if (cache_cRqRetryIndexQ_deqP$EN)
	  cache_cRqRetryIndexQ_deqP <= `BSV_ASSIGNMENT_DELAY
	      cache_cRqRetryIndexQ_deqP$D_IN;
	if (cache_cRqRetryIndexQ_deqReq_rl$EN)
	  cache_cRqRetryIndexQ_deqReq_rl <= `BSV_ASSIGNMENT_DELAY
	      cache_cRqRetryIndexQ_deqReq_rl$D_IN;
	if (cache_cRqRetryIndexQ_empty$EN)
	  cache_cRqRetryIndexQ_empty <= `BSV_ASSIGNMENT_DELAY
	      cache_cRqRetryIndexQ_empty$D_IN;
	if (cache_cRqRetryIndexQ_enqP$EN)
	  cache_cRqRetryIndexQ_enqP <= `BSV_ASSIGNMENT_DELAY
	      cache_cRqRetryIndexQ_enqP$D_IN;
	if (cache_cRqRetryIndexQ_enqReq_rl$EN)
	  cache_cRqRetryIndexQ_enqReq_rl <= `BSV_ASSIGNMENT_DELAY
	      cache_cRqRetryIndexQ_enqReq_rl$D_IN;
	if (cache_cRqRetryIndexQ_full$EN)
	  cache_cRqRetryIndexQ_full <= `BSV_ASSIGNMENT_DELAY
	      cache_cRqRetryIndexQ_full$D_IN;
	if (cache_doLdAfterReplace$EN)
	  cache_doLdAfterReplace <= `BSV_ASSIGNMENT_DELAY
	      cache_doLdAfterReplace$D_IN;
	if (cache_priorNewCRqSrc$EN)
	  cache_priorNewCRqSrc <= `BSV_ASSIGNMENT_DELAY
	      cache_priorNewCRqSrc$D_IN;
	if (cache_rqFromCQ_clearReq_rl$EN)
	  cache_rqFromCQ_clearReq_rl <= `BSV_ASSIGNMENT_DELAY
	      cache_rqFromCQ_clearReq_rl$D_IN;
	if (cache_rqFromCQ_data_0$EN)
	  cache_rqFromCQ_data_0 <= `BSV_ASSIGNMENT_DELAY
	      cache_rqFromCQ_data_0$D_IN;
	if (cache_rqFromCQ_data_1$EN)
	  cache_rqFromCQ_data_1 <= `BSV_ASSIGNMENT_DELAY
	      cache_rqFromCQ_data_1$D_IN;
	if (cache_rqFromCQ_deqP$EN)
	  cache_rqFromCQ_deqP <= `BSV_ASSIGNMENT_DELAY
	      cache_rqFromCQ_deqP$D_IN;
	if (cache_rqFromCQ_deqReq_rl$EN)
	  cache_rqFromCQ_deqReq_rl <= `BSV_ASSIGNMENT_DELAY
	      cache_rqFromCQ_deqReq_rl$D_IN;
	if (cache_rqFromCQ_empty$EN)
	  cache_rqFromCQ_empty <= `BSV_ASSIGNMENT_DELAY
	      cache_rqFromCQ_empty$D_IN;
	if (cache_rqFromCQ_enqP$EN)
	  cache_rqFromCQ_enqP <= `BSV_ASSIGNMENT_DELAY
	      cache_rqFromCQ_enqP$D_IN;
	if (cache_rqFromCQ_enqReq_rl$EN)
	  cache_rqFromCQ_enqReq_rl <= `BSV_ASSIGNMENT_DELAY
	      cache_rqFromCQ_enqReq_rl$D_IN;
	if (cache_rqFromCQ_full$EN)
	  cache_rqFromCQ_full <= `BSV_ASSIGNMENT_DELAY
	      cache_rqFromCQ_full$D_IN;
	if (cache_rqFromDmaQ_clearReq_rl$EN)
	  cache_rqFromDmaQ_clearReq_rl <= `BSV_ASSIGNMENT_DELAY
	      cache_rqFromDmaQ_clearReq_rl$D_IN;
	if (cache_rqFromDmaQ_data_0$EN)
	  cache_rqFromDmaQ_data_0 <= `BSV_ASSIGNMENT_DELAY
	      cache_rqFromDmaQ_data_0$D_IN;
	if (cache_rqFromDmaQ_data_1$EN)
	  cache_rqFromDmaQ_data_1 <= `BSV_ASSIGNMENT_DELAY
	      cache_rqFromDmaQ_data_1$D_IN;
	if (cache_rqFromDmaQ_deqP$EN)
	  cache_rqFromDmaQ_deqP <= `BSV_ASSIGNMENT_DELAY
	      cache_rqFromDmaQ_deqP$D_IN;
	if (cache_rqFromDmaQ_deqReq_rl$EN)
	  cache_rqFromDmaQ_deqReq_rl <= `BSV_ASSIGNMENT_DELAY
	      cache_rqFromDmaQ_deqReq_rl$D_IN;
	if (cache_rqFromDmaQ_empty$EN)
	  cache_rqFromDmaQ_empty <= `BSV_ASSIGNMENT_DELAY
	      cache_rqFromDmaQ_empty$D_IN;
	if (cache_rqFromDmaQ_enqP$EN)
	  cache_rqFromDmaQ_enqP <= `BSV_ASSIGNMENT_DELAY
	      cache_rqFromDmaQ_enqP$D_IN;
	if (cache_rqFromDmaQ_enqReq_rl$EN)
	  cache_rqFromDmaQ_enqReq_rl <= `BSV_ASSIGNMENT_DELAY
	      cache_rqFromDmaQ_enqReq_rl$D_IN;
	if (cache_rqFromDmaQ_full$EN)
	  cache_rqFromDmaQ_full <= `BSV_ASSIGNMENT_DELAY
	      cache_rqFromDmaQ_full$D_IN;
	if (cache_rsFromCQ_clearReq_rl$EN)
	  cache_rsFromCQ_clearReq_rl <= `BSV_ASSIGNMENT_DELAY
	      cache_rsFromCQ_clearReq_rl$D_IN;
	if (cache_rsFromCQ_data_0$EN)
	  cache_rsFromCQ_data_0 <= `BSV_ASSIGNMENT_DELAY
	      cache_rsFromCQ_data_0$D_IN;
	if (cache_rsFromCQ_data_1$EN)
	  cache_rsFromCQ_data_1 <= `BSV_ASSIGNMENT_DELAY
	      cache_rsFromCQ_data_1$D_IN;
	if (cache_rsFromCQ_deqP$EN)
	  cache_rsFromCQ_deqP <= `BSV_ASSIGNMENT_DELAY
	      cache_rsFromCQ_deqP$D_IN;
	if (cache_rsFromCQ_deqReq_rl$EN)
	  cache_rsFromCQ_deqReq_rl <= `BSV_ASSIGNMENT_DELAY
	      cache_rsFromCQ_deqReq_rl$D_IN;
	if (cache_rsFromCQ_empty$EN)
	  cache_rsFromCQ_empty <= `BSV_ASSIGNMENT_DELAY
	      cache_rsFromCQ_empty$D_IN;
	if (cache_rsFromCQ_enqP$EN)
	  cache_rsFromCQ_enqP <= `BSV_ASSIGNMENT_DELAY
	      cache_rsFromCQ_enqP$D_IN;
	if (cache_rsFromCQ_enqReq_rl$EN)
	  cache_rsFromCQ_enqReq_rl <= `BSV_ASSIGNMENT_DELAY
	      cache_rsFromCQ_enqReq_rl$D_IN;
	if (cache_rsFromCQ_full$EN)
	  cache_rsFromCQ_full <= `BSV_ASSIGNMENT_DELAY
	      cache_rsFromCQ_full$D_IN;
	if (cache_rsFromMQ_clearReq_rl$EN)
	  cache_rsFromMQ_clearReq_rl <= `BSV_ASSIGNMENT_DELAY
	      cache_rsFromMQ_clearReq_rl$D_IN;
	if (cache_rsFromMQ_data_0$EN)
	  cache_rsFromMQ_data_0 <= `BSV_ASSIGNMENT_DELAY
	      cache_rsFromMQ_data_0$D_IN;
	if (cache_rsFromMQ_data_1$EN)
	  cache_rsFromMQ_data_1 <= `BSV_ASSIGNMENT_DELAY
	      cache_rsFromMQ_data_1$D_IN;
	if (cache_rsFromMQ_deqP$EN)
	  cache_rsFromMQ_deqP <= `BSV_ASSIGNMENT_DELAY
	      cache_rsFromMQ_deqP$D_IN;
	if (cache_rsFromMQ_deqReq_rl$EN)
	  cache_rsFromMQ_deqReq_rl <= `BSV_ASSIGNMENT_DELAY
	      cache_rsFromMQ_deqReq_rl$D_IN;
	if (cache_rsFromMQ_empty$EN)
	  cache_rsFromMQ_empty <= `BSV_ASSIGNMENT_DELAY
	      cache_rsFromMQ_empty$D_IN;
	if (cache_rsFromMQ_enqP$EN)
	  cache_rsFromMQ_enqP <= `BSV_ASSIGNMENT_DELAY
	      cache_rsFromMQ_enqP$D_IN;
	if (cache_rsFromMQ_enqReq_rl$EN)
	  cache_rsFromMQ_enqReq_rl <= `BSV_ASSIGNMENT_DELAY
	      cache_rsFromMQ_enqReq_rl$D_IN;
	if (cache_rsFromMQ_full$EN)
	  cache_rsFromMQ_full <= `BSV_ASSIGNMENT_DELAY
	      cache_rsFromMQ_full$D_IN;
	if (cache_rsLdToDmaQ_clearReq_rl$EN)
	  cache_rsLdToDmaQ_clearReq_rl <= `BSV_ASSIGNMENT_DELAY
	      cache_rsLdToDmaQ_clearReq_rl$D_IN;
	if (cache_rsLdToDmaQ_data_0$EN)
	  cache_rsLdToDmaQ_data_0 <= `BSV_ASSIGNMENT_DELAY
	      cache_rsLdToDmaQ_data_0$D_IN;
	if (cache_rsLdToDmaQ_data_1$EN)
	  cache_rsLdToDmaQ_data_1 <= `BSV_ASSIGNMENT_DELAY
	      cache_rsLdToDmaQ_data_1$D_IN;
	if (cache_rsLdToDmaQ_deqP$EN)
	  cache_rsLdToDmaQ_deqP <= `BSV_ASSIGNMENT_DELAY
	      cache_rsLdToDmaQ_deqP$D_IN;
	if (cache_rsLdToDmaQ_deqReq_rl$EN)
	  cache_rsLdToDmaQ_deqReq_rl <= `BSV_ASSIGNMENT_DELAY
	      cache_rsLdToDmaQ_deqReq_rl$D_IN;
	if (cache_rsLdToDmaQ_empty$EN)
	  cache_rsLdToDmaQ_empty <= `BSV_ASSIGNMENT_DELAY
	      cache_rsLdToDmaQ_empty$D_IN;
	if (cache_rsLdToDmaQ_enqP$EN)
	  cache_rsLdToDmaQ_enqP <= `BSV_ASSIGNMENT_DELAY
	      cache_rsLdToDmaQ_enqP$D_IN;
	if (cache_rsLdToDmaQ_enqReq_rl$EN)
	  cache_rsLdToDmaQ_enqReq_rl <= `BSV_ASSIGNMENT_DELAY
	      cache_rsLdToDmaQ_enqReq_rl$D_IN;
	if (cache_rsLdToDmaQ_full$EN)
	  cache_rsLdToDmaQ_full <= `BSV_ASSIGNMENT_DELAY
	      cache_rsLdToDmaQ_full$D_IN;
	if (cache_rsStToDmaQ_clearReq_rl$EN)
	  cache_rsStToDmaQ_clearReq_rl <= `BSV_ASSIGNMENT_DELAY
	      cache_rsStToDmaQ_clearReq_rl$D_IN;
	if (cache_rsStToDmaQ_data_0$EN)
	  cache_rsStToDmaQ_data_0 <= `BSV_ASSIGNMENT_DELAY
	      cache_rsStToDmaQ_data_0$D_IN;
	if (cache_rsStToDmaQ_data_1$EN)
	  cache_rsStToDmaQ_data_1 <= `BSV_ASSIGNMENT_DELAY
	      cache_rsStToDmaQ_data_1$D_IN;
	if (cache_rsStToDmaQ_deqP$EN)
	  cache_rsStToDmaQ_deqP <= `BSV_ASSIGNMENT_DELAY
	      cache_rsStToDmaQ_deqP$D_IN;
	if (cache_rsStToDmaQ_deqReq_rl$EN)
	  cache_rsStToDmaQ_deqReq_rl <= `BSV_ASSIGNMENT_DELAY
	      cache_rsStToDmaQ_deqReq_rl$D_IN;
	if (cache_rsStToDmaQ_empty$EN)
	  cache_rsStToDmaQ_empty <= `BSV_ASSIGNMENT_DELAY
	      cache_rsStToDmaQ_empty$D_IN;
	if (cache_rsStToDmaQ_enqP$EN)
	  cache_rsStToDmaQ_enqP <= `BSV_ASSIGNMENT_DELAY
	      cache_rsStToDmaQ_enqP$D_IN;
	if (cache_rsStToDmaQ_enqReq_rl$EN)
	  cache_rsStToDmaQ_enqReq_rl <= `BSV_ASSIGNMENT_DELAY
	      cache_rsStToDmaQ_enqReq_rl$D_IN;
	if (cache_rsStToDmaQ_full$EN)
	  cache_rsStToDmaQ_full <= `BSV_ASSIGNMENT_DELAY
	      cache_rsStToDmaQ_full$D_IN;
	if (cache_rsToCIndexQ_clearReq_rl$EN)
	  cache_rsToCIndexQ_clearReq_rl <= `BSV_ASSIGNMENT_DELAY
	      cache_rsToCIndexQ_clearReq_rl$D_IN;
	if (cache_rsToCIndexQ_data_0$EN)
	  cache_rsToCIndexQ_data_0 <= `BSV_ASSIGNMENT_DELAY
	      cache_rsToCIndexQ_data_0$D_IN;
	if (cache_rsToCIndexQ_data_1$EN)
	  cache_rsToCIndexQ_data_1 <= `BSV_ASSIGNMENT_DELAY
	      cache_rsToCIndexQ_data_1$D_IN;
	if (cache_rsToCIndexQ_data_10$EN)
	  cache_rsToCIndexQ_data_10 <= `BSV_ASSIGNMENT_DELAY
	      cache_rsToCIndexQ_data_10$D_IN;
	if (cache_rsToCIndexQ_data_11$EN)
	  cache_rsToCIndexQ_data_11 <= `BSV_ASSIGNMENT_DELAY
	      cache_rsToCIndexQ_data_11$D_IN;
	if (cache_rsToCIndexQ_data_12$EN)
	  cache_rsToCIndexQ_data_12 <= `BSV_ASSIGNMENT_DELAY
	      cache_rsToCIndexQ_data_12$D_IN;
	if (cache_rsToCIndexQ_data_13$EN)
	  cache_rsToCIndexQ_data_13 <= `BSV_ASSIGNMENT_DELAY
	      cache_rsToCIndexQ_data_13$D_IN;
	if (cache_rsToCIndexQ_data_14$EN)
	  cache_rsToCIndexQ_data_14 <= `BSV_ASSIGNMENT_DELAY
	      cache_rsToCIndexQ_data_14$D_IN;
	if (cache_rsToCIndexQ_data_15$EN)
	  cache_rsToCIndexQ_data_15 <= `BSV_ASSIGNMENT_DELAY
	      cache_rsToCIndexQ_data_15$D_IN;
	if (cache_rsToCIndexQ_data_2$EN)
	  cache_rsToCIndexQ_data_2 <= `BSV_ASSIGNMENT_DELAY
	      cache_rsToCIndexQ_data_2$D_IN;
	if (cache_rsToCIndexQ_data_3$EN)
	  cache_rsToCIndexQ_data_3 <= `BSV_ASSIGNMENT_DELAY
	      cache_rsToCIndexQ_data_3$D_IN;
	if (cache_rsToCIndexQ_data_4$EN)
	  cache_rsToCIndexQ_data_4 <= `BSV_ASSIGNMENT_DELAY
	      cache_rsToCIndexQ_data_4$D_IN;
	if (cache_rsToCIndexQ_data_5$EN)
	  cache_rsToCIndexQ_data_5 <= `BSV_ASSIGNMENT_DELAY
	      cache_rsToCIndexQ_data_5$D_IN;
	if (cache_rsToCIndexQ_data_6$EN)
	  cache_rsToCIndexQ_data_6 <= `BSV_ASSIGNMENT_DELAY
	      cache_rsToCIndexQ_data_6$D_IN;
	if (cache_rsToCIndexQ_data_7$EN)
	  cache_rsToCIndexQ_data_7 <= `BSV_ASSIGNMENT_DELAY
	      cache_rsToCIndexQ_data_7$D_IN;
	if (cache_rsToCIndexQ_data_8$EN)
	  cache_rsToCIndexQ_data_8 <= `BSV_ASSIGNMENT_DELAY
	      cache_rsToCIndexQ_data_8$D_IN;
	if (cache_rsToCIndexQ_data_9$EN)
	  cache_rsToCIndexQ_data_9 <= `BSV_ASSIGNMENT_DELAY
	      cache_rsToCIndexQ_data_9$D_IN;
	if (cache_rsToCIndexQ_deqP$EN)
	  cache_rsToCIndexQ_deqP <= `BSV_ASSIGNMENT_DELAY
	      cache_rsToCIndexQ_deqP$D_IN;
	if (cache_rsToCIndexQ_deqReq_rl$EN)
	  cache_rsToCIndexQ_deqReq_rl <= `BSV_ASSIGNMENT_DELAY
	      cache_rsToCIndexQ_deqReq_rl$D_IN;
	if (cache_rsToCIndexQ_empty$EN)
	  cache_rsToCIndexQ_empty <= `BSV_ASSIGNMENT_DELAY
	      cache_rsToCIndexQ_empty$D_IN;
	if (cache_rsToCIndexQ_enqP$EN)
	  cache_rsToCIndexQ_enqP <= `BSV_ASSIGNMENT_DELAY
	      cache_rsToCIndexQ_enqP$D_IN;
	if (cache_rsToCIndexQ_enqReq_rl$EN)
	  cache_rsToCIndexQ_enqReq_rl <= `BSV_ASSIGNMENT_DELAY
	      cache_rsToCIndexQ_enqReq_rl$D_IN;
	if (cache_rsToCIndexQ_full$EN)
	  cache_rsToCIndexQ_full <= `BSV_ASSIGNMENT_DELAY
	      cache_rsToCIndexQ_full$D_IN;
	if (cache_toCQ_clearReq_rl$EN)
	  cache_toCQ_clearReq_rl <= `BSV_ASSIGNMENT_DELAY
	      cache_toCQ_clearReq_rl$D_IN;
	if (cache_toCQ_data_0$EN)
	  cache_toCQ_data_0 <= `BSV_ASSIGNMENT_DELAY cache_toCQ_data_0$D_IN;
	if (cache_toCQ_data_1$EN)
	  cache_toCQ_data_1 <= `BSV_ASSIGNMENT_DELAY cache_toCQ_data_1$D_IN;
	if (cache_toCQ_deqP$EN)
	  cache_toCQ_deqP <= `BSV_ASSIGNMENT_DELAY cache_toCQ_deqP$D_IN;
	if (cache_toCQ_deqReq_rl$EN)
	  cache_toCQ_deqReq_rl <= `BSV_ASSIGNMENT_DELAY
	      cache_toCQ_deqReq_rl$D_IN;
	if (cache_toCQ_empty$EN)
	  cache_toCQ_empty <= `BSV_ASSIGNMENT_DELAY cache_toCQ_empty$D_IN;
	if (cache_toCQ_enqP$EN)
	  cache_toCQ_enqP <= `BSV_ASSIGNMENT_DELAY cache_toCQ_enqP$D_IN;
	if (cache_toCQ_enqReq_rl$EN)
	  cache_toCQ_enqReq_rl <= `BSV_ASSIGNMENT_DELAY
	      cache_toCQ_enqReq_rl$D_IN;
	if (cache_toCQ_full$EN)
	  cache_toCQ_full <= `BSV_ASSIGNMENT_DELAY cache_toCQ_full$D_IN;
	if (cache_toMQ_clearReq_rl$EN)
	  cache_toMQ_clearReq_rl <= `BSV_ASSIGNMENT_DELAY
	      cache_toMQ_clearReq_rl$D_IN;
	if (cache_toMQ_data_0$EN)
	  cache_toMQ_data_0 <= `BSV_ASSIGNMENT_DELAY cache_toMQ_data_0$D_IN;
	if (cache_toMQ_data_1$EN)
	  cache_toMQ_data_1 <= `BSV_ASSIGNMENT_DELAY cache_toMQ_data_1$D_IN;
	if (cache_toMQ_deqP$EN)
	  cache_toMQ_deqP <= `BSV_ASSIGNMENT_DELAY cache_toMQ_deqP$D_IN;
	if (cache_toMQ_deqReq_rl$EN)
	  cache_toMQ_deqReq_rl <= `BSV_ASSIGNMENT_DELAY
	      cache_toMQ_deqReq_rl$D_IN;
	if (cache_toMQ_empty$EN)
	  cache_toMQ_empty <= `BSV_ASSIGNMENT_DELAY cache_toMQ_empty$D_IN;
	if (cache_toMQ_enqP$EN)
	  cache_toMQ_enqP <= `BSV_ASSIGNMENT_DELAY cache_toMQ_enqP$D_IN;
	if (cache_toMQ_enqReq_rl$EN)
	  cache_toMQ_enqReq_rl <= `BSV_ASSIGNMENT_DELAY
	      cache_toMQ_enqReq_rl$D_IN;
	if (cache_toMQ_full$EN)
	  cache_toMQ_full <= `BSV_ASSIGNMENT_DELAY cache_toMQ_full$D_IN;
	if (cache_whichCRq$EN)
	  cache_whichCRq <= `BSV_ASSIGNMENT_DELAY cache_whichCRq$D_IN;
	if (perfReqQ_clearReq_rl$EN)
	  perfReqQ_clearReq_rl <= `BSV_ASSIGNMENT_DELAY
	      perfReqQ_clearReq_rl$D_IN;
	if (perfReqQ_data_0$EN)
	  perfReqQ_data_0 <= `BSV_ASSIGNMENT_DELAY perfReqQ_data_0$D_IN;
	if (perfReqQ_deqReq_rl$EN)
	  perfReqQ_deqReq_rl <= `BSV_ASSIGNMENT_DELAY perfReqQ_deqReq_rl$D_IN;
	if (perfReqQ_empty$EN)
	  perfReqQ_empty <= `BSV_ASSIGNMENT_DELAY perfReqQ_empty$D_IN;
	if (perfReqQ_enqReq_rl$EN)
	  perfReqQ_enqReq_rl <= `BSV_ASSIGNMENT_DELAY perfReqQ_enqReq_rl$D_IN;
	if (perfReqQ_full$EN)
	  perfReqQ_full <= `BSV_ASSIGNMENT_DELAY perfReqQ_full$D_IN;
      end
  end
  // synopsys translate_off
  `ifdef BSV_NO_INITIAL_BLOCKS
  `else // not BSV_NO_INITIAL_BLOCKS
  initial
  begin
    cache_cRqRetryIndexQ_clearReq_rl = 1'h0;
    cache_cRqRetryIndexQ_data_0 = 4'hA;
    cache_cRqRetryIndexQ_data_1 = 4'hA;
    cache_cRqRetryIndexQ_data_10 = 4'hA;
    cache_cRqRetryIndexQ_data_11 = 4'hA;
    cache_cRqRetryIndexQ_data_12 = 4'hA;
    cache_cRqRetryIndexQ_data_13 = 4'hA;
    cache_cRqRetryIndexQ_data_14 = 4'hA;
    cache_cRqRetryIndexQ_data_15 = 4'hA;
    cache_cRqRetryIndexQ_data_2 = 4'hA;
    cache_cRqRetryIndexQ_data_3 = 4'hA;
    cache_cRqRetryIndexQ_data_4 = 4'hA;
    cache_cRqRetryIndexQ_data_5 = 4'hA;
    cache_cRqRetryIndexQ_data_6 = 4'hA;
    cache_cRqRetryIndexQ_data_7 = 4'hA;
    cache_cRqRetryIndexQ_data_8 = 4'hA;
    cache_cRqRetryIndexQ_data_9 = 4'hA;
    cache_cRqRetryIndexQ_deqP = 4'hA;
    cache_cRqRetryIndexQ_deqReq_rl = 1'h0;
    cache_cRqRetryIndexQ_empty = 1'h0;
    cache_cRqRetryIndexQ_enqP = 4'hA;
    cache_cRqRetryIndexQ_enqReq_rl = 5'h0A;
    cache_cRqRetryIndexQ_full = 1'h0;
    cache_doLdAfterReplace = 1'h0;
    cache_priorNewCRqSrc = 1'h0;
    cache_rqFromCQ_clearReq_rl = 1'h0;
    cache_rqFromCQ_data_0 = 74'h2AAAAAAAAAAAAAAAAAA;
    cache_rqFromCQ_data_1 = 74'h2AAAAAAAAAAAAAAAAAA;
    cache_rqFromCQ_deqP = 1'h0;
    cache_rqFromCQ_deqReq_rl = 1'h0;
    cache_rqFromCQ_empty = 1'h0;
    cache_rqFromCQ_enqP = 1'h0;
    cache_rqFromCQ_enqReq_rl = 75'h2AAAAAAAAAAAAAAAAAA;
    cache_rqFromCQ_full = 1'h0;
    cache_rqFromDmaQ_clearReq_rl = 1'h0;
    cache_rqFromDmaQ_data_0 =
	656'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
    cache_rqFromDmaQ_data_1 =
	656'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
    cache_rqFromDmaQ_deqP = 1'h0;
    cache_rqFromDmaQ_deqReq_rl = 1'h0;
    cache_rqFromDmaQ_empty = 1'h0;
    cache_rqFromDmaQ_enqP = 1'h0;
    cache_rqFromDmaQ_enqReq_rl =
	657'h0AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
    cache_rqFromDmaQ_full = 1'h0;
    cache_rsFromCQ_clearReq_rl = 1'h0;
    cache_rsFromCQ_data_0 =
	581'h0AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
    cache_rsFromCQ_data_1 =
	581'h0AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
    cache_rsFromCQ_deqP = 1'h0;
    cache_rsFromCQ_deqReq_rl = 1'h0;
    cache_rsFromCQ_empty = 1'h0;
    cache_rsFromCQ_enqP = 1'h0;
    cache_rsFromCQ_enqReq_rl =
	582'h2AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
    cache_rsFromCQ_full = 1'h0;
    cache_rsFromMQ_clearReq_rl = 1'h0;
    cache_rsFromMQ_data_0 =
	517'h0AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
    cache_rsFromMQ_data_1 =
	517'h0AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
    cache_rsFromMQ_deqP = 1'h0;
    cache_rsFromMQ_deqReq_rl = 1'h0;
    cache_rsFromMQ_empty = 1'h0;
    cache_rsFromMQ_enqP = 1'h0;
    cache_rsFromMQ_enqReq_rl =
	518'h2AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
    cache_rsFromMQ_full = 1'h0;
    cache_rsLdToDmaQ_clearReq_rl = 1'h0;
    cache_rsLdToDmaQ_data_0 =
	528'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
    cache_rsLdToDmaQ_data_1 =
	528'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
    cache_rsLdToDmaQ_deqP = 1'h0;
    cache_rsLdToDmaQ_deqReq_rl = 1'h0;
    cache_rsLdToDmaQ_empty = 1'h0;
    cache_rsLdToDmaQ_enqP = 1'h0;
    cache_rsLdToDmaQ_enqReq_rl =
	529'h0AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
    cache_rsLdToDmaQ_full = 1'h0;
    cache_rsStToDmaQ_clearReq_rl = 1'h0;
    cache_rsStToDmaQ_data_0 = 16'hAAAA;
    cache_rsStToDmaQ_data_1 = 16'hAAAA;
    cache_rsStToDmaQ_deqP = 1'h0;
    cache_rsStToDmaQ_deqReq_rl = 1'h0;
    cache_rsStToDmaQ_empty = 1'h0;
    cache_rsStToDmaQ_enqP = 1'h0;
    cache_rsStToDmaQ_enqReq_rl = 17'h0AAAA;
    cache_rsStToDmaQ_full = 1'h0;
    cache_rsToCIndexQ_clearReq_rl = 1'h0;
    cache_rsToCIndexQ_data_0 = 6'h2A;
    cache_rsToCIndexQ_data_1 = 6'h2A;
    cache_rsToCIndexQ_data_10 = 6'h2A;
    cache_rsToCIndexQ_data_11 = 6'h2A;
    cache_rsToCIndexQ_data_12 = 6'h2A;
    cache_rsToCIndexQ_data_13 = 6'h2A;
    cache_rsToCIndexQ_data_14 = 6'h2A;
    cache_rsToCIndexQ_data_15 = 6'h2A;
    cache_rsToCIndexQ_data_2 = 6'h2A;
    cache_rsToCIndexQ_data_3 = 6'h2A;
    cache_rsToCIndexQ_data_4 = 6'h2A;
    cache_rsToCIndexQ_data_5 = 6'h2A;
    cache_rsToCIndexQ_data_6 = 6'h2A;
    cache_rsToCIndexQ_data_7 = 6'h2A;
    cache_rsToCIndexQ_data_8 = 6'h2A;
    cache_rsToCIndexQ_data_9 = 6'h2A;
    cache_rsToCIndexQ_deqP = 4'hA;
    cache_rsToCIndexQ_deqReq_rl = 1'h0;
    cache_rsToCIndexQ_empty = 1'h0;
    cache_rsToCIndexQ_enqP = 4'hA;
    cache_rsToCIndexQ_enqReq_rl = 7'h2A;
    cache_rsToCIndexQ_full = 1'h0;
    cache_toCQ_clearReq_rl = 1'h0;
    cache_toCQ_data_0 =
	585'h0AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
    cache_toCQ_data_1 =
	585'h0AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
    cache_toCQ_deqP = 1'h0;
    cache_toCQ_deqReq_rl = 1'h0;
    cache_toCQ_empty = 1'h0;
    cache_toCQ_enqP = 1'h0;
    cache_toCQ_enqReq_rl =
	586'h2AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
    cache_toCQ_full = 1'h0;
    cache_toMQ_clearReq_rl = 1'h0;
    cache_toMQ_data_0 =
	641'h0AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
    cache_toMQ_data_1 =
	641'h0AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
    cache_toMQ_deqP = 1'h0;
    cache_toMQ_deqReq_rl = 1'h0;
    cache_toMQ_empty = 1'h0;
    cache_toMQ_enqP = 1'h0;
    cache_toMQ_enqReq_rl =
	642'h2AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
    cache_toMQ_full = 1'h0;
    cache_whichCRq = 4'hA;
    perfReqQ_clearReq_rl = 1'h0;
    perfReqQ_data_0 = 4'hA;
    perfReqQ_deqReq_rl = 1'h0;
    perfReqQ_empty = 1'h0;
    perfReqQ_enqReq_rl = 5'h0A;
    perfReqQ_full = 1'h0;
  end
  `endif // BSV_NO_INITIAL_BLOCKS
  // synopsys translate_on
  // handling of system tasks
  // synopsys translate_off
  always@(negedge CLK)
  begin
    #0;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_sendToM && cache_toMInfoQ$D_OUT[1:0] == 2'd0 &&
	  cache_cRqMshr$sendToM_getData[512])
	$display("Dynamic assertion failed: \"../../src_Core/Near_Mem_VM_WB_L1_L2/src_LLCache/coherence/src/LLBank.bsv\", line 560, column 38\ncannot have data");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_sendToM && cache_toMInfoQ$D_OUT[1:0] == 2'd0 &&
	  cache_cRqMshr$sendToM_getData[512])
	$finish(32'd0);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_sendToM && cache_toMInfoQ$D_OUT[1:0] == 2'd0 &&
	  cache_doLdAfterReplace)
	$display("Dynamic assertion failed: \"../../src_Core/Near_Mem_VM_WB_L1_L2/src_LLCache/coherence/src/LLBank.bsv\", line 561, column 41\ndoLdAfterReplace should be false");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_sendToM && cache_toMInfoQ$D_OUT[1:0] == 2'd0 &&
	  cache_doLdAfterReplace)
	$finish(32'd0);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_sendToM && cache_toMInfoQ$D_OUT[1:0] == 2'd1 &&
	  !cache_cRqMshr$sendToM_getRq[16])
	$display("Dynamic assertion failed: \"../../src_Core/Near_Mem_VM_WB_L1_L2/src_LLCache/coherence/src/LLBank.bsv\", line 585, column 43\nmust be dma write");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_sendToM && cache_toMInfoQ$D_OUT[1:0] == 2'd1 &&
	  !cache_cRqMshr$sendToM_getRq[16])
	$finish(32'd0);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_sendToM && cache_toMInfoQ$D_OUT[1:0] == 2'd1 &&
	  !cache_cRqMshr$sendToM_getData[512])
	$display("Dynamic assertion failed: \"../../src_Core/Near_Mem_VM_WB_L1_L2/src_LLCache/coherence/src/LLBank.bsv\", line 586, column 37\ndma write must have data");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_sendToM && cache_toMInfoQ$D_OUT[1:0] == 2'd1 &&
	  !cache_cRqMshr$sendToM_getData[512])
	$finish(32'd0);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_sendToM && cache_toMInfoQ$D_OUT[1:0] == 2'd1 &&
	  cache_doLdAfterReplace)
	$display("Dynamic assertion failed: \"../../src_Core/Near_Mem_VM_WB_L1_L2/src_LLCache/coherence/src/LLBank.bsv\", line 587, column 41\ndoLdAfterReplace should be false");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_sendToM && cache_toMInfoQ$D_OUT[1:0] == 2'd1 &&
	  cache_doLdAfterReplace)
	$finish(32'd0);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_sendToM && cache_toMInfoQ$D_OUT[1:0] == 2'd2 &&
	  cache_cRqMshr$sendToM_getRq[16])
	$display("Dynamic assertion failed: \"../../src_Core/Near_Mem_VM_WB_L1_L2/src_LLCache/coherence/src/LLBank.bsv\", line 626, column 41\nmust be child req");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_sendToM && cache_toMInfoQ$D_OUT[1:0] == 2'd2 &&
	  cache_cRqMshr$sendToM_getRq[16])
	$finish(32'd0);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_sendToM && cache_toMInfoQ$D_OUT[1:0] == 2'd2 &&
	  !cache_cRqMshr$sendToM_getData[512])
	$display("Dynamic assertion failed: \"../../src_Core/Near_Mem_VM_WB_L1_L2/src_LLCache/coherence/src/LLBank.bsv\", line 627, column 37\nreplace must have data");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_sendToM && cache_toMInfoQ$D_OUT[1:0] == 2'd2 &&
	  !cache_cRqMshr$sendToM_getData[512])
	$finish(32'd0);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_sendToM && cache_toMInfoQ$D_OUT[1:0] != 2'd0 &&
	  cache_toMInfoQ$D_OUT[1:0] != 2'd1 &&
	  cache_toMInfoQ$D_OUT[1:0] != 2'd2)
	$display("Dynamic assertion failed: \"../../src_Core/Near_Mem_VM_WB_L1_L2/src_LLCache/coherence/src/LLBank.bsv\", line 630, column 29\nunknown to mem type");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_sendToM && cache_toMInfoQ$D_OUT[1:0] != 2'd0 &&
	  cache_toMInfoQ$D_OUT[1:0] != 2'd1 &&
	  cache_toMInfoQ$D_OUT[1:0] != 2'd2)
	$finish(32'd0);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_sendRsToC &&
	  cache_cRqMshr$sendRsToDmaC_getRq[16])
	$display("Dynamic assertion failed: \"../../src_Core/Near_Mem_VM_WB_L1_L2/src_LLCache/coherence/src/LLBank.bsv\", line 697, column 37\ncRq should be child req");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_sendRsToC &&
	  cache_cRqMshr$sendRsToDmaC_getRq[16])
	$finish(32'd0);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_sendRqToC &&
	  cache_cRqMshr$sendRqToC_getState != 3'd3 &&
	  cache_cRqMshr$sendRqToC_getState != 3'd2)
	$display("Dynamic assertion failed: \"../../src_Core/Near_Mem_VM_WB_L1_L2/src_LLCache/coherence/src/LLBank.bsv\", line 761, column 13\nonly WaitSt and WaitOldTag needs req child");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_sendRqToC &&
	  cache_cRqMshr$sendRqToC_getState != 3'd3 &&
	  cache_cRqMshr$sendRqToC_getState != 3'd2)
	$finish(32'd0);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_sendRqToC &&
	  cache_cRqMshr$sendRqToC_getSlot[3:2] != 2'd1 &&
	  cache_cRqMshr$sendRqToC_getSlot[7:6] != 2'd1 &&
	  cache_cRqMshr$sendRqToC_getSlot[11:10] != 2'd1)
	$display("Dynamic assertion failed: \"../../src_Core/Near_Mem_VM_WB_L1_L2/src_LLCache/coherence/src/LLBank.bsv\", line 768, column 41\nshould have a child to downgrade");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_sendRqToC &&
	  cache_cRqMshr$sendRqToC_getSlot[3:2] != 2'd1 &&
	  cache_cRqMshr$sendRqToC_getSlot[7:6] != 2'd1 &&
	  cache_cRqMshr$sendRqToC_getSlot[11:10] != 2'd1)
	$finish(32'd0);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_sendRqToC &&
	  NOT_SEL_ARR_cache_cRqMshr_sendRqToC_getSlot_IF_ETC___d2508)
	$display("Dynamic assertion failed: \"../../src_Core/Near_Mem_VM_WB_L1_L2/src_LLCache/coherence/src/LLBank.bsv\", line 776, column 30\ndirPend should be ToSend");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_sendRqToC &&
	  NOT_SEL_ARR_cache_cRqMshr_sendRqToC_getSlot_IF_ETC___d2508)
	$finish(32'd0);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_sendRsLdToDma &&
	  !cache_cRqMshr$sendRsToDmaC_getData[512])
	$display("Dynamic assertion failed: \"../../src_Core/Near_Mem_VM_WB_L1_L2/src_LLCache/coherence/src/LLBank.bsv\", line 646, column 33\ndma read req always has valid data");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_sendRsLdToDma &&
	  !cache_cRqMshr$sendRsToDmaC_getData[512])
	$finish(32'd0);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_sendRsLdToDma &&
	  !cache_cRqMshr$sendRsToDmaC_getRq[16])
	$display("Dynamic assertion failed: \"../../src_Core/Near_Mem_VM_WB_L1_L2/src_LLCache/coherence/src/LLBank.bsv\", line 648, column 39\ncRq should be DMA req");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_sendRsLdToDma &&
	  !cache_cRqMshr$sendRsToDmaC_getRq[16])
	$finish(32'd0);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_sendRsLdToDma &&
	  (cache_cRqMshr$sendRsToDmaC_getRq[17] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[18] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[19] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[20] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[21] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[22] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[23] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[24] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[25] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[26] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[27] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[28] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[29] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[30] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[31] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[32] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[33] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[34] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[35] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[36] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[37] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[38] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[39] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[40] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[41] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[42] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[43] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[44] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[45] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[46] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[47] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[48] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[49] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[50] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[51] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[52] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[53] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[54] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[55] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[56] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[57] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[58] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[59] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[60] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[61] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[62] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[63] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[64] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[65] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[66] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[67] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[68] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[69] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[70] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[71] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[72] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[73] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[74] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[75] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[76] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[77] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[78] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[79] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[80] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[85:84] != 2'd1))
	$display("Dynamic assertion failed: \"../../src_Core/Near_Mem_VM_WB_L1_L2/src_LLCache/coherence/src/LLBank.bsv\", line 650, column 13\ncRq should be DMA read");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_sendRsLdToDma &&
	  (cache_cRqMshr$sendRsToDmaC_getRq[17] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[18] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[19] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[20] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[21] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[22] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[23] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[24] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[25] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[26] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[27] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[28] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[29] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[30] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[31] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[32] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[33] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[34] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[35] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[36] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[37] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[38] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[39] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[40] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[41] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[42] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[43] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[44] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[45] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[46] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[47] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[48] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[49] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[50] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[51] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[52] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[53] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[54] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[55] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[56] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[57] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[58] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[59] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[60] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[61] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[62] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[63] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[64] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[65] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[66] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[67] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[68] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[69] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[70] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[71] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[72] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[73] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[74] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[75] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[76] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[77] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[78] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[79] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[80] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[85:84] != 2'd1))
	$finish(32'd0);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_sendRsStToDma &&
	  !cache_cRqMshr$sendRsToDmaC_getRq[16])
	$display("Dynamic assertion failed: \"../../src_Core/Near_Mem_VM_WB_L1_L2/src_LLCache/coherence/src/LLBank.bsv\", line 671, column 39\ncRq should be DMA req");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_sendRsStToDma &&
	  !cache_cRqMshr$sendRsToDmaC_getRq[16])
	$finish(32'd0);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_sendRsStToDma &&
	  (!cache_cRqMshr$sendRsToDmaC_getRq[17] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[18] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[19] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[20] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[21] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[22] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[23] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[24] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[25] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[26] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[27] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[28] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[29] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[30] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[31] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[32] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[33] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[34] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[35] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[36] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[37] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[38] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[39] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[40] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[41] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[42] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[43] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[44] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[45] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[46] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[47] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[48] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[49] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[50] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[51] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[52] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[53] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[54] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[55] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[56] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[57] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[58] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[59] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[60] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[61] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[62] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[63] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[64] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[65] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[66] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[67] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[68] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[69] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[70] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[71] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[72] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[73] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[74] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[75] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[76] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[77] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[78] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[79] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[80] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[85:84] != 2'd3))
	$display("Dynamic assertion failed: \"../../src_Core/Near_Mem_VM_WB_L1_L2/src_LLCache/coherence/src/LLBank.bsv\", line 673, column 13\ncRq should be DMA write");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_sendRsStToDma &&
	  (!cache_cRqMshr$sendRsToDmaC_getRq[17] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[18] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[19] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[20] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[21] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[22] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[23] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[24] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[25] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[26] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[27] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[28] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[29] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[30] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[31] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[32] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[33] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[34] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[35] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[36] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[37] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[38] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[39] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[40] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[41] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[42] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[43] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[44] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[45] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[46] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[47] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[48] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[49] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[50] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[51] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[52] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[53] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[54] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[55] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[56] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[57] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[58] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[59] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[60] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[61] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[62] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[63] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[64] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[65] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[66] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[67] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[68] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[69] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[70] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[71] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[72] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[73] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[74] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[75] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[76] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[77] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[78] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[79] &&
	   !cache_cRqMshr$sendRsToDmaC_getRq[80] ||
	   cache_cRqMshr$sendRsToDmaC_getRq[85:84] != 2'd3))
	$finish(32'd0);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_cRq && cache_pipeline$first[517] &&
	  cache_pipeline_first__581_BITS_516_TO_513_583__ETC___d2588 &&
	  cache_cRqMshr$pipelineResp_getState != 3'd5)
	$display("Dynamic assertion failed: \"../../src_Core/Near_Mem_VM_WB_L1_L2/src_LLCache/coherence/src/LLBank.bsv\", line 1191, column 44\nowner is myself, must be swapped in");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_cRq && cache_pipeline$first[517] &&
	  cache_pipeline_first__581_BITS_516_TO_513_583__ETC___d2588 &&
	  cache_cRqMshr$pipelineResp_getState != 3'd5)
	$finish(32'd0);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_cRq && cache_pipeline$first[517] &&
	  cache_pipeline_first__581_BITS_516_TO_513_583__ETC___d2588 &&
	  (!cache_pipeline_first__581_BITS_573_TO_526_644__ETC___d2646 ||
	   cache_pipeline$first[525:524] == 2'd0))
	$display("Dynamic assertion failed: \"../../src_Core/Near_Mem_VM_WB_L1_L2/src_LLCache/coherence/src/LLBank.bsv\", line 1195, column 21\ncRq swapped in, tag must match, cs > I");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_cRq && cache_pipeline$first[517] &&
	  cache_pipeline_first__581_BITS_516_TO_513_583__ETC___d2588 &&
	  (!cache_pipeline_first__581_BITS_573_TO_526_644__ETC___d2646 ||
	   cache_pipeline$first[525:524] == 2'd0))
	$finish(32'd0);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_cRq &&
	  cache_pipeline_first__581_BIT_517_582_AND_cach_ETC___d3195)
	$display("Dynamic assertion failed: \"../../src_Core/Near_Mem_VM_WB_L1_L2/src_LLCache/coherence/src/LLBank.bsv\", line 893, column 38\nmust match pipe out cRq idx");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_cRq &&
	  cache_pipeline_first__581_BIT_517_582_AND_cach_ETC___d3195)
	$finish(32'd0);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_cRq &&
	  cache_pipeline_first__581_BIT_517_582_AND_cach_ETC___d3199)
	$display("Dynamic assertion failed: \"../../src_Core/Near_Mem_VM_WB_L1_L2/src_LLCache/coherence/src/LLBank.bsv\", line 896, column 13\ncRqHit but tag or cs incorrect");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_cRq &&
	  cache_pipeline_first__581_BIT_517_582_AND_cach_ETC___d3199)
	$finish(32'd0);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_cRq &&
	  cache_pipeline_first__581_BIT_517_582_AND_cach_ETC___d3268)
	$display("Dynamic assertion failed: \"../../src_Core/Near_Mem_VM_WB_L1_L2/src_LLCache/coherence/src/LLBank.bsv\", line 898, column 74\ntoState should match byteEn");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_cRq &&
	  cache_pipeline_first__581_BIT_517_582_AND_cach_ETC___d3268)
	$finish(32'd0);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_cRq &&
	  cache_pipeline_first__581_BIT_517_582_AND_cach_ETC___d3274)
	$display("Dynamic assertion failed: \"../../src_Core/Near_Mem_VM_WB_L1_L2/src_LLCache/coherence/src/LLBank.bsv\", line 907, column 13\ndma write should carry valid data");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_cRq &&
	  cache_pipeline_first__581_BIT_517_582_AND_cach_ETC___d3274)
	$finish(32'd0);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_cRq &&
	  cache_pipeline_first__581_BIT_517_582_AND_cach_ETC___d3278)
	$display("Dynamic assertion failed: \"../../src_Core/Near_Mem_VM_WB_L1_L2/src_LLCache/coherence/src/LLBank.bsv\", line 1082, column 17\ntag match and cs > I");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_cRq &&
	  cache_pipeline_first__581_BIT_517_582_AND_cach_ETC___d3278)
	$finish(32'd0);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_cRq &&
	  cache_pipeline_first__581_BIT_517_582_AND_cach_ETC___d3284)
	$display("Dynamic assertion failed: \"../../src_Core/Near_Mem_VM_WB_L1_L2/src_LLCache/coherence/src/LLBank.bsv\", line 1087, column 36\nwaitP must be false");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_cRq &&
	  cache_pipeline_first__581_BIT_517_582_AND_cach_ETC___d3284)
	$finish(32'd0);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_cRq && cache_pipeline$first[517] &&
	  cache_pipeline_first__581_BITS_516_TO_513_583__ETC___d3287)
	$display("Dynamic assertion failed: \"../../src_Core/Near_Mem_VM_WB_L1_L2/src_LLCache/coherence/src/LLBank.bsv\", line 835, column 38\nmust match pipe out cRq idx");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_cRq && cache_pipeline$first[517] &&
	  cache_pipeline_first__581_BITS_516_TO_513_583__ETC___d3287)
	$finish(32'd0);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_cRq && cache_pipeline$first[517] &&
	  cache_pipeline_first__581_BITS_516_TO_513_583__ETC___d2588 &&
	  NOT_cache_cRqMshr_pipelineResp_getRq_IF_cache__ETC___d3290)
	$display("Dynamic assertion failed: \"../../src_Core/Near_Mem_VM_WB_L1_L2/src_LLCache/coherence/src/LLBank.bsv\", line 841, column 14\ncRqHit but tag or cs incorrect");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_cRq && cache_pipeline$first[517] &&
	  cache_pipeline_first__581_BITS_516_TO_513_583__ETC___d2588 &&
	  NOT_cache_cRqMshr_pipelineResp_getRq_IF_cache__ETC___d3290)
	$finish(32'd0);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_cRq && cache_pipeline$first[517] &&
	  cache_pipeline_first__581_BITS_516_TO_513_583__ETC___d3295)
	$display("Dynamic assertion failed: \"../../src_Core/Near_Mem_VM_WB_L1_L2/src_LLCache/coherence/src/LLBank.bsv\", line 1047, column 36\nwaitP must be false");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_cRq && cache_pipeline$first[517] &&
	  cache_pipeline_first__581_BITS_516_TO_513_583__ETC___d3295)
	$finish(32'd0);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_cRq && cache_pipeline$first[517] &&
	  cache_pipeline_first__581_BITS_516_TO_513_583__ETC___d2588 &&
	  NOT_cache_cRqMshr_pipelineResp_getRq_IF_cache__ETC___d3299)
	$display("Dynamic assertion failed: \"../../src_Core/Near_Mem_VM_WB_L1_L2/src_LLCache/coherence/src/LLBank.bsv\", line 1054, column 56\ndir should be all I");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_cRq && cache_pipeline$first[517] &&
	  cache_pipeline_first__581_BITS_516_TO_513_583__ETC___d2588 &&
	  NOT_cache_cRqMshr_pipelineResp_getRq_IF_cache__ETC___d3299)
	$finish(32'd0);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_cRq && cache_pipeline$first[517] &&
	  !cache_pipeline_first__581_BITS_516_TO_513_583__ETC___d2588 &&
	  cache_cRqMshr$pipelineResp_getState != 3'd1)
	$display("Dynamic assertion failed: \"../../src_Core/Near_Mem_VM_WB_L1_L2/src_LLCache/coherence/src/LLBank.bsv\", line 1157, column 42\nowner is other, must first time go through tag match");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_cRq && cache_pipeline$first[517] &&
	  !cache_pipeline_first__581_BITS_516_TO_513_583__ETC___d2588 &&
	  cache_cRqMshr$pipelineResp_getState != 3'd1)
	$finish(32'd0);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_cRq && cache_pipeline$first[517] &&
	  !cache_pipeline_first__581_BITS_516_TO_513_583__ETC___d2588 &&
	  (cache_pipeline$first[525:524] == 2'd0 ||
	   !cache_pipeline_first__581_BITS_573_TO_526_644__ETC___d2646))
	$display("Dynamic assertion failed: \"../../src_Core/Near_Mem_VM_WB_L1_L2/src_LLCache/coherence/src/LLBank.bsv\", line 1160, column 22\ncRq should hit in tag match");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_cRq && cache_pipeline$first[517] &&
	  !cache_pipeline_first__581_BITS_516_TO_513_583__ETC___d2588 &&
	  (cache_pipeline$first[525:524] == 2'd0 ||
	   !cache_pipeline_first__581_BITS_573_TO_526_644__ETC___d2646))
	$finish(32'd0);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_cRq && cache_pipeline$first[517] &&
	  !cache_pipeline_first__581_BITS_516_TO_513_583__ETC___d2588 &&
	  !cache_cRqMshr$pipelineResp_searchEndOfChain[4] &&
	  !cache_pipeline$first[512])
	$display("Dynamic assertion failed: \"../../src_Core/Near_Mem_VM_WB_L1_L2/src_LLCache/coherence/src/LLBank.bsv\", line 1185, column 48\nline must be replacing");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_cRq && cache_pipeline$first[517] &&
	  !cache_pipeline_first__581_BITS_516_TO_513_583__ETC___d2588 &&
	  !cache_cRqMshr$pipelineResp_searchEndOfChain[4] &&
	  !cache_pipeline$first[512])
	$finish(32'd0);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_cRq &&
	  NOT_cache_pipeline_first__581_BIT_517_582_105__ETC___d3316)
	$display("Dynamic assertion failed: \"../../src_Core/Near_Mem_VM_WB_L1_L2/src_LLCache/coherence/src/LLBank.bsv\", line 893, column 38\nmust match pipe out cRq idx");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_cRq &&
	  NOT_cache_pipeline_first__581_BIT_517_582_105__ETC___d3316)
	$finish(32'd0);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_cRq &&
	  NOT_cache_pipeline_first__581_BIT_517_582_105__ETC___d3320)
	$display("Dynamic assertion failed: \"../../src_Core/Near_Mem_VM_WB_L1_L2/src_LLCache/coherence/src/LLBank.bsv\", line 898, column 74\ntoState should match byteEn");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_cRq &&
	  NOT_cache_pipeline_first__581_BIT_517_582_105__ETC___d3320)
	$finish(32'd0);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_cRq &&
	  NOT_cache_pipeline_first__581_BIT_517_582_105__ETC___d3324)
	$display("Dynamic assertion failed: \"../../src_Core/Near_Mem_VM_WB_L1_L2/src_LLCache/coherence/src/LLBank.bsv\", line 907, column 13\ndma write should carry valid data");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_cRq &&
	  NOT_cache_pipeline_first__581_BIT_517_582_105__ETC___d3324)
	$finish(32'd0);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_cRq &&
	  NOT_cache_pipeline_first__581_BIT_517_582_105__ETC___d3328)
	$display("Dynamic assertion failed: \"../../src_Core/Near_Mem_VM_WB_L1_L2/src_LLCache/coherence/src/LLBank.bsv\", line 1087, column 36\nwaitP must be false");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_cRq &&
	  NOT_cache_pipeline_first__581_BIT_517_582_105__ETC___d3328)
	$finish(32'd0);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_cRq &&
	  NOT_cache_pipeline_first__581_BIT_517_582_105__ETC___d3340)
	$display("Dynamic assertion failed: \"../../src_Core/Near_Mem_VM_WB_L1_L2/src_LLCache/coherence/src/LLBank.bsv\", line 1308, column 53\nshould not have any rep succ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_cRq &&
	  NOT_cache_pipeline_first__581_BIT_517_582_105__ETC___d3340)
	$finish(32'd0);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_cRq &&
	  NOT_cache_pipeline_first__581_BIT_517_582_105__ETC___d3345)
	$display("Dynamic assertion failed: \"../../src_Core/Near_Mem_VM_WB_L1_L2/src_LLCache/coherence/src/LLBank.bsv\", line 835, column 38\nmust match pipe out cRq idx");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_cRq &&
	  NOT_cache_pipeline_first__581_BIT_517_582_105__ETC___d3345)
	$finish(32'd0);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_cRq &&
	  NOT_cache_pipeline_first__581_BIT_517_582_105__ETC___d3351)
	$display("Dynamic assertion failed: \"../../src_Core/Near_Mem_VM_WB_L1_L2/src_LLCache/coherence/src/LLBank.bsv\", line 1047, column 36\nwaitP must be false");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_cRq &&
	  NOT_cache_pipeline_first__581_BIT_517_582_105__ETC___d3351)
	$finish(32'd0);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_cRq && !cache_pipeline$first[517] &&
	  NOT_cache_cRqMshr_pipelineResp_searchEndOfChai_ETC___d3353)
	$display("Dynamic assertion failed: \"../../src_Core/Near_Mem_VM_WB_L1_L2/src_LLCache/coherence/src/LLBank.bsv\", line 1054, column 56\ndir should be all I");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_cRq && !cache_pipeline$first[517] &&
	  NOT_cache_cRqMshr_pipelineResp_searchEndOfChai_ETC___d3353)
	$finish(32'd0);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_cRq &&
	  NOT_cache_pipeline_first__581_BIT_517_582_105__ETC___d3359)
	$display("Dynamic assertion failed: \"../../src_Core/Near_Mem_VM_WB_L1_L2/src_LLCache/coherence/src/LLBank.bsv\", line 1117, column 45\ncannot have rep succ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_cRq &&
	  NOT_cache_pipeline_first__581_BIT_517_582_105__ETC___d3359)
	$finish(32'd0);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_mRs && !cache_pipeline$first[517])
	$display("Dynamic assertion failed: \"../../src_Core/Near_Mem_VM_WB_L1_L2/src_LLCache/coherence/src/LLBank.bsv\", line 1318, column 43\nmRs owner must match some cRq");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_mRs && !cache_pipeline$first[517])
	$finish(32'd0);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_mRs &&
	  cache_cRqMshr$pipelineResp_getRq[16])
	$display("Dynamic assertion failed: \"../../src_Core/Near_Mem_VM_WB_L1_L2/src_LLCache/coherence/src/LLBank.bsv\", line 1329, column 37\nonly child req gets mem resp that refills the cache");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_mRs &&
	  cache_cRqMshr$pipelineResp_getRq[16])
	$finish(32'd0);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_mRs &&
	  (cache_pipeline$first[525:524] <
	   cache_cRqMshr$pipelineResp_getRq[85:84] ||
	   !cache_pipeline_first__581_BITS_573_TO_526_644__ETC___d2646))
	$display("Dynamic assertion failed: \"../../src_Core/Near_Mem_VM_WB_L1_L2/src_LLCache/coherence/src/LLBank.bsv\", line 1331, column 13\nmRs must be tag match & have enough cs");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_mRs &&
	  (cache_pipeline$first[525:524] <
	   cache_cRqMshr$pipelineResp_getRq[85:84] ||
	   !cache_pipeline_first__581_BITS_573_TO_526_644__ETC___d2646))
	$finish(32'd0);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_mRs &&
	  (cache_pipeline$first[519:518] != 2'd0 ||
	   cache_pipeline$first[521:520] != 2'd0 ||
	   cache_pipeline$first[523:522] != 2'd0))
	$display("Dynamic assertion failed: \"../../src_Core/Near_Mem_VM_WB_L1_L2/src_LLCache/coherence/src/LLBank.bsv\", line 1333, column 48\nall children must be I");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_mRs &&
	  (cache_pipeline$first[519:518] != 2'd0 ||
	   cache_pipeline$first[521:520] != 2'd0 ||
	   cache_pipeline$first[523:522] != 2'd0))
	$finish(32'd0);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_mRs && cache_pipeline$first[512])
	$display("Dynamic assertion failed: \"../../src_Core/Near_Mem_VM_WB_L1_L2/src_LLCache/coherence/src/LLBank.bsv\", line 1334, column 37\nmRs cannot hit on replacing line");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_mRs && cache_pipeline$first[512])
	$finish(32'd0);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_mRs &&
	  NOT_cache_cRqMshr_pipelineResp_getSlot_IF_cach_ETC___d3369)
	$display("Dynamic assertion failed: \"../../src_Core/Near_Mem_VM_WB_L1_L2/src_LLCache/coherence/src/LLBank.bsv\", line 1335, column 44\nmRs should hit on way in MSHR slot");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_mRs &&
	  NOT_cache_cRqMshr_pipelineResp_getSlot_IF_cach_ETC___d3369)
	$finish(32'd0);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_mRs &&
	  !cache_cRqMshr$pipelineResp_getSlot[12])
	$display("Dynamic assertion failed: \"../../src_Core/Near_Mem_VM_WB_L1_L2/src_LLCache/coherence/src/LLBank.bsv\", line 1336, column 31\nmRs should match cRq which is waiting for it");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_mRs &&
	  !cache_cRqMshr$pipelineResp_getSlot[12])
	$finish(32'd0);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_mRs &&
	  (cache_cRqMshr$pipelineResp_getSlot[3:2] != 2'd0 ||
	   cache_cRqMshr$pipelineResp_getSlot[7:6] != 2'd0 ||
	   cache_cRqMshr$pipelineResp_getSlot[11:10] != 2'd0))
	$display("Dynamic assertion failed: \"../../src_Core/Near_Mem_VM_WB_L1_L2/src_LLCache/coherence/src/LLBank.bsv\", line 1338, column 13\ncRq that needs mRs should not have children to wait for");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_mRs &&
	  (cache_cRqMshr$pipelineResp_getSlot[3:2] != 2'd0 ||
	   cache_cRqMshr$pipelineResp_getSlot[7:6] != 2'd0 ||
	   cache_cRqMshr$pipelineResp_getSlot[11:10] != 2'd0))
	$finish(32'd0);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_mRs &&
	  NOT_cache_pipeline_first__581_BITS_516_TO_513__ETC___d3798)
	$display("Dynamic assertion failed: \"../../src_Core/Near_Mem_VM_WB_L1_L2/src_LLCache/coherence/src/LLBank.bsv\", line 835, column 38\nmust match pipe out cRq idx");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_mRs &&
	  NOT_cache_pipeline_first__581_BITS_516_TO_513__ETC___d3798)
	$finish(32'd0);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_mRs &&
	  cache_cRqMshr$pipelineResp_getRq[16])
	$display("Dynamic assertion failed: \"../../src_Core/Near_Mem_VM_WB_L1_L2/src_LLCache/coherence/src/LLBank.bsv\", line 836, column 37\nshould be cRq from child");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_mRs &&
	  cache_cRqMshr$pipelineResp_getRq[16])
	$finish(32'd0);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_mRs &&
	  (!cache_pipeline_first__581_BITS_573_TO_526_644__ETC___d2646 ||
	   cache_pipeline$first[525:524] == 2'd0))
	$display("Dynamic assertion failed: \"../../src_Core/Near_Mem_VM_WB_L1_L2/src_LLCache/coherence/src/LLBank.bsv\", line 841, column 14\ncRqHit but tag or cs incorrect");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_mRs &&
	  (!cache_pipeline_first__581_BITS_573_TO_526_644__ETC___d2646 ||
	   cache_pipeline$first[525:524] == 2'd0))
	$finish(32'd0);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_cRs &&
	  cache_pipeline$first[525:524] == 2'd0)
	$display("Dynamic assertion failed: \"../../src_Core/Near_Mem_VM_WB_L1_L2/src_LLCache/coherence/src/LLBank.bsv\", line 1352, column 35\ncRs should hit on a line");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_cRs &&
	  cache_pipeline$first[525:524] == 2'd0)
	$finish(32'd0);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_cRs && cache_pipeline$first[517] &&
	  NOT_cache_cRqMshr_pipelineResp_getSlot_IF_cach_ETC___d3369)
	$display("Dynamic assertion failed: \"../../src_Core/Near_Mem_VM_WB_L1_L2/src_LLCache/coherence/src/LLBank.bsv\", line 1365, column 48\ncRs way should match MSHR slot");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_cRs && cache_pipeline$first[517] &&
	  NOT_cache_cRqMshr_pipelineResp_getSlot_IF_cach_ETC___d3369)
	$finish(32'd0);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_cRs && cache_pipeline$first[517] &&
	  cache_pipeline$first[512] &&
	  cache_cRqMshr$pipelineResp_getRq[16])
	$display("Dynamic assertion failed: \"../../src_Core/Near_Mem_VM_WB_L1_L2/src_LLCache/coherence/src/LLBank.bsv\", line 1369, column 45\nonly child req do replace");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_cRs && cache_pipeline$first[517] &&
	  cache_pipeline$first[512] &&
	  cache_cRqMshr$pipelineResp_getRq[16])
	$finish(32'd0);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_cRs && cache_pipeline$first[517] &&
	  cache_pipeline$first[512] &&
	  cache_cRqMshr$pipelineResp_getState != 3'd2)
	$display("Dynamic assertion failed: \"../../src_Core/Near_Mem_VM_WB_L1_L2/src_LLCache/coherence/src/LLBank.bsv\", line 1370, column 48\nmust be waiting for old tag");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_cRs && cache_pipeline$first[517] &&
	  cache_pipeline$first[512] &&
	  cache_cRqMshr$pipelineResp_getState != 3'd2)
	$finish(32'd0);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_cRs && cache_pipeline$first[517] &&
	  cache_pipeline$first[512] &&
	  cache_cRqMshr$pipelineResp_getSlot[12])
	$display("Dynamic assertion failed: \"../../src_Core/Near_Mem_VM_WB_L1_L2/src_LLCache/coherence/src/LLBank.bsv\", line 1371, column 40\ncannot wait for parent while replacing");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_cRs && cache_pipeline$first[517] &&
	  cache_pipeline$first[512] &&
	  cache_cRqMshr$pipelineResp_getSlot[12])
	$finish(32'd0);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_cRs && cache_pipeline$first[517] &&
	  cache_pipeline$first[512] &&
	  cache_cRqMshr$pipelineResp_getSlot[60:13] !=
	  cache_pipeline$first[573:526])
	$display("Dynamic assertion failed: \"../../src_Core/Near_Mem_VM_WB_L1_L2/src_LLCache/coherence/src/LLBank.bsv\", line 1372, column 56\nshould match replacing tag");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_cRs && cache_pipeline$first[517] &&
	  cache_pipeline$first[512] &&
	  cache_cRqMshr$pipelineResp_getSlot[60:13] !=
	  cache_pipeline$first[573:526])
	$finish(32'd0);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_cRs && cache_pipeline$first[517] &&
	  cache_pipeline$first[512] &&
	  IF_SEL_ARR_cache_pipeline_first__581_BITS_519__ETC___d3488 &&
	  cache_cRqMshr$pipelineResp_getRq[16])
	$display("Dynamic assertion failed: \"../../src_Core/Near_Mem_VM_WB_L1_L2/src_LLCache/coherence/src/LLBank.bsv\", line 953, column 37\nonly cRq from child can evict a line");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_cRs && cache_pipeline$first[517] &&
	  cache_pipeline$first[512] &&
	  IF_SEL_ARR_cache_pipeline_first__581_BITS_519__ETC___d3488 &&
	  cache_cRqMshr$pipelineResp_getRq[16])
	$finish(32'd0);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_cRs && cache_pipeline$first[517] &&
	  cache_pipeline$first[512] &&
	  IF_SEL_ARR_cache_pipeline_first__581_BITS_519__ETC___d3488 &&
	  (cache_pipeline$first[519:518] != 2'd0 ||
	   cache_pipeline$first[521:520] != 2'd0 ||
	   cache_pipeline$first[523:522] != 2'd0 ||
	   cache_pipeline$first[525:524] == 2'd0))
	$display("Dynamic assertion failed: \"../../src_Core/Near_Mem_VM_WB_L1_L2/src_LLCache/coherence/src/LLBank.bsv\", line 955, column 13\nonly evict valid line which has no children");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_cRs && cache_pipeline$first[517] &&
	  cache_pipeline$first[512] &&
	  IF_SEL_ARR_cache_pipeline_first__581_BITS_519__ETC___d3488 &&
	  (cache_pipeline$first[519:518] != 2'd0 ||
	   cache_pipeline$first[521:520] != 2'd0 ||
	   cache_pipeline$first[523:522] != 2'd0 ||
	   cache_pipeline$first[525:524] == 2'd0))
	$finish(32'd0);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_cRs && cache_pipeline$first[517] &&
	  !cache_pipeline$first[512] &&
	  cache_cRqMshr$pipelineResp_getState != 3'd3)
	$display("Dynamic assertion failed: \"../../src_Core/Near_Mem_VM_WB_L1_L2/src_LLCache/coherence/src/LLBank.bsv\", line 1405, column 44\nmust be waiting for child/parent state");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_cRs && cache_pipeline$first[517] &&
	  !cache_pipeline$first[512] &&
	  cache_cRqMshr$pipelineResp_getState != 3'd3)
	$finish(32'd0);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_cRs && cache_pipeline$first[517] &&
	  !cache_pipeline$first[512] &&
	  !cache_pipeline_first__581_BITS_573_TO_526_644__ETC___d2646)
	$display("Dynamic assertion failed: \"../../src_Core/Near_Mem_VM_WB_L1_L2/src_LLCache/coherence/src/LLBank.bsv\", line 1406, column 60\ncRq tag should match cRs hit line");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_cRs && cache_pipeline$first[517] &&
	  !cache_pipeline$first[512] &&
	  !cache_pipeline_first__581_BITS_573_TO_526_644__ETC___d2646)
	$finish(32'd0);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_cRs && cache_pipeline$first[517] &&
	  !cache_pipeline$first[512] &&
	  cache_cRqMshr$pipelineResp_getSlot[12])
	$display("Dynamic assertion failed: \"../../src_Core/Near_Mem_VM_WB_L1_L2/src_LLCache/coherence/src/LLBank.bsv\", line 1407, column 40\ncs > I, so cannot wait for memory");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_cRs && cache_pipeline$first[517] &&
	  !cache_pipeline$first[512] &&
	  cache_cRqMshr$pipelineResp_getSlot[12])
	$finish(32'd0);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_cRs && cache_pipeline$first[517] &&
	  NOT_cache_pipeline_first__581_BIT_512_308_309__ETC___d3801)
	$display("Dynamic assertion failed: \"../../src_Core/Near_Mem_VM_WB_L1_L2/src_LLCache/coherence/src/LLBank.bsv\", line 893, column 38\nmust match pipe out cRq idx");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_cRs && cache_pipeline$first[517] &&
	  NOT_cache_pipeline_first__581_BIT_512_308_309__ETC___d3801)
	$finish(32'd0);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_cRs && cache_pipeline$first[517] &&
	  !cache_pipeline$first[512] &&
	  IF_SEL_ARR_cache_cRqMshr_pipelineResp_getSlot__ETC___d3804)
	$display("Dynamic assertion failed: \"../../src_Core/Near_Mem_VM_WB_L1_L2/src_LLCache/coherence/src/LLBank.bsv\", line 896, column 13\ncRqHit but tag or cs incorrect");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_cRs && cache_pipeline$first[517] &&
	  !cache_pipeline$first[512] &&
	  IF_SEL_ARR_cache_cRqMshr_pipelineResp_getSlot__ETC___d3804)
	$finish(32'd0);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_cRs && cache_pipeline$first[517] &&
	  NOT_cache_pipeline_first__581_BIT_512_308_309__ETC___d3809)
	$display("Dynamic assertion failed: \"../../src_Core/Near_Mem_VM_WB_L1_L2/src_LLCache/coherence/src/LLBank.bsv\", line 898, column 74\ntoState should match byteEn");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_cRs && cache_pipeline$first[517] &&
	  NOT_cache_pipeline_first__581_BIT_512_308_309__ETC___d3809)
	$finish(32'd0);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_cRs && cache_pipeline$first[517] &&
	  !cache_pipeline$first[512] &&
	  IF_SEL_ARR_cache_cRqMshr_pipelineResp_getSlot__ETC___d3814)
	$display("Dynamic assertion failed: \"../../src_Core/Near_Mem_VM_WB_L1_L2/src_LLCache/coherence/src/LLBank.bsv\", line 907, column 13\ndma write should carry valid data");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_cRs && cache_pipeline$first[517] &&
	  !cache_pipeline$first[512] &&
	  IF_SEL_ARR_cache_cRqMshr_pipelineResp_getSlot__ETC___d3814)
	$finish(32'd0);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_cRs && cache_pipeline$first[517] &&
	  NOT_cache_pipeline_first__581_BIT_512_308_309__ETC___d3827)
	$display("Dynamic assertion failed: \"../../src_Core/Near_Mem_VM_WB_L1_L2/src_LLCache/coherence/src/LLBank.bsv\", line 835, column 38\nmust match pipe out cRq idx");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_cRs && cache_pipeline$first[517] &&
	  NOT_cache_pipeline_first__581_BIT_512_308_309__ETC___d3827)
	$finish(32'd0);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_cRs && cache_pipeline$first[517] &&
	  !cache_pipeline$first[512] &&
	  IF_SEL_ARR_cache_cRqMshr_pipelineResp_getSlot__ETC___d3830)
	$display("Dynamic assertion failed: \"../../src_Core/Near_Mem_VM_WB_L1_L2/src_LLCache/coherence/src/LLBank.bsv\", line 841, column 14\ncRqHit but tag or cs incorrect");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_pipelineResp_cRs && cache_pipeline$first[517] &&
	  !cache_pipeline$first[512] &&
	  IF_SEL_ARR_cache_cRqMshr_pipelineResp_getSlot__ETC___d3830)
	$finish(32'd0);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_mRsTransfer && cache_cRqMshr$transfer_getRq[16])
	$display("Dynamic assertion failed: \"../../src_Core/Near_Mem_VM_WB_L1_L2/src_LLCache/coherence/src/LLBank.bsv\", line 491, column 37\nrefill mem resp must be for child req");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_cache_mRsTransfer && cache_cRqMshr$transfer_getRq[16])
	$finish(32'd0);
  end
  // synopsys translate_on
endmodule