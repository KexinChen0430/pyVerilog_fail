module header
	// Internal signals
	// Generated Signal List
	// End of Generated Signal List
	// %COMPILER_OPTS%
	// Generated Signal Assignments
	// Generated Instances and Port Mappings
		// Generated Instance Port Map for inst_1
		inst_1_e inst_1 (
		);
		defparam inst_1.FOO = 16;
		// End of Generated Instance Port Map for inst_1
		// Generated Instance Port Map for inst_10
		inst_10_e inst_10 (
		);
		defparam inst_10.FOO = 32;
		// End of Generated Instance Port Map for inst_10
		// Generated Instance Port Map for inst_2
		inst_2_e inst_2 (
		);
		defparam inst_2.FOO = 16;
		// End of Generated Instance Port Map for inst_2
		// Generated Instance Port Map for inst_3
		inst_3_e inst_3 (
		);
		defparam inst_3.FOO = 16;
		// End of Generated Instance Port Map for inst_3
		// Generated Instance Port Map for inst_4
		inst_4_e inst_4 (
		);
		defparam inst_4.FOO = 16;
		// End of Generated Instance Port Map for inst_4
		// Generated Instance Port Map for inst_5
		inst_5_e inst_5 (
		);
		// End of Generated Instance Port Map for inst_5
		// Generated Instance Port Map for inst_6
		inst_6_e inst_6 (
		);
		// End of Generated Instance Port Map for inst_6
		// Generated Instance Port Map for inst_7
		inst_7_e inst_7 (
		);
		defparam inst_7.FOO = 32;
		// End of Generated Instance Port Map for inst_7
		// Generated Instance Port Map for inst_8
		inst_8_e inst_8 (
		);
		defparam inst_8.FOO = 32;
		// End of Generated Instance Port Map for inst_8
		// Generated Instance Port Map for inst_9
		inst_9_e inst_9 (
		);
		defparam inst_9.FOO = 32;
		// End of Generated Instance Port Map for inst_9
		// Generated Instance Port Map for inst_aa
		inst_aa_e inst_aa (
		);
		defparam inst_aa.NO_DEFAULT = "nodefault",
			inst_aa.NO_NAME = "noname",
			inst_aa.WIDTH = 15;
		// End of Generated Instance Port Map for inst_aa
		// Generated Instance Port Map for inst_ab
		inst_ab_e inst_ab (
		);
		defparam inst_ab.WIDTH = 31;
		// End of Generated Instance Port Map for inst_ab
		// Generated Instance Port Map for inst_ac
		inst_ac_e inst_ac (
		);
		// End of Generated Instance Port Map for inst_ac
		// Generated Instance Port Map for inst_ad
		inst_ad_e inst_ad (
		);
		// End of Generated Instance Port Map for inst_ad
		// Generated Instance Port Map for inst_ae
		inst_ae_e inst_ae (
		);
		// End of Generated Instance Port Map for inst_ae
		// Generated Instance Port Map for inst_m1
		inst_m_e inst_m1 (
		);
		defparam inst_m1.FOO = 15;
		// End of Generated Instance Port Map for inst_m1
		// Generated Instance Port Map for inst_m10
		inst_m_e inst_m10 (
		);
		defparam inst_m10.FOO = 30;
		// End of Generated Instance Port Map for inst_m10
		// Generated Instance Port Map for inst_m2
		inst_m_e inst_m2 (
		);
		defparam inst_m2.FOO = 15;
		// End of Generated Instance Port Map for inst_m2
		// Generated Instance Port Map for inst_m3
		inst_m_e inst_m3 (
		);
		defparam inst_m3.FOO = 15;
		// End of Generated Instance Port Map for inst_m3
		// Generated Instance Port Map for inst_m4
		inst_m_e inst_m4 (
		);
		defparam inst_m4.FOO = 15;
		// End of Generated Instance Port Map for inst_m4
		// Generated Instance Port Map for inst_m5
		inst_m_e inst_m5 (
		);
		defparam inst_m5.FOO = 15;
		// End of Generated Instance Port Map for inst_m5
		// Generated Instance Port Map for inst_m6
		inst_m_e inst_m6 (
		);
		defparam inst_m6.FOO = 30;
		// End of Generated Instance Port Map for inst_m6
		// Generated Instance Port Map for inst_m7
		inst_m_e inst_m7 (
		);
		defparam inst_m7.FOO = 30;
		// End of Generated Instance Port Map for inst_m7
		// Generated Instance Port Map for inst_m8
		inst_m_e inst_m8 (
		);
		defparam inst_m8.FOO = 30;
		// End of Generated Instance Port Map for inst_m8
		// Generated Instance Port Map for inst_m9
		inst_m_e inst_m9 (
		);
		defparam inst_m9.FOO = 30;
		// End of Generated Instance Port Map for inst_m9
endmodule