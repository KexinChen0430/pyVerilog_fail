module MEMORY(
    input [9:0] ADDR,
    input CLK,
    input RE,
    input INIT,
    output reg [10:0] DATAOUT = 0
    );
    reg[11:0] storage[0:1023];
    always @(posedge CLK)
    begin
        DATAOUT <= (RE) ? storage[ADDR] : DATAOUT;
        // Pythom help us
        storage[0] <= (INIT) ? 12'd2048 : storage[0];
        storage[1] <= (INIT) ? 12'd2060 : storage[1];
        storage[2] <= (INIT) ? 12'd2073 : storage[2];
        storage[3] <= (INIT) ? 12'd2086 : storage[3];
        storage[4] <= (INIT) ? 12'd2099 : storage[4];
        storage[5] <= (INIT) ? 12'd2112 : storage[5];
        storage[6] <= (INIT) ? 12'd2125 : storage[6];
        storage[7] <= (INIT) ? 12'd2138 : storage[7];
        storage[8] <= (INIT) ? 12'd2150 : storage[8];
        storage[9] <= (INIT) ? 12'd2163 : storage[9];
        storage[10] <= (INIT) ? 12'd2176 : storage[10];
        storage[11] <= (INIT) ? 12'd2189 : storage[11];
        storage[12] <= (INIT) ? 12'd2202 : storage[12];
        storage[13] <= (INIT) ? 12'd2215 : storage[13];
        storage[14] <= (INIT) ? 12'd2227 : storage[14];
        storage[15] <= (INIT) ? 12'd2240 : storage[15];
        storage[16] <= (INIT) ? 12'd2253 : storage[16];
        storage[17] <= (INIT) ? 12'd2266 : storage[17];
        storage[18] <= (INIT) ? 12'd2279 : storage[18];
        storage[19] <= (INIT) ? 12'd2291 : storage[19];
        storage[20] <= (INIT) ? 12'd2304 : storage[20];
        storage[21] <= (INIT) ? 12'd2317 : storage[21];
        storage[22] <= (INIT) ? 12'd2330 : storage[22];
        storage[23] <= (INIT) ? 12'd2342 : storage[23];
        storage[24] <= (INIT) ? 12'd2355 : storage[24];
        storage[25] <= (INIT) ? 12'd2368 : storage[25];
        storage[26] <= (INIT) ? 12'd2380 : storage[26];
        storage[27] <= (INIT) ? 12'd2393 : storage[27];
        storage[28] <= (INIT) ? 12'd2406 : storage[28];
        storage[29] <= (INIT) ? 12'd2418 : storage[29];
        storage[30] <= (INIT) ? 12'd2431 : storage[30];
        storage[31] <= (INIT) ? 12'd2444 : storage[31];
        storage[32] <= (INIT) ? 12'd2456 : storage[32];
        storage[33] <= (INIT) ? 12'd2469 : storage[33];
        storage[34] <= (INIT) ? 12'd2481 : storage[34];
        storage[35] <= (INIT) ? 12'd2494 : storage[35];
        storage[36] <= (INIT) ? 12'd2507 : storage[36];
        storage[37] <= (INIT) ? 12'd2519 : storage[37];
        storage[38] <= (INIT) ? 12'd2532 : storage[38];
        storage[39] <= (INIT) ? 12'd2544 : storage[39];
        storage[40] <= (INIT) ? 12'd2557 : storage[40];
        storage[41] <= (INIT) ? 12'd2569 : storage[41];
        storage[42] <= (INIT) ? 12'd2581 : storage[42];
        storage[43] <= (INIT) ? 12'd2594 : storage[43];
        storage[44] <= (INIT) ? 12'd2606 : storage[44];
        storage[45] <= (INIT) ? 12'd2619 : storage[45];
        storage[46] <= (INIT) ? 12'd2631 : storage[46];
        storage[47] <= (INIT) ? 12'd2643 : storage[47];
        storage[48] <= (INIT) ? 12'd2656 : storage[48];
        storage[49] <= (INIT) ? 12'd2668 : storage[49];
        storage[50] <= (INIT) ? 12'd2680 : storage[50];
        storage[51] <= (INIT) ? 12'd2692 : storage[51];
        storage[52] <= (INIT) ? 12'd2704 : storage[52];
        storage[53] <= (INIT) ? 12'd2717 : storage[53];
        storage[54] <= (INIT) ? 12'd2729 : storage[54];
        storage[55] <= (INIT) ? 12'd2741 : storage[55];
        storage[56] <= (INIT) ? 12'd2753 : storage[56];
        storage[57] <= (INIT) ? 12'd2765 : storage[57];
        storage[58] <= (INIT) ? 12'd2777 : storage[58];
        storage[59] <= (INIT) ? 12'd2789 : storage[59];
        storage[60] <= (INIT) ? 12'd2801 : storage[60];
        storage[61] <= (INIT) ? 12'd2813 : storage[61];
        storage[62] <= (INIT) ? 12'd2825 : storage[62];
        storage[63] <= (INIT) ? 12'd2837 : storage[63];
        storage[64] <= (INIT) ? 12'd2849 : storage[64];
        storage[65] <= (INIT) ? 12'd2860 : storage[65];
        storage[66] <= (INIT) ? 12'd2872 : storage[66];
        storage[67] <= (INIT) ? 12'd2884 : storage[67];
        storage[68] <= (INIT) ? 12'd2896 : storage[68];
        storage[69] <= (INIT) ? 12'd2907 : storage[69];
        storage[70] <= (INIT) ? 12'd2919 : storage[70];
        storage[71] <= (INIT) ? 12'd2931 : storage[71];
        storage[72] <= (INIT) ? 12'd2942 : storage[72];
        storage[73] <= (INIT) ? 12'd2954 : storage[73];
        storage[74] <= (INIT) ? 12'd2965 : storage[74];
        storage[75] <= (INIT) ? 12'd2977 : storage[75];
        storage[76] <= (INIT) ? 12'd2988 : storage[76];
        storage[77] <= (INIT) ? 12'd3000 : storage[77];
        storage[78] <= (INIT) ? 12'd3011 : storage[78];
        storage[79] <= (INIT) ? 12'd3022 : storage[79];
        storage[80] <= (INIT) ? 12'd3034 : storage[80];
        storage[81] <= (INIT) ? 12'd3045 : storage[81];
        storage[82] <= (INIT) ? 12'd3056 : storage[82];
        storage[83] <= (INIT) ? 12'd3067 : storage[83];
        storage[84] <= (INIT) ? 12'd3078 : storage[84];
        storage[85] <= (INIT) ? 12'd3090 : storage[85];
        storage[86] <= (INIT) ? 12'd3101 : storage[86];
        storage[87] <= (INIT) ? 12'd3112 : storage[87];
        storage[88] <= (INIT) ? 12'd3123 : storage[88];
        storage[89] <= (INIT) ? 12'd3133 : storage[89];
        storage[90] <= (INIT) ? 12'd3144 : storage[90];
        storage[91] <= (INIT) ? 12'd3155 : storage[91];
        storage[92] <= (INIT) ? 12'd3166 : storage[92];
        storage[93] <= (INIT) ? 12'd3177 : storage[93];
        storage[94] <= (INIT) ? 12'd3187 : storage[94];
        storage[95] <= (INIT) ? 12'd3198 : storage[95];
        storage[96] <= (INIT) ? 12'd3209 : storage[96];
        storage[97] <= (INIT) ? 12'd3219 : storage[97];
        storage[98] <= (INIT) ? 12'd3230 : storage[98];
        storage[99] <= (INIT) ? 12'd3240 : storage[99];
        storage[100] <= (INIT) ? 12'd3251 : storage[100];
        storage[101] <= (INIT) ? 12'd3261 : storage[101];
        storage[102] <= (INIT) ? 12'd3271 : storage[102];
        storage[103] <= (INIT) ? 12'd3282 : storage[103];
        storage[104] <= (INIT) ? 12'd3292 : storage[104];
        storage[105] <= (INIT) ? 12'd3302 : storage[105];
        storage[106] <= (INIT) ? 12'd3312 : storage[106];
        storage[107] <= (INIT) ? 12'd3322 : storage[107];
        storage[108] <= (INIT) ? 12'd3332 : storage[108];
        storage[109] <= (INIT) ? 12'd3342 : storage[109];
        storage[110] <= (INIT) ? 12'd3352 : storage[110];
        storage[111] <= (INIT) ? 12'd3362 : storage[111];
        storage[112] <= (INIT) ? 12'd3372 : storage[112];
        storage[113] <= (INIT) ? 12'd3382 : storage[113];
        storage[114] <= (INIT) ? 12'd3392 : storage[114];
        storage[115] <= (INIT) ? 12'd3401 : storage[115];
        storage[116] <= (INIT) ? 12'd3411 : storage[116];
        storage[117] <= (INIT) ? 12'd3420 : storage[117];
        storage[118] <= (INIT) ? 12'd3430 : storage[118];
        storage[119] <= (INIT) ? 12'd3439 : storage[119];
        storage[120] <= (INIT) ? 12'd3449 : storage[120];
        storage[121] <= (INIT) ? 12'd3458 : storage[121];
        storage[122] <= (INIT) ? 12'd3468 : storage[122];
        storage[123] <= (INIT) ? 12'd3477 : storage[123];
        storage[124] <= (INIT) ? 12'd3486 : storage[124];
        storage[125] <= (INIT) ? 12'd3495 : storage[125];
        storage[126] <= (INIT) ? 12'd3504 : storage[126];
        storage[127] <= (INIT) ? 12'd3513 : storage[127];
        storage[128] <= (INIT) ? 12'd3522 : storage[128];
        storage[129] <= (INIT) ? 12'd3531 : storage[129];
        storage[130] <= (INIT) ? 12'd3540 : storage[130];
        storage[131] <= (INIT) ? 12'd3549 : storage[131];
        storage[132] <= (INIT) ? 12'd3557 : storage[132];
        storage[133] <= (INIT) ? 12'd3566 : storage[133];
        storage[134] <= (INIT) ? 12'd3575 : storage[134];
        storage[135] <= (INIT) ? 12'd3583 : storage[135];
        storage[136] <= (INIT) ? 12'd3592 : storage[136];
        storage[137] <= (INIT) ? 12'd3600 : storage[137];
        storage[138] <= (INIT) ? 12'd3608 : storage[138];
        storage[139] <= (INIT) ? 12'd3617 : storage[139];
        storage[140] <= (INIT) ? 12'd3625 : storage[140];
        storage[141] <= (INIT) ? 12'd3633 : storage[141];
        storage[142] <= (INIT) ? 12'd3641 : storage[142];
        storage[143] <= (INIT) ? 12'd3649 : storage[143];
        storage[144] <= (INIT) ? 12'd3657 : storage[144];
        storage[145] <= (INIT) ? 12'd3665 : storage[145];
        storage[146] <= (INIT) ? 12'd3673 : storage[146];
        storage[147] <= (INIT) ? 12'd3681 : storage[147];
        storage[148] <= (INIT) ? 12'd3689 : storage[148];
        storage[149] <= (INIT) ? 12'd3696 : storage[149];
        storage[150] <= (INIT) ? 12'd3704 : storage[150];
        storage[151] <= (INIT) ? 12'd3711 : storage[151];
        storage[152] <= (INIT) ? 12'd3719 : storage[152];
        storage[153] <= (INIT) ? 12'd3726 : storage[153];
        storage[154] <= (INIT) ? 12'd3734 : storage[154];
        storage[155] <= (INIT) ? 12'd3741 : storage[155];
        storage[156] <= (INIT) ? 12'd3748 : storage[156];
        storage[157] <= (INIT) ? 12'd3755 : storage[157];
        storage[158] <= (INIT) ? 12'd3762 : storage[158];
        storage[159] <= (INIT) ? 12'd3769 : storage[159];
        storage[160] <= (INIT) ? 12'd3776 : storage[160];
        storage[161] <= (INIT) ? 12'd3783 : storage[161];
        storage[162] <= (INIT) ? 12'd3790 : storage[162];
        storage[163] <= (INIT) ? 12'd3797 : storage[163];
        storage[164] <= (INIT) ? 12'd3803 : storage[164];
        storage[165] <= (INIT) ? 12'd3810 : storage[165];
        storage[166] <= (INIT) ? 12'd3816 : storage[166];
        storage[167] <= (INIT) ? 12'd3823 : storage[167];
        storage[168] <= (INIT) ? 12'd3829 : storage[168];
        storage[169] <= (INIT) ? 12'd3835 : storage[169];
        storage[170] <= (INIT) ? 12'd3842 : storage[170];
        storage[171] <= (INIT) ? 12'd3848 : storage[171];
        storage[172] <= (INIT) ? 12'd3854 : storage[172];
        storage[173] <= (INIT) ? 12'd3860 : storage[173];
        storage[174] <= (INIT) ? 12'd3866 : storage[174];
        storage[175] <= (INIT) ? 12'd3872 : storage[175];
        storage[176] <= (INIT) ? 12'd3878 : storage[176];
        storage[177] <= (INIT) ? 12'd3883 : storage[177];
        storage[178] <= (INIT) ? 12'd3889 : storage[178];
        storage[179] <= (INIT) ? 12'd3895 : storage[179];
        storage[180] <= (INIT) ? 12'd3900 : storage[180];
        storage[181] <= (INIT) ? 12'd3906 : storage[181];
        storage[182] <= (INIT) ? 12'd3911 : storage[182];
        storage[183] <= (INIT) ? 12'd3916 : storage[183];
        storage[184] <= (INIT) ? 12'd3921 : storage[184];
        storage[185] <= (INIT) ? 12'd3927 : storage[185];
        storage[186] <= (INIT) ? 12'd3932 : storage[186];
        storage[187] <= (INIT) ? 12'd3937 : storage[187];
        storage[188] <= (INIT) ? 12'd3942 : storage[188];
        storage[189] <= (INIT) ? 12'd3946 : storage[189];
        storage[190] <= (INIT) ? 12'd3951 : storage[190];
        storage[191] <= (INIT) ? 12'd3956 : storage[191];
        storage[192] <= (INIT) ? 12'd3961 : storage[192];
        storage[193] <= (INIT) ? 12'd3965 : storage[193];
        storage[194] <= (INIT) ? 12'd3970 : storage[194];
        storage[195] <= (INIT) ? 12'd3974 : storage[195];
        storage[196] <= (INIT) ? 12'd3978 : storage[196];
        storage[197] <= (INIT) ? 12'd3983 : storage[197];
        storage[198] <= (INIT) ? 12'd3987 : storage[198];
        storage[199] <= (INIT) ? 12'd3991 : storage[199];
        storage[200] <= (INIT) ? 12'd3995 : storage[200];
        storage[201] <= (INIT) ? 12'd3999 : storage[201];
        storage[202] <= (INIT) ? 12'd4003 : storage[202];
        storage[203] <= (INIT) ? 12'd4006 : storage[203];
        storage[204] <= (INIT) ? 12'd4010 : storage[204];
        storage[205] <= (INIT) ? 12'd4014 : storage[205];
        storage[206] <= (INIT) ? 12'd4017 : storage[206];
        storage[207] <= (INIT) ? 12'd4021 : storage[207];
        storage[208] <= (INIT) ? 12'd4024 : storage[208];
        storage[209] <= (INIT) ? 12'd4028 : storage[209];
        storage[210] <= (INIT) ? 12'd4031 : storage[210];
        storage[211] <= (INIT) ? 12'd4034 : storage[211];
        storage[212] <= (INIT) ? 12'd4037 : storage[212];
        storage[213] <= (INIT) ? 12'd4040 : storage[213];
        storage[214] <= (INIT) ? 12'd4043 : storage[214];
        storage[215] <= (INIT) ? 12'd4046 : storage[215];
        storage[216] <= (INIT) ? 12'd4049 : storage[216];
        storage[217] <= (INIT) ? 12'd4051 : storage[217];
        storage[218] <= (INIT) ? 12'd4054 : storage[218];
        storage[219] <= (INIT) ? 12'd4056 : storage[219];
        storage[220] <= (INIT) ? 12'd4059 : storage[220];
        storage[221] <= (INIT) ? 12'd4061 : storage[221];
        storage[222] <= (INIT) ? 12'd4064 : storage[222];
        storage[223] <= (INIT) ? 12'd4066 : storage[223];
        storage[224] <= (INIT) ? 12'd4068 : storage[224];
        storage[225] <= (INIT) ? 12'd4070 : storage[225];
        storage[226] <= (INIT) ? 12'd4072 : storage[226];
        storage[227] <= (INIT) ? 12'd4074 : storage[227];
        storage[228] <= (INIT) ? 12'd4076 : storage[228];
        storage[229] <= (INIT) ? 12'd4078 : storage[229];
        storage[230] <= (INIT) ? 12'd4079 : storage[230];
        storage[231] <= (INIT) ? 12'd4081 : storage[231];
        storage[232] <= (INIT) ? 12'd4082 : storage[232];
        storage[233] <= (INIT) ? 12'd4084 : storage[233];
        storage[234] <= (INIT) ? 12'd4085 : storage[234];
        storage[235] <= (INIT) ? 12'd4086 : storage[235];
        storage[236] <= (INIT) ? 12'd4087 : storage[236];
        storage[237] <= (INIT) ? 12'd4089 : storage[237];
        storage[238] <= (INIT) ? 12'd4090 : storage[238];
        storage[239] <= (INIT) ? 12'd4091 : storage[239];
        storage[240] <= (INIT) ? 12'd4091 : storage[240];
        storage[241] <= (INIT) ? 12'd4092 : storage[241];
        storage[242] <= (INIT) ? 12'd4093 : storage[242];
        storage[243] <= (INIT) ? 12'd4093 : storage[243];
        storage[244] <= (INIT) ? 12'd4094 : storage[244];
        storage[245] <= (INIT) ? 12'd4094 : storage[245];
        storage[246] <= (INIT) ? 12'd4095 : storage[246];
        storage[247] <= (INIT) ? 12'd4095 : storage[247];
        storage[248] <= (INIT) ? 12'd4095 : storage[248];
        storage[249] <= (INIT) ? 12'd4095 : storage[249];
        storage[250] <= (INIT) ? 12'd4095 : storage[250];
        storage[251] <= (INIT) ? 12'd4095 : storage[251];
        storage[252] <= (INIT) ? 12'd4095 : storage[252];
        storage[253] <= (INIT) ? 12'd4095 : storage[253];
        storage[254] <= (INIT) ? 12'd4095 : storage[254];
        storage[255] <= (INIT) ? 12'd4095 : storage[255];
        storage[256] <= (INIT) ? 12'd4094 : storage[256];
        storage[257] <= (INIT) ? 12'd4094 : storage[257];
        storage[258] <= (INIT) ? 12'd4093 : storage[258];
        storage[259] <= (INIT) ? 12'd4092 : storage[259];
        storage[260] <= (INIT) ? 12'd4092 : storage[260];
        storage[261] <= (INIT) ? 12'd4091 : storage[261];
        storage[262] <= (INIT) ? 12'd4090 : storage[262];
        storage[263] <= (INIT) ? 12'd4089 : storage[263];
        storage[264] <= (INIT) ? 12'd4088 : storage[264];
        storage[265] <= (INIT) ? 12'd4087 : storage[265];
        storage[266] <= (INIT) ? 12'd4085 : storage[266];
        storage[267] <= (INIT) ? 12'd4084 : storage[267];
        storage[268] <= (INIT) ? 12'd4083 : storage[268];
        storage[269] <= (INIT) ? 12'd4081 : storage[269];
        storage[270] <= (INIT) ? 12'd4080 : storage[270];
        storage[271] <= (INIT) ? 12'd4078 : storage[271];
        storage[272] <= (INIT) ? 12'd4076 : storage[272];
        storage[273] <= (INIT) ? 12'd4074 : storage[273];
        storage[274] <= (INIT) ? 12'd4073 : storage[274];
        storage[275] <= (INIT) ? 12'd4071 : storage[275];
        storage[276] <= (INIT) ? 12'd4069 : storage[276];
        storage[277] <= (INIT) ? 12'd4066 : storage[277];
        storage[278] <= (INIT) ? 12'd4064 : storage[278];
        storage[279] <= (INIT) ? 12'd4062 : storage[279];
        storage[280] <= (INIT) ? 12'd4060 : storage[280];
        storage[281] <= (INIT) ? 12'd4057 : storage[281];
        storage[282] <= (INIT) ? 12'd4055 : storage[282];
        storage[283] <= (INIT) ? 12'd4052 : storage[283];
        storage[284] <= (INIT) ? 12'd4049 : storage[284];
        storage[285] <= (INIT) ? 12'd4047 : storage[285];
        storage[286] <= (INIT) ? 12'd4044 : storage[286];
        storage[287] <= (INIT) ? 12'd4041 : storage[287];
        storage[288] <= (INIT) ? 12'd4038 : storage[288];
        storage[289] <= (INIT) ? 12'd4035 : storage[289];
        storage[290] <= (INIT) ? 12'd4032 : storage[290];
        storage[291] <= (INIT) ? 12'd4028 : storage[291];
        storage[292] <= (INIT) ? 12'd4025 : storage[292];
        storage[293] <= (INIT) ? 12'd4022 : storage[293];
        storage[294] <= (INIT) ? 12'd4018 : storage[294];
        storage[295] <= (INIT) ? 12'd4015 : storage[295];
        storage[296] <= (INIT) ? 12'd4011 : storage[296];
        storage[297] <= (INIT) ? 12'd4007 : storage[297];
        storage[298] <= (INIT) ? 12'd4004 : storage[298];
        storage[299] <= (INIT) ? 12'd4000 : storage[299];
        storage[300] <= (INIT) ? 12'd3996 : storage[300];
        storage[301] <= (INIT) ? 12'd3992 : storage[301];
        storage[302] <= (INIT) ? 12'd3988 : storage[302];
        storage[303] <= (INIT) ? 12'd3984 : storage[303];
        storage[304] <= (INIT) ? 12'd3979 : storage[304];
        storage[305] <= (INIT) ? 12'd3975 : storage[305];
        storage[306] <= (INIT) ? 12'd3971 : storage[306];
        storage[307] <= (INIT) ? 12'd3966 : storage[307];
        storage[308] <= (INIT) ? 12'd3962 : storage[308];
        storage[309] <= (INIT) ? 12'd3957 : storage[309];
        storage[310] <= (INIT) ? 12'd3952 : storage[310];
        storage[311] <= (INIT) ? 12'd3948 : storage[311];
        storage[312] <= (INIT) ? 12'd3943 : storage[312];
        storage[313] <= (INIT) ? 12'd3938 : storage[313];
        storage[314] <= (INIT) ? 12'd3933 : storage[314];
        storage[315] <= (INIT) ? 12'd3928 : storage[315];
        storage[316] <= (INIT) ? 12'd3923 : storage[316];
        storage[317] <= (INIT) ? 12'd3918 : storage[317];
        storage[318] <= (INIT) ? 12'd3912 : storage[318];
        storage[319] <= (INIT) ? 12'd3907 : storage[319];
        storage[320] <= (INIT) ? 12'd3901 : storage[320];
        storage[321] <= (INIT) ? 12'd3896 : storage[321];
        storage[322] <= (INIT) ? 12'd3890 : storage[322];
        storage[323] <= (INIT) ? 12'd3885 : storage[323];
        storage[324] <= (INIT) ? 12'd3879 : storage[324];
        storage[325] <= (INIT) ? 12'd3873 : storage[325];
        storage[326] <= (INIT) ? 12'd3867 : storage[326];
        storage[327] <= (INIT) ? 12'd3861 : storage[327];
        storage[328] <= (INIT) ? 12'd3855 : storage[328];
        storage[329] <= (INIT) ? 12'd3849 : storage[329];
        storage[330] <= (INIT) ? 12'd3843 : storage[330];
        storage[331] <= (INIT) ? 12'd3837 : storage[331];
        storage[332] <= (INIT) ? 12'd3831 : storage[332];
        storage[333] <= (INIT) ? 12'd3824 : storage[333];
        storage[334] <= (INIT) ? 12'd3818 : storage[334];
        storage[335] <= (INIT) ? 12'd3811 : storage[335];
        storage[336] <= (INIT) ? 12'd3805 : storage[336];
        storage[337] <= (INIT) ? 12'd3798 : storage[337];
        storage[338] <= (INIT) ? 12'd3791 : storage[338];
        storage[339] <= (INIT) ? 12'd3785 : storage[339];
        storage[340] <= (INIT) ? 12'd3778 : storage[340];
        storage[341] <= (INIT) ? 12'd3771 : storage[341];
        storage[342] <= (INIT) ? 12'd3764 : storage[342];
        storage[343] <= (INIT) ? 12'd3757 : storage[343];
        storage[344] <= (INIT) ? 12'd3750 : storage[344];
        storage[345] <= (INIT) ? 12'd3743 : storage[345];
        storage[346] <= (INIT) ? 12'd3735 : storage[346];
        storage[347] <= (INIT) ? 12'd3728 : storage[347];
        storage[348] <= (INIT) ? 12'd3721 : storage[348];
        storage[349] <= (INIT) ? 12'd3713 : storage[349];
        storage[350] <= (INIT) ? 12'd3706 : storage[350];
        storage[351] <= (INIT) ? 12'd3698 : storage[351];
        storage[352] <= (INIT) ? 12'd3690 : storage[352];
        storage[353] <= (INIT) ? 12'd3683 : storage[353];
        storage[354] <= (INIT) ? 12'd3675 : storage[354];
        storage[355] <= (INIT) ? 12'd3667 : storage[355];
        storage[356] <= (INIT) ? 12'd3659 : storage[356];
        storage[357] <= (INIT) ? 12'd3651 : storage[357];
        storage[358] <= (INIT) ? 12'd3643 : storage[358];
        storage[359] <= (INIT) ? 12'd3635 : storage[359];
        storage[360] <= (INIT) ? 12'd3627 : storage[360];
        storage[361] <= (INIT) ? 12'd3619 : storage[361];
        storage[362] <= (INIT) ? 12'd3611 : storage[362];
        storage[363] <= (INIT) ? 12'd3602 : storage[363];
        storage[364] <= (INIT) ? 12'd3594 : storage[364];
        storage[365] <= (INIT) ? 12'd3585 : storage[365];
        storage[366] <= (INIT) ? 12'd3577 : storage[366];
        storage[367] <= (INIT) ? 12'd3568 : storage[367];
        storage[368] <= (INIT) ? 12'd3560 : storage[368];
        storage[369] <= (INIT) ? 12'd3551 : storage[369];
        storage[370] <= (INIT) ? 12'd3542 : storage[370];
        storage[371] <= (INIT) ? 12'd3533 : storage[371];
        storage[372] <= (INIT) ? 12'd3524 : storage[372];
        storage[373] <= (INIT) ? 12'd3515 : storage[373];
        storage[374] <= (INIT) ? 12'd3506 : storage[374];
        storage[375] <= (INIT) ? 12'd3497 : storage[375];
        storage[376] <= (INIT) ? 12'd3488 : storage[376];
        storage[377] <= (INIT) ? 12'd3479 : storage[377];
        storage[378] <= (INIT) ? 12'd3470 : storage[378];
        storage[379] <= (INIT) ? 12'd3461 : storage[379];
        storage[380] <= (INIT) ? 12'd3451 : storage[380];
        storage[381] <= (INIT) ? 12'd3442 : storage[381];
        storage[382] <= (INIT) ? 12'd3432 : storage[382];
        storage[383] <= (INIT) ? 12'd3423 : storage[383];
        storage[384] <= (INIT) ? 12'd3413 : storage[384];
        storage[385] <= (INIT) ? 12'd3404 : storage[385];
        storage[386] <= (INIT) ? 12'd3394 : storage[386];
        storage[387] <= (INIT) ? 12'd3384 : storage[387];
        storage[388] <= (INIT) ? 12'd3375 : storage[388];
        storage[389] <= (INIT) ? 12'd3365 : storage[389];
        storage[390] <= (INIT) ? 12'd3355 : storage[390];
        storage[391] <= (INIT) ? 12'd3345 : storage[391];
        storage[392] <= (INIT) ? 12'd3335 : storage[392];
        storage[393] <= (INIT) ? 12'd3325 : storage[393];
        storage[394] <= (INIT) ? 12'd3315 : storage[394];
        storage[395] <= (INIT) ? 12'd3305 : storage[395];
        storage[396] <= (INIT) ? 12'd3295 : storage[396];
        storage[397] <= (INIT) ? 12'd3284 : storage[397];
        storage[398] <= (INIT) ? 12'd3274 : storage[398];
        storage[399] <= (INIT) ? 12'd3264 : storage[399];
        storage[400] <= (INIT) ? 12'd3253 : storage[400];
        storage[401] <= (INIT) ? 12'd3243 : storage[401];
        storage[402] <= (INIT) ? 12'd3233 : storage[402];
        storage[403] <= (INIT) ? 12'd3222 : storage[403];
        storage[404] <= (INIT) ? 12'd3211 : storage[404];
        storage[405] <= (INIT) ? 12'd3201 : storage[405];
        storage[406] <= (INIT) ? 12'd3190 : storage[406];
        storage[407] <= (INIT) ? 12'd3179 : storage[407];
        storage[408] <= (INIT) ? 12'd3169 : storage[408];
        storage[409] <= (INIT) ? 12'd3158 : storage[409];
        storage[410] <= (INIT) ? 12'd3147 : storage[410];
        storage[411] <= (INIT) ? 12'd3136 : storage[411];
        storage[412] <= (INIT) ? 12'd3125 : storage[412];
        storage[413] <= (INIT) ? 12'd3114 : storage[413];
        storage[414] <= (INIT) ? 12'd3103 : storage[414];
        storage[415] <= (INIT) ? 12'd3092 : storage[415];
        storage[416] <= (INIT) ? 12'd3081 : storage[416];
        storage[417] <= (INIT) ? 12'd3070 : storage[417];
        storage[418] <= (INIT) ? 12'd3059 : storage[418];
        storage[419] <= (INIT) ? 12'd3048 : storage[419];
        storage[420] <= (INIT) ? 12'd3037 : storage[420];
        storage[421] <= (INIT) ? 12'd3025 : storage[421];
        storage[422] <= (INIT) ? 12'd3014 : storage[422];
        storage[423] <= (INIT) ? 12'd3003 : storage[423];
        storage[424] <= (INIT) ? 12'd2991 : storage[424];
        storage[425] <= (INIT) ? 12'd2980 : storage[425];
        storage[426] <= (INIT) ? 12'd2968 : storage[426];
        storage[427] <= (INIT) ? 12'd2957 : storage[427];
        storage[428] <= (INIT) ? 12'd2945 : storage[428];
        storage[429] <= (INIT) ? 12'd2934 : storage[429];
        storage[430] <= (INIT) ? 12'd2922 : storage[430];
        storage[431] <= (INIT) ? 12'd2910 : storage[431];
        storage[432] <= (INIT) ? 12'd2899 : storage[432];
        storage[433] <= (INIT) ? 12'd2887 : storage[433];
        storage[434] <= (INIT) ? 12'd2875 : storage[434];
        storage[435] <= (INIT) ? 12'd2863 : storage[435];
        storage[436] <= (INIT) ? 12'd2852 : storage[436];
        storage[437] <= (INIT) ? 12'd2840 : storage[437];
        storage[438] <= (INIT) ? 12'd2828 : storage[438];
        storage[439] <= (INIT) ? 12'd2816 : storage[439];
        storage[440] <= (INIT) ? 12'd2804 : storage[440];
        storage[441] <= (INIT) ? 12'd2792 : storage[441];
        storage[442] <= (INIT) ? 12'd2780 : storage[442];
        storage[443] <= (INIT) ? 12'd2768 : storage[443];
        storage[444] <= (INIT) ? 12'd2756 : storage[444];
        storage[445] <= (INIT) ? 12'd2744 : storage[445];
        storage[446] <= (INIT) ? 12'd2732 : storage[446];
        storage[447] <= (INIT) ? 12'd2720 : storage[447];
        storage[448] <= (INIT) ? 12'd2708 : storage[448];
        storage[449] <= (INIT) ? 12'd2695 : storage[449];
        storage[450] <= (INIT) ? 12'd2683 : storage[450];
        storage[451] <= (INIT) ? 12'd2671 : storage[451];
        storage[452] <= (INIT) ? 12'd2659 : storage[452];
        storage[453] <= (INIT) ? 12'd2646 : storage[453];
        storage[454] <= (INIT) ? 12'd2634 : storage[454];
        storage[455] <= (INIT) ? 12'd2622 : storage[455];
        storage[456] <= (INIT) ? 12'd2609 : storage[456];
        storage[457] <= (INIT) ? 12'd2597 : storage[457];
        storage[458] <= (INIT) ? 12'd2585 : storage[458];
        storage[459] <= (INIT) ? 12'd2572 : storage[459];
        storage[460] <= (INIT) ? 12'd2560 : storage[460];
        storage[461] <= (INIT) ? 12'd2547 : storage[461];
        storage[462] <= (INIT) ? 12'd2535 : storage[462];
        storage[463] <= (INIT) ? 12'd2522 : storage[463];
        storage[464] <= (INIT) ? 12'd2510 : storage[464];
        storage[465] <= (INIT) ? 12'd2497 : storage[465];
        storage[466] <= (INIT) ? 12'd2485 : storage[466];
        storage[467] <= (INIT) ? 12'd2472 : storage[467];
        storage[468] <= (INIT) ? 12'd2459 : storage[468];
        storage[469] <= (INIT) ? 12'd2447 : storage[469];
        storage[470] <= (INIT) ? 12'd2434 : storage[470];
        storage[471] <= (INIT) ? 12'd2422 : storage[471];
        storage[472] <= (INIT) ? 12'd2409 : storage[472];
        storage[473] <= (INIT) ? 12'd2396 : storage[473];
        storage[474] <= (INIT) ? 12'd2384 : storage[474];
        storage[475] <= (INIT) ? 12'd2371 : storage[475];
        storage[476] <= (INIT) ? 12'd2358 : storage[476];
        storage[477] <= (INIT) ? 12'd2346 : storage[477];
        storage[478] <= (INIT) ? 12'd2333 : storage[478];
        storage[479] <= (INIT) ? 12'd2320 : storage[479];
        storage[480] <= (INIT) ? 12'd2307 : storage[480];
        storage[481] <= (INIT) ? 12'd2295 : storage[481];
        storage[482] <= (INIT) ? 12'd2282 : storage[482];
        storage[483] <= (INIT) ? 12'd2269 : storage[483];
        storage[484] <= (INIT) ? 12'd2256 : storage[484];
        storage[485] <= (INIT) ? 12'd2243 : storage[485];
        storage[486] <= (INIT) ? 12'd2231 : storage[486];
        storage[487] <= (INIT) ? 12'd2218 : storage[487];
        storage[488] <= (INIT) ? 12'd2205 : storage[488];
        storage[489] <= (INIT) ? 12'd2192 : storage[489];
        storage[490] <= (INIT) ? 12'd2179 : storage[490];
        storage[491] <= (INIT) ? 12'd2166 : storage[491];
        storage[492] <= (INIT) ? 12'd2154 : storage[492];
        storage[493] <= (INIT) ? 12'd2141 : storage[493];
        storage[494] <= (INIT) ? 12'd2128 : storage[494];
        storage[495] <= (INIT) ? 12'd2115 : storage[495];
        storage[496] <= (INIT) ? 12'd2102 : storage[496];
        storage[497] <= (INIT) ? 12'd2089 : storage[497];
        storage[498] <= (INIT) ? 12'd2076 : storage[498];
        storage[499] <= (INIT) ? 12'd2064 : storage[499];
        storage[500] <= (INIT) ? 12'd2051 : storage[500];
        storage[501] <= (INIT) ? 12'd2038 : storage[501];
        storage[502] <= (INIT) ? 12'd2025 : storage[502];
        storage[503] <= (INIT) ? 12'd2012 : storage[503];
        storage[504] <= (INIT) ? 12'd1999 : storage[504];
        storage[505] <= (INIT) ? 12'd1986 : storage[505];
        storage[506] <= (INIT) ? 12'd1974 : storage[506];
        storage[507] <= (INIT) ? 12'd1961 : storage[507];
        storage[508] <= (INIT) ? 12'd1948 : storage[508];
        storage[509] <= (INIT) ? 12'd1935 : storage[509];
        storage[510] <= (INIT) ? 12'd1922 : storage[510];
        storage[511] <= (INIT) ? 12'd1909 : storage[511];
        storage[512] <= (INIT) ? 12'd1897 : storage[512];
        storage[513] <= (INIT) ? 12'd1884 : storage[513];
        storage[514] <= (INIT) ? 12'd1871 : storage[514];
        storage[515] <= (INIT) ? 12'd1858 : storage[515];
        storage[516] <= (INIT) ? 12'd1845 : storage[516];
        storage[517] <= (INIT) ? 12'd1833 : storage[517];
        storage[518] <= (INIT) ? 12'd1820 : storage[518];
        storage[519] <= (INIT) ? 12'd1807 : storage[519];
        storage[520] <= (INIT) ? 12'd1794 : storage[520];
        storage[521] <= (INIT) ? 12'd1781 : storage[521];
        storage[522] <= (INIT) ? 12'd1769 : storage[522];
        storage[523] <= (INIT) ? 12'd1756 : storage[523];
        storage[524] <= (INIT) ? 12'd1743 : storage[524];
        storage[525] <= (INIT) ? 12'd1731 : storage[525];
        storage[526] <= (INIT) ? 12'd1718 : storage[526];
        storage[527] <= (INIT) ? 12'd1705 : storage[527];
        storage[528] <= (INIT) ? 12'd1692 : storage[528];
        storage[529] <= (INIT) ? 12'd1680 : storage[529];
        storage[530] <= (INIT) ? 12'd1667 : storage[530];
        storage[531] <= (INIT) ? 12'd1655 : storage[531];
        storage[532] <= (INIT) ? 12'd1642 : storage[532];
        storage[533] <= (INIT) ? 12'd1629 : storage[533];
        storage[534] <= (INIT) ? 12'd1617 : storage[534];
        storage[535] <= (INIT) ? 12'd1604 : storage[535];
        storage[536] <= (INIT) ? 12'd1592 : storage[536];
        storage[537] <= (INIT) ? 12'd1579 : storage[537];
        storage[538] <= (INIT) ? 12'd1567 : storage[538];
        storage[539] <= (INIT) ? 12'd1554 : storage[539];
        storage[540] <= (INIT) ? 12'd1542 : storage[540];
        storage[541] <= (INIT) ? 12'd1529 : storage[541];
        storage[542] <= (INIT) ? 12'd1517 : storage[542];
        storage[543] <= (INIT) ? 12'd1504 : storage[543];
        storage[544] <= (INIT) ? 12'd1492 : storage[544];
        storage[545] <= (INIT) ? 12'd1480 : storage[545];
        storage[546] <= (INIT) ? 12'd1467 : storage[546];
        storage[547] <= (INIT) ? 12'd1455 : storage[547];
        storage[548] <= (INIT) ? 12'd1443 : storage[548];
        storage[549] <= (INIT) ? 12'd1430 : storage[549];
        storage[550] <= (INIT) ? 12'd1418 : storage[550];
        storage[551] <= (INIT) ? 12'd1406 : storage[551];
        storage[552] <= (INIT) ? 12'd1394 : storage[552];
        storage[553] <= (INIT) ? 12'd1381 : storage[553];
        storage[554] <= (INIT) ? 12'd1369 : storage[554];
        storage[555] <= (INIT) ? 12'd1357 : storage[555];
        storage[556] <= (INIT) ? 12'd1345 : storage[556];
        storage[557] <= (INIT) ? 12'd1333 : storage[557];
        storage[558] <= (INIT) ? 12'd1321 : storage[558];
        storage[559] <= (INIT) ? 12'd1309 : storage[559];
        storage[560] <= (INIT) ? 12'd1297 : storage[560];
        storage[561] <= (INIT) ? 12'd1285 : storage[561];
        storage[562] <= (INIT) ? 12'd1273 : storage[562];
        storage[563] <= (INIT) ? 12'd1261 : storage[563];
        storage[564] <= (INIT) ? 12'd1249 : storage[564];
        storage[565] <= (INIT) ? 12'd1238 : storage[565];
        storage[566] <= (INIT) ? 12'd1226 : storage[566];
        storage[567] <= (INIT) ? 12'd1214 : storage[567];
        storage[568] <= (INIT) ? 12'd1202 : storage[568];
        storage[569] <= (INIT) ? 12'd1191 : storage[569];
        storage[570] <= (INIT) ? 12'd1179 : storage[570];
        storage[571] <= (INIT) ? 12'd1167 : storage[571];
        storage[572] <= (INIT) ? 12'd1156 : storage[572];
        storage[573] <= (INIT) ? 12'd1144 : storage[573];
        storage[574] <= (INIT) ? 12'd1133 : storage[574];
        storage[575] <= (INIT) ? 12'd1121 : storage[575];
        storage[576] <= (INIT) ? 12'd1110 : storage[576];
        storage[577] <= (INIT) ? 12'd1098 : storage[577];
        storage[578] <= (INIT) ? 12'd1087 : storage[578];
        storage[579] <= (INIT) ? 12'd1075 : storage[579];
        storage[580] <= (INIT) ? 12'd1064 : storage[580];
        storage[581] <= (INIT) ? 12'd1053 : storage[581];
        storage[582] <= (INIT) ? 12'd1042 : storage[582];
        storage[583] <= (INIT) ? 12'd1031 : storage[583];
        storage[584] <= (INIT) ? 12'd1019 : storage[584];
        storage[585] <= (INIT) ? 12'd1008 : storage[585];
        storage[586] <= (INIT) ? 12'd997 : storage[586];
        storage[587] <= (INIT) ? 12'd986 : storage[587];
        storage[588] <= (INIT) ? 12'd975 : storage[588];
        storage[589] <= (INIT) ? 12'd964 : storage[589];
        storage[590] <= (INIT) ? 12'd953 : storage[590];
        storage[591] <= (INIT) ? 12'd943 : storage[591];
        storage[592] <= (INIT) ? 12'd932 : storage[592];
        storage[593] <= (INIT) ? 12'd921 : storage[593];
        storage[594] <= (INIT) ? 12'd910 : storage[594];
        storage[595] <= (INIT) ? 12'd900 : storage[595];
        storage[596] <= (INIT) ? 12'd889 : storage[596];
        storage[597] <= (INIT) ? 12'd878 : storage[597];
        storage[598] <= (INIT) ? 12'd868 : storage[598];
        storage[599] <= (INIT) ? 12'd857 : storage[599];
        storage[600] <= (INIT) ? 12'd847 : storage[600];
        storage[601] <= (INIT) ? 12'd836 : storage[601];
        storage[602] <= (INIT) ? 12'd826 : storage[602];
        storage[603] <= (INIT) ? 12'd816 : storage[603];
        storage[604] <= (INIT) ? 12'd806 : storage[604];
        storage[605] <= (INIT) ? 12'd795 : storage[605];
        storage[606] <= (INIT) ? 12'd785 : storage[606];
        storage[607] <= (INIT) ? 12'd775 : storage[607];
        storage[608] <= (INIT) ? 12'd765 : storage[608];
        storage[609] <= (INIT) ? 12'd755 : storage[609];
        storage[610] <= (INIT) ? 12'd745 : storage[610];
        storage[611] <= (INIT) ? 12'd735 : storage[611];
        storage[612] <= (INIT) ? 12'd725 : storage[612];
        storage[613] <= (INIT) ? 12'd716 : storage[613];
        storage[614] <= (INIT) ? 12'd706 : storage[614];
        storage[615] <= (INIT) ? 12'd696 : storage[615];
        storage[616] <= (INIT) ? 12'd687 : storage[616];
        storage[617] <= (INIT) ? 12'd677 : storage[617];
        storage[618] <= (INIT) ? 12'd667 : storage[618];
        storage[619] <= (INIT) ? 12'd658 : storage[619];
        storage[620] <= (INIT) ? 12'd648 : storage[620];
        storage[621] <= (INIT) ? 12'd639 : storage[621];
        storage[622] <= (INIT) ? 12'd630 : storage[622];
        storage[623] <= (INIT) ? 12'd621 : storage[623];
        storage[624] <= (INIT) ? 12'd611 : storage[624];
        storage[625] <= (INIT) ? 12'd602 : storage[625];
        storage[626] <= (INIT) ? 12'd593 : storage[626];
        storage[627] <= (INIT) ? 12'd584 : storage[627];
        storage[628] <= (INIT) ? 12'd575 : storage[628];
        storage[629] <= (INIT) ? 12'd566 : storage[629];
        storage[630] <= (INIT) ? 12'd557 : storage[630];
        storage[631] <= (INIT) ? 12'd549 : storage[631];
        storage[632] <= (INIT) ? 12'd540 : storage[632];
        storage[633] <= (INIT) ? 12'd531 : storage[633];
        storage[634] <= (INIT) ? 12'd523 : storage[634];
        storage[635] <= (INIT) ? 12'd514 : storage[635];
        storage[636] <= (INIT) ? 12'd506 : storage[636];
        storage[637] <= (INIT) ? 12'd497 : storage[637];
        storage[638] <= (INIT) ? 12'd489 : storage[638];
        storage[639] <= (INIT) ? 12'd480 : storage[639];
        storage[640] <= (INIT) ? 12'd472 : storage[640];
        storage[641] <= (INIT) ? 12'd464 : storage[641];
        storage[642] <= (INIT) ? 12'd456 : storage[642];
        storage[643] <= (INIT) ? 12'd448 : storage[643];
        storage[644] <= (INIT) ? 12'd440 : storage[644];
        storage[645] <= (INIT) ? 12'd432 : storage[645];
        storage[646] <= (INIT) ? 12'd424 : storage[646];
        storage[647] <= (INIT) ? 12'd416 : storage[647];
        storage[648] <= (INIT) ? 12'd408 : storage[648];
        storage[649] <= (INIT) ? 12'd401 : storage[649];
        storage[650] <= (INIT) ? 12'd393 : storage[650];
        storage[651] <= (INIT) ? 12'd386 : storage[651];
        storage[652] <= (INIT) ? 12'd378 : storage[652];
        storage[653] <= (INIT) ? 12'd371 : storage[653];
        storage[654] <= (INIT) ? 12'd363 : storage[654];
        storage[655] <= (INIT) ? 12'd356 : storage[655];
        storage[656] <= (INIT) ? 12'd349 : storage[656];
        storage[657] <= (INIT) ? 12'd342 : storage[657];
        storage[658] <= (INIT) ? 12'd335 : storage[658];
        storage[659] <= (INIT) ? 12'd328 : storage[659];
        storage[660] <= (INIT) ? 12'd321 : storage[660];
        storage[661] <= (INIT) ? 12'd314 : storage[661];
        storage[662] <= (INIT) ? 12'd307 : storage[662];
        storage[663] <= (INIT) ? 12'd300 : storage[663];
        storage[664] <= (INIT) ? 12'd294 : storage[664];
        storage[665] <= (INIT) ? 12'd287 : storage[665];
        storage[666] <= (INIT) ? 12'd280 : storage[666];
        storage[667] <= (INIT) ? 12'd274 : storage[667];
        storage[668] <= (INIT) ? 12'd268 : storage[668];
        storage[669] <= (INIT) ? 12'd261 : storage[669];
        storage[670] <= (INIT) ? 12'd255 : storage[670];
        storage[671] <= (INIT) ? 12'd249 : storage[671];
        storage[672] <= (INIT) ? 12'd243 : storage[672];
        storage[673] <= (INIT) ? 12'd237 : storage[673];
        storage[674] <= (INIT) ? 12'd231 : storage[674];
        storage[675] <= (INIT) ? 12'd225 : storage[675];
        storage[676] <= (INIT) ? 12'd219 : storage[676];
        storage[677] <= (INIT) ? 12'd213 : storage[677];
        storage[678] <= (INIT) ? 12'd207 : storage[678];
        storage[679] <= (INIT) ? 12'd202 : storage[679];
        storage[680] <= (INIT) ? 12'd196 : storage[680];
        storage[681] <= (INIT) ? 12'd191 : storage[681];
        storage[682] <= (INIT) ? 12'd185 : storage[682];
        storage[683] <= (INIT) ? 12'd180 : storage[683];
        storage[684] <= (INIT) ? 12'd175 : storage[684];
        storage[685] <= (INIT) ? 12'd170 : storage[685];
        storage[686] <= (INIT) ? 12'd165 : storage[686];
        storage[687] <= (INIT) ? 12'd160 : storage[687];
        storage[688] <= (INIT) ? 12'd155 : storage[688];
        storage[689] <= (INIT) ? 12'd150 : storage[689];
        storage[690] <= (INIT) ? 12'd145 : storage[690];
        storage[691] <= (INIT) ? 12'd140 : storage[691];
        storage[692] <= (INIT) ? 12'd136 : storage[692];
        storage[693] <= (INIT) ? 12'd131 : storage[693];
        storage[694] <= (INIT) ? 12'd127 : storage[694];
        storage[695] <= (INIT) ? 12'd122 : storage[695];
        storage[696] <= (INIT) ? 12'd118 : storage[696];
        storage[697] <= (INIT) ? 12'd114 : storage[697];
        storage[698] <= (INIT) ? 12'd109 : storage[698];
        storage[699] <= (INIT) ? 12'd105 : storage[699];
        storage[700] <= (INIT) ? 12'd101 : storage[700];
        storage[701] <= (INIT) ? 12'd97 : storage[701];
        storage[702] <= (INIT) ? 12'd93 : storage[702];
        storage[703] <= (INIT) ? 12'd89 : storage[703];
        storage[704] <= (INIT) ? 12'd86 : storage[704];
        storage[705] <= (INIT) ? 12'd82 : storage[705];
        storage[706] <= (INIT) ? 12'd79 : storage[706];
        storage[707] <= (INIT) ? 12'd75 : storage[707];
        storage[708] <= (INIT) ? 12'd72 : storage[708];
        storage[709] <= (INIT) ? 12'd68 : storage[709];
        storage[710] <= (INIT) ? 12'd65 : storage[710];
        storage[711] <= (INIT) ? 12'd62 : storage[711];
        storage[712] <= (INIT) ? 12'd59 : storage[712];
        storage[713] <= (INIT) ? 12'd56 : storage[713];
        storage[714] <= (INIT) ? 12'd53 : storage[714];
        storage[715] <= (INIT) ? 12'd50 : storage[715];
        storage[716] <= (INIT) ? 12'd47 : storage[716];
        storage[717] <= (INIT) ? 12'd44 : storage[717];
        storage[718] <= (INIT) ? 12'd42 : storage[718];
        storage[719] <= (INIT) ? 12'd39 : storage[719];
        storage[720] <= (INIT) ? 12'd37 : storage[720];
        storage[721] <= (INIT) ? 12'd34 : storage[721];
        storage[722] <= (INIT) ? 12'd32 : storage[722];
        storage[723] <= (INIT) ? 12'd30 : storage[723];
        storage[724] <= (INIT) ? 12'd28 : storage[724];
        storage[725] <= (INIT) ? 12'd25 : storage[725];
        storage[726] <= (INIT) ? 12'd23 : storage[726];
        storage[727] <= (INIT) ? 12'd22 : storage[727];
        storage[728] <= (INIT) ? 12'd20 : storage[728];
        storage[729] <= (INIT) ? 12'd18 : storage[729];
        storage[730] <= (INIT) ? 12'd16 : storage[730];
        storage[731] <= (INIT) ? 12'd15 : storage[731];
        storage[732] <= (INIT) ? 12'd13 : storage[732];
        storage[733] <= (INIT) ? 12'd12 : storage[733];
        storage[734] <= (INIT) ? 12'd10 : storage[734];
        storage[735] <= (INIT) ? 12'd9 : storage[735];
        storage[736] <= (INIT) ? 12'd8 : storage[736];
        storage[737] <= (INIT) ? 12'd7 : storage[737];
        storage[738] <= (INIT) ? 12'd6 : storage[738];
        storage[739] <= (INIT) ? 12'd5 : storage[739];
        storage[740] <= (INIT) ? 12'd4 : storage[740];
        storage[741] <= (INIT) ? 12'd3 : storage[741];
        storage[742] <= (INIT) ? 12'd2 : storage[742];
        storage[743] <= (INIT) ? 12'd2 : storage[743];
        storage[744] <= (INIT) ? 12'd1 : storage[744];
        storage[745] <= (INIT) ? 12'd1 : storage[745];
        storage[746] <= (INIT) ? 12'd0 : storage[746];
        storage[747] <= (INIT) ? 12'd0 : storage[747];
        storage[748] <= (INIT) ? 12'd0 : storage[748];
        storage[749] <= (INIT) ? 12'd0 : storage[749];
        storage[750] <= (INIT) ? 12'd0 : storage[750];
        storage[751] <= (INIT) ? 12'd0 : storage[751];
        storage[752] <= (INIT) ? 12'd0 : storage[752];
        storage[753] <= (INIT) ? 12'd0 : storage[753];
        storage[754] <= (INIT) ? 12'd0 : storage[754];
        storage[755] <= (INIT) ? 12'd0 : storage[755];
        storage[756] <= (INIT) ? 12'd1 : storage[756];
        storage[757] <= (INIT) ? 12'd1 : storage[757];
        storage[758] <= (INIT) ? 12'd2 : storage[758];
        storage[759] <= (INIT) ? 12'd2 : storage[759];
        storage[760] <= (INIT) ? 12'd3 : storage[760];
        storage[761] <= (INIT) ? 12'd4 : storage[761];
        storage[762] <= (INIT) ? 12'd5 : storage[762];
        storage[763] <= (INIT) ? 12'd6 : storage[763];
        storage[764] <= (INIT) ? 12'd7 : storage[764];
        storage[765] <= (INIT) ? 12'd8 : storage[765];
        storage[766] <= (INIT) ? 12'd9 : storage[766];
        storage[767] <= (INIT) ? 12'd11 : storage[767];
        storage[768] <= (INIT) ? 12'd12 : storage[768];
        storage[769] <= (INIT) ? 12'd13 : storage[769];
        storage[770] <= (INIT) ? 12'd15 : storage[770];
        storage[771] <= (INIT) ? 12'd17 : storage[771];
        storage[772] <= (INIT) ? 12'd18 : storage[772];
        storage[773] <= (INIT) ? 12'd20 : storage[773];
        storage[774] <= (INIT) ? 12'd22 : storage[774];
        storage[775] <= (INIT) ? 12'd24 : storage[775];
        storage[776] <= (INIT) ? 12'd26 : storage[776];
        storage[777] <= (INIT) ? 12'd28 : storage[777];
        storage[778] <= (INIT) ? 12'd30 : storage[778];
        storage[779] <= (INIT) ? 12'd32 : storage[779];
        storage[780] <= (INIT) ? 12'd35 : storage[780];
        storage[781] <= (INIT) ? 12'd37 : storage[781];
        storage[782] <= (INIT) ? 12'd40 : storage[782];
        storage[783] <= (INIT) ? 12'd42 : storage[783];
        storage[784] <= (INIT) ? 12'd45 : storage[784];
        storage[785] <= (INIT) ? 12'd48 : storage[785];
        storage[786] <= (INIT) ? 12'd51 : storage[786];
        storage[787] <= (INIT) ? 12'd53 : storage[787];
        storage[788] <= (INIT) ? 12'd56 : storage[788];
        storage[789] <= (INIT) ? 12'd59 : storage[789];
        storage[790] <= (INIT) ? 12'd63 : storage[790];
        storage[791] <= (INIT) ? 12'd66 : storage[791];
        storage[792] <= (INIT) ? 12'd69 : storage[792];
        storage[793] <= (INIT) ? 12'd72 : storage[793];
        storage[794] <= (INIT) ? 12'd76 : storage[794];
        storage[795] <= (INIT) ? 12'd79 : storage[795];
        storage[796] <= (INIT) ? 12'd83 : storage[796];
        storage[797] <= (INIT) ? 12'd87 : storage[797];
        storage[798] <= (INIT) ? 12'd90 : storage[798];
        storage[799] <= (INIT) ? 12'd94 : storage[799];
        storage[800] <= (INIT) ? 12'd98 : storage[800];
        storage[801] <= (INIT) ? 12'd102 : storage[801];
        storage[802] <= (INIT) ? 12'd106 : storage[802];
        storage[803] <= (INIT) ? 12'd110 : storage[803];
        storage[804] <= (INIT) ? 12'd115 : storage[804];
        storage[805] <= (INIT) ? 12'd119 : storage[805];
        storage[806] <= (INIT) ? 12'd123 : storage[806];
        storage[807] <= (INIT) ? 12'd128 : storage[807];
        storage[808] <= (INIT) ? 12'd132 : storage[808];
        storage[809] <= (INIT) ? 12'd137 : storage[809];
        storage[810] <= (INIT) ? 12'd141 : storage[810];
        storage[811] <= (INIT) ? 12'd146 : storage[811];
        storage[812] <= (INIT) ? 12'd151 : storage[812];
        storage[813] <= (INIT) ? 12'd156 : storage[813];
        storage[814] <= (INIT) ? 12'd161 : storage[814];
        storage[815] <= (INIT) ? 12'd166 : storage[815];
        storage[816] <= (INIT) ? 12'd171 : storage[816];
        storage[817] <= (INIT) ? 12'd176 : storage[817];
        storage[818] <= (INIT) ? 12'd181 : storage[818];
        storage[819] <= (INIT) ? 12'd187 : storage[819];
        storage[820] <= (INIT) ? 12'd192 : storage[820];
        storage[821] <= (INIT) ? 12'd198 : storage[821];
        storage[822] <= (INIT) ? 12'd203 : storage[822];
        storage[823] <= (INIT) ? 12'd209 : storage[823];
        storage[824] <= (INIT) ? 12'd215 : storage[824];
        storage[825] <= (INIT) ? 12'd220 : storage[825];
        storage[826] <= (INIT) ? 12'd226 : storage[826];
        storage[827] <= (INIT) ? 12'd232 : storage[827];
        storage[828] <= (INIT) ? 12'd238 : storage[828];
        storage[829] <= (INIT) ? 12'd244 : storage[829];
        storage[830] <= (INIT) ? 12'd250 : storage[830];
        storage[831] <= (INIT) ? 12'd256 : storage[831];
        storage[832] <= (INIT) ? 12'd263 : storage[832];
        storage[833] <= (INIT) ? 12'd269 : storage[833];
        storage[834] <= (INIT) ? 12'd275 : storage[834];
        storage[835] <= (INIT) ? 12'd282 : storage[835];
        storage[836] <= (INIT) ? 12'd288 : storage[836];
        storage[837] <= (INIT) ? 12'd295 : storage[837];
        storage[838] <= (INIT) ? 12'd302 : storage[838];
        storage[839] <= (INIT) ? 12'd309 : storage[839];
        storage[840] <= (INIT) ? 12'd315 : storage[840];
        storage[841] <= (INIT) ? 12'd322 : storage[841];
        storage[842] <= (INIT) ? 12'd329 : storage[842];
        storage[843] <= (INIT) ? 12'd336 : storage[843];
        storage[844] <= (INIT) ? 12'd343 : storage[844];
        storage[845] <= (INIT) ? 12'd351 : storage[845];
        storage[846] <= (INIT) ? 12'd358 : storage[846];
        storage[847] <= (INIT) ? 12'd365 : storage[847];
        storage[848] <= (INIT) ? 12'd372 : storage[848];
        storage[849] <= (INIT) ? 12'd380 : storage[849];
        storage[850] <= (INIT) ? 12'd387 : storage[850];
        storage[851] <= (INIT) ? 12'd395 : storage[851];
        storage[852] <= (INIT) ? 12'd403 : storage[852];
        storage[853] <= (INIT) ? 12'd410 : storage[853];
        storage[854] <= (INIT) ? 12'd418 : storage[854];
        storage[855] <= (INIT) ? 12'd426 : storage[855];
        storage[856] <= (INIT) ? 12'd434 : storage[856];
        storage[857] <= (INIT) ? 12'd442 : storage[857];
        storage[858] <= (INIT) ? 12'd450 : storage[858];
        storage[859] <= (INIT) ? 12'd458 : storage[859];
        storage[860] <= (INIT) ? 12'd466 : storage[860];
        storage[861] <= (INIT) ? 12'd474 : storage[861];
        storage[862] <= (INIT) ? 12'd482 : storage[862];
        storage[863] <= (INIT) ? 12'd491 : storage[863];
        storage[864] <= (INIT) ? 12'd499 : storage[864];
        storage[865] <= (INIT) ? 12'd508 : storage[865];
        storage[866] <= (INIT) ? 12'd516 : storage[866];
        storage[867] <= (INIT) ? 12'd525 : storage[867];
        storage[868] <= (INIT) ? 12'd533 : storage[868];
        storage[869] <= (INIT) ? 12'd542 : storage[869];
        storage[870] <= (INIT) ? 12'd551 : storage[870];
        storage[871] <= (INIT) ? 12'd560 : storage[871];
        storage[872] <= (INIT) ? 12'd568 : storage[872];
        storage[873] <= (INIT) ? 12'd577 : storage[873];
        storage[874] <= (INIT) ? 12'd586 : storage[874];
        storage[875] <= (INIT) ? 12'd595 : storage[875];
        storage[876] <= (INIT) ? 12'd604 : storage[876];
        storage[877] <= (INIT) ? 12'd614 : storage[877];
        storage[878] <= (INIT) ? 12'd623 : storage[878];
        storage[879] <= (INIT) ? 12'd632 : storage[879];
        storage[880] <= (INIT) ? 12'd641 : storage[880];
        storage[881] <= (INIT) ? 12'd651 : storage[881];
        storage[882] <= (INIT) ? 12'd660 : storage[882];
        storage[883] <= (INIT) ? 12'd670 : storage[883];
        storage[884] <= (INIT) ? 12'd679 : storage[884];
        storage[885] <= (INIT) ? 12'd689 : storage[885];
        storage[886] <= (INIT) ? 12'd698 : storage[886];
        storage[887] <= (INIT) ? 12'd708 : storage[887];
        storage[888] <= (INIT) ? 12'd718 : storage[888];
        storage[889] <= (INIT) ? 12'd728 : storage[889];
        storage[890] <= (INIT) ? 12'd738 : storage[890];
        storage[891] <= (INIT) ? 12'd747 : storage[891];
        storage[892] <= (INIT) ? 12'd757 : storage[892];
        storage[893] <= (INIT) ? 12'd767 : storage[893];
        storage[894] <= (INIT) ? 12'd778 : storage[894];
        storage[895] <= (INIT) ? 12'd788 : storage[895];
        storage[896] <= (INIT) ? 12'd798 : storage[896];
        storage[897] <= (INIT) ? 12'd808 : storage[897];
        storage[898] <= (INIT) ? 12'd818 : storage[898];
        storage[899] <= (INIT) ? 12'd829 : storage[899];
        storage[900] <= (INIT) ? 12'd839 : storage[900];
        storage[901] <= (INIT) ? 12'd849 : storage[901];
        storage[902] <= (INIT) ? 12'd860 : storage[902];
        storage[903] <= (INIT) ? 12'd870 : storage[903];
        storage[904] <= (INIT) ? 12'd881 : storage[904];
        storage[905] <= (INIT) ? 12'd891 : storage[905];
        storage[906] <= (INIT) ? 12'd902 : storage[906];
        storage[907] <= (INIT) ? 12'd913 : storage[907];
        storage[908] <= (INIT) ? 12'd924 : storage[908];
        storage[909] <= (INIT) ? 12'd934 : storage[909];
        storage[910] <= (INIT) ? 12'd945 : storage[910];
        storage[911] <= (INIT) ? 12'd956 : storage[911];
        storage[912] <= (INIT) ? 12'd967 : storage[912];
        storage[913] <= (INIT) ? 12'd978 : storage[913];
        storage[914] <= (INIT) ? 12'd989 : storage[914];
        storage[915] <= (INIT) ? 12'd1000 : storage[915];
        storage[916] <= (INIT) ? 12'd1011 : storage[916];
        storage[917] <= (INIT) ? 12'd1022 : storage[917];
        storage[918] <= (INIT) ? 12'd1033 : storage[918];
        storage[919] <= (INIT) ? 12'd1044 : storage[919];
        storage[920] <= (INIT) ? 12'd1056 : storage[920];
        storage[921] <= (INIT) ? 12'd1067 : storage[921];
        storage[922] <= (INIT) ? 12'd1078 : storage[922];
        storage[923] <= (INIT) ? 12'd1090 : storage[923];
        storage[924] <= (INIT) ? 12'd1101 : storage[924];
        storage[925] <= (INIT) ? 12'd1112 : storage[925];
        storage[926] <= (INIT) ? 12'd1124 : storage[926];
        storage[927] <= (INIT) ? 12'd1135 : storage[927];
        storage[928] <= (INIT) ? 12'd1147 : storage[928];
        storage[929] <= (INIT) ? 12'd1158 : storage[929];
        storage[930] <= (INIT) ? 12'd1170 : storage[930];
        storage[931] <= (INIT) ? 12'd1182 : storage[931];
        storage[932] <= (INIT) ? 12'd1193 : storage[932];
        storage[933] <= (INIT) ? 12'd1205 : storage[933];
        storage[934] <= (INIT) ? 12'd1217 : storage[934];
        storage[935] <= (INIT) ? 12'd1229 : storage[935];
        storage[936] <= (INIT) ? 12'd1240 : storage[936];
        storage[937] <= (INIT) ? 12'd1252 : storage[937];
        storage[938] <= (INIT) ? 12'd1264 : storage[938];
        storage[939] <= (INIT) ? 12'd1276 : storage[939];
        storage[940] <= (INIT) ? 12'd1288 : storage[940];
        storage[941] <= (INIT) ? 12'd1300 : storage[941];
        storage[942] <= (INIT) ? 12'd1312 : storage[942];
        storage[943] <= (INIT) ? 12'd1324 : storage[943];
        storage[944] <= (INIT) ? 12'd1336 : storage[944];
        storage[945] <= (INIT) ? 12'd1348 : storage[945];
        storage[946] <= (INIT) ? 12'd1360 : storage[946];
        storage[947] <= (INIT) ? 12'd1372 : storage[947];
        storage[948] <= (INIT) ? 12'd1384 : storage[948];
        storage[949] <= (INIT) ? 12'd1397 : storage[949];
        storage[950] <= (INIT) ? 12'd1409 : storage[950];
        storage[951] <= (INIT) ? 12'd1421 : storage[951];
        storage[952] <= (INIT) ? 12'd1433 : storage[952];
        storage[953] <= (INIT) ? 12'd1446 : storage[953];
        storage[954] <= (INIT) ? 12'd1458 : storage[954];
        storage[955] <= (INIT) ? 12'd1470 : storage[955];
        storage[956] <= (INIT) ? 12'd1482 : storage[956];
        storage[957] <= (INIT) ? 12'd1495 : storage[957];
        storage[958] <= (INIT) ? 12'd1507 : storage[958];
        storage[959] <= (INIT) ? 12'd1520 : storage[959];
        storage[960] <= (INIT) ? 12'd1532 : storage[960];
        storage[961] <= (INIT) ? 12'd1545 : storage[961];
        storage[962] <= (INIT) ? 12'd1557 : storage[962];
        storage[963] <= (INIT) ? 12'd1570 : storage[963];
        storage[964] <= (INIT) ? 12'd1582 : storage[964];
        storage[965] <= (INIT) ? 12'd1595 : storage[965];
        storage[966] <= (INIT) ? 12'd1607 : storage[966];
        storage[967] <= (INIT) ? 12'd1620 : storage[967];
        storage[968] <= (INIT) ? 12'd1632 : storage[968];
        storage[969] <= (INIT) ? 12'd1645 : storage[969];
        storage[970] <= (INIT) ? 12'd1658 : storage[970];
        storage[971] <= (INIT) ? 12'd1670 : storage[971];
        storage[972] <= (INIT) ? 12'd1683 : storage[972];
        storage[973] <= (INIT) ? 12'd1695 : storage[973];
        storage[974] <= (INIT) ? 12'd1708 : storage[974];
        storage[975] <= (INIT) ? 12'd1721 : storage[975];
        storage[976] <= (INIT) ? 12'd1734 : storage[976];
        storage[977] <= (INIT) ? 12'd1746 : storage[977];
        storage[978] <= (INIT) ? 12'd1759 : storage[978];
        storage[979] <= (INIT) ? 12'd1772 : storage[979];
        storage[980] <= (INIT) ? 12'd1784 : storage[980];
        storage[981] <= (INIT) ? 12'd1797 : storage[981];
        storage[982] <= (INIT) ? 12'd1810 : storage[982];
        storage[983] <= (INIT) ? 12'd1823 : storage[983];
        storage[984] <= (INIT) ? 12'd1836 : storage[984];
        storage[985] <= (INIT) ? 12'd1848 : storage[985];
        storage[986] <= (INIT) ? 12'd1861 : storage[986];
        storage[987] <= (INIT) ? 12'd1874 : storage[987];
        storage[988] <= (INIT) ? 12'd1887 : storage[988];
        storage[989] <= (INIT) ? 12'd1900 : storage[989];
        storage[990] <= (INIT) ? 12'd1912 : storage[990];
        storage[991] <= (INIT) ? 12'd1925 : storage[991];
        storage[992] <= (INIT) ? 12'd1938 : storage[992];
        storage[993] <= (INIT) ? 12'd1951 : storage[993];
        storage[994] <= (INIT) ? 12'd1964 : storage[994];
        storage[995] <= (INIT) ? 12'd1977 : storage[995];
        storage[996] <= (INIT) ? 12'd1990 : storage[996];
        storage[997] <= (INIT) ? 12'd2002 : storage[997];
        storage[998] <= (INIT) ? 12'd2015 : storage[998];
        storage[999] <= (INIT) ? 12'd2028 : storage[999];
        storage[1000] <= (INIT) ? 12'd0 : storage[1000];
        storage[1001] <= (INIT) ? 12'd0 : storage[1001];
        storage[1002] <= (INIT) ? 12'd0 : storage[1002];
        storage[1003] <= (INIT) ? 12'd0 : storage[1003];
        storage[1004] <= (INIT) ? 12'd0 : storage[1004];
        storage[1005] <= (INIT) ? 12'd0 : storage[1005];
        storage[1006] <= (INIT) ? 12'd0 : storage[1006];
        storage[1007] <= (INIT) ? 12'd0 : storage[1007];
        storage[1008] <= (INIT) ? 12'd0 : storage[1008];
        storage[1009] <= (INIT) ? 12'd0 : storage[1009];
        storage[1010] <= (INIT) ? 12'd0 : storage[1010];
        storage[1011] <= (INIT) ? 12'd0 : storage[1011];
        storage[1012] <= (INIT) ? 12'd0 : storage[1012];
        storage[1013] <= (INIT) ? 12'd0 : storage[1013];
        storage[1014] <= (INIT) ? 12'd0 : storage[1014];
        storage[1015] <= (INIT) ? 12'd0 : storage[1015];
        storage[1016] <= (INIT) ? 12'd0 : storage[1016];
        storage[1017] <= (INIT) ? 12'd0 : storage[1017];
        storage[1018] <= (INIT) ? 12'd0 : storage[1018];
        storage[1019] <= (INIT) ? 12'd0 : storage[1019];
        storage[1020] <= (INIT) ? 12'd0 : storage[1020];
        storage[1021] <= (INIT) ? 12'd0 : storage[1021];
        storage[1022] <= (INIT) ? 12'd0 : storage[1022];
        storage[1023] <= (INIT) ? 12'd0 : storage[1023];
    end
endmodule