module sky130_fd_sc_lp__iso0n (
    //# {{data|Data Signals}}
    input  A      ,
    output X      ,
    //# {{power|Power}}
    input  SLEEP_B,
    input  KAGND  ,
    input  VPB    ,
    input  VPWR   ,
    input  VNB
);
endmodule