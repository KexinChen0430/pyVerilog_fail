module
					nextState = s0;
				else
					nextState = s5;
			end
		endcase
	end
endmodule