module IB(
	(* iopad_external_pin *) input I,
	output O);
	assign O = I;
endmodule