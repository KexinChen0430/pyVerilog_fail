module XOR2_X1 (A, B, Z);
  input A;
  input B;
  output Z;
  xor(Z, A, B);
  specify
    if((B == 1'b0)) (A => Z) = (0.1, 0.1);
    if((B == 1'b1)) (A => Z) = (0.1, 0.1);
    if((A == 1'b0)) (B => Z) = (0.1, 0.1);
    if((A == 1'b1)) (B => Z) = (0.1, 0.1);
  endspecify
endmodule