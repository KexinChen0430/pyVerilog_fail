module ieee_ops (
  clk, ce, result, operation, a, b
)/* synthesis syn_black_box syn_noprune=1 */;
  input clk;
  input ce;
  output [31 : 0] result;
  input [5 : 0] operation;
  input [31 : 0] a;
  input [31 : 0] b;
  // synthesis translate_off
  wire sig00000001;
  wire sig00000002;
  wire sig00000003;
  wire sig00000004;
  wire sig00000005;
  wire sig00000006;
  wire sig00000007;
  wire sig00000008;
  wire sig00000009;
  wire sig0000000a;
  wire sig0000000b;
  wire sig0000000c;
  wire sig0000000d;
  wire sig0000000e;
  wire sig0000000f;
  wire sig00000010;
  wire sig00000011;
  wire sig00000012;
  wire sig00000013;
  wire sig00000014;
  wire sig00000015;
  wire sig00000016;
  wire sig00000017;
  wire sig00000018;
  wire sig00000019;
  wire sig0000001a;
  wire sig0000001b;
  wire sig0000001c;
  wire sig0000001d;
  wire sig0000001e;
  wire sig0000001f;
  wire sig00000020;
  wire sig00000021;
  wire sig00000022;
  wire sig00000023;
  wire sig00000024;
  wire sig00000025;
  wire sig00000026;
  wire sig00000027;
  wire sig00000028;
  wire sig00000029;
  wire sig0000002a;
  wire sig0000002b;
  wire sig0000002c;
  wire sig0000002d;
  wire sig0000002e;
  wire sig0000002f;
  wire sig00000030;
  wire sig00000031;
  wire sig00000032;
  wire sig00000033;
  wire sig00000034;
  wire sig00000035;
  wire sig00000036;
  wire sig00000037;
  wire sig00000038;
  wire sig00000039;
  wire sig0000003a;
  wire sig0000003b;
  wire sig0000003c;
  wire sig0000003d;
  wire sig0000003e;
  wire sig0000003f;
  wire sig00000040;
  wire sig00000041;
  wire sig00000042;
  wire sig00000043;
  wire sig00000044;
  wire sig00000045;
  wire sig00000046;
  wire sig00000047;
  wire sig00000048;
  wire sig00000049;
  wire sig0000004a;
  wire sig0000004b;
  wire sig0000004c;
  wire sig0000004d;
  wire sig0000004e;
  wire sig0000004f;
  wire sig00000050;
  wire sig00000051;
  wire sig00000052;
  wire sig00000053;
  wire sig00000054;
  wire sig00000055;
  wire sig00000056;
  wire sig00000057;
  wire sig00000058;
  wire sig00000059;
  wire sig0000005a;
  wire sig0000005b;
  wire sig0000005c;
  wire sig0000005d;
  wire sig0000005e;
  wire sig0000005f;
  wire sig00000060;
  wire sig00000061;
  wire sig00000062;
  wire sig00000063;
  wire sig00000064;
  wire sig00000065;
  wire sig00000066;
  wire sig00000067;
  wire sig00000068;
  wire sig00000069;
  wire sig0000006a;
  wire sig0000006b;
  wire sig0000006c;
  wire sig0000006d;
  wire sig0000006e;
  wire sig0000006f;
  wire sig00000070;
  wire sig00000071;
  wire sig00000072;
  wire sig00000073;
  wire sig00000074;
  wire sig00000075;
  wire sig00000076;
  wire sig00000077;
  wire sig00000078;
  wire sig00000079;
  wire sig0000007a;
  wire sig0000007b;
  wire sig0000007c;
  wire sig0000007d;
  wire sig0000007e;
  wire sig0000007f;
  wire sig00000080;
  wire sig00000081;
  wire sig00000082;
  wire sig00000083;
  wire sig00000084;
  wire sig00000085;
  wire sig00000086;
  wire sig00000087;
  wire sig00000088;
  wire sig00000089;
  wire sig0000008a;
  wire sig0000008b;
  wire sig0000008c;
  wire sig0000008d;
  wire sig0000008e;
  wire sig0000008f;
  wire sig00000090;
  wire sig00000091;
  wire sig00000092;
  wire sig00000093;
  wire sig00000094;
  wire sig00000095;
  wire sig00000096;
  wire sig00000097;
  wire sig00000098;
  wire sig00000099;
  wire sig0000009a;
  wire sig0000009b;
  wire sig0000009c;
  wire sig0000009d;
  wire sig0000009e;
  wire sig0000009f;
  wire sig000000a0;
  wire sig000000a1;
  wire sig000000a2;
  wire sig000000a3;
  wire sig000000a4;
  wire sig000000a5;
  wire sig000000a6;
  wire sig000000a7;
  wire sig000000a8;
  wire sig000000a9;
  wire sig000000aa;
  wire sig000000ab;
  wire sig000000ac;
  wire sig000000ad;
  wire sig000000ae;
  wire sig000000af;
  wire sig000000b0;
  wire sig000000b1;
  wire sig000000b2;
  wire sig000000b3;
  wire sig000000b4;
  wire sig000000b5;
  wire sig000000b6;
  wire sig000000b7;
  wire sig000000b8;
  wire sig000000b9;
  wire sig000000ba;
  wire sig000000bb;
  wire sig000000bc;
  wire sig000000bd;
  wire sig000000be;
  wire sig000000bf;
  wire sig000000c0;
  wire sig000000c1;
  wire sig000000c2;
  wire sig000000c3;
  wire sig000000c4;
  wire sig000000c5;
  wire sig000000c6;
  wire sig000000c7;
  wire sig000000c8;
  wire sig000000c9;
  wire sig000000ca;
  wire sig000000cb;
  wire sig000000cc;
  wire sig000000cd;
  wire sig000000ce;
  wire sig000000cf;
  wire sig000000d0;
  wire sig000000d1;
  wire sig000000d2;
  wire sig000000d3;
  wire sig000000d4;
  wire sig000000d5;
  wire sig000000d6;
  wire sig000000d7;
  wire sig000000d8;
  wire sig000000d9;
  wire sig000000da;
  wire sig000000db;
  wire sig000000dc;
  wire sig000000dd;
  wire sig000000de;
  wire sig000000df;
  wire sig000000e0;
  wire sig000000e1;
  wire sig000000e2;
  wire sig000000e3;
  wire sig000000e4;
  wire sig000000e5;
  wire sig000000e6;
  wire sig000000e7;
  wire sig000000e8;
  wire sig000000e9;
  wire sig000000ea;
  wire sig000000eb;
  wire sig000000ec;
  wire sig000000ed;
  wire sig000000ee;
  wire sig000000ef;
  wire sig000000f0;
  wire sig000000f1;
  wire sig000000f2;
  wire sig000000f3;
  wire sig000000f4;
  wire sig000000f5;
  wire sig000000f6;
  wire sig000000f7;
  wire sig000000f8;
  wire sig000000f9;
  wire sig000000fa;
  wire sig000000fb;
  wire sig000000fc;
  wire sig000000fd;
  wire sig000000fe;
  wire sig000000ff;
  wire sig00000100;
  wire sig00000101;
  wire sig00000102;
  wire sig00000103;
  wire sig00000104;
  wire sig00000105;
  wire sig00000106;
  wire sig00000107;
  wire sig00000108;
  wire sig00000109;
  wire sig0000010a;
  wire sig0000010b;
  wire sig0000010c;
  wire sig0000010d;
  wire sig0000010e;
  wire sig0000010f;
  wire sig00000110;
  wire sig00000111;
  wire sig00000112;
  wire sig00000113;
  wire sig00000114;
  wire sig00000115;
  wire sig00000116;
  wire sig00000117;
  wire sig00000118;
  wire sig00000119;
  wire sig0000011a;
  wire sig0000011b;
  wire sig0000011c;
  wire sig0000011d;
  wire sig0000011e;
  wire sig0000011f;
  wire sig00000120;
  wire sig00000121;
  wire sig00000122;
  wire sig00000123;
  wire sig00000124;
  wire sig00000125;
  wire sig00000126;
  wire sig00000127;
  wire sig00000128;
  wire sig00000129;
  wire sig0000012a;
  wire sig0000012b;
  wire sig0000012c;
  wire sig0000012d;
  wire sig0000012e;
  wire sig0000012f;
  wire sig00000130;
  wire sig00000131;
  wire sig00000132;
  wire sig00000133;
  wire sig00000134;
  wire sig00000135;
  wire sig00000136;
  wire sig00000137;
  wire sig00000138;
  wire sig00000139;
  wire sig0000013a;
  wire sig0000013b;
  wire sig0000013c;
  wire sig0000013d;
  wire sig0000013e;
  wire sig0000013f;
  wire sig00000140;
  wire sig00000141;
  wire sig00000142;
  wire sig00000143;
  wire sig00000144;
  wire sig00000145;
  wire sig00000146;
  wire sig00000147;
  wire sig00000148;
  wire sig00000149;
  wire sig0000014a;
  wire sig0000014b;
  wire sig0000014c;
  wire sig0000014d;
  wire sig0000014e;
  wire sig0000014f;
  wire sig00000150;
  wire sig00000151;
  wire sig00000152;
  wire sig00000153;
  wire sig00000154;
  wire sig00000155;
  wire sig00000156;
  wire sig00000157;
  wire sig00000158;
  wire sig00000159;
  wire sig0000015a;
  wire sig0000015b;
  wire sig0000015c;
  wire sig0000015d;
  wire sig0000015e;
  wire sig0000015f;
  wire sig00000160;
  wire sig00000161;
  wire sig00000162;
  wire sig00000163;
  wire sig00000164;
  wire sig00000165;
  wire sig00000166;
  wire sig00000167;
  wire sig00000168;
  wire sig00000169;
  wire sig0000016a;
  wire sig0000016b;
  wire sig0000016c;
  wire sig0000016d;
  wire sig0000016e;
  wire sig0000016f;
  wire sig00000170;
  wire sig00000171;
  wire sig00000172;
  wire sig00000173;
  wire sig00000174;
  wire sig00000175;
  wire sig00000176;
  wire sig00000177;
  wire sig00000178;
  wire sig00000179;
  wire sig0000017a;
  wire sig0000017b;
  wire sig0000017c;
  wire sig0000017d;
  wire sig0000017e;
  wire sig0000017f;
  wire sig00000180;
  wire sig00000181;
  wire sig00000182;
  wire sig00000183;
  wire sig00000184;
  wire sig00000185;
  wire sig00000186;
  wire sig00000187;
  wire sig00000188;
  wire sig00000189;
  wire sig0000018a;
  wire sig0000018b;
  wire sig0000018c;
  wire sig0000018d;
  wire sig0000018e;
  wire sig0000018f;
  wire sig00000190;
  wire sig00000191;
  wire sig00000192;
  wire sig00000193;
  wire sig00000194;
  wire sig00000195;
  wire sig00000196;
  wire sig00000197;
  wire sig00000198;
  wire sig00000199;
  wire sig0000019a;
  wire sig0000019b;
  wire sig0000019c;
  wire sig0000019d;
  wire sig0000019e;
  wire sig0000019f;
  wire sig000001a0;
  wire sig000001a1;
  wire sig000001a2;
  wire sig000001a3;
  wire sig000001a4;
  wire sig000001a5;
  wire sig000001a6;
  wire sig000001a7;
  wire sig000001a8;
  wire sig000001a9;
  wire sig000001aa;
  wire sig000001ab;
  wire sig000001ac;
  wire sig000001ad;
  wire sig000001ae;
  wire sig000001af;
  wire sig000001b0;
  wire sig000001b1;
  wire sig000001b2;
  wire sig000001b3;
  wire sig000001b4;
  wire sig000001b5;
  wire sig000001b6;
  wire sig000001b7;
  wire sig000001b8;
  wire sig000001b9;
  wire sig000001ba;
  wire sig000001bb;
  wire sig000001bc;
  wire sig000001bd;
  wire sig000001be;
  wire sig000001bf;
  wire sig000001c0;
  wire sig000001c1;
  wire sig000001c2;
  wire sig000001c3;
  wire sig000001c4;
  wire sig000001c5;
  wire sig000001c6;
  wire sig000001c7;
  wire sig000001c8;
  wire sig000001c9;
  wire sig000001ca;
  wire sig000001cb;
  wire sig000001cc;
  wire sig000001cd;
  wire sig000001ce;
  wire sig000001cf;
  wire sig000001d0;
  wire sig000001d1;
  wire sig000001d2;
  wire sig000001d3;
  wire sig000001d4;
  wire sig000001d5;
  wire sig000001d6;
  wire sig000001d7;
  wire sig000001d8;
  wire sig000001d9;
  wire sig000001da;
  wire sig000001db;
  wire sig000001dc;
  wire sig000001dd;
  wire sig000001de;
  wire sig000001df;
  wire sig000001e0;
  wire sig000001e1;
  wire sig000001e2;
  wire sig000001e3;
  wire sig000001e4;
  wire sig000001e5;
  wire sig000001e6;
  wire sig000001e7;
  wire sig000001e8;
  wire sig000001e9;
  wire sig000001ea;
  wire sig000001eb;
  wire sig000001ec;
  wire sig000001ed;
  wire sig000001ee;
  wire sig000001ef;
  wire sig000001f0;
  wire sig000001f1;
  wire sig000001f2;
  wire sig000001f3;
  wire sig000001f4;
  wire sig000001f5;
  wire sig000001f6;
  wire sig000001f7;
  wire sig000001f8;
  wire sig000001f9;
  wire sig000001fa;
  wire sig000001fb;
  wire sig000001fc;
  wire sig000001fd;
  wire sig000001fe;
  wire sig000001ff;
  wire sig00000200;
  wire sig00000201;
  wire sig00000202;
  wire sig00000203;
  wire sig00000204;
  wire sig00000205;
  wire sig00000206;
  wire sig00000207;
  wire sig00000208;
  wire sig00000209;
  wire sig0000020a;
  wire sig0000020b;
  wire sig0000020c;
  wire sig0000020d;
  wire sig0000020e;
  wire sig0000020f;
  wire sig00000210;
  wire sig00000211;
  wire sig00000212;
  wire sig00000213;
  wire sig00000214;
  wire sig00000215;
  wire sig00000216;
  wire sig00000217;
  wire sig00000218;
  wire sig00000219;
  wire sig0000021a;
  wire sig0000021b;
  wire sig0000021c;
  wire sig0000021d;
  wire sig0000021e;
  wire sig0000021f;
  wire sig00000220;
  wire sig00000221;
  wire sig00000222;
  wire sig00000223;
  wire sig00000224;
  wire sig00000225;
  wire sig00000226;
  wire sig00000227;
  wire sig00000228;
  wire sig00000229;
  wire sig0000022a;
  wire sig0000022b;
  wire sig0000022c;
  wire sig0000022d;
  wire sig0000022e;
  wire sig0000022f;
  wire sig00000230;
  wire sig00000231;
  wire sig00000232;
  wire sig00000233;
  wire sig00000234;
  wire sig00000235;
  wire sig00000236;
  wire sig00000237;
  wire sig00000238;
  wire sig00000239;
  wire sig0000023a;
  wire sig0000023b;
  wire sig0000023c;
  wire sig0000023d;
  wire sig0000023e;
  wire sig0000023f;
  wire sig00000240;
  wire sig00000241;
  wire sig00000242;
  wire sig00000243;
  wire sig00000244;
  wire sig00000245;
  wire sig00000246;
  wire sig00000247;
  wire sig00000248;
  wire sig00000249;
  wire sig0000024a;
  wire sig0000024b;
  wire sig0000024c;
  wire sig0000024d;
  wire sig0000024e;
  wire sig0000024f;
  wire sig00000250;
  wire sig00000251;
  wire sig00000252;
  wire sig00000253;
  wire sig00000254;
  wire sig00000255;
  wire sig00000256;
  wire sig00000257;
  wire sig00000258;
  wire sig00000259;
  wire sig0000025a;
  wire sig0000025b;
  wire sig0000025c;
  wire sig0000025d;
  wire sig0000025e;
  wire sig0000025f;
  wire sig00000260;
  wire sig00000261;
  wire sig00000262;
  wire sig00000263;
  wire sig00000264;
  wire sig00000265;
  wire sig00000266;
  wire sig00000267;
  wire sig00000268;
  wire sig00000269;
  wire sig0000026a;
  wire sig0000026b;
  wire sig0000026c;
  wire sig0000026d;
  wire sig0000026e;
  wire sig0000026f;
  wire sig00000270;
  wire sig00000271;
  wire sig00000272;
  wire sig00000273;
  wire sig00000274;
  wire sig00000275;
  wire sig00000276;
  wire sig00000277;
  wire sig00000278;
  wire sig00000279;
  wire sig0000027a;
  wire sig0000027b;
  wire sig0000027c;
  wire sig0000027d;
  wire sig0000027e;
  wire sig0000027f;
  wire sig00000280;
  wire sig00000281;
  wire sig00000282;
  wire sig00000283;
  wire sig00000284;
  wire sig00000285;
  wire sig00000286;
  wire sig00000287;
  wire sig00000288;
  wire sig00000289;
  wire sig0000028a;
  wire sig0000028b;
  wire sig0000028c;
  wire sig0000028d;
  wire sig0000028e;
  wire sig0000028f;
  wire sig00000290;
  wire sig00000291;
  wire sig00000292;
  wire sig00000293;
  wire sig00000294;
  wire sig00000295;
  wire sig00000296;
  wire sig00000297;
  wire sig00000298;
  wire sig00000299;
  wire sig0000029a;
  wire sig0000029b;
  wire sig0000029c;
  wire sig0000029d;
  wire sig0000029e;
  wire sig0000029f;
  wire sig000002a0;
  wire sig000002a1;
  wire sig000002a2;
  wire sig000002a3;
  wire sig000002a4;
  wire sig000002a5;
  wire sig000002a6;
  wire sig000002a7;
  wire sig000002a8;
  wire sig000002a9;
  wire sig000002aa;
  wire sig000002ab;
  wire sig000002ac;
  wire sig000002ad;
  wire sig000002ae;
  wire sig000002af;
  wire sig000002b0;
  wire sig000002b1;
  wire sig000002b2;
  wire sig000002b3;
  wire sig000002b4;
  wire sig000002b5;
  wire sig000002b6;
  wire sig000002b7;
  wire sig000002b8;
  wire sig000002b9;
  wire sig000002ba;
  wire sig000002bb;
  wire sig000002bc;
  wire sig000002bd;
  wire sig000002be;
  wire sig000002bf;
  wire sig000002c0;
  wire sig000002c1;
  wire sig000002c2;
  wire sig000002c3;
  wire sig000002c4;
  wire sig000002c5;
  wire sig000002c6;
  wire sig000002c7;
  wire sig000002c8;
  wire sig000002c9;
  wire sig000002ca;
  wire sig000002cb;
  wire sig000002cc;
  wire sig000002cd;
  wire sig000002ce;
  wire sig000002cf;
  wire sig000002d0;
  wire sig000002d1;
  wire sig000002d2;
  wire sig000002d3;
  wire sig000002d4;
  wire sig000002d5;
  wire sig000002d6;
  wire sig000002d7;
  wire sig000002d8;
  wire sig000002d9;
  wire sig000002da;
  wire sig000002db;
  wire sig000002dc;
  wire sig000002dd;
  wire sig000002de;
  wire sig000002df;
  wire sig000002e0;
  wire sig000002e1;
  wire sig000002e2;
  wire sig000002e3;
  wire sig000002e4;
  wire sig000002e5;
  wire sig000002e6;
  wire sig000002e7;
  wire sig000002e8;
  wire sig000002e9;
  wire sig000002ea;
  wire sig000002eb;
  wire sig000002ec;
  wire sig000002ed;
  wire sig000002ee;
  wire sig000002ef;
  wire sig000002f0;
  wire sig000002f1;
  wire sig000002f2;
  wire sig000002f3;
  wire sig000002f4;
  wire sig000002f5;
  wire sig000002f6;
  wire sig000002f7;
  wire sig000002f8;
  wire sig000002f9;
  wire sig000002fa;
  wire sig000002fb;
  wire sig000002fc;
  wire sig000002fd;
  wire sig000002fe;
  wire sig000002ff;
  wire sig00000300;
  wire sig00000301;
  wire sig00000302;
  wire sig00000303;
  wire sig00000304;
  wire sig00000305;
  wire sig00000306;
  wire sig00000307;
  wire sig00000308;
  wire sig00000309;
  wire sig0000030a;
  wire sig0000030b;
  wire sig0000030c;
  wire sig0000030d;
  wire sig0000030e;
  wire sig0000030f;
  wire sig00000310;
  wire sig00000311;
  wire sig00000312;
  wire sig00000313;
  wire sig00000314;
  wire sig00000315;
  wire sig00000316;
  wire sig00000317;
  wire sig00000318;
  wire sig00000319;
  wire sig0000031a;
  wire sig0000031b;
  wire sig0000031c;
  wire sig0000031d;
  wire sig0000031e;
  wire sig0000031f;
  wire sig00000320;
  wire sig00000321;
  wire sig00000322;
  wire sig00000323;
  wire sig00000324;
  wire sig00000325;
  wire sig00000326;
  wire sig00000327;
  wire sig00000328;
  wire sig00000329;
  wire sig0000032a;
  wire sig0000032b;
  wire sig0000032c;
  wire sig0000032d;
  wire sig0000032e;
  wire sig0000032f;
  wire sig00000330;
  wire sig00000331;
  wire sig00000332;
  wire sig00000333;
  wire sig00000334;
  wire sig00000335;
  wire sig00000336;
  wire sig00000337;
  wire sig00000338;
  wire sig00000339;
  wire sig0000033a;
  wire sig0000033b;
  wire sig0000033c;
  wire sig0000033d;
  wire sig0000033e;
  wire sig0000033f;
  wire sig00000340;
  wire sig00000341;
  wire sig00000342;
  wire sig00000343;
  wire sig00000344;
  wire sig00000345;
  wire sig00000346;
  wire sig00000347;
  wire sig00000348;
  wire sig00000349;
  wire sig0000034a;
  wire sig0000034b;
  wire sig0000034c;
  wire sig0000034d;
  wire sig0000034e;
  wire sig0000034f;
  wire sig00000350;
  wire sig00000351;
  wire sig00000352;
  wire sig00000353;
  wire sig00000354;
  wire sig00000355;
  wire sig00000356;
  wire sig00000357;
  wire sig00000358;
  wire sig00000359;
  wire sig0000035a;
  wire sig0000035b;
  wire sig0000035c;
  wire sig0000035d;
  wire sig0000035e;
  wire sig0000035f;
  wire sig00000360;
  wire sig00000361;
  wire sig00000362;
  wire sig00000363;
  wire sig00000364;
  wire sig00000365;
  wire sig00000366;
  wire sig00000367;
  wire sig00000368;
  wire sig00000369;
  wire sig0000036a;
  wire sig0000036b;
  wire sig0000036c;
  wire sig0000036d;
  wire sig0000036e;
  wire sig0000036f;
  wire sig00000370;
  wire sig00000371;
  wire sig00000372;
  wire sig00000373;
  wire sig00000374;
  wire sig00000375;
  wire sig00000376;
  wire sig00000377;
  wire sig00000378;
  wire sig00000379;
  wire sig0000037a;
  wire sig0000037b;
  wire sig0000037c;
  wire sig0000037d;
  wire sig0000037e;
  wire sig0000037f;
  wire sig00000380;
  wire sig00000381;
  wire sig00000382;
  wire sig00000383;
  wire sig00000384;
  wire sig00000385;
  wire sig00000386;
  wire sig00000387;
  wire sig00000388;
  wire sig00000389;
  wire sig0000038a;
  wire sig0000038b;
  wire sig0000038c;
  wire sig0000038d;
  wire sig0000038e;
  wire sig0000038f;
  wire sig00000390;
  wire sig00000391;
  wire sig00000392;
  wire sig00000393;
  wire sig00000394;
  wire sig00000395;
  wire sig00000396;
  wire sig00000397;
  wire sig00000398;
  wire sig00000399;
  wire sig0000039a;
  wire sig0000039b;
  wire sig0000039c;
  wire sig0000039d;
  wire sig0000039e;
  wire sig0000039f;
  wire sig000003a0;
  wire sig000003a1;
  wire sig000003a2;
  wire sig000003a3;
  wire sig000003a4;
  wire sig000003a5;
  wire sig000003a6;
  wire sig000003a7;
  wire sig000003a8;
  wire sig000003a9;
  wire sig000003aa;
  wire sig000003ab;
  wire sig000003ac;
  wire sig000003ad;
  wire sig000003ae;
  wire sig000003af;
  wire sig000003b0;
  wire sig000003b1;
  wire sig000003b2;
  wire sig000003b3;
  wire sig000003b4;
  wire sig000003b5;
  wire sig000003b6;
  wire sig000003b7;
  wire sig000003b8;
  wire sig000003b9;
  wire sig000003ba;
  wire sig000003bb;
  wire sig000003bc;
  wire sig000003bd;
  wire sig000003be;
  wire sig000003bf;
  wire sig000003c0;
  wire sig000003c1;
  wire sig000003c2;
  wire sig000003c3;
  wire sig000003c4;
  wire sig000003c5;
  wire sig000003c6;
  wire sig000003c7;
  wire sig000003c8;
  wire sig000003c9;
  wire sig000003ca;
  wire sig000003cb;
  wire sig000003cc;
  wire sig000003cd;
  wire sig000003ce;
  wire sig000003cf;
  wire sig000003d0;
  wire sig000003d1;
  wire sig000003d2;
  wire sig000003d3;
  wire sig000003d4;
  wire sig000003d5;
  wire sig000003d6;
  wire sig000003d7;
  wire sig000003d8;
  wire sig000003d9;
  wire sig000003da;
  wire sig000003db;
  wire sig000003dc;
  wire sig000003dd;
  wire sig000003de;
  wire sig000003df;
  wire sig000003e0;
  wire sig000003e1;
  wire sig000003e2;
  wire sig000003e3;
  wire sig000003e4;
  wire sig000003e5;
  wire sig000003e6;
  wire sig000003e7;
  wire sig000003e8;
  wire sig000003e9;
  wire sig000003ea;
  wire sig000003eb;
  wire sig000003ec;
  wire sig000003ed;
  wire sig000003ee;
  wire sig000003ef;
  wire sig000003f0;
  wire sig000003f1;
  wire sig000003f2;
  wire sig000003f3;
  wire sig000003f4;
  wire sig000003f5;
  wire sig000003f6;
  wire sig000003f7;
  wire sig000003f8;
  wire sig000003f9;
  wire sig000003fa;
  wire sig000003fb;
  wire sig000003fc;
  wire sig000003fd;
  wire sig000003fe;
  wire sig000003ff;
  wire sig00000400;
  wire sig00000401;
  wire sig00000402;
  wire sig00000403;
  wire sig00000404;
  wire sig00000405;
  wire sig00000406;
  wire sig00000407;
  wire sig00000408;
  wire sig00000409;
  wire sig0000040a;
  wire sig0000040b;
  wire sig0000040c;
  wire sig0000040d;
  wire sig0000040e;
  wire sig0000040f;
  wire sig00000410;
  wire sig00000411;
  wire sig00000412;
  wire sig00000413;
  wire sig00000414;
  wire sig00000415;
  wire sig00000416;
  wire sig00000417;
  wire sig00000418;
  wire sig00000419;
  wire sig0000041a;
  wire sig0000041b;
  wire sig0000041c;
  wire sig0000041d;
  wire sig0000041e;
  wire sig0000041f;
  wire sig00000420;
  wire sig00000421;
  wire sig00000422;
  wire sig00000423;
  wire sig00000424;
  wire sig00000425;
  wire sig00000426;
  wire sig00000427;
  wire sig00000428;
  wire sig00000429;
  wire sig0000042a;
  wire sig0000042b;
  wire sig0000042c;
  wire sig0000042d;
  wire sig0000042e;
  wire sig0000042f;
  wire sig00000430;
  wire sig00000431;
  wire sig00000432;
  wire sig00000433;
  wire sig00000434;
  wire sig00000435;
  wire sig00000436;
  wire sig00000437;
  wire sig00000438;
  wire sig00000439;
  wire sig0000043a;
  wire sig0000043b;
  wire sig0000043c;
  wire sig0000043d;
  wire sig0000043e;
  wire sig0000043f;
  wire sig00000440;
  wire sig00000441;
  wire sig00000442;
  wire sig00000443;
  wire sig00000444;
  wire sig00000445;
  wire sig00000446;
  wire sig00000447;
  wire sig00000448;
  wire sig00000449;
  wire sig0000044a;
  wire sig0000044b;
  wire sig0000044c;
  wire sig0000044d;
  wire sig0000044e;
  wire sig0000044f;
  wire sig00000450;
  wire sig00000451;
  wire sig00000452;
  wire sig00000453;
  wire sig00000454;
  wire sig00000455;
  wire sig00000456;
  wire sig00000457;
  wire sig00000458;
  wire sig00000459;
  wire sig0000045a;
  wire sig0000045b;
  wire sig0000045c;
  wire sig0000045d;
  wire sig0000045e;
  wire sig0000045f;
  wire sig00000460;
  wire sig00000461;
  wire sig00000462;
  wire sig00000463;
  wire sig00000464;
  wire sig00000465;
  wire sig00000466;
  wire sig00000467;
  wire sig00000468;
  wire sig00000469;
  wire sig0000046a;
  wire sig0000046b;
  wire sig0000046c;
  wire sig0000046d;
  wire sig0000046e;
  wire sig0000046f;
  wire sig00000470;
  wire sig00000471;
  wire sig00000472;
  wire sig00000473;
  wire sig00000474;
  wire sig00000475;
  wire sig00000476;
  wire sig00000477;
  wire sig00000478;
  wire sig00000479;
  wire sig0000047a;
  wire sig0000047b;
  wire sig0000047c;
  wire sig0000047d;
  wire sig0000047e;
  wire sig0000047f;
  wire sig00000480;
  wire sig00000481;
  wire sig00000482;
  wire sig00000483;
  wire sig00000484;
  wire sig00000485;
  wire sig00000486;
  wire sig00000487;
  wire sig00000488;
  wire sig00000489;
  wire sig0000048a;
  wire sig0000048b;
  wire sig0000048c;
  wire sig0000048d;
  wire sig0000048e;
  wire sig0000048f;
  wire sig00000490;
  wire sig00000491;
  wire sig00000492;
  wire sig00000493;
  wire sig00000494;
  wire sig00000495;
  wire sig00000496;
  wire sig00000497;
  wire sig00000498;
  wire sig00000499;
  wire sig0000049a;
  wire sig0000049b;
  wire sig0000049c;
  wire sig0000049d;
  wire sig0000049e;
  wire sig0000049f;
  wire sig000004a0;
  wire sig000004a1;
  wire sig000004a2;
  wire sig000004a3;
  wire sig000004a4;
  wire sig000004a5;
  wire sig000004a6;
  wire sig000004a7;
  wire sig000004a8;
  wire sig000004a9;
  wire sig000004aa;
  wire sig000004ab;
  wire sig000004ac;
  wire sig000004ad;
  wire sig000004ae;
  wire sig000004af;
  wire sig000004b0;
  wire sig000004b1;
  wire sig000004b2;
  wire sig000004b3;
  wire sig000004b4;
  wire sig000004b5;
  wire sig000004b6;
  wire sig000004b7;
  wire sig000004b8;
  wire sig000004b9;
  wire sig000004ba;
  wire sig000004bb;
  wire sig000004bc;
  wire sig000004bd;
  wire sig000004be;
  wire sig000004bf;
  wire sig000004c0;
  wire sig000004c1;
  wire sig000004c2;
  wire sig000004c3;
  wire sig000004c4;
  wire sig000004c5;
  wire sig000004c6;
  wire sig000004c7;
  wire sig000004c8;
  wire sig000004c9;
  wire sig000004ca;
  wire sig000004cb;
  wire sig000004cc;
  wire sig000004cd;
  wire sig000004ce;
  wire sig000004cf;
  wire sig000004d0;
  wire sig000004d1;
  wire sig000004d2;
  wire sig000004d3;
  wire sig000004d4;
  wire sig000004d5;
  wire sig000004d6;
  wire sig000004d7;
  wire sig000004d8;
  wire sig000004d9;
  wire sig000004da;
  wire sig000004db;
  wire sig000004dc;
  wire sig000004dd;
  wire sig000004de;
  wire sig000004df;
  wire sig000004e0;
  wire sig000004e1;
  wire sig000004e2;
  wire sig000004e3;
  wire sig000004e4;
  wire sig000004e5;
  wire sig000004e6;
  wire sig000004e7;
  wire sig000004e8;
  wire sig000004e9;
  wire sig000004ea;
  wire sig000004eb;
  wire sig000004ec;
  wire sig000004ed;
  wire sig000004ee;
  wire sig000004ef;
  wire sig000004f0;
  wire sig000004f1;
  wire sig000004f2;
  wire sig000004f3;
  wire sig000004f4;
  wire sig000004f5;
  wire sig000004f6;
  wire sig000004f7;
  wire sig000004f8;
  wire sig000004f9;
  wire sig000004fa;
  wire sig000004fb;
  wire sig000004fc;
  wire sig000004fd;
  wire sig000004fe;
  wire sig000004ff;
  wire sig00000500;
  wire sig00000501;
  wire sig00000502;
  wire sig00000503;
  wire sig00000504;
  wire sig00000505;
  wire sig00000506;
  wire sig00000507;
  wire sig00000508;
  wire sig00000509;
  wire sig0000050a;
  wire sig0000050b;
  wire sig0000050c;
  wire sig0000050d;
  wire sig0000050e;
  wire sig0000050f;
  wire sig00000510;
  wire sig00000511;
  wire sig00000512;
  wire sig00000513;
  wire sig00000514;
  wire sig00000515;
  wire sig00000516;
  wire sig00000517;
  wire sig00000518;
  wire sig00000519;
  wire sig0000051a;
  wire sig0000051b;
  wire sig0000051c;
  wire sig0000051d;
  wire sig0000051e;
  wire sig0000051f;
  wire sig00000520;
  wire sig00000521;
  wire sig00000522;
  wire sig00000523;
  wire sig00000524;
  wire sig00000525;
  wire sig00000526;
  wire sig00000527;
  wire sig00000528;
  wire sig00000529;
  wire sig0000052a;
  wire sig0000052b;
  wire sig0000052c;
  wire sig0000052d;
  wire sig0000052e;
  wire sig0000052f;
  wire sig00000530;
  wire sig00000531;
  wire sig00000532;
  wire sig00000533;
  wire sig00000534;
  wire sig00000535;
  wire sig00000536;
  wire sig00000537;
  wire sig00000538;
  wire sig00000539;
  wire sig0000053a;
  wire sig0000053b;
  wire sig0000053c;
  wire sig0000053d;
  wire sig0000053e;
  wire sig0000053f;
  wire sig00000540;
  wire sig00000541;
  wire sig00000542;
  wire sig00000543;
  wire sig00000544;
  wire sig00000545;
  wire sig00000546;
  wire sig00000547;
  wire sig00000548;
  wire sig00000549;
  wire sig0000054a;
  wire sig0000054b;
  wire sig0000054c;
  wire sig0000054d;
  wire sig0000054e;
  wire sig0000054f;
  wire sig00000550;
  wire sig00000551;
  wire sig00000552;
  wire sig00000553;
  wire sig00000554;
  wire sig00000555;
  wire sig00000556;
  wire sig00000557;
  wire sig00000558;
  wire sig00000559;
  wire sig0000055a;
  wire sig0000055b;
  wire sig0000055c;
  wire sig0000055d;
  wire sig0000055e;
  wire sig0000055f;
  wire sig00000560;
  wire sig00000561;
  wire sig00000562;
  wire sig00000563;
  wire sig00000564;
  wire sig00000565;
  wire sig00000566;
  wire sig00000567;
  wire sig00000568;
  wire sig00000569;
  wire sig0000056a;
  wire sig0000056b;
  wire sig0000056c;
  wire sig0000056d;
  wire sig0000056e;
  wire sig0000056f;
  wire sig00000570;
  wire sig00000571;
  wire sig00000572;
  wire sig00000573;
  wire sig00000574;
  wire sig00000575;
  wire sig00000576;
  wire sig00000577;
  wire sig00000578;
  wire sig00000579;
  wire sig0000057a;
  wire sig0000057b;
  wire sig0000057c;
  wire sig0000057d;
  wire sig0000057e;
  wire sig0000057f;
  wire sig00000580;
  wire sig00000581;
  wire sig00000582;
  wire sig00000583;
  wire sig00000584;
  wire sig00000585;
  wire sig00000586;
  wire sig00000587;
  wire sig00000588;
  wire sig00000589;
  wire sig0000058a;
  wire sig0000058b;
  wire sig0000058c;
  wire sig0000058d;
  wire sig0000058e;
  wire sig0000058f;
  wire sig00000590;
  wire sig00000591;
  wire sig00000592;
  wire sig00000593;
  wire sig00000594;
  wire sig00000595;
  wire sig00000596;
  wire sig00000597;
  wire sig00000598;
  wire sig00000599;
  wire sig0000059a;
  wire sig0000059b;
  wire sig0000059c;
  wire sig0000059d;
  wire sig0000059e;
  wire sig0000059f;
  wire sig000005a0;
  wire \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/sign_op ;
  wire sig000005a1;
  wire sig000005a2;
  wire sig000005a3;
  wire NLW_blk0000020d_O_UNCONNECTED;
  wire NLW_blk0000020e_O_UNCONNECTED;
  wire NLW_blk00000210_O_UNCONNECTED;
  wire NLW_blk00000212_O_UNCONNECTED;
  wire NLW_blk00000214_O_UNCONNECTED;
  wire NLW_blk00000216_O_UNCONNECTED;
  wire NLW_blk00000218_O_UNCONNECTED;
  wire NLW_blk0000021a_O_UNCONNECTED;
  wire NLW_blk0000027a_O_UNCONNECTED;
  wire [7 : 0] \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/exp_op ;
  wire [22 : 0] \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op ;
  assign
    result[31] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/sign_op ,
    result[30] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/exp_op [7],
    result[29] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/exp_op [6],
    result[28] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/exp_op [5],
    result[27] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/exp_op [4],
    result[26] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/exp_op [3],
    result[25] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/exp_op [2],
    result[24] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/exp_op [1],
    result[23] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/exp_op [0],
    result[22] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [22],
    result[21] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [21],
    result[20] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [20],
    result[19] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [19],
    result[18] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [18],
    result[17] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [17],
    result[16] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [16],
    result[15] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [15],
    result[14] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [14],
    result[13] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [13],
    result[12] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [12],
    result[11] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [11],
    result[10] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [10],
    result[9] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [9],
    result[8] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [8],
    result[7] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [7],
    result[6] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [6],
    result[5] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [5],
    result[4] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [4],
    result[3] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [3],
    result[2] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [2],
    result[1] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [1],
    result[0] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [0];
  GND   blk00000001 (
    .G(sig00000001)
  );
  VCC   blk00000002 (
    .P(sig00000002)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000003 (
    .C(clk),
    .CE(ce),
    .D(sig00000148),
    .Q(sig0000025d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000004 (
    .C(clk),
    .CE(ce),
    .D(sig0000025c),
    .Q(sig0000025b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000005 (
    .C(clk),
    .CE(ce),
    .D(sig000002a0),
    .Q(sig0000025c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000006 (
    .C(clk),
    .CE(ce),
    .D(sig000005a3),
    .Q(sig0000025f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000007 (
    .C(clk),
    .CE(ce),
    .D(sig000002a1),
    .Q(sig00000261)
  );
  MUXCY   blk00000008 (
    .CI(sig00000001),
    .DI(sig000002e1),
    .S(sig0000023a),
    .O(sig00000239)
  );
  XORCY   blk00000009 (
    .CI(sig00000001),
    .LI(sig0000023a),
    .O(sig00000269)
  );
  MUXCY   blk0000000a (
    .CI(sig00000239),
    .DI(sig00000001),
    .S(sig00000262),
    .O(sig0000023b)
  );
  XORCY   blk0000000b (
    .CI(sig00000239),
    .LI(sig00000262),
    .O(sig0000026a)
  );
  MUXCY   blk0000000c (
    .CI(sig0000023b),
    .DI(sig00000001),
    .S(sig00000263),
    .O(sig0000023c)
  );
  XORCY   blk0000000d (
    .CI(sig0000023b),
    .LI(sig00000263),
    .O(sig0000026b)
  );
  MUXCY   blk0000000e (
    .CI(sig0000023c),
    .DI(sig00000001),
    .S(sig00000264),
    .O(sig0000023d)
  );
  XORCY   blk0000000f (
    .CI(sig0000023c),
    .LI(sig00000264),
    .O(sig0000026c)
  );
  MUXCY   blk00000010 (
    .CI(sig0000023d),
    .DI(sig00000001),
    .S(sig00000265),
    .O(sig0000023e)
  );
  XORCY   blk00000011 (
    .CI(sig0000023d),
    .LI(sig00000265),
    .O(sig0000026d)
  );
  MUXCY   blk00000012 (
    .CI(sig0000023e),
    .DI(sig00000001),
    .S(sig00000266),
    .O(sig0000023f)
  );
  XORCY   blk00000013 (
    .CI(sig0000023e),
    .LI(sig00000266),
    .O(sig0000026e)
  );
  MUXCY   blk00000014 (
    .CI(sig0000023f),
    .DI(sig00000001),
    .S(sig00000267),
    .O(sig00000240)
  );
  XORCY   blk00000015 (
    .CI(sig0000023f),
    .LI(sig00000267),
    .O(sig0000026f)
  );
  XORCY   blk00000016 (
    .CI(sig00000240),
    .LI(sig00000268),
    .O(sig00000270)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000017 (
    .C(clk),
    .CE(ce),
    .D(sig00000002),
    .Q(sig00000251)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000018 (
    .C(clk),
    .CE(ce),
    .D(sig00000297),
    .Q(sig00000250)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000019 (
    .C(clk),
    .CE(ce),
    .D(sig00000296),
    .Q(sig0000024f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000001a (
    .C(clk),
    .CE(ce),
    .D(sig00000295),
    .Q(sig0000024e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000001b (
    .C(clk),
    .CE(ce),
    .D(sig00000293),
    .Q(sig0000024c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000001c (
    .C(clk),
    .CE(ce),
    .D(sig00000292),
    .Q(sig0000024b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000001d (
    .C(clk),
    .CE(ce),
    .D(sig00000291),
    .Q(sig0000024a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000001e (
    .C(clk),
    .CE(ce),
    .D(sig00000290),
    .Q(sig00000249)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000001f (
    .C(clk),
    .CE(ce),
    .D(sig0000028f),
    .Q(sig00000248)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000020 (
    .C(clk),
    .CE(ce),
    .D(sig0000028e),
    .Q(sig00000247)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000021 (
    .C(clk),
    .CE(ce),
    .D(sig0000028d),
    .Q(sig00000246)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000022 (
    .C(clk),
    .CE(ce),
    .D(sig0000028c),
    .Q(sig00000245)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000023 (
    .C(clk),
    .CE(ce),
    .D(sig0000028b),
    .Q(sig00000244)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000024 (
    .C(clk),
    .CE(ce),
    .D(sig0000028a),
    .Q(sig00000243)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000025 (
    .C(clk),
    .CE(ce),
    .D(sig0000029f),
    .Q(sig00000258)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000026 (
    .C(clk),
    .CE(ce),
    .D(sig0000029e),
    .Q(sig00000257)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000027 (
    .C(clk),
    .CE(ce),
    .D(sig0000029d),
    .Q(sig00000256)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000028 (
    .C(clk),
    .CE(ce),
    .D(sig0000029c),
    .Q(sig00000255)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000029 (
    .C(clk),
    .CE(ce),
    .D(sig0000029b),
    .Q(sig00000254)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000002a (
    .C(clk),
    .CE(ce),
    .D(sig0000029a),
    .Q(sig00000253)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000002b (
    .C(clk),
    .CE(ce),
    .D(sig00000299),
    .Q(sig00000252)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000002c (
    .C(clk),
    .CE(ce),
    .D(sig00000298),
    .Q(sig0000024d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000002d (
    .C(clk),
    .CE(ce),
    .D(sig00000294),
    .Q(sig00000242)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000002e (
    .C(clk),
    .CE(ce),
    .D(sig00000289),
    .Q(sig00000241)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000002f (
    .C(clk),
    .CE(ce),
    .D(sig00000270),
    .Q(sig0000008e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000030 (
    .C(clk),
    .CE(ce),
    .D(sig0000026f),
    .Q(sig0000008d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000031 (
    .C(clk),
    .CE(ce),
    .D(sig0000026e),
    .Q(sig0000008c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000032 (
    .C(clk),
    .CE(ce),
    .D(sig0000026d),
    .Q(sig0000008b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000033 (
    .C(clk),
    .CE(ce),
    .D(sig0000026c),
    .Q(sig0000008a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000034 (
    .C(clk),
    .CE(ce),
    .D(sig0000026b),
    .Q(sig00000089)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000035 (
    .C(clk),
    .CE(ce),
    .D(sig0000026a),
    .Q(sig00000088)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000036 (
    .C(clk),
    .CE(ce),
    .D(sig00000269),
    .Q(sig00000087)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000037 (
    .C(clk),
    .CE(ce),
    .D(sig00000117),
    .Q(sig0000008f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000038 (
    .C(clk),
    .CE(ce),
    .D(sig00000122),
    .Q(sig00000090)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000039 (
    .C(clk),
    .CE(ce),
    .D(sig00000129),
    .Q(sig0000009b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000003a (
    .C(clk),
    .CE(ce),
    .D(sig0000012a),
    .Q(sig000000a2)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000003b (
    .C(clk),
    .CE(ce),
    .D(sig0000012b),
    .Q(sig000000a3)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000003c (
    .C(clk),
    .CE(ce),
    .D(sig0000012c),
    .Q(sig000000a4)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000003d (
    .C(clk),
    .CE(ce),
    .D(sig0000012d),
    .Q(sig000000a5)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000003e (
    .C(clk),
    .CE(ce),
    .D(sig0000012e),
    .Q(sig000000a6)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000003f (
    .C(clk),
    .CE(ce),
    .D(sig0000012f),
    .Q(sig000000a7)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000040 (
    .C(clk),
    .CE(ce),
    .D(sig00000130),
    .Q(sig000000a8)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000041 (
    .C(clk),
    .CE(ce),
    .D(sig00000118),
    .Q(sig00000091)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000042 (
    .C(clk),
    .CE(ce),
    .D(sig00000119),
    .Q(sig00000092)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000043 (
    .C(clk),
    .CE(ce),
    .D(sig0000011a),
    .Q(sig00000093)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000044 (
    .C(clk),
    .CE(ce),
    .D(sig0000011b),
    .Q(sig00000094)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000045 (
    .C(clk),
    .CE(ce),
    .D(sig0000011c),
    .Q(sig00000095)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000046 (
    .C(clk),
    .CE(ce),
    .D(sig0000011d),
    .Q(sig00000096)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000047 (
    .C(clk),
    .CE(ce),
    .D(sig0000011e),
    .Q(sig00000097)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000048 (
    .C(clk),
    .CE(ce),
    .D(sig0000011f),
    .Q(sig00000098)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000049 (
    .C(clk),
    .CE(ce),
    .D(sig00000120),
    .Q(sig00000099)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000004a (
    .C(clk),
    .CE(ce),
    .D(sig00000121),
    .Q(sig0000009a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000004b (
    .C(clk),
    .CE(ce),
    .D(sig00000123),
    .Q(sig0000009c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000004c (
    .C(clk),
    .CE(ce),
    .D(sig00000124),
    .Q(sig0000009d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000004d (
    .C(clk),
    .CE(ce),
    .D(sig00000125),
    .Q(sig0000009e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000004e (
    .C(clk),
    .CE(ce),
    .D(sig00000126),
    .Q(sig0000009f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000004f (
    .C(clk),
    .CE(ce),
    .D(sig00000127),
    .Q(sig000000a0)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000050 (
    .C(clk),
    .CE(ce),
    .D(sig00000128),
    .Q(sig000000a1)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000051 (
    .C(clk),
    .CE(ce),
    .D(sig000000fd),
    .Q(sig000000a9)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000052 (
    .C(clk),
    .CE(ce),
    .D(sig00000108),
    .Q(sig000000aa)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000053 (
    .C(clk),
    .CE(ce),
    .D(sig0000010f),
    .Q(sig000000b5)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000054 (
    .C(clk),
    .CE(ce),
    .D(sig00000110),
    .Q(sig000000bc)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000055 (
    .C(clk),
    .CE(ce),
    .D(sig00000111),
    .Q(sig000000bd)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000056 (
    .C(clk),
    .CE(ce),
    .D(sig00000112),
    .Q(sig000000be)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000057 (
    .C(clk),
    .CE(ce),
    .D(sig00000113),
    .Q(sig000000bf)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000058 (
    .C(clk),
    .CE(ce),
    .D(sig00000114),
    .Q(sig000000c0)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000059 (
    .C(clk),
    .CE(ce),
    .D(sig00000115),
    .Q(sig000000c1)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000005a (
    .C(clk),
    .CE(ce),
    .D(sig00000116),
    .Q(sig000000c2)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000005b (
    .C(clk),
    .CE(ce),
    .D(sig000000fe),
    .Q(sig000000ab)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000005c (
    .C(clk),
    .CE(ce),
    .D(sig000000ff),
    .Q(sig000000ac)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000005d (
    .C(clk),
    .CE(ce),
    .D(sig00000100),
    .Q(sig000000ad)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000005e (
    .C(clk),
    .CE(ce),
    .D(sig00000101),
    .Q(sig000000ae)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000005f (
    .C(clk),
    .CE(ce),
    .D(sig00000102),
    .Q(sig000000af)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000060 (
    .C(clk),
    .CE(ce),
    .D(sig00000103),
    .Q(sig000000b0)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000061 (
    .C(clk),
    .CE(ce),
    .D(sig00000104),
    .Q(sig000000b1)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000062 (
    .C(clk),
    .CE(ce),
    .D(sig00000105),
    .Q(sig000000b2)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000063 (
    .C(clk),
    .CE(ce),
    .D(sig00000106),
    .Q(sig000000b3)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000064 (
    .C(clk),
    .CE(ce),
    .D(sig00000107),
    .Q(sig000000b4)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000065 (
    .C(clk),
    .CE(ce),
    .D(sig00000109),
    .Q(sig000000b6)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000066 (
    .C(clk),
    .CE(ce),
    .D(sig0000010a),
    .Q(sig000000b7)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000067 (
    .C(clk),
    .CE(ce),
    .D(sig0000010b),
    .Q(sig000000b8)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000068 (
    .C(clk),
    .CE(ce),
    .D(sig0000010c),
    .Q(sig000000b9)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000069 (
    .C(clk),
    .CE(ce),
    .D(sig0000010d),
    .Q(sig000000ba)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000006a (
    .C(clk),
    .CE(ce),
    .D(sig0000010e),
    .Q(sig000000bb)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000006b (
    .C(clk),
    .CE(ce),
    .D(sig000000e3),
    .Q(sig000000c5)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000006c (
    .C(clk),
    .CE(ce),
    .D(sig000000e4),
    .Q(sig000000c6)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000006d (
    .C(clk),
    .CE(ce),
    .D(sig000000ef),
    .Q(sig000000d1)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000006e (
    .C(clk),
    .CE(ce),
    .D(sig000000f6),
    .Q(sig000000d8)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000006f (
    .C(clk),
    .CE(ce),
    .D(sig000000f7),
    .Q(sig000000d9)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000070 (
    .C(clk),
    .CE(ce),
    .D(sig000000f8),
    .Q(sig000000da)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000071 (
    .C(clk),
    .CE(ce),
    .D(sig000000f9),
    .Q(sig000000db)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000072 (
    .C(clk),
    .CE(ce),
    .D(sig000000fa),
    .Q(sig000000dc)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000073 (
    .C(clk),
    .CE(ce),
    .D(sig000000fb),
    .Q(sig000000dd)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000074 (
    .C(clk),
    .CE(ce),
    .D(sig000000fc),
    .Q(sig000000de)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000075 (
    .C(clk),
    .CE(ce),
    .D(sig000000e5),
    .Q(sig000000c7)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000076 (
    .C(clk),
    .CE(ce),
    .D(sig000000e6),
    .Q(sig000000c8)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000077 (
    .C(clk),
    .CE(ce),
    .D(sig000000e7),
    .Q(sig000000c9)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000078 (
    .C(clk),
    .CE(ce),
    .D(sig000000e8),
    .Q(sig000000ca)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000079 (
    .C(clk),
    .CE(ce),
    .D(sig000000e9),
    .Q(sig000000cb)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000007a (
    .C(clk),
    .CE(ce),
    .D(sig000000ea),
    .Q(sig000000cc)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000007b (
    .C(clk),
    .CE(ce),
    .D(sig000000eb),
    .Q(sig000000cd)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000007c (
    .C(clk),
    .CE(ce),
    .D(sig000000ec),
    .Q(sig000000ce)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000007d (
    .C(clk),
    .CE(ce),
    .D(sig000000ed),
    .Q(sig000000cf)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000007e (
    .C(clk),
    .CE(ce),
    .D(sig000000ee),
    .Q(sig000000d0)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000007f (
    .C(clk),
    .CE(ce),
    .D(sig000000f0),
    .Q(sig000000d2)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000080 (
    .C(clk),
    .CE(ce),
    .D(sig000000f1),
    .Q(sig000000d3)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000081 (
    .C(clk),
    .CE(ce),
    .D(sig000000f2),
    .Q(sig000000d4)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000082 (
    .C(clk),
    .CE(ce),
    .D(sig000000f3),
    .Q(sig000000d5)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000083 (
    .C(clk),
    .CE(ce),
    .D(sig000000f4),
    .Q(sig000000d6)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000084 (
    .C(clk),
    .CE(ce),
    .D(sig000000f5),
    .Q(sig000000d7)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000085 (
    .C(clk),
    .CE(ce),
    .D(sig00000089),
    .Q(sig000000c3)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000086 (
    .C(clk),
    .CE(ce),
    .D(sig0000008a),
    .Q(sig000000c4)
  );
  MUXCY   blk00000087 (
    .CI(sig00000136),
    .DI(sig00000001),
    .S(sig0000013e),
    .O(sig00000137)
  );
  MUXCY   blk00000088 (
    .CI(sig00000135),
    .DI(sig00000001),
    .S(sig0000013d),
    .O(sig00000136)
  );
  MUXCY   blk00000089 (
    .CI(sig00000134),
    .DI(sig00000001),
    .S(sig0000013c),
    .O(sig00000135)
  );
  MUXCY   blk0000008a (
    .CI(sig00000133),
    .DI(sig00000001),
    .S(sig0000013b),
    .O(sig00000134)
  );
  MUXCY   blk0000008b (
    .CI(sig00000132),
    .DI(sig00000001),
    .S(sig0000013a),
    .O(sig00000133)
  );
  MUXCY   blk0000008c (
    .CI(sig00000131),
    .DI(sig00000001),
    .S(sig00000139),
    .O(sig00000132)
  );
  MUXCY   blk0000008d (
    .CI(sig00000002),
    .DI(sig00000001),
    .S(sig00000138),
    .O(sig00000131)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000008e (
    .C(clk),
    .CE(ce),
    .D(sig00000137),
    .Q(sig0000015a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000008f (
    .C(clk),
    .CE(ce),
    .D(sig00000136),
    .Q(sig00000159)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000090 (
    .C(clk),
    .CE(ce),
    .D(sig00000135),
    .Q(sig00000158)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000091 (
    .C(clk),
    .CE(ce),
    .D(sig00000134),
    .Q(sig00000157)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000092 (
    .C(clk),
    .CE(ce),
    .D(sig00000133),
    .Q(sig00000156)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000093 (
    .C(clk),
    .CE(ce),
    .D(sig00000132),
    .Q(sig00000155)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000094 (
    .C(clk),
    .CE(ce),
    .D(sig00000131),
    .Q(sig00000154)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000095 (
    .C(clk),
    .CE(ce),
    .D(sig0000015b),
    .Q(sig0000013f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000096 (
    .C(clk),
    .CE(ce),
    .D(sig0000015c),
    .Q(sig00000140)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000097 (
    .C(clk),
    .CE(ce),
    .D(sig0000015d),
    .Q(sig00000141)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000098 (
    .C(clk),
    .CE(ce),
    .D(sig0000015e),
    .Q(sig00000142)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000099 (
    .C(clk),
    .CE(ce),
    .D(sig0000015f),
    .Q(sig00000143)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000009a (
    .C(clk),
    .CE(ce),
    .D(sig00000160),
    .Q(sig00000144)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000009b (
    .C(clk),
    .CE(ce),
    .D(sig00000161),
    .Q(sig00000145)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000009c (
    .C(clk),
    .CE(ce),
    .D(sig00000162),
    .Q(sig00000146)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000009d (
    .C(clk),
    .CE(ce),
    .D(sig00000163),
    .Q(sig00000147)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000009e (
    .C(clk),
    .CE(ce),
    .D(sig00000164),
    .Q(sig00000148)
  );
  MUXF7   blk0000009f (
    .I0(sig00000152),
    .I1(sig00000153),
    .S(sig00000001),
    .O(sig00000164)
  );
  MUXF6   blk000000a0 (
    .I0(sig00000251),
    .I1(sig00000251),
    .S(sig0000014a),
    .O(sig00000153)
  );
  MUXF6   blk000000a1 (
    .I0(sig00000146),
    .I1(sig00000147),
    .S(sig0000014a),
    .O(sig00000152)
  );
  MUXF5   blk000000a2 (
    .I0(sig0000014c),
    .I1(sig0000014b),
    .S(sig000000c4),
    .O(sig00000162)
  );
  MUXF5   blk000000a3 (
    .I0(sig0000014e),
    .I1(sig0000014d),
    .S(sig000000c4),
    .O(sig00000163)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000a4 (
    .C(clk),
    .CE(ce),
    .D(sig000001e1),
    .Q(sig00000210)
  );
  MUXCY   blk000000a5 (
    .CI(sig0000020f),
    .DI(sig00000001),
    .S(sig00000211),
    .O(sig000001d8)
  );
  XORCY   blk000000a6 (
    .CI(sig0000020f),
    .LI(sig00000211),
    .O(sig000001e2)
  );
  MUXCY   blk000000a7 (
    .CI(sig000001d8),
    .DI(sig00000001),
    .S(sig00000212),
    .O(sig000001d9)
  );
  XORCY   blk000000a8 (
    .CI(sig000001d8),
    .LI(sig00000212),
    .O(sig000001e6)
  );
  MUXCY   blk000000a9 (
    .CI(sig000001d9),
    .DI(sig00000197),
    .S(sig00000225),
    .O(sig000001da)
  );
  XORCY   blk000000aa (
    .CI(sig000001d9),
    .LI(sig00000225),
    .O(sig000001e7)
  );
  MUXCY   blk000000ab (
    .CI(sig000001da),
    .DI(sig00000198),
    .S(sig00000226),
    .O(sig000001db)
  );
  XORCY   blk000000ac (
    .CI(sig000001da),
    .LI(sig00000226),
    .O(sig000001e8)
  );
  MUXCY   blk000000ad (
    .CI(sig000001db),
    .DI(sig0000019a),
    .S(sig00000227),
    .O(sig000001dc)
  );
  XORCY   blk000000ae (
    .CI(sig000001db),
    .LI(sig00000227),
    .O(sig000001e9)
  );
  MUXCY   blk000000af (
    .CI(sig000001dc),
    .DI(sig0000019b),
    .S(sig00000228),
    .O(sig000001dd)
  );
  XORCY   blk000000b0 (
    .CI(sig000001dc),
    .LI(sig00000228),
    .O(sig000001ea)
  );
  MUXCY   blk000000b1 (
    .CI(sig000001dd),
    .DI(sig0000019c),
    .S(sig00000229),
    .O(sig000001de)
  );
  XORCY   blk000000b2 (
    .CI(sig000001dd),
    .LI(sig00000229),
    .O(sig000001eb)
  );
  MUXCY   blk000000b3 (
    .CI(sig000001de),
    .DI(sig0000019d),
    .S(sig0000022a),
    .O(sig000001df)
  );
  XORCY   blk000000b4 (
    .CI(sig000001de),
    .LI(sig0000022a),
    .O(sig000001ec)
  );
  MUXCY   blk000000b5 (
    .CI(sig000001df),
    .DI(sig0000019e),
    .S(sig0000022b),
    .O(sig000001e0)
  );
  XORCY   blk000000b6 (
    .CI(sig000001df),
    .LI(sig0000022b),
    .O(sig000001ed)
  );
  MUXCY   blk000000b7 (
    .CI(sig000001e0),
    .DI(sig0000019f),
    .S(sig00000221),
    .O(sig000001d4)
  );
  XORCY   blk000000b8 (
    .CI(sig000001e0),
    .LI(sig00000221),
    .O(sig000001ee)
  );
  MUXCY   blk000000b9 (
    .CI(sig000001d4),
    .DI(sig000001a0),
    .S(sig00000222),
    .O(sig000001d5)
  );
  XORCY   blk000000ba (
    .CI(sig000001d4),
    .LI(sig00000222),
    .O(sig000001e3)
  );
  MUXCY   blk000000bb (
    .CI(sig000001d5),
    .DI(sig000001a1),
    .S(sig00000223),
    .O(sig000001d6)
  );
  XORCY   blk000000bc (
    .CI(sig000001d5),
    .LI(sig00000223),
    .O(sig000001e4)
  );
  MUXCY   blk000000bd (
    .CI(sig000001d6),
    .DI(sig00000199),
    .S(sig00000224),
    .O(sig000001d7)
  );
  XORCY   blk000000be (
    .CI(sig000001d6),
    .LI(sig00000224),
    .O(sig000001e5)
  );
  XORCY   blk000000bf (
    .CI(sig000001d7),
    .LI(sig00000001),
    .O(sig000001e1)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000c0 (
    .C(clk),
    .CE(ce),
    .D(sig000001cb),
    .Q(sig000001be)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000c1 (
    .C(clk),
    .CE(ce),
    .D(sig000001ca),
    .Q(sig000001bd)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000c2 (
    .C(clk),
    .CE(ce),
    .D(sig000001c9),
    .Q(sig000001bc)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000c3 (
    .C(clk),
    .CE(ce),
    .D(sig000001d3),
    .Q(sig000001c6)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000c4 (
    .C(clk),
    .CE(ce),
    .D(sig000001d2),
    .Q(sig000001c5)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000c5 (
    .C(clk),
    .CE(ce),
    .D(sig000001d1),
    .Q(sig000001c4)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000c6 (
    .C(clk),
    .CE(ce),
    .D(sig000001d0),
    .Q(sig000001c3)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000c7 (
    .C(clk),
    .CE(ce),
    .D(sig000001cf),
    .Q(sig000001c2)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000c8 (
    .C(clk),
    .CE(ce),
    .D(sig000001ce),
    .Q(sig000001c1)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000c9 (
    .C(clk),
    .CE(ce),
    .D(sig000001cd),
    .Q(sig000001c0)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000ca (
    .C(clk),
    .CE(ce),
    .D(sig000001cc),
    .Q(sig000001bf)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000cb (
    .C(clk),
    .CE(ce),
    .D(sig000001c8),
    .Q(sig000001bb)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000cc (
    .C(clk),
    .CE(ce),
    .D(sig000001c7),
    .Q(sig000001ba)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000cd (
    .C(clk),
    .CE(ce),
    .D(sig000001e5),
    .Q(sig000001cb)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000ce (
    .C(clk),
    .CE(ce),
    .D(sig000001e4),
    .Q(sig000001ca)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000cf (
    .C(clk),
    .CE(ce),
    .D(sig000001e3),
    .Q(sig000001c9)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000d0 (
    .C(clk),
    .CE(ce),
    .D(sig000001ee),
    .Q(sig000001d3)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000d1 (
    .C(clk),
    .CE(ce),
    .D(sig000001ed),
    .Q(sig000001d2)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000d2 (
    .C(clk),
    .CE(ce),
    .D(sig000001ec),
    .Q(sig000001d1)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000d3 (
    .C(clk),
    .CE(ce),
    .D(sig000001eb),
    .Q(sig000001d0)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000d4 (
    .C(clk),
    .CE(ce),
    .D(sig000001ea),
    .Q(sig000001cf)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000d5 (
    .C(clk),
    .CE(ce),
    .D(sig000001e9),
    .Q(sig000001ce)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000d6 (
    .C(clk),
    .CE(ce),
    .D(sig000001e8),
    .Q(sig000001cd)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000d7 (
    .C(clk),
    .CE(ce),
    .D(sig000001e7),
    .Q(sig000001cc)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000d8 (
    .C(clk),
    .CE(ce),
    .D(sig000001e6),
    .Q(sig000001c8)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000d9 (
    .C(clk),
    .CE(ce),
    .D(sig000001e2),
    .Q(sig000001c7)
  );
  MUXCY   blk000000da (
    .CI(sig00000210),
    .DI(sig0000017f),
    .S(sig0000022c),
    .O(sig000001f5)
  );
  XORCY   blk000000db (
    .CI(sig00000210),
    .LI(sig0000022c),
    .O(sig00000213)
  );
  MUXCY   blk000000dc (
    .CI(sig000001f5),
    .DI(sig00000180),
    .S(sig00000230),
    .O(sig000001f6)
  );
  XORCY   blk000000dd (
    .CI(sig000001f5),
    .LI(sig00000230),
    .O(sig00000218)
  );
  MUXCY   blk000000de (
    .CI(sig000001f6),
    .DI(sig00000184),
    .S(sig00000231),
    .O(sig000001f7)
  );
  XORCY   blk000000df (
    .CI(sig000001f6),
    .LI(sig00000231),
    .O(sig00000219)
  );
  MUXCY   blk000000e0 (
    .CI(sig000001f7),
    .DI(sig00000185),
    .S(sig00000232),
    .O(sig000001f8)
  );
  XORCY   blk000000e1 (
    .CI(sig000001f7),
    .LI(sig00000232),
    .O(sig0000021a)
  );
  MUXCY   blk000000e2 (
    .CI(sig000001f8),
    .DI(sig00000186),
    .S(sig00000233),
    .O(sig000001f9)
  );
  XORCY   blk000000e3 (
    .CI(sig000001f8),
    .LI(sig00000233),
    .O(sig0000021b)
  );
  MUXCY   blk000000e4 (
    .CI(sig000001f9),
    .DI(sig00000187),
    .S(sig00000234),
    .O(sig000001fa)
  );
  XORCY   blk000000e5 (
    .CI(sig000001f9),
    .LI(sig00000234),
    .O(sig0000021c)
  );
  MUXCY   blk000000e6 (
    .CI(sig000001fa),
    .DI(sig00000188),
    .S(sig00000235),
    .O(sig000001fb)
  );
  XORCY   blk000000e7 (
    .CI(sig000001fa),
    .LI(sig00000235),
    .O(sig0000021d)
  );
  MUXCY   blk000000e8 (
    .CI(sig000001fb),
    .DI(sig00000189),
    .S(sig00000236),
    .O(sig000001fc)
  );
  XORCY   blk000000e9 (
    .CI(sig000001fb),
    .LI(sig00000236),
    .O(sig0000021e)
  );
  MUXCY   blk000000ea (
    .CI(sig000001fc),
    .DI(sig0000018a),
    .S(sig00000237),
    .O(sig000001fd)
  );
  XORCY   blk000000eb (
    .CI(sig000001fc),
    .LI(sig00000237),
    .O(sig0000021f)
  );
  MUXCY   blk000000ec (
    .CI(sig000001fd),
    .DI(sig0000018b),
    .S(sig00000238),
    .O(sig000001f1)
  );
  XORCY   blk000000ed (
    .CI(sig000001fd),
    .LI(sig00000238),
    .O(sig00000220)
  );
  MUXCY   blk000000ee (
    .CI(sig000001f1),
    .DI(sig00000181),
    .S(sig0000022d),
    .O(sig000001f2)
  );
  XORCY   blk000000ef (
    .CI(sig000001f1),
    .LI(sig0000022d),
    .O(sig00000214)
  );
  MUXCY   blk000000f0 (
    .CI(sig000001f2),
    .DI(sig00000182),
    .S(sig0000022e),
    .O(sig000001f3)
  );
  XORCY   blk000000f1 (
    .CI(sig000001f2),
    .LI(sig0000022e),
    .O(sig00000215)
  );
  MUXCY   blk000000f2 (
    .CI(sig000001f3),
    .DI(sig00000183),
    .S(sig0000022f),
    .O(sig000001f4)
  );
  XORCY   blk000000f3 (
    .CI(sig000001f3),
    .LI(sig0000022f),
    .O(sig00000216)
  );
  XORCY   blk000000f4 (
    .CI(sig000001f4),
    .LI(sig000001f0),
    .O(sig00000217)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000f5 (
    .C(clk),
    .CE(ce),
    .D(sig00000213),
    .Q(sig000001ff)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000f6 (
    .C(clk),
    .CE(ce),
    .D(sig00000218),
    .Q(sig00000200)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000f7 (
    .C(clk),
    .CE(ce),
    .D(sig00000219),
    .Q(sig00000205)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000f8 (
    .C(clk),
    .CE(ce),
    .D(sig0000021a),
    .Q(sig00000206)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000f9 (
    .C(clk),
    .CE(ce),
    .D(sig0000021b),
    .Q(sig00000207)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000fa (
    .C(clk),
    .CE(ce),
    .D(sig0000021c),
    .Q(sig00000208)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000fb (
    .C(clk),
    .CE(ce),
    .D(sig0000021d),
    .Q(sig00000209)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000fc (
    .C(clk),
    .CE(ce),
    .D(sig0000021e),
    .Q(sig0000020a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000fd (
    .C(clk),
    .CE(ce),
    .D(sig0000021f),
    .Q(sig0000020b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000fe (
    .C(clk),
    .CE(ce),
    .D(sig00000220),
    .Q(sig0000020c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000ff (
    .C(clk),
    .CE(ce),
    .D(sig00000214),
    .Q(sig00000201)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000100 (
    .C(clk),
    .CE(ce),
    .D(sig00000215),
    .Q(sig00000202)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000101 (
    .C(clk),
    .CE(ce),
    .D(sig00000216),
    .Q(sig00000203)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000102 (
    .C(clk),
    .CE(ce),
    .D(sig00000217),
    .Q(sig00000204)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000103 (
    .C(clk),
    .CE(ce),
    .D(sig000000ca),
    .Q(sig000001ad)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000104 (
    .C(clk),
    .CE(ce),
    .D(sig000000cb),
    .Q(sig000001ae)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000105 (
    .C(clk),
    .CE(ce),
    .D(sig000000cc),
    .Q(sig000001b2)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000106 (
    .C(clk),
    .CE(ce),
    .D(sig000000cd),
    .Q(sig000001b3)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000107 (
    .C(clk),
    .CE(ce),
    .D(sig000000ce),
    .Q(sig000001b4)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000108 (
    .C(clk),
    .CE(ce),
    .D(sig000000cf),
    .Q(sig000001b5)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000109 (
    .C(clk),
    .CE(ce),
    .D(sig000000d0),
    .Q(sig000001b6)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000010a (
    .C(clk),
    .CE(ce),
    .D(sig000000d2),
    .Q(sig000001b7)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000010b (
    .C(clk),
    .CE(ce),
    .D(sig000000d3),
    .Q(sig000001b8)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000010c (
    .C(clk),
    .CE(ce),
    .D(sig000000d4),
    .Q(sig000001b9)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000010d (
    .C(clk),
    .CE(ce),
    .D(sig000000d5),
    .Q(sig000001af)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000010e (
    .C(clk),
    .CE(ce),
    .D(sig000000d6),
    .Q(sig000001b0)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000010f (
    .C(clk),
    .CE(ce),
    .D(sig000000d7),
    .Q(sig000001b1)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000110 (
    .C(clk),
    .CE(ce),
    .D(sig00000273),
    .Q(sig00000172)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000111 (
    .C(clk),
    .CE(ce),
    .D(sig00000274),
    .Q(sig00000173)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000112 (
    .C(clk),
    .CE(ce),
    .D(sig00000275),
    .Q(sig00000177)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000113 (
    .C(clk),
    .CE(ce),
    .D(sig00000276),
    .Q(sig00000178)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000114 (
    .C(clk),
    .CE(ce),
    .D(sig00000277),
    .Q(sig00000179)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000115 (
    .C(clk),
    .CE(ce),
    .D(sig00000278),
    .Q(sig0000017a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000116 (
    .C(clk),
    .CE(ce),
    .D(sig00000279),
    .Q(sig0000017b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000117 (
    .C(clk),
    .CE(ce),
    .D(sig0000027a),
    .Q(sig0000017c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000118 (
    .C(clk),
    .CE(ce),
    .D(sig0000027b),
    .Q(sig0000017d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000119 (
    .C(clk),
    .CE(ce),
    .D(sig0000027d),
    .Q(sig0000017e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000011a (
    .C(clk),
    .CE(ce),
    .D(sig0000027e),
    .Q(sig00000174)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000011b (
    .C(clk),
    .CE(ce),
    .D(sig0000027f),
    .Q(sig00000175)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000011c (
    .C(clk),
    .CE(ce),
    .D(sig00000280),
    .Q(sig00000176)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000011d (
    .C(clk),
    .CE(ce),
    .D(sig00000271),
    .Q(sig000001a2)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000011e (
    .C(clk),
    .CE(ce),
    .D(sig0000027c),
    .Q(sig000001a3)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000011f (
    .C(clk),
    .CE(ce),
    .D(sig00000281),
    .Q(sig000001a5)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000120 (
    .C(clk),
    .CE(ce),
    .D(sig00000282),
    .Q(sig000001a6)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000121 (
    .C(clk),
    .CE(ce),
    .D(sig00000283),
    .Q(sig000001a7)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000122 (
    .C(clk),
    .CE(ce),
    .D(sig00000284),
    .Q(sig000001a8)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000123 (
    .C(clk),
    .CE(ce),
    .D(sig00000285),
    .Q(sig000001a9)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000124 (
    .C(clk),
    .CE(ce),
    .D(sig00000286),
    .Q(sig000001aa)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000125 (
    .C(clk),
    .CE(ce),
    .D(sig00000287),
    .Q(sig000001ab)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000126 (
    .C(clk),
    .CE(ce),
    .D(sig00000288),
    .Q(sig000001ac)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000127 (
    .C(clk),
    .CE(ce),
    .D(sig00000272),
    .Q(sig000001a4)
  );
  MUXCY   blk00000128 (
    .CI(sig0000020e),
    .DI(sig00000001),
    .S(sig000001ef),
    .O(sig0000020f)
  );
  MUXCY   blk00000129 (
    .CI(sig0000025a),
    .DI(sig00000001),
    .S(sig00000002),
    .O(sig0000020e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000012a (
    .C(clk),
    .CE(ce),
    .D(sig0000025a),
    .Q(sig000001fe)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000012b (
    .C(clk),
    .CE(ce),
    .D(sig00000261),
    .Q(sig0000020d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000012c (
    .C(clk),
    .CE(ce),
    .D(sig00000419),
    .Q(sig00000386)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000012d (
    .C(clk),
    .CE(ce),
    .D(sig0000041e),
    .Q(sig000003da)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000012e (
    .C(clk),
    .CE(ce),
    .D(sig000003e8),
    .Q(sig000002ea)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000012f (
    .C(clk),
    .CE(ce),
    .D(a[31]),
    .Q(sig000002d8)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000130 (
    .C(clk),
    .CE(ce),
    .D(sig000002ec),
    .Q(sig000002eb)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000131 (
    .C(clk),
    .CE(ce),
    .D(sig00000439),
    .Q(sig000002ec)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000132 (
    .C(clk),
    .CE(ce),
    .D(sig0000041b),
    .Q(sig000003d9)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000133 (
    .C(clk),
    .CE(ce),
    .D(sig0000040b),
    .Q(sig0000037c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000134 (
    .C(clk),
    .CE(ce),
    .D(sig0000040a),
    .Q(sig0000037d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000135 (
    .C(clk),
    .CE(ce),
    .D(sig0000041a),
    .Q(sig00000348)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000136 (
    .C(clk),
    .CE(ce),
    .D(sig000003dc),
    .Q(sig00000343)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000137 (
    .C(clk),
    .CE(ce),
    .D(sig000003e1),
    .Q(sig00000341)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000138 (
    .C(clk),
    .CE(ce),
    .D(sig000003e3),
    .Q(sig00000344)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000139 (
    .C(clk),
    .CE(ce),
    .D(sig000003e0),
    .Q(sig00000340)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000013a (
    .C(clk),
    .CE(ce),
    .D(sig000003db),
    .Q(sig0000033e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000013b (
    .C(clk),
    .CE(ce),
    .D(sig000003e2),
    .Q(sig00000342)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000013c (
    .C(clk),
    .CE(ce),
    .D(sig000005a2),
    .Q(sig0000033f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000013d (
    .C(clk),
    .CE(ce),
    .D(sig00000204),
    .Q(sig0000037a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000013e (
    .C(clk),
    .CE(ce),
    .D(sig00000302),
    .Q(sig000003e5)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000013f (
    .C(clk),
    .CE(ce),
    .D(sig00000306),
    .Q(sig000003e6)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000140 (
    .C(clk),
    .CE(ce),
    .D(sig000002ee),
    .Q(sig000003dd)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000141 (
    .C(clk),
    .CE(ce),
    .D(sig000002f2),
    .Q(sig000003de)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000142 (
    .I0(b[23]),
    .I1(a[23]),
    .O(sig00000361)
  );
  MUXCY   blk00000143 (
    .CI(sig00000002),
    .DI(b[23]),
    .S(sig00000361),
    .O(sig00000359)
  );
  XORCY   blk00000144 (
    .CI(sig00000002),
    .LI(sig00000361),
    .O(sig000003e9)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000145 (
    .I0(b[24]),
    .I1(a[24]),
    .O(sig00000362)
  );
  MUXCY   blk00000146 (
    .CI(sig00000359),
    .DI(b[24]),
    .S(sig00000362),
    .O(sig0000035a)
  );
  XORCY   blk00000147 (
    .CI(sig00000359),
    .LI(sig00000362),
    .O(sig000003ea)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000148 (
    .I0(b[25]),
    .I1(a[25]),
    .O(sig00000363)
  );
  MUXCY   blk00000149 (
    .CI(sig0000035a),
    .DI(b[25]),
    .S(sig00000363),
    .O(sig0000035b)
  );
  XORCY   blk0000014a (
    .CI(sig0000035a),
    .LI(sig00000363),
    .O(sig000003eb)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk0000014b (
    .I0(b[26]),
    .I1(a[26]),
    .O(sig00000364)
  );
  MUXCY   blk0000014c (
    .CI(sig0000035b),
    .DI(b[26]),
    .S(sig00000364),
    .O(sig0000035c)
  );
  XORCY   blk0000014d (
    .CI(sig0000035b),
    .LI(sig00000364),
    .O(sig000003ec)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk0000014e (
    .I0(b[27]),
    .I1(a[27]),
    .O(sig00000365)
  );
  MUXCY   blk0000014f (
    .CI(sig0000035c),
    .DI(b[27]),
    .S(sig00000365),
    .O(sig0000035d)
  );
  XORCY   blk00000150 (
    .CI(sig0000035c),
    .LI(sig00000365),
    .O(sig000003ed)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000151 (
    .I0(b[28]),
    .I1(a[28]),
    .O(sig00000366)
  );
  MUXCY   blk00000152 (
    .CI(sig0000035d),
    .DI(b[28]),
    .S(sig00000366),
    .O(sig0000035e)
  );
  XORCY   blk00000153 (
    .CI(sig0000035d),
    .LI(sig00000366),
    .O(sig000003ee)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000154 (
    .I0(b[29]),
    .I1(a[29]),
    .O(sig00000367)
  );
  MUXCY   blk00000155 (
    .CI(sig0000035e),
    .DI(b[29]),
    .S(sig00000367),
    .O(sig0000035f)
  );
  XORCY   blk00000156 (
    .CI(sig0000035e),
    .LI(sig00000367),
    .O(sig000003ef)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000157 (
    .I0(b[30]),
    .I1(a[30]),
    .O(sig00000368)
  );
  MUXCY   blk00000158 (
    .CI(sig0000035f),
    .DI(b[30]),
    .S(sig00000368),
    .O(sig00000360)
  );
  XORCY   blk00000159 (
    .CI(sig0000035f),
    .LI(sig00000368),
    .O(sig000003f0)
  );
  XORCY   blk0000015a (
    .CI(sig00000360),
    .LI(sig00000002),
    .O(sig000003f1)
  );
  MUXCY   blk0000015b (
    .CI(sig00000002),
    .DI(sig00000333),
    .S(sig00000371),
    .O(sig00000369)
  );
  XORCY   blk0000015c (
    .CI(sig00000002),
    .LI(sig00000371),
    .O(sig00000411)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk0000015d (
    .I0(sig00000334),
    .I1(sig0000045e),
    .O(sig00000372)
  );
  MUXCY   blk0000015e (
    .CI(sig00000369),
    .DI(sig00000334),
    .S(sig00000372),
    .O(sig0000036a)
  );
  XORCY   blk0000015f (
    .CI(sig00000369),
    .LI(sig00000372),
    .O(sig00000412)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000160 (
    .I0(sig00000335),
    .I1(sig0000045d),
    .O(sig00000373)
  );
  MUXCY   blk00000161 (
    .CI(sig0000036a),
    .DI(sig00000335),
    .S(sig00000373),
    .O(sig0000036b)
  );
  XORCY   blk00000162 (
    .CI(sig0000036a),
    .LI(sig00000373),
    .O(sig00000413)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000163 (
    .I0(sig00000336),
    .I1(sig0000043d),
    .O(sig00000374)
  );
  MUXCY   blk00000164 (
    .CI(sig0000036b),
    .DI(sig00000336),
    .S(sig00000374),
    .O(sig0000036c)
  );
  XORCY   blk00000165 (
    .CI(sig0000036b),
    .LI(sig00000374),
    .O(sig00000414)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000166 (
    .I0(sig00000337),
    .I1(sig0000043c),
    .O(sig00000375)
  );
  MUXCY   blk00000167 (
    .CI(sig0000036c),
    .DI(sig00000337),
    .S(sig00000375),
    .O(sig0000036d)
  );
  XORCY   blk00000168 (
    .CI(sig0000036c),
    .LI(sig00000375),
    .O(sig00000415)
  );
  MUXCY   blk00000169 (
    .CI(sig0000036d),
    .DI(sig00000338),
    .S(sig00000376),
    .O(sig0000036e)
  );
  XORCY   blk0000016a (
    .CI(sig0000036d),
    .LI(sig00000376),
    .O(sig00000416)
  );
  MUXCY   blk0000016b (
    .CI(sig0000036e),
    .DI(sig00000339),
    .S(sig00000377),
    .O(sig0000036f)
  );
  XORCY   blk0000016c (
    .CI(sig0000036e),
    .LI(sig00000377),
    .O(sig00000417)
  );
  MUXCY   blk0000016d (
    .CI(sig0000036f),
    .DI(sig0000033a),
    .S(sig00000378),
    .O(sig00000370)
  );
  XORCY   blk0000016e (
    .CI(sig0000036f),
    .LI(sig00000378),
    .O(sig00000418)
  );
  XORCY   blk0000016f (
    .CI(sig00000370),
    .LI(sig00000002),
    .O(sig00000419)
  );
  MUXCY   blk00000170 (
    .CI(sig00000301),
    .DI(sig00000001),
    .S(sig00000304),
    .O(sig00000302)
  );
  MUXCY   blk00000171 (
    .CI(sig00000002),
    .DI(sig00000001),
    .S(sig00000303),
    .O(sig00000301)
  );
  MUXCY   blk00000172 (
    .CI(sig00000305),
    .DI(sig00000001),
    .S(sig00000308),
    .O(sig00000306)
  );
  MUXCY   blk00000173 (
    .CI(sig00000002),
    .DI(sig00000001),
    .S(sig00000307),
    .O(sig00000305)
  );
  MUXCY   blk00000174 (
    .CI(sig000002ed),
    .DI(sig00000001),
    .S(sig000002f0),
    .O(sig000002ee)
  );
  MUXCY   blk00000175 (
    .CI(sig00000002),
    .DI(sig00000001),
    .S(sig000002ef),
    .O(sig000002ed)
  );
  MUXCY   blk00000176 (
    .CI(sig000002f1),
    .DI(sig00000001),
    .S(sig000002f4),
    .O(sig000002f2)
  );
  MUXCY   blk00000177 (
    .CI(sig00000002),
    .DI(sig00000001),
    .S(sig000002f3),
    .O(sig000002f1)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000178 (
    .C(clk),
    .CE(ce),
    .D(sig00000357),
    .Q(sig00000319)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000179 (
    .C(clk),
    .CE(ce),
    .D(sig0000041d),
    .Q(sig00000318)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000017a (
    .C(clk),
    .CE(ce),
    .D(sig000003f3),
    .Q(sig00000317)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000017b (
    .C(clk),
    .CE(ce),
    .D(sig000003f2),
    .Q(sig00000316)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000017c (
    .C(clk),
    .CE(ce),
    .D(sig0000041c),
    .Q(sig00000315)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000017d (
    .C(clk),
    .CE(ce),
    .D(sig000002fa),
    .Q(sig000003df)
  );
  MUXCY   blk0000017e (
    .CI(sig00000002),
    .DI(sig00000001),
    .S(sig000002fb),
    .O(sig000002f5)
  );
  MUXCY   blk0000017f (
    .CI(sig000002f5),
    .DI(sig00000001),
    .S(sig000002fc),
    .O(sig000002f6)
  );
  MUXCY   blk00000180 (
    .CI(sig000002f6),
    .DI(sig00000001),
    .S(sig000002fd),
    .O(sig000002f7)
  );
  MUXCY   blk00000181 (
    .CI(sig000002f7),
    .DI(sig00000001),
    .S(sig000002fe),
    .O(sig000002f8)
  );
  MUXCY   blk00000182 (
    .CI(sig000002f8),
    .DI(sig00000001),
    .S(sig000002ff),
    .O(sig000002f9)
  );
  MUXCY   blk00000183 (
    .CI(sig000002f9),
    .DI(sig00000001),
    .S(sig00000300),
    .O(sig000002fa)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000184 (
    .C(clk),
    .CE(ce),
    .D(sig0000030e),
    .Q(sig000003e7)
  );
  MUXCY   blk00000185 (
    .CI(sig00000002),
    .DI(sig00000001),
    .S(sig0000030f),
    .O(sig00000309)
  );
  MUXCY   blk00000186 (
    .CI(sig00000309),
    .DI(sig00000001),
    .S(sig00000310),
    .O(sig0000030a)
  );
  MUXCY   blk00000187 (
    .CI(sig0000030a),
    .DI(sig00000001),
    .S(sig00000311),
    .O(sig0000030b)
  );
  MUXCY   blk00000188 (
    .CI(sig0000030b),
    .DI(sig00000001),
    .S(sig00000312),
    .O(sig0000030c)
  );
  MUXCY   blk00000189 (
    .CI(sig0000030c),
    .DI(sig00000001),
    .S(sig00000313),
    .O(sig0000030d)
  );
  MUXCY   blk0000018a (
    .CI(sig0000030d),
    .DI(sig00000001),
    .S(sig00000314),
    .O(sig0000030e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000018b (
    .C(clk),
    .CE(ce),
    .D(sig00000385),
    .Q(sig00000356)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000018c (
    .C(clk),
    .CE(ce),
    .D(sig00000384),
    .Q(sig00000355)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000018d (
    .C(clk),
    .CE(ce),
    .D(sig00000383),
    .Q(sig00000354)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000018e (
    .C(clk),
    .CE(ce),
    .D(sig00000382),
    .Q(sig00000353)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000018f (
    .C(clk),
    .CE(ce),
    .D(sig00000381),
    .Q(sig00000352)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000190 (
    .C(clk),
    .CE(ce),
    .D(sig00000380),
    .Q(sig00000351)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000191 (
    .C(clk),
    .CE(ce),
    .D(sig0000037f),
    .Q(sig00000350)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000192 (
    .C(clk),
    .CE(ce),
    .D(sig0000037e),
    .Q(sig0000034f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000193 (
    .C(clk),
    .CE(ce),
    .D(sig00000418),
    .Q(sig00000385)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000194 (
    .C(clk),
    .CE(ce),
    .D(sig00000417),
    .Q(sig00000384)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000195 (
    .C(clk),
    .CE(ce),
    .D(sig00000416),
    .Q(sig00000383)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000196 (
    .C(clk),
    .CE(ce),
    .D(sig00000415),
    .Q(sig00000382)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000197 (
    .C(clk),
    .CE(ce),
    .D(sig00000414),
    .Q(sig00000381)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000198 (
    .C(clk),
    .CE(ce),
    .D(sig00000413),
    .Q(sig00000380)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000199 (
    .C(clk),
    .CE(ce),
    .D(sig00000412),
    .Q(sig0000037f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000019a (
    .C(clk),
    .CE(ce),
    .D(sig00000411),
    .Q(sig0000037e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000019b (
    .C(clk),
    .CE(ce),
    .D(b[30]),
    .Q(sig000002e9)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000019c (
    .C(clk),
    .CE(ce),
    .D(b[29]),
    .Q(sig000002e8)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000019d (
    .C(clk),
    .CE(ce),
    .D(b[28]),
    .Q(sig000002e7)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000019e (
    .C(clk),
    .CE(ce),
    .D(b[27]),
    .Q(sig000002e6)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000019f (
    .C(clk),
    .CE(ce),
    .D(b[26]),
    .Q(sig000002e5)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001a0 (
    .C(clk),
    .CE(ce),
    .D(b[25]),
    .Q(sig000002e4)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001a1 (
    .C(clk),
    .CE(ce),
    .D(b[24]),
    .Q(sig000002e3)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001a2 (
    .C(clk),
    .CE(ce),
    .D(b[23]),
    .Q(sig000002e2)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001a3 (
    .C(clk),
    .CE(ce),
    .D(a[30]),
    .Q(sig000002d7)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001a4 (
    .C(clk),
    .CE(ce),
    .D(a[29]),
    .Q(sig000002d6)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001a5 (
    .C(clk),
    .CE(ce),
    .D(a[28]),
    .Q(sig000002d5)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001a6 (
    .C(clk),
    .CE(ce),
    .D(a[27]),
    .Q(sig000002d4)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001a7 (
    .C(clk),
    .CE(ce),
    .D(a[26]),
    .Q(sig000002d3)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001a8 (
    .C(clk),
    .CE(ce),
    .D(a[25]),
    .Q(sig000002d2)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001a9 (
    .C(clk),
    .CE(ce),
    .D(a[24]),
    .Q(sig000002d1)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001aa (
    .C(clk),
    .CE(ce),
    .D(a[23]),
    .Q(sig000002d0)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001ab (
    .C(clk),
    .CE(ce),
    .D(sig000003f1),
    .Q(sig000002e1)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001ac (
    .C(clk),
    .CE(ce),
    .D(sig000003f0),
    .Q(sig000002e0)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001ad (
    .C(clk),
    .CE(ce),
    .D(sig000003ef),
    .Q(sig000002df)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001ae (
    .C(clk),
    .CE(ce),
    .D(sig000003ee),
    .Q(sig000002de)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001af (
    .C(clk),
    .CE(ce),
    .D(sig000003ed),
    .Q(sig000002dd)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001b0 (
    .C(clk),
    .CE(ce),
    .D(sig000003ec),
    .Q(sig000002dc)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001b1 (
    .C(clk),
    .CE(ce),
    .D(sig000003eb),
    .Q(sig000002db)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001b2 (
    .C(clk),
    .CE(ce),
    .D(sig000003ea),
    .Q(sig000002da)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001b3 (
    .C(clk),
    .CE(ce),
    .D(sig000003e9),
    .Q(sig000002d9)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001b4 (
    .C(clk),
    .CE(ce),
    .D(sig000003f9),
    .Q(sig0000034e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001b5 (
    .C(clk),
    .CE(ce),
    .D(sig000003f8),
    .Q(sig0000034d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001b6 (
    .C(clk),
    .CE(ce),
    .D(sig000003f4),
    .Q(sig00000347)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001b7 (
    .C(clk),
    .CE(ce),
    .D(sig00000402),
    .Q(sig0000032a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001b8 (
    .C(clk),
    .CE(ce),
    .D(sig00000401),
    .Q(sig00000329)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001b9 (
    .C(clk),
    .CE(ce),
    .D(sig00000400),
    .Q(sig00000328)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001ba (
    .C(clk),
    .CE(ce),
    .D(sig000003ff),
    .Q(sig00000327)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001bb (
    .C(clk),
    .CE(ce),
    .D(sig000003fe),
    .Q(sig00000326)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001bc (
    .C(clk),
    .CE(ce),
    .D(sig000003fd),
    .Q(sig00000325)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001bd (
    .C(clk),
    .CE(ce),
    .D(sig000003fc),
    .Q(sig00000324)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001be (
    .C(clk),
    .CE(ce),
    .D(sig000003fb),
    .Q(sig00000323)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001bf (
    .C(clk),
    .CE(ce),
    .D(sig000003fa),
    .Q(sig00000322)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001c0 (
    .C(clk),
    .CE(ce),
    .D(sig0000040e),
    .Q(sig0000033c)
  );
  XORCY   blk000001c1 (
    .CI(sig00000321),
    .LI(sig00000001),
    .O(sig00000402)
  );
  XORCY   blk000001c2 (
    .CI(sig00000320),
    .LI(sig00000409),
    .O(sig00000401)
  );
  MUXCY   blk000001c3 (
    .CI(sig00000320),
    .DI(sig00000001),
    .S(sig00000409),
    .O(sig00000321)
  );
  XORCY   blk000001c4 (
    .CI(sig0000031f),
    .LI(sig00000408),
    .O(sig00000400)
  );
  MUXCY   blk000001c5 (
    .CI(sig0000031f),
    .DI(sig00000001),
    .S(sig00000408),
    .O(sig00000320)
  );
  XORCY   blk000001c6 (
    .CI(sig0000031e),
    .LI(sig00000407),
    .O(sig000003ff)
  );
  MUXCY   blk000001c7 (
    .CI(sig0000031e),
    .DI(sig00000001),
    .S(sig00000407),
    .O(sig0000031f)
  );
  XORCY   blk000001c8 (
    .CI(sig0000031d),
    .LI(sig00000406),
    .O(sig000003fe)
  );
  MUXCY   blk000001c9 (
    .CI(sig0000031d),
    .DI(sig00000001),
    .S(sig00000406),
    .O(sig0000031e)
  );
  XORCY   blk000001ca (
    .CI(sig0000031c),
    .LI(sig00000405),
    .O(sig000003fd)
  );
  MUXCY   blk000001cb (
    .CI(sig0000031c),
    .DI(sig00000001),
    .S(sig00000405),
    .O(sig0000031d)
  );
  XORCY   blk000001cc (
    .CI(sig0000031b),
    .LI(sig00000404),
    .O(sig000003fc)
  );
  MUXCY   blk000001cd (
    .CI(sig0000031b),
    .DI(sig00000001),
    .S(sig00000404),
    .O(sig0000031c)
  );
  XORCY   blk000001ce (
    .CI(sig0000031a),
    .LI(sig00000403),
    .O(sig000003fb)
  );
  MUXCY   blk000001cf (
    .CI(sig0000031a),
    .DI(sig00000001),
    .S(sig00000403),
    .O(sig0000031b)
  );
  XORCY   blk000001d0 (
    .CI(sig00000001),
    .LI(sig000003e4),
    .O(sig000003fa)
  );
  MUXCY   blk000001d1 (
    .CI(sig00000001),
    .DI(sig00000002),
    .S(sig000003e4),
    .O(sig0000031a)
  );
  MUXCY   blk000001d2 (
    .CI(sig000003cc),
    .DI(sig00000001),
    .S(sig00000002),
    .O(sig000003cd)
  );
  MUXCY   blk000001d3 (
    .CI(sig000003cb),
    .DI(a[30]),
    .S(sig000003c5),
    .O(sig000003cc)
  );
  MUXCY   blk000001d4 (
    .CI(sig000003ca),
    .DI(a[29]),
    .S(sig000003c4),
    .O(sig000003cb)
  );
  MUXCY   blk000001d5 (
    .CI(sig000003c9),
    .DI(a[28]),
    .S(sig000003c3),
    .O(sig000003ca)
  );
  MUXCY   blk000001d6 (
    .CI(sig000003c8),
    .DI(a[27]),
    .S(sig000003c1),
    .O(sig000003c9)
  );
  MUXCY   blk000001d7 (
    .CI(sig000003c7),
    .DI(a[26]),
    .S(sig000003c0),
    .O(sig000003c8)
  );
  MUXCY   blk000001d8 (
    .CI(sig000003d6),
    .DI(a[25]),
    .S(sig000003be),
    .O(sig000003c7)
  );
  MUXCY   blk000001d9 (
    .CI(sig000003d5),
    .DI(a[24]),
    .S(sig000003bd),
    .O(sig000003d6)
  );
  MUXCY   blk000001da (
    .CI(sig000003d4),
    .DI(a[23]),
    .S(sig000003bb),
    .O(sig000003d5)
  );
  MUXCY   blk000001db (
    .CI(sig000003d3),
    .DI(a[22]),
    .S(sig000003ba),
    .O(sig000003d4)
  );
  MUXCY   blk000001dc (
    .CI(sig000003d2),
    .DI(a[21]),
    .S(sig000003b8),
    .O(sig000003d3)
  );
  MUXCY   blk000001dd (
    .CI(sig000003d1),
    .DI(a[20]),
    .S(sig000003b7),
    .O(sig000003d2)
  );
  MUXCY   blk000001de (
    .CI(sig000003d0),
    .DI(a[19]),
    .S(sig000003b5),
    .O(sig000003d1)
  );
  MUXCY   blk000001df (
    .CI(sig000003cf),
    .DI(a[18]),
    .S(sig000003b4),
    .O(sig000003d0)
  );
  MUXCY   blk000001e0 (
    .CI(sig000003ce),
    .DI(a[17]),
    .S(sig000003b2),
    .O(sig000003cf)
  );
  MUXCY   blk000001e1 (
    .CI(sig00000002),
    .DI(a[16]),
    .S(sig000003b1),
    .O(sig000003ce)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001e2 (
    .C(clk),
    .CE(ce),
    .D(sig000003cd),
    .Q(sig000003d7)
  );
  MUXCY   blk000001e3 (
    .CI(sig0000038c),
    .DI(a[15]),
    .S(sig0000039d),
    .O(sig0000038d)
  );
  MUXCY   blk000001e4 (
    .CI(sig0000038b),
    .DI(a[14]),
    .S(sig0000039c),
    .O(sig0000038c)
  );
  MUXCY   blk000001e5 (
    .CI(sig0000038a),
    .DI(a[13]),
    .S(sig0000039b),
    .O(sig0000038b)
  );
  MUXCY   blk000001e6 (
    .CI(sig00000389),
    .DI(a[12]),
    .S(sig0000039a),
    .O(sig0000038a)
  );
  MUXCY   blk000001e7 (
    .CI(sig00000388),
    .DI(a[11]),
    .S(sig00000399),
    .O(sig00000389)
  );
  MUXCY   blk000001e8 (
    .CI(sig00000387),
    .DI(a[10]),
    .S(sig00000398),
    .O(sig00000388)
  );
  MUXCY   blk000001e9 (
    .CI(sig00000396),
    .DI(a[9]),
    .S(sig000003a6),
    .O(sig00000387)
  );
  MUXCY   blk000001ea (
    .CI(sig00000395),
    .DI(a[8]),
    .S(sig000003a5),
    .O(sig00000396)
  );
  MUXCY   blk000001eb (
    .CI(sig00000394),
    .DI(a[7]),
    .S(sig000003a4),
    .O(sig00000395)
  );
  MUXCY   blk000001ec (
    .CI(sig00000393),
    .DI(a[6]),
    .S(sig000003a3),
    .O(sig00000394)
  );
  MUXCY   blk000001ed (
    .CI(sig00000392),
    .DI(a[5]),
    .S(sig000003a2),
    .O(sig00000393)
  );
  MUXCY   blk000001ee (
    .CI(sig00000391),
    .DI(a[4]),
    .S(sig000003a1),
    .O(sig00000392)
  );
  MUXCY   blk000001ef (
    .CI(sig00000390),
    .DI(a[3]),
    .S(sig000003a0),
    .O(sig00000391)
  );
  MUXCY   blk000001f0 (
    .CI(sig0000038f),
    .DI(a[2]),
    .S(sig0000039f),
    .O(sig00000390)
  );
  MUXCY   blk000001f1 (
    .CI(sig0000038e),
    .DI(a[1]),
    .S(sig0000039e),
    .O(sig0000038f)
  );
  MUXCY   blk000001f2 (
    .CI(sig00000002),
    .DI(a[0]),
    .S(sig00000397),
    .O(sig0000038e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001f3 (
    .C(clk),
    .CE(ce),
    .D(sig0000038d),
    .Q(sig000003a7)
  );
  MUXCY   blk000001f4 (
    .CI(sig000003ae),
    .DI(sig00000001),
    .S(sig000003c6),
    .O(sig000003af)
  );
  MUXCY   blk000001f5 (
    .CI(sig000003ad),
    .DI(sig00000001),
    .S(sig000003c2),
    .O(sig000003ae)
  );
  MUXCY   blk000001f6 (
    .CI(sig000003ac),
    .DI(sig00000001),
    .S(sig000003bf),
    .O(sig000003ad)
  );
  MUXCY   blk000001f7 (
    .CI(sig000003ab),
    .DI(sig00000001),
    .S(sig000003bc),
    .O(sig000003ac)
  );
  MUXCY   blk000001f8 (
    .CI(sig000003aa),
    .DI(sig00000001),
    .S(sig000003b9),
    .O(sig000003ab)
  );
  MUXCY   blk000001f9 (
    .CI(sig000003a9),
    .DI(sig00000001),
    .S(sig000003b6),
    .O(sig000003aa)
  );
  MUXCY   blk000001fa (
    .CI(sig000003a8),
    .DI(sig00000001),
    .S(sig000003b3),
    .O(sig000003a9)
  );
  MUXCY   blk000001fb (
    .CI(sig00000002),
    .DI(sig00000001),
    .S(sig000003b0),
    .O(sig000003a8)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001fc (
    .C(clk),
    .CE(ce),
    .D(sig000003af),
    .Q(sig000003d8)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001fd (
    .C(clk),
    .CE(ce),
    .D(sig00000582),
    .Q(sig00000560)
  );
  MUXCY   blk000001fe (
    .CI(sig00000002),
    .DI(sig00000001),
    .S(sig00000563),
    .O(sig00000561)
  );
  MUXCY   blk000001ff (
    .CI(sig00000561),
    .DI(sig00000002),
    .S(sig00000566),
    .O(sig00000562)
  );
  MUXCY   blk00000200 (
    .CI(sig00000562),
    .DI(sig00000001),
    .S(sig00000565),
    .O(sig0000057f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000201 (
    .C(clk),
    .CE(ce),
    .D(sig000004a9),
    .Q(sig00000557)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000202 (
    .C(clk),
    .CE(ce),
    .D(sig000004b4),
    .Q(sig00000556)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000203 (
    .C(clk),
    .CE(ce),
    .D(sig000004bc),
    .Q(sig00000555)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000204 (
    .C(clk),
    .CE(ce),
    .D(sig000004bd),
    .Q(sig00000554)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000205 (
    .C(clk),
    .CE(ce),
    .D(sig000004be),
    .Q(sig0000055f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000206 (
    .C(clk),
    .CE(ce),
    .D(sig000004bf),
    .Q(sig0000055e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000207 (
    .C(clk),
    .CE(ce),
    .D(sig000004c0),
    .Q(sig0000055d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000208 (
    .C(clk),
    .CE(ce),
    .D(sig000004c1),
    .Q(sig0000055c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000209 (
    .C(clk),
    .CE(ce),
    .D(sig000004c2),
    .Q(sig0000055b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000020a (
    .C(clk),
    .CE(ce),
    .D(sig000004aa),
    .Q(sig0000055a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000020b (
    .C(clk),
    .CE(ce),
    .D(sig000004ab),
    .Q(sig00000559)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000020c (
    .C(clk),
    .CE(ce),
    .D(sig000004ac),
    .Q(sig00000558)
  );
  XORCY   blk0000020d (
    .CI(sig000004fd),
    .LI(sig00000001),
    .O(NLW_blk0000020d_O_UNCONNECTED)
  );
  XORCY   blk0000020e (
    .CI(sig000004fc),
    .LI(sig00000001),
    .O(NLW_blk0000020e_O_UNCONNECTED)
  );
  MUXCY   blk0000020f (
    .CI(sig000004fc),
    .DI(sig00000001),
    .S(sig00000001),
    .O(sig000004fd)
  );
  XORCY   blk00000210 (
    .CI(sig000004fb),
    .LI(sig00000001),
    .O(NLW_blk00000210_O_UNCONNECTED)
  );
  MUXCY   blk00000211 (
    .CI(sig000004fb),
    .DI(sig00000001),
    .S(sig00000001),
    .O(sig000004fc)
  );
  XORCY   blk00000212 (
    .CI(sig000004fa),
    .LI(sig00000001),
    .O(NLW_blk00000212_O_UNCONNECTED)
  );
  MUXCY   blk00000213 (
    .CI(sig000004fa),
    .DI(sig00000001),
    .S(sig00000001),
    .O(sig000004fb)
  );
  XORCY   blk00000214 (
    .CI(sig000004f9),
    .LI(sig00000001),
    .O(NLW_blk00000214_O_UNCONNECTED)
  );
  MUXCY   blk00000215 (
    .CI(sig000004f9),
    .DI(sig00000001),
    .S(sig00000001),
    .O(sig000004fa)
  );
  XORCY   blk00000216 (
    .CI(sig000004f8),
    .LI(sig00000001),
    .O(NLW_blk00000216_O_UNCONNECTED)
  );
  MUXCY   blk00000217 (
    .CI(sig000004f8),
    .DI(sig00000001),
    .S(sig00000001),
    .O(sig000004f9)
  );
  XORCY   blk00000218 (
    .CI(sig000004f7),
    .LI(sig00000001),
    .O(NLW_blk00000218_O_UNCONNECTED)
  );
  MUXCY   blk00000219 (
    .CI(sig000004f7),
    .DI(sig00000001),
    .S(sig00000001),
    .O(sig000004f8)
  );
  XORCY   blk0000021a (
    .CI(sig00000567),
    .LI(sig00000001),
    .O(NLW_blk0000021a_O_UNCONNECTED)
  );
  MUXCY   blk0000021b (
    .CI(sig00000567),
    .DI(sig00000001),
    .S(sig00000001),
    .O(sig000004f7)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000021c (
    .C(clk),
    .CE(ce),
    .D(sig00000523),
    .Q(sig0000050a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000021d (
    .C(clk),
    .CE(ce),
    .D(sig00000526),
    .Q(sig0000050b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000021e (
    .C(clk),
    .CE(ce),
    .D(sig00000527),
    .Q(sig0000050e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000021f (
    .C(clk),
    .CE(ce),
    .D(sig00000528),
    .Q(sig0000050f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000220 (
    .C(clk),
    .CE(ce),
    .D(sig00000529),
    .Q(sig00000510)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000221 (
    .C(clk),
    .CE(ce),
    .D(sig0000052a),
    .Q(sig00000511)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000222 (
    .C(clk),
    .CE(ce),
    .D(sig0000052b),
    .Q(sig00000512)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000223 (
    .C(clk),
    .CE(ce),
    .D(sig0000052c),
    .Q(sig00000513)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000224 (
    .C(clk),
    .CE(ce),
    .D(sig0000052d),
    .Q(sig00000514)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000225 (
    .C(clk),
    .CE(ce),
    .D(sig0000052e),
    .Q(sig00000515)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000226 (
    .C(clk),
    .CE(ce),
    .D(sig00000524),
    .Q(sig0000050c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000227 (
    .C(clk),
    .CE(ce),
    .D(sig00000525),
    .Q(sig0000050d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000228 (
    .C(clk),
    .CE(ce),
    .D(sig0000050a),
    .Q(sig000004fe)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000229 (
    .C(clk),
    .CE(ce),
    .D(sig0000050b),
    .Q(sig000004ff)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000022a (
    .C(clk),
    .CE(ce),
    .D(sig0000050e),
    .Q(sig00000502)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000022b (
    .C(clk),
    .CE(ce),
    .D(sig0000050f),
    .Q(sig00000503)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000022c (
    .C(clk),
    .CE(ce),
    .D(sig00000510),
    .Q(sig00000504)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000022d (
    .C(clk),
    .CE(ce),
    .D(sig00000511),
    .Q(sig00000505)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000022e (
    .C(clk),
    .CE(ce),
    .D(sig00000512),
    .Q(sig00000506)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000022f (
    .C(clk),
    .CE(ce),
    .D(sig00000513),
    .Q(sig00000507)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000230 (
    .C(clk),
    .CE(ce),
    .D(sig00000514),
    .Q(sig00000508)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000231 (
    .C(clk),
    .CE(ce),
    .D(sig00000515),
    .Q(sig00000509)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000232 (
    .C(clk),
    .CE(ce),
    .D(sig0000050c),
    .Q(sig00000500)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000233 (
    .C(clk),
    .CE(ce),
    .D(sig0000050d),
    .Q(sig00000501)
  );
  XORCY   blk00000234 (
    .CI(sig00000518),
    .LI(sig00000001),
    .O(sig00000522)
  );
  XORCY   blk00000235 (
    .CI(sig00000517),
    .LI(sig0000056a),
    .O(sig00000525)
  );
  MUXCY   blk00000236 (
    .CI(sig00000517),
    .DI(sig00000001),
    .S(sig0000056a),
    .O(sig00000518)
  );
  XORCY   blk00000237 (
    .CI(sig00000516),
    .LI(sig00000569),
    .O(sig00000524)
  );
  MUXCY   blk00000238 (
    .CI(sig00000516),
    .DI(sig00000001),
    .S(sig00000569),
    .O(sig00000517)
  );
  XORCY   blk00000239 (
    .CI(sig00000521),
    .LI(sig00000573),
    .O(sig0000052e)
  );
  MUXCY   blk0000023a (
    .CI(sig00000521),
    .DI(sig00000001),
    .S(sig00000573),
    .O(sig00000516)
  );
  XORCY   blk0000023b (
    .CI(sig00000520),
    .LI(sig00000572),
    .O(sig0000052d)
  );
  MUXCY   blk0000023c (
    .CI(sig00000520),
    .DI(sig00000001),
    .S(sig00000572),
    .O(sig00000521)
  );
  XORCY   blk0000023d (
    .CI(sig0000051f),
    .LI(sig00000571),
    .O(sig0000052c)
  );
  MUXCY   blk0000023e (
    .CI(sig0000051f),
    .DI(sig00000001),
    .S(sig00000571),
    .O(sig00000520)
  );
  XORCY   blk0000023f (
    .CI(sig0000051e),
    .LI(sig00000570),
    .O(sig0000052b)
  );
  MUXCY   blk00000240 (
    .CI(sig0000051e),
    .DI(sig00000001),
    .S(sig00000570),
    .O(sig0000051f)
  );
  XORCY   blk00000241 (
    .CI(sig0000051d),
    .LI(sig0000056f),
    .O(sig0000052a)
  );
  MUXCY   blk00000242 (
    .CI(sig0000051d),
    .DI(sig00000001),
    .S(sig0000056f),
    .O(sig0000051e)
  );
  XORCY   blk00000243 (
    .CI(sig0000051c),
    .LI(sig0000056e),
    .O(sig00000529)
  );
  MUXCY   blk00000244 (
    .CI(sig0000051c),
    .DI(sig00000001),
    .S(sig0000056e),
    .O(sig0000051d)
  );
  XORCY   blk00000245 (
    .CI(sig0000051b),
    .LI(sig0000056d),
    .O(sig00000528)
  );
  MUXCY   blk00000246 (
    .CI(sig0000051b),
    .DI(sig00000001),
    .S(sig0000056d),
    .O(sig0000051c)
  );
  XORCY   blk00000247 (
    .CI(sig0000051a),
    .LI(sig0000056c),
    .O(sig00000527)
  );
  MUXCY   blk00000248 (
    .CI(sig0000051a),
    .DI(sig00000001),
    .S(sig0000056c),
    .O(sig0000051b)
  );
  XORCY   blk00000249 (
    .CI(sig00000519),
    .LI(sig0000056b),
    .O(sig00000526)
  );
  MUXCY   blk0000024a (
    .CI(sig00000519),
    .DI(sig00000001),
    .S(sig0000056b),
    .O(sig0000051a)
  );
  XORCY   blk0000024b (
    .CI(sig0000057f),
    .LI(sig00000564),
    .O(sig00000523)
  );
  MUXCY   blk0000024c (
    .CI(sig0000057f),
    .DI(sig00000001),
    .S(sig00000564),
    .O(sig00000519)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000024d (
    .C(clk),
    .CE(ce),
    .D(sig00000522),
    .Q(sig00000568)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000024e (
    .C(clk),
    .CE(ce),
    .D(sig00000548),
    .Q(sig0000052f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000024f (
    .C(clk),
    .CE(ce),
    .D(sig0000054b),
    .Q(sig00000530)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000250 (
    .C(clk),
    .CE(ce),
    .D(sig0000054c),
    .Q(sig00000533)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000251 (
    .C(clk),
    .CE(ce),
    .D(sig0000054d),
    .Q(sig00000534)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000252 (
    .C(clk),
    .CE(ce),
    .D(sig0000054e),
    .Q(sig00000535)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000253 (
    .C(clk),
    .CE(ce),
    .D(sig0000054f),
    .Q(sig00000536)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000254 (
    .C(clk),
    .CE(ce),
    .D(sig00000550),
    .Q(sig00000537)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000255 (
    .C(clk),
    .CE(ce),
    .D(sig00000551),
    .Q(sig00000538)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000256 (
    .C(clk),
    .CE(ce),
    .D(sig00000552),
    .Q(sig00000539)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000257 (
    .C(clk),
    .CE(ce),
    .D(sig00000553),
    .Q(sig0000053a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000258 (
    .C(clk),
    .CE(ce),
    .D(sig00000549),
    .Q(sig00000531)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000259 (
    .C(clk),
    .CE(ce),
    .D(sig0000054a),
    .Q(sig00000532)
  );
  XORCY   blk0000025a (
    .CI(sig0000053d),
    .LI(sig00000001),
    .O(sig00000547)
  );
  XORCY   blk0000025b (
    .CI(sig0000053c),
    .LI(sig00000002),
    .O(sig0000054a)
  );
  MUXCY   blk0000025c (
    .CI(sig0000053c),
    .DI(sig00000001),
    .S(sig00000002),
    .O(sig0000053d)
  );
  XORCY   blk0000025d (
    .CI(sig0000053b),
    .LI(sig00000575),
    .O(sig00000549)
  );
  MUXCY   blk0000025e (
    .CI(sig0000053b),
    .DI(sig00000001),
    .S(sig00000575),
    .O(sig0000053c)
  );
  XORCY   blk0000025f (
    .CI(sig00000546),
    .LI(sig0000057e),
    .O(sig00000553)
  );
  MUXCY   blk00000260 (
    .CI(sig00000546),
    .DI(sig00000001),
    .S(sig0000057e),
    .O(sig0000053b)
  );
  XORCY   blk00000261 (
    .CI(sig00000545),
    .LI(sig0000057d),
    .O(sig00000552)
  );
  MUXCY   blk00000262 (
    .CI(sig00000545),
    .DI(sig00000001),
    .S(sig0000057d),
    .O(sig00000546)
  );
  XORCY   blk00000263 (
    .CI(sig00000544),
    .LI(sig0000057c),
    .O(sig00000551)
  );
  MUXCY   blk00000264 (
    .CI(sig00000544),
    .DI(sig00000001),
    .S(sig0000057c),
    .O(sig00000545)
  );
  XORCY   blk00000265 (
    .CI(sig00000543),
    .LI(sig0000057b),
    .O(sig00000550)
  );
  MUXCY   blk00000266 (
    .CI(sig00000543),
    .DI(sig00000001),
    .S(sig0000057b),
    .O(sig00000544)
  );
  XORCY   blk00000267 (
    .CI(sig00000542),
    .LI(sig0000057a),
    .O(sig0000054f)
  );
  MUXCY   blk00000268 (
    .CI(sig00000542),
    .DI(sig00000001),
    .S(sig0000057a),
    .O(sig00000543)
  );
  XORCY   blk00000269 (
    .CI(sig00000541),
    .LI(sig00000579),
    .O(sig0000054e)
  );
  MUXCY   blk0000026a (
    .CI(sig00000541),
    .DI(sig00000001),
    .S(sig00000579),
    .O(sig00000542)
  );
  XORCY   blk0000026b (
    .CI(sig00000540),
    .LI(sig00000578),
    .O(sig0000054d)
  );
  MUXCY   blk0000026c (
    .CI(sig00000540),
    .DI(sig00000001),
    .S(sig00000578),
    .O(sig00000541)
  );
  XORCY   blk0000026d (
    .CI(sig0000053f),
    .LI(sig00000577),
    .O(sig0000054c)
  );
  MUXCY   blk0000026e (
    .CI(sig0000053f),
    .DI(sig00000001),
    .S(sig00000577),
    .O(sig00000540)
  );
  XORCY   blk0000026f (
    .CI(sig0000053e),
    .LI(sig00000576),
    .O(sig0000054b)
  );
  MUXCY   blk00000270 (
    .CI(sig0000053e),
    .DI(sig00000001),
    .S(sig00000576),
    .O(sig0000053f)
  );
  XORCY   blk00000271 (
    .CI(sig00000568),
    .LI(sig00000574),
    .O(sig00000548)
  );
  MUXCY   blk00000272 (
    .CI(sig00000568),
    .DI(sig00000001),
    .S(sig00000574),
    .O(sig0000053e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000273 (
    .C(clk),
    .CE(ce),
    .D(sig00000547),
    .Q(sig00000567)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000274 (
    .C(clk),
    .CE(ce),
    .D(sig00000473),
    .Q(sig00000439)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000275 (
    .C(clk),
    .CE(ce),
    .D(sig00000583),
    .Q(sig0000045e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000276 (
    .C(clk),
    .CE(ce),
    .D(sig0000044f),
    .Q(sig0000045d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000277 (
    .C(clk),
    .CE(ce),
    .D(sig0000043b),
    .Q(sig0000043d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000278 (
    .C(clk),
    .CE(ce),
    .D(sig00000584),
    .Q(sig0000043b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000279 (
    .C(clk),
    .CE(ce),
    .D(sig00000462),
    .Q(sig0000045f)
  );
  MUXF5   blk0000027a (
    .I0(sig00000463),
    .I1(sig00000464),
    .S(sig0000044f),
    .O(NLW_blk0000027a_O_UNCONNECTED)
  );
  MUXF5   blk0000027b (
    .I0(sig00000460),
    .I1(sig00000461),
    .S(sig0000044f),
    .O(sig00000462)
  );
  MUXCY   blk0000027c (
    .CI(sig0000046b),
    .DI(sig00000001),
    .S(sig0000048c),
    .O(sig0000046c)
  );
  MUXCY   blk0000027d (
    .CI(sig0000046a),
    .DI(sig00000001),
    .S(sig0000048b),
    .O(sig0000046b)
  );
  MUXCY   blk0000027e (
    .CI(sig00000469),
    .DI(sig00000001),
    .S(sig0000048a),
    .O(sig0000046a)
  );
  MUXCY   blk0000027f (
    .CI(sig00000468),
    .DI(sig00000001),
    .S(sig00000489),
    .O(sig00000469)
  );
  MUXCY   blk00000280 (
    .CI(sig00000467),
    .DI(sig00000001),
    .S(sig00000488),
    .O(sig00000468)
  );
  MUXCY   blk00000281 (
    .CI(sig00000466),
    .DI(sig00000001),
    .S(sig00000487),
    .O(sig00000467)
  );
  MUXCY   blk00000282 (
    .CI(sig00000465),
    .DI(sig00000001),
    .S(sig00000486),
    .O(sig00000466)
  );
  MUXCY   blk00000283 (
    .CI(sig00000002),
    .DI(sig00000001),
    .S(sig00000481),
    .O(sig00000465)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000284 (
    .C(clk),
    .CE(ce),
    .D(sig0000046c),
    .Q(sig00000585)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000285 (
    .C(clk),
    .CE(ce),
    .D(sig0000046b),
    .Q(sig0000047e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000286 (
    .C(clk),
    .CE(ce),
    .D(sig0000046a),
    .Q(sig0000047d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000287 (
    .C(clk),
    .CE(ce),
    .D(sig00000469),
    .Q(sig0000047c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000288 (
    .C(clk),
    .CE(ce),
    .D(sig00000468),
    .Q(sig0000047b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000289 (
    .C(clk),
    .CE(ce),
    .D(sig00000467),
    .Q(sig0000047a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000028a (
    .C(clk),
    .CE(ce),
    .D(sig00000466),
    .Q(sig00000479)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000028b (
    .C(clk),
    .CE(ce),
    .D(sig00000465),
    .Q(sig00000474)
  );
  MUXCY   blk0000028c (
    .CI(sig00000471),
    .DI(sig00000001),
    .S(sig00000485),
    .O(sig00000472)
  );
  MUXCY   blk0000028d (
    .CI(sig00000470),
    .DI(sig00000001),
    .S(sig00000484),
    .O(sig00000471)
  );
  MUXCY   blk0000028e (
    .CI(sig0000046f),
    .DI(sig00000001),
    .S(sig00000483),
    .O(sig00000470)
  );
  MUXCY   blk0000028f (
    .CI(sig0000046e),
    .DI(sig00000001),
    .S(sig00000482),
    .O(sig0000046f)
  );
  MUXCY   blk00000290 (
    .CI(sig0000046d),
    .DI(sig00000001),
    .S(sig0000048e),
    .O(sig0000046e)
  );
  MUXCY   blk00000291 (
    .CI(sig00000002),
    .DI(sig00000001),
    .S(sig0000048d),
    .O(sig0000046d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000292 (
    .C(clk),
    .CE(ce),
    .D(sig00000472),
    .Q(sig00000478)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000293 (
    .C(clk),
    .CE(ce),
    .D(sig00000471),
    .Q(sig00000477)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000294 (
    .C(clk),
    .CE(ce),
    .D(sig00000470),
    .Q(sig00000476)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000295 (
    .C(clk),
    .CE(ce),
    .D(sig0000046f),
    .Q(sig00000475)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000296 (
    .C(clk),
    .CE(ce),
    .D(sig0000046e),
    .Q(sig00000480)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000297 (
    .C(clk),
    .CE(ce),
    .D(sig0000046d),
    .Q(sig0000047f)
  );
  MUXF5   blk00000298 (
    .I0(sig00000455),
    .I1(sig00000001),
    .S(sig00000585),
    .O(sig0000045c)
  );
  MUXF5   blk00000299 (
    .I0(sig00000454),
    .I1(sig00000458),
    .S(sig00000585),
    .O(sig0000045b)
  );
  MUXF5   blk0000029a (
    .I0(sig00000453),
    .I1(sig00000457),
    .S(sig00000585),
    .O(sig0000045a)
  );
  MUXF5   blk0000029b (
    .I0(sig00000452),
    .I1(sig00000456),
    .S(sig00000585),
    .O(sig00000459)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000029c (
    .C(clk),
    .CE(ce),
    .D(sig00000459),
    .Q(sig0000044e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000029d (
    .C(clk),
    .CE(ce),
    .D(sig0000045a),
    .Q(sig0000044f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000029e (
    .C(clk),
    .CE(ce),
    .D(sig0000045b),
    .Q(sig00000450)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000029f (
    .C(clk),
    .CE(ce),
    .D(sig0000045c),
    .Q(sig00000451)
  );
  MUXF5   blk000002a0 (
    .I0(sig00000445),
    .I1(sig00000449),
    .S(sig00000585),
    .O(sig0000044d)
  );
  MUXF5   blk000002a1 (
    .I0(sig00000444),
    .I1(sig00000448),
    .S(sig00000585),
    .O(sig0000044c)
  );
  MUXF5   blk000002a2 (
    .I0(sig00000443),
    .I1(sig00000447),
    .S(sig00000585),
    .O(sig0000044b)
  );
  MUXF5   blk000002a3 (
    .I0(sig00000442),
    .I1(sig00000446),
    .S(sig00000585),
    .O(sig0000044a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002a4 (
    .C(clk),
    .CE(ce),
    .D(sig0000044a),
    .Q(sig0000043e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002a5 (
    .C(clk),
    .CE(ce),
    .D(sig0000044b),
    .Q(sig0000043f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002a6 (
    .C(clk),
    .CE(ce),
    .D(sig0000044c),
    .Q(sig00000440)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002a7 (
    .C(clk),
    .CE(ce),
    .D(sig0000044d),
    .Q(sig00000441)
  );
  FDRSE   blk000002a8 (
    .C(clk),
    .CE(ce),
    .D(sig00000500),
    .R(sig0000059e),
    .S(sig00000001),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [10])
  );
  FDRSE   blk000002a9 (
    .C(clk),
    .CE(ce),
    .D(sig00000501),
    .R(sig0000059e),
    .S(sig00000001),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [11])
  );
  FDRSE   blk000002aa (
    .C(clk),
    .CE(ce),
    .D(sig0000052f),
    .R(sig0000059e),
    .S(sig00000001),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [12])
  );
  FDRSE   blk000002ab (
    .C(clk),
    .CE(ce),
    .D(sig00000530),
    .R(sig0000059e),
    .S(sig00000001),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [13])
  );
  FDRSE   blk000002ac (
    .C(clk),
    .CE(ce),
    .D(sig00000533),
    .R(sig0000059e),
    .S(sig00000001),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [14])
  );
  FDRSE   blk000002ad (
    .C(clk),
    .CE(ce),
    .D(sig00000539),
    .R(sig0000059e),
    .S(sig00000001),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [20])
  );
  FDRSE   blk000002ae (
    .C(clk),
    .CE(ce),
    .D(sig00000534),
    .R(sig0000059e),
    .S(sig00000001),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [15])
  );
  FDRSE   blk000002af (
    .C(clk),
    .CE(ce),
    .D(sig0000053a),
    .R(sig0000059e),
    .S(sig00000001),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [21])
  );
  FDRSE   blk000002b0 (
    .C(clk),
    .CE(ce),
    .D(sig00000535),
    .R(sig0000059e),
    .S(sig00000001),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [16])
  );
  FDRSE   blk000002b1 (
    .C(clk),
    .CE(ce),
    .D(sig00000536),
    .R(sig0000059e),
    .S(sig00000001),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [17])
  );
  FDRSE   blk000002b2 (
    .C(clk),
    .CE(ce),
    .D(sig00000531),
    .R(sig0000059f),
    .S(sig000005a0),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [22])
  );
  FDRSE   blk000002b3 (
    .C(clk),
    .CE(ce),
    .D(sig00000537),
    .R(sig0000059e),
    .S(sig00000001),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [18])
  );
  FDRSE   blk000002b4 (
    .C(clk),
    .CE(ce),
    .D(sig00000538),
    .R(sig0000059e),
    .S(sig00000001),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [19])
  );
  FDRSE   blk000002b5 (
    .C(clk),
    .CE(ce),
    .D(sig000004fe),
    .R(sig0000059e),
    .S(sig00000001),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [0])
  );
  FDRSE   blk000002b6 (
    .C(clk),
    .CE(ce),
    .D(sig000004ff),
    .R(sig0000059e),
    .S(sig00000001),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [1])
  );
  FDRSE   blk000002b7 (
    .C(clk),
    .CE(ce),
    .D(sig00000504),
    .R(sig0000059e),
    .S(sig00000001),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [4])
  );
  FDRSE   blk000002b8 (
    .C(clk),
    .CE(ce),
    .D(sig00000502),
    .R(sig0000059e),
    .S(sig00000001),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [2])
  );
  FDRSE   blk000002b9 (
    .C(clk),
    .CE(ce),
    .D(sig00000503),
    .R(sig0000059e),
    .S(sig00000001),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [3])
  );
  FDRSE   blk000002ba (
    .C(clk),
    .CE(ce),
    .D(sig00000505),
    .R(sig0000059e),
    .S(sig00000001),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [5])
  );
  FDRSE   blk000002bb (
    .C(clk),
    .CE(ce),
    .D(sig00000506),
    .R(sig0000059e),
    .S(sig00000001),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [6])
  );
  FDRSE   blk000002bc (
    .C(clk),
    .CE(ce),
    .D(sig00000507),
    .R(sig0000059e),
    .S(sig00000001),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [7])
  );
  FDRSE   blk000002bd (
    .C(clk),
    .CE(ce),
    .D(sig00000508),
    .R(sig0000059e),
    .S(sig00000001),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [8])
  );
  FDRSE   blk000002be (
    .C(clk),
    .CE(ce),
    .D(sig00000509),
    .R(sig0000059e),
    .S(sig00000001),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [9])
  );
  FDRSE   blk000002bf (
    .C(clk),
    .CE(ce),
    .D(sig000003d9),
    .R(sig00000001),
    .S(sig00000001),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/sign_op )
  );
  FDE   blk000002c0 (
    .C(clk),
    .CE(ce),
    .D(sig00000596),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/exp_op [0])
  );
  FDE   blk000002c1 (
    .C(clk),
    .CE(ce),
    .D(sig00000597),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/exp_op [1])
  );
  FDE   blk000002c2 (
    .C(clk),
    .CE(ce),
    .D(sig00000598),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/exp_op [2])
  );
  FDE   blk000002c3 (
    .C(clk),
    .CE(ce),
    .D(sig00000599),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/exp_op [3])
  );
  FDE   blk000002c4 (
    .C(clk),
    .CE(ce),
    .D(sig0000059a),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/exp_op [4])
  );
  FDE   blk000002c5 (
    .C(clk),
    .CE(ce),
    .D(sig0000059b),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/exp_op [5])
  );
  FDE   blk000002c6 (
    .C(clk),
    .CE(ce),
    .D(sig0000059c),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/exp_op [6])
  );
  FDE   blk000002c7 (
    .C(clk),
    .CE(ce),
    .D(sig0000059d),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/exp_op [7])
  );
  MUXCY   blk000002c8 (
    .CI(sig00000001),
    .DI(sig0000058e),
    .S(sig0000058d),
    .O(sig00000586)
  );
  XORCY   blk000002c9 (
    .CI(sig00000001),
    .LI(sig0000058d),
    .O(sig00000596)
  );
  MUXCY   blk000002ca (
    .CI(sig00000586),
    .DI(sig00000001),
    .S(sig0000058f),
    .O(sig00000587)
  );
  XORCY   blk000002cb (
    .CI(sig00000586),
    .LI(sig0000058f),
    .O(sig00000597)
  );
  MUXCY   blk000002cc (
    .CI(sig00000587),
    .DI(sig00000001),
    .S(sig00000590),
    .O(sig00000588)
  );
  XORCY   blk000002cd (
    .CI(sig00000587),
    .LI(sig00000590),
    .O(sig00000598)
  );
  MUXCY   blk000002ce (
    .CI(sig00000588),
    .DI(sig00000001),
    .S(sig00000591),
    .O(sig00000589)
  );
  XORCY   blk000002cf (
    .CI(sig00000588),
    .LI(sig00000591),
    .O(sig00000599)
  );
  MUXCY   blk000002d0 (
    .CI(sig00000589),
    .DI(sig00000001),
    .S(sig00000592),
    .O(sig0000058a)
  );
  XORCY   blk000002d1 (
    .CI(sig00000589),
    .LI(sig00000592),
    .O(sig0000059a)
  );
  MUXCY   blk000002d2 (
    .CI(sig0000058a),
    .DI(sig00000001),
    .S(sig00000593),
    .O(sig0000058b)
  );
  XORCY   blk000002d3 (
    .CI(sig0000058a),
    .LI(sig00000593),
    .O(sig0000059b)
  );
  MUXCY   blk000002d4 (
    .CI(sig0000058b),
    .DI(sig00000001),
    .S(sig00000594),
    .O(sig0000058c)
  );
  XORCY   blk000002d5 (
    .CI(sig0000058b),
    .LI(sig00000594),
    .O(sig0000059c)
  );
  XORCY   blk000002d6 (
    .CI(sig0000058c),
    .LI(sig00000595),
    .O(sig0000059d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002d7 (
    .C(clk),
    .CE(ce),
    .D(sig000004e7),
    .Q(sig0000048f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002d8 (
    .C(clk),
    .CE(ce),
    .D(sig000004ef),
    .Q(sig0000049a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002d9 (
    .C(clk),
    .CE(ce),
    .D(sig000004f0),
    .Q(sig000004a2)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002da (
    .C(clk),
    .CE(ce),
    .D(sig000004f1),
    .Q(sig000004a3)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002db (
    .C(clk),
    .CE(ce),
    .D(sig000004f2),
    .Q(sig000004a4)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002dc (
    .C(clk),
    .CE(ce),
    .D(sig000004f3),
    .Q(sig000004a5)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002dd (
    .C(clk),
    .CE(ce),
    .D(sig000004f4),
    .Q(sig000004a6)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002de (
    .C(clk),
    .CE(ce),
    .D(sig000004f5),
    .Q(sig000004a7)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002df (
    .C(clk),
    .CE(ce),
    .D(sig000004f6),
    .Q(sig000004a8)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002e0 (
    .C(clk),
    .CE(ce),
    .D(sig000004dd),
    .Q(sig00000490)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002e1 (
    .C(clk),
    .CE(ce),
    .D(sig000004de),
    .Q(sig00000491)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002e2 (
    .C(clk),
    .CE(ce),
    .D(sig000004df),
    .Q(sig00000492)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002e3 (
    .C(clk),
    .CE(ce),
    .D(sig000004e0),
    .Q(sig00000493)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002e4 (
    .C(clk),
    .CE(ce),
    .D(sig000004e1),
    .Q(sig00000494)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002e5 (
    .C(clk),
    .CE(ce),
    .D(sig000004e2),
    .Q(sig00000495)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002e6 (
    .C(clk),
    .CE(ce),
    .D(sig000004e3),
    .Q(sig00000496)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002e7 (
    .C(clk),
    .CE(ce),
    .D(sig000004e4),
    .Q(sig00000497)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002e8 (
    .C(clk),
    .CE(ce),
    .D(sig000004e5),
    .Q(sig00000498)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002e9 (
    .C(clk),
    .CE(ce),
    .D(sig000004e6),
    .Q(sig00000499)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002ea (
    .C(clk),
    .CE(ce),
    .D(sig000004e8),
    .Q(sig0000049b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002eb (
    .C(clk),
    .CE(ce),
    .D(sig000004e9),
    .Q(sig0000049c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002ec (
    .C(clk),
    .CE(ce),
    .D(sig000004ea),
    .Q(sig0000049d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002ed (
    .C(clk),
    .CE(ce),
    .D(sig000004eb),
    .Q(sig0000049e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002ee (
    .C(clk),
    .CE(ce),
    .D(sig000004ec),
    .Q(sig0000049f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002ef (
    .C(clk),
    .CE(ce),
    .D(sig000004ed),
    .Q(sig000004a0)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002f0 (
    .C(clk),
    .CE(ce),
    .D(sig000004ee),
    .Q(sig000004a1)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002f1 (
    .C(clk),
    .CE(ce),
    .D(sig000004cd),
    .Q(sig000004a9)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002f2 (
    .C(clk),
    .CE(ce),
    .D(sig000004d5),
    .Q(sig000004b4)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002f3 (
    .C(clk),
    .CE(ce),
    .D(sig000004d6),
    .Q(sig000004bc)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002f4 (
    .C(clk),
    .CE(ce),
    .D(sig000004d7),
    .Q(sig000004bd)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002f5 (
    .C(clk),
    .CE(ce),
    .D(sig000004d8),
    .Q(sig000004be)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002f6 (
    .C(clk),
    .CE(ce),
    .D(sig000004d9),
    .Q(sig000004bf)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002f7 (
    .C(clk),
    .CE(ce),
    .D(sig000004da),
    .Q(sig000004c0)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002f8 (
    .C(clk),
    .CE(ce),
    .D(sig000004db),
    .Q(sig000004c1)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002f9 (
    .C(clk),
    .CE(ce),
    .D(sig000004dc),
    .Q(sig000004c2)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002fa (
    .C(clk),
    .CE(ce),
    .D(sig000004c3),
    .Q(sig000004aa)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002fb (
    .C(clk),
    .CE(ce),
    .D(sig000004c4),
    .Q(sig000004ab)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002fc (
    .C(clk),
    .CE(ce),
    .D(sig000004c5),
    .Q(sig000004ac)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002fd (
    .C(clk),
    .CE(ce),
    .D(sig000004c6),
    .Q(sig000004ad)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002fe (
    .C(clk),
    .CE(ce),
    .D(sig000004c7),
    .Q(sig000004ae)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002ff (
    .C(clk),
    .CE(ce),
    .D(sig000004c8),
    .Q(sig000004af)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000300 (
    .C(clk),
    .CE(ce),
    .D(sig000004c9),
    .Q(sig000004b0)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000301 (
    .C(clk),
    .CE(ce),
    .D(sig000004ca),
    .Q(sig000004b1)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000302 (
    .C(clk),
    .CE(ce),
    .D(sig000004cb),
    .Q(sig000004b2)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000303 (
    .C(clk),
    .CE(ce),
    .D(sig000004cc),
    .Q(sig000004b3)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000304 (
    .C(clk),
    .CE(ce),
    .D(sig000004ce),
    .Q(sig000004b5)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000305 (
    .C(clk),
    .CE(ce),
    .D(sig000004cf),
    .Q(sig000004b6)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000306 (
    .C(clk),
    .CE(ce),
    .D(sig000004d0),
    .Q(sig000004b7)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000307 (
    .C(clk),
    .CE(ce),
    .D(sig000004d1),
    .Q(sig000004b8)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000308 (
    .C(clk),
    .CE(ce),
    .D(sig000004d2),
    .Q(sig000004b9)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000309 (
    .C(clk),
    .CE(ce),
    .D(sig000004d3),
    .Q(sig000004ba)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000030a (
    .C(clk),
    .CE(ce),
    .D(sig000004d4),
    .Q(sig000004bb)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000030b (
    .C(clk),
    .CE(ce),
    .D(sig000001ba),
    .Q(sig0000041f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000030c (
    .C(clk),
    .CE(ce),
    .D(sig000001bb),
    .Q(sig00000420)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000030d (
    .C(clk),
    .CE(ce),
    .D(sig000001bf),
    .Q(sig0000042b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000030e (
    .C(clk),
    .CE(ce),
    .D(sig000001c0),
    .Q(sig00000432)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000030f (
    .C(clk),
    .CE(ce),
    .D(sig000001c1),
    .Q(sig00000433)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000310 (
    .C(clk),
    .CE(ce),
    .D(sig000001c2),
    .Q(sig00000434)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000311 (
    .C(clk),
    .CE(ce),
    .D(sig000001c3),
    .Q(sig00000435)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000312 (
    .C(clk),
    .CE(ce),
    .D(sig000001c4),
    .Q(sig00000436)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000313 (
    .C(clk),
    .CE(ce),
    .D(sig000001c5),
    .Q(sig00000437)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000314 (
    .C(clk),
    .CE(ce),
    .D(sig000001c6),
    .Q(sig00000438)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000315 (
    .C(clk),
    .CE(ce),
    .D(sig000001bc),
    .Q(sig00000421)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000316 (
    .C(clk),
    .CE(ce),
    .D(sig000001bd),
    .Q(sig00000422)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000317 (
    .C(clk),
    .CE(ce),
    .D(sig000001be),
    .Q(sig00000423)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000318 (
    .C(clk),
    .CE(ce),
    .D(sig000001ff),
    .Q(sig00000424)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000319 (
    .C(clk),
    .CE(ce),
    .D(sig00000200),
    .Q(sig00000425)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000031a (
    .C(clk),
    .CE(ce),
    .D(sig00000205),
    .Q(sig00000426)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000031b (
    .C(clk),
    .CE(ce),
    .D(sig00000206),
    .Q(sig00000427)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000031c (
    .C(clk),
    .CE(ce),
    .D(sig00000207),
    .Q(sig00000428)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000031d (
    .C(clk),
    .CE(ce),
    .D(sig00000208),
    .Q(sig00000429)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000031e (
    .C(clk),
    .CE(ce),
    .D(sig00000209),
    .Q(sig0000042a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000031f (
    .C(clk),
    .CE(ce),
    .D(sig0000020a),
    .Q(sig0000042c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000320 (
    .C(clk),
    .CE(ce),
    .D(sig0000020b),
    .Q(sig0000042d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000321 (
    .C(clk),
    .CE(ce),
    .D(sig0000020c),
    .Q(sig0000042e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000322 (
    .C(clk),
    .CE(ce),
    .D(sig00000201),
    .Q(sig0000042f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000323 (
    .C(clk),
    .CE(ce),
    .D(sig00000202),
    .Q(sig00000430)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000324 (
    .C(clk),
    .CE(ce),
    .D(sig00000203),
    .Q(sig00000431)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000325 (
    .C(clk),
    .CE(ce),
    .D(a[0]),
    .Q(sig000002a2)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000326 (
    .C(clk),
    .CE(ce),
    .D(a[1]),
    .Q(sig000002a3)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000327 (
    .C(clk),
    .CE(ce),
    .D(a[2]),
    .Q(sig000002ae)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000328 (
    .C(clk),
    .CE(ce),
    .D(a[3]),
    .Q(sig000002b2)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000329 (
    .C(clk),
    .CE(ce),
    .D(a[4]),
    .Q(sig000002b3)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000032a (
    .C(clk),
    .CE(ce),
    .D(a[5]),
    .Q(sig000002b4)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000032b (
    .C(clk),
    .CE(ce),
    .D(a[6]),
    .Q(sig000002b5)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000032c (
    .C(clk),
    .CE(ce),
    .D(a[7]),
    .Q(sig000002b6)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000032d (
    .C(clk),
    .CE(ce),
    .D(a[8]),
    .Q(sig000002b7)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000032e (
    .C(clk),
    .CE(ce),
    .D(a[9]),
    .Q(sig000002b8)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000032f (
    .C(clk),
    .CE(ce),
    .D(a[10]),
    .Q(sig000002a4)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000330 (
    .C(clk),
    .CE(ce),
    .D(a[11]),
    .Q(sig000002a5)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000331 (
    .C(clk),
    .CE(ce),
    .D(a[12]),
    .Q(sig000002a6)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000332 (
    .C(clk),
    .CE(ce),
    .D(a[13]),
    .Q(sig000002a7)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000333 (
    .C(clk),
    .CE(ce),
    .D(a[14]),
    .Q(sig000002a8)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000334 (
    .C(clk),
    .CE(ce),
    .D(a[15]),
    .Q(sig000002a9)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000335 (
    .C(clk),
    .CE(ce),
    .D(a[16]),
    .Q(sig000002aa)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000336 (
    .C(clk),
    .CE(ce),
    .D(a[17]),
    .Q(sig000002ab)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000337 (
    .C(clk),
    .CE(ce),
    .D(a[18]),
    .Q(sig000002ac)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000338 (
    .C(clk),
    .CE(ce),
    .D(a[19]),
    .Q(sig000002ad)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000339 (
    .C(clk),
    .CE(ce),
    .D(a[20]),
    .Q(sig000002af)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000033a (
    .C(clk),
    .CE(ce),
    .D(a[21]),
    .Q(sig000002b0)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000033b (
    .C(clk),
    .CE(ce),
    .D(a[22]),
    .Q(sig000002b1)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000033c (
    .C(clk),
    .CE(ce),
    .D(b[0]),
    .Q(sig000002b9)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000033d (
    .C(clk),
    .CE(ce),
    .D(b[1]),
    .Q(sig000002ba)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000033e (
    .C(clk),
    .CE(ce),
    .D(b[2]),
    .Q(sig000002c5)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000033f (
    .C(clk),
    .CE(ce),
    .D(b[3]),
    .Q(sig000002c9)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000340 (
    .C(clk),
    .CE(ce),
    .D(b[4]),
    .Q(sig000002ca)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000341 (
    .C(clk),
    .CE(ce),
    .D(b[5]),
    .Q(sig000002cb)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000342 (
    .C(clk),
    .CE(ce),
    .D(b[6]),
    .Q(sig000002cc)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000343 (
    .C(clk),
    .CE(ce),
    .D(b[7]),
    .Q(sig000002cd)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000344 (
    .C(clk),
    .CE(ce),
    .D(b[8]),
    .Q(sig000002ce)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000345 (
    .C(clk),
    .CE(ce),
    .D(b[9]),
    .Q(sig000002cf)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000346 (
    .C(clk),
    .CE(ce),
    .D(b[10]),
    .Q(sig000002bb)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000347 (
    .C(clk),
    .CE(ce),
    .D(b[11]),
    .Q(sig000002bc)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000348 (
    .C(clk),
    .CE(ce),
    .D(b[12]),
    .Q(sig000002bd)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000349 (
    .C(clk),
    .CE(ce),
    .D(b[13]),
    .Q(sig000002be)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000034a (
    .C(clk),
    .CE(ce),
    .D(b[14]),
    .Q(sig000002bf)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000034b (
    .C(clk),
    .CE(ce),
    .D(b[15]),
    .Q(sig000002c0)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000034c (
    .C(clk),
    .CE(ce),
    .D(b[16]),
    .Q(sig000002c1)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000034d (
    .C(clk),
    .CE(ce),
    .D(b[17]),
    .Q(sig000002c2)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000034e (
    .C(clk),
    .CE(ce),
    .D(b[18]),
    .Q(sig000002c3)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000034f (
    .C(clk),
    .CE(ce),
    .D(b[19]),
    .Q(sig000002c4)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000350 (
    .C(clk),
    .CE(ce),
    .D(b[20]),
    .Q(sig000002c6)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000351 (
    .C(clk),
    .CE(ce),
    .D(b[21]),
    .Q(sig000002c7)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000352 (
    .C(clk),
    .CE(ce),
    .D(b[22]),
    .Q(sig000002c8)
  );
  LUT2 #(
    .INIT ( 4'h8 ))
  blk00000353 (
    .I0(sig00000450),
    .I1(sig00000451),
    .O(sig00000464)
  );
  LUT2 #(
    .INIT ( 4'h8 ))
  blk00000354 (
    .I0(sig0000044e),
    .I1(sig0000044f),
    .O(sig00000463)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000355 (
    .I0(b[31]),
    .I1(operation[0]),
    .O(sig000003e8)
  );
  LUT3 #(
    .INIT ( 8'h96 ))
  blk00000356 (
    .I0(operation[0]),
    .I1(b[31]),
    .I2(a[31]),
    .O(sig0000041e)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000357 (
    .I0(a[15]),
    .I1(b[15]),
    .O(sig0000039d)
  );
  LUT3 #(
    .INIT ( 8'h01 ))
  blk00000358 (
    .I0(b[22]),
    .I1(b[21]),
    .I2(b[20]),
    .O(sig00000314)
  );
  LUT3 #(
    .INIT ( 8'h01 ))
  blk00000359 (
    .I0(a[22]),
    .I1(a[21]),
    .I2(a[20]),
    .O(sig00000300)
  );
  LUT4 #(
    .INIT ( 16'h0001 ))
  blk0000035a (
    .I0(b[28]),
    .I1(b[27]),
    .I2(b[30]),
    .I3(b[29]),
    .O(sig00000308)
  );
  LUT4 #(
    .INIT ( 16'h8000 ))
  blk0000035b (
    .I0(b[28]),
    .I1(b[27]),
    .I2(b[30]),
    .I3(b[29]),
    .O(sig00000304)
  );
  LUT4 #(
    .INIT ( 16'h0001 ))
  blk0000035c (
    .I0(a[28]),
    .I1(a[27]),
    .I2(a[30]),
    .I3(a[29]),
    .O(sig000002f4)
  );
  LUT4 #(
    .INIT ( 16'h8000 ))
  blk0000035d (
    .I0(a[28]),
    .I1(a[27]),
    .I2(a[30]),
    .I3(a[29]),
    .O(sig000002f0)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk0000035e (
    .I0(b[30]),
    .I1(a[30]),
    .O(sig000003c5)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk0000035f (
    .I0(a[14]),
    .I1(b[14]),
    .O(sig0000039c)
  );
  LUT4 #(
    .INIT ( 16'h0001 ))
  blk00000360 (
    .I0(b[17]),
    .I1(b[16]),
    .I2(b[19]),
    .I3(b[18]),
    .O(sig00000313)
  );
  LUT4 #(
    .INIT ( 16'h0001 ))
  blk00000361 (
    .I0(b[24]),
    .I1(b[23]),
    .I2(b[26]),
    .I3(b[25]),
    .O(sig00000307)
  );
  LUT4 #(
    .INIT ( 16'h8000 ))
  blk00000362 (
    .I0(b[24]),
    .I1(b[23]),
    .I2(b[26]),
    .I3(b[25]),
    .O(sig00000303)
  );
  LUT4 #(
    .INIT ( 16'h0001 ))
  blk00000363 (
    .I0(a[17]),
    .I1(a[16]),
    .I2(a[19]),
    .I3(a[18]),
    .O(sig000002ff)
  );
  LUT4 #(
    .INIT ( 16'h0001 ))
  blk00000364 (
    .I0(a[24]),
    .I1(a[23]),
    .I2(a[26]),
    .I3(a[25]),
    .O(sig000002f3)
  );
  LUT4 #(
    .INIT ( 16'h8000 ))
  blk00000365 (
    .I0(a[24]),
    .I1(a[23]),
    .I2(a[26]),
    .I3(a[25]),
    .O(sig000002ef)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000366 (
    .I0(a[13]),
    .I1(b[13]),
    .O(sig0000039b)
  );
  LUT4 #(
    .INIT ( 16'h0001 ))
  blk00000367 (
    .I0(b[13]),
    .I1(b[12]),
    .I2(b[15]),
    .I3(b[14]),
    .O(sig00000312)
  );
  LUT4 #(
    .INIT ( 16'h0001 ))
  blk00000368 (
    .I0(a[13]),
    .I1(a[12]),
    .I2(a[15]),
    .I3(a[14]),
    .O(sig000002fe)
  );
  LUT2 #(
    .INIT ( 4'h8 ))
  blk00000369 (
    .I0(sig00000585),
    .I1(sig00000478),
    .O(sig00000473)
  );
  LUT2 #(
    .INIT ( 4'h8 ))
  blk0000036a (
    .I0(sig0000033d),
    .I1(sig0000037b),
    .O(sig0000040a)
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  blk0000036b (
    .I0(sig0000034c),
    .I1(sig0000034b),
    .O(sig000003f3)
  );
  LUT2 #(
    .INIT ( 4'h8 ))
  blk0000036c (
    .I0(sig000002d8),
    .I1(sig000002ea),
    .O(sig000003dc)
  );
  LUT2 #(
    .INIT ( 4'hE ))
  blk0000036d (
    .I0(sig000003e6),
    .I1(sig000003de),
    .O(sig000005a3)
  );
  LUT2 #(
    .INIT ( 4'hE ))
  blk0000036e (
    .I0(sig0000025b),
    .I1(sig00000260),
    .O(sig000002a1)
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  blk0000036f (
    .I0(sig0000008b),
    .I1(sig00000248),
    .O(sig0000011f)
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  blk00000370 (
    .I0(sig0000008b),
    .I1(sig00000247),
    .O(sig0000011e)
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  blk00000371 (
    .I0(sig0000008b),
    .I1(sig00000246),
    .O(sig0000011d)
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  blk00000372 (
    .I0(sig0000008b),
    .I1(sig00000245),
    .O(sig0000011c)
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  blk00000373 (
    .I0(sig0000008b),
    .I1(sig00000244),
    .O(sig0000011b)
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  blk00000374 (
    .I0(sig0000008b),
    .I1(sig00000243),
    .O(sig0000011a)
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  blk00000375 (
    .I0(sig0000008b),
    .I1(sig00000258),
    .O(sig00000119)
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  blk00000376 (
    .I0(sig0000008b),
    .I1(sig00000257),
    .O(sig00000118)
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  blk00000377 (
    .I0(sig0000008b),
    .I1(sig00000251),
    .O(sig00000128)
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  blk00000378 (
    .I0(sig0000008b),
    .I1(sig00000250),
    .O(sig00000127)
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  blk00000379 (
    .I0(sig0000008b),
    .I1(sig0000024f),
    .O(sig00000126)
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  blk0000037a (
    .I0(sig0000008b),
    .I1(sig0000024e),
    .O(sig00000125)
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  blk0000037b (
    .I0(sig0000008b),
    .I1(sig0000024c),
    .O(sig00000124)
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  blk0000037c (
    .I0(sig0000008b),
    .I1(sig0000024b),
    .O(sig00000123)
  );
  LUT2 #(
    .INIT ( 4'h8 ))
  blk0000037d (
    .I0(sig0000008b),
    .I1(sig00000248),
    .O(sig00000122)
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  blk0000037e (
    .I0(sig0000008b),
    .I1(sig0000024a),
    .O(sig00000121)
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  blk0000037f (
    .I0(sig0000008b),
    .I1(sig00000249),
    .O(sig00000120)
  );
  LUT2 #(
    .INIT ( 4'h8 ))
  blk00000380 (
    .I0(sig0000008b),
    .I1(sig00000247),
    .O(sig00000117)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000381 (
    .I0(sig000002ea),
    .I1(sig000002d8),
    .O(sig000003e3)
  );
  LUT3 #(
    .INIT ( 8'h7F ))
  blk00000382 (
    .I0(sig00000087),
    .I1(sig00000088),
    .I2(sig00000241),
    .O(sig0000015b)
  );
  LUT3 #(
    .INIT ( 8'h10 ))
  blk00000383 (
    .I0(sig000000e2),
    .I1(sig000000e1),
    .I2(sig000000bb),
    .O(sig000000f5)
  );
  LUT3 #(
    .INIT ( 8'h10 ))
  blk00000384 (
    .I0(sig000000c3),
    .I1(sig000000c4),
    .I2(sig000000a1),
    .O(sig0000010e)
  );
  LUT3 #(
    .INIT ( 8'h10 ))
  blk00000385 (
    .I0(sig000000c3),
    .I1(sig000000c4),
    .I2(sig000000a0),
    .O(sig0000010d)
  );
  LUT3 #(
    .INIT ( 8'h10 ))
  blk00000386 (
    .I0(sig000000c3),
    .I1(sig000000c4),
    .I2(sig0000009f),
    .O(sig0000010c)
  );
  LUT3 #(
    .INIT ( 8'h10 ))
  blk00000387 (
    .I0(sig000000c3),
    .I1(sig000000c4),
    .I2(sig0000009e),
    .O(sig0000010b)
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  blk00000388 (
    .I0(sig0000008b),
    .I1(sig00000256),
    .I2(sig00000251),
    .O(sig00000130)
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  blk00000389 (
    .I0(sig0000008b),
    .I1(sig00000255),
    .I2(sig00000250),
    .O(sig0000012f)
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  blk0000038a (
    .I0(sig0000008b),
    .I1(sig00000254),
    .I2(sig0000024f),
    .O(sig0000012e)
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  blk0000038b (
    .I0(sig0000008b),
    .I1(sig00000253),
    .I2(sig0000024e),
    .O(sig0000012d)
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  blk0000038c (
    .I0(sig0000008b),
    .I1(sig00000252),
    .I2(sig0000024c),
    .O(sig0000012c)
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  blk0000038d (
    .I0(sig0000008b),
    .I1(sig0000024d),
    .I2(sig0000024b),
    .O(sig0000012b)
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  blk0000038e (
    .I0(sig0000008b),
    .I1(sig00000242),
    .I2(sig0000024a),
    .O(sig0000012a)
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  blk0000038f (
    .I0(sig0000008b),
    .I1(sig00000241),
    .I2(sig00000249),
    .O(sig00000129)
  );
  LUT4 #(
    .INIT ( 16'hA8AA ))
  blk00000390 (
    .I0(sig00000346),
    .I1(sig0000034c),
    .I2(sig0000034b),
    .I3(sig000002eb),
    .O(sig0000041b)
  );
  LUT4 #(
    .INIT ( 16'h5554 ))
  blk00000391 (
    .I0(sig0000033f),
    .I1(sig00000342),
    .I2(sig00000340),
    .I3(sig0000033e),
    .O(sig000003f8)
  );
  LUT4 #(
    .INIT ( 16'h22F2 ))
  blk00000392 (
    .I0(sig000003dd),
    .I1(sig000003df),
    .I2(sig000003e5),
    .I3(sig000003e7),
    .O(sig000003e2)
  );
  LUT4 #(
    .INIT ( 16'hF888 ))
  blk00000393 (
    .I0(sig000003e5),
    .I1(sig000003e7),
    .I2(sig000003dd),
    .I3(sig000003df),
    .O(sig000003e0)
  );
  LUT4 #(
    .INIT ( 16'h8000 ))
  blk00000394 (
    .I0(sig000003e7),
    .I1(sig000003e5),
    .I2(sig000003df),
    .I3(sig000003dd),
    .O(sig000003db)
  );
  LUT4 #(
    .INIT ( 16'h151F ))
  blk00000395 (
    .I0(sig00000088),
    .I1(sig00000087),
    .I2(sig00000250),
    .I3(sig00000251),
    .O(sig00000161)
  );
  LUT4 #(
    .INIT ( 16'h0E04 ))
  blk00000396 (
    .I0(sig000000e1),
    .I1(sig000000ba),
    .I2(sig000000e2),
    .I3(sig000000bb),
    .O(sig000000f4)
  );
  LUT4 #(
    .INIT ( 16'h0E04 ))
  blk00000397 (
    .I0(sig000000c3),
    .I1(sig0000009d),
    .I2(sig000000c4),
    .I3(sig000000a1),
    .O(sig0000010a)
  );
  LUT4 #(
    .INIT ( 16'h0E04 ))
  blk00000398 (
    .I0(sig000000c3),
    .I1(sig0000009c),
    .I2(sig000000c4),
    .I3(sig000000a0),
    .O(sig00000109)
  );
  LUT4 #(
    .INIT ( 16'h0E04 ))
  blk00000399 (
    .I0(sig000000c3),
    .I1(sig0000009a),
    .I2(sig000000c4),
    .I3(sig0000009f),
    .O(sig00000107)
  );
  LUT4 #(
    .INIT ( 16'h0E04 ))
  blk0000039a (
    .I0(sig000000c3),
    .I1(sig00000099),
    .I2(sig000000c4),
    .I3(sig0000009e),
    .O(sig00000106)
  );
  LUT4 #(
    .INIT ( 16'hEC4C ))
  blk0000039b (
    .I0(sig000003df),
    .I1(sig000002ea),
    .I2(sig000003dd),
    .I3(sig000002d8),
    .O(sig000003e1)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk0000039c (
    .I0(a[12]),
    .I1(b[12]),
    .O(sig0000039a)
  );
  LUT4 #(
    .INIT ( 16'h0001 ))
  blk0000039d (
    .I0(b[9]),
    .I1(b[8]),
    .I2(b[11]),
    .I3(b[10]),
    .O(sig00000311)
  );
  LUT4 #(
    .INIT ( 16'h0001 ))
  blk0000039e (
    .I0(a[9]),
    .I1(a[8]),
    .I2(a[11]),
    .I3(a[10]),
    .O(sig000002fd)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk0000039f (
    .I0(a[11]),
    .I1(b[11]),
    .O(sig00000399)
  );
  LUT4 #(
    .INIT ( 16'h0001 ))
  blk000003a0 (
    .I0(b[5]),
    .I1(b[4]),
    .I2(b[7]),
    .I3(b[6]),
    .O(sig00000310)
  );
  LUT4 #(
    .INIT ( 16'h0001 ))
  blk000003a1 (
    .I0(a[5]),
    .I1(a[4]),
    .I2(a[7]),
    .I3(a[6]),
    .O(sig000002fc)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk000003a2 (
    .I0(a[10]),
    .I1(b[10]),
    .O(sig00000398)
  );
  LUT4 #(
    .INIT ( 16'h0001 ))
  blk000003a3 (
    .I0(b[1]),
    .I1(b[0]),
    .I2(b[3]),
    .I3(b[2]),
    .O(sig0000030f)
  );
  LUT4 #(
    .INIT ( 16'h0001 ))
  blk000003a4 (
    .I0(a[1]),
    .I1(a[0]),
    .I2(a[3]),
    .I3(a[2]),
    .O(sig000002fb)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk000003a5 (
    .I0(a[9]),
    .I1(b[9]),
    .O(sig000003a6)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk000003a6 (
    .I0(a[8]),
    .I1(b[8]),
    .O(sig000003a5)
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  blk000003a7 (
    .I0(sig00000476),
    .I1(sig00000475),
    .O(sig00000458)
  );
  LUT2 #(
    .INIT ( 4'h8 ))
  blk000003a8 (
    .I0(sig0000047b),
    .I1(sig00000585),
    .O(sig00000455)
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  blk000003a9 (
    .I0(sig00000476),
    .I1(sig00000433),
    .O(sig00000449)
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  blk000003aa (
    .I0(sig00000476),
    .I1(sig00000435),
    .O(sig00000448)
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  blk000003ab (
    .I0(sig00000450),
    .I1(sig00000440),
    .I2(sig00000441),
    .O(sig00000461)
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  blk000003ac (
    .I0(sig0000044e),
    .I1(sig0000043e),
    .I2(sig0000043f),
    .O(sig00000460)
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  blk000003ad (
    .I0(sig00000476),
    .I1(sig00000480),
    .I2(sig00000478),
    .O(sig00000457)
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  blk000003ae (
    .I0(sig00000476),
    .I1(sig0000047f),
    .I2(sig00000477),
    .O(sig00000456)
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  blk000003af (
    .I0(sig0000047b),
    .I1(sig0000047a),
    .I2(sig0000047e),
    .O(sig00000454)
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  blk000003b0 (
    .I0(sig0000047b),
    .I1(sig00000479),
    .I2(sig0000047d),
    .O(sig00000453)
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  blk000003b1 (
    .I0(sig0000047b),
    .I1(sig00000474),
    .I2(sig0000047c),
    .O(sig00000452)
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  blk000003b2 (
    .I0(sig00000476),
    .I1(sig00000437),
    .I2(sig0000041f),
    .O(sig00000447)
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  blk000003b3 (
    .I0(sig00000476),
    .I1(sig00000421),
    .I2(sig0000042b),
    .O(sig00000446)
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  blk000003b4 (
    .I0(sig0000047b),
    .I1(sig0000042c),
    .I2(sig00000423),
    .O(sig00000445)
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  blk000003b5 (
    .I0(sig0000047b),
    .I1(sig0000042e),
    .I2(sig00000425),
    .O(sig00000444)
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  blk000003b6 (
    .I0(sig0000047b),
    .I1(sig00000430),
    .I2(sig00000427),
    .O(sig00000443)
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  blk000003b7 (
    .I0(sig0000047b),
    .I1(sig0000037a),
    .I2(sig00000429),
    .O(sig00000442)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk000003b8 (
    .I0(a[7]),
    .I1(b[7]),
    .O(sig000003a4)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk000003b9 (
    .I0(a[6]),
    .I1(b[6]),
    .O(sig000003a3)
  );
  LUT4 #(
    .INIT ( 16'hFFFE ))
  blk000003ba (
    .I0(sig0000008e),
    .I1(sig0000008d),
    .I2(sig0000008c),
    .I3(sig0000002e),
    .O(sig000002a0)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk000003bb (
    .I0(a[5]),
    .I1(b[5]),
    .O(sig000003a2)
  );
  LUT2 #(
    .INIT ( 4'h1 ))
  blk000003bc (
    .I0(sig000001be),
    .I1(sig000001bd),
    .O(sig0000048c)
  );
  LUT2 #(
    .INIT ( 4'h1 ))
  blk000003bd (
    .I0(sig00000250),
    .I1(sig00000251),
    .O(sig0000013e)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk000003be (
    .I0(a[4]),
    .I1(b[4]),
    .O(sig000003a1)
  );
  LUT2 #(
    .INIT ( 4'h1 ))
  blk000003bf (
    .I0(sig00000200),
    .I1(sig000001ff),
    .O(sig0000048b)
  );
  LUT2 #(
    .INIT ( 4'h1 ))
  blk000003c0 (
    .I0(sig000001bf),
    .I1(sig000001bb),
    .O(sig00000484)
  );
  LUT4 #(
    .INIT ( 16'h0001 ))
  blk000003c1 (
    .I0(sig0000024c),
    .I1(sig0000024b),
    .I2(sig0000024f),
    .I3(sig0000024e),
    .O(sig0000013d)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk000003c2 (
    .I0(sig000002e1),
    .I1(sig000002e0),
    .O(sig00000268)
  );
  LUT3 #(
    .INIT ( 8'h32 ))
  blk000003c3 (
    .I0(sig00000315),
    .I1(sig00000316),
    .I2(sig00000356),
    .O(sig00000595)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk000003c4 (
    .I0(a[3]),
    .I1(b[3]),
    .O(sig000003a0)
  );
  LUT2 #(
    .INIT ( 4'h1 ))
  blk000003c5 (
    .I0(sig00000206),
    .I1(sig00000205),
    .O(sig0000048a)
  );
  LUT2 #(
    .INIT ( 4'h1 ))
  blk000003c6 (
    .I0(sig000001c1),
    .I1(sig000001c0),
    .O(sig00000483)
  );
  LUT4 #(
    .INIT ( 16'h0001 ))
  blk000003c7 (
    .I0(sig00000248),
    .I1(sig00000247),
    .I2(sig0000024a),
    .I3(sig00000249),
    .O(sig0000013c)
  );
  LUT2 #(
    .INIT ( 4'h8 ))
  blk000003c8 (
    .I0(sig00000317),
    .I1(ce),
    .O(sig000005a0)
  );
  LUT2 #(
    .INIT ( 4'h8 ))
  blk000003c9 (
    .I0(sig00000318),
    .I1(ce),
    .O(sig0000059f)
  );
  LUT2 #(
    .INIT ( 4'h8 ))
  blk000003ca (
    .I0(sig00000319),
    .I1(ce),
    .O(sig0000059e)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk000003cb (
    .I0(a[2]),
    .I1(b[2]),
    .O(sig0000039f)
  );
  LUT2 #(
    .INIT ( 4'h1 ))
  blk000003cc (
    .I0(sig00000208),
    .I1(sig00000207),
    .O(sig00000489)
  );
  LUT2 #(
    .INIT ( 4'h1 ))
  blk000003cd (
    .I0(sig000001c3),
    .I1(sig000001c2),
    .O(sig00000482)
  );
  LUT4 #(
    .INIT ( 16'h0001 ))
  blk000003ce (
    .I0(sig00000244),
    .I1(sig00000243),
    .I2(sig00000246),
    .I3(sig00000245),
    .O(sig0000013b)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk000003cf (
    .I0(a[1]),
    .I1(b[1]),
    .O(sig0000039e)
  );
  LUT2 #(
    .INIT ( 4'h1 ))
  blk000003d0 (
    .I0(sig000001c5),
    .I1(sig000001c4),
    .O(sig0000048e)
  );
  LUT2 #(
    .INIT ( 4'h1 ))
  blk000003d1 (
    .I0(sig0000020a),
    .I1(sig00000209),
    .O(sig00000488)
  );
  LUT4 #(
    .INIT ( 16'h0001 ))
  blk000003d2 (
    .I0(sig00000256),
    .I1(sig00000255),
    .I2(sig00000258),
    .I3(sig00000257),
    .O(sig0000013a)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk000003d3 (
    .I0(a[0]),
    .I1(b[0]),
    .O(sig00000397)
  );
  LUT2 #(
    .INIT ( 4'h1 ))
  blk000003d4 (
    .I0(sig000001bc),
    .I1(sig000001c6),
    .O(sig0000048d)
  );
  LUT2 #(
    .INIT ( 4'h1 ))
  blk000003d5 (
    .I0(sig0000020c),
    .I1(sig0000020b),
    .O(sig00000487)
  );
  LUT4 #(
    .INIT ( 16'h0001 ))
  blk000003d6 (
    .I0(sig00000252),
    .I1(sig0000024d),
    .I2(sig00000254),
    .I3(sig00000253),
    .O(sig00000139)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk000003d7 (
    .I0(b[29]),
    .I1(a[29]),
    .O(sig000003c4)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk000003d8 (
    .I0(b[28]),
    .I1(a[28]),
    .O(sig000003c3)
  );
  LUT2 #(
    .INIT ( 4'h1 ))
  blk000003d9 (
    .I0(sig00000202),
    .I1(sig00000201),
    .O(sig00000486)
  );
  LUT2 #(
    .INIT ( 4'h1 ))
  blk000003da (
    .I0(sig00000241),
    .I1(sig00000242),
    .O(sig00000138)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk000003db (
    .I0(b[27]),
    .I1(a[27]),
    .O(sig000003c1)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk000003dc (
    .I0(b[26]),
    .I1(a[26]),
    .O(sig000003c0)
  );
  LUT2 #(
    .INIT ( 4'h1 ))
  blk000003dd (
    .I0(sig00000204),
    .I1(sig00000203),
    .O(sig00000481)
  );
  LUT2 #(
    .INIT ( 4'h8 ))
  blk000003de (
    .I0(sig000003e6),
    .I1(sig000003de),
    .O(sig000005a2)
  );
  LUT3 #(
    .INIT ( 8'h32 ))
  blk000003df (
    .I0(sig0000034c),
    .I1(sig0000034b),
    .I2(sig00000358),
    .O(sig000003f2)
  );
  LUT3 #(
    .INIT ( 8'hAC ))
  blk000003e0 (
    .I0(sig00000450),
    .I1(sig0000044e),
    .I2(sig0000044f),
    .O(sig00000583)
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  blk000003e1 (
    .I0(sig00000585),
    .I1(sig0000047b),
    .I2(sig00000476),
    .O(sig00000584)
  );
  LUT3 #(
    .INIT ( 8'hAC ))
  blk000003e2 (
    .I0(sig000002ea),
    .I1(sig000002d8),
    .I2(sig00000047),
    .O(sig0000041a)
  );
  LUT3 #(
    .INIT ( 8'hAC ))
  blk000003e3 (
    .I0(sig000002b8),
    .I1(sig000002cf),
    .I2(sig000005a1),
    .O(sig0000029f)
  );
  LUT3 #(
    .INIT ( 8'hAC ))
  blk000003e4 (
    .I0(sig000002b7),
    .I1(sig000002ce),
    .I2(sig000005a1),
    .O(sig0000029e)
  );
  LUT3 #(
    .INIT ( 8'hAC ))
  blk000003e5 (
    .I0(sig000002b6),
    .I1(sig000002cd),
    .I2(sig000005a1),
    .O(sig0000029d)
  );
  LUT3 #(
    .INIT ( 8'hAC ))
  blk000003e6 (
    .I0(sig000002b5),
    .I1(sig000002cc),
    .I2(sig000005a1),
    .O(sig0000029c)
  );
  LUT3 #(
    .INIT ( 8'hAC ))
  blk000003e7 (
    .I0(sig000002b4),
    .I1(sig000002cb),
    .I2(sig000005a1),
    .O(sig0000029b)
  );
  LUT3 #(
    .INIT ( 8'hAC ))
  blk000003e8 (
    .I0(sig000002b3),
    .I1(sig000002ca),
    .I2(sig000005a1),
    .O(sig0000029a)
  );
  LUT3 #(
    .INIT ( 8'hAC ))
  blk000003e9 (
    .I0(sig000002b2),
    .I1(sig000002c9),
    .I2(sig000005a1),
    .O(sig00000299)
  );
  LUT3 #(
    .INIT ( 8'hAC ))
  blk000003ea (
    .I0(sig000002ae),
    .I1(sig000002c5),
    .I2(sig000005a1),
    .O(sig00000298)
  );
  LUT3 #(
    .INIT ( 8'hAC ))
  blk000003eb (
    .I0(sig000002b1),
    .I1(sig000002c8),
    .I2(sig000005a1),
    .O(sig00000297)
  );
  LUT3 #(
    .INIT ( 8'hAC ))
  blk000003ec (
    .I0(sig000002b0),
    .I1(sig000002c7),
    .I2(sig000005a1),
    .O(sig00000296)
  );
  LUT3 #(
    .INIT ( 8'hAC ))
  blk000003ed (
    .I0(sig000002af),
    .I1(sig000002c6),
    .I2(sig000005a1),
    .O(sig00000295)
  );
  LUT3 #(
    .INIT ( 8'hAC ))
  blk000003ee (
    .I0(sig000002a3),
    .I1(sig000002ba),
    .I2(sig000005a1),
    .O(sig00000294)
  );
  LUT3 #(
    .INIT ( 8'hAC ))
  blk000003ef (
    .I0(sig000002ad),
    .I1(sig000002c4),
    .I2(sig000005a1),
    .O(sig00000293)
  );
  LUT3 #(
    .INIT ( 8'hAC ))
  blk000003f0 (
    .I0(sig000002ac),
    .I1(sig000002c3),
    .I2(sig000005a1),
    .O(sig00000292)
  );
  LUT3 #(
    .INIT ( 8'hAC ))
  blk000003f1 (
    .I0(sig000002ab),
    .I1(sig000002c2),
    .I2(sig000005a1),
    .O(sig00000291)
  );
  LUT3 #(
    .INIT ( 8'hAC ))
  blk000003f2 (
    .I0(sig000002aa),
    .I1(sig000002c1),
    .I2(sig000005a1),
    .O(sig00000290)
  );
  LUT3 #(
    .INIT ( 8'hAC ))
  blk000003f3 (
    .I0(sig000002a9),
    .I1(sig000002c0),
    .I2(sig000005a1),
    .O(sig0000028f)
  );
  LUT3 #(
    .INIT ( 8'hAC ))
  blk000003f4 (
    .I0(sig000002a8),
    .I1(sig000002bf),
    .I2(sig000005a1),
    .O(sig0000028e)
  );
  LUT3 #(
    .INIT ( 8'hAC ))
  blk000003f5 (
    .I0(sig000002a7),
    .I1(sig000002be),
    .I2(sig000005a1),
    .O(sig0000028d)
  );
  LUT3 #(
    .INIT ( 8'hAC ))
  blk000003f6 (
    .I0(sig000002a6),
    .I1(sig000002bd),
    .I2(sig000005a1),
    .O(sig0000028c)
  );
  LUT3 #(
    .INIT ( 8'hAC ))
  blk000003f7 (
    .I0(sig000002a5),
    .I1(sig000002bc),
    .I2(sig000005a1),
    .O(sig0000028b)
  );
  LUT3 #(
    .INIT ( 8'hAC ))
  blk000003f8 (
    .I0(sig000002a4),
    .I1(sig000002bb),
    .I2(sig000005a1),
    .O(sig0000028a)
  );
  LUT3 #(
    .INIT ( 8'hAC ))
  blk000003f9 (
    .I0(sig000002a2),
    .I1(sig000002b9),
    .I2(sig000005a1),
    .O(sig00000289)
  );
  LUT4 #(
    .INIT ( 16'hFF04 ))
  blk000003fa (
    .I0(sig00000048),
    .I1(sig0000037d),
    .I2(sig0000034c),
    .I3(sig0000034b),
    .O(sig0000041c)
  );
  LUT4 #(
    .INIT ( 16'hFFFE ))
  blk000003fb (
    .I0(sig0000034c),
    .I1(sig0000034b),
    .I2(sig00000358),
    .I3(sig0000037d),
    .O(sig00000357)
  );
  LUT4 #(
    .INIT ( 16'h00AC ))
  blk000003fc (
    .I0(sig000002cf),
    .I1(sig000002b8),
    .I2(sig000005a1),
    .I3(sig000005a2),
    .O(sig00000288)
  );
  LUT4 #(
    .INIT ( 16'h00AC ))
  blk000003fd (
    .I0(sig000002ce),
    .I1(sig000002b7),
    .I2(sig000005a1),
    .I3(sig000005a2),
    .O(sig00000287)
  );
  LUT4 #(
    .INIT ( 16'h00AC ))
  blk000003fe (
    .I0(sig000002cd),
    .I1(sig000002b6),
    .I2(sig000005a1),
    .I3(sig000005a2),
    .O(sig00000286)
  );
  LUT4 #(
    .INIT ( 16'h00AC ))
  blk000003ff (
    .I0(sig000002cc),
    .I1(sig000002b5),
    .I2(sig000005a1),
    .I3(sig000005a2),
    .O(sig00000285)
  );
  LUT4 #(
    .INIT ( 16'h00AC ))
  blk00000400 (
    .I0(sig000002cb),
    .I1(sig000002b4),
    .I2(sig000005a1),
    .I3(sig000005a2),
    .O(sig00000284)
  );
  LUT4 #(
    .INIT ( 16'h00AC ))
  blk00000401 (
    .I0(sig000002ca),
    .I1(sig000002b3),
    .I2(sig000005a1),
    .I3(sig000005a2),
    .O(sig00000283)
  );
  LUT4 #(
    .INIT ( 16'h00AC ))
  blk00000402 (
    .I0(sig000002c9),
    .I1(sig000002b2),
    .I2(sig000005a1),
    .I3(sig000005a2),
    .O(sig00000282)
  );
  LUT4 #(
    .INIT ( 16'h00AC ))
  blk00000403 (
    .I0(sig000002c5),
    .I1(sig000002ae),
    .I2(sig000005a1),
    .I3(sig000005a2),
    .O(sig00000281)
  );
  LUT4 #(
    .INIT ( 16'h00AC ))
  blk00000404 (
    .I0(sig000002c8),
    .I1(sig000002b1),
    .I2(sig000005a1),
    .I3(sig000005a2),
    .O(sig0000027f)
  );
  LUT4 #(
    .INIT ( 16'h00AC ))
  blk00000405 (
    .I0(sig000002c7),
    .I1(sig000002b0),
    .I2(sig000005a1),
    .I3(sig000005a2),
    .O(sig0000027e)
  );
  LUT4 #(
    .INIT ( 16'h00AC ))
  blk00000406 (
    .I0(sig000002c6),
    .I1(sig000002af),
    .I2(sig000005a1),
    .I3(sig000005a2),
    .O(sig0000027d)
  );
  LUT4 #(
    .INIT ( 16'h00AC ))
  blk00000407 (
    .I0(sig000002ba),
    .I1(sig000002a3),
    .I2(sig000005a1),
    .I3(sig000005a2),
    .O(sig0000027c)
  );
  LUT4 #(
    .INIT ( 16'h00AC ))
  blk00000408 (
    .I0(sig000002c4),
    .I1(sig000002ad),
    .I2(sig000005a1),
    .I3(sig000005a2),
    .O(sig0000027b)
  );
  LUT4 #(
    .INIT ( 16'h00AC ))
  blk00000409 (
    .I0(sig000002c3),
    .I1(sig000002ac),
    .I2(sig000005a1),
    .I3(sig000005a2),
    .O(sig0000027a)
  );
  LUT4 #(
    .INIT ( 16'h00AC ))
  blk0000040a (
    .I0(sig000002c2),
    .I1(sig000002ab),
    .I2(sig000005a1),
    .I3(sig000005a2),
    .O(sig00000279)
  );
  LUT4 #(
    .INIT ( 16'h00AC ))
  blk0000040b (
    .I0(sig000002c1),
    .I1(sig000002aa),
    .I2(sig000005a1),
    .I3(sig000005a2),
    .O(sig00000278)
  );
  LUT4 #(
    .INIT ( 16'h00AC ))
  blk0000040c (
    .I0(sig000002c0),
    .I1(sig000002a9),
    .I2(sig000005a1),
    .I3(sig000005a2),
    .O(sig00000277)
  );
  LUT4 #(
    .INIT ( 16'h00AC ))
  blk0000040d (
    .I0(sig000002bf),
    .I1(sig000002a8),
    .I2(sig000005a1),
    .I3(sig000005a2),
    .O(sig00000276)
  );
  LUT4 #(
    .INIT ( 16'h00AC ))
  blk0000040e (
    .I0(sig000002be),
    .I1(sig000002a7),
    .I2(sig000005a1),
    .I3(sig000005a2),
    .O(sig00000275)
  );
  LUT4 #(
    .INIT ( 16'h00AC ))
  blk0000040f (
    .I0(sig000002bd),
    .I1(sig000002a6),
    .I2(sig000005a1),
    .I3(sig000005a2),
    .O(sig00000274)
  );
  LUT4 #(
    .INIT ( 16'h00AC ))
  blk00000410 (
    .I0(sig000002bc),
    .I1(sig000002a5),
    .I2(sig000005a1),
    .I3(sig000005a2),
    .O(sig00000273)
  );
  LUT4 #(
    .INIT ( 16'h00AC ))
  blk00000411 (
    .I0(sig000002bb),
    .I1(sig000002a4),
    .I2(sig000005a1),
    .I3(sig000005a2),
    .O(sig00000272)
  );
  LUT4 #(
    .INIT ( 16'h00AC ))
  blk00000412 (
    .I0(sig000002b9),
    .I1(sig000002a2),
    .I2(sig000005a1),
    .I3(sig000005a2),
    .O(sig00000271)
  );
  LUT4 #(
    .INIT ( 16'hFF32 ))
  blk00000413 (
    .I0(sig0000037d),
    .I1(sig0000034b),
    .I2(sig00000358),
    .I3(sig0000034c),
    .O(sig0000041d)
  );
  LUT3 #(
    .INIT ( 8'hF4 ))
  blk00000414 (
    .I0(sig00000342),
    .I1(sig00000070),
    .I2(sig0000033f),
    .O(sig000003f9)
  );
  LUT4 #(
    .INIT ( 16'h085D ))
  blk00000415 (
    .I0(sig000000e2),
    .I1(sig000000bb),
    .I2(sig000000e1),
    .I3(sig00000050),
    .O(sig000000f3)
  );
  LUT4 #(
    .INIT ( 16'h085D ))
  blk00000416 (
    .I0(sig000000c4),
    .I1(sig000000a0),
    .I2(sig000000c3),
    .I3(sig00000065),
    .O(sig00000104)
  );
  LUT4 #(
    .INIT ( 16'h085D ))
  blk00000417 (
    .I0(sig000000c4),
    .I1(sig0000009f),
    .I2(sig000000c3),
    .I3(sig0000006d),
    .O(sig00000103)
  );
  LUT4 #(
    .INIT ( 16'h085D ))
  blk00000418 (
    .I0(sig000000c4),
    .I1(sig0000009e),
    .I2(sig000000c3),
    .I3(sig0000006e),
    .O(sig00000102)
  );
  LUT4 #(
    .INIT ( 16'h085D ))
  blk00000419 (
    .I0(sig000000c4),
    .I1(sig000000a1),
    .I2(sig000000c3),
    .I3(sig0000006f),
    .O(sig00000105)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk0000041a (
    .I0(sig00000498),
    .I1(sig0000049d),
    .I2(sig0000044f),
    .O(sig00000072)
  );
  LUT3 #(
    .INIT ( 8'hAC ))
  blk0000041b (
    .I0(sig00000072),
    .I1(sig00000071),
    .I2(sig00000583),
    .O(sig000004c9)
  );
  LUT3 #(
    .INIT ( 8'hAC ))
  blk0000041c (
    .I0(sig0000004b),
    .I1(sig00000073),
    .I2(sig00000583),
    .O(sig000004c8)
  );
  LUT3 #(
    .INIT ( 8'hAC ))
  blk0000041d (
    .I0(sig00000049),
    .I1(sig00000075),
    .I2(sig00000583),
    .O(sig000004c7)
  );
  LUT3 #(
    .INIT ( 8'hAC ))
  blk0000041e (
    .I0(sig0000004a),
    .I1(sig00000076),
    .I2(sig00000583),
    .O(sig000004c6)
  );
  LUT3 #(
    .INIT ( 8'hAC ))
  blk0000041f (
    .I0(sig0000004c),
    .I1(sig00000077),
    .I2(sig00000583),
    .O(sig000004c5)
  );
  LUT3 #(
    .INIT ( 8'hAC ))
  blk00000420 (
    .I0(sig0000004d),
    .I1(sig00000078),
    .I2(sig00000583),
    .O(sig000004c4)
  );
  LUT3 #(
    .INIT ( 8'hAC ))
  blk00000421 (
    .I0(sig0000004f),
    .I1(sig00000079),
    .I2(sig00000583),
    .O(sig000004dc)
  );
  LUT3 #(
    .INIT ( 8'hAC ))
  blk00000422 (
    .I0(sig00000053),
    .I1(sig0000007a),
    .I2(sig00000583),
    .O(sig000004db)
  );
  LUT3 #(
    .INIT ( 8'hAC ))
  blk00000423 (
    .I0(sig0000004e),
    .I1(sig0000007b),
    .I2(sig00000583),
    .O(sig000004c3)
  );
  LUT3 #(
    .INIT ( 8'hAC ))
  blk00000424 (
    .I0(sig00000051),
    .I1(sig0000007c),
    .I2(sig00000583),
    .O(sig000004da)
  );
  LUT3 #(
    .INIT ( 8'hAC ))
  blk00000425 (
    .I0(sig00000052),
    .I1(sig0000007d),
    .I2(sig00000583),
    .O(sig000004d9)
  );
  LUT3 #(
    .INIT ( 8'hAC ))
  blk00000426 (
    .I0(sig00000054),
    .I1(sig0000007e),
    .I2(sig00000583),
    .O(sig000004d8)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000427 (
    .I0(sig000004a3),
    .I1(sig000004a7),
    .I2(sig0000044f),
    .O(sig0000007f)
  );
  LUT3 #(
    .INIT ( 8'hAC ))
  blk00000428 (
    .I0(sig00000055),
    .I1(sig0000007f),
    .I2(sig00000583),
    .O(sig000004d7)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000429 (
    .I0(sig000004a2),
    .I1(sig000004a6),
    .I2(sig0000044f),
    .O(sig00000080)
  );
  LUT3 #(
    .INIT ( 8'hAC ))
  blk0000042a (
    .I0(sig00000056),
    .I1(sig00000080),
    .I2(sig00000583),
    .O(sig000004d6)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk0000042b (
    .I0(sig00000081),
    .I1(sig0000007f),
    .I2(sig00000583),
    .O(sig000004d5)
  );
  LUT3 #(
    .INIT ( 8'hAC ))
  blk0000042c (
    .I0(sig00000083),
    .I1(sig00000082),
    .I2(sig00000583),
    .O(sig000004ce)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk0000042d (
    .I0(sig0000048f),
    .I1(sig000004a4),
    .I2(sig0000044f),
    .O(sig00000084)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk0000042e (
    .I0(sig00000084),
    .I1(sig00000080),
    .I2(sig00000583),
    .O(sig000004cd)
  );
  LUT3 #(
    .INIT ( 8'hAC ))
  blk0000042f (
    .I0(sig00000086),
    .I1(sig00000085),
    .I2(sig00000583),
    .O(sig000004cc)
  );
  LUT3 #(
    .INIT ( 8'hAC ))
  blk00000430 (
    .I0(sig00000057),
    .I1(sig00000072),
    .I2(sig00000583),
    .O(sig000004cb)
  );
  LUT3 #(
    .INIT ( 8'hAC ))
  blk00000431 (
    .I0(sig00000058),
    .I1(sig00000074),
    .I2(sig00000583),
    .O(sig000004ca)
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  blk00000432 (
    .I0(sig000000e2),
    .I1(sig00000059),
    .I2(sig00000004),
    .O(sig000000fc)
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  blk00000433 (
    .I0(sig000000e2),
    .I1(sig0000005b),
    .I2(sig00000006),
    .O(sig000000fb)
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  blk00000434 (
    .I0(sig000000e2),
    .I1(sig00000007),
    .I2(sig00000008),
    .O(sig000000e3)
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  blk00000435 (
    .I0(sig000000e2),
    .I1(sig0000005e),
    .I2(sig00000003),
    .O(sig000000fa)
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  blk00000436 (
    .I0(sig000000e2),
    .I1(sig0000005f),
    .I2(sig00000005),
    .O(sig000000f9)
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  blk00000437 (
    .I0(sig000000e2),
    .I1(sig00000060),
    .I2(sig00000009),
    .O(sig000000f8)
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  blk00000438 (
    .I0(sig000000e2),
    .I1(sig00000061),
    .I2(sig0000000a),
    .O(sig000000f7)
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  blk00000439 (
    .I0(sig000000e2),
    .I1(sig00000062),
    .I2(sig0000000b),
    .O(sig000000f6)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk0000043a (
    .I0(sig000000b8),
    .I1(sig000000b9),
    .I2(sig000000e1),
    .O(sig0000000e)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk0000043b (
    .I0(sig000000e2),
    .I1(sig0000000f),
    .I2(sig0000000e),
    .O(sig000000f2)
  );
  LUT3 #(
    .INIT ( 8'hAC ))
  blk0000043c (
    .I0(sig000000b8),
    .I1(sig000000b7),
    .I2(sig000000e1),
    .O(sig00000010)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk0000043d (
    .I0(sig000000e2),
    .I1(sig00000011),
    .I2(sig00000010),
    .O(sig000000f1)
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  blk0000043e (
    .I0(sig000000e2),
    .I1(sig00000063),
    .I2(sig0000000e),
    .O(sig000000f0)
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  blk0000043f (
    .I0(sig000000e2),
    .I1(sig0000005d),
    .I2(sig0000000c),
    .O(sig000000ef)
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  blk00000440 (
    .I0(sig000000e2),
    .I1(sig00000064),
    .I2(sig00000010),
    .O(sig000000ee)
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  blk00000441 (
    .I0(sig000000e2),
    .I1(sig00000066),
    .I2(sig00000012),
    .O(sig000000ed)
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  blk00000442 (
    .I0(sig000000e2),
    .I1(sig00000067),
    .I2(sig00000013),
    .O(sig000000ec)
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  blk00000443 (
    .I0(sig000000e2),
    .I1(sig00000068),
    .I2(sig00000014),
    .O(sig000000eb)
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  blk00000444 (
    .I0(sig000000e2),
    .I1(sig00000069),
    .I2(sig00000015),
    .O(sig000000ea)
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  blk00000445 (
    .I0(sig000000e2),
    .I1(sig0000006a),
    .I2(sig00000016),
    .O(sig000000e9)
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  blk00000446 (
    .I0(sig000000e2),
    .I1(sig0000006b),
    .I2(sig00000017),
    .O(sig000000e8)
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  blk00000447 (
    .I0(sig000000e2),
    .I1(sig0000006c),
    .I2(sig00000018),
    .O(sig000000e7)
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  blk00000448 (
    .I0(sig000000e2),
    .I1(sig0000005a),
    .I2(sig00000019),
    .O(sig000000e6)
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  blk00000449 (
    .I0(sig000000e2),
    .I1(sig0000005c),
    .I2(sig0000001a),
    .O(sig000000e5)
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  blk0000044a (
    .I0(sig000000e2),
    .I1(sig0000001b),
    .I2(sig0000000d),
    .O(sig000000e4)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk0000044b (
    .I0(sig00000094),
    .I1(sig00000098),
    .I2(sig000000c3),
    .O(sig0000001c)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk0000044c (
    .I0(sig000000c4),
    .I1(sig0000001d),
    .I2(sig0000001c),
    .O(sig00000101)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk0000044d (
    .I0(sig00000093),
    .I1(sig00000097),
    .I2(sig000000c3),
    .O(sig0000001e)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk0000044e (
    .I0(sig000000c4),
    .I1(sig0000001f),
    .I2(sig0000001e),
    .O(sig00000100)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk0000044f (
    .I0(sig00000092),
    .I1(sig00000096),
    .I2(sig000000c3),
    .O(sig00000020)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk00000450 (
    .I0(sig000000c4),
    .I1(sig00000021),
    .I2(sig00000020),
    .O(sig000000ff)
  );
  LUT3 #(
    .INIT ( 8'hAC ))
  blk00000451 (
    .I0(sig00000094),
    .I1(sig000000a8),
    .I2(sig000000c3),
    .O(sig00000022)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk00000452 (
    .I0(sig000000c4),
    .I1(sig00000023),
    .I2(sig00000022),
    .O(sig00000116)
  );
  LUT3 #(
    .INIT ( 8'hAC ))
  blk00000453 (
    .I0(sig00000093),
    .I1(sig000000a7),
    .I2(sig000000c3),
    .O(sig00000024)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk00000454 (
    .I0(sig000000c4),
    .I1(sig00000025),
    .I2(sig00000024),
    .O(sig00000115)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000455 (
    .I0(sig00000096),
    .I1(sig0000009a),
    .I2(sig000000c3),
    .O(sig00000027)
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  blk00000456 (
    .I0(sig000000c4),
    .I1(sig00000026),
    .I2(sig00000027),
    .O(sig00000114)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000457 (
    .I0(sig00000095),
    .I1(sig00000099),
    .I2(sig000000c3),
    .O(sig00000029)
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  blk00000458 (
    .I0(sig000000c4),
    .I1(sig00000028),
    .I2(sig00000029),
    .O(sig00000113)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000459 (
    .I0(sig00000091),
    .I1(sig00000095),
    .I2(sig000000c3),
    .O(sig0000002a)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk0000045a (
    .I0(sig000000c4),
    .I1(sig0000002b),
    .I2(sig0000002a),
    .O(sig000000fe)
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  blk0000045b (
    .I0(sig000000c4),
    .I1(sig0000002c),
    .I2(sig0000001c),
    .O(sig00000112)
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  blk0000045c (
    .I0(sig000000c4),
    .I1(sig0000002d),
    .I2(sig0000001e),
    .O(sig00000111)
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  blk0000045d (
    .I0(sig000000c4),
    .I1(sig0000002f),
    .I2(sig00000020),
    .O(sig00000110)
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  blk0000045e (
    .I0(sig000000c4),
    .I1(sig00000030),
    .I2(sig0000002a),
    .O(sig0000010f)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk0000045f (
    .I0(sig0000008f),
    .I1(sig000000a3),
    .I2(sig000000c3),
    .O(sig00000031)
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  blk00000460 (
    .I0(sig000000c4),
    .I1(sig00000031),
    .I2(sig00000024),
    .O(sig000000fd)
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  blk00000461 (
    .I0(sig000000c4),
    .I1(sig00000032),
    .I2(sig00000022),
    .O(sig00000108)
  );
  LUT3 #(
    .INIT ( 8'h80 ))
  blk00000462 (
    .I0(sig00000322),
    .I1(sig00000326),
    .I2(sig00000327),
    .O(sig00000410)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000463 (
    .I0(b[25]),
    .I1(a[25]),
    .O(sig000003be)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000464 (
    .I0(b[24]),
    .I1(a[24]),
    .O(sig000003bd)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000465 (
    .I0(b[23]),
    .I1(a[23]),
    .O(sig000003bb)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000466 (
    .I0(b[22]),
    .I1(a[22]),
    .O(sig000003ba)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000467 (
    .I0(b[21]),
    .I1(a[21]),
    .O(sig000003b8)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000468 (
    .I0(b[20]),
    .I1(a[20]),
    .O(sig000003b7)
  );
  LUT2 #(
    .INIT ( 4'h8 ))
  blk00000469 (
    .I0(sig00000143),
    .I1(sig00000157),
    .O(sig00000151)
  );
  LUT2 #(
    .INIT ( 4'h8 ))
  blk0000046a (
    .I0(sig00000145),
    .I1(sig00000159),
    .O(sig00000150)
  );
  LUT2 #(
    .INIT ( 4'h8 ))
  blk0000046b (
    .I0(sig00000141),
    .I1(sig00000155),
    .O(sig0000014f)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk0000046c (
    .I0(b[19]),
    .I1(a[19]),
    .O(sig000003b5)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk0000046d (
    .I0(b[18]),
    .I1(a[18]),
    .O(sig000003b4)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk0000046e (
    .I0(b[17]),
    .I1(a[17]),
    .O(sig000003b2)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk0000046f (
    .I0(b[16]),
    .I1(a[16]),
    .O(sig000003b1)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000470 (
    .I0(sig000002e1),
    .I1(sig000002df),
    .O(sig00000267)
  );
  LUT3 #(
    .INIT ( 8'h32 ))
  blk00000471 (
    .I0(sig00000315),
    .I1(sig00000316),
    .I2(sig00000355),
    .O(sig00000594)
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  blk00000472 (
    .I0(sig0000045f),
    .I1(sig000004ad),
    .I2(sig000004ac),
    .O(sig0000056a)
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  blk00000473 (
    .I0(sig000002e1),
    .I1(sig000002e9),
    .I2(sig000002d7),
    .O(sig00000409)
  );
  LUT4 #(
    .INIT ( 16'h6696 ))
  blk00000474 (
    .I0(sig00000183),
    .I1(sig000001fe),
    .I2(sig000001b1),
    .I3(sig0000020d),
    .O(sig0000022f)
  );
  LUT4 #(
    .INIT ( 16'h6696 ))
  blk00000475 (
    .I0(sig00000199),
    .I1(sig0000025a),
    .I2(sig000000c9),
    .I3(sig00000261),
    .O(sig00000224)
  );
  LUT4 #(
    .INIT ( 16'h151F ))
  blk00000476 (
    .I0(sig0000024b),
    .I1(sig00000033),
    .I2(sig00000088),
    .I3(sig00000087),
    .O(sig00000160)
  );
  LUT4 #(
    .INIT ( 16'h151F ))
  blk00000477 (
    .I0(sig00000247),
    .I1(sig00000034),
    .I2(sig00000088),
    .I3(sig00000087),
    .O(sig0000015f)
  );
  LUT4 #(
    .INIT ( 16'h151F ))
  blk00000478 (
    .I0(sig00000088),
    .I1(sig00000087),
    .I2(sig00000243),
    .I3(sig00000035),
    .O(sig0000015e)
  );
  LUT4 #(
    .INIT ( 16'h151F ))
  blk00000479 (
    .I0(sig00000088),
    .I1(sig00000087),
    .I2(sig00000255),
    .I3(sig00000036),
    .O(sig0000015d)
  );
  LUT4 #(
    .INIT ( 16'h151F ))
  blk0000047a (
    .I0(sig00000088),
    .I1(sig00000087),
    .I2(sig0000024d),
    .I3(sig00000037),
    .O(sig0000015c)
  );
  LUT4 #(
    .INIT ( 16'h9009 ))
  blk0000047b (
    .I0(sig00000334),
    .I1(sig0000045e),
    .I2(sig00000335),
    .I3(sig0000045d),
    .O(sig0000040c)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk0000047c (
    .I0(sig000002e1),
    .I1(sig000002de),
    .O(sig00000266)
  );
  LUT3 #(
    .INIT ( 8'h32 ))
  blk0000047d (
    .I0(sig00000315),
    .I1(sig00000316),
    .I2(sig00000354),
    .O(sig00000593)
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  blk0000047e (
    .I0(sig00000560),
    .I1(sig00000557),
    .I2(sig00000556),
    .O(sig00000575)
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  blk0000047f (
    .I0(sig0000045f),
    .I1(sig000004ae),
    .I2(sig000004ad),
    .O(sig00000569)
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  blk00000480 (
    .I0(sig000002e1),
    .I1(sig000002e8),
    .I2(sig000002d6),
    .O(sig00000408)
  );
  LUT4 #(
    .INIT ( 16'h6696 ))
  blk00000481 (
    .I0(sig00000182),
    .I1(sig000001fe),
    .I2(sig000001b0),
    .I3(sig0000020d),
    .O(sig0000022e)
  );
  LUT4 #(
    .INIT ( 16'h6696 ))
  blk00000482 (
    .I0(sig000001a1),
    .I1(sig0000025a),
    .I2(sig000000c8),
    .I3(sig00000261),
    .O(sig00000223)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000483 (
    .I0(sig000002e1),
    .I1(sig000002dd),
    .O(sig00000265)
  );
  LUT3 #(
    .INIT ( 8'h32 ))
  blk00000484 (
    .I0(sig00000315),
    .I1(sig00000316),
    .I2(sig00000353),
    .O(sig00000592)
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  blk00000485 (
    .I0(sig00000560),
    .I1(sig00000556),
    .I2(sig00000555),
    .O(sig0000057e)
  );
  LUT3 #(
    .INIT ( 8'hAC ))
  blk00000486 (
    .I0(sig000004ae),
    .I1(sig000004af),
    .I2(sig0000045f),
    .O(sig00000573)
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  blk00000487 (
    .I0(sig000002e1),
    .I1(sig000002e7),
    .I2(sig000002d5),
    .O(sig00000407)
  );
  LUT4 #(
    .INIT ( 16'h6696 ))
  blk00000488 (
    .I0(sig00000181),
    .I1(sig000001fe),
    .I2(sig000001af),
    .I3(sig0000020d),
    .O(sig0000022d)
  );
  LUT4 #(
    .INIT ( 16'h6696 ))
  blk00000489 (
    .I0(sig000001a0),
    .I1(sig0000025a),
    .I2(sig000000c7),
    .I3(sig00000261),
    .O(sig00000222)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk0000048a (
    .I0(sig000002dc),
    .I1(sig000002e1),
    .O(sig00000264)
  );
  LUT3 #(
    .INIT ( 8'h32 ))
  blk0000048b (
    .I0(sig00000315),
    .I1(sig00000316),
    .I2(sig00000352),
    .O(sig00000591)
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  blk0000048c (
    .I0(sig00000560),
    .I1(sig00000555),
    .I2(sig00000554),
    .O(sig0000057d)
  );
  LUT3 #(
    .INIT ( 8'hAC ))
  blk0000048d (
    .I0(sig000004af),
    .I1(sig000004b0),
    .I2(sig0000045f),
    .O(sig00000572)
  );
  LUT3 #(
    .INIT ( 8'hAC ))
  blk0000048e (
    .I0(sig000002d4),
    .I1(sig000002e6),
    .I2(sig000002e1),
    .O(sig00000406)
  );
  LUT4 #(
    .INIT ( 16'h6696 ))
  blk0000048f (
    .I0(sig0000018b),
    .I1(sig000001fe),
    .I2(sig000001b9),
    .I3(sig0000020d),
    .O(sig00000238)
  );
  LUT4 #(
    .INIT ( 16'h6696 ))
  blk00000490 (
    .I0(sig0000019f),
    .I1(sig0000025a),
    .I2(sig000000de),
    .I3(sig00000261),
    .O(sig00000221)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000491 (
    .I0(sig000002db),
    .I1(sig000002e1),
    .O(sig00000263)
  );
  LUT3 #(
    .INIT ( 8'h32 ))
  blk00000492 (
    .I0(sig00000315),
    .I1(sig00000316),
    .I2(sig00000351),
    .O(sig00000590)
  );
  LUT3 #(
    .INIT ( 8'hAC ))
  blk00000493 (
    .I0(sig0000055f),
    .I1(sig00000554),
    .I2(sig00000560),
    .O(sig0000057c)
  );
  LUT3 #(
    .INIT ( 8'hAC ))
  blk00000494 (
    .I0(sig000004b0),
    .I1(sig000004b1),
    .I2(sig0000045f),
    .O(sig00000571)
  );
  LUT3 #(
    .INIT ( 8'hAC ))
  blk00000495 (
    .I0(sig000002d3),
    .I1(sig000002e5),
    .I2(sig000002e1),
    .O(sig00000405)
  );
  LUT4 #(
    .INIT ( 16'h6696 ))
  blk00000496 (
    .I0(sig0000018a),
    .I1(sig000001fe),
    .I2(sig000001b8),
    .I3(sig0000020d),
    .O(sig00000237)
  );
  LUT4 #(
    .INIT ( 16'h39C6 ))
  blk00000497 (
    .I0(sig000000dd),
    .I1(sig0000019e),
    .I2(sig00000261),
    .I3(sig0000025a),
    .O(sig0000022b)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000498 (
    .I0(sig000002da),
    .I1(sig000002e1),
    .O(sig00000262)
  );
  LUT3 #(
    .INIT ( 8'h32 ))
  blk00000499 (
    .I0(sig00000315),
    .I1(sig00000316),
    .I2(sig00000350),
    .O(sig0000058f)
  );
  LUT3 #(
    .INIT ( 8'hAC ))
  blk0000049a (
    .I0(sig0000055e),
    .I1(sig0000055f),
    .I2(sig00000560),
    .O(sig0000057b)
  );
  LUT3 #(
    .INIT ( 8'hAC ))
  blk0000049b (
    .I0(sig000004b1),
    .I1(sig000004b2),
    .I2(sig0000045f),
    .O(sig00000570)
  );
  LUT3 #(
    .INIT ( 8'hAC ))
  blk0000049c (
    .I0(sig000002d2),
    .I1(sig000002e4),
    .I2(sig000002e1),
    .O(sig00000404)
  );
  LUT4 #(
    .INIT ( 16'h39C6 ))
  blk0000049d (
    .I0(sig000001b7),
    .I1(sig00000189),
    .I2(sig0000020d),
    .I3(sig000001fe),
    .O(sig00000236)
  );
  LUT4 #(
    .INIT ( 16'h39C6 ))
  blk0000049e (
    .I0(sig000000dc),
    .I1(sig0000019d),
    .I2(sig00000261),
    .I3(sig0000025a),
    .O(sig0000022a)
  );
  LUT3 #(
    .INIT ( 8'hAC ))
  blk0000049f (
    .I0(sig0000055d),
    .I1(sig0000055e),
    .I2(sig00000560),
    .O(sig0000057a)
  );
  LUT3 #(
    .INIT ( 8'hAC ))
  blk000004a0 (
    .I0(sig000004b2),
    .I1(sig000004b3),
    .I2(sig0000045f),
    .O(sig0000056f)
  );
  LUT3 #(
    .INIT ( 8'hAC ))
  blk000004a1 (
    .I0(sig000002d1),
    .I1(sig000002e3),
    .I2(sig000002e1),
    .O(sig00000403)
  );
  LUT4 #(
    .INIT ( 16'h39C6 ))
  blk000004a2 (
    .I0(sig000001b6),
    .I1(sig00000188),
    .I2(sig0000020d),
    .I3(sig000001fe),
    .O(sig00000235)
  );
  LUT4 #(
    .INIT ( 16'h39C6 ))
  blk000004a3 (
    .I0(sig000000db),
    .I1(sig0000019c),
    .I2(sig00000261),
    .I3(sig0000025a),
    .O(sig00000229)
  );
  LUT3 #(
    .INIT ( 8'hAC ))
  blk000004a4 (
    .I0(sig0000055c),
    .I1(sig0000055d),
    .I2(sig00000560),
    .O(sig00000579)
  );
  LUT3 #(
    .INIT ( 8'hAC ))
  blk000004a5 (
    .I0(sig000004b3),
    .I1(sig000004b5),
    .I2(sig0000045f),
    .O(sig0000056e)
  );
  LUT3 #(
    .INIT ( 8'h53 ))
  blk000004a6 (
    .I0(sig000002d0),
    .I1(sig000002e2),
    .I2(sig000002e1),
    .O(sig000003e4)
  );
  LUT4 #(
    .INIT ( 16'h39C6 ))
  blk000004a7 (
    .I0(sig000001b5),
    .I1(sig00000187),
    .I2(sig0000020d),
    .I3(sig000001fe),
    .O(sig00000234)
  );
  LUT4 #(
    .INIT ( 16'h39C6 ))
  blk000004a8 (
    .I0(sig000000da),
    .I1(sig0000019b),
    .I2(sig00000261),
    .I3(sig0000025a),
    .O(sig00000228)
  );
  LUT3 #(
    .INIT ( 8'hAC ))
  blk000004a9 (
    .I0(sig0000055b),
    .I1(sig0000055c),
    .I2(sig00000560),
    .O(sig00000578)
  );
  LUT3 #(
    .INIT ( 8'hAC ))
  blk000004aa (
    .I0(sig000004b5),
    .I1(sig000004b6),
    .I2(sig0000045f),
    .O(sig0000056d)
  );
  LUT4 #(
    .INIT ( 16'h39C6 ))
  blk000004ab (
    .I0(sig000001b4),
    .I1(sig00000186),
    .I2(sig0000020d),
    .I3(sig000001fe),
    .O(sig00000233)
  );
  LUT4 #(
    .INIT ( 16'h39C6 ))
  blk000004ac (
    .I0(sig000000d9),
    .I1(sig0000019a),
    .I2(sig00000261),
    .I3(sig0000025a),
    .O(sig00000227)
  );
  LUT4 #(
    .INIT ( 16'h00AC ))
  blk000004ad (
    .I0(sig00000341),
    .I1(sig00000348),
    .I2(sig00000340),
    .I3(sig0000033e),
    .O(sig000003f5)
  );
  LUT3 #(
    .INIT ( 8'hAC ))
  blk000004ae (
    .I0(sig0000055a),
    .I1(sig0000055b),
    .I2(sig00000560),
    .O(sig00000577)
  );
  LUT3 #(
    .INIT ( 8'hAC ))
  blk000004af (
    .I0(sig000004b6),
    .I1(sig000004b7),
    .I2(sig0000045f),
    .O(sig0000056c)
  );
  LUT4 #(
    .INIT ( 16'h39C6 ))
  blk000004b0 (
    .I0(sig000001b3),
    .I1(sig00000185),
    .I2(sig0000020d),
    .I3(sig000001fe),
    .O(sig00000232)
  );
  LUT4 #(
    .INIT ( 16'h39C6 ))
  blk000004b1 (
    .I0(sig000000d8),
    .I1(sig00000198),
    .I2(sig00000261),
    .I3(sig0000025a),
    .O(sig00000226)
  );
  LUT3 #(
    .INIT ( 8'hAC ))
  blk000004b2 (
    .I0(sig00000559),
    .I1(sig0000055a),
    .I2(sig00000560),
    .O(sig00000576)
  );
  LUT3 #(
    .INIT ( 8'hAC ))
  blk000004b3 (
    .I0(sig000004b7),
    .I1(sig000004b8),
    .I2(sig0000045f),
    .O(sig0000056b)
  );
  LUT4 #(
    .INIT ( 16'h39C6 ))
  blk000004b4 (
    .I0(sig000001b2),
    .I1(sig00000184),
    .I2(sig0000020d),
    .I3(sig000001fe),
    .O(sig00000231)
  );
  LUT4 #(
    .INIT ( 16'h39C6 ))
  blk000004b5 (
    .I0(sig000000d1),
    .I1(sig00000197),
    .I2(sig00000261),
    .I3(sig0000025a),
    .O(sig00000225)
  );
  LUT3 #(
    .INIT ( 8'hAC ))
  blk000004b6 (
    .I0(sig00000558),
    .I1(sig00000559),
    .I2(sig00000560),
    .O(sig00000574)
  );
  LUT3 #(
    .INIT ( 8'hD2 ))
  blk000004b7 (
    .I0(sig000000c6),
    .I1(sig00000261),
    .I2(sig0000025a),
    .O(sig00000212)
  );
  LUT4 #(
    .INIT ( 16'h39C6 ))
  blk000004b8 (
    .I0(sig000001ae),
    .I1(sig00000180),
    .I2(sig0000020d),
    .I3(sig000001fe),
    .O(sig00000230)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000004b9 (
    .I0(sig000004ba),
    .I1(sig000004b9),
    .I2(sig0000045f),
    .O(sig00000565)
  );
  LUT3 #(
    .INIT ( 8'hD2 ))
  blk000004ba (
    .I0(sig000000c5),
    .I1(sig00000261),
    .I2(sig0000025a),
    .O(sig00000211)
  );
  LUT4 #(
    .INIT ( 16'h39C6 ))
  blk000004bb (
    .I0(sig000001ad),
    .I1(sig0000017f),
    .I2(sig0000020d),
    .I3(sig000001fe),
    .O(sig0000022c)
  );
  LUT4 #(
    .INIT ( 16'h0222 ))
  blk000004bc (
    .I0(sig00000581),
    .I1(sig000004bb),
    .I2(sig000004ba),
    .I3(sig0000045f),
    .O(sig00000566)
  );
  LUT3 #(
    .INIT ( 8'hAC ))
  blk000004bd (
    .I0(sig000004b8),
    .I1(sig000004b9),
    .I2(sig0000045f),
    .O(sig00000563)
  );
  LUT3 #(
    .INIT ( 8'h32 ))
  blk000004be (
    .I0(sig0000034f),
    .I1(sig00000316),
    .I2(sig00000315),
    .O(sig0000058e)
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  blk000004bf (
    .I0(sig00000148),
    .O(sig000001ef)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk000004c0 (
    .I0(b[30]),
    .I1(a[30]),
    .O(sig000003c6)
  );
  LUT3 #(
    .INIT ( 8'hAC ))
  blk000004c1 (
    .I0(sig000004b8),
    .I1(sig000004b9),
    .I2(sig0000045f),
    .O(sig00000564)
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  blk000004c2 (
    .I0(sig000001fe),
    .O(sig000001f0)
  );
  LUT4 #(
    .INIT ( 16'hFE01 ))
  blk000004c3 (
    .I0(sig00000532),
    .I1(sig00000315),
    .I2(sig00000316),
    .I3(sig0000058e),
    .O(sig0000058d)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk000004c4 (
    .I0(sig00000333),
    .I1(sig0000045f),
    .O(sig00000371)
  );
  LUT4 #(
    .INIT ( 16'hD580 ))
  blk000004c5 (
    .I0(sig000000c3),
    .I1(sig00000140),
    .I2(sig00000154),
    .I3(sig0000013f),
    .O(sig0000014c)
  );
  LUT4 #(
    .INIT ( 16'hD580 ))
  blk000004c6 (
    .I0(sig000000c3),
    .I1(sig00000142),
    .I2(sig00000156),
    .I3(sig0000014f),
    .O(sig0000014b)
  );
  LUT4 #(
    .INIT ( 16'hD580 ))
  blk000004c7 (
    .I0(sig000000c3),
    .I1(sig00000251),
    .I2(sig0000015a),
    .I3(sig00000150),
    .O(sig0000014d)
  );
  LUT4 #(
    .INIT ( 16'hD580 ))
  blk000004c8 (
    .I0(sig000000c3),
    .I1(sig00000144),
    .I2(sig00000158),
    .I3(sig00000151),
    .O(sig0000014e)
  );
  LUT4 #(
    .INIT ( 16'h0800 ))
  blk000004c9 (
    .I0(sig0000040f),
    .I1(sig00000410),
    .I2(sig0000032a),
    .I3(sig00000323),
    .O(sig0000040e)
  );
  LUT4 #(
    .INIT ( 16'hEFFF ))
  blk000004ca (
    .I0(sig0000033a),
    .I1(sig00000339),
    .I2(sig0000040d),
    .I3(sig0000040c),
    .O(sig00000038)
  );
  LUT4 #(
    .INIT ( 16'h0006 ))
  blk000004cb (
    .I0(sig00000333),
    .I1(sig0000045f),
    .I2(sig00000338),
    .I3(sig00000038),
    .O(sig0000040b)
  );
  LUT3 #(
    .INIT ( 8'h10 ))
  blk000004cc (
    .I0(sig00000585),
    .I1(sig0000047b),
    .I2(sig0000041f),
    .O(sig000004ee)
  );
  LUT3 #(
    .INIT ( 8'h10 ))
  blk000004cd (
    .I0(sig00000585),
    .I1(sig0000047b),
    .I2(sig00000420),
    .O(sig000004ed)
  );
  LUT3 #(
    .INIT ( 8'h10 ))
  blk000004ce (
    .I0(sig00000585),
    .I1(sig0000047b),
    .I2(sig0000042b),
    .O(sig000004ec)
  );
  LUT3 #(
    .INIT ( 8'h10 ))
  blk000004cf (
    .I0(sig00000585),
    .I1(sig0000047b),
    .I2(sig00000432),
    .O(sig000004eb)
  );
  LUT3 #(
    .INIT ( 8'h10 ))
  blk000004d0 (
    .I0(sig00000585),
    .I1(sig0000047b),
    .I2(sig00000433),
    .O(sig000004ea)
  );
  LUT3 #(
    .INIT ( 8'h10 ))
  blk000004d1 (
    .I0(sig00000585),
    .I1(sig0000047b),
    .I2(sig00000434),
    .O(sig000004e9)
  );
  LUT3 #(
    .INIT ( 8'h10 ))
  blk000004d2 (
    .I0(sig00000585),
    .I1(sig0000047b),
    .I2(sig00000435),
    .O(sig000004e8)
  );
  LUT3 #(
    .INIT ( 8'h10 ))
  blk000004d3 (
    .I0(sig00000585),
    .I1(sig0000047b),
    .I2(sig00000436),
    .O(sig000004e6)
  );
  LUT3 #(
    .INIT ( 8'h10 ))
  blk000004d4 (
    .I0(sig0000044f),
    .I1(sig0000044e),
    .I2(sig000004a1),
    .O(sig000004d4)
  );
  LUT3 #(
    .INIT ( 8'h10 ))
  blk000004d5 (
    .I0(sig0000044f),
    .I1(sig0000044e),
    .I2(sig000004a0),
    .O(sig000004d3)
  );
  LUT4 #(
    .INIT ( 16'h0E04 ))
  blk000004d6 (
    .I0(sig0000047b),
    .I1(sig00000425),
    .I2(sig00000585),
    .I3(sig00000435),
    .O(sig000004df)
  );
  LUT4 #(
    .INIT ( 16'h0E04 ))
  blk000004d7 (
    .I0(sig0000047b),
    .I1(sig00000426),
    .I2(sig00000585),
    .I3(sig00000436),
    .O(sig000004de)
  );
  LUT4 #(
    .INIT ( 16'h0E04 ))
  blk000004d8 (
    .I0(sig0000047b),
    .I1(sig00000437),
    .I2(sig00000585),
    .I3(sig0000041f),
    .O(sig000004e5)
  );
  LUT4 #(
    .INIT ( 16'h0E04 ))
  blk000004d9 (
    .I0(sig0000047b),
    .I1(sig00000438),
    .I2(sig00000585),
    .I3(sig00000420),
    .O(sig000004e4)
  );
  LUT4 #(
    .INIT ( 16'h0E04 ))
  blk000004da (
    .I0(sig0000047b),
    .I1(sig00000421),
    .I2(sig00000585),
    .I3(sig0000042b),
    .O(sig000004e3)
  );
  LUT4 #(
    .INIT ( 16'h0E04 ))
  blk000004db (
    .I0(sig0000047b),
    .I1(sig00000422),
    .I2(sig00000585),
    .I3(sig00000432),
    .O(sig000004e2)
  );
  LUT4 #(
    .INIT ( 16'h0E04 ))
  blk000004dc (
    .I0(sig0000047b),
    .I1(sig00000423),
    .I2(sig00000585),
    .I3(sig00000433),
    .O(sig000004e1)
  );
  LUT4 #(
    .INIT ( 16'h0E04 ))
  blk000004dd (
    .I0(sig0000047b),
    .I1(sig00000424),
    .I2(sig00000585),
    .I3(sig00000434),
    .O(sig000004e0)
  );
  LUT4 #(
    .INIT ( 16'h0E04 ))
  blk000004de (
    .I0(sig0000044e),
    .I1(sig0000049f),
    .I2(sig0000044f),
    .I3(sig000004a1),
    .O(sig000004d2)
  );
  LUT4 #(
    .INIT ( 16'h0E04 ))
  blk000004df (
    .I0(sig0000044e),
    .I1(sig0000049e),
    .I2(sig0000044f),
    .I3(sig000004a0),
    .O(sig000004d1)
  );
  LUT2 #(
    .INIT ( 4'h7 ))
  blk000004e0 (
    .I0(sig000003e6),
    .I1(sig000003de),
    .O(sig00000280)
  );
  LUT3 #(
    .INIT ( 8'h1B ))
  blk000004e1 (
    .I0(sig0000047b),
    .I1(sig00000428),
    .I2(sig00000438),
    .O(sig00000039)
  );
  LUT4 #(
    .INIT ( 16'h085D ))
  blk000004e2 (
    .I0(sig00000585),
    .I1(sig00000420),
    .I2(sig00000476),
    .I3(sig00000039),
    .O(sig000004f6)
  );
  LUT4 #(
    .INIT ( 16'h085D ))
  blk000004e3 (
    .I0(sig00000585),
    .I1(sig0000042b),
    .I2(sig00000476),
    .I3(sig0000003a),
    .O(sig000004f5)
  );
  LUT4 #(
    .INIT ( 16'h085D ))
  blk000004e4 (
    .I0(sig00000585),
    .I1(sig0000041f),
    .I2(sig00000476),
    .I3(sig0000003b),
    .O(sig000004dd)
  );
  LUT4 #(
    .INIT ( 16'h085D ))
  blk000004e5 (
    .I0(sig00000585),
    .I1(sig00000432),
    .I2(sig00000476),
    .I3(sig0000003c),
    .O(sig000004f4)
  );
  LUT4 #(
    .INIT ( 16'h085D ))
  blk000004e6 (
    .I0(sig00000585),
    .I1(sig00000433),
    .I2(sig00000476),
    .I3(sig0000003d),
    .O(sig000004f3)
  );
  LUT4 #(
    .INIT ( 16'h085D ))
  blk000004e7 (
    .I0(sig00000585),
    .I1(sig00000434),
    .I2(sig00000476),
    .I3(sig0000003e),
    .O(sig000004f2)
  );
  LUT4 #(
    .INIT ( 16'h085D ))
  blk000004e8 (
    .I0(sig00000585),
    .I1(sig00000435),
    .I2(sig00000476),
    .I3(sig0000003f),
    .O(sig000004f1)
  );
  LUT4 #(
    .INIT ( 16'h085D ))
  blk000004e9 (
    .I0(sig00000585),
    .I1(sig00000436),
    .I2(sig00000476),
    .I3(sig00000040),
    .O(sig000004f0)
  );
  LUT4 #(
    .INIT ( 16'h085D ))
  blk000004ea (
    .I0(sig0000044f),
    .I1(sig000004a1),
    .I2(sig00000450),
    .I3(sig00000041),
    .O(sig000004d0)
  );
  LUT4 #(
    .INIT ( 16'h085D ))
  blk000004eb (
    .I0(sig0000044f),
    .I1(sig000004a0),
    .I2(sig00000450),
    .I3(sig00000042),
    .O(sig000004cf)
  );
  LUT4 #(
    .INIT ( 16'h9009 ))
  blk000004ec (
    .I0(a[28]),
    .I1(b[28]),
    .I2(a[29]),
    .I3(b[29]),
    .O(sig000003c2)
  );
  LUT4 #(
    .INIT ( 16'h9009 ))
  blk000004ed (
    .I0(a[26]),
    .I1(b[26]),
    .I2(a[27]),
    .I3(b[27]),
    .O(sig000003bf)
  );
  LUT4 #(
    .INIT ( 16'h9009 ))
  blk000004ee (
    .I0(a[24]),
    .I1(b[24]),
    .I2(a[25]),
    .I3(b[25]),
    .O(sig000003bc)
  );
  LUT4 #(
    .INIT ( 16'h9009 ))
  blk000004ef (
    .I0(a[22]),
    .I1(b[22]),
    .I2(a[23]),
    .I3(b[23]),
    .O(sig000003b9)
  );
  LUT4 #(
    .INIT ( 16'h9009 ))
  blk000004f0 (
    .I0(a[20]),
    .I1(b[20]),
    .I2(a[21]),
    .I3(b[21]),
    .O(sig000003b6)
  );
  LUT4 #(
    .INIT ( 16'h9009 ))
  blk000004f1 (
    .I0(a[18]),
    .I1(b[18]),
    .I2(a[19]),
    .I3(b[19]),
    .O(sig000003b3)
  );
  LUT4 #(
    .INIT ( 16'h9009 ))
  blk000004f2 (
    .I0(a[16]),
    .I1(b[16]),
    .I2(a[17]),
    .I3(b[17]),
    .O(sig000003b0)
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  blk000004f3 (
    .I0(sig000002d9),
    .O(sig0000023a)
  );
  INV   blk000004f4 (
    .I(sig000001ba),
    .O(sig00000485)
  );
  INV   blk000004f5 (
    .I(sig0000045f),
    .O(sig00000582)
  );
  INV   blk000004f6 (
    .I(sig00000338),
    .O(sig00000376)
  );
  INV   blk000004f7 (
    .I(sig00000339),
    .O(sig00000377)
  );
  INV   blk000004f8 (
    .I(sig0000033a),
    .O(sig00000378)
  );
  MUXF5   blk000004f9 (
    .I0(sig00000043),
    .I1(sig00000044),
    .S(sig00000585),
    .O(sig000004ef)
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  blk000004fa (
    .I0(sig0000047b),
    .I1(sig00000430),
    .I2(sig00000427),
    .O(sig00000043)
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  blk000004fb (
    .I0(sig00000476),
    .I1(sig00000437),
    .I2(sig0000041f),
    .O(sig00000044)
  );
  MUXF5   blk000004fc (
    .I0(sig00000045),
    .I1(sig00000046),
    .S(sig00000585),
    .O(sig000004e7)
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  blk000004fd (
    .I0(sig0000047b),
    .I1(sig00000431),
    .I2(sig00000428),
    .O(sig00000045)
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  blk000004fe (
    .I0(sig00000476),
    .I1(sig00000438),
    .I2(sig00000420),
    .O(sig00000046)
  );
  LUT4 #(
    .INIT ( 16'hFF32 ))
  blk000004ff (
    .I0(sig0000033e),
    .I1(sig00000342),
    .I2(sig000003f5),
    .I3(sig0000033f),
    .O(sig000003f6)
  );
  LUT3 #(
    .INIT ( 8'h10 ))
  blk00000500 (
    .I0(sig0000033f),
    .I1(sig00000342),
    .I2(sig000003f5),
    .O(sig000003f7)
  );
  MUXF5   blk00000501 (
    .I0(sig000003f7),
    .I1(sig000003f6),
    .S(sig00000343),
    .O(sig000003f4)
  );
  LUT4_L #(
    .INIT ( 16'h8880 ))
  blk00000502 (
    .I0(sig0000008b),
    .I1(sig0000008a),
    .I2(sig00000089),
    .I3(sig00000088),
    .LO(sig0000002e)
  );
  LUT3_D #(
    .INIT ( 8'h5D ))
  blk00000503 (
    .I0(sig000003d7),
    .I1(sig000003d8),
    .I2(sig000003a7),
    .LO(sig00000047),
    .O(sig000005a1)
  );
  LUT3_D #(
    .INIT ( 8'hFE ))
  blk00000504 (
    .I0(sig00000386),
    .I1(sig0000037c),
    .I2(sig000002eb),
    .LO(sig00000048),
    .O(sig00000358)
  );
  LUT3_L #(
    .INIT ( 8'h2E ))
  blk00000505 (
    .I0(sig00000340),
    .I1(sig0000033e),
    .I2(sig00000344),
    .LO(sig00000070)
  );
  LUT3_L #(
    .INIT ( 8'h1B ))
  blk00000506 (
    .I0(sig000000e1),
    .I1(sig000000b9),
    .I2(sig000000ba),
    .LO(sig00000050)
  );
  LUT3_L #(
    .INIT ( 8'h1B ))
  blk00000507 (
    .I0(sig000000c3),
    .I1(sig00000097),
    .I2(sig0000009c),
    .LO(sig00000065)
  );
  LUT3_L #(
    .INIT ( 8'h1B ))
  blk00000508 (
    .I0(sig000000c3),
    .I1(sig00000096),
    .I2(sig0000009a),
    .LO(sig0000006d)
  );
  LUT3_L #(
    .INIT ( 8'h1B ))
  blk00000509 (
    .I0(sig000000c3),
    .I1(sig00000095),
    .I2(sig00000099),
    .LO(sig0000006e)
  );
  LUT3_L #(
    .INIT ( 8'h1B ))
  blk0000050a (
    .I0(sig000000c3),
    .I1(sig00000098),
    .I2(sig0000009d),
    .LO(sig0000006f)
  );
  LUT3_D #(
    .INIT ( 8'hAC ))
  blk0000050b (
    .I0(sig0000049b),
    .I1(sig00000496),
    .I2(sig0000044f),
    .LO(sig00000049),
    .O(sig00000071)
  );
  LUT3_D #(
    .INIT ( 8'hAC ))
  blk0000050c (
    .I0(sig00000499),
    .I1(sig00000495),
    .I2(sig0000044f),
    .LO(sig0000004a),
    .O(sig00000073)
  );
  LUT3_D #(
    .INIT ( 8'hCA ))
  blk0000050d (
    .I0(sig00000497),
    .I1(sig0000049c),
    .I2(sig0000044f),
    .LO(sig0000004b),
    .O(sig00000074)
  );
  LUT3_D #(
    .INIT ( 8'hAC ))
  blk0000050e (
    .I0(sig00000498),
    .I1(sig00000494),
    .I2(sig0000044f),
    .LO(sig0000004c),
    .O(sig00000075)
  );
  LUT3_D #(
    .INIT ( 8'hAC ))
  blk0000050f (
    .I0(sig00000497),
    .I1(sig00000493),
    .I2(sig0000044f),
    .LO(sig0000004d),
    .O(sig00000076)
  );
  LUT3_D #(
    .INIT ( 8'hAC ))
  blk00000510 (
    .I0(sig00000496),
    .I1(sig00000492),
    .I2(sig0000044f),
    .LO(sig0000004e),
    .O(sig00000077)
  );
  LUT3_D #(
    .INIT ( 8'hAC ))
  blk00000511 (
    .I0(sig00000495),
    .I1(sig00000491),
    .I2(sig0000044f),
    .LO(sig0000004f),
    .O(sig00000078)
  );
  LUT3_D #(
    .INIT ( 8'hAC ))
  blk00000512 (
    .I0(sig00000493),
    .I1(sig000004a8),
    .I2(sig0000044f),
    .LO(sig00000051),
    .O(sig00000079)
  );
  LUT3_D #(
    .INIT ( 8'hAC ))
  blk00000513 (
    .I0(sig00000492),
    .I1(sig000004a7),
    .I2(sig0000044f),
    .LO(sig00000052),
    .O(sig0000007a)
  );
  LUT3_D #(
    .INIT ( 8'hAC ))
  blk00000514 (
    .I0(sig00000494),
    .I1(sig00000490),
    .I2(sig0000044f),
    .LO(sig00000053),
    .O(sig0000007b)
  );
  LUT3_D #(
    .INIT ( 8'hAC ))
  blk00000515 (
    .I0(sig00000491),
    .I1(sig000004a6),
    .I2(sig0000044f),
    .LO(sig00000054),
    .O(sig0000007c)
  );
  LUT3_D #(
    .INIT ( 8'hAC ))
  blk00000516 (
    .I0(sig00000490),
    .I1(sig000004a5),
    .I2(sig0000044f),
    .LO(sig00000055),
    .O(sig0000007d)
  );
  LUT3_D #(
    .INIT ( 8'hAC ))
  blk00000517 (
    .I0(sig000004a8),
    .I1(sig000004a4),
    .I2(sig0000044f),
    .LO(sig00000056),
    .O(sig0000007e)
  );
  LUT3_L #(
    .INIT ( 8'hCA ))
  blk00000518 (
    .I0(sig0000049a),
    .I1(sig000004a5),
    .I2(sig0000044f),
    .LO(sig00000081)
  );
  LUT3_D #(
    .INIT ( 8'hCA ))
  blk00000519 (
    .I0(sig0000049b),
    .I1(sig0000049f),
    .I2(sig0000044f),
    .LO(sig00000057),
    .O(sig00000082)
  );
  LUT3_L #(
    .INIT ( 8'hCA ))
  blk0000051a (
    .I0(sig0000049d),
    .I1(sig000004a1),
    .I2(sig0000044f),
    .LO(sig00000083)
  );
  LUT3_D #(
    .INIT ( 8'hCA ))
  blk0000051b (
    .I0(sig00000499),
    .I1(sig0000049e),
    .I2(sig0000044f),
    .LO(sig00000058),
    .O(sig00000085)
  );
  LUT3_L #(
    .INIT ( 8'hCA ))
  blk0000051c (
    .I0(sig0000049c),
    .I1(sig000004a0),
    .I2(sig0000044f),
    .LO(sig00000086)
  );
  LUT3_D #(
    .INIT ( 8'hAC ))
  blk0000051d (
    .I0(sig000000ab),
    .I1(sig000000c2),
    .I2(sig000000e1),
    .LO(sig00000059),
    .O(sig00000003)
  );
  LUT3_D #(
    .INIT ( 8'hAC ))
  blk0000051e (
    .I0(sig000000ad),
    .I1(sig000000ac),
    .I2(sig000000e1),
    .LO(sig0000005a),
    .O(sig00000004)
  );
  LUT3_D #(
    .INIT ( 8'hAC ))
  blk0000051f (
    .I0(sig000000c2),
    .I1(sig000000c1),
    .I2(sig000000e1),
    .LO(sig0000005b),
    .O(sig00000005)
  );
  LUT3_D #(
    .INIT ( 8'hAC ))
  blk00000520 (
    .I0(sig000000ac),
    .I1(sig000000ab),
    .I2(sig000000e1),
    .LO(sig0000005c),
    .O(sig00000006)
  );
  LUT3_L #(
    .INIT ( 8'hCA ))
  blk00000521 (
    .I0(sig000000a9),
    .I1(sig000000aa),
    .I2(sig000000e1),
    .LO(sig00000007)
  );
  LUT3_D #(
    .INIT ( 8'hAC ))
  blk00000522 (
    .I0(sig000000bc),
    .I1(sig000000b5),
    .I2(sig000000e1),
    .LO(sig0000005d),
    .O(sig00000008)
  );
  LUT3_D #(
    .INIT ( 8'hAC ))
  blk00000523 (
    .I0(sig000000c1),
    .I1(sig000000c0),
    .I2(sig000000e1),
    .LO(sig0000005e),
    .O(sig00000009)
  );
  LUT3_D #(
    .INIT ( 8'hAC ))
  blk00000524 (
    .I0(sig000000c0),
    .I1(sig000000bf),
    .I2(sig000000e1),
    .LO(sig0000005f),
    .O(sig0000000a)
  );
  LUT3_D #(
    .INIT ( 8'hAC ))
  blk00000525 (
    .I0(sig000000bf),
    .I1(sig000000be),
    .I2(sig000000e1),
    .LO(sig00000060),
    .O(sig0000000b)
  );
  LUT3_D #(
    .INIT ( 8'hAC ))
  blk00000526 (
    .I0(sig000000be),
    .I1(sig000000bd),
    .I2(sig000000e1),
    .LO(sig00000061),
    .O(sig0000000c)
  );
  LUT3_D #(
    .INIT ( 8'hAC ))
  blk00000527 (
    .I0(sig000000bd),
    .I1(sig000000bc),
    .I2(sig000000e1),
    .LO(sig00000062),
    .O(sig0000000d)
  );
  LUT3_L #(
    .INIT ( 8'hE4 ))
  blk00000528 (
    .I0(sig000000e1),
    .I1(sig000000ba),
    .I2(sig000000bb),
    .LO(sig0000000f)
  );
  LUT3_L #(
    .INIT ( 8'hE4 ))
  blk00000529 (
    .I0(sig000000e1),
    .I1(sig000000b9),
    .I2(sig000000ba),
    .LO(sig00000011)
  );
  LUT3_D #(
    .INIT ( 8'hAC ))
  blk0000052a (
    .I0(sig000000b7),
    .I1(sig000000b6),
    .I2(sig000000e1),
    .LO(sig00000063),
    .O(sig00000012)
  );
  LUT3_D #(
    .INIT ( 8'hAC ))
  blk0000052b (
    .I0(sig000000b6),
    .I1(sig000000b4),
    .I2(sig000000e1),
    .LO(sig00000064),
    .O(sig00000013)
  );
  LUT3_D #(
    .INIT ( 8'hAC ))
  blk0000052c (
    .I0(sig000000b4),
    .I1(sig000000b3),
    .I2(sig000000e1),
    .LO(sig00000066),
    .O(sig00000014)
  );
  LUT3_D #(
    .INIT ( 8'hAC ))
  blk0000052d (
    .I0(sig000000b3),
    .I1(sig000000b2),
    .I2(sig000000e1),
    .LO(sig00000067),
    .O(sig00000015)
  );
  LUT3_D #(
    .INIT ( 8'hAC ))
  blk0000052e (
    .I0(sig000000b2),
    .I1(sig000000b1),
    .I2(sig000000e1),
    .LO(sig00000068),
    .O(sig00000016)
  );
  LUT3_D #(
    .INIT ( 8'hAC ))
  blk0000052f (
    .I0(sig000000b1),
    .I1(sig000000b0),
    .I2(sig000000e1),
    .LO(sig00000069),
    .O(sig00000017)
  );
  LUT3_D #(
    .INIT ( 8'hAC ))
  blk00000530 (
    .I0(sig000000b0),
    .I1(sig000000af),
    .I2(sig000000e1),
    .LO(sig0000006a),
    .O(sig00000018)
  );
  LUT3_D #(
    .INIT ( 8'hAC ))
  blk00000531 (
    .I0(sig000000af),
    .I1(sig000000ae),
    .I2(sig000000e1),
    .LO(sig0000006b),
    .O(sig00000019)
  );
  LUT3_D #(
    .INIT ( 8'hAC ))
  blk00000532 (
    .I0(sig000000ae),
    .I1(sig000000ad),
    .I2(sig000000e1),
    .LO(sig0000006c),
    .O(sig0000001a)
  );
  LUT3_L #(
    .INIT ( 8'hAC ))
  blk00000533 (
    .I0(sig000000b5),
    .I1(sig000000aa),
    .I2(sig000000e1),
    .LO(sig0000001b)
  );
  LUT3_L #(
    .INIT ( 8'hAC ))
  blk00000534 (
    .I0(sig000000a1),
    .I1(sig0000009d),
    .I2(sig000000c3),
    .LO(sig0000001d)
  );
  LUT3_L #(
    .INIT ( 8'hAC ))
  blk00000535 (
    .I0(sig000000a0),
    .I1(sig0000009c),
    .I2(sig000000c3),
    .LO(sig0000001f)
  );
  LUT3_L #(
    .INIT ( 8'hAC ))
  blk00000536 (
    .I0(sig0000009f),
    .I1(sig0000009a),
    .I2(sig000000c3),
    .LO(sig00000021)
  );
  LUT3_L #(
    .INIT ( 8'hCA ))
  blk00000537 (
    .I0(sig00000098),
    .I1(sig0000009d),
    .I2(sig000000c3),
    .LO(sig00000023)
  );
  LUT3_L #(
    .INIT ( 8'hCA ))
  blk00000538 (
    .I0(sig00000097),
    .I1(sig0000009c),
    .I2(sig000000c3),
    .LO(sig00000025)
  );
  LUT3_L #(
    .INIT ( 8'hAC ))
  blk00000539 (
    .I0(sig00000092),
    .I1(sig000000a6),
    .I2(sig000000c3),
    .LO(sig00000026)
  );
  LUT3_L #(
    .INIT ( 8'hAC ))
  blk0000053a (
    .I0(sig00000091),
    .I1(sig000000a5),
    .I2(sig000000c3),
    .LO(sig00000028)
  );
  LUT3_L #(
    .INIT ( 8'hAC ))
  blk0000053b (
    .I0(sig0000009e),
    .I1(sig00000099),
    .I2(sig000000c3),
    .LO(sig0000002b)
  );
  LUT3_L #(
    .INIT ( 8'hAC ))
  blk0000053c (
    .I0(sig000000a8),
    .I1(sig000000a4),
    .I2(sig000000c3),
    .LO(sig0000002c)
  );
  LUT3_L #(
    .INIT ( 8'hAC ))
  blk0000053d (
    .I0(sig000000a7),
    .I1(sig000000a3),
    .I2(sig000000c3),
    .LO(sig0000002d)
  );
  LUT3_L #(
    .INIT ( 8'hCA ))
  blk0000053e (
    .I0(sig000000a2),
    .I1(sig000000a6),
    .I2(sig000000c3),
    .LO(sig0000002f)
  );
  LUT3_L #(
    .INIT ( 8'hCA ))
  blk0000053f (
    .I0(sig0000009b),
    .I1(sig000000a5),
    .I2(sig000000c3),
    .LO(sig00000030)
  );
  LUT3_L #(
    .INIT ( 8'hCA ))
  blk00000540 (
    .I0(sig00000090),
    .I1(sig000000a4),
    .I2(sig000000c3),
    .LO(sig00000032)
  );
  LUT4_L #(
    .INIT ( 16'h8000 ))
  blk00000541 (
    .I0(sig00000328),
    .I1(sig00000329),
    .I2(sig00000324),
    .I3(sig00000325),
    .LO(sig0000040f)
  );
  LUT3_L #(
    .INIT ( 8'hEA ))
  blk00000542 (
    .I0(sig0000024c),
    .I1(sig0000024e),
    .I2(sig00000087),
    .LO(sig00000033)
  );
  LUT3_L #(
    .INIT ( 8'hEA ))
  blk00000543 (
    .I0(sig00000248),
    .I1(sig00000249),
    .I2(sig00000087),
    .LO(sig00000034)
  );
  LUT3_L #(
    .INIT ( 8'hEA ))
  blk00000544 (
    .I0(sig00000244),
    .I1(sig00000245),
    .I2(sig00000087),
    .LO(sig00000035)
  );
  LUT3_L #(
    .INIT ( 8'hEA ))
  blk00000545 (
    .I0(sig00000256),
    .I1(sig00000257),
    .I2(sig00000087),
    .LO(sig00000036)
  );
  LUT3_L #(
    .INIT ( 8'hEA ))
  blk00000546 (
    .I0(sig00000252),
    .I1(sig00000253),
    .I2(sig00000087),
    .LO(sig00000037)
  );
  LUT4_L #(
    .INIT ( 16'h9009 ))
  blk00000547 (
    .I0(sig00000336),
    .I1(sig0000043d),
    .I2(sig00000337),
    .I3(sig0000043c),
    .LO(sig0000040d)
  );
  LUT3_L #(
    .INIT ( 8'h1B ))
  blk00000548 (
    .I0(sig0000047b),
    .I1(sig00000429),
    .I2(sig00000421),
    .LO(sig0000003a)
  );
  LUT3_L #(
    .INIT ( 8'h1B ))
  blk00000549 (
    .I0(sig0000047b),
    .I1(sig00000427),
    .I2(sig00000437),
    .LO(sig0000003b)
  );
  LUT3_L #(
    .INIT ( 8'h1B ))
  blk0000054a (
    .I0(sig0000047b),
    .I1(sig0000042a),
    .I2(sig00000422),
    .LO(sig0000003c)
  );
  LUT3_L #(
    .INIT ( 8'h1B ))
  blk0000054b (
    .I0(sig0000047b),
    .I1(sig0000042c),
    .I2(sig00000423),
    .LO(sig0000003d)
  );
  LUT3_L #(
    .INIT ( 8'h1B ))
  blk0000054c (
    .I0(sig0000047b),
    .I1(sig0000042d),
    .I2(sig00000424),
    .LO(sig0000003e)
  );
  LUT3_L #(
    .INIT ( 8'h1B ))
  blk0000054d (
    .I0(sig0000047b),
    .I1(sig0000042e),
    .I2(sig00000425),
    .LO(sig0000003f)
  );
  LUT3_L #(
    .INIT ( 8'h1B ))
  blk0000054e (
    .I0(sig0000047b),
    .I1(sig0000042f),
    .I2(sig00000426),
    .LO(sig00000040)
  );
  LUT3_L #(
    .INIT ( 8'h1B ))
  blk0000054f (
    .I0(sig0000044e),
    .I1(sig0000049d),
    .I2(sig0000049f),
    .LO(sig00000041)
  );
  LUT3_L #(
    .INIT ( 8'h1B ))
  blk00000550 (
    .I0(sig0000044e),
    .I1(sig0000049c),
    .I2(sig0000049e),
    .LO(sig00000042)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000551 (
    .A0(sig00000001),
    .A1(sig00000001),
    .A2(sig00000001),
    .A3(sig00000001),
    .CE(ce),
    .CLK(clk),
    .D(sig00000087),
    .Q(sig000000df)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000552 (
    .C(clk),
    .CE(ce),
    .D(sig000000df),
    .Q(sig000000e1)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000553 (
    .A0(sig00000001),
    .A1(sig00000002),
    .A2(sig00000001),
    .A3(sig00000001),
    .CE(ce),
    .CLK(clk),
    .D(sig000003da),
    .Q(sig00000259)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000554 (
    .C(clk),
    .CE(ce),
    .D(sig00000259),
    .Q(sig0000025a)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000555 (
    .A0(sig00000001),
    .A1(sig00000001),
    .A2(sig00000001),
    .A3(sig00000001),
    .CE(ce),
    .CLK(clk),
    .D(sig0000025f),
    .Q(sig0000025e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000556 (
    .C(clk),
    .CE(ce),
    .D(sig0000025e),
    .Q(sig00000260)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000557 (
    .A0(sig00000001),
    .A1(sig00000002),
    .A2(sig00000001),
    .A3(sig00000001),
    .CE(ce),
    .CLK(clk),
    .D(sig00000172),
    .Q(sig00000165)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000558 (
    .C(clk),
    .CE(ce),
    .D(sig00000165),
    .Q(sig0000017f)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000559 (
    .A0(sig00000001),
    .A1(sig00000001),
    .A2(sig00000001),
    .A3(sig00000001),
    .CE(ce),
    .CLK(clk),
    .D(sig00000088),
    .Q(sig000000e0)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000055a (
    .C(clk),
    .CE(ce),
    .D(sig000000e0),
    .Q(sig000000e2)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000055b (
    .A0(sig00000001),
    .A1(sig00000001),
    .A2(sig00000001),
    .A3(sig00000001),
    .CE(ce),
    .CLK(clk),
    .D(sig0000008b),
    .Q(sig00000149)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000055c (
    .C(clk),
    .CE(ce),
    .D(sig00000149),
    .Q(sig0000014a)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000055d (
    .A0(sig00000001),
    .A1(sig00000002),
    .A2(sig00000001),
    .A3(sig00000001),
    .CE(ce),
    .CLK(clk),
    .D(sig00000178),
    .Q(sig0000016b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000055e (
    .C(clk),
    .CE(ce),
    .D(sig0000016b),
    .Q(sig00000185)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000055f (
    .A0(sig00000001),
    .A1(sig00000002),
    .A2(sig00000001),
    .A3(sig00000001),
    .CE(ce),
    .CLK(clk),
    .D(sig00000173),
    .Q(sig00000166)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000560 (
    .C(clk),
    .CE(ce),
    .D(sig00000166),
    .Q(sig00000180)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000561 (
    .A0(sig00000001),
    .A1(sig00000002),
    .A2(sig00000001),
    .A3(sig00000001),
    .CE(ce),
    .CLK(clk),
    .D(sig00000177),
    .Q(sig0000016a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000562 (
    .C(clk),
    .CE(ce),
    .D(sig0000016a),
    .Q(sig00000184)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000563 (
    .A0(sig00000001),
    .A1(sig00000002),
    .A2(sig00000001),
    .A3(sig00000001),
    .CE(ce),
    .CLK(clk),
    .D(sig00000179),
    .Q(sig0000016c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000564 (
    .C(clk),
    .CE(ce),
    .D(sig0000016c),
    .Q(sig00000186)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000565 (
    .A0(sig00000001),
    .A1(sig00000002),
    .A2(sig00000001),
    .A3(sig00000001),
    .CE(ce),
    .CLK(clk),
    .D(sig0000017a),
    .Q(sig0000016d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000566 (
    .C(clk),
    .CE(ce),
    .D(sig0000016d),
    .Q(sig00000187)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000567 (
    .A0(sig00000001),
    .A1(sig00000002),
    .A2(sig00000001),
    .A3(sig00000001),
    .CE(ce),
    .CLK(clk),
    .D(sig0000017d),
    .Q(sig00000170)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000568 (
    .C(clk),
    .CE(ce),
    .D(sig00000170),
    .Q(sig0000018a)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000569 (
    .A0(sig00000001),
    .A1(sig00000002),
    .A2(sig00000001),
    .A3(sig00000001),
    .CE(ce),
    .CLK(clk),
    .D(sig0000017b),
    .Q(sig0000016e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000056a (
    .C(clk),
    .CE(ce),
    .D(sig0000016e),
    .Q(sig00000188)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000056b (
    .A0(sig00000001),
    .A1(sig00000002),
    .A2(sig00000001),
    .A3(sig00000001),
    .CE(ce),
    .CLK(clk),
    .D(sig0000017c),
    .Q(sig0000016f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000056c (
    .C(clk),
    .CE(ce),
    .D(sig0000016f),
    .Q(sig00000189)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000056d (
    .A0(sig00000001),
    .A1(sig00000002),
    .A2(sig00000001),
    .A3(sig00000001),
    .CE(ce),
    .CLK(clk),
    .D(sig00000175),
    .Q(sig00000168)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000056e (
    .C(clk),
    .CE(ce),
    .D(sig00000168),
    .Q(sig00000182)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000056f (
    .A0(sig00000001),
    .A1(sig00000002),
    .A2(sig00000001),
    .A3(sig00000001),
    .CE(ce),
    .CLK(clk),
    .D(sig0000017e),
    .Q(sig00000171)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000570 (
    .C(clk),
    .CE(ce),
    .D(sig00000171),
    .Q(sig0000018b)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000571 (
    .A0(sig00000001),
    .A1(sig00000002),
    .A2(sig00000001),
    .A3(sig00000001),
    .CE(ce),
    .CLK(clk),
    .D(sig00000174),
    .Q(sig00000167)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000572 (
    .C(clk),
    .CE(ce),
    .D(sig00000167),
    .Q(sig00000181)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000573 (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000001),
    .A3(sig00000001),
    .CE(ce),
    .CLK(clk),
    .D(sig000001a3),
    .Q(sig0000018d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000574 (
    .C(clk),
    .CE(ce),
    .D(sig0000018d),
    .Q(sig00000198)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000575 (
    .A0(sig00000001),
    .A1(sig00000002),
    .A2(sig00000001),
    .A3(sig00000001),
    .CE(ce),
    .CLK(clk),
    .D(sig00000176),
    .Q(sig00000169)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000576 (
    .C(clk),
    .CE(ce),
    .D(sig00000169),
    .Q(sig00000183)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000577 (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000001),
    .A3(sig00000001),
    .CE(ce),
    .CLK(clk),
    .D(sig000001a2),
    .Q(sig0000018c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000578 (
    .C(clk),
    .CE(ce),
    .D(sig0000018c),
    .Q(sig00000197)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000579 (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000001),
    .A3(sig00000001),
    .CE(ce),
    .CLK(clk),
    .D(sig000001a5),
    .Q(sig0000018f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000057a (
    .C(clk),
    .CE(ce),
    .D(sig0000018f),
    .Q(sig0000019a)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000057b (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000001),
    .A3(sig00000001),
    .CE(ce),
    .CLK(clk),
    .D(sig000001a6),
    .Q(sig00000190)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000057c (
    .C(clk),
    .CE(ce),
    .D(sig00000190),
    .Q(sig0000019b)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000057d (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000001),
    .A3(sig00000001),
    .CE(ce),
    .CLK(clk),
    .D(sig000001a9),
    .Q(sig00000193)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000057e (
    .C(clk),
    .CE(ce),
    .D(sig00000193),
    .Q(sig0000019e)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000057f (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000001),
    .A3(sig00000001),
    .CE(ce),
    .CLK(clk),
    .D(sig000001a7),
    .Q(sig00000191)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000580 (
    .C(clk),
    .CE(ce),
    .D(sig00000191),
    .Q(sig0000019c)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000581 (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000001),
    .A3(sig00000001),
    .CE(ce),
    .CLK(clk),
    .D(sig000001a8),
    .Q(sig00000192)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000582 (
    .C(clk),
    .CE(ce),
    .D(sig00000192),
    .Q(sig0000019d)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000583 (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000001),
    .A3(sig00000001),
    .CE(ce),
    .CLK(clk),
    .D(sig000001ac),
    .Q(sig00000196)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000584 (
    .C(clk),
    .CE(ce),
    .D(sig00000196),
    .Q(sig000001a1)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000585 (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000001),
    .A3(sig00000001),
    .CE(ce),
    .CLK(clk),
    .D(sig000001aa),
    .Q(sig00000194)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000586 (
    .C(clk),
    .CE(ce),
    .D(sig00000194),
    .Q(sig0000019f)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000587 (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000001),
    .A3(sig00000001),
    .CE(ce),
    .CLK(clk),
    .D(sig000001ab),
    .Q(sig00000195)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000588 (
    .C(clk),
    .CE(ce),
    .D(sig00000195),
    .Q(sig000001a0)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000589 (
    .A0(sig00000001),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000001),
    .CE(ce),
    .CLK(clk),
    .D(sig0000034e),
    .Q(sig0000034a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000058a (
    .C(clk),
    .CE(ce),
    .D(sig0000034a),
    .Q(sig0000034c)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000058b (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000001),
    .A3(sig00000001),
    .CE(ce),
    .CLK(clk),
    .D(sig000001a4),
    .Q(sig0000018e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000058c (
    .C(clk),
    .CE(ce),
    .D(sig0000018e),
    .Q(sig00000199)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000058d (
    .A0(sig00000001),
    .A1(sig00000001),
    .A2(sig00000001),
    .A3(sig00000001),
    .CE(ce),
    .CLK(clk),
    .D(sig0000037a),
    .Q(sig00000379)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000058e (
    .C(clk),
    .CE(ce),
    .D(sig00000379),
    .Q(sig0000037b)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000058f (
    .A0(sig00000001),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000001),
    .CE(ce),
    .CLK(clk),
    .D(sig0000034d),
    .Q(sig00000349)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000590 (
    .C(clk),
    .CE(ce),
    .D(sig00000349),
    .Q(sig0000034b)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000591 (
    .A0(sig00000001),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000001),
    .CE(ce),
    .CLK(clk),
    .D(sig00000347),
    .Q(sig00000345)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000592 (
    .C(clk),
    .CE(ce),
    .D(sig00000345),
    .Q(sig00000346)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000593 (
    .A0(sig00000001),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000001),
    .CE(ce),
    .CLK(clk),
    .D(sig00000327),
    .Q(sig00000330)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000594 (
    .C(clk),
    .CE(ce),
    .D(sig00000330),
    .Q(sig00000338)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000595 (
    .A0(sig00000001),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000001),
    .CE(ce),
    .CLK(clk),
    .D(sig00000329),
    .Q(sig00000332)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000596 (
    .C(clk),
    .CE(ce),
    .D(sig00000332),
    .Q(sig0000033a)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000597 (
    .A0(sig00000001),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000001),
    .CE(ce),
    .CLK(clk),
    .D(sig00000328),
    .Q(sig00000331)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000598 (
    .C(clk),
    .CE(ce),
    .D(sig00000331),
    .Q(sig00000339)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000599 (
    .A0(sig00000001),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000001),
    .CE(ce),
    .CLK(clk),
    .D(sig00000324),
    .Q(sig0000032d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000059a (
    .C(clk),
    .CE(ce),
    .D(sig0000032d),
    .Q(sig00000335)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000059b (
    .A0(sig00000001),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000001),
    .CE(ce),
    .CLK(clk),
    .D(sig00000326),
    .Q(sig0000032f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000059c (
    .C(clk),
    .CE(ce),
    .D(sig0000032f),
    .Q(sig00000337)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000059d (
    .A0(sig00000001),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000001),
    .CE(ce),
    .CLK(clk),
    .D(sig00000325),
    .Q(sig0000032e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000059e (
    .C(clk),
    .CE(ce),
    .D(sig0000032e),
    .Q(sig00000336)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000059f (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000001),
    .CE(ce),
    .CLK(clk),
    .D(sig0000033c),
    .Q(sig0000033b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000005a0 (
    .C(clk),
    .CE(ce),
    .D(sig0000033b),
    .Q(sig0000033d)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000005a1 (
    .A0(sig00000001),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000001),
    .CE(ce),
    .CLK(clk),
    .D(sig00000323),
    .Q(sig0000032c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000005a2 (
    .C(clk),
    .CE(ce),
    .D(sig0000032c),
    .Q(sig00000334)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000005a3 (
    .A0(sig00000001),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000001),
    .CE(ce),
    .CLK(clk),
    .D(sig00000322),
    .Q(sig0000032b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000005a4 (
    .C(clk),
    .CE(ce),
    .D(sig0000032b),
    .Q(sig00000333)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000005a5 (
    .A0(sig00000001),
    .A1(sig00000001),
    .A2(sig00000001),
    .A3(sig00000001),
    .CE(ce),
    .CLK(clk),
    .D(sig00000585),
    .Q(sig0000043a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000005a6 (
    .C(clk),
    .CE(ce),
    .D(sig0000043a),
    .Q(sig0000043c)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000005a7 (
    .A0(sig00000001),
    .A1(sig00000002),
    .A2(sig00000001),
    .A3(sig00000001),
    .CE(ce),
    .CLK(clk),
    .D(sig0000025d),
    .Q(sig00000580)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000005a8 (
    .C(clk),
    .CE(ce),
    .D(sig00000580),
    .Q(sig00000581)
  );
// synthesis translate_on
endmodule