module header
    // Internal signals
		// Generated Signal List
		// End of Generated Signal List
    // %COMPILER_OPTS%
	// Generated Signal Assignments
    // Generated Instances
    // wiring ...
	// Generated Instances and Port Mappings
		// Generated Instance Port Map for inst_a
		inst_a_e inst_a(
			.p_mix_sig_in_01_gi(sig_in_01),
			.p_mix_sig_in_03_gi(sig_in_03),
			.p_mix_sig_io_05_gc(sig_io_05),
			.p_mix_sig_io_06_gc(sig_io_06),
			.p_mix_sig_out_02_go(sig_out_02),
			.p_mix_sig_out_04_go(sig_out_04)
		);
		// End of Generated Instance Port Map for inst_a
endmodule