module top(
	output reg serial_tx,
	input serial_rx,
	input cpu_reset,
	(* dont_touch = "true" *)	input clk100,
	output [13:0] ddram_a,
	output [2:0] ddram_ba,
	output ddram_ras_n,
	output ddram_cas_n,
	output ddram_we_n,
	output ddram_cs_n,
	output [1:0] ddram_dm,
	inout [15:0] ddram_dq,
	output [1:0] ddram_dqs_p,
	output [1:0] ddram_dqs_n,
	output ddram_clk_p,
	output ddram_clk_n,
	output ddram_cke,
	output ddram_odt,
	output ddram_reset_n,
	output [3:0] led
);
wire [3:0] led;
assign led[0] = main_locked;
assign led[1] = idelayctl_rdy;
assign led[2] = 0;
assign led[3] = 0;
// Manually inserted OBUFs
wire [13:0] ddram_a_iob;
wire [ 2:0] ddram_ba_iob;
wire        ddram_ras_n_iob;
wire        ddram_cas_n_iob;
wire        ddram_we_n_iob;
wire        ddram_cs_n_iob;
wire [ 1:0] ddram_dm_iob;
wire        ddram_cke_iob;
wire        ddram_odt_iob;
wire        ddram_reset_n_iob;
OBUF #(.IOSTANDARD("SSTL135"), .SLEW("FAST")) obuf_a0  (.I(ddram_a_iob[ 0]), .O(ddram_a[ 0]));
OBUF #(.IOSTANDARD("SSTL135"), .SLEW("FAST")) obuf_a1  (.I(ddram_a_iob[ 1]), .O(ddram_a[ 1]));
OBUF #(.IOSTANDARD("SSTL135"), .SLEW("FAST")) obuf_a2  (.I(ddram_a_iob[ 2]), .O(ddram_a[ 2]));
OBUF #(.IOSTANDARD("SSTL135"), .SLEW("FAST")) obuf_a3  (.I(ddram_a_iob[ 3]), .O(ddram_a[ 3]));
OBUF #(.IOSTANDARD("SSTL135"), .SLEW("FAST")) obuf_a4  (.I(ddram_a_iob[ 4]), .O(ddram_a[ 4]));
OBUF #(.IOSTANDARD("SSTL135"), .SLEW("FAST")) obuf_a5  (.I(ddram_a_iob[ 5]), .O(ddram_a[ 5]));
OBUF #(.IOSTANDARD("SSTL135"), .SLEW("FAST")) obuf_a6  (.I(ddram_a_iob[ 6]), .O(ddram_a[ 6]));
OBUF #(.IOSTANDARD("SSTL135"), .SLEW("FAST")) obuf_a7  (.I(ddram_a_iob[ 7]), .O(ddram_a[ 7]));
OBUF #(.IOSTANDARD("SSTL135"), .SLEW("FAST")) obuf_a8  (.I(ddram_a_iob[ 8]), .O(ddram_a[ 8]));
OBUF #(.IOSTANDARD("SSTL135"), .SLEW("FAST")) obuf_a9  (.I(ddram_a_iob[ 9]), .O(ddram_a[ 9]));
OBUF #(.IOSTANDARD("SSTL135"), .SLEW("FAST")) obuf_a10 (.I(ddram_a_iob[10]), .O(ddram_a[10]));
OBUF #(.IOSTANDARD("SSTL135"), .SLEW("FAST")) obuf_a11 (.I(ddram_a_iob[11]), .O(ddram_a[11]));
OBUF #(.IOSTANDARD("SSTL135"), .SLEW("FAST")) obuf_a12 (.I(ddram_a_iob[12]), .O(ddram_a[12]));
OBUF #(.IOSTANDARD("SSTL135"), .SLEW("FAST")) obuf_a13 (.I(ddram_a_iob[13]), .O(ddram_a[13]));
OBUF #(.IOSTANDARD("SSTL135"), .SLEW("FAST")) obuf_ba0 (.I(ddram_ba_iob[0]), .O(ddram_ba[0]));
OBUF #(.IOSTANDARD("SSTL135"), .SLEW("FAST")) obuf_ba1 (.I(ddram_ba_iob[1]), .O(ddram_ba[1]));
OBUF #(.IOSTANDARD("SSTL135"), .SLEW("FAST")) obuf_ba2 (.I(ddram_ba_iob[2]), .O(ddram_ba[2]));
OBUF #(.IOSTANDARD("SSTL135"), .SLEW("FAST")) obuf_dm0 (.I(ddram_dm_iob[0]), .O(ddram_dm[0]));
OBUF #(.IOSTANDARD("SSTL135"), .SLEW("FAST")) obuf_dm1 (.I(ddram_dm_iob[1]), .O(ddram_dm[1]));
OBUF #(.IOSTANDARD("SSTL135"), .SLEW("FAST")) obuf_ras (.I(ddram_ras_n_iob), .O(ddram_ras_n));
OBUF #(.IOSTANDARD("SSTL135"), .SLEW("FAST")) obuf_cas (.I(ddram_cas_n_iob), .O(ddram_cas_n));
OBUF #(.IOSTANDARD("SSTL135"), .SLEW("FAST")) obuf_we  (.I(ddram_we_n_iob),  .O(ddram_we_n));
OBUF #(.IOSTANDARD("SSTL135"), .SLEW("FAST")) obuf_cs  (.I(ddram_cs_n_iob),  .O(ddram_cs_n));
OBUF #(.IOSTANDARD("SSTL135"), .SLEW("FAST")) obuf_cke (.I(ddram_cke_iob),  .O(ddram_cke));
OBUF #(.IOSTANDARD("SSTL135"), .SLEW("FAST")) obuf_odt (.I(ddram_odt_iob),  .O(ddram_odt));
OBUF #(.IOSTANDARD("SSTL135"), .SLEW("FAST")) obuf_rst (.I(ddram_reset_n_iob),.O(ddram_reset_n));
// End manually inserted OBUFs
wire idelayctl_rdy;
reg main_ctrl_reset_storage = 1'd0;
reg main_ctrl_reset_re = 1'd0;
reg [31:0] main_ctrl_scratch_storage = 32'd305419896;
reg main_ctrl_scratch_re = 1'd0;
wire [31:0] main_ctrl_bus_errors_status;
wire main_ctrl_bus_errors_we;
wire main_ctrl_reset;
wire main_ctrl_bus_error;
reg [31:0] main_ctrl_bus_errors = 32'd0;
wire [29:0] main_sram_bus_adr;
wire [31:0] main_sram_bus_dat_w;
wire [31:0] main_sram_bus_dat_r;
wire [3:0] main_sram_bus_sel;
wire main_sram_bus_cyc;
wire main_sram_bus_stb;
reg main_sram_bus_ack = 1'd0;
wire main_sram_bus_we;
wire [2:0] main_sram_bus_cti;
wire [1:0] main_sram_bus_bte;
reg main_sram_bus_err = 1'd0;
wire [9:0] main_sram_adr;
wire [31:0] main_sram_dat_r;
reg [3:0] main_sram_we = 4'd0;
wire [31:0] main_sram_dat_w;
reg [31:0] main_uart_storage = 32'd9895604;
reg main_uart_sink_valid = 1'd0;
reg main_uart_sink_ready = 1'd0;
wire main_uart_sink_last;
reg [7:0] main_uart_sink_payload_data = 8'd0;
reg main_uart_uart_clk_txen = 1'd0;
reg [31:0] main_uart_phase_accumulator_tx = 32'd0;
reg [7:0] main_uart_tx_reg = 8'd0;
reg [3:0] main_uart_tx_bitcount = 4'd0;
reg main_uart_tx_busy = 1'd0;
reg main_uart_source_valid = 1'd0;
wire main_uart_source_ready;
reg [7:0] main_uart_source_payload_data = 8'd0;
reg main_uart_uart_clk_rxen = 1'd0;
reg [31:0] main_uart_phase_accumulator_rx = 32'd0;
wire main_uart_rx;
reg main_uart_rx_r = 1'd0;
reg [7:0] main_uart_rx_reg = 8'd0;
reg [3:0] main_uart_rx_bitcount = 4'd0;
reg main_uart_rx_busy = 1'd0;
wire [29:0] main_uart_wishbone_adr;
wire [31:0] main_uart_wishbone_dat_w;
wire [31:0] main_uart_wishbone_dat_r;
wire [3:0] main_uart_wishbone_sel;
reg main_uart_wishbone_cyc = 1'd0;
reg main_uart_wishbone_stb = 1'd0;
wire main_uart_wishbone_ack;
reg main_uart_wishbone_we = 1'd0;
reg [2:0] main_uart_wishbone_cti = 3'd0;
reg [1:0] main_uart_wishbone_bte = 2'd0;
wire main_uart_wishbone_err;
reg [2:0] main_uart_byte_counter = 3'd0;
reg main_uart_byte_counter_reset = 1'd0;
reg main_uart_byte_counter_ce = 1'd0;
reg [2:0] main_uart_word_counter = 3'd0;
reg main_uart_word_counter_reset = 1'd0;
reg main_uart_word_counter_ce = 1'd0;
reg [7:0] main_uart_cmd = 8'd0;
reg main_uart_cmd_ce = 1'd0;
reg [7:0] main_uart_length = 8'd0;
reg main_uart_length_ce = 1'd0;
reg [31:0] main_uart_address = 32'd0;
reg main_uart_address_ce = 1'd0;
reg [31:0] main_uart_data = 32'd0;
reg main_uart_rx_data_ce = 1'd0;
reg main_uart_tx_data_ce = 1'd0;
wire main_uart_reset;
wire main_uart_wait;
wire main_uart_done;
reg [22:0] main_uart_count = 23'd5000000;
reg main_uart_is_ongoing = 1'd0;
reg [31:0] main_load_storage = 32'd0;
reg main_load_re = 1'd0;
reg [31:0] main_reload_storage = 32'd0;
reg main_reload_re = 1'd0;
reg main_en_storage = 1'd0;
reg main_en_re = 1'd0;
reg main_update_value_storage = 1'd0;
reg main_update_value_re = 1'd0;
reg [31:0] main_value_status = 32'd0;
wire main_value_we;
wire main_irq;
wire main_zero_status;
reg main_zero_pending = 1'd0;
wire main_zero_trigger;
reg main_zero_clear = 1'd0;
reg main_zero_old_trigger = 1'd0;
wire main_eventmanager_status_re;
wire main_eventmanager_status_r;
wire main_eventmanager_status_we;
wire main_eventmanager_status_w;
wire main_eventmanager_pending_re;
wire main_eventmanager_pending_r;
wire main_eventmanager_pending_we;
wire main_eventmanager_pending_w;
reg main_eventmanager_storage = 1'd0;
reg main_eventmanager_re = 1'd0;
reg [31:0] main_value = 32'd0;
reg [13:0] main_interface_adr = 14'd0;
reg main_interface_we = 1'd0;
wire [7:0] main_interface_dat_w;
wire [7:0] main_interface_dat_r;
wire [29:0] main_bus_wishbone_adr;
wire [31:0] main_bus_wishbone_dat_w;
wire [31:0] main_bus_wishbone_dat_r;
wire [3:0] main_bus_wishbone_sel;
wire main_bus_wishbone_cyc;
wire main_bus_wishbone_stb;
reg main_bus_wishbone_ack = 1'd0;
wire main_bus_wishbone_we;
wire [2:0] main_bus_wishbone_cti;
wire [1:0] main_bus_wishbone_bte;
reg main_bus_wishbone_err = 1'd0;
wire [29:0] main_interface0_wb_sdram_adr;
wire [31:0] main_interface0_wb_sdram_dat_w;
reg [31:0] main_interface0_wb_sdram_dat_r = 32'd0;
wire [3:0] main_interface0_wb_sdram_sel;
wire main_interface0_wb_sdram_cyc;
wire main_interface0_wb_sdram_stb;
reg main_interface0_wb_sdram_ack = 1'd0;
wire main_interface0_wb_sdram_we;
wire [2:0] main_interface0_wb_sdram_cti;
wire [1:0] main_interface0_wb_sdram_bte;
reg main_interface0_wb_sdram_err = 1'd0;
wire sys_clk;
wire sys_rst;
wire sys4x_clk;
wire sys4x_clkb;
wire sys4x_dqs_clk;
wire clk200_clk;
wire clk200_rst;
wire main_reset;
wire main_locked;
wire main_pll_clkin;
wire main_clkout0;
wire main_clkout_buf0;
wire main_clkout1;
wire main_clkout_buf1;
wire main_clkout2;
wire main_clkout_buf2;
wire main_clkout3;
wire main_clkout_buf3;
wire main_clkout_buf4;
reg [3:0] main_reset_counter = 4'd15;
reg main_ic_reset = 1'd1;
reg [4:0] main_a7ddrphy_half_sys8x_taps_storage = 5'd16;
reg main_a7ddrphy_half_sys8x_taps_re = 1'd0;
wire main_a7ddrphy_cdly_rst_re;
wire main_a7ddrphy_cdly_rst_r;
wire main_a7ddrphy_cdly_rst_we;
reg main_a7ddrphy_cdly_rst_w = 1'd0;
wire main_a7ddrphy_cdly_inc_re;
wire main_a7ddrphy_cdly_inc_r;
wire main_a7ddrphy_cdly_inc_we;
reg main_a7ddrphy_cdly_inc_w = 1'd0;
reg [1:0] main_a7ddrphy_dly_sel_storage = 2'd0;
reg main_a7ddrphy_dly_sel_re = 1'd0;
wire main_a7ddrphy_rdly_dq_rst_re;
wire main_a7ddrphy_rdly_dq_rst_r;
wire main_a7ddrphy_rdly_dq_rst_we;
reg main_a7ddrphy_rdly_dq_rst_w = 1'd0;
wire main_a7ddrphy_rdly_dq_inc_re;
wire main_a7ddrphy_rdly_dq_inc_r;
wire main_a7ddrphy_rdly_dq_inc_we;
reg main_a7ddrphy_rdly_dq_inc_w = 1'd0;
wire main_a7ddrphy_rdly_dq_bitslip_rst_re;
wire main_a7ddrphy_rdly_dq_bitslip_rst_r;
wire main_a7ddrphy_rdly_dq_bitslip_rst_we;
reg main_a7ddrphy_rdly_dq_bitslip_rst_w = 1'd0;
wire main_a7ddrphy_rdly_dq_bitslip_re;
wire main_a7ddrphy_rdly_dq_bitslip_r;
wire main_a7ddrphy_rdly_dq_bitslip_we;
reg main_a7ddrphy_rdly_dq_bitslip_w = 1'd0;
wire [13:0] main_a7ddrphy_dfi_p0_address;
wire [2:0] main_a7ddrphy_dfi_p0_bank;
wire main_a7ddrphy_dfi_p0_cas_n;
wire main_a7ddrphy_dfi_p0_cs_n;
wire main_a7ddrphy_dfi_p0_ras_n;
wire main_a7ddrphy_dfi_p0_we_n;
wire main_a7ddrphy_dfi_p0_cke;
wire main_a7ddrphy_dfi_p0_odt;
wire main_a7ddrphy_dfi_p0_reset_n;
wire main_a7ddrphy_dfi_p0_act_n;
wire [31:0] main_a7ddrphy_dfi_p0_wrdata;
wire main_a7ddrphy_dfi_p0_wrdata_en;
wire [3:0] main_a7ddrphy_dfi_p0_wrdata_mask;
wire main_a7ddrphy_dfi_p0_rddata_en;
reg [31:0] main_a7ddrphy_dfi_p0_rddata = 32'd0;
reg main_a7ddrphy_dfi_p0_rddata_valid = 1'd0;
wire [13:0] main_a7ddrphy_dfi_p1_address;
wire [2:0] main_a7ddrphy_dfi_p1_bank;
wire main_a7ddrphy_dfi_p1_cas_n;
wire main_a7ddrphy_dfi_p1_cs_n;
wire main_a7ddrphy_dfi_p1_ras_n;
wire main_a7ddrphy_dfi_p1_we_n;
wire main_a7ddrphy_dfi_p1_cke;
wire main_a7ddrphy_dfi_p1_odt;
wire main_a7ddrphy_dfi_p1_reset_n;
wire main_a7ddrphy_dfi_p1_act_n;
wire [31:0] main_a7ddrphy_dfi_p1_wrdata;
wire main_a7ddrphy_dfi_p1_wrdata_en;
wire [3:0] main_a7ddrphy_dfi_p1_wrdata_mask;
wire main_a7ddrphy_dfi_p1_rddata_en;
reg [31:0] main_a7ddrphy_dfi_p1_rddata = 32'd0;
reg main_a7ddrphy_dfi_p1_rddata_valid = 1'd0;
wire [13:0] main_a7ddrphy_dfi_p2_address;
wire [2:0] main_a7ddrphy_dfi_p2_bank;
wire main_a7ddrphy_dfi_p2_cas_n;
wire main_a7ddrphy_dfi_p2_cs_n;
wire main_a7ddrphy_dfi_p2_ras_n;
wire main_a7ddrphy_dfi_p2_we_n;
wire main_a7ddrphy_dfi_p2_cke;
wire main_a7ddrphy_dfi_p2_odt;
wire main_a7ddrphy_dfi_p2_reset_n;
wire main_a7ddrphy_dfi_p2_act_n;
wire [31:0] main_a7ddrphy_dfi_p2_wrdata;
wire main_a7ddrphy_dfi_p2_wrdata_en;
wire [3:0] main_a7ddrphy_dfi_p2_wrdata_mask;
wire main_a7ddrphy_dfi_p2_rddata_en;
reg [31:0] main_a7ddrphy_dfi_p2_rddata = 32'd0;
reg main_a7ddrphy_dfi_p2_rddata_valid = 1'd0;
wire [13:0] main_a7ddrphy_dfi_p3_address;
wire [2:0] main_a7ddrphy_dfi_p3_bank;
wire main_a7ddrphy_dfi_p3_cas_n;
wire main_a7ddrphy_dfi_p3_cs_n;
wire main_a7ddrphy_dfi_p3_ras_n;
wire main_a7ddrphy_dfi_p3_we_n;
wire main_a7ddrphy_dfi_p3_cke;
wire main_a7ddrphy_dfi_p3_odt;
wire main_a7ddrphy_dfi_p3_reset_n;
wire main_a7ddrphy_dfi_p3_act_n;
wire [31:0] main_a7ddrphy_dfi_p3_wrdata;
wire main_a7ddrphy_dfi_p3_wrdata_en;
wire [3:0] main_a7ddrphy_dfi_p3_wrdata_mask;
wire main_a7ddrphy_dfi_p3_rddata_en;
reg [31:0] main_a7ddrphy_dfi_p3_rddata = 32'd0;
reg main_a7ddrphy_dfi_p3_rddata_valid = 1'd0;
wire main_a7ddrphy_sd_clk_se_nodelay;
reg main_a7ddrphy_oe_dqs = 1'd0;
wire main_a7ddrphy_dqs_preamble;
wire main_a7ddrphy_dqs_postamble;
reg [7:0] main_a7ddrphy_dqs_serdes_pattern = 8'd85;
wire main_a7ddrphy_dqs_nodelay0;
wire main_a7ddrphy_dqs_t0;
wire main_a7ddrphy0;
wire main_a7ddrphy_dqs_nodelay1;
wire main_a7ddrphy_dqs_t1;
wire main_a7ddrphy1;
reg main_a7ddrphy_oe_dq = 1'd0;
wire main_a7ddrphy_dq_o_nodelay0;
wire main_a7ddrphy_dq_i_nodelay0;
wire main_a7ddrphy_dq_i_delayed0;
wire main_a7ddrphy_dq_t0;
wire [7:0] main_a7ddrphy_dq_i_data0;
wire [7:0] main_a7ddrphy_bitslip0_i;
reg [7:0] main_a7ddrphy_bitslip0_o = 8'd0;
reg [2:0] main_a7ddrphy_bitslip0_value = 3'd0;
reg [15:0] main_a7ddrphy_bitslip0_r = 16'd0;
wire main_a7ddrphy_dq_o_nodelay1;
wire main_a7ddrphy_dq_i_nodelay1;
wire main_a7ddrphy_dq_i_delayed1;
wire main_a7ddrphy_dq_t1;
wire [7:0] main_a7ddrphy_dq_i_data1;
wire [7:0] main_a7ddrphy_bitslip1_i;
reg [7:0] main_a7ddrphy_bitslip1_o = 8'd0;
reg [2:0] main_a7ddrphy_bitslip1_value = 3'd0;
reg [15:0] main_a7ddrphy_bitslip1_r = 16'd0;
wire main_a7ddrphy_dq_o_nodelay2;
wire main_a7ddrphy_dq_i_nodelay2;
wire main_a7ddrphy_dq_i_delayed2;
wire main_a7ddrphy_dq_t2;
wire [7:0] main_a7ddrphy_dq_i_data2;
wire [7:0] main_a7ddrphy_bitslip2_i;
reg [7:0] main_a7ddrphy_bitslip2_o = 8'd0;
reg [2:0] main_a7ddrphy_bitslip2_value = 3'd0;
reg [15:0] main_a7ddrphy_bitslip2_r = 16'd0;
wire main_a7ddrphy_dq_o_nodelay3;
wire main_a7ddrphy_dq_i_nodelay3;
wire main_a7ddrphy_dq_i_delayed3;
wire main_a7ddrphy_dq_t3;
wire [7:0] main_a7ddrphy_dq_i_data3;
wire [7:0] main_a7ddrphy_bitslip3_i;
reg [7:0] main_a7ddrphy_bitslip3_o = 8'd0;
reg [2:0] main_a7ddrphy_bitslip3_value = 3'd0;
reg [15:0] main_a7ddrphy_bitslip3_r = 16'd0;
wire main_a7ddrphy_dq_o_nodelay4;
wire main_a7ddrphy_dq_i_nodelay4;
wire main_a7ddrphy_dq_i_delayed4;
wire main_a7ddrphy_dq_t4;
wire [7:0] main_a7ddrphy_dq_i_data4;
wire [7:0] main_a7ddrphy_bitslip4_i;
reg [7:0] main_a7ddrphy_bitslip4_o = 8'd0;
reg [2:0] main_a7ddrphy_bitslip4_value = 3'd0;
reg [15:0] main_a7ddrphy_bitslip4_r = 16'd0;
wire main_a7ddrphy_dq_o_nodelay5;
wire main_a7ddrphy_dq_i_nodelay5;
wire main_a7ddrphy_dq_i_delayed5;
wire main_a7ddrphy_dq_t5;
wire [7:0] main_a7ddrphy_dq_i_data5;
wire [7:0] main_a7ddrphy_bitslip5_i;
reg [7:0] main_a7ddrphy_bitslip5_o = 8'd0;
reg [2:0] main_a7ddrphy_bitslip5_value = 3'd0;
reg [15:0] main_a7ddrphy_bitslip5_r = 16'd0;
wire main_a7ddrphy_dq_o_nodelay6;
wire main_a7ddrphy_dq_i_nodelay6;
wire main_a7ddrphy_dq_i_delayed6;
wire main_a7ddrphy_dq_t6;
wire [7:0] main_a7ddrphy_dq_i_data6;
wire [7:0] main_a7ddrphy_bitslip6_i;
reg [7:0] main_a7ddrphy_bitslip6_o = 8'd0;
reg [2:0] main_a7ddrphy_bitslip6_value = 3'd0;
reg [15:0] main_a7ddrphy_bitslip6_r = 16'd0;
wire main_a7ddrphy_dq_o_nodelay7;
wire main_a7ddrphy_dq_i_nodelay7;
wire main_a7ddrphy_dq_i_delayed7;
wire main_a7ddrphy_dq_t7;
wire [7:0] main_a7ddrphy_dq_i_data7;
wire [7:0] main_a7ddrphy_bitslip7_i;
reg [7:0] main_a7ddrphy_bitslip7_o = 8'd0;
reg [2:0] main_a7ddrphy_bitslip7_value = 3'd0;
reg [15:0] main_a7ddrphy_bitslip7_r = 16'd0;
wire main_a7ddrphy_dq_o_nodelay8;
wire main_a7ddrphy_dq_i_nodelay8;
wire main_a7ddrphy_dq_i_delayed8;
wire main_a7ddrphy_dq_t8;
wire [7:0] main_a7ddrphy_dq_i_data8;
wire [7:0] main_a7ddrphy_bitslip8_i;
reg [7:0] main_a7ddrphy_bitslip8_o = 8'd0;
reg [2:0] main_a7ddrphy_bitslip8_value = 3'd0;
reg [15:0] main_a7ddrphy_bitslip8_r = 16'd0;
wire main_a7ddrphy_dq_o_nodelay9;
wire main_a7ddrphy_dq_i_nodelay9;
wire main_a7ddrphy_dq_i_delayed9;
wire main_a7ddrphy_dq_t9;
wire [7:0] main_a7ddrphy_dq_i_data9;
wire [7:0] main_a7ddrphy_bitslip9_i;
reg [7:0] main_a7ddrphy_bitslip9_o = 8'd0;
reg [2:0] main_a7ddrphy_bitslip9_value = 3'd0;
reg [15:0] main_a7ddrphy_bitslip9_r = 16'd0;
wire main_a7ddrphy_dq_o_nodelay10;
wire main_a7ddrphy_dq_i_nodelay10;
wire main_a7ddrphy_dq_i_delayed10;
wire main_a7ddrphy_dq_t10;
wire [7:0] main_a7ddrphy_dq_i_data10;
wire [7:0] main_a7ddrphy_bitslip10_i;
reg [7:0] main_a7ddrphy_bitslip10_o = 8'd0;
reg [2:0] main_a7ddrphy_bitslip10_value = 3'd0;
reg [15:0] main_a7ddrphy_bitslip10_r = 16'd0;
wire main_a7ddrphy_dq_o_nodelay11;
wire main_a7ddrphy_dq_i_nodelay11;
wire main_a7ddrphy_dq_i_delayed11;
wire main_a7ddrphy_dq_t11;
wire [7:0] main_a7ddrphy_dq_i_data11;
wire [7:0] main_a7ddrphy_bitslip11_i;
reg [7:0] main_a7ddrphy_bitslip11_o = 8'd0;
reg [2:0] main_a7ddrphy_bitslip11_value = 3'd0;
reg [15:0] main_a7ddrphy_bitslip11_r = 16'd0;
wire main_a7ddrphy_dq_o_nodelay12;
wire main_a7ddrphy_dq_i_nodelay12;
wire main_a7ddrphy_dq_i_delayed12;
wire main_a7ddrphy_dq_t12;
wire [7:0] main_a7ddrphy_dq_i_data12;
wire [7:0] main_a7ddrphy_bitslip12_i;
reg [7:0] main_a7ddrphy_bitslip12_o = 8'd0;
reg [2:0] main_a7ddrphy_bitslip12_value = 3'd0;
reg [15:0] main_a7ddrphy_bitslip12_r = 16'd0;
wire main_a7ddrphy_dq_o_nodelay13;
wire main_a7ddrphy_dq_i_nodelay13;
wire main_a7ddrphy_dq_i_delayed13;
wire main_a7ddrphy_dq_t13;
wire [7:0] main_a7ddrphy_dq_i_data13;
wire [7:0] main_a7ddrphy_bitslip13_i;
reg [7:0] main_a7ddrphy_bitslip13_o = 8'd0;
reg [2:0] main_a7ddrphy_bitslip13_value = 3'd0;
reg [15:0] main_a7ddrphy_bitslip13_r = 16'd0;
wire main_a7ddrphy_dq_o_nodelay14;
wire main_a7ddrphy_dq_i_nodelay14;
wire main_a7ddrphy_dq_i_delayed14;
wire main_a7ddrphy_dq_t14;
wire [7:0] main_a7ddrphy_dq_i_data14;
wire [7:0] main_a7ddrphy_bitslip14_i;
reg [7:0] main_a7ddrphy_bitslip14_o = 8'd0;
reg [2:0] main_a7ddrphy_bitslip14_value = 3'd0;
reg [15:0] main_a7ddrphy_bitslip14_r = 16'd0;
wire main_a7ddrphy_dq_o_nodelay15;
wire main_a7ddrphy_dq_i_nodelay15;
wire main_a7ddrphy_dq_i_delayed15;
wire main_a7ddrphy_dq_t15;
wire [7:0] main_a7ddrphy_dq_i_data15;
wire [7:0] main_a7ddrphy_bitslip15_i;
reg [7:0] main_a7ddrphy_bitslip15_o = 8'd0;
reg [2:0] main_a7ddrphy_bitslip15_value = 3'd0;
reg [15:0] main_a7ddrphy_bitslip15_r = 16'd0;
reg main_a7ddrphy_n_rddata_en0 = 1'd0;
reg main_a7ddrphy_n_rddata_en1 = 1'd0;
reg main_a7ddrphy_n_rddata_en2 = 1'd0;
reg main_a7ddrphy_n_rddata_en3 = 1'd0;
reg main_a7ddrphy_n_rddata_en4 = 1'd0;
reg main_a7ddrphy_n_rddata_en5 = 1'd0;
reg main_a7ddrphy_n_rddata_en6 = 1'd0;
reg main_a7ddrphy_n_rddata_en7 = 1'd0;
wire main_a7ddrphy_oe;
reg [3:0] main_a7ddrphy_last_wrdata_en = 4'd0;
wire [13:0] main_sdram_inti_p0_address;
wire [2:0] main_sdram_inti_p0_bank;
reg main_sdram_inti_p0_cas_n = 1'd1;
reg main_sdram_inti_p0_cs_n = 1'd1;
reg main_sdram_inti_p0_ras_n = 1'd1;
reg main_sdram_inti_p0_we_n = 1'd1;
wire main_sdram_inti_p0_cke;
wire main_sdram_inti_p0_odt;
wire main_sdram_inti_p0_reset_n;
reg main_sdram_inti_p0_act_n = 1'd1;
wire [31:0] main_sdram_inti_p0_wrdata;
wire main_sdram_inti_p0_wrdata_en;
wire [3:0] main_sdram_inti_p0_wrdata_mask;
wire main_sdram_inti_p0_rddata_en;
reg [31:0] main_sdram_inti_p0_rddata = 32'd0;
reg main_sdram_inti_p0_rddata_valid = 1'd0;
wire [13:0] main_sdram_inti_p1_address;
wire [2:0] main_sdram_inti_p1_bank;
reg main_sdram_inti_p1_cas_n = 1'd1;
reg main_sdram_inti_p1_cs_n = 1'd1;
reg main_sdram_inti_p1_ras_n = 1'd1;
reg main_sdram_inti_p1_we_n = 1'd1;
wire main_sdram_inti_p1_cke;
wire main_sdram_inti_p1_odt;
wire main_sdram_inti_p1_reset_n;
reg main_sdram_inti_p1_act_n = 1'd1;
wire [31:0] main_sdram_inti_p1_wrdata;
wire main_sdram_inti_p1_wrdata_en;
wire [3:0] main_sdram_inti_p1_wrdata_mask;
wire main_sdram_inti_p1_rddata_en;
reg [31:0] main_sdram_inti_p1_rddata = 32'd0;
reg main_sdram_inti_p1_rddata_valid = 1'd0;
wire [13:0] main_sdram_inti_p2_address;
wire [2:0] main_sdram_inti_p2_bank;
reg main_sdram_inti_p2_cas_n = 1'd1;
reg main_sdram_inti_p2_cs_n = 1'd1;
reg main_sdram_inti_p2_ras_n = 1'd1;
reg main_sdram_inti_p2_we_n = 1'd1;
wire main_sdram_inti_p2_cke;
wire main_sdram_inti_p2_odt;
wire main_sdram_inti_p2_reset_n;
reg main_sdram_inti_p2_act_n = 1'd1;
wire [31:0] main_sdram_inti_p2_wrdata;
wire main_sdram_inti_p2_wrdata_en;
wire [3:0] main_sdram_inti_p2_wrdata_mask;
wire main_sdram_inti_p2_rddata_en;
reg [31:0] main_sdram_inti_p2_rddata = 32'd0;
reg main_sdram_inti_p2_rddata_valid = 1'd0;
wire [13:0] main_sdram_inti_p3_address;
wire [2:0] main_sdram_inti_p3_bank;
reg main_sdram_inti_p3_cas_n = 1'd1;
reg main_sdram_inti_p3_cs_n = 1'd1;
reg main_sdram_inti_p3_ras_n = 1'd1;
reg main_sdram_inti_p3_we_n = 1'd1;
wire main_sdram_inti_p3_cke;
wire main_sdram_inti_p3_odt;
wire main_sdram_inti_p3_reset_n;
reg main_sdram_inti_p3_act_n = 1'd1;
wire [31:0] main_sdram_inti_p3_wrdata;
wire main_sdram_inti_p3_wrdata_en;
wire [3:0] main_sdram_inti_p3_wrdata_mask;
wire main_sdram_inti_p3_rddata_en;
reg [31:0] main_sdram_inti_p3_rddata = 32'd0;
reg main_sdram_inti_p3_rddata_valid = 1'd0;
wire [13:0] main_sdram_slave_p0_address;
wire [2:0] main_sdram_slave_p0_bank;
wire main_sdram_slave_p0_cas_n;
wire main_sdram_slave_p0_cs_n;
wire main_sdram_slave_p0_ras_n;
wire main_sdram_slave_p0_we_n;
wire main_sdram_slave_p0_cke;
wire main_sdram_slave_p0_odt;
wire main_sdram_slave_p0_reset_n;
wire main_sdram_slave_p0_act_n;
wire [31:0] main_sdram_slave_p0_wrdata;
wire main_sdram_slave_p0_wrdata_en;
wire [3:0] main_sdram_slave_p0_wrdata_mask;
wire main_sdram_slave_p0_rddata_en;
reg [31:0] main_sdram_slave_p0_rddata = 32'd0;
reg main_sdram_slave_p0_rddata_valid = 1'd0;
wire [13:0] main_sdram_slave_p1_address;
wire [2:0] main_sdram_slave_p1_bank;
wire main_sdram_slave_p1_cas_n;
wire main_sdram_slave_p1_cs_n;
wire main_sdram_slave_p1_ras_n;
wire main_sdram_slave_p1_we_n;
wire main_sdram_slave_p1_cke;
wire main_sdram_slave_p1_odt;
wire main_sdram_slave_p1_reset_n;
wire main_sdram_slave_p1_act_n;
wire [31:0] main_sdram_slave_p1_wrdata;
wire main_sdram_slave_p1_wrdata_en;
wire [3:0] main_sdram_slave_p1_wrdata_mask;
wire main_sdram_slave_p1_rddata_en;
reg [31:0] main_sdram_slave_p1_rddata = 32'd0;
reg main_sdram_slave_p1_rddata_valid = 1'd0;
wire [13:0] main_sdram_slave_p2_address;
wire [2:0] main_sdram_slave_p2_bank;
wire main_sdram_slave_p2_cas_n;
wire main_sdram_slave_p2_cs_n;
wire main_sdram_slave_p2_ras_n;
wire main_sdram_slave_p2_we_n;
wire main_sdram_slave_p2_cke;
wire main_sdram_slave_p2_odt;
wire main_sdram_slave_p2_reset_n;
wire main_sdram_slave_p2_act_n;
wire [31:0] main_sdram_slave_p2_wrdata;
wire main_sdram_slave_p2_wrdata_en;
wire [3:0] main_sdram_slave_p2_wrdata_mask;
wire main_sdram_slave_p2_rddata_en;
reg [31:0] main_sdram_slave_p2_rddata = 32'd0;
reg main_sdram_slave_p2_rddata_valid = 1'd0;
wire [13:0] main_sdram_slave_p3_address;
wire [2:0] main_sdram_slave_p3_bank;
wire main_sdram_slave_p3_cas_n;
wire main_sdram_slave_p3_cs_n;
wire main_sdram_slave_p3_ras_n;
wire main_sdram_slave_p3_we_n;
wire main_sdram_slave_p3_cke;
wire main_sdram_slave_p3_odt;
wire main_sdram_slave_p3_reset_n;
wire main_sdram_slave_p3_act_n;
wire [31:0] main_sdram_slave_p3_wrdata;
wire main_sdram_slave_p3_wrdata_en;
wire [3:0] main_sdram_slave_p3_wrdata_mask;
wire main_sdram_slave_p3_rddata_en;
reg [31:0] main_sdram_slave_p3_rddata = 32'd0;
reg main_sdram_slave_p3_rddata_valid = 1'd0;
reg [13:0] main_sdram_master_p0_address = 14'd0;
reg [2:0] main_sdram_master_p0_bank = 3'd0;
reg main_sdram_master_p0_cas_n = 1'd1;
reg main_sdram_master_p0_cs_n = 1'd1;
reg main_sdram_master_p0_ras_n = 1'd1;
reg main_sdram_master_p0_we_n = 1'd1;
reg main_sdram_master_p0_cke = 1'd0;
reg main_sdram_master_p0_odt = 1'd0;
reg main_sdram_master_p0_reset_n = 1'd0;
reg main_sdram_master_p0_act_n = 1'd1;
reg [31:0] main_sdram_master_p0_wrdata = 32'd0;
reg main_sdram_master_p0_wrdata_en = 1'd0;
reg [3:0] main_sdram_master_p0_wrdata_mask = 4'd0;
reg main_sdram_master_p0_rddata_en = 1'd0;
wire [31:0] main_sdram_master_p0_rddata;
wire main_sdram_master_p0_rddata_valid;
reg [13:0] main_sdram_master_p1_address = 14'd0;
reg [2:0] main_sdram_master_p1_bank = 3'd0;
reg main_sdram_master_p1_cas_n = 1'd1;
reg main_sdram_master_p1_cs_n = 1'd1;
reg main_sdram_master_p1_ras_n = 1'd1;
reg main_sdram_master_p1_we_n = 1'd1;
reg main_sdram_master_p1_cke = 1'd0;
reg main_sdram_master_p1_odt = 1'd0;
reg main_sdram_master_p1_reset_n = 1'd0;
reg main_sdram_master_p1_act_n = 1'd1;
reg [31:0] main_sdram_master_p1_wrdata = 32'd0;
reg main_sdram_master_p1_wrdata_en = 1'd0;
reg [3:0] main_sdram_master_p1_wrdata_mask = 4'd0;
reg main_sdram_master_p1_rddata_en = 1'd0;
wire [31:0] main_sdram_master_p1_rddata;
wire main_sdram_master_p1_rddata_valid;
reg [13:0] main_sdram_master_p2_address = 14'd0;
reg [2:0] main_sdram_master_p2_bank = 3'd0;
reg main_sdram_master_p2_cas_n = 1'd1;
reg main_sdram_master_p2_cs_n = 1'd1;
reg main_sdram_master_p2_ras_n = 1'd1;
reg main_sdram_master_p2_we_n = 1'd1;
reg main_sdram_master_p2_cke = 1'd0;
reg main_sdram_master_p2_odt = 1'd0;
reg main_sdram_master_p2_reset_n = 1'd0;
reg main_sdram_master_p2_act_n = 1'd1;
reg [31:0] main_sdram_master_p2_wrdata = 32'd0;
reg main_sdram_master_p2_wrdata_en = 1'd0;
reg [3:0] main_sdram_master_p2_wrdata_mask = 4'd0;
reg main_sdram_master_p2_rddata_en = 1'd0;
wire [31:0] main_sdram_master_p2_rddata;
wire main_sdram_master_p2_rddata_valid;
reg [13:0] main_sdram_master_p3_address = 14'd0;
reg [2:0] main_sdram_master_p3_bank = 3'd0;
reg main_sdram_master_p3_cas_n = 1'd1;
reg main_sdram_master_p3_cs_n = 1'd1;
reg main_sdram_master_p3_ras_n = 1'd1;
reg main_sdram_master_p3_we_n = 1'd1;
reg main_sdram_master_p3_cke = 1'd0;
reg main_sdram_master_p3_odt = 1'd0;
reg main_sdram_master_p3_reset_n = 1'd0;
reg main_sdram_master_p3_act_n = 1'd1;
reg [31:0] main_sdram_master_p3_wrdata = 32'd0;
reg main_sdram_master_p3_wrdata_en = 1'd0;
reg [3:0] main_sdram_master_p3_wrdata_mask = 4'd0;
reg main_sdram_master_p3_rddata_en = 1'd0;
wire [31:0] main_sdram_master_p3_rddata;
wire main_sdram_master_p3_rddata_valid;
reg [3:0] main_sdram_storage = 4'd0;
reg main_sdram_re = 1'd0;
reg [5:0] main_sdram_phaseinjector0_command_storage = 6'd0;
reg main_sdram_phaseinjector0_command_re = 1'd0;
wire main_sdram_phaseinjector0_command_issue_re;
wire main_sdram_phaseinjector0_command_issue_r;
wire main_sdram_phaseinjector0_command_issue_we;
reg main_sdram_phaseinjector0_command_issue_w = 1'd0;
reg [13:0] main_sdram_phaseinjector0_address_storage = 14'd0;
reg main_sdram_phaseinjector0_address_re = 1'd0;
reg [2:0] main_sdram_phaseinjector0_baddress_storage = 3'd0;
reg main_sdram_phaseinjector0_baddress_re = 1'd0;
reg [31:0] main_sdram_phaseinjector0_wrdata_storage = 32'd0;
reg main_sdram_phaseinjector0_wrdata_re = 1'd0;
reg [31:0] main_sdram_phaseinjector0_status = 32'd0;
wire main_sdram_phaseinjector0_we;
reg [5:0] main_sdram_phaseinjector1_command_storage = 6'd0;
reg main_sdram_phaseinjector1_command_re = 1'd0;
wire main_sdram_phaseinjector1_command_issue_re;
wire main_sdram_phaseinjector1_command_issue_r;
wire main_sdram_phaseinjector1_command_issue_we;
reg main_sdram_phaseinjector1_command_issue_w = 1'd0;
reg [13:0] main_sdram_phaseinjector1_address_storage = 14'd0;
reg main_sdram_phaseinjector1_address_re = 1'd0;
reg [2:0] main_sdram_phaseinjector1_baddress_storage = 3'd0;
reg main_sdram_phaseinjector1_baddress_re = 1'd0;
reg [31:0] main_sdram_phaseinjector1_wrdata_storage = 32'd0;
reg main_sdram_phaseinjector1_wrdata_re = 1'd0;
reg [31:0] main_sdram_phaseinjector1_status = 32'd0;
wire main_sdram_phaseinjector1_we;
reg [5:0] main_sdram_phaseinjector2_command_storage = 6'd0;
reg main_sdram_phaseinjector2_command_re = 1'd0;
wire main_sdram_phaseinjector2_command_issue_re;
wire main_sdram_phaseinjector2_command_issue_r;
wire main_sdram_phaseinjector2_command_issue_we;
reg main_sdram_phaseinjector2_command_issue_w = 1'd0;
reg [13:0] main_sdram_phaseinjector2_address_storage = 14'd0;
reg main_sdram_phaseinjector2_address_re = 1'd0;
reg [2:0] main_sdram_phaseinjector2_baddress_storage = 3'd0;
reg main_sdram_phaseinjector2_baddress_re = 1'd0;
reg [31:0] main_sdram_phaseinjector2_wrdata_storage = 32'd0;
reg main_sdram_phaseinjector2_wrdata_re = 1'd0;
reg [31:0] main_sdram_phaseinjector2_status = 32'd0;
wire main_sdram_phaseinjector2_we;
reg [5:0] main_sdram_phaseinjector3_command_storage = 6'd0;
reg main_sdram_phaseinjector3_command_re = 1'd0;
wire main_sdram_phaseinjector3_command_issue_re;
wire main_sdram_phaseinjector3_command_issue_r;
wire main_sdram_phaseinjector3_command_issue_we;
reg main_sdram_phaseinjector3_command_issue_w = 1'd0;
reg [13:0] main_sdram_phaseinjector3_address_storage = 14'd0;
reg main_sdram_phaseinjector3_address_re = 1'd0;
reg [2:0] main_sdram_phaseinjector3_baddress_storage = 3'd0;
reg main_sdram_phaseinjector3_baddress_re = 1'd0;
reg [31:0] main_sdram_phaseinjector3_wrdata_storage = 32'd0;
reg main_sdram_phaseinjector3_wrdata_re = 1'd0;
reg [31:0] main_sdram_phaseinjector3_status = 32'd0;
wire main_sdram_phaseinjector3_we;
wire main_sdram_interface_bank0_valid;
wire main_sdram_interface_bank0_ready;
wire main_sdram_interface_bank0_we;
wire [20:0] main_sdram_interface_bank0_addr;
wire main_sdram_interface_bank0_lock;
wire main_sdram_interface_bank0_wdata_ready;
wire main_sdram_interface_bank0_rdata_valid;
wire main_sdram_interface_bank1_valid;
wire main_sdram_interface_bank1_ready;
wire main_sdram_interface_bank1_we;
wire [20:0] main_sdram_interface_bank1_addr;
wire main_sdram_interface_bank1_lock;
wire main_sdram_interface_bank1_wdata_ready;
wire main_sdram_interface_bank1_rdata_valid;
wire main_sdram_interface_bank2_valid;
wire main_sdram_interface_bank2_ready;
wire main_sdram_interface_bank2_we;
wire [20:0] main_sdram_interface_bank2_addr;
wire main_sdram_interface_bank2_lock;
wire main_sdram_interface_bank2_wdata_ready;
wire main_sdram_interface_bank2_rdata_valid;
wire main_sdram_interface_bank3_valid;
wire main_sdram_interface_bank3_ready;
wire main_sdram_interface_bank3_we;
wire [20:0] main_sdram_interface_bank3_addr;
wire main_sdram_interface_bank3_lock;
wire main_sdram_interface_bank3_wdata_ready;
wire main_sdram_interface_bank3_rdata_valid;
wire main_sdram_interface_bank4_valid;
wire main_sdram_interface_bank4_ready;
wire main_sdram_interface_bank4_we;
wire [20:0] main_sdram_interface_bank4_addr;
wire main_sdram_interface_bank4_lock;
wire main_sdram_interface_bank4_wdata_ready;
wire main_sdram_interface_bank4_rdata_valid;
wire main_sdram_interface_bank5_valid;
wire main_sdram_interface_bank5_ready;
wire main_sdram_interface_bank5_we;
wire [20:0] main_sdram_interface_bank5_addr;
wire main_sdram_interface_bank5_lock;
wire main_sdram_interface_bank5_wdata_ready;
wire main_sdram_interface_bank5_rdata_valid;
wire main_sdram_interface_bank6_valid;
wire main_sdram_interface_bank6_ready;
wire main_sdram_interface_bank6_we;
wire [20:0] main_sdram_interface_bank6_addr;
wire main_sdram_interface_bank6_lock;
wire main_sdram_interface_bank6_wdata_ready;
wire main_sdram_interface_bank6_rdata_valid;
wire main_sdram_interface_bank7_valid;
wire main_sdram_interface_bank7_ready;
wire main_sdram_interface_bank7_we;
wire [20:0] main_sdram_interface_bank7_addr;
wire main_sdram_interface_bank7_lock;
wire main_sdram_interface_bank7_wdata_ready;
wire main_sdram_interface_bank7_rdata_valid;
reg [127:0] main_sdram_interface_wdata = 128'd0;
reg [15:0] main_sdram_interface_wdata_we = 16'd0;
wire [127:0] main_sdram_interface_rdata;
reg [13:0] main_sdram_dfi_p0_address = 14'd0;
reg [2:0] main_sdram_dfi_p0_bank = 3'd0;
reg main_sdram_dfi_p0_cas_n = 1'd1;
reg main_sdram_dfi_p0_cs_n = 1'd1;
reg main_sdram_dfi_p0_ras_n = 1'd1;
reg main_sdram_dfi_p0_we_n = 1'd1;
wire main_sdram_dfi_p0_cke;
wire main_sdram_dfi_p0_odt;
wire main_sdram_dfi_p0_reset_n;
reg main_sdram_dfi_p0_act_n = 1'd1;
wire [31:0] main_sdram_dfi_p0_wrdata;
reg main_sdram_dfi_p0_wrdata_en = 1'd0;
wire [3:0] main_sdram_dfi_p0_wrdata_mask;
reg main_sdram_dfi_p0_rddata_en = 1'd0;
wire [31:0] main_sdram_dfi_p0_rddata;
wire main_sdram_dfi_p0_rddata_valid;
reg [13:0] main_sdram_dfi_p1_address = 14'd0;
reg [2:0] main_sdram_dfi_p1_bank = 3'd0;
reg main_sdram_dfi_p1_cas_n = 1'd1;
reg main_sdram_dfi_p1_cs_n = 1'd1;
reg main_sdram_dfi_p1_ras_n = 1'd1;
reg main_sdram_dfi_p1_we_n = 1'd1;
wire main_sdram_dfi_p1_cke;
wire main_sdram_dfi_p1_odt;
wire main_sdram_dfi_p1_reset_n;
reg main_sdram_dfi_p1_act_n = 1'd1;
wire [31:0] main_sdram_dfi_p1_wrdata;
reg main_sdram_dfi_p1_wrdata_en = 1'd0;
wire [3:0] main_sdram_dfi_p1_wrdata_mask;
reg main_sdram_dfi_p1_rddata_en = 1'd0;
wire [31:0] main_sdram_dfi_p1_rddata;
wire main_sdram_dfi_p1_rddata_valid;
reg [13:0] main_sdram_dfi_p2_address = 14'd0;
reg [2:0] main_sdram_dfi_p2_bank = 3'd0;
reg main_sdram_dfi_p2_cas_n = 1'd1;
reg main_sdram_dfi_p2_cs_n = 1'd1;
reg main_sdram_dfi_p2_ras_n = 1'd1;
reg main_sdram_dfi_p2_we_n = 1'd1;
wire main_sdram_dfi_p2_cke;
wire main_sdram_dfi_p2_odt;
wire main_sdram_dfi_p2_reset_n;
reg main_sdram_dfi_p2_act_n = 1'd1;
wire [31:0] main_sdram_dfi_p2_wrdata;
reg main_sdram_dfi_p2_wrdata_en = 1'd0;
wire [3:0] main_sdram_dfi_p2_wrdata_mask;
reg main_sdram_dfi_p2_rddata_en = 1'd0;
wire [31:0] main_sdram_dfi_p2_rddata;
wire main_sdram_dfi_p2_rddata_valid;
reg [13:0] main_sdram_dfi_p3_address = 14'd0;
reg [2:0] main_sdram_dfi_p3_bank = 3'd0;
reg main_sdram_dfi_p3_cas_n = 1'd1;
reg main_sdram_dfi_p3_cs_n = 1'd1;
reg main_sdram_dfi_p3_ras_n = 1'd1;
reg main_sdram_dfi_p3_we_n = 1'd1;
wire main_sdram_dfi_p3_cke;
wire main_sdram_dfi_p3_odt;
wire main_sdram_dfi_p3_reset_n;
reg main_sdram_dfi_p3_act_n = 1'd1;
wire [31:0] main_sdram_dfi_p3_wrdata;
reg main_sdram_dfi_p3_wrdata_en = 1'd0;
wire [3:0] main_sdram_dfi_p3_wrdata_mask;
reg main_sdram_dfi_p3_rddata_en = 1'd0;
wire [31:0] main_sdram_dfi_p3_rddata;
wire main_sdram_dfi_p3_rddata_valid;
reg main_sdram_cmd_valid = 1'd0;
reg main_sdram_cmd_ready = 1'd0;
reg main_sdram_cmd_last = 1'd0;
reg [13:0] main_sdram_cmd_payload_a = 14'd0;
reg [2:0] main_sdram_cmd_payload_ba = 3'd0;
reg main_sdram_cmd_payload_cas = 1'd0;
reg main_sdram_cmd_payload_ras = 1'd0;
reg main_sdram_cmd_payload_we = 1'd0;
reg main_sdram_cmd_payload_is_read = 1'd0;
reg main_sdram_cmd_payload_is_write = 1'd0;
wire main_sdram_wants_refresh;
wire main_sdram_wants_zqcs;
wire main_sdram_timer_wait;
wire main_sdram_timer_done0;
wire [8:0] main_sdram_timer_count0;
wire main_sdram_timer_done1;
reg [8:0] main_sdram_timer_count1 = 9'd390;
wire main_sdram_postponer_req_i;
reg main_sdram_postponer_req_o = 1'd0;
reg main_sdram_postponer_count = 1'd0;
reg main_sdram_sequencer_start0 = 1'd0;
wire main_sdram_sequencer_done0;
wire main_sdram_sequencer_start1;
reg main_sdram_sequencer_done1 = 1'd0;
reg [5:0] main_sdram_sequencer_counter = 6'd0;
reg main_sdram_sequencer_count = 1'd0;
wire main_sdram_zqcs_timer_wait;
wire main_sdram_zqcs_timer_done0;
wire [25:0] main_sdram_zqcs_timer_count0;
wire main_sdram_zqcs_timer_done1;
reg [25:0] main_sdram_zqcs_timer_count1 = 26'd49999999;
reg main_sdram_zqcs_executer_start = 1'd0;
reg main_sdram_zqcs_executer_done = 1'd0;
reg [4:0] main_sdram_zqcs_executer_counter = 5'd0;
wire main_sdram_bankmachine0_req_valid;
wire main_sdram_bankmachine0_req_ready;
wire main_sdram_bankmachine0_req_we;
wire [20:0] main_sdram_bankmachine0_req_addr;
wire main_sdram_bankmachine0_req_lock;
reg main_sdram_bankmachine0_req_wdata_ready = 1'd0;
reg main_sdram_bankmachine0_req_rdata_valid = 1'd0;
wire main_sdram_bankmachine0_refresh_req;
reg main_sdram_bankmachine0_refresh_gnt = 1'd0;
reg main_sdram_bankmachine0_cmd_valid = 1'd0;
reg main_sdram_bankmachine0_cmd_ready = 1'd0;
reg [13:0] main_sdram_bankmachine0_cmd_payload_a = 14'd0;
wire [2:0] main_sdram_bankmachine0_cmd_payload_ba;
reg main_sdram_bankmachine0_cmd_payload_cas = 1'd0;
reg main_sdram_bankmachine0_cmd_payload_ras = 1'd0;
reg main_sdram_bankmachine0_cmd_payload_we = 1'd0;
reg main_sdram_bankmachine0_cmd_payload_is_cmd = 1'd0;
reg main_sdram_bankmachine0_cmd_payload_is_read = 1'd0;
reg main_sdram_bankmachine0_cmd_payload_is_write = 1'd0;
reg main_sdram_bankmachine0_auto_precharge = 1'd0;
wire main_sdram_bankmachine0_cmd_buffer_lookahead_sink_valid;
wire main_sdram_bankmachine0_cmd_buffer_lookahead_sink_ready;
reg main_sdram_bankmachine0_cmd_buffer_lookahead_sink_first = 1'd0;
reg main_sdram_bankmachine0_cmd_buffer_lookahead_sink_last = 1'd0;
wire main_sdram_bankmachine0_cmd_buffer_lookahead_sink_payload_we;
wire [20:0] main_sdram_bankmachine0_cmd_buffer_lookahead_sink_payload_addr;
wire main_sdram_bankmachine0_cmd_buffer_lookahead_source_valid;
wire main_sdram_bankmachine0_cmd_buffer_lookahead_source_ready;
wire main_sdram_bankmachine0_cmd_buffer_lookahead_source_first;
wire main_sdram_bankmachine0_cmd_buffer_lookahead_source_last;
wire main_sdram_bankmachine0_cmd_buffer_lookahead_source_payload_we;
wire [20:0] main_sdram_bankmachine0_cmd_buffer_lookahead_source_payload_addr;
wire main_sdram_bankmachine0_cmd_buffer_lookahead_syncfifo0_we;
wire main_sdram_bankmachine0_cmd_buffer_lookahead_syncfifo0_writable;
wire main_sdram_bankmachine0_cmd_buffer_lookahead_syncfifo0_re;
wire main_sdram_bankmachine0_cmd_buffer_lookahead_syncfifo0_readable;
wire [23:0] main_sdram_bankmachine0_cmd_buffer_lookahead_syncfifo0_din;
wire [23:0] main_sdram_bankmachine0_cmd_buffer_lookahead_syncfifo0_dout;
reg [3:0] main_sdram_bankmachine0_cmd_buffer_lookahead_level = 4'd0;
reg main_sdram_bankmachine0_cmd_buffer_lookahead_replace = 1'd0;
reg [2:0] main_sdram_bankmachine0_cmd_buffer_lookahead_produce = 3'd0;
reg [2:0] main_sdram_bankmachine0_cmd_buffer_lookahead_consume = 3'd0;
reg [2:0] main_sdram_bankmachine0_cmd_buffer_lookahead_wrport_adr = 3'd0;
wire [23:0] main_sdram_bankmachine0_cmd_buffer_lookahead_wrport_dat_r;
wire main_sdram_bankmachine0_cmd_buffer_lookahead_wrport_we;
wire [23:0] main_sdram_bankmachine0_cmd_buffer_lookahead_wrport_dat_w;
wire main_sdram_bankmachine0_cmd_buffer_lookahead_do_read;
wire [2:0] main_sdram_bankmachine0_cmd_buffer_lookahead_rdport_adr;
wire [23:0] main_sdram_bankmachine0_cmd_buffer_lookahead_rdport_dat_r;
wire main_sdram_bankmachine0_cmd_buffer_lookahead_fifo_in_payload_we;
wire [20:0] main_sdram_bankmachine0_cmd_buffer_lookahead_fifo_in_payload_addr;
wire main_sdram_bankmachine0_cmd_buffer_lookahead_fifo_in_first;
wire main_sdram_bankmachine0_cmd_buffer_lookahead_fifo_in_last;
wire main_sdram_bankmachine0_cmd_buffer_lookahead_fifo_out_payload_we;
wire [20:0] main_sdram_bankmachine0_cmd_buffer_lookahead_fifo_out_payload_addr;
wire main_sdram_bankmachine0_cmd_buffer_lookahead_fifo_out_first;
wire main_sdram_bankmachine0_cmd_buffer_lookahead_fifo_out_last;
wire main_sdram_bankmachine0_cmd_buffer_sink_valid;
wire main_sdram_bankmachine0_cmd_buffer_sink_ready;
wire main_sdram_bankmachine0_cmd_buffer_sink_first;
wire main_sdram_bankmachine0_cmd_buffer_sink_last;
wire main_sdram_bankmachine0_cmd_buffer_sink_payload_we;
wire [20:0] main_sdram_bankmachine0_cmd_buffer_sink_payload_addr;
reg main_sdram_bankmachine0_cmd_buffer_source_valid = 1'd0;
wire main_sdram_bankmachine0_cmd_buffer_source_ready;
reg main_sdram_bankmachine0_cmd_buffer_source_first = 1'd0;
reg main_sdram_bankmachine0_cmd_buffer_source_last = 1'd0;
reg main_sdram_bankmachine0_cmd_buffer_source_payload_we = 1'd0;
reg [20:0] main_sdram_bankmachine0_cmd_buffer_source_payload_addr = 21'd0;
reg [13:0] main_sdram_bankmachine0_row = 14'd0;
reg main_sdram_bankmachine0_row_opened = 1'd0;
wire main_sdram_bankmachine0_row_hit;
reg main_sdram_bankmachine0_row_open = 1'd0;
reg main_sdram_bankmachine0_row_close = 1'd0;
reg main_sdram_bankmachine0_row_col_n_addr_sel = 1'd0;
wire main_sdram_bankmachine0_twtpcon_valid;
(* dont_touch = "true" *) reg main_sdram_bankmachine0_twtpcon_ready = 1'd1;
reg [2:0] main_sdram_bankmachine0_twtpcon_count = 3'd0;
wire main_sdram_bankmachine0_trccon_valid;
(* dont_touch = "true" *) reg main_sdram_bankmachine0_trccon_ready = 1'd1;
reg [1:0] main_sdram_bankmachine0_trccon_count = 2'd0;
wire main_sdram_bankmachine0_trascon_valid;
(* dont_touch = "true" *) reg main_sdram_bankmachine0_trascon_ready = 1'd1;
reg [1:0] main_sdram_bankmachine0_trascon_count = 2'd0;
wire main_sdram_bankmachine1_req_valid;
wire main_sdram_bankmachine1_req_ready;
wire main_sdram_bankmachine1_req_we;
wire [20:0] main_sdram_bankmachine1_req_addr;
wire main_sdram_bankmachine1_req_lock;
reg main_sdram_bankmachine1_req_wdata_ready = 1'd0;
reg main_sdram_bankmachine1_req_rdata_valid = 1'd0;
wire main_sdram_bankmachine1_refresh_req;
reg main_sdram_bankmachine1_refresh_gnt = 1'd0;
reg main_sdram_bankmachine1_cmd_valid = 1'd0;
reg main_sdram_bankmachine1_cmd_ready = 1'd0;
reg [13:0] main_sdram_bankmachine1_cmd_payload_a = 14'd0;
wire [2:0] main_sdram_bankmachine1_cmd_payload_ba;
reg main_sdram_bankmachine1_cmd_payload_cas = 1'd0;
reg main_sdram_bankmachine1_cmd_payload_ras = 1'd0;
reg main_sdram_bankmachine1_cmd_payload_we = 1'd0;
reg main_sdram_bankmachine1_cmd_payload_is_cmd = 1'd0;
reg main_sdram_bankmachine1_cmd_payload_is_read = 1'd0;
reg main_sdram_bankmachine1_cmd_payload_is_write = 1'd0;
reg main_sdram_bankmachine1_auto_precharge = 1'd0;
wire main_sdram_bankmachine1_cmd_buffer_lookahead_sink_valid;
wire main_sdram_bankmachine1_cmd_buffer_lookahead_sink_ready;
reg main_sdram_bankmachine1_cmd_buffer_lookahead_sink_first = 1'd0;
reg main_sdram_bankmachine1_cmd_buffer_lookahead_sink_last = 1'd0;
wire main_sdram_bankmachine1_cmd_buffer_lookahead_sink_payload_we;
wire [20:0] main_sdram_bankmachine1_cmd_buffer_lookahead_sink_payload_addr;
wire main_sdram_bankmachine1_cmd_buffer_lookahead_source_valid;
wire main_sdram_bankmachine1_cmd_buffer_lookahead_source_ready;
wire main_sdram_bankmachine1_cmd_buffer_lookahead_source_first;
wire main_sdram_bankmachine1_cmd_buffer_lookahead_source_last;
wire main_sdram_bankmachine1_cmd_buffer_lookahead_source_payload_we;
wire [20:0] main_sdram_bankmachine1_cmd_buffer_lookahead_source_payload_addr;
wire main_sdram_bankmachine1_cmd_buffer_lookahead_syncfifo1_we;
wire main_sdram_bankmachine1_cmd_buffer_lookahead_syncfifo1_writable;
wire main_sdram_bankmachine1_cmd_buffer_lookahead_syncfifo1_re;
wire main_sdram_bankmachine1_cmd_buffer_lookahead_syncfifo1_readable;
wire [23:0] main_sdram_bankmachine1_cmd_buffer_lookahead_syncfifo1_din;
wire [23:0] main_sdram_bankmachine1_cmd_buffer_lookahead_syncfifo1_dout;
reg [3:0] main_sdram_bankmachine1_cmd_buffer_lookahead_level = 4'd0;
reg main_sdram_bankmachine1_cmd_buffer_lookahead_replace = 1'd0;
reg [2:0] main_sdram_bankmachine1_cmd_buffer_lookahead_produce = 3'd0;
reg [2:0] main_sdram_bankmachine1_cmd_buffer_lookahead_consume = 3'd0;
reg [2:0] main_sdram_bankmachine1_cmd_buffer_lookahead_wrport_adr = 3'd0;
wire [23:0] main_sdram_bankmachine1_cmd_buffer_lookahead_wrport_dat_r;
wire main_sdram_bankmachine1_cmd_buffer_lookahead_wrport_we;
wire [23:0] main_sdram_bankmachine1_cmd_buffer_lookahead_wrport_dat_w;
wire main_sdram_bankmachine1_cmd_buffer_lookahead_do_read;
wire [2:0] main_sdram_bankmachine1_cmd_buffer_lookahead_rdport_adr;
wire [23:0] main_sdram_bankmachine1_cmd_buffer_lookahead_rdport_dat_r;
wire main_sdram_bankmachine1_cmd_buffer_lookahead_fifo_in_payload_we;
wire [20:0] main_sdram_bankmachine1_cmd_buffer_lookahead_fifo_in_payload_addr;
wire main_sdram_bankmachine1_cmd_buffer_lookahead_fifo_in_first;
wire main_sdram_bankmachine1_cmd_buffer_lookahead_fifo_in_last;
wire main_sdram_bankmachine1_cmd_buffer_lookahead_fifo_out_payload_we;
wire [20:0] main_sdram_bankmachine1_cmd_buffer_lookahead_fifo_out_payload_addr;
wire main_sdram_bankmachine1_cmd_buffer_lookahead_fifo_out_first;
wire main_sdram_bankmachine1_cmd_buffer_lookahead_fifo_out_last;
wire main_sdram_bankmachine1_cmd_buffer_sink_valid;
wire main_sdram_bankmachine1_cmd_buffer_sink_ready;
wire main_sdram_bankmachine1_cmd_buffer_sink_first;
wire main_sdram_bankmachine1_cmd_buffer_sink_last;
wire main_sdram_bankmachine1_cmd_buffer_sink_payload_we;
wire [20:0] main_sdram_bankmachine1_cmd_buffer_sink_payload_addr;
reg main_sdram_bankmachine1_cmd_buffer_source_valid = 1'd0;
wire main_sdram_bankmachine1_cmd_buffer_source_ready;
reg main_sdram_bankmachine1_cmd_buffer_source_first = 1'd0;
reg main_sdram_bankmachine1_cmd_buffer_source_last = 1'd0;
reg main_sdram_bankmachine1_cmd_buffer_source_payload_we = 1'd0;
reg [20:0] main_sdram_bankmachine1_cmd_buffer_source_payload_addr = 21'd0;
reg [13:0] main_sdram_bankmachine1_row = 14'd0;
reg main_sdram_bankmachine1_row_opened = 1'd0;
wire main_sdram_bankmachine1_row_hit;
reg main_sdram_bankmachine1_row_open = 1'd0;
reg main_sdram_bankmachine1_row_close = 1'd0;
reg main_sdram_bankmachine1_row_col_n_addr_sel = 1'd0;
wire main_sdram_bankmachine1_twtpcon_valid;
(* dont_touch = "true" *) reg main_sdram_bankmachine1_twtpcon_ready = 1'd1;
reg [2:0] main_sdram_bankmachine1_twtpcon_count = 3'd0;
wire main_sdram_bankmachine1_trccon_valid;
(* dont_touch = "true" *) reg main_sdram_bankmachine1_trccon_ready = 1'd1;
reg [1:0] main_sdram_bankmachine1_trccon_count = 2'd0;
wire main_sdram_bankmachine1_trascon_valid;
(* dont_touch = "true" *) reg main_sdram_bankmachine1_trascon_ready = 1'd1;
reg [1:0] main_sdram_bankmachine1_trascon_count = 2'd0;
wire main_sdram_bankmachine2_req_valid;
wire main_sdram_bankmachine2_req_ready;
wire main_sdram_bankmachine2_req_we;
wire [20:0] main_sdram_bankmachine2_req_addr;
wire main_sdram_bankmachine2_req_lock;
reg main_sdram_bankmachine2_req_wdata_ready = 1'd0;
reg main_sdram_bankmachine2_req_rdata_valid = 1'd0;
wire main_sdram_bankmachine2_refresh_req;
reg main_sdram_bankmachine2_refresh_gnt = 1'd0;
reg main_sdram_bankmachine2_cmd_valid = 1'd0;
reg main_sdram_bankmachine2_cmd_ready = 1'd0;
reg [13:0] main_sdram_bankmachine2_cmd_payload_a = 14'd0;
wire [2:0] main_sdram_bankmachine2_cmd_payload_ba;
reg main_sdram_bankmachine2_cmd_payload_cas = 1'd0;
reg main_sdram_bankmachine2_cmd_payload_ras = 1'd0;
reg main_sdram_bankmachine2_cmd_payload_we = 1'd0;
reg main_sdram_bankmachine2_cmd_payload_is_cmd = 1'd0;
reg main_sdram_bankmachine2_cmd_payload_is_read = 1'd0;
reg main_sdram_bankmachine2_cmd_payload_is_write = 1'd0;
reg main_sdram_bankmachine2_auto_precharge = 1'd0;
wire main_sdram_bankmachine2_cmd_buffer_lookahead_sink_valid;
wire main_sdram_bankmachine2_cmd_buffer_lookahead_sink_ready;
reg main_sdram_bankmachine2_cmd_buffer_lookahead_sink_first = 1'd0;
reg main_sdram_bankmachine2_cmd_buffer_lookahead_sink_last = 1'd0;
wire main_sdram_bankmachine2_cmd_buffer_lookahead_sink_payload_we;
wire [20:0] main_sdram_bankmachine2_cmd_buffer_lookahead_sink_payload_addr;
wire main_sdram_bankmachine2_cmd_buffer_lookahead_source_valid;
wire main_sdram_bankmachine2_cmd_buffer_lookahead_source_ready;
wire main_sdram_bankmachine2_cmd_buffer_lookahead_source_first;
wire main_sdram_bankmachine2_cmd_buffer_lookahead_source_last;
wire main_sdram_bankmachine2_cmd_buffer_lookahead_source_payload_we;
wire [20:0] main_sdram_bankmachine2_cmd_buffer_lookahead_source_payload_addr;
wire main_sdram_bankmachine2_cmd_buffer_lookahead_syncfifo2_we;
wire main_sdram_bankmachine2_cmd_buffer_lookahead_syncfifo2_writable;
wire main_sdram_bankmachine2_cmd_buffer_lookahead_syncfifo2_re;
wire main_sdram_bankmachine2_cmd_buffer_lookahead_syncfifo2_readable;
wire [23:0] main_sdram_bankmachine2_cmd_buffer_lookahead_syncfifo2_din;
wire [23:0] main_sdram_bankmachine2_cmd_buffer_lookahead_syncfifo2_dout;
reg [3:0] main_sdram_bankmachine2_cmd_buffer_lookahead_level = 4'd0;
reg main_sdram_bankmachine2_cmd_buffer_lookahead_replace = 1'd0;
reg [2:0] main_sdram_bankmachine2_cmd_buffer_lookahead_produce = 3'd0;
reg [2:0] main_sdram_bankmachine2_cmd_buffer_lookahead_consume = 3'd0;
reg [2:0] main_sdram_bankmachine2_cmd_buffer_lookahead_wrport_adr = 3'd0;
wire [23:0] main_sdram_bankmachine2_cmd_buffer_lookahead_wrport_dat_r;
wire main_sdram_bankmachine2_cmd_buffer_lookahead_wrport_we;
wire [23:0] main_sdram_bankmachine2_cmd_buffer_lookahead_wrport_dat_w;
wire main_sdram_bankmachine2_cmd_buffer_lookahead_do_read;
wire [2:0] main_sdram_bankmachine2_cmd_buffer_lookahead_rdport_adr;
wire [23:0] main_sdram_bankmachine2_cmd_buffer_lookahead_rdport_dat_r;
wire main_sdram_bankmachine2_cmd_buffer_lookahead_fifo_in_payload_we;
wire [20:0] main_sdram_bankmachine2_cmd_buffer_lookahead_fifo_in_payload_addr;
wire main_sdram_bankmachine2_cmd_buffer_lookahead_fifo_in_first;
wire main_sdram_bankmachine2_cmd_buffer_lookahead_fifo_in_last;
wire main_sdram_bankmachine2_cmd_buffer_lookahead_fifo_out_payload_we;
wire [20:0] main_sdram_bankmachine2_cmd_buffer_lookahead_fifo_out_payload_addr;
wire main_sdram_bankmachine2_cmd_buffer_lookahead_fifo_out_first;
wire main_sdram_bankmachine2_cmd_buffer_lookahead_fifo_out_last;
wire main_sdram_bankmachine2_cmd_buffer_sink_valid;
wire main_sdram_bankmachine2_cmd_buffer_sink_ready;
wire main_sdram_bankmachine2_cmd_buffer_sink_first;
wire main_sdram_bankmachine2_cmd_buffer_sink_last;
wire main_sdram_bankmachine2_cmd_buffer_sink_payload_we;
wire [20:0] main_sdram_bankmachine2_cmd_buffer_sink_payload_addr;
reg main_sdram_bankmachine2_cmd_buffer_source_valid = 1'd0;
wire main_sdram_bankmachine2_cmd_buffer_source_ready;
reg main_sdram_bankmachine2_cmd_buffer_source_first = 1'd0;
reg main_sdram_bankmachine2_cmd_buffer_source_last = 1'd0;
reg main_sdram_bankmachine2_cmd_buffer_source_payload_we = 1'd0;
reg [20:0] main_sdram_bankmachine2_cmd_buffer_source_payload_addr = 21'd0;
reg [13:0] main_sdram_bankmachine2_row = 14'd0;
reg main_sdram_bankmachine2_row_opened = 1'd0;
wire main_sdram_bankmachine2_row_hit;
reg main_sdram_bankmachine2_row_open = 1'd0;
reg main_sdram_bankmachine2_row_close = 1'd0;
reg main_sdram_bankmachine2_row_col_n_addr_sel = 1'd0;
wire main_sdram_bankmachine2_twtpcon_valid;
(* dont_touch = "true" *) reg main_sdram_bankmachine2_twtpcon_ready = 1'd1;
reg [2:0] main_sdram_bankmachine2_twtpcon_count = 3'd0;
wire main_sdram_bankmachine2_trccon_valid;
(* dont_touch = "true" *) reg main_sdram_bankmachine2_trccon_ready = 1'd1;
reg [1:0] main_sdram_bankmachine2_trccon_count = 2'd0;
wire main_sdram_bankmachine2_trascon_valid;
(* dont_touch = "true" *) reg main_sdram_bankmachine2_trascon_ready = 1'd1;
reg [1:0] main_sdram_bankmachine2_trascon_count = 2'd0;
wire main_sdram_bankmachine3_req_valid;
wire main_sdram_bankmachine3_req_ready;
wire main_sdram_bankmachine3_req_we;
wire [20:0] main_sdram_bankmachine3_req_addr;
wire main_sdram_bankmachine3_req_lock;
reg main_sdram_bankmachine3_req_wdata_ready = 1'd0;
reg main_sdram_bankmachine3_req_rdata_valid = 1'd0;
wire main_sdram_bankmachine3_refresh_req;
reg main_sdram_bankmachine3_refresh_gnt = 1'd0;
reg main_sdram_bankmachine3_cmd_valid = 1'd0;
reg main_sdram_bankmachine3_cmd_ready = 1'd0;
reg [13:0] main_sdram_bankmachine3_cmd_payload_a = 14'd0;
wire [2:0] main_sdram_bankmachine3_cmd_payload_ba;
reg main_sdram_bankmachine3_cmd_payload_cas = 1'd0;
reg main_sdram_bankmachine3_cmd_payload_ras = 1'd0;
reg main_sdram_bankmachine3_cmd_payload_we = 1'd0;
reg main_sdram_bankmachine3_cmd_payload_is_cmd = 1'd0;
reg main_sdram_bankmachine3_cmd_payload_is_read = 1'd0;
reg main_sdram_bankmachine3_cmd_payload_is_write = 1'd0;
reg main_sdram_bankmachine3_auto_precharge = 1'd0;
wire main_sdram_bankmachine3_cmd_buffer_lookahead_sink_valid;
wire main_sdram_bankmachine3_cmd_buffer_lookahead_sink_ready;
reg main_sdram_bankmachine3_cmd_buffer_lookahead_sink_first = 1'd0;
reg main_sdram_bankmachine3_cmd_buffer_lookahead_sink_last = 1'd0;
wire main_sdram_bankmachine3_cmd_buffer_lookahead_sink_payload_we;
wire [20:0] main_sdram_bankmachine3_cmd_buffer_lookahead_sink_payload_addr;
wire main_sdram_bankmachine3_cmd_buffer_lookahead_source_valid;
wire main_sdram_bankmachine3_cmd_buffer_lookahead_source_ready;
wire main_sdram_bankmachine3_cmd_buffer_lookahead_source_first;
wire main_sdram_bankmachine3_cmd_buffer_lookahead_source_last;
wire main_sdram_bankmachine3_cmd_buffer_lookahead_source_payload_we;
wire [20:0] main_sdram_bankmachine3_cmd_buffer_lookahead_source_payload_addr;
wire main_sdram_bankmachine3_cmd_buffer_lookahead_syncfifo3_we;
wire main_sdram_bankmachine3_cmd_buffer_lookahead_syncfifo3_writable;
wire main_sdram_bankmachine3_cmd_buffer_lookahead_syncfifo3_re;
wire main_sdram_bankmachine3_cmd_buffer_lookahead_syncfifo3_readable;
wire [23:0] main_sdram_bankmachine3_cmd_buffer_lookahead_syncfifo3_din;
wire [23:0] main_sdram_bankmachine3_cmd_buffer_lookahead_syncfifo3_dout;
reg [3:0] main_sdram_bankmachine3_cmd_buffer_lookahead_level = 4'd0;
reg main_sdram_bankmachine3_cmd_buffer_lookahead_replace = 1'd0;
reg [2:0] main_sdram_bankmachine3_cmd_buffer_lookahead_produce = 3'd0;
reg [2:0] main_sdram_bankmachine3_cmd_buffer_lookahead_consume = 3'd0;
reg [2:0] main_sdram_bankmachine3_cmd_buffer_lookahead_wrport_adr = 3'd0;
wire [23:0] main_sdram_bankmachine3_cmd_buffer_lookahead_wrport_dat_r;
wire main_sdram_bankmachine3_cmd_buffer_lookahead_wrport_we;
wire [23:0] main_sdram_bankmachine3_cmd_buffer_lookahead_wrport_dat_w;
wire main_sdram_bankmachine3_cmd_buffer_lookahead_do_read;
wire [2:0] main_sdram_bankmachine3_cmd_buffer_lookahead_rdport_adr;
wire [23:0] main_sdram_bankmachine3_cmd_buffer_lookahead_rdport_dat_r;
wire main_sdram_bankmachine3_cmd_buffer_lookahead_fifo_in_payload_we;
wire [20:0] main_sdram_bankmachine3_cmd_buffer_lookahead_fifo_in_payload_addr;
wire main_sdram_bankmachine3_cmd_buffer_lookahead_fifo_in_first;
wire main_sdram_bankmachine3_cmd_buffer_lookahead_fifo_in_last;
wire main_sdram_bankmachine3_cmd_buffer_lookahead_fifo_out_payload_we;
wire [20:0] main_sdram_bankmachine3_cmd_buffer_lookahead_fifo_out_payload_addr;
wire main_sdram_bankmachine3_cmd_buffer_lookahead_fifo_out_first;
wire main_sdram_bankmachine3_cmd_buffer_lookahead_fifo_out_last;
wire main_sdram_bankmachine3_cmd_buffer_sink_valid;
wire main_sdram_bankmachine3_cmd_buffer_sink_ready;
wire main_sdram_bankmachine3_cmd_buffer_sink_first;
wire main_sdram_bankmachine3_cmd_buffer_sink_last;
wire main_sdram_bankmachine3_cmd_buffer_sink_payload_we;
wire [20:0] main_sdram_bankmachine3_cmd_buffer_sink_payload_addr;
reg main_sdram_bankmachine3_cmd_buffer_source_valid = 1'd0;
wire main_sdram_bankmachine3_cmd_buffer_source_ready;
reg main_sdram_bankmachine3_cmd_buffer_source_first = 1'd0;
reg main_sdram_bankmachine3_cmd_buffer_source_last = 1'd0;
reg main_sdram_bankmachine3_cmd_buffer_source_payload_we = 1'd0;
reg [20:0] main_sdram_bankmachine3_cmd_buffer_source_payload_addr = 21'd0;
reg [13:0] main_sdram_bankmachine3_row = 14'd0;
reg main_sdram_bankmachine3_row_opened = 1'd0;
wire main_sdram_bankmachine3_row_hit;
reg main_sdram_bankmachine3_row_open = 1'd0;
reg main_sdram_bankmachine3_row_close = 1'd0;
reg main_sdram_bankmachine3_row_col_n_addr_sel = 1'd0;
wire main_sdram_bankmachine3_twtpcon_valid;
(* dont_touch = "true" *) reg main_sdram_bankmachine3_twtpcon_ready = 1'd1;
reg [2:0] main_sdram_bankmachine3_twtpcon_count = 3'd0;
wire main_sdram_bankmachine3_trccon_valid;
(* dont_touch = "true" *) reg main_sdram_bankmachine3_trccon_ready = 1'd1;
reg [1:0] main_sdram_bankmachine3_trccon_count = 2'd0;
wire main_sdram_bankmachine3_trascon_valid;
(* dont_touch = "true" *) reg main_sdram_bankmachine3_trascon_ready = 1'd1;
reg [1:0] main_sdram_bankmachine3_trascon_count = 2'd0;
wire main_sdram_bankmachine4_req_valid;
wire main_sdram_bankmachine4_req_ready;
wire main_sdram_bankmachine4_req_we;
wire [20:0] main_sdram_bankmachine4_req_addr;
wire main_sdram_bankmachine4_req_lock;
reg main_sdram_bankmachine4_req_wdata_ready = 1'd0;
reg main_sdram_bankmachine4_req_rdata_valid = 1'd0;
wire main_sdram_bankmachine4_refresh_req;
reg main_sdram_bankmachine4_refresh_gnt = 1'd0;
reg main_sdram_bankmachine4_cmd_valid = 1'd0;
reg main_sdram_bankmachine4_cmd_ready = 1'd0;
reg [13:0] main_sdram_bankmachine4_cmd_payload_a = 14'd0;
wire [2:0] main_sdram_bankmachine4_cmd_payload_ba;
reg main_sdram_bankmachine4_cmd_payload_cas = 1'd0;
reg main_sdram_bankmachine4_cmd_payload_ras = 1'd0;
reg main_sdram_bankmachine4_cmd_payload_we = 1'd0;
reg main_sdram_bankmachine4_cmd_payload_is_cmd = 1'd0;
reg main_sdram_bankmachine4_cmd_payload_is_read = 1'd0;
reg main_sdram_bankmachine4_cmd_payload_is_write = 1'd0;
reg main_sdram_bankmachine4_auto_precharge = 1'd0;
wire main_sdram_bankmachine4_cmd_buffer_lookahead_sink_valid;
wire main_sdram_bankmachine4_cmd_buffer_lookahead_sink_ready;
reg main_sdram_bankmachine4_cmd_buffer_lookahead_sink_first = 1'd0;
reg main_sdram_bankmachine4_cmd_buffer_lookahead_sink_last = 1'd0;
wire main_sdram_bankmachine4_cmd_buffer_lookahead_sink_payload_we;
wire [20:0] main_sdram_bankmachine4_cmd_buffer_lookahead_sink_payload_addr;
wire main_sdram_bankmachine4_cmd_buffer_lookahead_source_valid;
wire main_sdram_bankmachine4_cmd_buffer_lookahead_source_ready;
wire main_sdram_bankmachine4_cmd_buffer_lookahead_source_first;
wire main_sdram_bankmachine4_cmd_buffer_lookahead_source_last;
wire main_sdram_bankmachine4_cmd_buffer_lookahead_source_payload_we;
wire [20:0] main_sdram_bankmachine4_cmd_buffer_lookahead_source_payload_addr;
wire main_sdram_bankmachine4_cmd_buffer_lookahead_syncfifo4_we;
wire main_sdram_bankmachine4_cmd_buffer_lookahead_syncfifo4_writable;
wire main_sdram_bankmachine4_cmd_buffer_lookahead_syncfifo4_re;
wire main_sdram_bankmachine4_cmd_buffer_lookahead_syncfifo4_readable;
wire [23:0] main_sdram_bankmachine4_cmd_buffer_lookahead_syncfifo4_din;
wire [23:0] main_sdram_bankmachine4_cmd_buffer_lookahead_syncfifo4_dout;
reg [3:0] main_sdram_bankmachine4_cmd_buffer_lookahead_level = 4'd0;
reg main_sdram_bankmachine4_cmd_buffer_lookahead_replace = 1'd0;
reg [2:0] main_sdram_bankmachine4_cmd_buffer_lookahead_produce = 3'd0;
reg [2:0] main_sdram_bankmachine4_cmd_buffer_lookahead_consume = 3'd0;
reg [2:0] main_sdram_bankmachine4_cmd_buffer_lookahead_wrport_adr = 3'd0;
wire [23:0] main_sdram_bankmachine4_cmd_buffer_lookahead_wrport_dat_r;
wire main_sdram_bankmachine4_cmd_buffer_lookahead_wrport_we;
wire [23:0] main_sdram_bankmachine4_cmd_buffer_lookahead_wrport_dat_w;
wire main_sdram_bankmachine4_cmd_buffer_lookahead_do_read;
wire [2:0] main_sdram_bankmachine4_cmd_buffer_lookahead_rdport_adr;
wire [23:0] main_sdram_bankmachine4_cmd_buffer_lookahead_rdport_dat_r;
wire main_sdram_bankmachine4_cmd_buffer_lookahead_fifo_in_payload_we;
wire [20:0] main_sdram_bankmachine4_cmd_buffer_lookahead_fifo_in_payload_addr;
wire main_sdram_bankmachine4_cmd_buffer_lookahead_fifo_in_first;
wire main_sdram_bankmachine4_cmd_buffer_lookahead_fifo_in_last;
wire main_sdram_bankmachine4_cmd_buffer_lookahead_fifo_out_payload_we;
wire [20:0] main_sdram_bankmachine4_cmd_buffer_lookahead_fifo_out_payload_addr;
wire main_sdram_bankmachine4_cmd_buffer_lookahead_fifo_out_first;
wire main_sdram_bankmachine4_cmd_buffer_lookahead_fifo_out_last;
wire main_sdram_bankmachine4_cmd_buffer_sink_valid;
wire main_sdram_bankmachine4_cmd_buffer_sink_ready;
wire main_sdram_bankmachine4_cmd_buffer_sink_first;
wire main_sdram_bankmachine4_cmd_buffer_sink_last;
wire main_sdram_bankmachine4_cmd_buffer_sink_payload_we;
wire [20:0] main_sdram_bankmachine4_cmd_buffer_sink_payload_addr;
reg main_sdram_bankmachine4_cmd_buffer_source_valid = 1'd0;
wire main_sdram_bankmachine4_cmd_buffer_source_ready;
reg main_sdram_bankmachine4_cmd_buffer_source_first = 1'd0;
reg main_sdram_bankmachine4_cmd_buffer_source_last = 1'd0;
reg main_sdram_bankmachine4_cmd_buffer_source_payload_we = 1'd0;
reg [20:0] main_sdram_bankmachine4_cmd_buffer_source_payload_addr = 21'd0;
reg [13:0] main_sdram_bankmachine4_row = 14'd0;
reg main_sdram_bankmachine4_row_opened = 1'd0;
wire main_sdram_bankmachine4_row_hit;
reg main_sdram_bankmachine4_row_open = 1'd0;
reg main_sdram_bankmachine4_row_close = 1'd0;
reg main_sdram_bankmachine4_row_col_n_addr_sel = 1'd0;
wire main_sdram_bankmachine4_twtpcon_valid;
(* dont_touch = "true" *) reg main_sdram_bankmachine4_twtpcon_ready = 1'd1;
reg [2:0] main_sdram_bankmachine4_twtpcon_count = 3'd0;
wire main_sdram_bankmachine4_trccon_valid;
(* dont_touch = "true" *) reg main_sdram_bankmachine4_trccon_ready = 1'd1;
reg [1:0] main_sdram_bankmachine4_trccon_count = 2'd0;
wire main_sdram_bankmachine4_trascon_valid;
(* dont_touch = "true" *) reg main_sdram_bankmachine4_trascon_ready = 1'd1;
reg [1:0] main_sdram_bankmachine4_trascon_count = 2'd0;
wire main_sdram_bankmachine5_req_valid;
wire main_sdram_bankmachine5_req_ready;
wire main_sdram_bankmachine5_req_we;
wire [20:0] main_sdram_bankmachine5_req_addr;
wire main_sdram_bankmachine5_req_lock;
reg main_sdram_bankmachine5_req_wdata_ready = 1'd0;
reg main_sdram_bankmachine5_req_rdata_valid = 1'd0;
wire main_sdram_bankmachine5_refresh_req;
reg main_sdram_bankmachine5_refresh_gnt = 1'd0;
reg main_sdram_bankmachine5_cmd_valid = 1'd0;
reg main_sdram_bankmachine5_cmd_ready = 1'd0;
reg [13:0] main_sdram_bankmachine5_cmd_payload_a = 14'd0;
wire [2:0] main_sdram_bankmachine5_cmd_payload_ba;
reg main_sdram_bankmachine5_cmd_payload_cas = 1'd0;
reg main_sdram_bankmachine5_cmd_payload_ras = 1'd0;
reg main_sdram_bankmachine5_cmd_payload_we = 1'd0;
reg main_sdram_bankmachine5_cmd_payload_is_cmd = 1'd0;
reg main_sdram_bankmachine5_cmd_payload_is_read = 1'd0;
reg main_sdram_bankmachine5_cmd_payload_is_write = 1'd0;
reg main_sdram_bankmachine5_auto_precharge = 1'd0;
wire main_sdram_bankmachine5_cmd_buffer_lookahead_sink_valid;
wire main_sdram_bankmachine5_cmd_buffer_lookahead_sink_ready;
reg main_sdram_bankmachine5_cmd_buffer_lookahead_sink_first = 1'd0;
reg main_sdram_bankmachine5_cmd_buffer_lookahead_sink_last = 1'd0;
wire main_sdram_bankmachine5_cmd_buffer_lookahead_sink_payload_we;
wire [20:0] main_sdram_bankmachine5_cmd_buffer_lookahead_sink_payload_addr;
wire main_sdram_bankmachine5_cmd_buffer_lookahead_source_valid;
wire main_sdram_bankmachine5_cmd_buffer_lookahead_source_ready;
wire main_sdram_bankmachine5_cmd_buffer_lookahead_source_first;
wire main_sdram_bankmachine5_cmd_buffer_lookahead_source_last;
wire main_sdram_bankmachine5_cmd_buffer_lookahead_source_payload_we;
wire [20:0] main_sdram_bankmachine5_cmd_buffer_lookahead_source_payload_addr;
wire main_sdram_bankmachine5_cmd_buffer_lookahead_syncfifo5_we;
wire main_sdram_bankmachine5_cmd_buffer_lookahead_syncfifo5_writable;
wire main_sdram_bankmachine5_cmd_buffer_lookahead_syncfifo5_re;
wire main_sdram_bankmachine5_cmd_buffer_lookahead_syncfifo5_readable;
wire [23:0] main_sdram_bankmachine5_cmd_buffer_lookahead_syncfifo5_din;
wire [23:0] main_sdram_bankmachine5_cmd_buffer_lookahead_syncfifo5_dout;
reg [3:0] main_sdram_bankmachine5_cmd_buffer_lookahead_level = 4'd0;
reg main_sdram_bankmachine5_cmd_buffer_lookahead_replace = 1'd0;
reg [2:0] main_sdram_bankmachine5_cmd_buffer_lookahead_produce = 3'd0;
reg [2:0] main_sdram_bankmachine5_cmd_buffer_lookahead_consume = 3'd0;
reg [2:0] main_sdram_bankmachine5_cmd_buffer_lookahead_wrport_adr = 3'd0;
wire [23:0] main_sdram_bankmachine5_cmd_buffer_lookahead_wrport_dat_r;
wire main_sdram_bankmachine5_cmd_buffer_lookahead_wrport_we;
wire [23:0] main_sdram_bankmachine5_cmd_buffer_lookahead_wrport_dat_w;
wire main_sdram_bankmachine5_cmd_buffer_lookahead_do_read;
wire [2:0] main_sdram_bankmachine5_cmd_buffer_lookahead_rdport_adr;
wire [23:0] main_sdram_bankmachine5_cmd_buffer_lookahead_rdport_dat_r;
wire main_sdram_bankmachine5_cmd_buffer_lookahead_fifo_in_payload_we;
wire [20:0] main_sdram_bankmachine5_cmd_buffer_lookahead_fifo_in_payload_addr;
wire main_sdram_bankmachine5_cmd_buffer_lookahead_fifo_in_first;
wire main_sdram_bankmachine5_cmd_buffer_lookahead_fifo_in_last;
wire main_sdram_bankmachine5_cmd_buffer_lookahead_fifo_out_payload_we;
wire [20:0] main_sdram_bankmachine5_cmd_buffer_lookahead_fifo_out_payload_addr;
wire main_sdram_bankmachine5_cmd_buffer_lookahead_fifo_out_first;
wire main_sdram_bankmachine5_cmd_buffer_lookahead_fifo_out_last;
wire main_sdram_bankmachine5_cmd_buffer_sink_valid;
wire main_sdram_bankmachine5_cmd_buffer_sink_ready;
wire main_sdram_bankmachine5_cmd_buffer_sink_first;
wire main_sdram_bankmachine5_cmd_buffer_sink_last;
wire main_sdram_bankmachine5_cmd_buffer_sink_payload_we;
wire [20:0] main_sdram_bankmachine5_cmd_buffer_sink_payload_addr;
reg main_sdram_bankmachine5_cmd_buffer_source_valid = 1'd0;
wire main_sdram_bankmachine5_cmd_buffer_source_ready;
reg main_sdram_bankmachine5_cmd_buffer_source_first = 1'd0;
reg main_sdram_bankmachine5_cmd_buffer_source_last = 1'd0;
reg main_sdram_bankmachine5_cmd_buffer_source_payload_we = 1'd0;
reg [20:0] main_sdram_bankmachine5_cmd_buffer_source_payload_addr = 21'd0;
reg [13:0] main_sdram_bankmachine5_row = 14'd0;
reg main_sdram_bankmachine5_row_opened = 1'd0;
wire main_sdram_bankmachine5_row_hit;
reg main_sdram_bankmachine5_row_open = 1'd0;
reg main_sdram_bankmachine5_row_close = 1'd0;
reg main_sdram_bankmachine5_row_col_n_addr_sel = 1'd0;
wire main_sdram_bankmachine5_twtpcon_valid;
(* dont_touch = "true" *) reg main_sdram_bankmachine5_twtpcon_ready = 1'd1;
reg [2:0] main_sdram_bankmachine5_twtpcon_count = 3'd0;
wire main_sdram_bankmachine5_trccon_valid;
(* dont_touch = "true" *) reg main_sdram_bankmachine5_trccon_ready = 1'd1;
reg [1:0] main_sdram_bankmachine5_trccon_count = 2'd0;
wire main_sdram_bankmachine5_trascon_valid;
(* dont_touch = "true" *) reg main_sdram_bankmachine5_trascon_ready = 1'd1;
reg [1:0] main_sdram_bankmachine5_trascon_count = 2'd0;
wire main_sdram_bankmachine6_req_valid;
wire main_sdram_bankmachine6_req_ready;
wire main_sdram_bankmachine6_req_we;
wire [20:0] main_sdram_bankmachine6_req_addr;
wire main_sdram_bankmachine6_req_lock;
reg main_sdram_bankmachine6_req_wdata_ready = 1'd0;
reg main_sdram_bankmachine6_req_rdata_valid = 1'd0;
wire main_sdram_bankmachine6_refresh_req;
reg main_sdram_bankmachine6_refresh_gnt = 1'd0;
reg main_sdram_bankmachine6_cmd_valid = 1'd0;
reg main_sdram_bankmachine6_cmd_ready = 1'd0;
reg [13:0] main_sdram_bankmachine6_cmd_payload_a = 14'd0;
wire [2:0] main_sdram_bankmachine6_cmd_payload_ba;
reg main_sdram_bankmachine6_cmd_payload_cas = 1'd0;
reg main_sdram_bankmachine6_cmd_payload_ras = 1'd0;
reg main_sdram_bankmachine6_cmd_payload_we = 1'd0;
reg main_sdram_bankmachine6_cmd_payload_is_cmd = 1'd0;
reg main_sdram_bankmachine6_cmd_payload_is_read = 1'd0;
reg main_sdram_bankmachine6_cmd_payload_is_write = 1'd0;
reg main_sdram_bankmachine6_auto_precharge = 1'd0;
wire main_sdram_bankmachine6_cmd_buffer_lookahead_sink_valid;
wire main_sdram_bankmachine6_cmd_buffer_lookahead_sink_ready;
reg main_sdram_bankmachine6_cmd_buffer_lookahead_sink_first = 1'd0;
reg main_sdram_bankmachine6_cmd_buffer_lookahead_sink_last = 1'd0;
wire main_sdram_bankmachine6_cmd_buffer_lookahead_sink_payload_we;
wire [20:0] main_sdram_bankmachine6_cmd_buffer_lookahead_sink_payload_addr;
wire main_sdram_bankmachine6_cmd_buffer_lookahead_source_valid;
wire main_sdram_bankmachine6_cmd_buffer_lookahead_source_ready;
wire main_sdram_bankmachine6_cmd_buffer_lookahead_source_first;
wire main_sdram_bankmachine6_cmd_buffer_lookahead_source_last;
wire main_sdram_bankmachine6_cmd_buffer_lookahead_source_payload_we;
wire [20:0] main_sdram_bankmachine6_cmd_buffer_lookahead_source_payload_addr;
wire main_sdram_bankmachine6_cmd_buffer_lookahead_syncfifo6_we;
wire main_sdram_bankmachine6_cmd_buffer_lookahead_syncfifo6_writable;
wire main_sdram_bankmachine6_cmd_buffer_lookahead_syncfifo6_re;
wire main_sdram_bankmachine6_cmd_buffer_lookahead_syncfifo6_readable;
wire [23:0] main_sdram_bankmachine6_cmd_buffer_lookahead_syncfifo6_din;
wire [23:0] main_sdram_bankmachine6_cmd_buffer_lookahead_syncfifo6_dout;
reg [3:0] main_sdram_bankmachine6_cmd_buffer_lookahead_level = 4'd0;
reg main_sdram_bankmachine6_cmd_buffer_lookahead_replace = 1'd0;
reg [2:0] main_sdram_bankmachine6_cmd_buffer_lookahead_produce = 3'd0;
reg [2:0] main_sdram_bankmachine6_cmd_buffer_lookahead_consume = 3'd0;
reg [2:0] main_sdram_bankmachine6_cmd_buffer_lookahead_wrport_adr = 3'd0;
wire [23:0] main_sdram_bankmachine6_cmd_buffer_lookahead_wrport_dat_r;
wire main_sdram_bankmachine6_cmd_buffer_lookahead_wrport_we;
wire [23:0] main_sdram_bankmachine6_cmd_buffer_lookahead_wrport_dat_w;
wire main_sdram_bankmachine6_cmd_buffer_lookahead_do_read;
wire [2:0] main_sdram_bankmachine6_cmd_buffer_lookahead_rdport_adr;
wire [23:0] main_sdram_bankmachine6_cmd_buffer_lookahead_rdport_dat_r;
wire main_sdram_bankmachine6_cmd_buffer_lookahead_fifo_in_payload_we;
wire [20:0] main_sdram_bankmachine6_cmd_buffer_lookahead_fifo_in_payload_addr;
wire main_sdram_bankmachine6_cmd_buffer_lookahead_fifo_in_first;
wire main_sdram_bankmachine6_cmd_buffer_lookahead_fifo_in_last;
wire main_sdram_bankmachine6_cmd_buffer_lookahead_fifo_out_payload_we;
wire [20:0] main_sdram_bankmachine6_cmd_buffer_lookahead_fifo_out_payload_addr;
wire main_sdram_bankmachine6_cmd_buffer_lookahead_fifo_out_first;
wire main_sdram_bankmachine6_cmd_buffer_lookahead_fifo_out_last;
wire main_sdram_bankmachine6_cmd_buffer_sink_valid;
wire main_sdram_bankmachine6_cmd_buffer_sink_ready;
wire main_sdram_bankmachine6_cmd_buffer_sink_first;
wire main_sdram_bankmachine6_cmd_buffer_sink_last;
wire main_sdram_bankmachine6_cmd_buffer_sink_payload_we;
wire [20:0] main_sdram_bankmachine6_cmd_buffer_sink_payload_addr;
reg main_sdram_bankmachine6_cmd_buffer_source_valid = 1'd0;
wire main_sdram_bankmachine6_cmd_buffer_source_ready;
reg main_sdram_bankmachine6_cmd_buffer_source_first = 1'd0;
reg main_sdram_bankmachine6_cmd_buffer_source_last = 1'd0;
reg main_sdram_bankmachine6_cmd_buffer_source_payload_we = 1'd0;
reg [20:0] main_sdram_bankmachine6_cmd_buffer_source_payload_addr = 21'd0;
reg [13:0] main_sdram_bankmachine6_row = 14'd0;
reg main_sdram_bankmachine6_row_opened = 1'd0;
wire main_sdram_bankmachine6_row_hit;
reg main_sdram_bankmachine6_row_open = 1'd0;
reg main_sdram_bankmachine6_row_close = 1'd0;
reg main_sdram_bankmachine6_row_col_n_addr_sel = 1'd0;
wire main_sdram_bankmachine6_twtpcon_valid;
(* dont_touch = "true" *) reg main_sdram_bankmachine6_twtpcon_ready = 1'd1;
reg [2:0] main_sdram_bankmachine6_twtpcon_count = 3'd0;
wire main_sdram_bankmachine6_trccon_valid;
(* dont_touch = "true" *) reg main_sdram_bankmachine6_trccon_ready = 1'd1;
reg [1:0] main_sdram_bankmachine6_trccon_count = 2'd0;
wire main_sdram_bankmachine6_trascon_valid;
(* dont_touch = "true" *) reg main_sdram_bankmachine6_trascon_ready = 1'd1;
reg [1:0] main_sdram_bankmachine6_trascon_count = 2'd0;
wire main_sdram_bankmachine7_req_valid;
wire main_sdram_bankmachine7_req_ready;
wire main_sdram_bankmachine7_req_we;
wire [20:0] main_sdram_bankmachine7_req_addr;
wire main_sdram_bankmachine7_req_lock;
reg main_sdram_bankmachine7_req_wdata_ready = 1'd0;
reg main_sdram_bankmachine7_req_rdata_valid = 1'd0;
wire main_sdram_bankmachine7_refresh_req;
reg main_sdram_bankmachine7_refresh_gnt = 1'd0;
reg main_sdram_bankmachine7_cmd_valid = 1'd0;
reg main_sdram_bankmachine7_cmd_ready = 1'd0;
reg [13:0] main_sdram_bankmachine7_cmd_payload_a = 14'd0;
wire [2:0] main_sdram_bankmachine7_cmd_payload_ba;
reg main_sdram_bankmachine7_cmd_payload_cas = 1'd0;
reg main_sdram_bankmachine7_cmd_payload_ras = 1'd0;
reg main_sdram_bankmachine7_cmd_payload_we = 1'd0;
reg main_sdram_bankmachine7_cmd_payload_is_cmd = 1'd0;
reg main_sdram_bankmachine7_cmd_payload_is_read = 1'd0;
reg main_sdram_bankmachine7_cmd_payload_is_write = 1'd0;
reg main_sdram_bankmachine7_auto_precharge = 1'd0;
wire main_sdram_bankmachine7_cmd_buffer_lookahead_sink_valid;
wire main_sdram_bankmachine7_cmd_buffer_lookahead_sink_ready;
reg main_sdram_bankmachine7_cmd_buffer_lookahead_sink_first = 1'd0;
reg main_sdram_bankmachine7_cmd_buffer_lookahead_sink_last = 1'd0;
wire main_sdram_bankmachine7_cmd_buffer_lookahead_sink_payload_we;
wire [20:0] main_sdram_bankmachine7_cmd_buffer_lookahead_sink_payload_addr;
wire main_sdram_bankmachine7_cmd_buffer_lookahead_source_valid;
wire main_sdram_bankmachine7_cmd_buffer_lookahead_source_ready;
wire main_sdram_bankmachine7_cmd_buffer_lookahead_source_first;
wire main_sdram_bankmachine7_cmd_buffer_lookahead_source_last;
wire main_sdram_bankmachine7_cmd_buffer_lookahead_source_payload_we;
wire [20:0] main_sdram_bankmachine7_cmd_buffer_lookahead_source_payload_addr;
wire main_sdram_bankmachine7_cmd_buffer_lookahead_syncfifo7_we;
wire main_sdram_bankmachine7_cmd_buffer_lookahead_syncfifo7_writable;
wire main_sdram_bankmachine7_cmd_buffer_lookahead_syncfifo7_re;
wire main_sdram_bankmachine7_cmd_buffer_lookahead_syncfifo7_readable;
wire [23:0] main_sdram_bankmachine7_cmd_buffer_lookahead_syncfifo7_din;
wire [23:0] main_sdram_bankmachine7_cmd_buffer_lookahead_syncfifo7_dout;
reg [3:0] main_sdram_bankmachine7_cmd_buffer_lookahead_level = 4'd0;
reg main_sdram_bankmachine7_cmd_buffer_lookahead_replace = 1'd0;
reg [2:0] main_sdram_bankmachine7_cmd_buffer_lookahead_produce = 3'd0;
reg [2:0] main_sdram_bankmachine7_cmd_buffer_lookahead_consume = 3'd0;
reg [2:0] main_sdram_bankmachine7_cmd_buffer_lookahead_wrport_adr = 3'd0;
wire [23:0] main_sdram_bankmachine7_cmd_buffer_lookahead_wrport_dat_r;
wire main_sdram_bankmachine7_cmd_buffer_lookahead_wrport_we;
wire [23:0] main_sdram_bankmachine7_cmd_buffer_lookahead_wrport_dat_w;
wire main_sdram_bankmachine7_cmd_buffer_lookahead_do_read;
wire [2:0] main_sdram_bankmachine7_cmd_buffer_lookahead_rdport_adr;
wire [23:0] main_sdram_bankmachine7_cmd_buffer_lookahead_rdport_dat_r;
wire main_sdram_bankmachine7_cmd_buffer_lookahead_fifo_in_payload_we;
wire [20:0] main_sdram_bankmachine7_cmd_buffer_lookahead_fifo_in_payload_addr;
wire main_sdram_bankmachine7_cmd_buffer_lookahead_fifo_in_first;
wire main_sdram_bankmachine7_cmd_buffer_lookahead_fifo_in_last;
wire main_sdram_bankmachine7_cmd_buffer_lookahead_fifo_out_payload_we;
wire [20:0] main_sdram_bankmachine7_cmd_buffer_lookahead_fifo_out_payload_addr;
wire main_sdram_bankmachine7_cmd_buffer_lookahead_fifo_out_first;
wire main_sdram_bankmachine7_cmd_buffer_lookahead_fifo_out_last;
wire main_sdram_bankmachine7_cmd_buffer_sink_valid;
wire main_sdram_bankmachine7_cmd_buffer_sink_ready;
wire main_sdram_bankmachine7_cmd_buffer_sink_first;
wire main_sdram_bankmachine7_cmd_buffer_sink_last;
wire main_sdram_bankmachine7_cmd_buffer_sink_payload_we;
wire [20:0] main_sdram_bankmachine7_cmd_buffer_sink_payload_addr;
reg main_sdram_bankmachine7_cmd_buffer_source_valid = 1'd0;
wire main_sdram_bankmachine7_cmd_buffer_source_ready;
reg main_sdram_bankmachine7_cmd_buffer_source_first = 1'd0;
reg main_sdram_bankmachine7_cmd_buffer_source_last = 1'd0;
reg main_sdram_bankmachine7_cmd_buffer_source_payload_we = 1'd0;
reg [20:0] main_sdram_bankmachine7_cmd_buffer_source_payload_addr = 21'd0;
reg [13:0] main_sdram_bankmachine7_row = 14'd0;
reg main_sdram_bankmachine7_row_opened = 1'd0;
wire main_sdram_bankmachine7_row_hit;
reg main_sdram_bankmachine7_row_open = 1'd0;
reg main_sdram_bankmachine7_row_close = 1'd0;
reg main_sdram_bankmachine7_row_col_n_addr_sel = 1'd0;
wire main_sdram_bankmachine7_twtpcon_valid;
(* dont_touch = "true" *) reg main_sdram_bankmachine7_twtpcon_ready = 1'd1;
reg [2:0] main_sdram_bankmachine7_twtpcon_count = 3'd0;
wire main_sdram_bankmachine7_trccon_valid;
(* dont_touch = "true" *) reg main_sdram_bankmachine7_trccon_ready = 1'd1;
reg [1:0] main_sdram_bankmachine7_trccon_count = 2'd0;
wire main_sdram_bankmachine7_trascon_valid;
(* dont_touch = "true" *) reg main_sdram_bankmachine7_trascon_ready = 1'd1;
reg [1:0] main_sdram_bankmachine7_trascon_count = 2'd0;
wire main_sdram_ras_allowed;
wire main_sdram_cas_allowed;
reg main_sdram_choose_cmd_want_reads = 1'd0;
reg main_sdram_choose_cmd_want_writes = 1'd0;
reg main_sdram_choose_cmd_want_cmds = 1'd0;
reg main_sdram_choose_cmd_want_activates = 1'd0;
wire main_sdram_choose_cmd_cmd_valid;
reg main_sdram_choose_cmd_cmd_ready = 1'd0;
wire [13:0] main_sdram_choose_cmd_cmd_payload_a;
wire [2:0] main_sdram_choose_cmd_cmd_payload_ba;
reg main_sdram_choose_cmd_cmd_payload_cas = 1'd0;
reg main_sdram_choose_cmd_cmd_payload_ras = 1'd0;
reg main_sdram_choose_cmd_cmd_payload_we = 1'd0;
wire main_sdram_choose_cmd_cmd_payload_is_cmd;
wire main_sdram_choose_cmd_cmd_payload_is_read;
wire main_sdram_choose_cmd_cmd_payload_is_write;
reg [7:0] main_sdram_choose_cmd_valids = 8'd0;
wire [7:0] main_sdram_choose_cmd_request;
reg [2:0] main_sdram_choose_cmd_grant = 3'd0;
wire main_sdram_choose_cmd_ce;
reg main_sdram_choose_req_want_reads = 1'd0;
reg main_sdram_choose_req_want_writes = 1'd0;
reg main_sdram_choose_req_want_cmds = 1'd0;
reg main_sdram_choose_req_want_activates = 1'd0;
wire main_sdram_choose_req_cmd_valid;
reg main_sdram_choose_req_cmd_ready = 1'd0;
wire [13:0] main_sdram_choose_req_cmd_payload_a;
wire [2:0] main_sdram_choose_req_cmd_payload_ba;
reg main_sdram_choose_req_cmd_payload_cas = 1'd0;
reg main_sdram_choose_req_cmd_payload_ras = 1'd0;
reg main_sdram_choose_req_cmd_payload_we = 1'd0;
wire main_sdram_choose_req_cmd_payload_is_cmd;
wire main_sdram_choose_req_cmd_payload_is_read;
wire main_sdram_choose_req_cmd_payload_is_write;
reg [7:0] main_sdram_choose_req_valids = 8'd0;
wire [7:0] main_sdram_choose_req_request;
reg [2:0] main_sdram_choose_req_grant = 3'd0;
wire main_sdram_choose_req_ce;
reg [13:0] main_sdram_nop_a = 14'd0;
reg [2:0] main_sdram_nop_ba = 3'd0;
reg [1:0] main_sdram_steerer_sel0 = 2'd0;
reg [1:0] main_sdram_steerer_sel1 = 2'd0;
reg [1:0] main_sdram_steerer_sel2 = 2'd0;
reg [1:0] main_sdram_steerer_sel3 = 2'd0;
reg main_sdram_steerer0 = 1'd1;
reg main_sdram_steerer1 = 1'd1;
reg main_sdram_steerer2 = 1'd1;
reg main_sdram_steerer3 = 1'd1;
reg main_sdram_steerer4 = 1'd1;
reg main_sdram_steerer5 = 1'd1;
reg main_sdram_steerer6 = 1'd1;
reg main_sdram_steerer7 = 1'd1;
wire main_sdram_trrdcon_valid;
(* dont_touch = "true" *) reg main_sdram_trrdcon_ready = 1'd1;
reg main_sdram_trrdcon_count = 1'd0;
wire main_sdram_tfawcon_valid;
(* dont_touch = "true" *) reg main_sdram_tfawcon_ready = 1'd1;
wire [1:0] main_sdram_tfawcon_count;
reg [2:0] main_sdram_tfawcon_window = 3'd0;
wire main_sdram_tccdcon_valid;
(* dont_touch = "true" *) reg main_sdram_tccdcon_ready = 1'd1;
reg main_sdram_tccdcon_count = 1'd0;
wire main_sdram_twtrcon_valid;
(* dont_touch = "true" *) reg main_sdram_twtrcon_ready = 1'd1;
reg [2:0] main_sdram_twtrcon_count = 3'd0;
wire main_sdram_read_available;
wire main_sdram_write_available;
reg main_sdram_en0 = 1'd0;
wire main_sdram_max_time0;
reg [4:0] main_sdram_time0 = 5'd0;
reg main_sdram_en1 = 1'd0;
wire main_sdram_max_time1;
reg [3:0] main_sdram_time1 = 4'd0;
wire main_sdram_go_to_refresh;
reg main_port_cmd_valid = 1'd0;
wire main_port_cmd_ready;
reg main_port_cmd_payload_we = 1'd0;
reg [23:0] main_port_cmd_payload_addr = 24'd0;
wire main_port_wdata_valid;
wire main_port_wdata_ready;
wire main_port_wdata_first;
wire main_port_wdata_last;
wire [127:0] main_port_wdata_payload_data;
wire [15:0] main_port_wdata_payload_we;
wire main_port_rdata_valid;
wire main_port_rdata_ready;
reg main_port_rdata_first = 1'd0;
reg main_port_rdata_last = 1'd0;
wire [127:0] main_port_rdata_payload_data;
wire [29:0] main_interface1_wb_sdram_adr;
wire [31:0] main_interface1_wb_sdram_dat_w;
wire [31:0] main_interface1_wb_sdram_dat_r;
wire [3:0] main_interface1_wb_sdram_sel;
wire main_interface1_wb_sdram_cyc;
wire main_interface1_wb_sdram_stb;
wire main_interface1_wb_sdram_ack;
wire main_interface1_wb_sdram_we;
wire [2:0] main_interface1_wb_sdram_cti;
wire [1:0] main_interface1_wb_sdram_bte;
wire main_interface1_wb_sdram_err;
wire [29:0] main_adr;
wire [127:0] main_dat_w;
wire [127:0] main_dat_r;
wire [15:0] main_sel;
reg main_cyc = 1'd0;
reg main_stb = 1'd0;
reg main_ack = 1'd0;
reg main_we = 1'd0;
wire main_data_port_adr;
wire [127:0] main_data_port_dat_r;
reg [15:0] main_data_port_we = 16'd0;
reg [127:0] main_data_port_dat_w = 128'd0;
reg main_write_from_slave = 1'd0;
reg [1:0] main_adr_offset_r = 2'd0;
wire main_tag_port_adr;
wire [31:0] main_tag_port_dat_r;
reg main_tag_port_we = 1'd0;
wire [31:0] main_tag_port_dat_w;
wire [30:0] main_tag_do_tag;
wire main_tag_do_dirty;
wire [30:0] main_tag_di_tag;
reg main_tag_di_dirty = 1'd0;
reg main_word_clr = 1'd0;
reg main_word_inc = 1'd0;
wire main_wdata_converter_sink_valid;
wire main_wdata_converter_sink_ready;
reg main_wdata_converter_sink_first = 1'd0;
reg main_wdata_converter_sink_last = 1'd0;
wire [127:0] main_wdata_converter_sink_payload_data;
wire [15:0] main_wdata_converter_sink_payload_we;
wire main_wdata_converter_source_valid;
wire main_wdata_converter_source_ready;
wire main_wdata_converter_source_first;
wire main_wdata_converter_source_last;
wire [127:0] main_wdata_converter_source_payload_data;
wire [15:0] main_wdata_converter_source_payload_we;
wire main_wdata_converter_converter_sink_valid;
wire main_wdata_converter_converter_sink_ready;
wire main_wdata_converter_converter_sink_first;
wire main_wdata_converter_converter_sink_last;
wire [143:0] main_wdata_converter_converter_sink_payload_data;
wire main_wdata_converter_converter_source_valid;
wire main_wdata_converter_converter_source_ready;
wire main_wdata_converter_converter_source_first;
wire main_wdata_converter_converter_source_last;
wire [143:0] main_wdata_converter_converter_source_payload_data;
wire main_wdata_converter_converter_source_payload_valid_token_count;
wire main_wdata_converter_source_source_valid;
wire main_wdata_converter_source_source_ready;
wire main_wdata_converter_source_source_first;
wire main_wdata_converter_source_source_last;
wire [143:0] main_wdata_converter_source_source_payload_data;
wire main_rdata_converter_sink_valid;
wire main_rdata_converter_sink_ready;
wire main_rdata_converter_sink_first;
wire main_rdata_converter_sink_last;
wire [127:0] main_rdata_converter_sink_payload_data;
wire main_rdata_converter_source_valid;
wire main_rdata_converter_source_ready;
wire main_rdata_converter_source_first;
wire main_rdata_converter_source_last;
wire [127:0] main_rdata_converter_source_payload_data;
wire main_rdata_converter_converter_sink_valid;
wire main_rdata_converter_converter_sink_ready;
wire main_rdata_converter_converter_sink_first;
wire main_rdata_converter_converter_sink_last;
wire [127:0] main_rdata_converter_converter_sink_payload_data;
wire main_rdata_converter_converter_source_valid;
wire main_rdata_converter_converter_source_ready;
wire main_rdata_converter_converter_source_first;
wire main_rdata_converter_converter_source_last;
wire [127:0] main_rdata_converter_converter_source_payload_data;
wire main_rdata_converter_converter_source_payload_valid_token_count;
wire main_rdata_converter_source_source_valid;
wire main_rdata_converter_source_source_ready;
wire main_rdata_converter_source_source_first;
wire main_rdata_converter_source_source_last;
wire [127:0] main_rdata_converter_source_source_payload_data;
reg main_count = 1'd0;
reg [2:0] builder_uartwishbonebridge_state = 3'd0;
reg [2:0] builder_uartwishbonebridge_next_state = 3'd0;
reg builder_wb2csr_state = 1'd0;
reg builder_wb2csr_next_state = 1'd0;
wire builder_pll_fb;
reg [1:0] builder_refresher_state = 2'd0;
reg [1:0] builder_refresher_next_state = 2'd0;
reg [2:0] builder_bankmachine0_state = 3'd0;
reg [2:0] builder_bankmachine0_next_state = 3'd0;
reg [2:0] builder_bankmachine1_state = 3'd0;
reg [2:0] builder_bankmachine1_next_state = 3'd0;
reg [2:0] builder_bankmachine2_state = 3'd0;
reg [2:0] builder_bankmachine2_next_state = 3'd0;
reg [2:0] builder_bankmachine3_state = 3'd0;
reg [2:0] builder_bankmachine3_next_state = 3'd0;
reg [2:0] builder_bankmachine4_state = 3'd0;
reg [2:0] builder_bankmachine4_next_state = 3'd0;
reg [2:0] builder_bankmachine5_state = 3'd0;
reg [2:0] builder_bankmachine5_next_state = 3'd0;
reg [2:0] builder_bankmachine6_state = 3'd0;
reg [2:0] builder_bankmachine6_next_state = 3'd0;
reg [2:0] builder_bankmachine7_state = 3'd0;
reg [2:0] builder_bankmachine7_next_state = 3'd0;
reg [3:0] builder_multiplexer_state = 4'd0;
reg [3:0] builder_multiplexer_next_state = 4'd0;
wire builder_roundrobin0_request;
wire builder_roundrobin0_grant;
wire builder_roundrobin0_ce;
wire builder_roundrobin1_request;
wire builder_roundrobin1_grant;
wire builder_roundrobin1_ce;
wire builder_roundrobin2_request;
wire builder_roundrobin2_grant;
wire builder_roundrobin2_ce;
wire builder_roundrobin3_request;
wire builder_roundrobin3_grant;
wire builder_roundrobin3_ce;
wire builder_roundrobin4_request;
wire builder_roundrobin4_grant;
wire builder_roundrobin4_ce;
wire builder_roundrobin5_request;
wire builder_roundrobin5_grant;
wire builder_roundrobin5_ce;
wire builder_roundrobin6_request;
wire builder_roundrobin6_grant;
wire builder_roundrobin6_ce;
wire builder_roundrobin7_request;
wire builder_roundrobin7_grant;
wire builder_roundrobin7_ce;
reg [2:0] builder_rbank = 3'd0;
reg [2:0] builder_wbank = 3'd0;
reg builder_locked0 = 1'd0;
reg builder_locked1 = 1'd0;
reg builder_locked2 = 1'd0;
reg builder_locked3 = 1'd0;
reg builder_locked4 = 1'd0;
reg builder_locked5 = 1'd0;
reg builder_locked6 = 1'd0;
reg builder_locked7 = 1'd0;
reg builder_new_master_wdata_ready0 = 1'd0;
reg builder_new_master_wdata_ready1 = 1'd0;
reg builder_new_master_wdata_ready2 = 1'd0;
reg builder_new_master_rdata_valid0 = 1'd0;
reg builder_new_master_rdata_valid1 = 1'd0;
reg builder_new_master_rdata_valid2 = 1'd0;
reg builder_new_master_rdata_valid3 = 1'd0;
reg builder_new_master_rdata_valid4 = 1'd0;
reg builder_new_master_rdata_valid5 = 1'd0;
reg builder_new_master_rdata_valid6 = 1'd0;
reg builder_new_master_rdata_valid7 = 1'd0;
reg builder_new_master_rdata_valid8 = 1'd0;
reg builder_new_master_rdata_valid9 = 1'd0;
reg [1:0] builder_fullmemorywe_state = 2'd0;
reg [1:0] builder_fullmemorywe_next_state = 2'd0;
reg [1:0] builder_litedramwishbone2native_state = 2'd0;
reg [1:0] builder_litedramwishbone2native_next_state = 2'd0;
reg main_count_next_value = 1'd0;
reg main_count_next_value_ce = 1'd0;
wire builder_wb_sdram_con_request;
wire builder_wb_sdram_con_grant;
wire [29:0] builder_basesoc_shared_adr;
wire [31:0] builder_basesoc_shared_dat_w;
reg [31:0] builder_basesoc_shared_dat_r = 32'd0;
wire [3:0] builder_basesoc_shared_sel;
wire builder_basesoc_shared_cyc;
wire builder_basesoc_shared_stb;
reg builder_basesoc_shared_ack = 1'd0;
wire builder_basesoc_shared_we;
wire [2:0] builder_basesoc_shared_cti;
wire [1:0] builder_basesoc_shared_bte;
wire builder_basesoc_shared_err;
wire builder_basesoc_request;
wire builder_basesoc_grant;
reg [2:0] builder_basesoc_slave_sel = 3'd0;
reg [2:0] builder_basesoc_slave_sel_r = 3'd0;
reg builder_basesoc_error = 1'd0;
wire builder_basesoc_wait;
wire builder_basesoc_done;
reg [19:0] builder_basesoc_count = 20'd1000000;
wire [13:0] builder_basesoc_csrbankarray_interface0_bank_bus_adr;
wire builder_basesoc_csrbankarray_interface0_bank_bus_we;
wire [7:0] builder_basesoc_csrbankarray_interface0_bank_bus_dat_w;
reg [7:0] builder_basesoc_csrbankarray_interface0_bank_bus_dat_r = 8'd0;
wire builder_basesoc_csrbankarray_csrbank0_reset0_re;
wire builder_basesoc_csrbankarray_csrbank0_reset0_r;
wire builder_basesoc_csrbankarray_csrbank0_reset0_we;
wire builder_basesoc_csrbankarray_csrbank0_reset0_w;
wire builder_basesoc_csrbankarray_csrbank0_scratch3_re;
wire [7:0] builder_basesoc_csrbankarray_csrbank0_scratch3_r;
wire builder_basesoc_csrbankarray_csrbank0_scratch3_we;
wire [7:0] builder_basesoc_csrbankarray_csrbank0_scratch3_w;
wire builder_basesoc_csrbankarray_csrbank0_scratch2_re;
wire [7:0] builder_basesoc_csrbankarray_csrbank0_scratch2_r;
wire builder_basesoc_csrbankarray_csrbank0_scratch2_we;
wire [7:0] builder_basesoc_csrbankarray_csrbank0_scratch2_w;
wire builder_basesoc_csrbankarray_csrbank0_scratch1_re;
wire [7:0] builder_basesoc_csrbankarray_csrbank0_scratch1_r;
wire builder_basesoc_csrbankarray_csrbank0_scratch1_we;
wire [7:0] builder_basesoc_csrbankarray_csrbank0_scratch1_w;
wire builder_basesoc_csrbankarray_csrbank0_scratch0_re;
wire [7:0] builder_basesoc_csrbankarray_csrbank0_scratch0_r;
wire builder_basesoc_csrbankarray_csrbank0_scratch0_we;
wire [7:0] builder_basesoc_csrbankarray_csrbank0_scratch0_w;
wire builder_basesoc_csrbankarray_csrbank0_bus_errors3_re;
wire [7:0] builder_basesoc_csrbankarray_csrbank0_bus_errors3_r;
wire builder_basesoc_csrbankarray_csrbank0_bus_errors3_we;
wire [7:0] builder_basesoc_csrbankarray_csrbank0_bus_errors3_w;
wire builder_basesoc_csrbankarray_csrbank0_bus_errors2_re;
wire [7:0] builder_basesoc_csrbankarray_csrbank0_bus_errors2_r;
wire builder_basesoc_csrbankarray_csrbank0_bus_errors2_we;
wire [7:0] builder_basesoc_csrbankarray_csrbank0_bus_errors2_w;
wire builder_basesoc_csrbankarray_csrbank0_bus_errors1_re;
wire [7:0] builder_basesoc_csrbankarray_csrbank0_bus_errors1_r;
wire builder_basesoc_csrbankarray_csrbank0_bus_errors1_we;
wire [7:0] builder_basesoc_csrbankarray_csrbank0_bus_errors1_w;
wire builder_basesoc_csrbankarray_csrbank0_bus_errors0_re;
wire [7:0] builder_basesoc_csrbankarray_csrbank0_bus_errors0_r;
wire builder_basesoc_csrbankarray_csrbank0_bus_errors0_we;
wire [7:0] builder_basesoc_csrbankarray_csrbank0_bus_errors0_w;
wire builder_basesoc_csrbankarray_csrbank0_sel;
wire [13:0] builder_basesoc_csrbankarray_interface1_bank_bus_adr;
wire builder_basesoc_csrbankarray_interface1_bank_bus_we;
wire [7:0] builder_basesoc_csrbankarray_interface1_bank_bus_dat_w;
reg [7:0] builder_basesoc_csrbankarray_interface1_bank_bus_dat_r = 8'd0;
wire builder_basesoc_csrbankarray_csrbank1_half_sys8x_taps0_re;
wire [4:0] builder_basesoc_csrbankarray_csrbank1_half_sys8x_taps0_r;
wire builder_basesoc_csrbankarray_csrbank1_half_sys8x_taps0_we;
wire [4:0] builder_basesoc_csrbankarray_csrbank1_half_sys8x_taps0_w;
wire builder_basesoc_csrbankarray_csrbank1_dly_sel0_re;
wire [1:0] builder_basesoc_csrbankarray_csrbank1_dly_sel0_r;
wire builder_basesoc_csrbankarray_csrbank1_dly_sel0_we;
wire [1:0] builder_basesoc_csrbankarray_csrbank1_dly_sel0_w;
wire builder_basesoc_csrbankarray_csrbank1_sel;
wire [13:0] builder_basesoc_csrbankarray_sram_bus_adr;
wire builder_basesoc_csrbankarray_sram_bus_we;
wire [7:0] builder_basesoc_csrbankarray_sram_bus_dat_w;
reg [7:0] builder_basesoc_csrbankarray_sram_bus_dat_r = 8'd0;
wire [6:0] builder_basesoc_csrbankarray_adr;
wire [7:0] builder_basesoc_csrbankarray_dat_r;
wire builder_basesoc_csrbankarray_sel;
reg builder_basesoc_csrbankarray_sel_r = 1'd0;
wire [13:0] builder_basesoc_csrbankarray_interface2_bank_bus_adr;
wire builder_basesoc_csrbankarray_interface2_bank_bus_we;
wire [7:0] builder_basesoc_csrbankarray_interface2_bank_bus_dat_w;
reg [7:0] builder_basesoc_csrbankarray_interface2_bank_bus_dat_r = 8'd0;
wire builder_basesoc_csrbankarray_csrbank2_dfii_control0_re;
wire [3:0] builder_basesoc_csrbankarray_csrbank2_dfii_control0_r;
wire builder_basesoc_csrbankarray_csrbank2_dfii_control0_we;
wire [3:0] builder_basesoc_csrbankarray_csrbank2_dfii_control0_w;
wire builder_basesoc_csrbankarray_csrbank2_dfii_pi0_command0_re;
wire [5:0] builder_basesoc_csrbankarray_csrbank2_dfii_pi0_command0_r;
wire builder_basesoc_csrbankarray_csrbank2_dfii_pi0_command0_we;
wire [5:0] builder_basesoc_csrbankarray_csrbank2_dfii_pi0_command0_w;
wire builder_basesoc_csrbankarray_csrbank2_dfii_pi0_address1_re;
wire [5:0] builder_basesoc_csrbankarray_csrbank2_dfii_pi0_address1_r;
wire builder_basesoc_csrbankarray_csrbank2_dfii_pi0_address1_we;
wire [5:0] builder_basesoc_csrbankarray_csrbank2_dfii_pi0_address1_w;
wire builder_basesoc_csrbankarray_csrbank2_dfii_pi0_address0_re;
wire [7:0] builder_basesoc_csrbankarray_csrbank2_dfii_pi0_address0_r;
wire builder_basesoc_csrbankarray_csrbank2_dfii_pi0_address0_we;
wire [7:0] builder_basesoc_csrbankarray_csrbank2_dfii_pi0_address0_w;
wire builder_basesoc_csrbankarray_csrbank2_dfii_pi0_baddress0_re;
wire [2:0] builder_basesoc_csrbankarray_csrbank2_dfii_pi0_baddress0_r;
wire builder_basesoc_csrbankarray_csrbank2_dfii_pi0_baddress0_we;
wire [2:0] builder_basesoc_csrbankarray_csrbank2_dfii_pi0_baddress0_w;
wire builder_basesoc_csrbankarray_csrbank2_dfii_pi0_wrdata3_re;
wire [7:0] builder_basesoc_csrbankarray_csrbank2_dfii_pi0_wrdata3_r;
wire builder_basesoc_csrbankarray_csrbank2_dfii_pi0_wrdata3_we;
wire [7:0] builder_basesoc_csrbankarray_csrbank2_dfii_pi0_wrdata3_w;
wire builder_basesoc_csrbankarray_csrbank2_dfii_pi0_wrdata2_re;
wire [7:0] builder_basesoc_csrbankarray_csrbank2_dfii_pi0_wrdata2_r;
wire builder_basesoc_csrbankarray_csrbank2_dfii_pi0_wrdata2_we;
wire [7:0] builder_basesoc_csrbankarray_csrbank2_dfii_pi0_wrdata2_w;
wire builder_basesoc_csrbankarray_csrbank2_dfii_pi0_wrdata1_re;
wire [7:0] builder_basesoc_csrbankarray_csrbank2_dfii_pi0_wrdata1_r;
wire builder_basesoc_csrbankarray_csrbank2_dfii_pi0_wrdata1_we;
wire [7:0] builder_basesoc_csrbankarray_csrbank2_dfii_pi0_wrdata1_w;
wire builder_basesoc_csrbankarray_csrbank2_dfii_pi0_wrdata0_re;
wire [7:0] builder_basesoc_csrbankarray_csrbank2_dfii_pi0_wrdata0_r;
wire builder_basesoc_csrbankarray_csrbank2_dfii_pi0_wrdata0_we;
wire [7:0] builder_basesoc_csrbankarray_csrbank2_dfii_pi0_wrdata0_w;
wire builder_basesoc_csrbankarray_csrbank2_dfii_pi0_rddata3_re;
wire [7:0] builder_basesoc_csrbankarray_csrbank2_dfii_pi0_rddata3_r;
wire builder_basesoc_csrbankarray_csrbank2_dfii_pi0_rddata3_we;
wire [7:0] builder_basesoc_csrbankarray_csrbank2_dfii_pi0_rddata3_w;
wire builder_basesoc_csrbankarray_csrbank2_dfii_pi0_rddata2_re;
wire [7:0] builder_basesoc_csrbankarray_csrbank2_dfii_pi0_rddata2_r;
wire builder_basesoc_csrbankarray_csrbank2_dfii_pi0_rddata2_we;
wire [7:0] builder_basesoc_csrbankarray_csrbank2_dfii_pi0_rddata2_w;
wire builder_basesoc_csrbankarray_csrbank2_dfii_pi0_rddata1_re;
wire [7:0] builder_basesoc_csrbankarray_csrbank2_dfii_pi0_rddata1_r;
wire builder_basesoc_csrbankarray_csrbank2_dfii_pi0_rddata1_we;
wire [7:0] builder_basesoc_csrbankarray_csrbank2_dfii_pi0_rddata1_w;
wire builder_basesoc_csrbankarray_csrbank2_dfii_pi0_rddata0_re;
wire [7:0] builder_basesoc_csrbankarray_csrbank2_dfii_pi0_rddata0_r;
wire builder_basesoc_csrbankarray_csrbank2_dfii_pi0_rddata0_we;
wire [7:0] builder_basesoc_csrbankarray_csrbank2_dfii_pi0_rddata0_w;
wire builder_basesoc_csrbankarray_csrbank2_dfii_pi1_command0_re;
wire [5:0] builder_basesoc_csrbankarray_csrbank2_dfii_pi1_command0_r;
wire builder_basesoc_csrbankarray_csrbank2_dfii_pi1_command0_we;
wire [5:0] builder_basesoc_csrbankarray_csrbank2_dfii_pi1_command0_w;
wire builder_basesoc_csrbankarray_csrbank2_dfii_pi1_address1_re;
wire [5:0] builder_basesoc_csrbankarray_csrbank2_dfii_pi1_address1_r;
wire builder_basesoc_csrbankarray_csrbank2_dfii_pi1_address1_we;
wire [5:0] builder_basesoc_csrbankarray_csrbank2_dfii_pi1_address1_w;
wire builder_basesoc_csrbankarray_csrbank2_dfii_pi1_address0_re;
wire [7:0] builder_basesoc_csrbankarray_csrbank2_dfii_pi1_address0_r;
wire builder_basesoc_csrbankarray_csrbank2_dfii_pi1_address0_we;
wire [7:0] builder_basesoc_csrbankarray_csrbank2_dfii_pi1_address0_w;
wire builder_basesoc_csrbankarray_csrbank2_dfii_pi1_baddress0_re;
wire [2:0] builder_basesoc_csrbankarray_csrbank2_dfii_pi1_baddress0_r;
wire builder_basesoc_csrbankarray_csrbank2_dfii_pi1_baddress0_we;
wire [2:0] builder_basesoc_csrbankarray_csrbank2_dfii_pi1_baddress0_w;
wire builder_basesoc_csrbankarray_csrbank2_dfii_pi1_wrdata3_re;
wire [7:0] builder_basesoc_csrbankarray_csrbank2_dfii_pi1_wrdata3_r;
wire builder_basesoc_csrbankarray_csrbank2_dfii_pi1_wrdata3_we;
wire [7:0] builder_basesoc_csrbankarray_csrbank2_dfii_pi1_wrdata3_w;
wire builder_basesoc_csrbankarray_csrbank2_dfii_pi1_wrdata2_re;
wire [7:0] builder_basesoc_csrbankarray_csrbank2_dfii_pi1_wrdata2_r;
wire builder_basesoc_csrbankarray_csrbank2_dfii_pi1_wrdata2_we;
wire [7:0] builder_basesoc_csrbankarray_csrbank2_dfii_pi1_wrdata2_w;
wire builder_basesoc_csrbankarray_csrbank2_dfii_pi1_wrdata1_re;
wire [7:0] builder_basesoc_csrbankarray_csrbank2_dfii_pi1_wrdata1_r;
wire builder_basesoc_csrbankarray_csrbank2_dfii_pi1_wrdata1_we;
wire [7:0] builder_basesoc_csrbankarray_csrbank2_dfii_pi1_wrdata1_w;
wire builder_basesoc_csrbankarray_csrbank2_dfii_pi1_wrdata0_re;
wire [7:0] builder_basesoc_csrbankarray_csrbank2_dfii_pi1_wrdata0_r;
wire builder_basesoc_csrbankarray_csrbank2_dfii_pi1_wrdata0_we;
wire [7:0] builder_basesoc_csrbankarray_csrbank2_dfii_pi1_wrdata0_w;
wire builder_basesoc_csrbankarray_csrbank2_dfii_pi1_rddata3_re;
wire [7:0] builder_basesoc_csrbankarray_csrbank2_dfii_pi1_rddata3_r;
wire builder_basesoc_csrbankarray_csrbank2_dfii_pi1_rddata3_we;
wire [7:0] builder_basesoc_csrbankarray_csrbank2_dfii_pi1_rddata3_w;
wire builder_basesoc_csrbankarray_csrbank2_dfii_pi1_rddata2_re;
wire [7:0] builder_basesoc_csrbankarray_csrbank2_dfii_pi1_rddata2_r;
wire builder_basesoc_csrbankarray_csrbank2_dfii_pi1_rddata2_we;
wire [7:0] builder_basesoc_csrbankarray_csrbank2_dfii_pi1_rddata2_w;
wire builder_basesoc_csrbankarray_csrbank2_dfii_pi1_rddata1_re;
wire [7:0] builder_basesoc_csrbankarray_csrbank2_dfii_pi1_rddata1_r;
wire builder_basesoc_csrbankarray_csrbank2_dfii_pi1_rddata1_we;
wire [7:0] builder_basesoc_csrbankarray_csrbank2_dfii_pi1_rddata1_w;
wire builder_basesoc_csrbankarray_csrbank2_dfii_pi1_rddata0_re;
wire [7:0] builder_basesoc_csrbankarray_csrbank2_dfii_pi1_rddata0_r;
wire builder_basesoc_csrbankarray_csrbank2_dfii_pi1_rddata0_we;
wire [7:0] builder_basesoc_csrbankarray_csrbank2_dfii_pi1_rddata0_w;
wire builder_basesoc_csrbankarray_csrbank2_dfii_pi2_command0_re;
wire [5:0] builder_basesoc_csrbankarray_csrbank2_dfii_pi2_command0_r;
wire builder_basesoc_csrbankarray_csrbank2_dfii_pi2_command0_we;
wire [5:0] builder_basesoc_csrbankarray_csrbank2_dfii_pi2_command0_w;
wire builder_basesoc_csrbankarray_csrbank2_dfii_pi2_address1_re;
wire [5:0] builder_basesoc_csrbankarray_csrbank2_dfii_pi2_address1_r;
wire builder_basesoc_csrbankarray_csrbank2_dfii_pi2_address1_we;
wire [5:0] builder_basesoc_csrbankarray_csrbank2_dfii_pi2_address1_w;
wire builder_basesoc_csrbankarray_csrbank2_dfii_pi2_address0_re;
wire [7:0] builder_basesoc_csrbankarray_csrbank2_dfii_pi2_address0_r;
wire builder_basesoc_csrbankarray_csrbank2_dfii_pi2_address0_we;
wire [7:0] builder_basesoc_csrbankarray_csrbank2_dfii_pi2_address0_w;
wire builder_basesoc_csrbankarray_csrbank2_dfii_pi2_baddress0_re;
wire [2:0] builder_basesoc_csrbankarray_csrbank2_dfii_pi2_baddress0_r;
wire builder_basesoc_csrbankarray_csrbank2_dfii_pi2_baddress0_we;
wire [2:0] builder_basesoc_csrbankarray_csrbank2_dfii_pi2_baddress0_w;
wire builder_basesoc_csrbankarray_csrbank2_dfii_pi2_wrdata3_re;
wire [7:0] builder_basesoc_csrbankarray_csrbank2_dfii_pi2_wrdata3_r;
wire builder_basesoc_csrbankarray_csrbank2_dfii_pi2_wrdata3_we;
wire [7:0] builder_basesoc_csrbankarray_csrbank2_dfii_pi2_wrdata3_w;
wire builder_basesoc_csrbankarray_csrbank2_dfii_pi2_wrdata2_re;
wire [7:0] builder_basesoc_csrbankarray_csrbank2_dfii_pi2_wrdata2_r;
wire builder_basesoc_csrbankarray_csrbank2_dfii_pi2_wrdata2_we;
wire [7:0] builder_basesoc_csrbankarray_csrbank2_dfii_pi2_wrdata2_w;
wire builder_basesoc_csrbankarray_csrbank2_dfii_pi2_wrdata1_re;
wire [7:0] builder_basesoc_csrbankarray_csrbank2_dfii_pi2_wrdata1_r;
wire builder_basesoc_csrbankarray_csrbank2_dfii_pi2_wrdata1_we;
wire [7:0] builder_basesoc_csrbankarray_csrbank2_dfii_pi2_wrdata1_w;
wire builder_basesoc_csrbankarray_csrbank2_dfii_pi2_wrdata0_re;
wire [7:0] builder_basesoc_csrbankarray_csrbank2_dfii_pi2_wrdata0_r;
wire builder_basesoc_csrbankarray_csrbank2_dfii_pi2_wrdata0_we;
wire [7:0] builder_basesoc_csrbankarray_csrbank2_dfii_pi2_wrdata0_w;
wire builder_basesoc_csrbankarray_csrbank2_dfii_pi2_rddata3_re;
wire [7:0] builder_basesoc_csrbankarray_csrbank2_dfii_pi2_rddata3_r;
wire builder_basesoc_csrbankarray_csrbank2_dfii_pi2_rddata3_we;
wire [7:0] builder_basesoc_csrbankarray_csrbank2_dfii_pi2_rddata3_w;
wire builder_basesoc_csrbankarray_csrbank2_dfii_pi2_rddata2_re;
wire [7:0] builder_basesoc_csrbankarray_csrbank2_dfii_pi2_rddata2_r;
wire builder_basesoc_csrbankarray_csrbank2_dfii_pi2_rddata2_we;
wire [7:0] builder_basesoc_csrbankarray_csrbank2_dfii_pi2_rddata2_w;
wire builder_basesoc_csrbankarray_csrbank2_dfii_pi2_rddata1_re;
wire [7:0] builder_basesoc_csrbankarray_csrbank2_dfii_pi2_rddata1_r;
wire builder_basesoc_csrbankarray_csrbank2_dfii_pi2_rddata1_we;
wire [7:0] builder_basesoc_csrbankarray_csrbank2_dfii_pi2_rddata1_w;
wire builder_basesoc_csrbankarray_csrbank2_dfii_pi2_rddata0_re;
wire [7:0] builder_basesoc_csrbankarray_csrbank2_dfii_pi2_rddata0_r;
wire builder_basesoc_csrbankarray_csrbank2_dfii_pi2_rddata0_we;
wire [7:0] builder_basesoc_csrbankarray_csrbank2_dfii_pi2_rddata0_w;
wire builder_basesoc_csrbankarray_csrbank2_dfii_pi3_command0_re;
wire [5:0] builder_basesoc_csrbankarray_csrbank2_dfii_pi3_command0_r;
wire builder_basesoc_csrbankarray_csrbank2_dfii_pi3_command0_we;
wire [5:0] builder_basesoc_csrbankarray_csrbank2_dfii_pi3_command0_w;
wire builder_basesoc_csrbankarray_csrbank2_dfii_pi3_address1_re;
wire [5:0] builder_basesoc_csrbankarray_csrbank2_dfii_pi3_address1_r;
wire builder_basesoc_csrbankarray_csrbank2_dfii_pi3_address1_we;
wire [5:0] builder_basesoc_csrbankarray_csrbank2_dfii_pi3_address1_w;
wire builder_basesoc_csrbankarray_csrbank2_dfii_pi3_address0_re;
wire [7:0] builder_basesoc_csrbankarray_csrbank2_dfii_pi3_address0_r;
wire builder_basesoc_csrbankarray_csrbank2_dfii_pi3_address0_we;
wire [7:0] builder_basesoc_csrbankarray_csrbank2_dfii_pi3_address0_w;
wire builder_basesoc_csrbankarray_csrbank2_dfii_pi3_baddress0_re;
wire [2:0] builder_basesoc_csrbankarray_csrbank2_dfii_pi3_baddress0_r;
wire builder_basesoc_csrbankarray_csrbank2_dfii_pi3_baddress0_we;
wire [2:0] builder_basesoc_csrbankarray_csrbank2_dfii_pi3_baddress0_w;
wire builder_basesoc_csrbankarray_csrbank2_dfii_pi3_wrdata3_re;
wire [7:0] builder_basesoc_csrbankarray_csrbank2_dfii_pi3_wrdata3_r;
wire builder_basesoc_csrbankarray_csrbank2_dfii_pi3_wrdata3_we;
wire [7:0] builder_basesoc_csrbankarray_csrbank2_dfii_pi3_wrdata3_w;
wire builder_basesoc_csrbankarray_csrbank2_dfii_pi3_wrdata2_re;
wire [7:0] builder_basesoc_csrbankarray_csrbank2_dfii_pi3_wrdata2_r;
wire builder_basesoc_csrbankarray_csrbank2_dfii_pi3_wrdata2_we;
wire [7:0] builder_basesoc_csrbankarray_csrbank2_dfii_pi3_wrdata2_w;
wire builder_basesoc_csrbankarray_csrbank2_dfii_pi3_wrdata1_re;
wire [7:0] builder_basesoc_csrbankarray_csrbank2_dfii_pi3_wrdata1_r;
wire builder_basesoc_csrbankarray_csrbank2_dfii_pi3_wrdata1_we;
wire [7:0] builder_basesoc_csrbankarray_csrbank2_dfii_pi3_wrdata1_w;
wire builder_basesoc_csrbankarray_csrbank2_dfii_pi3_wrdata0_re;
wire [7:0] builder_basesoc_csrbankarray_csrbank2_dfii_pi3_wrdata0_r;
wire builder_basesoc_csrbankarray_csrbank2_dfii_pi3_wrdata0_we;
wire [7:0] builder_basesoc_csrbankarray_csrbank2_dfii_pi3_wrdata0_w;
wire builder_basesoc_csrbankarray_csrbank2_dfii_pi3_rddata3_re;
wire [7:0] builder_basesoc_csrbankarray_csrbank2_dfii_pi3_rddata3_r;
wire builder_basesoc_csrbankarray_csrbank2_dfii_pi3_rddata3_we;
wire [7:0] builder_basesoc_csrbankarray_csrbank2_dfii_pi3_rddata3_w;
wire builder_basesoc_csrbankarray_csrbank2_dfii_pi3_rddata2_re;
wire [7:0] builder_basesoc_csrbankarray_csrbank2_dfii_pi3_rddata2_r;
wire builder_basesoc_csrbankarray_csrbank2_dfii_pi3_rddata2_we;
wire [7:0] builder_basesoc_csrbankarray_csrbank2_dfii_pi3_rddata2_w;
wire builder_basesoc_csrbankarray_csrbank2_dfii_pi3_rddata1_re;
wire [7:0] builder_basesoc_csrbankarray_csrbank2_dfii_pi3_rddata1_r;
wire builder_basesoc_csrbankarray_csrbank2_dfii_pi3_rddata1_we;
wire [7:0] builder_basesoc_csrbankarray_csrbank2_dfii_pi3_rddata1_w;
wire builder_basesoc_csrbankarray_csrbank2_dfii_pi3_rddata0_re;
wire [7:0] builder_basesoc_csrbankarray_csrbank2_dfii_pi3_rddata0_r;
wire builder_basesoc_csrbankarray_csrbank2_dfii_pi3_rddata0_we;
wire [7:0] builder_basesoc_csrbankarray_csrbank2_dfii_pi3_rddata0_w;
wire builder_basesoc_csrbankarray_csrbank2_sel;
wire [13:0] builder_basesoc_csrbankarray_interface3_bank_bus_adr;
wire builder_basesoc_csrbankarray_interface3_bank_bus_we;
wire [7:0] builder_basesoc_csrbankarray_interface3_bank_bus_dat_w;
reg [7:0] builder_basesoc_csrbankarray_interface3_bank_bus_dat_r = 8'd0;
wire builder_basesoc_csrbankarray_csrbank3_load3_re;
wire [7:0] builder_basesoc_csrbankarray_csrbank3_load3_r;
wire builder_basesoc_csrbankarray_csrbank3_load3_we;
wire [7:0] builder_basesoc_csrbankarray_csrbank3_load3_w;
wire builder_basesoc_csrbankarray_csrbank3_load2_re;
wire [7:0] builder_basesoc_csrbankarray_csrbank3_load2_r;
wire builder_basesoc_csrbankarray_csrbank3_load2_we;
wire [7:0] builder_basesoc_csrbankarray_csrbank3_load2_w;
wire builder_basesoc_csrbankarray_csrbank3_load1_re;
wire [7:0] builder_basesoc_csrbankarray_csrbank3_load1_r;
wire builder_basesoc_csrbankarray_csrbank3_load1_we;
wire [7:0] builder_basesoc_csrbankarray_csrbank3_load1_w;
wire builder_basesoc_csrbankarray_csrbank3_load0_re;
wire [7:0] builder_basesoc_csrbankarray_csrbank3_load0_r;
wire builder_basesoc_csrbankarray_csrbank3_load0_we;
wire [7:0] builder_basesoc_csrbankarray_csrbank3_load0_w;
wire builder_basesoc_csrbankarray_csrbank3_reload3_re;
wire [7:0] builder_basesoc_csrbankarray_csrbank3_reload3_r;
wire builder_basesoc_csrbankarray_csrbank3_reload3_we;
wire [7:0] builder_basesoc_csrbankarray_csrbank3_reload3_w;
wire builder_basesoc_csrbankarray_csrbank3_reload2_re;
wire [7:0] builder_basesoc_csrbankarray_csrbank3_reload2_r;
wire builder_basesoc_csrbankarray_csrbank3_reload2_we;
wire [7:0] builder_basesoc_csrbankarray_csrbank3_reload2_w;
wire builder_basesoc_csrbankarray_csrbank3_reload1_re;
wire [7:0] builder_basesoc_csrbankarray_csrbank3_reload1_r;
wire builder_basesoc_csrbankarray_csrbank3_reload1_we;
wire [7:0] builder_basesoc_csrbankarray_csrbank3_reload1_w;
wire builder_basesoc_csrbankarray_csrbank3_reload0_re;
wire [7:0] builder_basesoc_csrbankarray_csrbank3_reload0_r;
wire builder_basesoc_csrbankarray_csrbank3_reload0_we;
wire [7:0] builder_basesoc_csrbankarray_csrbank3_reload0_w;
wire builder_basesoc_csrbankarray_csrbank3_en0_re;
wire builder_basesoc_csrbankarray_csrbank3_en0_r;
wire builder_basesoc_csrbankarray_csrbank3_en0_we;
wire builder_basesoc_csrbankarray_csrbank3_en0_w;
wire builder_basesoc_csrbankarray_csrbank3_update_value0_re;
wire builder_basesoc_csrbankarray_csrbank3_update_value0_r;
wire builder_basesoc_csrbankarray_csrbank3_update_value0_we;
wire builder_basesoc_csrbankarray_csrbank3_update_value0_w;
wire builder_basesoc_csrbankarray_csrbank3_value3_re;
wire [7:0] builder_basesoc_csrbankarray_csrbank3_value3_r;
wire builder_basesoc_csrbankarray_csrbank3_value3_we;
wire [7:0] builder_basesoc_csrbankarray_csrbank3_value3_w;
wire builder_basesoc_csrbankarray_csrbank3_value2_re;
wire [7:0] builder_basesoc_csrbankarray_csrbank3_value2_r;
wire builder_basesoc_csrbankarray_csrbank3_value2_we;
wire [7:0] builder_basesoc_csrbankarray_csrbank3_value2_w;
wire builder_basesoc_csrbankarray_csrbank3_value1_re;
wire [7:0] builder_basesoc_csrbankarray_csrbank3_value1_r;
wire builder_basesoc_csrbankarray_csrbank3_value1_we;
wire [7:0] builder_basesoc_csrbankarray_csrbank3_value1_w;
wire builder_basesoc_csrbankarray_csrbank3_value0_re;
wire [7:0] builder_basesoc_csrbankarray_csrbank3_value0_r;
wire builder_basesoc_csrbankarray_csrbank3_value0_we;
wire [7:0] builder_basesoc_csrbankarray_csrbank3_value0_w;
wire builder_basesoc_csrbankarray_csrbank3_ev_enable0_re;
wire builder_basesoc_csrbankarray_csrbank3_ev_enable0_r;
wire builder_basesoc_csrbankarray_csrbank3_ev_enable0_we;
wire builder_basesoc_csrbankarray_csrbank3_ev_enable0_w;
wire builder_basesoc_csrbankarray_csrbank3_sel;
wire [13:0] builder_basesoc_csrcon_adr;
wire builder_basesoc_csrcon_we;
wire [7:0] builder_basesoc_csrcon_dat_w;
wire [7:0] builder_basesoc_csrcon_dat_r;
reg builder_rhs_array_muxed0 = 1'd0;
reg [13:0] builder_rhs_array_muxed1 = 14'd0;
reg [2:0] builder_rhs_array_muxed2 = 3'd0;
reg builder_rhs_array_muxed3 = 1'd0;
reg builder_rhs_array_muxed4 = 1'd0;
reg builder_rhs_array_muxed5 = 1'd0;
reg builder_t_array_muxed0 = 1'd0;
reg builder_t_array_muxed1 = 1'd0;
reg builder_t_array_muxed2 = 1'd0;
reg builder_rhs_array_muxed6 = 1'd0;
reg [13:0] builder_rhs_array_muxed7 = 14'd0;
reg [2:0] builder_rhs_array_muxed8 = 3'd0;
reg builder_rhs_array_muxed9 = 1'd0;
reg builder_rhs_array_muxed10 = 1'd0;
reg builder_rhs_array_muxed11 = 1'd0;
reg builder_t_array_muxed3 = 1'd0;
reg builder_t_array_muxed4 = 1'd0;
reg builder_t_array_muxed5 = 1'd0;
reg [20:0] builder_rhs_array_muxed12 = 21'd0;
reg builder_rhs_array_muxed13 = 1'd0;
reg builder_rhs_array_muxed14 = 1'd0;
reg [20:0] builder_rhs_array_muxed15 = 21'd0;
reg builder_rhs_array_muxed16 = 1'd0;
reg builder_rhs_array_muxed17 = 1'd0;
reg [20:0] builder_rhs_array_muxed18 = 21'd0;
reg builder_rhs_array_muxed19 = 1'd0;
reg builder_rhs_array_muxed20 = 1'd0;
reg [20:0] builder_rhs_array_muxed21 = 21'd0;
reg builder_rhs_array_muxed22 = 1'd0;
reg builder_rhs_array_muxed23 = 1'd0;
reg [20:0] builder_rhs_array_muxed24 = 21'd0;
reg builder_rhs_array_muxed25 = 1'd0;
reg builder_rhs_array_muxed26 = 1'd0;
reg [20:0] builder_rhs_array_muxed27 = 21'd0;
reg builder_rhs_array_muxed28 = 1'd0;
reg builder_rhs_array_muxed29 = 1'd0;
reg [20:0] builder_rhs_array_muxed30 = 21'd0;
reg builder_rhs_array_muxed31 = 1'd0;
reg builder_rhs_array_muxed32 = 1'd0;
reg [20:0] builder_rhs_array_muxed33 = 21'd0;
reg builder_rhs_array_muxed34 = 1'd0;
reg builder_rhs_array_muxed35 = 1'd0;
reg [29:0] builder_rhs_array_muxed36 = 30'd0;
reg [31:0] builder_rhs_array_muxed37 = 32'd0;
reg [3:0] builder_rhs_array_muxed38 = 4'd0;
reg builder_rhs_array_muxed39 = 1'd0;
reg builder_rhs_array_muxed40 = 1'd0;
reg builder_rhs_array_muxed41 = 1'd0;
reg [2:0] builder_rhs_array_muxed42 = 3'd0;
reg [1:0] builder_rhs_array_muxed43 = 2'd0;
reg [29:0] builder_rhs_array_muxed44 = 30'd0;
reg [31:0] builder_rhs_array_muxed45 = 32'd0;
reg [3:0] builder_rhs_array_muxed46 = 4'd0;
reg builder_rhs_array_muxed47 = 1'd0;
reg builder_rhs_array_muxed48 = 1'd0;
reg builder_rhs_array_muxed49 = 1'd0;
reg [2:0] builder_rhs_array_muxed50 = 3'd0;
reg [1:0] builder_rhs_array_muxed51 = 2'd0;
reg [2:0] builder_array_muxed0 = 3'd0;
reg [13:0] builder_array_muxed1 = 14'd0;
reg builder_array_muxed2 = 1'd0;
reg builder_array_muxed3 = 1'd0;
reg builder_array_muxed4 = 1'd0;
reg builder_array_muxed5 = 1'd0;
reg builder_array_muxed6 = 1'd0;
reg [2:0] builder_array_muxed7 = 3'd0;
reg [13:0] builder_array_muxed8 = 14'd0;
reg builder_array_muxed9 = 1'd0;
reg builder_array_muxed10 = 1'd0;
reg builder_array_muxed11 = 1'd0;
reg builder_array_muxed12 = 1'd0;
reg builder_array_muxed13 = 1'd0;
reg [2:0] builder_array_muxed14 = 3'd0;
reg [13:0] builder_array_muxed15 = 14'd0;
reg builder_array_muxed16 = 1'd0;
reg builder_array_muxed17 = 1'd0;
reg builder_array_muxed18 = 1'd0;
reg builder_array_muxed19 = 1'd0;
reg builder_array_muxed20 = 1'd0;
reg [2:0] builder_array_muxed21 = 3'd0;
reg [13:0] builder_array_muxed22 = 14'd0;
reg builder_array_muxed23 = 1'd0;
reg builder_array_muxed24 = 1'd0;
reg builder_array_muxed25 = 1'd0;
reg builder_array_muxed26 = 1'd0;
reg builder_array_muxed27 = 1'd0;
(* async_reg = "true", mr_ff = "true", dont_touch = "true" *) reg builder_regs0 = 1'd0;
(* async_reg = "true", dont_touch = "true" *) reg builder_regs1 = 1'd0;
wire builder_xilinxasyncresetsynchronizerimpl0;
wire builder_xilinxasyncresetsynchronizerimpl0_rst_meta;
wire builder_xilinxasyncresetsynchronizerimpl1;
wire builder_xilinxasyncresetsynchronizerimpl1_rst_meta;
wire builder_xilinxasyncresetsynchronizerimpl1_expr;
wire builder_xilinxasyncresetsynchronizerimpl2;
wire builder_xilinxasyncresetsynchronizerimpl2_rst_meta;
wire builder_xilinxasyncresetsynchronizerimpl2_expr;
wire builder_xilinxasyncresetsynchronizerimpl3;
wire builder_xilinxasyncresetsynchronizerimpl3_rst_meta;
assign main_ctrl_bus_error = builder_basesoc_error;
assign main_ctrl_reset = main_ctrl_reset_re;
assign main_ctrl_bus_errors_status = main_ctrl_bus_errors;
always @(*) begin
	main_sram_we <= 4'd0;
	main_sram_we[0] <= (((main_sram_bus_cyc & main_sram_bus_stb) & main_sram_bus_we) & main_sram_bus_sel[0]);
	main_sram_we[1] <= (((main_sram_bus_cyc & main_sram_bus_stb) & main_sram_bus_we) & main_sram_bus_sel[1]);
	main_sram_we[2] <= (((main_sram_bus_cyc & main_sram_bus_stb) & main_sram_bus_we) & main_sram_bus_sel[2]);
	main_sram_we[3] <= (((main_sram_bus_cyc & main_sram_bus_stb) & main_sram_bus_we) & main_sram_bus_sel[3]);
end
assign main_sram_adr = main_sram_bus_adr[9:0];
assign main_sram_bus_dat_r = main_sram_dat_r;
assign main_sram_dat_w = main_sram_bus_dat_w;
assign main_uart_reset = main_uart_done;
assign main_uart_source_ready = 1'd1;
assign main_uart_wishbone_adr = (main_uart_address + main_uart_word_counter);
assign main_uart_wishbone_dat_w = main_uart_data;
assign main_uart_wishbone_sel = 4'd15;
always @(*) begin
	main_uart_sink_payload_data <= 8'd0;
	case (main_uart_byte_counter)
		1'd0: begin
			main_uart_sink_payload_data <= main_uart_data[31:24];
		end
		1'd1: begin
			main_uart_sink_payload_data <= main_uart_data[23:16];
		end
		2'd2: begin
			main_uart_sink_payload_data <= main_uart_data[15:8];
		end
		default: begin
			main_uart_sink_payload_data <= main_uart_data[7:0];
		end
	endcase
end
assign main_uart_wait = (~main_uart_is_ongoing);
assign main_uart_sink_last = ((main_uart_byte_counter == 2'd3) & (main_uart_word_counter == (main_uart_length - 1'd1)));
always @(*) begin
	main_uart_word_counter_ce <= 1'd0;
	builder_uartwishbonebridge_next_state <= 3'd0;
	main_uart_wishbone_cyc <= 1'd0;
	main_uart_cmd_ce <= 1'd0;
	main_uart_wishbone_stb <= 1'd0;
	main_uart_length_ce <= 1'd0;
	main_uart_wishbone_we <= 1'd0;
	main_uart_address_ce <= 1'd0;
	main_uart_rx_data_ce <= 1'd0;
	main_uart_byte_counter_reset <= 1'd0;
	main_uart_tx_data_ce <= 1'd0;
	main_uart_byte_counter_ce <= 1'd0;
	main_uart_word_counter_reset <= 1'd0;
	main_uart_is_ongoing <= 1'd0;
	main_uart_sink_valid <= 1'd0;
	builder_uartwishbonebridge_next_state <= builder_uartwishbonebridge_state;
	case (builder_uartwishbonebridge_state)
		1'd1: begin
			if (main_uart_source_valid) begin
				main_uart_length_ce <= 1'd1;
				builder_uartwishbonebridge_next_state <= 2'd2;
			end
		end
		2'd2: begin
			if (main_uart_source_valid) begin
				main_uart_address_ce <= 1'd1;
				main_uart_byte_counter_ce <= 1'd1;
				if ((main_uart_byte_counter == 2'd3)) begin
					if ((main_uart_cmd == 1'd1)) begin
						builder_uartwishbonebridge_next_state <= 2'd3;
					end else begin
						if ((main_uart_cmd == 2'd2)) begin
							builder_uartwishbonebridge_next_state <= 3'd5;
						end
					end
					main_uart_byte_counter_reset <= 1'd1;
				end
			end
		end
		2'd3: begin
			if (main_uart_source_valid) begin
				main_uart_rx_data_ce <= 1'd1;
				main_uart_byte_counter_ce <= 1'd1;
				if ((main_uart_byte_counter == 2'd3)) begin
					builder_uartwishbonebridge_next_state <= 3'd4;
					main_uart_byte_counter_reset <= 1'd1;
				end
			end
		end
		3'd4: begin
			main_uart_wishbone_stb <= 1'd1;
			main_uart_wishbone_we <= 1'd1;
			main_uart_wishbone_cyc <= 1'd1;
			if (main_uart_wishbone_ack) begin
				main_uart_word_counter_ce <= 1'd1;
				if ((main_uart_word_counter == (main_uart_length - 1'd1))) begin
					builder_uartwishbonebridge_next_state <= 1'd0;
				end else begin
					builder_uartwishbonebridge_next_state <= 2'd3;
				end
			end
		end
		3'd5: begin
			main_uart_wishbone_stb <= 1'd1;
			main_uart_wishbone_we <= 1'd0;
			main_uart_wishbone_cyc <= 1'd1;
			if (main_uart_wishbone_ack) begin
				main_uart_tx_data_ce <= 1'd1;
				builder_uartwishbonebridge_next_state <= 3'd6;
			end
		end
		3'd6: begin
			main_uart_sink_valid <= 1'd1;
			if (main_uart_sink_ready) begin
				main_uart_byte_counter_ce <= 1'd1;
				if ((main_uart_byte_counter == 2'd3)) begin
					main_uart_word_counter_ce <= 1'd1;
					if ((main_uart_word_counter == (main_uart_length - 1'd1))) begin
						builder_uartwishbonebridge_next_state <= 1'd0;
					end else begin
						builder_uartwishbonebridge_next_state <= 3'd5;
						main_uart_byte_counter_reset <= 1'd1;
					end
				end
			end
		end
		default: begin
			if (main_uart_source_valid) begin
				main_uart_cmd_ce <= 1'd1;
				if (((main_uart_source_payload_data == 1'd1) | (main_uart_source_payload_data == 2'd2))) begin
					builder_uartwishbonebridge_next_state <= 1'd1;
				end
				main_uart_byte_counter_reset <= 1'd1;
				main_uart_word_counter_reset <= 1'd1;
			end
			main_uart_is_ongoing <= 1'd1;
		end
	endcase
end
assign main_uart_done = (main_uart_count == 1'd0);
assign main_zero_trigger = (main_value != 1'd0);
assign main_eventmanager_status_w = main_zero_status;
always @(*) begin
	main_zero_clear <= 1'd0;
	if ((main_eventmanager_pending_re & main_eventmanager_pending_r)) begin
		main_zero_clear <= 1'd1;
	end
end
assign main_eventmanager_pending_w = main_zero_pending;
assign main_irq = (main_eventmanager_pending_w & main_eventmanager_storage);
assign main_zero_status = main_zero_trigger;
assign main_interface_dat_w = main_bus_wishbone_dat_w;
assign main_bus_wishbone_dat_r = main_interface_dat_r;
always @(*) begin
	builder_wb2csr_next_state <= 1'd0;
	main_interface_adr <= 14'd0;
	main_interface_we <= 1'd0;
	main_bus_wishbone_ack <= 1'd0;
	builder_wb2csr_next_state <= builder_wb2csr_state;
	case (builder_wb2csr_state)
		1'd1: begin
			main_bus_wishbone_ack <= 1'd1;
			builder_wb2csr_next_state <= 1'd0;
		end
		default: begin
			if ((main_bus_wishbone_cyc & main_bus_wishbone_stb)) begin
				main_interface_adr <= main_bus_wishbone_adr;
				main_interface_we <= main_bus_wishbone_we;
				builder_wb2csr_next_state <= 1'd1;
			end
		end
	endcase
end
assign main_reset = (~cpu_reset);
assign sys_clk = main_clkout_buf0;
assign sys4x_clk = main_clkout_buf1;
assign sys4x_clkb = main_clkout_buf4;
assign sys4x_dqs_clk = main_clkout_buf2;
assign clk200_clk = main_clkout_buf3;
always @(*) begin
	main_a7ddrphy_dqs_serdes_pattern <= 8'd85;
	main_a7ddrphy_dqs_serdes_pattern <= 7'd85;
	if ((main_a7ddrphy_dqs_preamble | main_a7ddrphy_dqs_postamble)) begin
		main_a7ddrphy_dqs_serdes_pattern <= 1'd0;
	end
end
assign main_a7ddrphy_bitslip0_i = main_a7ddrphy_dq_i_data0;
assign main_a7ddrphy_bitslip1_i = main_a7ddrphy_dq_i_data1;
assign main_a7ddrphy_bitslip2_i = main_a7ddrphy_dq_i_data2;
assign main_a7ddrphy_bitslip3_i = main_a7ddrphy_dq_i_data3;
assign main_a7ddrphy_bitslip4_i = main_a7ddrphy_dq_i_data4;
assign main_a7ddrphy_bitslip5_i = main_a7ddrphy_dq_i_data5;
assign main_a7ddrphy_bitslip6_i = main_a7ddrphy_dq_i_data6;
assign main_a7ddrphy_bitslip7_i = main_a7ddrphy_dq_i_data7;
assign main_a7ddrphy_bitslip8_i = main_a7ddrphy_dq_i_data8;
assign main_a7ddrphy_bitslip9_i = main_a7ddrphy_dq_i_data9;
assign main_a7ddrphy_bitslip10_i = main_a7ddrphy_dq_i_data10;
assign main_a7ddrphy_bitslip11_i = main_a7ddrphy_dq_i_data11;
assign main_a7ddrphy_bitslip12_i = main_a7ddrphy_dq_i_data12;
assign main_a7ddrphy_bitslip13_i = main_a7ddrphy_dq_i_data13;
assign main_a7ddrphy_bitslip14_i = main_a7ddrphy_dq_i_data14;
assign main_a7ddrphy_bitslip15_i = main_a7ddrphy_dq_i_data15;
always @(*) begin
	main_a7ddrphy_dfi_p0_rddata <= 32'd0;
	main_a7ddrphy_dfi_p0_rddata[0] <= main_a7ddrphy_bitslip0_o[0];
	main_a7ddrphy_dfi_p0_rddata[16] <= main_a7ddrphy_bitslip0_o[1];
	main_a7ddrphy_dfi_p0_rddata[1] <= main_a7ddrphy_bitslip1_o[0];
	main_a7ddrphy_dfi_p0_rddata[17] <= main_a7ddrphy_bitslip1_o[1];
	main_a7ddrphy_dfi_p0_rddata[2] <= main_a7ddrphy_bitslip2_o[0];
	main_a7ddrphy_dfi_p0_rddata[18] <= main_a7ddrphy_bitslip2_o[1];
	main_a7ddrphy_dfi_p0_rddata[3] <= main_a7ddrphy_bitslip3_o[0];
	main_a7ddrphy_dfi_p0_rddata[19] <= main_a7ddrphy_bitslip3_o[1];
	main_a7ddrphy_dfi_p0_rddata[4] <= main_a7ddrphy_bitslip4_o[0];
	main_a7ddrphy_dfi_p0_rddata[20] <= main_a7ddrphy_bitslip4_o[1];
	main_a7ddrphy_dfi_p0_rddata[5] <= main_a7ddrphy_bitslip5_o[0];
	main_a7ddrphy_dfi_p0_rddata[21] <= main_a7ddrphy_bitslip5_o[1];
	main_a7ddrphy_dfi_p0_rddata[6] <= main_a7ddrphy_bitslip6_o[0];
	main_a7ddrphy_dfi_p0_rddata[22] <= main_a7ddrphy_bitslip6_o[1];
	main_a7ddrphy_dfi_p0_rddata[7] <= main_a7ddrphy_bitslip7_o[0];
	main_a7ddrphy_dfi_p0_rddata[23] <= main_a7ddrphy_bitslip7_o[1];
	main_a7ddrphy_dfi_p0_rddata[8] <= main_a7ddrphy_bitslip8_o[0];
	main_a7ddrphy_dfi_p0_rddata[24] <= main_a7ddrphy_bitslip8_o[1];
	main_a7ddrphy_dfi_p0_rddata[9] <= main_a7ddrphy_bitslip9_o[0];
	main_a7ddrphy_dfi_p0_rddata[25] <= main_a7ddrphy_bitslip9_o[1];
	main_a7ddrphy_dfi_p0_rddata[10] <= main_a7ddrphy_bitslip10_o[0];
	main_a7ddrphy_dfi_p0_rddata[26] <= main_a7ddrphy_bitslip10_o[1];
	main_a7ddrphy_dfi_p0_rddata[11] <= main_a7ddrphy_bitslip11_o[0];
	main_a7ddrphy_dfi_p0_rddata[27] <= main_a7ddrphy_bitslip11_o[1];
	main_a7ddrphy_dfi_p0_rddata[12] <= main_a7ddrphy_bitslip12_o[0];
	main_a7ddrphy_dfi_p0_rddata[28] <= main_a7ddrphy_bitslip12_o[1];
	main_a7ddrphy_dfi_p0_rddata[13] <= main_a7ddrphy_bitslip13_o[0];
	main_a7ddrphy_dfi_p0_rddata[29] <= main_a7ddrphy_bitslip13_o[1];
	main_a7ddrphy_dfi_p0_rddata[14] <= main_a7ddrphy_bitslip14_o[0];
	main_a7ddrphy_dfi_p0_rddata[30] <= main_a7ddrphy_bitslip14_o[1];
	main_a7ddrphy_dfi_p0_rddata[15] <= main_a7ddrphy_bitslip15_o[0];
	main_a7ddrphy_dfi_p0_rddata[31] <= main_a7ddrphy_bitslip15_o[1];
end
always @(*) begin
	main_a7ddrphy_dfi_p1_rddata <= 32'd0;
	main_a7ddrphy_dfi_p1_rddata[0] <= main_a7ddrphy_bitslip0_o[2];
	main_a7ddrphy_dfi_p1_rddata[16] <= main_a7ddrphy_bitslip0_o[3];
	main_a7ddrphy_dfi_p1_rddata[1] <= main_a7ddrphy_bitslip1_o[2];
	main_a7ddrphy_dfi_p1_rddata[17] <= main_a7ddrphy_bitslip1_o[3];
	main_a7ddrphy_dfi_p1_rddata[2] <= main_a7ddrphy_bitslip2_o[2];
	main_a7ddrphy_dfi_p1_rddata[18] <= main_a7ddrphy_bitslip2_o[3];
	main_a7ddrphy_dfi_p1_rddata[3] <= main_a7ddrphy_bitslip3_o[2];
	main_a7ddrphy_dfi_p1_rddata[19] <= main_a7ddrphy_bitslip3_o[3];
	main_a7ddrphy_dfi_p1_rddata[4] <= main_a7ddrphy_bitslip4_o[2];
	main_a7ddrphy_dfi_p1_rddata[20] <= main_a7ddrphy_bitslip4_o[3];
	main_a7ddrphy_dfi_p1_rddata[5] <= main_a7ddrphy_bitslip5_o[2];
	main_a7ddrphy_dfi_p1_rddata[21] <= main_a7ddrphy_bitslip5_o[3];
	main_a7ddrphy_dfi_p1_rddata[6] <= main_a7ddrphy_bitslip6_o[2];
	main_a7ddrphy_dfi_p1_rddata[22] <= main_a7ddrphy_bitslip6_o[3];
	main_a7ddrphy_dfi_p1_rddata[7] <= main_a7ddrphy_bitslip7_o[2];
	main_a7ddrphy_dfi_p1_rddata[23] <= main_a7ddrphy_bitslip7_o[3];
	main_a7ddrphy_dfi_p1_rddata[8] <= main_a7ddrphy_bitslip8_o[2];
	main_a7ddrphy_dfi_p1_rddata[24] <= main_a7ddrphy_bitslip8_o[3];
	main_a7ddrphy_dfi_p1_rddata[9] <= main_a7ddrphy_bitslip9_o[2];
	main_a7ddrphy_dfi_p1_rddata[25] <= main_a7ddrphy_bitslip9_o[3];
	main_a7ddrphy_dfi_p1_rddata[10] <= main_a7ddrphy_bitslip10_o[2];
	main_a7ddrphy_dfi_p1_rddata[26] <= main_a7ddrphy_bitslip10_o[3];
	main_a7ddrphy_dfi_p1_rddata[11] <= main_a7ddrphy_bitslip11_o[2];
	main_a7ddrphy_dfi_p1_rddata[27] <= main_a7ddrphy_bitslip11_o[3];
	main_a7ddrphy_dfi_p1_rddata[12] <= main_a7ddrphy_bitslip12_o[2];
	main_a7ddrphy_dfi_p1_rddata[28] <= main_a7ddrphy_bitslip12_o[3];
	main_a7ddrphy_dfi_p1_rddata[13] <= main_a7ddrphy_bitslip13_o[2];
	main_a7ddrphy_dfi_p1_rddata[29] <= main_a7ddrphy_bitslip13_o[3];
	main_a7ddrphy_dfi_p1_rddata[14] <= main_a7ddrphy_bitslip14_o[2];
	main_a7ddrphy_dfi_p1_rddata[30] <= main_a7ddrphy_bitslip14_o[3];
	main_a7ddrphy_dfi_p1_rddata[15] <= main_a7ddrphy_bitslip15_o[2];
	main_a7ddrphy_dfi_p1_rddata[31] <= main_a7ddrphy_bitslip15_o[3];
end
always @(*) begin
	main_a7ddrphy_dfi_p2_rddata <= 32'd0;
	main_a7ddrphy_dfi_p2_rddata[0] <= main_a7ddrphy_bitslip0_o[4];
	main_a7ddrphy_dfi_p2_rddata[16] <= main_a7ddrphy_bitslip0_o[5];
	main_a7ddrphy_dfi_p2_rddata[1] <= main_a7ddrphy_bitslip1_o[4];
	main_a7ddrphy_dfi_p2_rddata[17] <= main_a7ddrphy_bitslip1_o[5];
	main_a7ddrphy_dfi_p2_rddata[2] <= main_a7ddrphy_bitslip2_o[4];
	main_a7ddrphy_dfi_p2_rddata[18] <= main_a7ddrphy_bitslip2_o[5];
	main_a7ddrphy_dfi_p2_rddata[3] <= main_a7ddrphy_bitslip3_o[4];
	main_a7ddrphy_dfi_p2_rddata[19] <= main_a7ddrphy_bitslip3_o[5];
	main_a7ddrphy_dfi_p2_rddata[4] <= main_a7ddrphy_bitslip4_o[4];
	main_a7ddrphy_dfi_p2_rddata[20] <= main_a7ddrphy_bitslip4_o[5];
	main_a7ddrphy_dfi_p2_rddata[5] <= main_a7ddrphy_bitslip5_o[4];
	main_a7ddrphy_dfi_p2_rddata[21] <= main_a7ddrphy_bitslip5_o[5];
	main_a7ddrphy_dfi_p2_rddata[6] <= main_a7ddrphy_bitslip6_o[4];
	main_a7ddrphy_dfi_p2_rddata[22] <= main_a7ddrphy_bitslip6_o[5];
	main_a7ddrphy_dfi_p2_rddata[7] <= main_a7ddrphy_bitslip7_o[4];
	main_a7ddrphy_dfi_p2_rddata[23] <= main_a7ddrphy_bitslip7_o[5];
	main_a7ddrphy_dfi_p2_rddata[8] <= main_a7ddrphy_bitslip8_o[4];
	main_a7ddrphy_dfi_p2_rddata[24] <= main_a7ddrphy_bitslip8_o[5];
	main_a7ddrphy_dfi_p2_rddata[9] <= main_a7ddrphy_bitslip9_o[4];
	main_a7ddrphy_dfi_p2_rddata[25] <= main_a7ddrphy_bitslip9_o[5];
	main_a7ddrphy_dfi_p2_rddata[10] <= main_a7ddrphy_bitslip10_o[4];
	main_a7ddrphy_dfi_p2_rddata[26] <= main_a7ddrphy_bitslip10_o[5];
	main_a7ddrphy_dfi_p2_rddata[11] <= main_a7ddrphy_bitslip11_o[4];
	main_a7ddrphy_dfi_p2_rddata[27] <= main_a7ddrphy_bitslip11_o[5];
	main_a7ddrphy_dfi_p2_rddata[12] <= main_a7ddrphy_bitslip12_o[4];
	main_a7ddrphy_dfi_p2_rddata[28] <= main_a7ddrphy_bitslip12_o[5];
	main_a7ddrphy_dfi_p2_rddata[13] <= main_a7ddrphy_bitslip13_o[4];
	main_a7ddrphy_dfi_p2_rddata[29] <= main_a7ddrphy_bitslip13_o[5];
	main_a7ddrphy_dfi_p2_rddata[14] <= main_a7ddrphy_bitslip14_o[4];
	main_a7ddrphy_dfi_p2_rddata[30] <= main_a7ddrphy_bitslip14_o[5];
	main_a7ddrphy_dfi_p2_rddata[15] <= main_a7ddrphy_bitslip15_o[4];
	main_a7ddrphy_dfi_p2_rddata[31] <= main_a7ddrphy_bitslip15_o[5];
end
always @(*) begin
	main_a7ddrphy_dfi_p3_rddata <= 32'd0;
	main_a7ddrphy_dfi_p3_rddata[0] <= main_a7ddrphy_bitslip0_o[6];
	main_a7ddrphy_dfi_p3_rddata[16] <= main_a7ddrphy_bitslip0_o[7];
	main_a7ddrphy_dfi_p3_rddata[1] <= main_a7ddrphy_bitslip1_o[6];
	main_a7ddrphy_dfi_p3_rddata[17] <= main_a7ddrphy_bitslip1_o[7];
	main_a7ddrphy_dfi_p3_rddata[2] <= main_a7ddrphy_bitslip2_o[6];
	main_a7ddrphy_dfi_p3_rddata[18] <= main_a7ddrphy_bitslip2_o[7];
	main_a7ddrphy_dfi_p3_rddata[3] <= main_a7ddrphy_bitslip3_o[6];
	main_a7ddrphy_dfi_p3_rddata[19] <= main_a7ddrphy_bitslip3_o[7];
	main_a7ddrphy_dfi_p3_rddata[4] <= main_a7ddrphy_bitslip4_o[6];
	main_a7ddrphy_dfi_p3_rddata[20] <= main_a7ddrphy_bitslip4_o[7];
	main_a7ddrphy_dfi_p3_rddata[5] <= main_a7ddrphy_bitslip5_o[6];
	main_a7ddrphy_dfi_p3_rddata[21] <= main_a7ddrphy_bitslip5_o[7];
	main_a7ddrphy_dfi_p3_rddata[6] <= main_a7ddrphy_bitslip6_o[6];
	main_a7ddrphy_dfi_p3_rddata[22] <= main_a7ddrphy_bitslip6_o[7];
	main_a7ddrphy_dfi_p3_rddata[7] <= main_a7ddrphy_bitslip7_o[6];
	main_a7ddrphy_dfi_p3_rddata[23] <= main_a7ddrphy_bitslip7_o[7];
	main_a7ddrphy_dfi_p3_rddata[8] <= main_a7ddrphy_bitslip8_o[6];
	main_a7ddrphy_dfi_p3_rddata[24] <= main_a7ddrphy_bitslip8_o[7];
	main_a7ddrphy_dfi_p3_rddata[9] <= main_a7ddrphy_bitslip9_o[6];
	main_a7ddrphy_dfi_p3_rddata[25] <= main_a7ddrphy_bitslip9_o[7];
	main_a7ddrphy_dfi_p3_rddata[10] <= main_a7ddrphy_bitslip10_o[6];
	main_a7ddrphy_dfi_p3_rddata[26] <= main_a7ddrphy_bitslip10_o[7];
	main_a7ddrphy_dfi_p3_rddata[11] <= main_a7ddrphy_bitslip11_o[6];
	main_a7ddrphy_dfi_p3_rddata[27] <= main_a7ddrphy_bitslip11_o[7];
	main_a7ddrphy_dfi_p3_rddata[12] <= main_a7ddrphy_bitslip12_o[6];
	main_a7ddrphy_dfi_p3_rddata[28] <= main_a7ddrphy_bitslip12_o[7];
	main_a7ddrphy_dfi_p3_rddata[13] <= main_a7ddrphy_bitslip13_o[6];
	main_a7ddrphy_dfi_p3_rddata[29] <= main_a7ddrphy_bitslip13_o[7];
	main_a7ddrphy_dfi_p3_rddata[14] <= main_a7ddrphy_bitslip14_o[6];
	main_a7ddrphy_dfi_p3_rddata[30] <= main_a7ddrphy_bitslip14_o[7];
	main_a7ddrphy_dfi_p3_rddata[15] <= main_a7ddrphy_bitslip15_o[6];
	main_a7ddrphy_dfi_p3_rddata[31] <= main_a7ddrphy_bitslip15_o[7];
end
assign main_a7ddrphy_oe = ((main_a7ddrphy_last_wrdata_en[1] | main_a7ddrphy_last_wrdata_en[2]) | main_a7ddrphy_last_wrdata_en[3]);
assign main_a7ddrphy_dqs_preamble = (main_a7ddrphy_last_wrdata_en[1] & (~main_a7ddrphy_last_wrdata_en[2]));
assign main_a7ddrphy_dqs_postamble = (main_a7ddrphy_last_wrdata_en[3] & (~main_a7ddrphy_last_wrdata_en[2]));
assign main_a7ddrphy_dfi_p0_address = main_sdram_master_p0_address;
assign main_a7ddrphy_dfi_p0_bank = main_sdram_master_p0_bank;
assign main_a7ddrphy_dfi_p0_cas_n = main_sdram_master_p0_cas_n;
assign main_a7ddrphy_dfi_p0_cs_n = main_sdram_master_p0_cs_n;
assign main_a7ddrphy_dfi_p0_ras_n = main_sdram_master_p0_ras_n;
assign main_a7ddrphy_dfi_p0_we_n = main_sdram_master_p0_we_n;
assign main_a7ddrphy_dfi_p0_cke = main_sdram_master_p0_cke;
assign main_a7ddrphy_dfi_p0_odt = main_sdram_master_p0_odt;
assign main_a7ddrphy_dfi_p0_reset_n = main_sdram_master_p0_reset_n;
assign main_a7ddrphy_dfi_p0_act_n = main_sdram_master_p0_act_n;
assign main_a7ddrphy_dfi_p0_wrdata = main_sdram_master_p0_wrdata;
assign main_a7ddrphy_dfi_p0_wrdata_en = main_sdram_master_p0_wrdata_en;
assign main_a7ddrphy_dfi_p0_wrdata_mask = main_sdram_master_p0_wrdata_mask;
assign main_a7ddrphy_dfi_p0_rddata_en = main_sdram_master_p0_rddata_en;
assign main_sdram_master_p0_rddata = main_a7ddrphy_dfi_p0_rddata;
assign main_sdram_master_p0_rddata_valid = main_a7ddrphy_dfi_p0_rddata_valid;
assign main_a7ddrphy_dfi_p1_address = main_sdram_master_p1_address;
assign main_a7ddrphy_dfi_p1_bank = main_sdram_master_p1_bank;
assign main_a7ddrphy_dfi_p1_cas_n = main_sdram_master_p1_cas_n;
assign main_a7ddrphy_dfi_p1_cs_n = main_sdram_master_p1_cs_n;
assign main_a7ddrphy_dfi_p1_ras_n = main_sdram_master_p1_ras_n;
assign main_a7ddrphy_dfi_p1_we_n = main_sdram_master_p1_we_n;
assign main_a7ddrphy_dfi_p1_cke = main_sdram_master_p1_cke;
assign main_a7ddrphy_dfi_p1_odt = main_sdram_master_p1_odt;
assign main_a7ddrphy_dfi_p1_reset_n = main_sdram_master_p1_reset_n;
assign main_a7ddrphy_dfi_p1_act_n = main_sdram_master_p1_act_n;
assign main_a7ddrphy_dfi_p1_wrdata = main_sdram_master_p1_wrdata;
assign main_a7ddrphy_dfi_p1_wrdata_en = main_sdram_master_p1_wrdata_en;
assign main_a7ddrphy_dfi_p1_wrdata_mask = main_sdram_master_p1_wrdata_mask;
assign main_a7ddrphy_dfi_p1_rddata_en = main_sdram_master_p1_rddata_en;
assign main_sdram_master_p1_rddata = main_a7ddrphy_dfi_p1_rddata;
assign main_sdram_master_p1_rddata_valid = main_a7ddrphy_dfi_p1_rddata_valid;
assign main_a7ddrphy_dfi_p2_address = main_sdram_master_p2_address;
assign main_a7ddrphy_dfi_p2_bank = main_sdram_master_p2_bank;
assign main_a7ddrphy_dfi_p2_cas_n = main_sdram_master_p2_cas_n;
assign main_a7ddrphy_dfi_p2_cs_n = main_sdram_master_p2_cs_n;
assign main_a7ddrphy_dfi_p2_ras_n = main_sdram_master_p2_ras_n;
assign main_a7ddrphy_dfi_p2_we_n = main_sdram_master_p2_we_n;
assign main_a7ddrphy_dfi_p2_cke = main_sdram_master_p2_cke;
assign main_a7ddrphy_dfi_p2_odt = main_sdram_master_p2_odt;
assign main_a7ddrphy_dfi_p2_reset_n = main_sdram_master_p2_reset_n;
assign main_a7ddrphy_dfi_p2_act_n = main_sdram_master_p2_act_n;
assign main_a7ddrphy_dfi_p2_wrdata = main_sdram_master_p2_wrdata;
assign main_a7ddrphy_dfi_p2_wrdata_en = main_sdram_master_p2_wrdata_en;
assign main_a7ddrphy_dfi_p2_wrdata_mask = main_sdram_master_p2_wrdata_mask;
assign main_a7ddrphy_dfi_p2_rddata_en = main_sdram_master_p2_rddata_en;
assign main_sdram_master_p2_rddata = main_a7ddrphy_dfi_p2_rddata;
assign main_sdram_master_p2_rddata_valid = main_a7ddrphy_dfi_p2_rddata_valid;
assign main_a7ddrphy_dfi_p3_address = main_sdram_master_p3_address;
assign main_a7ddrphy_dfi_p3_bank = main_sdram_master_p3_bank;
assign main_a7ddrphy_dfi_p3_cas_n = main_sdram_master_p3_cas_n;
assign main_a7ddrphy_dfi_p3_cs_n = main_sdram_master_p3_cs_n;
assign main_a7ddrphy_dfi_p3_ras_n = main_sdram_master_p3_ras_n;
assign main_a7ddrphy_dfi_p3_we_n = main_sdram_master_p3_we_n;
assign main_a7ddrphy_dfi_p3_cke = main_sdram_master_p3_cke;
assign main_a7ddrphy_dfi_p3_odt = main_sdram_master_p3_odt;
assign main_a7ddrphy_dfi_p3_reset_n = main_sdram_master_p3_reset_n;
assign main_a7ddrphy_dfi_p3_act_n = main_sdram_master_p3_act_n;
assign main_a7ddrphy_dfi_p3_wrdata = main_sdram_master_p3_wrdata;
assign main_a7ddrphy_dfi_p3_wrdata_en = main_sdram_master_p3_wrdata_en;
assign main_a7ddrphy_dfi_p3_wrdata_mask = main_sdram_master_p3_wrdata_mask;
assign main_a7ddrphy_dfi_p3_rddata_en = main_sdram_master_p3_rddata_en;
assign main_sdram_master_p3_rddata = main_a7ddrphy_dfi_p3_rddata;
assign main_sdram_master_p3_rddata_valid = main_a7ddrphy_dfi_p3_rddata_valid;
assign main_sdram_slave_p0_address = main_sdram_dfi_p0_address;
assign main_sdram_slave_p0_bank = main_sdram_dfi_p0_bank;
assign main_sdram_slave_p0_cas_n = main_sdram_dfi_p0_cas_n;
assign main_sdram_slave_p0_cs_n = main_sdram_dfi_p0_cs_n;
assign main_sdram_slave_p0_ras_n = main_sdram_dfi_p0_ras_n;
assign main_sdram_slave_p0_we_n = main_sdram_dfi_p0_we_n;
assign main_sdram_slave_p0_cke = main_sdram_dfi_p0_cke;
assign main_sdram_slave_p0_odt = main_sdram_dfi_p0_odt;
assign main_sdram_slave_p0_reset_n = main_sdram_dfi_p0_reset_n;
assign main_sdram_slave_p0_act_n = main_sdram_dfi_p0_act_n;
assign main_sdram_slave_p0_wrdata = main_sdram_dfi_p0_wrdata;
assign main_sdram_slave_p0_wrdata_en = main_sdram_dfi_p0_wrdata_en;
assign main_sdram_slave_p0_wrdata_mask = main_sdram_dfi_p0_wrdata_mask;
assign main_sdram_slave_p0_rddata_en = main_sdram_dfi_p0_rddata_en;
assign main_sdram_dfi_p0_rddata = main_sdram_slave_p0_rddata;
assign main_sdram_dfi_p0_rddata_valid = main_sdram_slave_p0_rddata_valid;
assign main_sdram_slave_p1_address = main_sdram_dfi_p1_address;
assign main_sdram_slave_p1_bank = main_sdram_dfi_p1_bank;
assign main_sdram_slave_p1_cas_n = main_sdram_dfi_p1_cas_n;
assign main_sdram_slave_p1_cs_n = main_sdram_dfi_p1_cs_n;
assign main_sdram_slave_p1_ras_n = main_sdram_dfi_p1_ras_n;
assign main_sdram_slave_p1_we_n = main_sdram_dfi_p1_we_n;
assign main_sdram_slave_p1_cke = main_sdram_dfi_p1_cke;
assign main_sdram_slave_p1_odt = main_sdram_dfi_p1_odt;
assign main_sdram_slave_p1_reset_n = main_sdram_dfi_p1_reset_n;
assign main_sdram_slave_p1_act_n = main_sdram_dfi_p1_act_n;
assign main_sdram_slave_p1_wrdata = main_sdram_dfi_p1_wrdata;
assign main_sdram_slave_p1_wrdata_en = main_sdram_dfi_p1_wrdata_en;
assign main_sdram_slave_p1_wrdata_mask = main_sdram_dfi_p1_wrdata_mask;
assign main_sdram_slave_p1_rddata_en = main_sdram_dfi_p1_rddata_en;
assign main_sdram_dfi_p1_rddata = main_sdram_slave_p1_rddata;
assign main_sdram_dfi_p1_rddata_valid = main_sdram_slave_p1_rddata_valid;
assign main_sdram_slave_p2_address = main_sdram_dfi_p2_address;
assign main_sdram_slave_p2_bank = main_sdram_dfi_p2_bank;
assign main_sdram_slave_p2_cas_n = main_sdram_dfi_p2_cas_n;
assign main_sdram_slave_p2_cs_n = main_sdram_dfi_p2_cs_n;
assign main_sdram_slave_p2_ras_n = main_sdram_dfi_p2_ras_n;
assign main_sdram_slave_p2_we_n = main_sdram_dfi_p2_we_n;
assign main_sdram_slave_p2_cke = main_sdram_dfi_p2_cke;
assign main_sdram_slave_p2_odt = main_sdram_dfi_p2_odt;
assign main_sdram_slave_p2_reset_n = main_sdram_dfi_p2_reset_n;
assign main_sdram_slave_p2_act_n = main_sdram_dfi_p2_act_n;
assign main_sdram_slave_p2_wrdata = main_sdram_dfi_p2_wrdata;
assign main_sdram_slave_p2_wrdata_en = main_sdram_dfi_p2_wrdata_en;
assign main_sdram_slave_p2_wrdata_mask = main_sdram_dfi_p2_wrdata_mask;
assign main_sdram_slave_p2_rddata_en = main_sdram_dfi_p2_rddata_en;
assign main_sdram_dfi_p2_rddata = main_sdram_slave_p2_rddata;
assign main_sdram_dfi_p2_rddata_valid = main_sdram_slave_p2_rddata_valid;
assign main_sdram_slave_p3_address = main_sdram_dfi_p3_address;
assign main_sdram_slave_p3_bank = main_sdram_dfi_p3_bank;
assign main_sdram_slave_p3_cas_n = main_sdram_dfi_p3_cas_n;
assign main_sdram_slave_p3_cs_n = main_sdram_dfi_p3_cs_n;
assign main_sdram_slave_p3_ras_n = main_sdram_dfi_p3_ras_n;
assign main_sdram_slave_p3_we_n = main_sdram_dfi_p3_we_n;
assign main_sdram_slave_p3_cke = main_sdram_dfi_p3_cke;
assign main_sdram_slave_p3_odt = main_sdram_dfi_p3_odt;
assign main_sdram_slave_p3_reset_n = main_sdram_dfi_p3_reset_n;
assign main_sdram_slave_p3_act_n = main_sdram_dfi_p3_act_n;
assign main_sdram_slave_p3_wrdata = main_sdram_dfi_p3_wrdata;
assign main_sdram_slave_p3_wrdata_en = main_sdram_dfi_p3_wrdata_en;
assign main_sdram_slave_p3_wrdata_mask = main_sdram_dfi_p3_wrdata_mask;
assign main_sdram_slave_p3_rddata_en = main_sdram_dfi_p3_rddata_en;
assign main_sdram_dfi_p3_rddata = main_sdram_slave_p3_rddata;
assign main_sdram_dfi_p3_rddata_valid = main_sdram_slave_p3_rddata_valid;
always @(*) begin
	main_sdram_master_p0_address <= 14'd0;
	main_sdram_master_p0_bank <= 3'd0;
	main_sdram_master_p0_cas_n <= 1'd1;
	main_sdram_master_p0_cs_n <= 1'd1;
	main_sdram_master_p0_ras_n <= 1'd1;
	main_sdram_master_p0_we_n <= 1'd1;
	main_sdram_master_p0_cke <= 1'd0;
	main_sdram_master_p0_odt <= 1'd0;
	main_sdram_master_p0_reset_n <= 1'd0;
	main_sdram_master_p0_act_n <= 1'd1;
	main_sdram_master_p0_wrdata <= 32'd0;
	main_sdram_inti_p1_rddata <= 32'd0;
	main_sdram_master_p0_wrdata_en <= 1'd0;
	main_sdram_inti_p1_rddata_valid <= 1'd0;
	main_sdram_master_p0_wrdata_mask <= 4'd0;
	main_sdram_master_p0_rddata_en <= 1'd0;
	main_sdram_master_p1_address <= 14'd0;
	main_sdram_master_p1_bank <= 3'd0;
	main_sdram_master_p1_cas_n <= 1'd1;
	main_sdram_master_p1_cs_n <= 1'd1;
	main_sdram_master_p1_ras_n <= 1'd1;
	main_sdram_master_p1_we_n <= 1'd1;
	main_sdram_master_p1_cke <= 1'd0;
	main_sdram_master_p1_odt <= 1'd0;
	main_sdram_master_p1_reset_n <= 1'd0;
	main_sdram_master_p1_act_n <= 1'd1;
	main_sdram_master_p1_wrdata <= 32'd0;
	main_sdram_inti_p2_rddata <= 32'd0;
	main_sdram_master_p1_wrdata_en <= 1'd0;
	main_sdram_inti_p2_rddata_valid <= 1'd0;
	main_sdram_master_p1_wrdata_mask <= 4'd0;
	main_sdram_master_p1_rddata_en <= 1'd0;
	main_sdram_master_p2_address <= 14'd0;
	main_sdram_master_p2_bank <= 3'd0;
	main_sdram_master_p2_cas_n <= 1'd1;
	main_sdram_master_p2_cs_n <= 1'd1;
	main_sdram_master_p2_ras_n <= 1'd1;
	main_sdram_master_p2_we_n <= 1'd1;
	main_sdram_master_p2_cke <= 1'd0;
	main_sdram_master_p2_odt <= 1'd0;
	main_sdram_master_p2_reset_n <= 1'd0;
	main_sdram_master_p2_act_n <= 1'd1;
	main_sdram_master_p2_wrdata <= 32'd0;
	main_sdram_inti_p3_rddata <= 32'd0;
	main_sdram_master_p2_wrdata_en <= 1'd0;
	main_sdram_inti_p3_rddata_valid <= 1'd0;
	main_sdram_master_p2_wrdata_mask <= 4'd0;
	main_sdram_master_p2_rddata_en <= 1'd0;
	main_sdram_master_p3_address <= 14'd0;
	main_sdram_master_p3_bank <= 3'd0;
	main_sdram_master_p3_cas_n <= 1'd1;
	main_sdram_master_p3_cs_n <= 1'd1;
	main_sdram_master_p3_ras_n <= 1'd1;
	main_sdram_master_p3_we_n <= 1'd1;
	main_sdram_master_p3_cke <= 1'd0;
	main_sdram_master_p3_odt <= 1'd0;
	main_sdram_master_p3_reset_n <= 1'd0;
	main_sdram_master_p3_act_n <= 1'd1;
	main_sdram_master_p3_wrdata <= 32'd0;
	main_sdram_master_p3_wrdata_en <= 1'd0;
	main_sdram_master_p3_wrdata_mask <= 4'd0;
	main_sdram_master_p3_rddata_en <= 1'd0;
	main_sdram_slave_p0_rddata <= 32'd0;
	main_sdram_slave_p0_rddata_valid <= 1'd0;
	main_sdram_slave_p1_rddata <= 32'd0;
	main_sdram_slave_p1_rddata_valid <= 1'd0;
	main_sdram_slave_p2_rddata <= 32'd0;
	main_sdram_slave_p2_rddata_valid <= 1'd0;
	main_sdram_slave_p3_rddata <= 32'd0;
	main_sdram_slave_p3_rddata_valid <= 1'd0;
	main_sdram_inti_p0_rddata <= 32'd0;
	main_sdram_inti_p0_rddata_valid <= 1'd0;
	if (main_sdram_storage[0]) begin
		main_sdram_master_p0_address <= main_sdram_slave_p0_address;
		main_sdram_master_p0_bank <= main_sdram_slave_p0_bank;
		main_sdram_master_p0_cas_n <= main_sdram_slave_p0_cas_n;
		main_sdram_master_p0_cs_n <= main_sdram_slave_p0_cs_n;
		main_sdram_master_p0_ras_n <= main_sdram_slave_p0_ras_n;
		main_sdram_master_p0_we_n <= main_sdram_slave_p0_we_n;
		main_sdram_master_p0_cke <= main_sdram_slave_p0_cke;
		main_sdram_master_p0_odt <= main_sdram_slave_p0_odt;
		main_sdram_master_p0_reset_n <= main_sdram_slave_p0_reset_n;
		main_sdram_master_p0_act_n <= main_sdram_slave_p0_act_n;
		main_sdram_master_p0_wrdata <= main_sdram_slave_p0_wrdata;
		main_sdram_master_p0_wrdata_en <= main_sdram_slave_p0_wrdata_en;
		main_sdram_master_p0_wrdata_mask <= main_sdram_slave_p0_wrdata_mask;
		main_sdram_master_p0_rddata_en <= main_sdram_slave_p0_rddata_en;
		main_sdram_slave_p0_rddata <= main_sdram_master_p0_rddata;
		main_sdram_slave_p0_rddata_valid <= main_sdram_master_p0_rddata_valid;
		main_sdram_master_p1_address <= main_sdram_slave_p1_address;
		main_sdram_master_p1_bank <= main_sdram_slave_p1_bank;
		main_sdram_master_p1_cas_n <= main_sdram_slave_p1_cas_n;
		main_sdram_master_p1_cs_n <= main_sdram_slave_p1_cs_n;
		main_sdram_master_p1_ras_n <= main_sdram_slave_p1_ras_n;
		main_sdram_master_p1_we_n <= main_sdram_slave_p1_we_n;
		main_sdram_master_p1_cke <= main_sdram_slave_p1_cke;
		main_sdram_master_p1_odt <= main_sdram_slave_p1_odt;
		main_sdram_master_p1_reset_n <= main_sdram_slave_p1_reset_n;
		main_sdram_master_p1_act_n <= main_sdram_slave_p1_act_n;
		main_sdram_master_p1_wrdata <= main_sdram_slave_p1_wrdata;
		main_sdram_master_p1_wrdata_en <= main_sdram_slave_p1_wrdata_en;
		main_sdram_master_p1_wrdata_mask <= main_sdram_slave_p1_wrdata_mask;
		main_sdram_master_p1_rddata_en <= main_sdram_slave_p1_rddata_en;
		main_sdram_slave_p1_rddata <= main_sdram_master_p1_rddata;
		main_sdram_slave_p1_rddata_valid <= main_sdram_master_p1_rddata_valid;
		main_sdram_master_p2_address <= main_sdram_slave_p2_address;
		main_sdram_master_p2_bank <= main_sdram_slave_p2_bank;
		main_sdram_master_p2_cas_n <= main_sdram_slave_p2_cas_n;
		main_sdram_master_p2_cs_n <= main_sdram_slave_p2_cs_n;
		main_sdram_master_p2_ras_n <= main_sdram_slave_p2_ras_n;
		main_sdram_master_p2_we_n <= main_sdram_slave_p2_we_n;
		main_sdram_master_p2_cke <= main_sdram_slave_p2_cke;
		main_sdram_master_p2_odt <= main_sdram_slave_p2_odt;
		main_sdram_master_p2_reset_n <= main_sdram_slave_p2_reset_n;
		main_sdram_master_p2_act_n <= main_sdram_slave_p2_act_n;
		main_sdram_master_p2_wrdata <= main_sdram_slave_p2_wrdata;
		main_sdram_master_p2_wrdata_en <= main_sdram_slave_p2_wrdata_en;
		main_sdram_master_p2_wrdata_mask <= main_sdram_slave_p2_wrdata_mask;
		main_sdram_master_p2_rddata_en <= main_sdram_slave_p2_rddata_en;
		main_sdram_slave_p2_rddata <= main_sdram_master_p2_rddata;
		main_sdram_slave_p2_rddata_valid <= main_sdram_master_p2_rddata_valid;
		main_sdram_master_p3_address <= main_sdram_slave_p3_address;
		main_sdram_master_p3_bank <= main_sdram_slave_p3_bank;
		main_sdram_master_p3_cas_n <= main_sdram_slave_p3_cas_n;
		main_sdram_master_p3_cs_n <= main_sdram_slave_p3_cs_n;
		main_sdram_master_p3_ras_n <= main_sdram_slave_p3_ras_n;
		main_sdram_master_p3_we_n <= main_sdram_slave_p3_we_n;
		main_sdram_master_p3_cke <= main_sdram_slave_p3_cke;
		main_sdram_master_p3_odt <= main_sdram_slave_p3_odt;
		main_sdram_master_p3_reset_n <= main_sdram_slave_p3_reset_n;
		main_sdram_master_p3_act_n <= main_sdram_slave_p3_act_n;
		main_sdram_master_p3_wrdata <= main_sdram_slave_p3_wrdata;
		main_sdram_master_p3_wrdata_en <= main_sdram_slave_p3_wrdata_en;
		main_sdram_master_p3_wrdata_mask <= main_sdram_slave_p3_wrdata_mask;
		main_sdram_master_p3_rddata_en <= main_sdram_slave_p3_rddata_en;
		main_sdram_slave_p3_rddata <= main_sdram_master_p3_rddata;
		main_sdram_slave_p3_rddata_valid <= main_sdram_master_p3_rddata_valid;
	end else begin
		main_sdram_master_p0_address <= main_sdram_inti_p0_address;
		main_sdram_master_p0_bank <= main_sdram_inti_p0_bank;
		main_sdram_master_p0_cas_n <= main_sdram_inti_p0_cas_n;
		main_sdram_master_p0_cs_n <= main_sdram_inti_p0_cs_n;
		main_sdram_master_p0_ras_n <= main_sdram_inti_p0_ras_n;
		main_sdram_master_p0_we_n <= main_sdram_inti_p0_we_n;
		main_sdram_master_p0_cke <= main_sdram_inti_p0_cke;
		main_sdram_master_p0_odt <= main_sdram_inti_p0_odt;
		main_sdram_master_p0_reset_n <= main_sdram_inti_p0_reset_n;
		main_sdram_master_p0_act_n <= main_sdram_inti_p0_act_n;
		main_sdram_master_p0_wrdata <= main_sdram_inti_p0_wrdata;
		main_sdram_master_p0_wrdata_en <= main_sdram_inti_p0_wrdata_en;
		main_sdram_master_p0_wrdata_mask <= main_sdram_inti_p0_wrdata_mask;
		main_sdram_master_p0_rddata_en <= main_sdram_inti_p0_rddata_en;
		main_sdram_inti_p0_rddata <= main_sdram_master_p0_rddata;
		main_sdram_inti_p0_rddata_valid <= main_sdram_master_p0_rddata_valid;
		main_sdram_master_p1_address <= main_sdram_inti_p1_address;
		main_sdram_master_p1_bank <= main_sdram_inti_p1_bank;
		main_sdram_master_p1_cas_n <= main_sdram_inti_p1_cas_n;
		main_sdram_master_p1_cs_n <= main_sdram_inti_p1_cs_n;
		main_sdram_master_p1_ras_n <= main_sdram_inti_p1_ras_n;
		main_sdram_master_p1_we_n <= main_sdram_inti_p1_we_n;
		main_sdram_master_p1_cke <= main_sdram_inti_p1_cke;
		main_sdram_master_p1_odt <= main_sdram_inti_p1_odt;
		main_sdram_master_p1_reset_n <= main_sdram_inti_p1_reset_n;
		main_sdram_master_p1_act_n <= main_sdram_inti_p1_act_n;
		main_sdram_master_p1_wrdata <= main_sdram_inti_p1_wrdata;
		main_sdram_master_p1_wrdata_en <= main_sdram_inti_p1_wrdata_en;
		main_sdram_master_p1_wrdata_mask <= main_sdram_inti_p1_wrdata_mask;
		main_sdram_master_p1_rddata_en <= main_sdram_inti_p1_rddata_en;
		main_sdram_inti_p1_rddata <= main_sdram_master_p1_rddata;
		main_sdram_inti_p1_rddata_valid <= main_sdram_master_p1_rddata_valid;
		main_sdram_master_p2_address <= main_sdram_inti_p2_address;
		main_sdram_master_p2_bank <= main_sdram_inti_p2_bank;
		main_sdram_master_p2_cas_n <= main_sdram_inti_p2_cas_n;
		main_sdram_master_p2_cs_n <= main_sdram_inti_p2_cs_n;
		main_sdram_master_p2_ras_n <= main_sdram_inti_p2_ras_n;
		main_sdram_master_p2_we_n <= main_sdram_inti_p2_we_n;
		main_sdram_master_p2_cke <= main_sdram_inti_p2_cke;
		main_sdram_master_p2_odt <= main_sdram_inti_p2_odt;
		main_sdram_master_p2_reset_n <= main_sdram_inti_p2_reset_n;
		main_sdram_master_p2_act_n <= main_sdram_inti_p2_act_n;
		main_sdram_master_p2_wrdata <= main_sdram_inti_p2_wrdata;
		main_sdram_master_p2_wrdata_en <= main_sdram_inti_p2_wrdata_en;
		main_sdram_master_p2_wrdata_mask <= main_sdram_inti_p2_wrdata_mask;
		main_sdram_master_p2_rddata_en <= main_sdram_inti_p2_rddata_en;
		main_sdram_inti_p2_rddata <= main_sdram_master_p2_rddata;
		main_sdram_inti_p2_rddata_valid <= main_sdram_master_p2_rddata_valid;
		main_sdram_master_p3_address <= main_sdram_inti_p3_address;
		main_sdram_master_p3_bank <= main_sdram_inti_p3_bank;
		main_sdram_master_p3_cas_n <= main_sdram_inti_p3_cas_n;
		main_sdram_master_p3_cs_n <= main_sdram_inti_p3_cs_n;
		main_sdram_master_p3_ras_n <= main_sdram_inti_p3_ras_n;
		main_sdram_master_p3_we_n <= main_sdram_inti_p3_we_n;
		main_sdram_master_p3_cke <= main_sdram_inti_p3_cke;
		main_sdram_master_p3_odt <= main_sdram_inti_p3_odt;
		main_sdram_master_p3_reset_n <= main_sdram_inti_p3_reset_n;
		main_sdram_master_p3_act_n <= main_sdram_inti_p3_act_n;
		main_sdram_master_p3_wrdata <= main_sdram_inti_p3_wrdata;
		main_sdram_master_p3_wrdata_en <= main_sdram_inti_p3_wrdata_en;
		main_sdram_master_p3_wrdata_mask <= main_sdram_inti_p3_wrdata_mask;
		main_sdram_master_p3_rddata_en <= main_sdram_inti_p3_rddata_en;
		main_sdram_inti_p3_rddata <= main_sdram_master_p3_rddata;
		main_sdram_inti_p3_rddata_valid <= main_sdram_master_p3_rddata_valid;
	end
end
assign main_sdram_inti_p0_cke = main_sdram_storage[1];
assign main_sdram_inti_p1_cke = main_sdram_storage[1];
assign main_sdram_inti_p2_cke = main_sdram_storage[1];
assign main_sdram_inti_p3_cke = main_sdram_storage[1];
assign main_sdram_inti_p0_odt = main_sdram_storage[2];
assign main_sdram_inti_p1_odt = main_sdram_storage[2];
assign main_sdram_inti_p2_odt = main_sdram_storage[2];
assign main_sdram_inti_p3_odt = main_sdram_storage[2];
assign main_sdram_inti_p0_reset_n = main_sdram_storage[3];
assign main_sdram_inti_p1_reset_n = main_sdram_storage[3];
assign main_sdram_inti_p2_reset_n = main_sdram_storage[3];
assign main_sdram_inti_p3_reset_n = main_sdram_storage[3];
always @(*) begin
	main_sdram_inti_p0_cs_n <= 1'd1;
	main_sdram_inti_p0_ras_n <= 1'd1;
	main_sdram_inti_p0_we_n <= 1'd1;
	main_sdram_inti_p0_cas_n <= 1'd1;
	if (main_sdram_phaseinjector0_command_issue_re) begin
		main_sdram_inti_p0_cs_n <= {1{(~main_sdram_phaseinjector0_command_storage[0])}};
		main_sdram_inti_p0_we_n <= (~main_sdram_phaseinjector0_command_storage[1]);
		main_sdram_inti_p0_cas_n <= (~main_sdram_phaseinjector0_command_storage[2]);
		main_sdram_inti_p0_ras_n <= (~main_sdram_phaseinjector0_command_storage[3]);
	end else begin
		main_sdram_inti_p0_cs_n <= {1{1'd1}};
		main_sdram_inti_p0_we_n <= 1'd1;
		main_sdram_inti_p0_cas_n <= 1'd1;
		main_sdram_inti_p0_ras_n <= 1'd1;
	end
end
assign main_sdram_inti_p0_address = main_sdram_phaseinjector0_address_storage;
assign main_sdram_inti_p0_bank = main_sdram_phaseinjector0_baddress_storage;
assign main_sdram_inti_p0_wrdata_en = (main_sdram_phaseinjector0_command_issue_re & main_sdram_phaseinjector0_command_storage[4]);
assign main_sdram_inti_p0_rddata_en = (main_sdram_phaseinjector0_command_issue_re & main_sdram_phaseinjector0_command_storage[5]);
assign main_sdram_inti_p0_wrdata = main_sdram_phaseinjector0_wrdata_storage;
assign main_sdram_inti_p0_wrdata_mask = 1'd0;
always @(*) begin
	main_sdram_inti_p1_cs_n <= 1'd1;
	main_sdram_inti_p1_ras_n <= 1'd1;
	main_sdram_inti_p1_we_n <= 1'd1;
	main_sdram_inti_p1_cas_n <= 1'd1;
	if (main_sdram_phaseinjector1_command_issue_re) begin
		main_sdram_inti_p1_cs_n <= {1{(~main_sdram_phaseinjector1_command_storage[0])}};
		main_sdram_inti_p1_we_n <= (~main_sdram_phaseinjector1_command_storage[1]);
		main_sdram_inti_p1_cas_n <= (~main_sdram_phaseinjector1_command_storage[2]);
		main_sdram_inti_p1_ras_n <= (~main_sdram_phaseinjector1_command_storage[3]);
	end else begin
		main_sdram_inti_p1_cs_n <= {1{1'd1}};
		main_sdram_inti_p1_we_n <= 1'd1;
		main_sdram_inti_p1_cas_n <= 1'd1;
		main_sdram_inti_p1_ras_n <= 1'd1;
	end
end
assign main_sdram_inti_p1_address = main_sdram_phaseinjector1_address_storage;
assign main_sdram_inti_p1_bank = main_sdram_phaseinjector1_baddress_storage;
assign main_sdram_inti_p1_wrdata_en = (main_sdram_phaseinjector1_command_issue_re & main_sdram_phaseinjector1_command_storage[4]);
assign main_sdram_inti_p1_rddata_en = (main_sdram_phaseinjector1_command_issue_re & main_sdram_phaseinjector1_command_storage[5]);
assign main_sdram_inti_p1_wrdata = main_sdram_phaseinjector1_wrdata_storage;
assign main_sdram_inti_p1_wrdata_mask = 1'd0;
always @(*) begin
	main_sdram_inti_p2_cs_n <= 1'd1;
	main_sdram_inti_p2_ras_n <= 1'd1;
	main_sdram_inti_p2_we_n <= 1'd1;
	main_sdram_inti_p2_cas_n <= 1'd1;
	if (main_sdram_phaseinjector2_command_issue_re) begin
		main_sdram_inti_p2_cs_n <= {1{(~main_sdram_phaseinjector2_command_storage[0])}};
		main_sdram_inti_p2_we_n <= (~main_sdram_phaseinjector2_command_storage[1]);
		main_sdram_inti_p2_cas_n <= (~main_sdram_phaseinjector2_command_storage[2]);
		main_sdram_inti_p2_ras_n <= (~main_sdram_phaseinjector2_command_storage[3]);
	end else begin
		main_sdram_inti_p2_cs_n <= {1{1'd1}};
		main_sdram_inti_p2_we_n <= 1'd1;
		main_sdram_inti_p2_cas_n <= 1'd1;
		main_sdram_inti_p2_ras_n <= 1'd1;
	end
end
assign main_sdram_inti_p2_address = main_sdram_phaseinjector2_address_storage;
assign main_sdram_inti_p2_bank = main_sdram_phaseinjector2_baddress_storage;
assign main_sdram_inti_p2_wrdata_en = (main_sdram_phaseinjector2_command_issue_re & main_sdram_phaseinjector2_command_storage[4]);
assign main_sdram_inti_p2_rddata_en = (main_sdram_phaseinjector2_command_issue_re & main_sdram_phaseinjector2_command_storage[5]);
assign main_sdram_inti_p2_wrdata = main_sdram_phaseinjector2_wrdata_storage;
assign main_sdram_inti_p2_wrdata_mask = 1'd0;
always @(*) begin
	main_sdram_inti_p3_cs_n <= 1'd1;
	main_sdram_inti_p3_ras_n <= 1'd1;
	main_sdram_inti_p3_we_n <= 1'd1;
	main_sdram_inti_p3_cas_n <= 1'd1;
	if (main_sdram_phaseinjector3_command_issue_re) begin
		main_sdram_inti_p3_cs_n <= {1{(~main_sdram_phaseinjector3_command_storage[0])}};
		main_sdram_inti_p3_we_n <= (~main_sdram_phaseinjector3_command_storage[1]);
		main_sdram_inti_p3_cas_n <= (~main_sdram_phaseinjector3_command_storage[2]);
		main_sdram_inti_p3_ras_n <= (~main_sdram_phaseinjector3_command_storage[3]);
	end else begin
		main_sdram_inti_p3_cs_n <= {1{1'd1}};
		main_sdram_inti_p3_we_n <= 1'd1;
		main_sdram_inti_p3_cas_n <= 1'd1;
		main_sdram_inti_p3_ras_n <= 1'd1;
	end
end
assign main_sdram_inti_p3_address = main_sdram_phaseinjector3_address_storage;
assign main_sdram_inti_p3_bank = main_sdram_phaseinjector3_baddress_storage;
assign main_sdram_inti_p3_wrdata_en = (main_sdram_phaseinjector3_command_issue_re & main_sdram_phaseinjector3_command_storage[4]);
assign main_sdram_inti_p3_rddata_en = (main_sdram_phaseinjector3_command_issue_re & main_sdram_phaseinjector3_command_storage[5]);
assign main_sdram_inti_p3_wrdata = main_sdram_phaseinjector3_wrdata_storage;
assign main_sdram_inti_p3_wrdata_mask = 1'd0;
assign main_sdram_bankmachine0_req_valid = main_sdram_interface_bank0_valid;
assign main_sdram_interface_bank0_ready = main_sdram_bankmachine0_req_ready;
assign main_sdram_bankmachine0_req_we = main_sdram_interface_bank0_we;
assign main_sdram_bankmachine0_req_addr = main_sdram_interface_bank0_addr;
assign main_sdram_interface_bank0_lock = main_sdram_bankmachine0_req_lock;
assign main_sdram_interface_bank0_wdata_ready = main_sdram_bankmachine0_req_wdata_ready;
assign main_sdram_interface_bank0_rdata_valid = main_sdram_bankmachine0_req_rdata_valid;
assign main_sdram_bankmachine1_req_valid = main_sdram_interface_bank1_valid;
assign main_sdram_interface_bank1_ready = main_sdram_bankmachine1_req_ready;
assign main_sdram_bankmachine1_req_we = main_sdram_interface_bank1_we;
assign main_sdram_bankmachine1_req_addr = main_sdram_interface_bank1_addr;
assign main_sdram_interface_bank1_lock = main_sdram_bankmachine1_req_lock;
assign main_sdram_interface_bank1_wdata_ready = main_sdram_bankmachine1_req_wdata_ready;
assign main_sdram_interface_bank1_rdata_valid = main_sdram_bankmachine1_req_rdata_valid;
assign main_sdram_bankmachine2_req_valid = main_sdram_interface_bank2_valid;
assign main_sdram_interface_bank2_ready = main_sdram_bankmachine2_req_ready;
assign main_sdram_bankmachine2_req_we = main_sdram_interface_bank2_we;
assign main_sdram_bankmachine2_req_addr = main_sdram_interface_bank2_addr;
assign main_sdram_interface_bank2_lock = main_sdram_bankmachine2_req_lock;
assign main_sdram_interface_bank2_wdata_ready = main_sdram_bankmachine2_req_wdata_ready;
assign main_sdram_interface_bank2_rdata_valid = main_sdram_bankmachine2_req_rdata_valid;
assign main_sdram_bankmachine3_req_valid = main_sdram_interface_bank3_valid;
assign main_sdram_interface_bank3_ready = main_sdram_bankmachine3_req_ready;
assign main_sdram_bankmachine3_req_we = main_sdram_interface_bank3_we;
assign main_sdram_bankmachine3_req_addr = main_sdram_interface_bank3_addr;
assign main_sdram_interface_bank3_lock = main_sdram_bankmachine3_req_lock;
assign main_sdram_interface_bank3_wdata_ready = main_sdram_bankmachine3_req_wdata_ready;
assign main_sdram_interface_bank3_rdata_valid = main_sdram_bankmachine3_req_rdata_valid;
assign main_sdram_bankmachine4_req_valid = main_sdram_interface_bank4_valid;
assign main_sdram_interface_bank4_ready = main_sdram_bankmachine4_req_ready;
assign main_sdram_bankmachine4_req_we = main_sdram_interface_bank4_we;
assign main_sdram_bankmachine4_req_addr = main_sdram_interface_bank4_addr;
assign main_sdram_interface_bank4_lock = main_sdram_bankmachine4_req_lock;
assign main_sdram_interface_bank4_wdata_ready = main_sdram_bankmachine4_req_wdata_ready;
assign main_sdram_interface_bank4_rdata_valid = main_sdram_bankmachine4_req_rdata_valid;
assign main_sdram_bankmachine5_req_valid = main_sdram_interface_bank5_valid;
assign main_sdram_interface_bank5_ready = main_sdram_bankmachine5_req_ready;
assign main_sdram_bankmachine5_req_we = main_sdram_interface_bank5_we;
assign main_sdram_bankmachine5_req_addr = main_sdram_interface_bank5_addr;
assign main_sdram_interface_bank5_lock = main_sdram_bankmachine5_req_lock;
assign main_sdram_interface_bank5_wdata_ready = main_sdram_bankmachine5_req_wdata_ready;
assign main_sdram_interface_bank5_rdata_valid = main_sdram_bankmachine5_req_rdata_valid;
assign main_sdram_bankmachine6_req_valid = main_sdram_interface_bank6_valid;
assign main_sdram_interface_bank6_ready = main_sdram_bankmachine6_req_ready;
assign main_sdram_bankmachine6_req_we = main_sdram_interface_bank6_we;
assign main_sdram_bankmachine6_req_addr = main_sdram_interface_bank6_addr;
assign main_sdram_interface_bank6_lock = main_sdram_bankmachine6_req_lock;
assign main_sdram_interface_bank6_wdata_ready = main_sdram_bankmachine6_req_wdata_ready;
assign main_sdram_interface_bank6_rdata_valid = main_sdram_bankmachine6_req_rdata_valid;
assign main_sdram_bankmachine7_req_valid = main_sdram_interface_bank7_valid;
assign main_sdram_interface_bank7_ready = main_sdram_bankmachine7_req_ready;
assign main_sdram_bankmachine7_req_we = main_sdram_interface_bank7_we;
assign main_sdram_bankmachine7_req_addr = main_sdram_interface_bank7_addr;
assign main_sdram_interface_bank7_lock = main_sdram_bankmachine7_req_lock;
assign main_sdram_interface_bank7_wdata_ready = main_sdram_bankmachine7_req_wdata_ready;
assign main_sdram_interface_bank7_rdata_valid = main_sdram_bankmachine7_req_rdata_valid;
assign main_sdram_timer_wait = (~main_sdram_timer_done0);
assign main_sdram_postponer_req_i = main_sdram_timer_done0;
assign main_sdram_wants_refresh = main_sdram_postponer_req_o;
assign main_sdram_wants_zqcs = main_sdram_zqcs_timer_done0;
assign main_sdram_zqcs_timer_wait = (~main_sdram_zqcs_executer_done);
assign main_sdram_timer_done1 = (main_sdram_timer_count1 == 1'd0);
assign main_sdram_timer_done0 = main_sdram_timer_done1;
assign main_sdram_timer_count0 = main_sdram_timer_count1;
assign main_sdram_sequencer_start1 = (main_sdram_sequencer_start0 | (main_sdram_sequencer_count != 1'd0));
assign main_sdram_sequencer_done0 = (main_sdram_sequencer_done1 & (main_sdram_sequencer_count == 1'd0));
assign main_sdram_zqcs_timer_done1 = (main_sdram_zqcs_timer_count1 == 1'd0);
assign main_sdram_zqcs_timer_done0 = main_sdram_zqcs_timer_done1;
assign main_sdram_zqcs_timer_count0 = main_sdram_zqcs_timer_count1;
always @(*) begin
	main_sdram_zqcs_executer_start <= 1'd0;
	main_sdram_cmd_last <= 1'd0;
	main_sdram_sequencer_start0 <= 1'd0;
	main_sdram_cmd_valid <= 1'd0;
	builder_refresher_next_state <= 2'd0;
	builder_refresher_next_state <= builder_refresher_state;
	case (builder_refresher_state)
		1'd1: begin
			main_sdram_cmd_valid <= 1'd1;
			if (main_sdram_cmd_ready) begin
				main_sdram_sequencer_start0 <= 1'd1;
				builder_refresher_next_state <= 2'd2;
			end
		end
		2'd2: begin
			main_sdram_cmd_valid <= 1'd1;
			if (main_sdram_sequencer_done0) begin
				if (main_sdram_wants_zqcs) begin
					main_sdram_zqcs_executer_start <= 1'd1;
					builder_refresher_next_state <= 2'd3;
				end else begin
					main_sdram_cmd_valid <= 1'd0;
					main_sdram_cmd_last <= 1'd1;
					builder_refresher_next_state <= 1'd0;
				end
			end
		end
		2'd3: begin
			main_sdram_cmd_valid <= 1'd1;
			if (main_sdram_zqcs_executer_done) begin
				main_sdram_cmd_valid <= 1'd0;
				main_sdram_cmd_last <= 1'd1;
				builder_refresher_next_state <= 1'd0;
			end
		end
		default: begin
			if (1'd1) begin
				if (main_sdram_wants_refresh) begin
					builder_refresher_next_state <= 1'd1;
				end
			end
		end
	endcase
end
assign main_sdram_bankmachine0_cmd_buffer_lookahead_sink_valid = main_sdram_bankmachine0_req_valid;
assign main_sdram_bankmachine0_req_ready = main_sdram_bankmachine0_cmd_buffer_lookahead_sink_ready;
assign main_sdram_bankmachine0_cmd_buffer_lookahead_sink_payload_we = main_sdram_bankmachine0_req_we;
assign main_sdram_bankmachine0_cmd_buffer_lookahead_sink_payload_addr = main_sdram_bankmachine0_req_addr;
assign main_sdram_bankmachine0_cmd_buffer_sink_valid = main_sdram_bankmachine0_cmd_buffer_lookahead_source_valid;
assign main_sdram_bankmachine0_cmd_buffer_lookahead_source_ready = main_sdram_bankmachine0_cmd_buffer_sink_ready;
assign main_sdram_bankmachine0_cmd_buffer_sink_first = main_sdram_bankmachine0_cmd_buffer_lookahead_source_first;
assign main_sdram_bankmachine0_cmd_buffer_sink_last = main_sdram_bankmachine0_cmd_buffer_lookahead_source_last;
assign main_sdram_bankmachine0_cmd_buffer_sink_payload_we = main_sdram_bankmachine0_cmd_buffer_lookahead_source_payload_we;
assign main_sdram_bankmachine0_cmd_buffer_sink_payload_addr = main_sdram_bankmachine0_cmd_buffer_lookahead_source_payload_addr;
assign main_sdram_bankmachine0_cmd_buffer_source_ready = (main_sdram_bankmachine0_req_wdata_ready | main_sdram_bankmachine0_req_rdata_valid);
assign main_sdram_bankmachine0_req_lock = (main_sdram_bankmachine0_cmd_buffer_lookahead_source_valid | main_sdram_bankmachine0_cmd_buffer_source_valid);
assign main_sdram_bankmachine0_row_hit = (main_sdram_bankmachine0_row == main_sdram_bankmachine0_cmd_buffer_source_payload_addr[20:7]);
assign main_sdram_bankmachine0_cmd_payload_ba = 1'd0;
always @(*) begin
	main_sdram_bankmachine0_cmd_payload_a <= 14'd0;
	if (main_sdram_bankmachine0_row_col_n_addr_sel) begin
		main_sdram_bankmachine0_cmd_payload_a <= main_sdram_bankmachine0_cmd_buffer_source_payload_addr[20:7];
	end else begin
		main_sdram_bankmachine0_cmd_payload_a <= ((main_sdram_bankmachine0_auto_precharge <<< 4'd10) | {main_sdram_bankmachine0_cmd_buffer_source_payload_addr[6:0], {3{1'd0}}});
	end
end
assign main_sdram_bankmachine0_twtpcon_valid = ((main_sdram_bankmachine0_cmd_valid & main_sdram_bankmachine0_cmd_ready) & main_sdram_bankmachine0_cmd_payload_is_write);
assign main_sdram_bankmachine0_trccon_valid = ((main_sdram_bankmachine0_cmd_valid & main_sdram_bankmachine0_cmd_ready) & main_sdram_bankmachine0_row_open);
assign main_sdram_bankmachine0_trascon_valid = ((main_sdram_bankmachine0_cmd_valid & main_sdram_bankmachine0_cmd_ready) & main_sdram_bankmachine0_row_open);
always @(*) begin
	main_sdram_bankmachine0_auto_precharge <= 1'd0;
	if ((main_sdram_bankmachine0_cmd_buffer_lookahead_source_valid & main_sdram_bankmachine0_cmd_buffer_source_valid)) begin
		if ((main_sdram_bankmachine0_cmd_buffer_lookahead_source_payload_addr[20:7] != main_sdram_bankmachine0_cmd_buffer_source_payload_addr[20:7])) begin
			main_sdram_bankmachine0_auto_precharge <= (main_sdram_bankmachine0_row_close == 1'd0);
		end
	end
end
assign main_sdram_bankmachine0_cmd_buffer_lookahead_syncfifo0_din = {main_sdram_bankmachine0_cmd_buffer_lookahead_fifo_in_last, main_sdram_bankmachine0_cmd_buffer_lookahead_fifo_in_first, main_sdram_bankmachine0_cmd_buffer_lookahead_fifo_in_payload_addr, main_sdram_bankmachine0_cmd_buffer_lookahead_fifo_in_payload_we};
assign {main_sdram_bankmachine0_cmd_buffer_lookahead_fifo_out_last, main_sdram_bankmachine0_cmd_buffer_lookahead_fifo_out_first, main_sdram_bankmachine0_cmd_buffer_lookahead_fifo_out_payload_addr, main_sdram_bankmachine0_cmd_buffer_lookahead_fifo_out_payload_we} = main_sdram_bankmachine0_cmd_buffer_lookahead_syncfifo0_dout;
assign main_sdram_bankmachine0_cmd_buffer_lookahead_sink_ready = main_sdram_bankmachine0_cmd_buffer_lookahead_syncfifo0_writable;
assign main_sdram_bankmachine0_cmd_buffer_lookahead_syncfifo0_we = main_sdram_bankmachine0_cmd_buffer_lookahead_sink_valid;
assign main_sdram_bankmachine0_cmd_buffer_lookahead_fifo_in_first = main_sdram_bankmachine0_cmd_buffer_lookahead_sink_first;
assign main_sdram_bankmachine0_cmd_buffer_lookahead_fifo_in_last = main_sdram_bankmachine0_cmd_buffer_lookahead_sink_last;
assign main_sdram_bankmachine0_cmd_buffer_lookahead_fifo_in_payload_we = main_sdram_bankmachine0_cmd_buffer_lookahead_sink_payload_we;
assign main_sdram_bankmachine0_cmd_buffer_lookahead_fifo_in_payload_addr = main_sdram_bankmachine0_cmd_buffer_lookahead_sink_payload_addr;
assign main_sdram_bankmachine0_cmd_buffer_lookahead_source_valid = main_sdram_bankmachine0_cmd_buffer_lookahead_syncfifo0_readable;
assign main_sdram_bankmachine0_cmd_buffer_lookahead_source_first = main_sdram_bankmachine0_cmd_buffer_lookahead_fifo_out_first;
assign main_sdram_bankmachine0_cmd_buffer_lookahead_source_last = main_sdram_bankmachine0_cmd_buffer_lookahead_fifo_out_last;
assign main_sdram_bankmachine0_cmd_buffer_lookahead_source_payload_we = main_sdram_bankmachine0_cmd_buffer_lookahead_fifo_out_payload_we;
assign main_sdram_bankmachine0_cmd_buffer_lookahead_source_payload_addr = main_sdram_bankmachine0_cmd_buffer_lookahead_fifo_out_payload_addr;
assign main_sdram_bankmachine0_cmd_buffer_lookahead_syncfifo0_re = main_sdram_bankmachine0_cmd_buffer_lookahead_source_ready;
always @(*) begin
	main_sdram_bankmachine0_cmd_buffer_lookahead_wrport_adr <= 3'd0;
	if (main_sdram_bankmachine0_cmd_buffer_lookahead_replace) begin
		main_sdram_bankmachine0_cmd_buffer_lookahead_wrport_adr <= (main_sdram_bankmachine0_cmd_buffer_lookahead_produce - 1'd1);
	end else begin
		main_sdram_bankmachine0_cmd_buffer_lookahead_wrport_adr <= main_sdram_bankmachine0_cmd_buffer_lookahead_produce;
	end
end
assign main_sdram_bankmachine0_cmd_buffer_lookahead_wrport_dat_w = main_sdram_bankmachine0_cmd_buffer_lookahead_syncfifo0_din;
assign main_sdram_bankmachine0_cmd_buffer_lookahead_wrport_we = (main_sdram_bankmachine0_cmd_buffer_lookahead_syncfifo0_we & (main_sdram_bankmachine0_cmd_buffer_lookahead_syncfifo0_writable | main_sdram_bankmachine0_cmd_buffer_lookahead_replace));
assign main_sdram_bankmachine0_cmd_buffer_lookahead_do_read = (main_sdram_bankmachine0_cmd_buffer_lookahead_syncfifo0_readable & main_sdram_bankmachine0_cmd_buffer_lookahead_syncfifo0_re);
assign main_sdram_bankmachine0_cmd_buffer_lookahead_rdport_adr = main_sdram_bankmachine0_cmd_buffer_lookahead_consume;
assign main_sdram_bankmachine0_cmd_buffer_lookahead_syncfifo0_dout = main_sdram_bankmachine0_cmd_buffer_lookahead_rdport_dat_r;
assign main_sdram_bankmachine0_cmd_buffer_lookahead_syncfifo0_writable = (main_sdram_bankmachine0_cmd_buffer_lookahead_level != 4'd8);
assign main_sdram_bankmachine0_cmd_buffer_lookahead_syncfifo0_readable = (main_sdram_bankmachine0_cmd_buffer_lookahead_level != 1'd0);
assign main_sdram_bankmachine0_cmd_buffer_sink_ready = ((~main_sdram_bankmachine0_cmd_buffer_source_valid) | main_sdram_bankmachine0_cmd_buffer_source_ready);
always @(*) begin
	main_sdram_bankmachine0_cmd_payload_cas <= 1'd0;
	main_sdram_bankmachine0_cmd_payload_ras <= 1'd0;
	main_sdram_bankmachine0_cmd_payload_we <= 1'd0;
	main_sdram_bankmachine0_row_col_n_addr_sel <= 1'd0;
	main_sdram_bankmachine0_cmd_payload_is_cmd <= 1'd0;
	main_sdram_bankmachine0_cmd_payload_is_read <= 1'd0;
	main_sdram_bankmachine0_cmd_payload_is_write <= 1'd0;
	main_sdram_bankmachine0_req_wdata_ready <= 1'd0;
	builder_bankmachine0_next_state <= 3'd0;
	main_sdram_bankmachine0_req_rdata_valid <= 1'd0;
	main_sdram_bankmachine0_refresh_gnt <= 1'd0;
	main_sdram_bankmachine0_cmd_valid <= 1'd0;
	main_sdram_bankmachine0_row_open <= 1'd0;
	main_sdram_bankmachine0_row_close <= 1'd0;
	builder_bankmachine0_next_state <= builder_bankmachine0_state;
	case (builder_bankmachine0_state)
		1'd1: begin
			if ((main_sdram_bankmachine0_twtpcon_ready & main_sdram_bankmachine0_trascon_ready)) begin
				main_sdram_bankmachine0_cmd_valid <= 1'd1;
				if (main_sdram_bankmachine0_cmd_ready) begin
					builder_bankmachine0_next_state <= 3'd5;
				end
				main_sdram_bankmachine0_cmd_payload_ras <= 1'd1;
				main_sdram_bankmachine0_cmd_payload_we <= 1'd1;
				main_sdram_bankmachine0_cmd_payload_is_cmd <= 1'd1;
			end
			main_sdram_bankmachine0_row_close <= 1'd1;
		end
		2'd2: begin
			if ((main_sdram_bankmachine0_twtpcon_ready & main_sdram_bankmachine0_trascon_ready)) begin
				builder_bankmachine0_next_state <= 3'd5;
			end
			main_sdram_bankmachine0_row_close <= 1'd1;
		end
		2'd3: begin
			if (main_sdram_bankmachine0_trccon_ready) begin
				main_sdram_bankmachine0_row_col_n_addr_sel <= 1'd1;
				main_sdram_bankmachine0_row_open <= 1'd1;
				main_sdram_bankmachine0_cmd_valid <= 1'd1;
				main_sdram_bankmachine0_cmd_payload_is_cmd <= 1'd1;
				if (main_sdram_bankmachine0_cmd_ready) begin
					builder_bankmachine0_next_state <= 3'd6;
				end
				main_sdram_bankmachine0_cmd_payload_ras <= 1'd1;
			end
		end
		3'd4: begin
			if (main_sdram_bankmachine0_twtpcon_ready) begin
				main_sdram_bankmachine0_refresh_gnt <= 1'd1;
			end
			main_sdram_bankmachine0_row_close <= 1'd1;
			main_sdram_bankmachine0_cmd_payload_is_cmd <= 1'd1;
			if ((~main_sdram_bankmachine0_refresh_req)) begin
				builder_bankmachine0_next_state <= 1'd0;
			end
		end
		3'd5: begin
			builder_bankmachine0_next_state <= 2'd3;
		end
		3'd6: begin
			builder_bankmachine0_next_state <= 1'd0;
		end
		default: begin
			if (main_sdram_bankmachine0_refresh_req) begin
				builder_bankmachine0_next_state <= 3'd4;
			end else begin
				if (main_sdram_bankmachine0_cmd_buffer_source_valid) begin
					if (main_sdram_bankmachine0_row_opened) begin
						if (main_sdram_bankmachine0_row_hit) begin
							main_sdram_bankmachine0_cmd_valid <= 1'd1;
							if (main_sdram_bankmachine0_cmd_buffer_source_payload_we) begin
								main_sdram_bankmachine0_req_wdata_ready <= main_sdram_bankmachine0_cmd_ready;
								main_sdram_bankmachine0_cmd_payload_is_write <= 1'd1;
								main_sdram_bankmachine0_cmd_payload_we <= 1'd1;
							end else begin
								main_sdram_bankmachine0_req_rdata_valid <= main_sdram_bankmachine0_cmd_ready;
								main_sdram_bankmachine0_cmd_payload_is_read <= 1'd1;
							end
							main_sdram_bankmachine0_cmd_payload_cas <= 1'd1;
							if ((main_sdram_bankmachine0_cmd_ready & main_sdram_bankmachine0_auto_precharge)) begin
								builder_bankmachine0_next_state <= 2'd2;
							end
						end else begin
							builder_bankmachine0_next_state <= 1'd1;
						end
					end else begin
						builder_bankmachine0_next_state <= 2'd3;
					end
				end
			end
		end
	endcase
end
assign main_sdram_bankmachine1_cmd_buffer_lookahead_sink_valid = main_sdram_bankmachine1_req_valid;
assign main_sdram_bankmachine1_req_ready = main_sdram_bankmachine1_cmd_buffer_lookahead_sink_ready;
assign main_sdram_bankmachine1_cmd_buffer_lookahead_sink_payload_we = main_sdram_bankmachine1_req_we;
assign main_sdram_bankmachine1_cmd_buffer_lookahead_sink_payload_addr = main_sdram_bankmachine1_req_addr;
assign main_sdram_bankmachine1_cmd_buffer_sink_valid = main_sdram_bankmachine1_cmd_buffer_lookahead_source_valid;
assign main_sdram_bankmachine1_cmd_buffer_lookahead_source_ready = main_sdram_bankmachine1_cmd_buffer_sink_ready;
assign main_sdram_bankmachine1_cmd_buffer_sink_first = main_sdram_bankmachine1_cmd_buffer_lookahead_source_first;
assign main_sdram_bankmachine1_cmd_buffer_sink_last = main_sdram_bankmachine1_cmd_buffer_lookahead_source_last;
assign main_sdram_bankmachine1_cmd_buffer_sink_payload_we = main_sdram_bankmachine1_cmd_buffer_lookahead_source_payload_we;
assign main_sdram_bankmachine1_cmd_buffer_sink_payload_addr = main_sdram_bankmachine1_cmd_buffer_lookahead_source_payload_addr;
assign main_sdram_bankmachine1_cmd_buffer_source_ready = (main_sdram_bankmachine1_req_wdata_ready | main_sdram_bankmachine1_req_rdata_valid);
assign main_sdram_bankmachine1_req_lock = (main_sdram_bankmachine1_cmd_buffer_lookahead_source_valid | main_sdram_bankmachine1_cmd_buffer_source_valid);
assign main_sdram_bankmachine1_row_hit = (main_sdram_bankmachine1_row == main_sdram_bankmachine1_cmd_buffer_source_payload_addr[20:7]);
assign main_sdram_bankmachine1_cmd_payload_ba = 1'd1;
always @(*) begin
	main_sdram_bankmachine1_cmd_payload_a <= 14'd0;
	if (main_sdram_bankmachine1_row_col_n_addr_sel) begin
		main_sdram_bankmachine1_cmd_payload_a <= main_sdram_bankmachine1_cmd_buffer_source_payload_addr[20:7];
	end else begin
		main_sdram_bankmachine1_cmd_payload_a <= ((main_sdram_bankmachine1_auto_precharge <<< 4'd10) | {main_sdram_bankmachine1_cmd_buffer_source_payload_addr[6:0], {3{1'd0}}});
	end
end
assign main_sdram_bankmachine1_twtpcon_valid = ((main_sdram_bankmachine1_cmd_valid & main_sdram_bankmachine1_cmd_ready) & main_sdram_bankmachine1_cmd_payload_is_write);
assign main_sdram_bankmachine1_trccon_valid = ((main_sdram_bankmachine1_cmd_valid & main_sdram_bankmachine1_cmd_ready) & main_sdram_bankmachine1_row_open);
assign main_sdram_bankmachine1_trascon_valid = ((main_sdram_bankmachine1_cmd_valid & main_sdram_bankmachine1_cmd_ready) & main_sdram_bankmachine1_row_open);
always @(*) begin
	main_sdram_bankmachine1_auto_precharge <= 1'd0;
	if ((main_sdram_bankmachine1_cmd_buffer_lookahead_source_valid & main_sdram_bankmachine1_cmd_buffer_source_valid)) begin
		if ((main_sdram_bankmachine1_cmd_buffer_lookahead_source_payload_addr[20:7] != main_sdram_bankmachine1_cmd_buffer_source_payload_addr[20:7])) begin
			main_sdram_bankmachine1_auto_precharge <= (main_sdram_bankmachine1_row_close == 1'd0);
		end
	end
end
assign main_sdram_bankmachine1_cmd_buffer_lookahead_syncfifo1_din = {main_sdram_bankmachine1_cmd_buffer_lookahead_fifo_in_last, main_sdram_bankmachine1_cmd_buffer_lookahead_fifo_in_first, main_sdram_bankmachine1_cmd_buffer_lookahead_fifo_in_payload_addr, main_sdram_bankmachine1_cmd_buffer_lookahead_fifo_in_payload_we};
assign {main_sdram_bankmachine1_cmd_buffer_lookahead_fifo_out_last, main_sdram_bankmachine1_cmd_buffer_lookahead_fifo_out_first, main_sdram_bankmachine1_cmd_buffer_lookahead_fifo_out_payload_addr, main_sdram_bankmachine1_cmd_buffer_lookahead_fifo_out_payload_we} = main_sdram_bankmachine1_cmd_buffer_lookahead_syncfifo1_dout;
assign main_sdram_bankmachine1_cmd_buffer_lookahead_sink_ready = main_sdram_bankmachine1_cmd_buffer_lookahead_syncfifo1_writable;
assign main_sdram_bankmachine1_cmd_buffer_lookahead_syncfifo1_we = main_sdram_bankmachine1_cmd_buffer_lookahead_sink_valid;
assign main_sdram_bankmachine1_cmd_buffer_lookahead_fifo_in_first = main_sdram_bankmachine1_cmd_buffer_lookahead_sink_first;
assign main_sdram_bankmachine1_cmd_buffer_lookahead_fifo_in_last = main_sdram_bankmachine1_cmd_buffer_lookahead_sink_last;
assign main_sdram_bankmachine1_cmd_buffer_lookahead_fifo_in_payload_we = main_sdram_bankmachine1_cmd_buffer_lookahead_sink_payload_we;
assign main_sdram_bankmachine1_cmd_buffer_lookahead_fifo_in_payload_addr = main_sdram_bankmachine1_cmd_buffer_lookahead_sink_payload_addr;
assign main_sdram_bankmachine1_cmd_buffer_lookahead_source_valid = main_sdram_bankmachine1_cmd_buffer_lookahead_syncfifo1_readable;
assign main_sdram_bankmachine1_cmd_buffer_lookahead_source_first = main_sdram_bankmachine1_cmd_buffer_lookahead_fifo_out_first;
assign main_sdram_bankmachine1_cmd_buffer_lookahead_source_last = main_sdram_bankmachine1_cmd_buffer_lookahead_fifo_out_last;
assign main_sdram_bankmachine1_cmd_buffer_lookahead_source_payload_we = main_sdram_bankmachine1_cmd_buffer_lookahead_fifo_out_payload_we;
assign main_sdram_bankmachine1_cmd_buffer_lookahead_source_payload_addr = main_sdram_bankmachine1_cmd_buffer_lookahead_fifo_out_payload_addr;
assign main_sdram_bankmachine1_cmd_buffer_lookahead_syncfifo1_re = main_sdram_bankmachine1_cmd_buffer_lookahead_source_ready;
always @(*) begin
	main_sdram_bankmachine1_cmd_buffer_lookahead_wrport_adr <= 3'd0;
	if (main_sdram_bankmachine1_cmd_buffer_lookahead_replace) begin
		main_sdram_bankmachine1_cmd_buffer_lookahead_wrport_adr <= (main_sdram_bankmachine1_cmd_buffer_lookahead_produce - 1'd1);
	end else begin
		main_sdram_bankmachine1_cmd_buffer_lookahead_wrport_adr <= main_sdram_bankmachine1_cmd_buffer_lookahead_produce;
	end
end
assign main_sdram_bankmachine1_cmd_buffer_lookahead_wrport_dat_w = main_sdram_bankmachine1_cmd_buffer_lookahead_syncfifo1_din;
assign main_sdram_bankmachine1_cmd_buffer_lookahead_wrport_we = (main_sdram_bankmachine1_cmd_buffer_lookahead_syncfifo1_we & (main_sdram_bankmachine1_cmd_buffer_lookahead_syncfifo1_writable | main_sdram_bankmachine1_cmd_buffer_lookahead_replace));
assign main_sdram_bankmachine1_cmd_buffer_lookahead_do_read = (main_sdram_bankmachine1_cmd_buffer_lookahead_syncfifo1_readable & main_sdram_bankmachine1_cmd_buffer_lookahead_syncfifo1_re);
assign main_sdram_bankmachine1_cmd_buffer_lookahead_rdport_adr = main_sdram_bankmachine1_cmd_buffer_lookahead_consume;
assign main_sdram_bankmachine1_cmd_buffer_lookahead_syncfifo1_dout = main_sdram_bankmachine1_cmd_buffer_lookahead_rdport_dat_r;
assign main_sdram_bankmachine1_cmd_buffer_lookahead_syncfifo1_writable = (main_sdram_bankmachine1_cmd_buffer_lookahead_level != 4'd8);
assign main_sdram_bankmachine1_cmd_buffer_lookahead_syncfifo1_readable = (main_sdram_bankmachine1_cmd_buffer_lookahead_level != 1'd0);
assign main_sdram_bankmachine1_cmd_buffer_sink_ready = ((~main_sdram_bankmachine1_cmd_buffer_source_valid) | main_sdram_bankmachine1_cmd_buffer_source_ready);
always @(*) begin
	main_sdram_bankmachine1_cmd_payload_cas <= 1'd0;
	main_sdram_bankmachine1_cmd_payload_ras <= 1'd0;
	main_sdram_bankmachine1_cmd_payload_we <= 1'd0;
	main_sdram_bankmachine1_row_col_n_addr_sel <= 1'd0;
	main_sdram_bankmachine1_cmd_payload_is_cmd <= 1'd0;
	main_sdram_bankmachine1_cmd_payload_is_read <= 1'd0;
	builder_bankmachine1_next_state <= 3'd0;
	main_sdram_bankmachine1_cmd_payload_is_write <= 1'd0;
	main_sdram_bankmachine1_req_wdata_ready <= 1'd0;
	main_sdram_bankmachine1_req_rdata_valid <= 1'd0;
	main_sdram_bankmachine1_refresh_gnt <= 1'd0;
	main_sdram_bankmachine1_cmd_valid <= 1'd0;
	main_sdram_bankmachine1_row_open <= 1'd0;
	main_sdram_bankmachine1_row_close <= 1'd0;
	builder_bankmachine1_next_state <= builder_bankmachine1_state;
	case (builder_bankmachine1_state)
		1'd1: begin
			if ((main_sdram_bankmachine1_twtpcon_ready & main_sdram_bankmachine1_trascon_ready)) begin
				main_sdram_bankmachine1_cmd_valid <= 1'd1;
				if (main_sdram_bankmachine1_cmd_ready) begin
					builder_bankmachine1_next_state <= 3'd5;
				end
				main_sdram_bankmachine1_cmd_payload_ras <= 1'd1;
				main_sdram_bankmachine1_cmd_payload_we <= 1'd1;
				main_sdram_bankmachine1_cmd_payload_is_cmd <= 1'd1;
			end
			main_sdram_bankmachine1_row_close <= 1'd1;
		end
		2'd2: begin
			if ((main_sdram_bankmachine1_twtpcon_ready & main_sdram_bankmachine1_trascon_ready)) begin
				builder_bankmachine1_next_state <= 3'd5;
			end
			main_sdram_bankmachine1_row_close <= 1'd1;
		end
		2'd3: begin
			if (main_sdram_bankmachine1_trccon_ready) begin
				main_sdram_bankmachine1_row_col_n_addr_sel <= 1'd1;
				main_sdram_bankmachine1_row_open <= 1'd1;
				main_sdram_bankmachine1_cmd_valid <= 1'd1;
				main_sdram_bankmachine1_cmd_payload_is_cmd <= 1'd1;
				if (main_sdram_bankmachine1_cmd_ready) begin
					builder_bankmachine1_next_state <= 3'd6;
				end
				main_sdram_bankmachine1_cmd_payload_ras <= 1'd1;
			end
		end
		3'd4: begin
			if (main_sdram_bankmachine1_twtpcon_ready) begin
				main_sdram_bankmachine1_refresh_gnt <= 1'd1;
			end
			main_sdram_bankmachine1_row_close <= 1'd1;
			main_sdram_bankmachine1_cmd_payload_is_cmd <= 1'd1;
			if ((~main_sdram_bankmachine1_refresh_req)) begin
				builder_bankmachine1_next_state <= 1'd0;
			end
		end
		3'd5: begin
			builder_bankmachine1_next_state <= 2'd3;
		end
		3'd6: begin
			builder_bankmachine1_next_state <= 1'd0;
		end
		default: begin
			if (main_sdram_bankmachine1_refresh_req) begin
				builder_bankmachine1_next_state <= 3'd4;
			end else begin
				if (main_sdram_bankmachine1_cmd_buffer_source_valid) begin
					if (main_sdram_bankmachine1_row_opened) begin
						if (main_sdram_bankmachine1_row_hit) begin
							main_sdram_bankmachine1_cmd_valid <= 1'd1;
							if (main_sdram_bankmachine1_cmd_buffer_source_payload_we) begin
								main_sdram_bankmachine1_req_wdata_ready <= main_sdram_bankmachine1_cmd_ready;
								main_sdram_bankmachine1_cmd_payload_is_write <= 1'd1;
								main_sdram_bankmachine1_cmd_payload_we <= 1'd1;
							end else begin
								main_sdram_bankmachine1_req_rdata_valid <= main_sdram_bankmachine1_cmd_ready;
								main_sdram_bankmachine1_cmd_payload_is_read <= 1'd1;
							end
							main_sdram_bankmachine1_cmd_payload_cas <= 1'd1;
							if ((main_sdram_bankmachine1_cmd_ready & main_sdram_bankmachine1_auto_precharge)) begin
								builder_bankmachine1_next_state <= 2'd2;
							end
						end else begin
							builder_bankmachine1_next_state <= 1'd1;
						end
					end else begin
						builder_bankmachine1_next_state <= 2'd3;
					end
				end
			end
		end
	endcase
end
assign main_sdram_bankmachine2_cmd_buffer_lookahead_sink_valid = main_sdram_bankmachine2_req_valid;
assign main_sdram_bankmachine2_req_ready = main_sdram_bankmachine2_cmd_buffer_lookahead_sink_ready;
assign main_sdram_bankmachine2_cmd_buffer_lookahead_sink_payload_we = main_sdram_bankmachine2_req_we;
assign main_sdram_bankmachine2_cmd_buffer_lookahead_sink_payload_addr = main_sdram_bankmachine2_req_addr;
assign main_sdram_bankmachine2_cmd_buffer_sink_valid = main_sdram_bankmachine2_cmd_buffer_lookahead_source_valid;
assign main_sdram_bankmachine2_cmd_buffer_lookahead_source_ready = main_sdram_bankmachine2_cmd_buffer_sink_ready;
assign main_sdram_bankmachine2_cmd_buffer_sink_first = main_sdram_bankmachine2_cmd_buffer_lookahead_source_first;
assign main_sdram_bankmachine2_cmd_buffer_sink_last = main_sdram_bankmachine2_cmd_buffer_lookahead_source_last;
assign main_sdram_bankmachine2_cmd_buffer_sink_payload_we = main_sdram_bankmachine2_cmd_buffer_lookahead_source_payload_we;
assign main_sdram_bankmachine2_cmd_buffer_sink_payload_addr = main_sdram_bankmachine2_cmd_buffer_lookahead_source_payload_addr;
assign main_sdram_bankmachine2_cmd_buffer_source_ready = (main_sdram_bankmachine2_req_wdata_ready | main_sdram_bankmachine2_req_rdata_valid);
assign main_sdram_bankmachine2_req_lock = (main_sdram_bankmachine2_cmd_buffer_lookahead_source_valid | main_sdram_bankmachine2_cmd_buffer_source_valid);
assign main_sdram_bankmachine2_row_hit = (main_sdram_bankmachine2_row == main_sdram_bankmachine2_cmd_buffer_source_payload_addr[20:7]);
assign main_sdram_bankmachine2_cmd_payload_ba = 2'd2;
always @(*) begin
	main_sdram_bankmachine2_cmd_payload_a <= 14'd0;
	if (main_sdram_bankmachine2_row_col_n_addr_sel) begin
		main_sdram_bankmachine2_cmd_payload_a <= main_sdram_bankmachine2_cmd_buffer_source_payload_addr[20:7];
	end else begin
		main_sdram_bankmachine2_cmd_payload_a <= ((main_sdram_bankmachine2_auto_precharge <<< 4'd10) | {main_sdram_bankmachine2_cmd_buffer_source_payload_addr[6:0], {3{1'd0}}});
	end
end
assign main_sdram_bankmachine2_twtpcon_valid = ((main_sdram_bankmachine2_cmd_valid & main_sdram_bankmachine2_cmd_ready) & main_sdram_bankmachine2_cmd_payload_is_write);
assign main_sdram_bankmachine2_trccon_valid = ((main_sdram_bankmachine2_cmd_valid & main_sdram_bankmachine2_cmd_ready) & main_sdram_bankmachine2_row_open);
assign main_sdram_bankmachine2_trascon_valid = ((main_sdram_bankmachine2_cmd_valid & main_sdram_bankmachine2_cmd_ready) & main_sdram_bankmachine2_row_open);
always @(*) begin
	main_sdram_bankmachine2_auto_precharge <= 1'd0;
	if ((main_sdram_bankmachine2_cmd_buffer_lookahead_source_valid & main_sdram_bankmachine2_cmd_buffer_source_valid)) begin
		if ((main_sdram_bankmachine2_cmd_buffer_lookahead_source_payload_addr[20:7] != main_sdram_bankmachine2_cmd_buffer_source_payload_addr[20:7])) begin
			main_sdram_bankmachine2_auto_precharge <= (main_sdram_bankmachine2_row_close == 1'd0);
		end
	end
end
assign main_sdram_bankmachine2_cmd_buffer_lookahead_syncfifo2_din = {main_sdram_bankmachine2_cmd_buffer_lookahead_fifo_in_last, main_sdram_bankmachine2_cmd_buffer_lookahead_fifo_in_first, main_sdram_bankmachine2_cmd_buffer_lookahead_fifo_in_payload_addr, main_sdram_bankmachine2_cmd_buffer_lookahead_fifo_in_payload_we};
assign {main_sdram_bankmachine2_cmd_buffer_lookahead_fifo_out_last, main_sdram_bankmachine2_cmd_buffer_lookahead_fifo_out_first, main_sdram_bankmachine2_cmd_buffer_lookahead_fifo_out_payload_addr, main_sdram_bankmachine2_cmd_buffer_lookahead_fifo_out_payload_we} = main_sdram_bankmachine2_cmd_buffer_lookahead_syncfifo2_dout;
assign main_sdram_bankmachine2_cmd_buffer_lookahead_sink_ready = main_sdram_bankmachine2_cmd_buffer_lookahead_syncfifo2_writable;
assign main_sdram_bankmachine2_cmd_buffer_lookahead_syncfifo2_we = main_sdram_bankmachine2_cmd_buffer_lookahead_sink_valid;
assign main_sdram_bankmachine2_cmd_buffer_lookahead_fifo_in_first = main_sdram_bankmachine2_cmd_buffer_lookahead_sink_first;
assign main_sdram_bankmachine2_cmd_buffer_lookahead_fifo_in_last = main_sdram_bankmachine2_cmd_buffer_lookahead_sink_last;
assign main_sdram_bankmachine2_cmd_buffer_lookahead_fifo_in_payload_we = main_sdram_bankmachine2_cmd_buffer_lookahead_sink_payload_we;
assign main_sdram_bankmachine2_cmd_buffer_lookahead_fifo_in_payload_addr = main_sdram_bankmachine2_cmd_buffer_lookahead_sink_payload_addr;
assign main_sdram_bankmachine2_cmd_buffer_lookahead_source_valid = main_sdram_bankmachine2_cmd_buffer_lookahead_syncfifo2_readable;
assign main_sdram_bankmachine2_cmd_buffer_lookahead_source_first = main_sdram_bankmachine2_cmd_buffer_lookahead_fifo_out_first;
assign main_sdram_bankmachine2_cmd_buffer_lookahead_source_last = main_sdram_bankmachine2_cmd_buffer_lookahead_fifo_out_last;
assign main_sdram_bankmachine2_cmd_buffer_lookahead_source_payload_we = main_sdram_bankmachine2_cmd_buffer_lookahead_fifo_out_payload_we;
assign main_sdram_bankmachine2_cmd_buffer_lookahead_source_payload_addr = main_sdram_bankmachine2_cmd_buffer_lookahead_fifo_out_payload_addr;
assign main_sdram_bankmachine2_cmd_buffer_lookahead_syncfifo2_re = main_sdram_bankmachine2_cmd_buffer_lookahead_source_ready;
always @(*) begin
	main_sdram_bankmachine2_cmd_buffer_lookahead_wrport_adr <= 3'd0;
	if (main_sdram_bankmachine2_cmd_buffer_lookahead_replace) begin
		main_sdram_bankmachine2_cmd_buffer_lookahead_wrport_adr <= (main_sdram_bankmachine2_cmd_buffer_lookahead_produce - 1'd1);
	end else begin
		main_sdram_bankmachine2_cmd_buffer_lookahead_wrport_adr <= main_sdram_bankmachine2_cmd_buffer_lookahead_produce;
	end
end
assign main_sdram_bankmachine2_cmd_buffer_lookahead_wrport_dat_w = main_sdram_bankmachine2_cmd_buffer_lookahead_syncfifo2_din;
assign main_sdram_bankmachine2_cmd_buffer_lookahead_wrport_we = (main_sdram_bankmachine2_cmd_buffer_lookahead_syncfifo2_we & (main_sdram_bankmachine2_cmd_buffer_lookahead_syncfifo2_writable | main_sdram_bankmachine2_cmd_buffer_lookahead_replace));
assign main_sdram_bankmachine2_cmd_buffer_lookahead_do_read = (main_sdram_bankmachine2_cmd_buffer_lookahead_syncfifo2_readable & main_sdram_bankmachine2_cmd_buffer_lookahead_syncfifo2_re);
assign main_sdram_bankmachine2_cmd_buffer_lookahead_rdport_adr = main_sdram_bankmachine2_cmd_buffer_lookahead_consume;
assign main_sdram_bankmachine2_cmd_buffer_lookahead_syncfifo2_dout = main_sdram_bankmachine2_cmd_buffer_lookahead_rdport_dat_r;
assign main_sdram_bankmachine2_cmd_buffer_lookahead_syncfifo2_writable = (main_sdram_bankmachine2_cmd_buffer_lookahead_level != 4'd8);
assign main_sdram_bankmachine2_cmd_buffer_lookahead_syncfifo2_readable = (main_sdram_bankmachine2_cmd_buffer_lookahead_level != 1'd0);
assign main_sdram_bankmachine2_cmd_buffer_sink_ready = ((~main_sdram_bankmachine2_cmd_buffer_source_valid) | main_sdram_bankmachine2_cmd_buffer_source_ready);
always @(*) begin
	main_sdram_bankmachine2_cmd_payload_cas <= 1'd0;
	main_sdram_bankmachine2_cmd_payload_ras <= 1'd0;
	main_sdram_bankmachine2_cmd_payload_we <= 1'd0;
	builder_bankmachine2_next_state <= 3'd0;
	main_sdram_bankmachine2_cmd_payload_is_cmd <= 1'd0;
	main_sdram_bankmachine2_row_col_n_addr_sel <= 1'd0;
	main_sdram_bankmachine2_cmd_payload_is_read <= 1'd0;
	main_sdram_bankmachine2_cmd_payload_is_write <= 1'd0;
	main_sdram_bankmachine2_req_wdata_ready <= 1'd0;
	main_sdram_bankmachine2_req_rdata_valid <= 1'd0;
	main_sdram_bankmachine2_refresh_gnt <= 1'd0;
	main_sdram_bankmachine2_cmd_valid <= 1'd0;
	main_sdram_bankmachine2_row_open <= 1'd0;
	main_sdram_bankmachine2_row_close <= 1'd0;
	builder_bankmachine2_next_state <= builder_bankmachine2_state;
	case (builder_bankmachine2_state)
		1'd1: begin
			if ((main_sdram_bankmachine2_twtpcon_ready & main_sdram_bankmachine2_trascon_ready)) begin
				main_sdram_bankmachine2_cmd_valid <= 1'd1;
				if (main_sdram_bankmachine2_cmd_ready) begin
					builder_bankmachine2_next_state <= 3'd5;
				end
				main_sdram_bankmachine2_cmd_payload_ras <= 1'd1;
				main_sdram_bankmachine2_cmd_payload_we <= 1'd1;
				main_sdram_bankmachine2_cmd_payload_is_cmd <= 1'd1;
			end
			main_sdram_bankmachine2_row_close <= 1'd1;
		end
		2'd2: begin
			if ((main_sdram_bankmachine2_twtpcon_ready & main_sdram_bankmachine2_trascon_ready)) begin
				builder_bankmachine2_next_state <= 3'd5;
			end
			main_sdram_bankmachine2_row_close <= 1'd1;
		end
		2'd3: begin
			if (main_sdram_bankmachine2_trccon_ready) begin
				main_sdram_bankmachine2_row_col_n_addr_sel <= 1'd1;
				main_sdram_bankmachine2_row_open <= 1'd1;
				main_sdram_bankmachine2_cmd_valid <= 1'd1;
				main_sdram_bankmachine2_cmd_payload_is_cmd <= 1'd1;
				if (main_sdram_bankmachine2_cmd_ready) begin
					builder_bankmachine2_next_state <= 3'd6;
				end
				main_sdram_bankmachine2_cmd_payload_ras <= 1'd1;
			end
		end
		3'd4: begin
			if (main_sdram_bankmachine2_twtpcon_ready) begin
				main_sdram_bankmachine2_refresh_gnt <= 1'd1;
			end
			main_sdram_bankmachine2_row_close <= 1'd1;
			main_sdram_bankmachine2_cmd_payload_is_cmd <= 1'd1;
			if ((~main_sdram_bankmachine2_refresh_req)) begin
				builder_bankmachine2_next_state <= 1'd0;
			end
		end
		3'd5: begin
			builder_bankmachine2_next_state <= 2'd3;
		end
		3'd6: begin
			builder_bankmachine2_next_state <= 1'd0;
		end
		default: begin
			if (main_sdram_bankmachine2_refresh_req) begin
				builder_bankmachine2_next_state <= 3'd4;
			end else begin
				if (main_sdram_bankmachine2_cmd_buffer_source_valid) begin
					if (main_sdram_bankmachine2_row_opened) begin
						if (main_sdram_bankmachine2_row_hit) begin
							main_sdram_bankmachine2_cmd_valid <= 1'd1;
							if (main_sdram_bankmachine2_cmd_buffer_source_payload_we) begin
								main_sdram_bankmachine2_req_wdata_ready <= main_sdram_bankmachine2_cmd_ready;
								main_sdram_bankmachine2_cmd_payload_is_write <= 1'd1;
								main_sdram_bankmachine2_cmd_payload_we <= 1'd1;
							end else begin
								main_sdram_bankmachine2_req_rdata_valid <= main_sdram_bankmachine2_cmd_ready;
								main_sdram_bankmachine2_cmd_payload_is_read <= 1'd1;
							end
							main_sdram_bankmachine2_cmd_payload_cas <= 1'd1;
							if ((main_sdram_bankmachine2_cmd_ready & main_sdram_bankmachine2_auto_precharge)) begin
								builder_bankmachine2_next_state <= 2'd2;
							end
						end else begin
							builder_bankmachine2_next_state <= 1'd1;
						end
					end else begin
						builder_bankmachine2_next_state <= 2'd3;
					end
				end
			end
		end
	endcase
end
assign main_sdram_bankmachine3_cmd_buffer_lookahead_sink_valid = main_sdram_bankmachine3_req_valid;
assign main_sdram_bankmachine3_req_ready = main_sdram_bankmachine3_cmd_buffer_lookahead_sink_ready;
assign main_sdram_bankmachine3_cmd_buffer_lookahead_sink_payload_we = main_sdram_bankmachine3_req_we;
assign main_sdram_bankmachine3_cmd_buffer_lookahead_sink_payload_addr = main_sdram_bankmachine3_req_addr;
assign main_sdram_bankmachine3_cmd_buffer_sink_valid = main_sdram_bankmachine3_cmd_buffer_lookahead_source_valid;
assign main_sdram_bankmachine3_cmd_buffer_lookahead_source_ready = main_sdram_bankmachine3_cmd_buffer_sink_ready;
assign main_sdram_bankmachine3_cmd_buffer_sink_first = main_sdram_bankmachine3_cmd_buffer_lookahead_source_first;
assign main_sdram_bankmachine3_cmd_buffer_sink_last = main_sdram_bankmachine3_cmd_buffer_lookahead_source_last;
assign main_sdram_bankmachine3_cmd_buffer_sink_payload_we = main_sdram_bankmachine3_cmd_buffer_lookahead_source_payload_we;
assign main_sdram_bankmachine3_cmd_buffer_sink_payload_addr = main_sdram_bankmachine3_cmd_buffer_lookahead_source_payload_addr;
assign main_sdram_bankmachine3_cmd_buffer_source_ready = (main_sdram_bankmachine3_req_wdata_ready | main_sdram_bankmachine3_req_rdata_valid);
assign main_sdram_bankmachine3_req_lock = (main_sdram_bankmachine3_cmd_buffer_lookahead_source_valid | main_sdram_bankmachine3_cmd_buffer_source_valid);
assign main_sdram_bankmachine3_row_hit = (main_sdram_bankmachine3_row == main_sdram_bankmachine3_cmd_buffer_source_payload_addr[20:7]);
assign main_sdram_bankmachine3_cmd_payload_ba = 2'd3;
always @(*) begin
	main_sdram_bankmachine3_cmd_payload_a <= 14'd0;
	if (main_sdram_bankmachine3_row_col_n_addr_sel) begin
		main_sdram_bankmachine3_cmd_payload_a <= main_sdram_bankmachine3_cmd_buffer_source_payload_addr[20:7];
	end else begin
		main_sdram_bankmachine3_cmd_payload_a <= ((main_sdram_bankmachine3_auto_precharge <<< 4'd10) | {main_sdram_bankmachine3_cmd_buffer_source_payload_addr[6:0], {3{1'd0}}});
	end
end
assign main_sdram_bankmachine3_twtpcon_valid = ((main_sdram_bankmachine3_cmd_valid & main_sdram_bankmachine3_cmd_ready) & main_sdram_bankmachine3_cmd_payload_is_write);
assign main_sdram_bankmachine3_trccon_valid = ((main_sdram_bankmachine3_cmd_valid & main_sdram_bankmachine3_cmd_ready) & main_sdram_bankmachine3_row_open);
assign main_sdram_bankmachine3_trascon_valid = ((main_sdram_bankmachine3_cmd_valid & main_sdram_bankmachine3_cmd_ready) & main_sdram_bankmachine3_row_open);
always @(*) begin
	main_sdram_bankmachine3_auto_precharge <= 1'd0;
	if ((main_sdram_bankmachine3_cmd_buffer_lookahead_source_valid & main_sdram_bankmachine3_cmd_buffer_source_valid)) begin
		if ((main_sdram_bankmachine3_cmd_buffer_lookahead_source_payload_addr[20:7] != main_sdram_bankmachine3_cmd_buffer_source_payload_addr[20:7])) begin
			main_sdram_bankmachine3_auto_precharge <= (main_sdram_bankmachine3_row_close == 1'd0);
		end
	end
end
assign main_sdram_bankmachine3_cmd_buffer_lookahead_syncfifo3_din = {main_sdram_bankmachine3_cmd_buffer_lookahead_fifo_in_last, main_sdram_bankmachine3_cmd_buffer_lookahead_fifo_in_first, main_sdram_bankmachine3_cmd_buffer_lookahead_fifo_in_payload_addr, main_sdram_bankmachine3_cmd_buffer_lookahead_fifo_in_payload_we};
assign {main_sdram_bankmachine3_cmd_buffer_lookahead_fifo_out_last, main_sdram_bankmachine3_cmd_buffer_lookahead_fifo_out_first, main_sdram_bankmachine3_cmd_buffer_lookahead_fifo_out_payload_addr, main_sdram_bankmachine3_cmd_buffer_lookahead_fifo_out_payload_we} = main_sdram_bankmachine3_cmd_buffer_lookahead_syncfifo3_dout;
assign main_sdram_bankmachine3_cmd_buffer_lookahead_sink_ready = main_sdram_bankmachine3_cmd_buffer_lookahead_syncfifo3_writable;
assign main_sdram_bankmachine3_cmd_buffer_lookahead_syncfifo3_we = main_sdram_bankmachine3_cmd_buffer_lookahead_sink_valid;
assign main_sdram_bankmachine3_cmd_buffer_lookahead_fifo_in_first = main_sdram_bankmachine3_cmd_buffer_lookahead_sink_first;
assign main_sdram_bankmachine3_cmd_buffer_lookahead_fifo_in_last = main_sdram_bankmachine3_cmd_buffer_lookahead_sink_last;
assign main_sdram_bankmachine3_cmd_buffer_lookahead_fifo_in_payload_we = main_sdram_bankmachine3_cmd_buffer_lookahead_sink_payload_we;
assign main_sdram_bankmachine3_cmd_buffer_lookahead_fifo_in_payload_addr = main_sdram_bankmachine3_cmd_buffer_lookahead_sink_payload_addr;
assign main_sdram_bankmachine3_cmd_buffer_lookahead_source_valid = main_sdram_bankmachine3_cmd_buffer_lookahead_syncfifo3_readable;
assign main_sdram_bankmachine3_cmd_buffer_lookahead_source_first = main_sdram_bankmachine3_cmd_buffer_lookahead_fifo_out_first;
assign main_sdram_bankmachine3_cmd_buffer_lookahead_source_last = main_sdram_bankmachine3_cmd_buffer_lookahead_fifo_out_last;
assign main_sdram_bankmachine3_cmd_buffer_lookahead_source_payload_we = main_sdram_bankmachine3_cmd_buffer_lookahead_fifo_out_payload_we;
assign main_sdram_bankmachine3_cmd_buffer_lookahead_source_payload_addr = main_sdram_bankmachine3_cmd_buffer_lookahead_fifo_out_payload_addr;
assign main_sdram_bankmachine3_cmd_buffer_lookahead_syncfifo3_re = main_sdram_bankmachine3_cmd_buffer_lookahead_source_ready;
always @(*) begin
	main_sdram_bankmachine3_cmd_buffer_lookahead_wrport_adr <= 3'd0;
	if (main_sdram_bankmachine3_cmd_buffer_lookahead_replace) begin
		main_sdram_bankmachine3_cmd_buffer_lookahead_wrport_adr <= (main_sdram_bankmachine3_cmd_buffer_lookahead_produce - 1'd1);
	end else begin
		main_sdram_bankmachine3_cmd_buffer_lookahead_wrport_adr <= main_sdram_bankmachine3_cmd_buffer_lookahead_produce;
	end
end
assign main_sdram_bankmachine3_cmd_buffer_lookahead_wrport_dat_w = main_sdram_bankmachine3_cmd_buffer_lookahead_syncfifo3_din;
assign main_sdram_bankmachine3_cmd_buffer_lookahead_wrport_we = (main_sdram_bankmachine3_cmd_buffer_lookahead_syncfifo3_we & (main_sdram_bankmachine3_cmd_buffer_lookahead_syncfifo3_writable | main_sdram_bankmachine3_cmd_buffer_lookahead_replace));
assign main_sdram_bankmachine3_cmd_buffer_lookahead_do_read = (main_sdram_bankmachine3_cmd_buffer_lookahead_syncfifo3_readable & main_sdram_bankmachine3_cmd_buffer_lookahead_syncfifo3_re);
assign main_sdram_bankmachine3_cmd_buffer_lookahead_rdport_adr = main_sdram_bankmachine3_cmd_buffer_lookahead_consume;
assign main_sdram_bankmachine3_cmd_buffer_lookahead_syncfifo3_dout = main_sdram_bankmachine3_cmd_buffer_lookahead_rdport_dat_r;
assign main_sdram_bankmachine3_cmd_buffer_lookahead_syncfifo3_writable = (main_sdram_bankmachine3_cmd_buffer_lookahead_level != 4'd8);
assign main_sdram_bankmachine3_cmd_buffer_lookahead_syncfifo3_readable = (main_sdram_bankmachine3_cmd_buffer_lookahead_level != 1'd0);
assign main_sdram_bankmachine3_cmd_buffer_sink_ready = ((~main_sdram_bankmachine3_cmd_buffer_source_valid) | main_sdram_bankmachine3_cmd_buffer_source_ready);
always @(*) begin
	main_sdram_bankmachine3_cmd_payload_cas <= 1'd0;
	builder_bankmachine3_next_state <= 3'd0;
	main_sdram_bankmachine3_cmd_payload_ras <= 1'd0;
	main_sdram_bankmachine3_cmd_payload_we <= 1'd0;
	main_sdram_bankmachine3_row_col_n_addr_sel <= 1'd0;
	main_sdram_bankmachine3_cmd_payload_is_cmd <= 1'd0;
	main_sdram_bankmachine3_cmd_payload_is_read <= 1'd0;
	main_sdram_bankmachine3_cmd_payload_is_write <= 1'd0;
	main_sdram_bankmachine3_req_wdata_ready <= 1'd0;
	main_sdram_bankmachine3_req_rdata_valid <= 1'd0;
	main_sdram_bankmachine3_refresh_gnt <= 1'd0;
	main_sdram_bankmachine3_cmd_valid <= 1'd0;
	main_sdram_bankmachine3_row_open <= 1'd0;
	main_sdram_bankmachine3_row_close <= 1'd0;
	builder_bankmachine3_next_state <= builder_bankmachine3_state;
	case (builder_bankmachine3_state)
		1'd1: begin
			if ((main_sdram_bankmachine3_twtpcon_ready & main_sdram_bankmachine3_trascon_ready)) begin
				main_sdram_bankmachine3_cmd_valid <= 1'd1;
				if (main_sdram_bankmachine3_cmd_ready) begin
					builder_bankmachine3_next_state <= 3'd5;
				end
				main_sdram_bankmachine3_cmd_payload_ras <= 1'd1;
				main_sdram_bankmachine3_cmd_payload_we <= 1'd1;
				main_sdram_bankmachine3_cmd_payload_is_cmd <= 1'd1;
			end
			main_sdram_bankmachine3_row_close <= 1'd1;
		end
		2'd2: begin
			if ((main_sdram_bankmachine3_twtpcon_ready & main_sdram_bankmachine3_trascon_ready)) begin
				builder_bankmachine3_next_state <= 3'd5;
			end
			main_sdram_bankmachine3_row_close <= 1'd1;
		end
		2'd3: begin
			if (main_sdram_bankmachine3_trccon_ready) begin
				main_sdram_bankmachine3_row_col_n_addr_sel <= 1'd1;
				main_sdram_bankmachine3_row_open <= 1'd1;
				main_sdram_bankmachine3_cmd_valid <= 1'd1;
				main_sdram_bankmachine3_cmd_payload_is_cmd <= 1'd1;
				if (main_sdram_bankmachine3_cmd_ready) begin
					builder_bankmachine3_next_state <= 3'd6;
				end
				main_sdram_bankmachine3_cmd_payload_ras <= 1'd1;
			end
		end
		3'd4: begin
			if (main_sdram_bankmachine3_twtpcon_ready) begin
				main_sdram_bankmachine3_refresh_gnt <= 1'd1;
			end
			main_sdram_bankmachine3_row_close <= 1'd1;
			main_sdram_bankmachine3_cmd_payload_is_cmd <= 1'd1;
			if ((~main_sdram_bankmachine3_refresh_req)) begin
				builder_bankmachine3_next_state <= 1'd0;
			end
		end
		3'd5: begin
			builder_bankmachine3_next_state <= 2'd3;
		end
		3'd6: begin
			builder_bankmachine3_next_state <= 1'd0;
		end
		default: begin
			if (main_sdram_bankmachine3_refresh_req) begin
				builder_bankmachine3_next_state <= 3'd4;
			end else begin
				if (main_sdram_bankmachine3_cmd_buffer_source_valid) begin
					if (main_sdram_bankmachine3_row_opened) begin
						if (main_sdram_bankmachine3_row_hit) begin
							main_sdram_bankmachine3_cmd_valid <= 1'd1;
							if (main_sdram_bankmachine3_cmd_buffer_source_payload_we) begin
								main_sdram_bankmachine3_req_wdata_ready <= main_sdram_bankmachine3_cmd_ready;
								main_sdram_bankmachine3_cmd_payload_is_write <= 1'd1;
								main_sdram_bankmachine3_cmd_payload_we <= 1'd1;
							end else begin
								main_sdram_bankmachine3_req_rdata_valid <= main_sdram_bankmachine3_cmd_ready;
								main_sdram_bankmachine3_cmd_payload_is_read <= 1'd1;
							end
							main_sdram_bankmachine3_cmd_payload_cas <= 1'd1;
							if ((main_sdram_bankmachine3_cmd_ready & main_sdram_bankmachine3_auto_precharge)) begin
								builder_bankmachine3_next_state <= 2'd2;
							end
						end else begin
							builder_bankmachine3_next_state <= 1'd1;
						end
					end else begin
						builder_bankmachine3_next_state <= 2'd3;
					end
				end
			end
		end
	endcase
end
assign main_sdram_bankmachine4_cmd_buffer_lookahead_sink_valid = main_sdram_bankmachine4_req_valid;
assign main_sdram_bankmachine4_req_ready = main_sdram_bankmachine4_cmd_buffer_lookahead_sink_ready;
assign main_sdram_bankmachine4_cmd_buffer_lookahead_sink_payload_we = main_sdram_bankmachine4_req_we;
assign main_sdram_bankmachine4_cmd_buffer_lookahead_sink_payload_addr = main_sdram_bankmachine4_req_addr;
assign main_sdram_bankmachine4_cmd_buffer_sink_valid = main_sdram_bankmachine4_cmd_buffer_lookahead_source_valid;
assign main_sdram_bankmachine4_cmd_buffer_lookahead_source_ready = main_sdram_bankmachine4_cmd_buffer_sink_ready;
assign main_sdram_bankmachine4_cmd_buffer_sink_first = main_sdram_bankmachine4_cmd_buffer_lookahead_source_first;
assign main_sdram_bankmachine4_cmd_buffer_sink_last = main_sdram_bankmachine4_cmd_buffer_lookahead_source_last;
assign main_sdram_bankmachine4_cmd_buffer_sink_payload_we = main_sdram_bankmachine4_cmd_buffer_lookahead_source_payload_we;
assign main_sdram_bankmachine4_cmd_buffer_sink_payload_addr = main_sdram_bankmachine4_cmd_buffer_lookahead_source_payload_addr;
assign main_sdram_bankmachine4_cmd_buffer_source_ready = (main_sdram_bankmachine4_req_wdata_ready | main_sdram_bankmachine4_req_rdata_valid);
assign main_sdram_bankmachine4_req_lock = (main_sdram_bankmachine4_cmd_buffer_lookahead_source_valid | main_sdram_bankmachine4_cmd_buffer_source_valid);
assign main_sdram_bankmachine4_row_hit = (main_sdram_bankmachine4_row == main_sdram_bankmachine4_cmd_buffer_source_payload_addr[20:7]);
assign main_sdram_bankmachine4_cmd_payload_ba = 3'd4;
always @(*) begin
	main_sdram_bankmachine4_cmd_payload_a <= 14'd0;
	if (main_sdram_bankmachine4_row_col_n_addr_sel) begin
		main_sdram_bankmachine4_cmd_payload_a <= main_sdram_bankmachine4_cmd_buffer_source_payload_addr[20:7];
	end else begin
		main_sdram_bankmachine4_cmd_payload_a <= ((main_sdram_bankmachine4_auto_precharge <<< 4'd10) | {main_sdram_bankmachine4_cmd_buffer_source_payload_addr[6:0], {3{1'd0}}});
	end
end
assign main_sdram_bankmachine4_twtpcon_valid = ((main_sdram_bankmachine4_cmd_valid & main_sdram_bankmachine4_cmd_ready) & main_sdram_bankmachine4_cmd_payload_is_write);
assign main_sdram_bankmachine4_trccon_valid = ((main_sdram_bankmachine4_cmd_valid & main_sdram_bankmachine4_cmd_ready) & main_sdram_bankmachine4_row_open);
assign main_sdram_bankmachine4_trascon_valid = ((main_sdram_bankmachine4_cmd_valid & main_sdram_bankmachine4_cmd_ready) & main_sdram_bankmachine4_row_open);
always @(*) begin
	main_sdram_bankmachine4_auto_precharge <= 1'd0;
	if ((main_sdram_bankmachine4_cmd_buffer_lookahead_source_valid & main_sdram_bankmachine4_cmd_buffer_source_valid)) begin
		if ((main_sdram_bankmachine4_cmd_buffer_lookahead_source_payload_addr[20:7] != main_sdram_bankmachine4_cmd_buffer_source_payload_addr[20:7])) begin
			main_sdram_bankmachine4_auto_precharge <= (main_sdram_bankmachine4_row_close == 1'd0);
		end
	end
end
assign main_sdram_bankmachine4_cmd_buffer_lookahead_syncfifo4_din = {main_sdram_bankmachine4_cmd_buffer_lookahead_fifo_in_last, main_sdram_bankmachine4_cmd_buffer_lookahead_fifo_in_first, main_sdram_bankmachine4_cmd_buffer_lookahead_fifo_in_payload_addr, main_sdram_bankmachine4_cmd_buffer_lookahead_fifo_in_payload_we};
assign {main_sdram_bankmachine4_cmd_buffer_lookahead_fifo_out_last, main_sdram_bankmachine4_cmd_buffer_lookahead_fifo_out_first, main_sdram_bankmachine4_cmd_buffer_lookahead_fifo_out_payload_addr, main_sdram_bankmachine4_cmd_buffer_lookahead_fifo_out_payload_we} = main_sdram_bankmachine4_cmd_buffer_lookahead_syncfifo4_dout;
assign main_sdram_bankmachine4_cmd_buffer_lookahead_sink_ready = main_sdram_bankmachine4_cmd_buffer_lookahead_syncfifo4_writable;
assign main_sdram_bankmachine4_cmd_buffer_lookahead_syncfifo4_we = main_sdram_bankmachine4_cmd_buffer_lookahead_sink_valid;
assign main_sdram_bankmachine4_cmd_buffer_lookahead_fifo_in_first = main_sdram_bankmachine4_cmd_buffer_lookahead_sink_first;
assign main_sdram_bankmachine4_cmd_buffer_lookahead_fifo_in_last = main_sdram_bankmachine4_cmd_buffer_lookahead_sink_last;
assign main_sdram_bankmachine4_cmd_buffer_lookahead_fifo_in_payload_we = main_sdram_bankmachine4_cmd_buffer_lookahead_sink_payload_we;
assign main_sdram_bankmachine4_cmd_buffer_lookahead_fifo_in_payload_addr = main_sdram_bankmachine4_cmd_buffer_lookahead_sink_payload_addr;
assign main_sdram_bankmachine4_cmd_buffer_lookahead_source_valid = main_sdram_bankmachine4_cmd_buffer_lookahead_syncfifo4_readable;
assign main_sdram_bankmachine4_cmd_buffer_lookahead_source_first = main_sdram_bankmachine4_cmd_buffer_lookahead_fifo_out_first;
assign main_sdram_bankmachine4_cmd_buffer_lookahead_source_last = main_sdram_bankmachine4_cmd_buffer_lookahead_fifo_out_last;
assign main_sdram_bankmachine4_cmd_buffer_lookahead_source_payload_we = main_sdram_bankmachine4_cmd_buffer_lookahead_fifo_out_payload_we;
assign main_sdram_bankmachine4_cmd_buffer_lookahead_source_payload_addr = main_sdram_bankmachine4_cmd_buffer_lookahead_fifo_out_payload_addr;
assign main_sdram_bankmachine4_cmd_buffer_lookahead_syncfifo4_re = main_sdram_bankmachine4_cmd_buffer_lookahead_source_ready;
always @(*) begin
	main_sdram_bankmachine4_cmd_buffer_lookahead_wrport_adr <= 3'd0;
	if (main_sdram_bankmachine4_cmd_buffer_lookahead_replace) begin
		main_sdram_bankmachine4_cmd_buffer_lookahead_wrport_adr <= (main_sdram_bankmachine4_cmd_buffer_lookahead_produce - 1'd1);
	end else begin
		main_sdram_bankmachine4_cmd_buffer_lookahead_wrport_adr <= main_sdram_bankmachine4_cmd_buffer_lookahead_produce;
	end
end
assign main_sdram_bankmachine4_cmd_buffer_lookahead_wrport_dat_w = main_sdram_bankmachine4_cmd_buffer_lookahead_syncfifo4_din;
assign main_sdram_bankmachine4_cmd_buffer_lookahead_wrport_we = (main_sdram_bankmachine4_cmd_buffer_lookahead_syncfifo4_we & (main_sdram_bankmachine4_cmd_buffer_lookahead_syncfifo4_writable | main_sdram_bankmachine4_cmd_buffer_lookahead_replace));
assign main_sdram_bankmachine4_cmd_buffer_lookahead_do_read = (main_sdram_bankmachine4_cmd_buffer_lookahead_syncfifo4_readable & main_sdram_bankmachine4_cmd_buffer_lookahead_syncfifo4_re);
assign main_sdram_bankmachine4_cmd_buffer_lookahead_rdport_adr = main_sdram_bankmachine4_cmd_buffer_lookahead_consume;
assign main_sdram_bankmachine4_cmd_buffer_lookahead_syncfifo4_dout = main_sdram_bankmachine4_cmd_buffer_lookahead_rdport_dat_r;
assign main_sdram_bankmachine4_cmd_buffer_lookahead_syncfifo4_writable = (main_sdram_bankmachine4_cmd_buffer_lookahead_level != 4'd8);
assign main_sdram_bankmachine4_cmd_buffer_lookahead_syncfifo4_readable = (main_sdram_bankmachine4_cmd_buffer_lookahead_level != 1'd0);
assign main_sdram_bankmachine4_cmd_buffer_sink_ready = ((~main_sdram_bankmachine4_cmd_buffer_source_valid) | main_sdram_bankmachine4_cmd_buffer_source_ready);
always @(*) begin
	main_sdram_bankmachine4_cmd_payload_cas <= 1'd0;
	main_sdram_bankmachine4_row_close <= 1'd0;
	main_sdram_bankmachine4_cmd_payload_ras <= 1'd0;
	main_sdram_bankmachine4_cmd_payload_we <= 1'd0;
	main_sdram_bankmachine4_row_col_n_addr_sel <= 1'd0;
	main_sdram_bankmachine4_cmd_payload_is_cmd <= 1'd0;
	main_sdram_bankmachine4_cmd_payload_is_read <= 1'd0;
	main_sdram_bankmachine4_cmd_payload_is_write <= 1'd0;
	main_sdram_bankmachine4_req_wdata_ready <= 1'd0;
	main_sdram_bankmachine4_req_rdata_valid <= 1'd0;
	main_sdram_bankmachine4_refresh_gnt <= 1'd0;
	main_sdram_bankmachine4_cmd_valid <= 1'd0;
	main_sdram_bankmachine4_row_open <= 1'd0;
	builder_bankmachine4_next_state <= 3'd0;
	builder_bankmachine4_next_state <= builder_bankmachine4_state;
	case (builder_bankmachine4_state)
		1'd1: begin
			if ((main_sdram_bankmachine4_twtpcon_ready & main_sdram_bankmachine4_trascon_ready)) begin
				main_sdram_bankmachine4_cmd_valid <= 1'd1;
				if (main_sdram_bankmachine4_cmd_ready) begin
					builder_bankmachine4_next_state <= 3'd5;
				end
				main_sdram_bankmachine4_cmd_payload_ras <= 1'd1;
				main_sdram_bankmachine4_cmd_payload_we <= 1'd1;
				main_sdram_bankmachine4_cmd_payload_is_cmd <= 1'd1;
			end
			main_sdram_bankmachine4_row_close <= 1'd1;
		end
		2'd2: begin
			if ((main_sdram_bankmachine4_twtpcon_ready & main_sdram_bankmachine4_trascon_ready)) begin
				builder_bankmachine4_next_state <= 3'd5;
			end
			main_sdram_bankmachine4_row_close <= 1'd1;
		end
		2'd3: begin
			if (main_sdram_bankmachine4_trccon_ready) begin
				main_sdram_bankmachine4_row_col_n_addr_sel <= 1'd1;
				main_sdram_bankmachine4_row_open <= 1'd1;
				main_sdram_bankmachine4_cmd_valid <= 1'd1;
				main_sdram_bankmachine4_cmd_payload_is_cmd <= 1'd1;
				if (main_sdram_bankmachine4_cmd_ready) begin
					builder_bankmachine4_next_state <= 3'd6;
				end
				main_sdram_bankmachine4_cmd_payload_ras <= 1'd1;
			end
		end
		3'd4: begin
			if (main_sdram_bankmachine4_twtpcon_ready) begin
				main_sdram_bankmachine4_refresh_gnt <= 1'd1;
			end
			main_sdram_bankmachine4_row_close <= 1'd1;
			main_sdram_bankmachine4_cmd_payload_is_cmd <= 1'd1;
			if ((~main_sdram_bankmachine4_refresh_req)) begin
				builder_bankmachine4_next_state <= 1'd0;
			end
		end
		3'd5: begin
			builder_bankmachine4_next_state <= 2'd3;
		end
		3'd6: begin
			builder_bankmachine4_next_state <= 1'd0;
		end
		default: begin
			if (main_sdram_bankmachine4_refresh_req) begin
				builder_bankmachine4_next_state <= 3'd4;
			end else begin
				if (main_sdram_bankmachine4_cmd_buffer_source_valid) begin
					if (main_sdram_bankmachine4_row_opened) begin
						if (main_sdram_bankmachine4_row_hit) begin
							main_sdram_bankmachine4_cmd_valid <= 1'd1;
							if (main_sdram_bankmachine4_cmd_buffer_source_payload_we) begin
								main_sdram_bankmachine4_req_wdata_ready <= main_sdram_bankmachine4_cmd_ready;
								main_sdram_bankmachine4_cmd_payload_is_write <= 1'd1;
								main_sdram_bankmachine4_cmd_payload_we <= 1'd1;
							end else begin
								main_sdram_bankmachine4_req_rdata_valid <= main_sdram_bankmachine4_cmd_ready;
								main_sdram_bankmachine4_cmd_payload_is_read <= 1'd1;
							end
							main_sdram_bankmachine4_cmd_payload_cas <= 1'd1;
							if ((main_sdram_bankmachine4_cmd_ready & main_sdram_bankmachine4_auto_precharge)) begin
								builder_bankmachine4_next_state <= 2'd2;
							end
						end else begin
							builder_bankmachine4_next_state <= 1'd1;
						end
					end else begin
						builder_bankmachine4_next_state <= 2'd3;
					end
				end
			end
		end
	endcase
end
assign main_sdram_bankmachine5_cmd_buffer_lookahead_sink_valid = main_sdram_bankmachine5_req_valid;
assign main_sdram_bankmachine5_req_ready = main_sdram_bankmachine5_cmd_buffer_lookahead_sink_ready;
assign main_sdram_bankmachine5_cmd_buffer_lookahead_sink_payload_we = main_sdram_bankmachine5_req_we;
assign main_sdram_bankmachine5_cmd_buffer_lookahead_sink_payload_addr = main_sdram_bankmachine5_req_addr;
assign main_sdram_bankmachine5_cmd_buffer_sink_valid = main_sdram_bankmachine5_cmd_buffer_lookahead_source_valid;
assign main_sdram_bankmachine5_cmd_buffer_lookahead_source_ready = main_sdram_bankmachine5_cmd_buffer_sink_ready;
assign main_sdram_bankmachine5_cmd_buffer_sink_first = main_sdram_bankmachine5_cmd_buffer_lookahead_source_first;
assign main_sdram_bankmachine5_cmd_buffer_sink_last = main_sdram_bankmachine5_cmd_buffer_lookahead_source_last;
assign main_sdram_bankmachine5_cmd_buffer_sink_payload_we = main_sdram_bankmachine5_cmd_buffer_lookahead_source_payload_we;
assign main_sdram_bankmachine5_cmd_buffer_sink_payload_addr = main_sdram_bankmachine5_cmd_buffer_lookahead_source_payload_addr;
assign main_sdram_bankmachine5_cmd_buffer_source_ready = (main_sdram_bankmachine5_req_wdata_ready | main_sdram_bankmachine5_req_rdata_valid);
assign main_sdram_bankmachine5_req_lock = (main_sdram_bankmachine5_cmd_buffer_lookahead_source_valid | main_sdram_bankmachine5_cmd_buffer_source_valid);
assign main_sdram_bankmachine5_row_hit = (main_sdram_bankmachine5_row == main_sdram_bankmachine5_cmd_buffer_source_payload_addr[20:7]);
assign main_sdram_bankmachine5_cmd_payload_ba = 3'd5;
always @(*) begin
	main_sdram_bankmachine5_cmd_payload_a <= 14'd0;
	if (main_sdram_bankmachine5_row_col_n_addr_sel) begin
		main_sdram_bankmachine5_cmd_payload_a <= main_sdram_bankmachine5_cmd_buffer_source_payload_addr[20:7];
	end else begin
		main_sdram_bankmachine5_cmd_payload_a <= ((main_sdram_bankmachine5_auto_precharge <<< 4'd10) | {main_sdram_bankmachine5_cmd_buffer_source_payload_addr[6:0], {3{1'd0}}});
	end
end
assign main_sdram_bankmachine5_twtpcon_valid = ((main_sdram_bankmachine5_cmd_valid & main_sdram_bankmachine5_cmd_ready) & main_sdram_bankmachine5_cmd_payload_is_write);
assign main_sdram_bankmachine5_trccon_valid = ((main_sdram_bankmachine5_cmd_valid & main_sdram_bankmachine5_cmd_ready) & main_sdram_bankmachine5_row_open);
assign main_sdram_bankmachine5_trascon_valid = ((main_sdram_bankmachine5_cmd_valid & main_sdram_bankmachine5_cmd_ready) & main_sdram_bankmachine5_row_open);
always @(*) begin
	main_sdram_bankmachine5_auto_precharge <= 1'd0;
	if ((main_sdram_bankmachine5_cmd_buffer_lookahead_source_valid & main_sdram_bankmachine5_cmd_buffer_source_valid)) begin
		if ((main_sdram_bankmachine5_cmd_buffer_lookahead_source_payload_addr[20:7] != main_sdram_bankmachine5_cmd_buffer_source_payload_addr[20:7])) begin
			main_sdram_bankmachine5_auto_precharge <= (main_sdram_bankmachine5_row_close == 1'd0);
		end
	end
end
assign main_sdram_bankmachine5_cmd_buffer_lookahead_syncfifo5_din = {main_sdram_bankmachine5_cmd_buffer_lookahead_fifo_in_last, main_sdram_bankmachine5_cmd_buffer_lookahead_fifo_in_first, main_sdram_bankmachine5_cmd_buffer_lookahead_fifo_in_payload_addr, main_sdram_bankmachine5_cmd_buffer_lookahead_fifo_in_payload_we};
assign {main_sdram_bankmachine5_cmd_buffer_lookahead_fifo_out_last, main_sdram_bankmachine5_cmd_buffer_lookahead_fifo_out_first, main_sdram_bankmachine5_cmd_buffer_lookahead_fifo_out_payload_addr, main_sdram_bankmachine5_cmd_buffer_lookahead_fifo_out_payload_we} = main_sdram_bankmachine5_cmd_buffer_lookahead_syncfifo5_dout;
assign main_sdram_bankmachine5_cmd_buffer_lookahead_sink_ready = main_sdram_bankmachine5_cmd_buffer_lookahead_syncfifo5_writable;
assign main_sdram_bankmachine5_cmd_buffer_lookahead_syncfifo5_we = main_sdram_bankmachine5_cmd_buffer_lookahead_sink_valid;
assign main_sdram_bankmachine5_cmd_buffer_lookahead_fifo_in_first = main_sdram_bankmachine5_cmd_buffer_lookahead_sink_first;
assign main_sdram_bankmachine5_cmd_buffer_lookahead_fifo_in_last = main_sdram_bankmachine5_cmd_buffer_lookahead_sink_last;
assign main_sdram_bankmachine5_cmd_buffer_lookahead_fifo_in_payload_we = main_sdram_bankmachine5_cmd_buffer_lookahead_sink_payload_we;
assign main_sdram_bankmachine5_cmd_buffer_lookahead_fifo_in_payload_addr = main_sdram_bankmachine5_cmd_buffer_lookahead_sink_payload_addr;
assign main_sdram_bankmachine5_cmd_buffer_lookahead_source_valid = main_sdram_bankmachine5_cmd_buffer_lookahead_syncfifo5_readable;
assign main_sdram_bankmachine5_cmd_buffer_lookahead_source_first = main_sdram_bankmachine5_cmd_buffer_lookahead_fifo_out_first;
assign main_sdram_bankmachine5_cmd_buffer_lookahead_source_last = main_sdram_bankmachine5_cmd_buffer_lookahead_fifo_out_last;
assign main_sdram_bankmachine5_cmd_buffer_lookahead_source_payload_we = main_sdram_bankmachine5_cmd_buffer_lookahead_fifo_out_payload_we;
assign main_sdram_bankmachine5_cmd_buffer_lookahead_source_payload_addr = main_sdram_bankmachine5_cmd_buffer_lookahead_fifo_out_payload_addr;
assign main_sdram_bankmachine5_cmd_buffer_lookahead_syncfifo5_re = main_sdram_bankmachine5_cmd_buffer_lookahead_source_ready;
always @(*) begin
	main_sdram_bankmachine5_cmd_buffer_lookahead_wrport_adr <= 3'd0;
	if (main_sdram_bankmachine5_cmd_buffer_lookahead_replace) begin
		main_sdram_bankmachine5_cmd_buffer_lookahead_wrport_adr <= (main_sdram_bankmachine5_cmd_buffer_lookahead_produce - 1'd1);
	end else begin
		main_sdram_bankmachine5_cmd_buffer_lookahead_wrport_adr <= main_sdram_bankmachine5_cmd_buffer_lookahead_produce;
	end
end
assign main_sdram_bankmachine5_cmd_buffer_lookahead_wrport_dat_w = main_sdram_bankmachine5_cmd_buffer_lookahead_syncfifo5_din;
assign main_sdram_bankmachine5_cmd_buffer_lookahead_wrport_we = (main_sdram_bankmachine5_cmd_buffer_lookahead_syncfifo5_we & (main_sdram_bankmachine5_cmd_buffer_lookahead_syncfifo5_writable | main_sdram_bankmachine5_cmd_buffer_lookahead_replace));
assign main_sdram_bankmachine5_cmd_buffer_lookahead_do_read = (main_sdram_bankmachine5_cmd_buffer_lookahead_syncfifo5_readable & main_sdram_bankmachine5_cmd_buffer_lookahead_syncfifo5_re);
assign main_sdram_bankmachine5_cmd_buffer_lookahead_rdport_adr = main_sdram_bankmachine5_cmd_buffer_lookahead_consume;
assign main_sdram_bankmachine5_cmd_buffer_lookahead_syncfifo5_dout = main_sdram_bankmachine5_cmd_buffer_lookahead_rdport_dat_r;
assign main_sdram_bankmachine5_cmd_buffer_lookahead_syncfifo5_writable = (main_sdram_bankmachine5_cmd_buffer_lookahead_level != 4'd8);
assign main_sdram_bankmachine5_cmd_buffer_lookahead_syncfifo5_readable = (main_sdram_bankmachine5_cmd_buffer_lookahead_level != 1'd0);
assign main_sdram_bankmachine5_cmd_buffer_sink_ready = ((~main_sdram_bankmachine5_cmd_buffer_source_valid) | main_sdram_bankmachine5_cmd_buffer_source_ready);
always @(*) begin
	main_sdram_bankmachine5_cmd_payload_cas <= 1'd0;
	main_sdram_bankmachine5_cmd_payload_ras <= 1'd0;
	main_sdram_bankmachine5_cmd_payload_we <= 1'd0;
	main_sdram_bankmachine5_row_col_n_addr_sel <= 1'd0;
	main_sdram_bankmachine5_cmd_payload_is_cmd <= 1'd0;
	main_sdram_bankmachine5_cmd_payload_is_read <= 1'd0;
	main_sdram_bankmachine5_cmd_payload_is_write <= 1'd0;
	main_sdram_bankmachine5_req_wdata_ready <= 1'd0;
	main_sdram_bankmachine5_req_rdata_valid <= 1'd0;
	main_sdram_bankmachine5_refresh_gnt <= 1'd0;
	main_sdram_bankmachine5_cmd_valid <= 1'd0;
	builder_bankmachine5_next_state <= 3'd0;
	main_sdram_bankmachine5_row_open <= 1'd0;
	main_sdram_bankmachine5_row_close <= 1'd0;
	builder_bankmachine5_next_state <= builder_bankmachine5_state;
	case (builder_bankmachine5_state)
		1'd1: begin
			if ((main_sdram_bankmachine5_twtpcon_ready & main_sdram_bankmachine5_trascon_ready)) begin
				main_sdram_bankmachine5_cmd_valid <= 1'd1;
				if (main_sdram_bankmachine5_cmd_ready) begin
					builder_bankmachine5_next_state <= 3'd5;
				end
				main_sdram_bankmachine5_cmd_payload_ras <= 1'd1;
				main_sdram_bankmachine5_cmd_payload_we <= 1'd1;
				main_sdram_bankmachine5_cmd_payload_is_cmd <= 1'd1;
			end
			main_sdram_bankmachine5_row_close <= 1'd1;
		end
		2'd2: begin
			if ((main_sdram_bankmachine5_twtpcon_ready & main_sdram_bankmachine5_trascon_ready)) begin
				builder_bankmachine5_next_state <= 3'd5;
			end
			main_sdram_bankmachine5_row_close <= 1'd1;
		end
		2'd3: begin
			if (main_sdram_bankmachine5_trccon_ready) begin
				main_sdram_bankmachine5_row_col_n_addr_sel <= 1'd1;
				main_sdram_bankmachine5_row_open <= 1'd1;
				main_sdram_bankmachine5_cmd_valid <= 1'd1;
				main_sdram_bankmachine5_cmd_payload_is_cmd <= 1'd1;
				if (main_sdram_bankmachine5_cmd_ready) begin
					builder_bankmachine5_next_state <= 3'd6;
				end
				main_sdram_bankmachine5_cmd_payload_ras <= 1'd1;
			end
		end
		3'd4: begin
			if (main_sdram_bankmachine5_twtpcon_ready) begin
				main_sdram_bankmachine5_refresh_gnt <= 1'd1;
			end
			main_sdram_bankmachine5_row_close <= 1'd1;
			main_sdram_bankmachine5_cmd_payload_is_cmd <= 1'd1;
			if ((~main_sdram_bankmachine5_refresh_req)) begin
				builder_bankmachine5_next_state <= 1'd0;
			end
		end
		3'd5: begin
			builder_bankmachine5_next_state <= 2'd3;
		end
		3'd6: begin
			builder_bankmachine5_next_state <= 1'd0;
		end
		default: begin
			if (main_sdram_bankmachine5_refresh_req) begin
				builder_bankmachine5_next_state <= 3'd4;
			end else begin
				if (main_sdram_bankmachine5_cmd_buffer_source_valid) begin
					if (main_sdram_bankmachine5_row_opened) begin
						if (main_sdram_bankmachine5_row_hit) begin
							main_sdram_bankmachine5_cmd_valid <= 1'd1;
							if (main_sdram_bankmachine5_cmd_buffer_source_payload_we) begin
								main_sdram_bankmachine5_req_wdata_ready <= main_sdram_bankmachine5_cmd_ready;
								main_sdram_bankmachine5_cmd_payload_is_write <= 1'd1;
								main_sdram_bankmachine5_cmd_payload_we <= 1'd1;
							end else begin
								main_sdram_bankmachine5_req_rdata_valid <= main_sdram_bankmachine5_cmd_ready;
								main_sdram_bankmachine5_cmd_payload_is_read <= 1'd1;
							end
							main_sdram_bankmachine5_cmd_payload_cas <= 1'd1;
							if ((main_sdram_bankmachine5_cmd_ready & main_sdram_bankmachine5_auto_precharge)) begin
								builder_bankmachine5_next_state <= 2'd2;
							end
						end else begin
							builder_bankmachine5_next_state <= 1'd1;
						end
					end else begin
						builder_bankmachine5_next_state <= 2'd3;
					end
				end
			end
		end
	endcase
end
assign main_sdram_bankmachine6_cmd_buffer_lookahead_sink_valid = main_sdram_bankmachine6_req_valid;
assign main_sdram_bankmachine6_req_ready = main_sdram_bankmachine6_cmd_buffer_lookahead_sink_ready;
assign main_sdram_bankmachine6_cmd_buffer_lookahead_sink_payload_we = main_sdram_bankmachine6_req_we;
assign main_sdram_bankmachine6_cmd_buffer_lookahead_sink_payload_addr = main_sdram_bankmachine6_req_addr;
assign main_sdram_bankmachine6_cmd_buffer_sink_valid = main_sdram_bankmachine6_cmd_buffer_lookahead_source_valid;
assign main_sdram_bankmachine6_cmd_buffer_lookahead_source_ready = main_sdram_bankmachine6_cmd_buffer_sink_ready;
assign main_sdram_bankmachine6_cmd_buffer_sink_first = main_sdram_bankmachine6_cmd_buffer_lookahead_source_first;
assign main_sdram_bankmachine6_cmd_buffer_sink_last = main_sdram_bankmachine6_cmd_buffer_lookahead_source_last;
assign main_sdram_bankmachine6_cmd_buffer_sink_payload_we = main_sdram_bankmachine6_cmd_buffer_lookahead_source_payload_we;
assign main_sdram_bankmachine6_cmd_buffer_sink_payload_addr = main_sdram_bankmachine6_cmd_buffer_lookahead_source_payload_addr;
assign main_sdram_bankmachine6_cmd_buffer_source_ready = (main_sdram_bankmachine6_req_wdata_ready | main_sdram_bankmachine6_req_rdata_valid);
assign main_sdram_bankmachine6_req_lock = (main_sdram_bankmachine6_cmd_buffer_lookahead_source_valid | main_sdram_bankmachine6_cmd_buffer_source_valid);
assign main_sdram_bankmachine6_row_hit = (main_sdram_bankmachine6_row == main_sdram_bankmachine6_cmd_buffer_source_payload_addr[20:7]);
assign main_sdram_bankmachine6_cmd_payload_ba = 3'd6;
always @(*) begin
	main_sdram_bankmachine6_cmd_payload_a <= 14'd0;
	if (main_sdram_bankmachine6_row_col_n_addr_sel) begin
		main_sdram_bankmachine6_cmd_payload_a <= main_sdram_bankmachine6_cmd_buffer_source_payload_addr[20:7];
	end else begin
		main_sdram_bankmachine6_cmd_payload_a <= ((main_sdram_bankmachine6_auto_precharge <<< 4'd10) | {main_sdram_bankmachine6_cmd_buffer_source_payload_addr[6:0], {3{1'd0}}});
	end
end
assign main_sdram_bankmachine6_twtpcon_valid = ((main_sdram_bankmachine6_cmd_valid & main_sdram_bankmachine6_cmd_ready) & main_sdram_bankmachine6_cmd_payload_is_write);
assign main_sdram_bankmachine6_trccon_valid = ((main_sdram_bankmachine6_cmd_valid & main_sdram_bankmachine6_cmd_ready) & main_sdram_bankmachine6_row_open);
assign main_sdram_bankmachine6_trascon_valid = ((main_sdram_bankmachine6_cmd_valid & main_sdram_bankmachine6_cmd_ready) & main_sdram_bankmachine6_row_open);
always @(*) begin
	main_sdram_bankmachine6_auto_precharge <= 1'd0;
	if ((main_sdram_bankmachine6_cmd_buffer_lookahead_source_valid & main_sdram_bankmachine6_cmd_buffer_source_valid)) begin
		if ((main_sdram_bankmachine6_cmd_buffer_lookahead_source_payload_addr[20:7] != main_sdram_bankmachine6_cmd_buffer_source_payload_addr[20:7])) begin
			main_sdram_bankmachine6_auto_precharge <= (main_sdram_bankmachine6_row_close == 1'd0);
		end
	end
end
assign main_sdram_bankmachine6_cmd_buffer_lookahead_syncfifo6_din = {main_sdram_bankmachine6_cmd_buffer_lookahead_fifo_in_last, main_sdram_bankmachine6_cmd_buffer_lookahead_fifo_in_first, main_sdram_bankmachine6_cmd_buffer_lookahead_fifo_in_payload_addr, main_sdram_bankmachine6_cmd_buffer_lookahead_fifo_in_payload_we};
assign {main_sdram_bankmachine6_cmd_buffer_lookahead_fifo_out_last, main_sdram_bankmachine6_cmd_buffer_lookahead_fifo_out_first, main_sdram_bankmachine6_cmd_buffer_lookahead_fifo_out_payload_addr, main_sdram_bankmachine6_cmd_buffer_lookahead_fifo_out_payload_we} = main_sdram_bankmachine6_cmd_buffer_lookahead_syncfifo6_dout;
assign main_sdram_bankmachine6_cmd_buffer_lookahead_sink_ready = main_sdram_bankmachine6_cmd_buffer_lookahead_syncfifo6_writable;
assign main_sdram_bankmachine6_cmd_buffer_lookahead_syncfifo6_we = main_sdram_bankmachine6_cmd_buffer_lookahead_sink_valid;
assign main_sdram_bankmachine6_cmd_buffer_lookahead_fifo_in_first = main_sdram_bankmachine6_cmd_buffer_lookahead_sink_first;
assign main_sdram_bankmachine6_cmd_buffer_lookahead_fifo_in_last = main_sdram_bankmachine6_cmd_buffer_lookahead_sink_last;
assign main_sdram_bankmachine6_cmd_buffer_lookahead_fifo_in_payload_we = main_sdram_bankmachine6_cmd_buffer_lookahead_sink_payload_we;
assign main_sdram_bankmachine6_cmd_buffer_lookahead_fifo_in_payload_addr = main_sdram_bankmachine6_cmd_buffer_lookahead_sink_payload_addr;
assign main_sdram_bankmachine6_cmd_buffer_lookahead_source_valid = main_sdram_bankmachine6_cmd_buffer_lookahead_syncfifo6_readable;
assign main_sdram_bankmachine6_cmd_buffer_lookahead_source_first = main_sdram_bankmachine6_cmd_buffer_lookahead_fifo_out_first;
assign main_sdram_bankmachine6_cmd_buffer_lookahead_source_last = main_sdram_bankmachine6_cmd_buffer_lookahead_fifo_out_last;
assign main_sdram_bankmachine6_cmd_buffer_lookahead_source_payload_we = main_sdram_bankmachine6_cmd_buffer_lookahead_fifo_out_payload_we;
assign main_sdram_bankmachine6_cmd_buffer_lookahead_source_payload_addr = main_sdram_bankmachine6_cmd_buffer_lookahead_fifo_out_payload_addr;
assign main_sdram_bankmachine6_cmd_buffer_lookahead_syncfifo6_re = main_sdram_bankmachine6_cmd_buffer_lookahead_source_ready;
always @(*) begin
	main_sdram_bankmachine6_cmd_buffer_lookahead_wrport_adr <= 3'd0;
	if (main_sdram_bankmachine6_cmd_buffer_lookahead_replace) begin
		main_sdram_bankmachine6_cmd_buffer_lookahead_wrport_adr <= (main_sdram_bankmachine6_cmd_buffer_lookahead_produce - 1'd1);
	end else begin
		main_sdram_bankmachine6_cmd_buffer_lookahead_wrport_adr <= main_sdram_bankmachine6_cmd_buffer_lookahead_produce;
	end
end
assign main_sdram_bankmachine6_cmd_buffer_lookahead_wrport_dat_w = main_sdram_bankmachine6_cmd_buffer_lookahead_syncfifo6_din;
assign main_sdram_bankmachine6_cmd_buffer_lookahead_wrport_we = (main_sdram_bankmachine6_cmd_buffer_lookahead_syncfifo6_we & (main_sdram_bankmachine6_cmd_buffer_lookahead_syncfifo6_writable | main_sdram_bankmachine6_cmd_buffer_lookahead_replace));
assign main_sdram_bankmachine6_cmd_buffer_lookahead_do_read = (main_sdram_bankmachine6_cmd_buffer_lookahead_syncfifo6_readable & main_sdram_bankmachine6_cmd_buffer_lookahead_syncfifo6_re);
assign main_sdram_bankmachine6_cmd_buffer_lookahead_rdport_adr = main_sdram_bankmachine6_cmd_buffer_lookahead_consume;
assign main_sdram_bankmachine6_cmd_buffer_lookahead_syncfifo6_dout = main_sdram_bankmachine6_cmd_buffer_lookahead_rdport_dat_r;
assign main_sdram_bankmachine6_cmd_buffer_lookahead_syncfifo6_writable = (main_sdram_bankmachine6_cmd_buffer_lookahead_level != 4'd8);
assign main_sdram_bankmachine6_cmd_buffer_lookahead_syncfifo6_readable = (main_sdram_bankmachine6_cmd_buffer_lookahead_level != 1'd0);
assign main_sdram_bankmachine6_cmd_buffer_sink_ready = ((~main_sdram_bankmachine6_cmd_buffer_source_valid) | main_sdram_bankmachine6_cmd_buffer_source_ready);
always @(*) begin
	main_sdram_bankmachine6_cmd_payload_cas <= 1'd0;
	main_sdram_bankmachine6_cmd_payload_ras <= 1'd0;
	main_sdram_bankmachine6_cmd_payload_we <= 1'd0;
	main_sdram_bankmachine6_row_col_n_addr_sel <= 1'd0;
	main_sdram_bankmachine6_cmd_payload_is_cmd <= 1'd0;
	main_sdram_bankmachine6_cmd_payload_is_read <= 1'd0;
	main_sdram_bankmachine6_cmd_payload_is_write <= 1'd0;
	main_sdram_bankmachine6_req_wdata_ready <= 1'd0;
	main_sdram_bankmachine6_req_rdata_valid <= 1'd0;
	main_sdram_bankmachine6_refresh_gnt <= 1'd0;
	main_sdram_bankmachine6_cmd_valid <= 1'd0;
	builder_bankmachine6_next_state <= 3'd0;
	main_sdram_bankmachine6_row_open <= 1'd0;
	main_sdram_bankmachine6_row_close <= 1'd0;
	builder_bankmachine6_next_state <= builder_bankmachine6_state;
	case (builder_bankmachine6_state)
		1'd1: begin
			if ((main_sdram_bankmachine6_twtpcon_ready & main_sdram_bankmachine6_trascon_ready)) begin
				main_sdram_bankmachine6_cmd_valid <= 1'd1;
				if (main_sdram_bankmachine6_cmd_ready) begin
					builder_bankmachine6_next_state <= 3'd5;
				end
				main_sdram_bankmachine6_cmd_payload_ras <= 1'd1;
				main_sdram_bankmachine6_cmd_payload_we <= 1'd1;
				main_sdram_bankmachine6_cmd_payload_is_cmd <= 1'd1;
			end
			main_sdram_bankmachine6_row_close <= 1'd1;
		end
		2'd2: begin
			if ((main_sdram_bankmachine6_twtpcon_ready & main_sdram_bankmachine6_trascon_ready)) begin
				builder_bankmachine6_next_state <= 3'd5;
			end
			main_sdram_bankmachine6_row_close <= 1'd1;
		end
		2'd3: begin
			if (main_sdram_bankmachine6_trccon_ready) begin
				main_sdram_bankmachine6_row_col_n_addr_sel <= 1'd1;
				main_sdram_bankmachine6_row_open <= 1'd1;
				main_sdram_bankmachine6_cmd_valid <= 1'd1;
				main_sdram_bankmachine6_cmd_payload_is_cmd <= 1'd1;
				if (main_sdram_bankmachine6_cmd_ready) begin
					builder_bankmachine6_next_state <= 3'd6;
				end
				main_sdram_bankmachine6_cmd_payload_ras <= 1'd1;
			end
		end
		3'd4: begin
			if (main_sdram_bankmachine6_twtpcon_ready) begin
				main_sdram_bankmachine6_refresh_gnt <= 1'd1;
			end
			main_sdram_bankmachine6_row_close <= 1'd1;
			main_sdram_bankmachine6_cmd_payload_is_cmd <= 1'd1;
			if ((~main_sdram_bankmachine6_refresh_req)) begin
				builder_bankmachine6_next_state <= 1'd0;
			end
		end
		3'd5: begin
			builder_bankmachine6_next_state <= 2'd3;
		end
		3'd6: begin
			builder_bankmachine6_next_state <= 1'd0;
		end
		default: begin
			if (main_sdram_bankmachine6_refresh_req) begin
				builder_bankmachine6_next_state <= 3'd4;
			end else begin
				if (main_sdram_bankmachine6_cmd_buffer_source_valid) begin
					if (main_sdram_bankmachine6_row_opened) begin
						if (main_sdram_bankmachine6_row_hit) begin
							main_sdram_bankmachine6_cmd_valid <= 1'd1;
							if (main_sdram_bankmachine6_cmd_buffer_source_payload_we) begin
								main_sdram_bankmachine6_req_wdata_ready <= main_sdram_bankmachine6_cmd_ready;
								main_sdram_bankmachine6_cmd_payload_is_write <= 1'd1;
								main_sdram_bankmachine6_cmd_payload_we <= 1'd1;
							end else begin
								main_sdram_bankmachine6_req_rdata_valid <= main_sdram_bankmachine6_cmd_ready;
								main_sdram_bankmachine6_cmd_payload_is_read <= 1'd1;
							end
							main_sdram_bankmachine6_cmd_payload_cas <= 1'd1;
							if ((main_sdram_bankmachine6_cmd_ready & main_sdram_bankmachine6_auto_precharge)) begin
								builder_bankmachine6_next_state <= 2'd2;
							end
						end else begin
							builder_bankmachine6_next_state <= 1'd1;
						end
					end else begin
						builder_bankmachine6_next_state <= 2'd3;
					end
				end
			end
		end
	endcase
end
assign main_sdram_bankmachine7_cmd_buffer_lookahead_sink_valid = main_sdram_bankmachine7_req_valid;
assign main_sdram_bankmachine7_req_ready = main_sdram_bankmachine7_cmd_buffer_lookahead_sink_ready;
assign main_sdram_bankmachine7_cmd_buffer_lookahead_sink_payload_we = main_sdram_bankmachine7_req_we;
assign main_sdram_bankmachine7_cmd_buffer_lookahead_sink_payload_addr = main_sdram_bankmachine7_req_addr;
assign main_sdram_bankmachine7_cmd_buffer_sink_valid = main_sdram_bankmachine7_cmd_buffer_lookahead_source_valid;
assign main_sdram_bankmachine7_cmd_buffer_lookahead_source_ready = main_sdram_bankmachine7_cmd_buffer_sink_ready;
assign main_sdram_bankmachine7_cmd_buffer_sink_first = main_sdram_bankmachine7_cmd_buffer_lookahead_source_first;
assign main_sdram_bankmachine7_cmd_buffer_sink_last = main_sdram_bankmachine7_cmd_buffer_lookahead_source_last;
assign main_sdram_bankmachine7_cmd_buffer_sink_payload_we = main_sdram_bankmachine7_cmd_buffer_lookahead_source_payload_we;
assign main_sdram_bankmachine7_cmd_buffer_sink_payload_addr = main_sdram_bankmachine7_cmd_buffer_lookahead_source_payload_addr;
assign main_sdram_bankmachine7_cmd_buffer_source_ready = (main_sdram_bankmachine7_req_wdata_ready | main_sdram_bankmachine7_req_rdata_valid);
assign main_sdram_bankmachine7_req_lock = (main_sdram_bankmachine7_cmd_buffer_lookahead_source_valid | main_sdram_bankmachine7_cmd_buffer_source_valid);
assign main_sdram_bankmachine7_row_hit = (main_sdram_bankmachine7_row == main_sdram_bankmachine7_cmd_buffer_source_payload_addr[20:7]);
assign main_sdram_bankmachine7_cmd_payload_ba = 3'd7;
always @(*) begin
	main_sdram_bankmachine7_cmd_payload_a <= 14'd0;
	if (main_sdram_bankmachine7_row_col_n_addr_sel) begin
		main_sdram_bankmachine7_cmd_payload_a <= main_sdram_bankmachine7_cmd_buffer_source_payload_addr[20:7];
	end else begin
		main_sdram_bankmachine7_cmd_payload_a <= ((main_sdram_bankmachine7_auto_precharge <<< 4'd10) | {main_sdram_bankmachine7_cmd_buffer_source_payload_addr[6:0], {3{1'd0}}});
	end
end
assign main_sdram_bankmachine7_twtpcon_valid = ((main_sdram_bankmachine7_cmd_valid & main_sdram_bankmachine7_cmd_ready) & main_sdram_bankmachine7_cmd_payload_is_write);
assign main_sdram_bankmachine7_trccon_valid = ((main_sdram_bankmachine7_cmd_valid & main_sdram_bankmachine7_cmd_ready) & main_sdram_bankmachine7_row_open);
assign main_sdram_bankmachine7_trascon_valid = ((main_sdram_bankmachine7_cmd_valid & main_sdram_bankmachine7_cmd_ready) & main_sdram_bankmachine7_row_open);
always @(*) begin
	main_sdram_bankmachine7_auto_precharge <= 1'd0;
	if ((main_sdram_bankmachine7_cmd_buffer_lookahead_source_valid & main_sdram_bankmachine7_cmd_buffer_source_valid)) begin
		if ((main_sdram_bankmachine7_cmd_buffer_lookahead_source_payload_addr[20:7] != main_sdram_bankmachine7_cmd_buffer_source_payload_addr[20:7])) begin
			main_sdram_bankmachine7_auto_precharge <= (main_sdram_bankmachine7_row_close == 1'd0);
		end
	end
end
assign main_sdram_bankmachine7_cmd_buffer_lookahead_syncfifo7_din = {main_sdram_bankmachine7_cmd_buffer_lookahead_fifo_in_last, main_sdram_bankmachine7_cmd_buffer_lookahead_fifo_in_first, main_sdram_bankmachine7_cmd_buffer_lookahead_fifo_in_payload_addr, main_sdram_bankmachine7_cmd_buffer_lookahead_fifo_in_payload_we};
assign {main_sdram_bankmachine7_cmd_buffer_lookahead_fifo_out_last, main_sdram_bankmachine7_cmd_buffer_lookahead_fifo_out_first, main_sdram_bankmachine7_cmd_buffer_lookahead_fifo_out_payload_addr, main_sdram_bankmachine7_cmd_buffer_lookahead_fifo_out_payload_we} = main_sdram_bankmachine7_cmd_buffer_lookahead_syncfifo7_dout;
assign main_sdram_bankmachine7_cmd_buffer_lookahead_sink_ready = main_sdram_bankmachine7_cmd_buffer_lookahead_syncfifo7_writable;
assign main_sdram_bankmachine7_cmd_buffer_lookahead_syncfifo7_we = main_sdram_bankmachine7_cmd_buffer_lookahead_sink_valid;
assign main_sdram_bankmachine7_cmd_buffer_lookahead_fifo_in_first = main_sdram_bankmachine7_cmd_buffer_lookahead_sink_first;
assign main_sdram_bankmachine7_cmd_buffer_lookahead_fifo_in_last = main_sdram_bankmachine7_cmd_buffer_lookahead_sink_last;
assign main_sdram_bankmachine7_cmd_buffer_lookahead_fifo_in_payload_we = main_sdram_bankmachine7_cmd_buffer_lookahead_sink_payload_we;
assign main_sdram_bankmachine7_cmd_buffer_lookahead_fifo_in_payload_addr = main_sdram_bankmachine7_cmd_buffer_lookahead_sink_payload_addr;
assign main_sdram_bankmachine7_cmd_buffer_lookahead_source_valid = main_sdram_bankmachine7_cmd_buffer_lookahead_syncfifo7_readable;
assign main_sdram_bankmachine7_cmd_buffer_lookahead_source_first = main_sdram_bankmachine7_cmd_buffer_lookahead_fifo_out_first;
assign main_sdram_bankmachine7_cmd_buffer_lookahead_source_last = main_sdram_bankmachine7_cmd_buffer_lookahead_fifo_out_last;
assign main_sdram_bankmachine7_cmd_buffer_lookahead_source_payload_we = main_sdram_bankmachine7_cmd_buffer_lookahead_fifo_out_payload_we;
assign main_sdram_bankmachine7_cmd_buffer_lookahead_source_payload_addr = main_sdram_bankmachine7_cmd_buffer_lookahead_fifo_out_payload_addr;
assign main_sdram_bankmachine7_cmd_buffer_lookahead_syncfifo7_re = main_sdram_bankmachine7_cmd_buffer_lookahead_source_ready;
always @(*) begin
	main_sdram_bankmachine7_cmd_buffer_lookahead_wrport_adr <= 3'd0;
	if (main_sdram_bankmachine7_cmd_buffer_lookahead_replace) begin
		main_sdram_bankmachine7_cmd_buffer_lookahead_wrport_adr <= (main_sdram_bankmachine7_cmd_buffer_lookahead_produce - 1'd1);
	end else begin
		main_sdram_bankmachine7_cmd_buffer_lookahead_wrport_adr <= main_sdram_bankmachine7_cmd_buffer_lookahead_produce;
	end
end
assign main_sdram_bankmachine7_cmd_buffer_lookahead_wrport_dat_w = main_sdram_bankmachine7_cmd_buffer_lookahead_syncfifo7_din;
assign main_sdram_bankmachine7_cmd_buffer_lookahead_wrport_we = (main_sdram_bankmachine7_cmd_buffer_lookahead_syncfifo7_we & (main_sdram_bankmachine7_cmd_buffer_lookahead_syncfifo7_writable | main_sdram_bankmachine7_cmd_buffer_lookahead_replace));
assign main_sdram_bankmachine7_cmd_buffer_lookahead_do_read = (main_sdram_bankmachine7_cmd_buffer_lookahead_syncfifo7_readable & main_sdram_bankmachine7_cmd_buffer_lookahead_syncfifo7_re);
assign main_sdram_bankmachine7_cmd_buffer_lookahead_rdport_adr = main_sdram_bankmachine7_cmd_buffer_lookahead_consume;
assign main_sdram_bankmachine7_cmd_buffer_lookahead_syncfifo7_dout = main_sdram_bankmachine7_cmd_buffer_lookahead_rdport_dat_r;
assign main_sdram_bankmachine7_cmd_buffer_lookahead_syncfifo7_writable = (main_sdram_bankmachine7_cmd_buffer_lookahead_level != 4'd8);
assign main_sdram_bankmachine7_cmd_buffer_lookahead_syncfifo7_readable = (main_sdram_bankmachine7_cmd_buffer_lookahead_level != 1'd0);
assign main_sdram_bankmachine7_cmd_buffer_sink_ready = ((~main_sdram_bankmachine7_cmd_buffer_source_valid) | main_sdram_bankmachine7_cmd_buffer_source_ready);
always @(*) begin
	main_sdram_bankmachine7_cmd_payload_cas <= 1'd0;
	main_sdram_bankmachine7_cmd_payload_ras <= 1'd0;
	main_sdram_bankmachine7_cmd_payload_we <= 1'd0;
	main_sdram_bankmachine7_row_col_n_addr_sel <= 1'd0;
	main_sdram_bankmachine7_cmd_payload_is_cmd <= 1'd0;
	main_sdram_bankmachine7_cmd_payload_is_read <= 1'd0;
	main_sdram_bankmachine7_cmd_payload_is_write <= 1'd0;
	main_sdram_bankmachine7_req_wdata_ready <= 1'd0;
	main_sdram_bankmachine7_req_rdata_valid <= 1'd0;
	builder_bankmachine7_next_state <= 3'd0;
	main_sdram_bankmachine7_refresh_gnt <= 1'd0;
	main_sdram_bankmachine7_cmd_valid <= 1'd0;
	main_sdram_bankmachine7_row_open <= 1'd0;
	main_sdram_bankmachine7_row_close <= 1'd0;
	builder_bankmachine7_next_state <= builder_bankmachine7_state;
	case (builder_bankmachine7_state)
		1'd1: begin
			if ((main_sdram_bankmachine7_twtpcon_ready & main_sdram_bankmachine7_trascon_ready)) begin
				main_sdram_bankmachine7_cmd_valid <= 1'd1;
				if (main_sdram_bankmachine7_cmd_ready) begin
					builder_bankmachine7_next_state <= 3'd5;
				end
				main_sdram_bankmachine7_cmd_payload_ras <= 1'd1;
				main_sdram_bankmachine7_cmd_payload_we <= 1'd1;
				main_sdram_bankmachine7_cmd_payload_is_cmd <= 1'd1;
			end
			main_sdram_bankmachine7_row_close <= 1'd1;
		end
		2'd2: begin
			if ((main_sdram_bankmachine7_twtpcon_ready & main_sdram_bankmachine7_trascon_ready)) begin
				builder_bankmachine7_next_state <= 3'd5;
			end
			main_sdram_bankmachine7_row_close <= 1'd1;
		end
		2'd3: begin
			if (main_sdram_bankmachine7_trccon_ready) begin
				main_sdram_bankmachine7_row_col_n_addr_sel <= 1'd1;
				main_sdram_bankmachine7_row_open <= 1'd1;
				main_sdram_bankmachine7_cmd_valid <= 1'd1;
				main_sdram_bankmachine7_cmd_payload_is_cmd <= 1'd1;
				if (main_sdram_bankmachine7_cmd_ready) begin
					builder_bankmachine7_next_state <= 3'd6;
				end
				main_sdram_bankmachine7_cmd_payload_ras <= 1'd1;
			end
		end
		3'd4: begin
			if (main_sdram_bankmachine7_twtpcon_ready) begin
				main_sdram_bankmachine7_refresh_gnt <= 1'd1;
			end
			main_sdram_bankmachine7_row_close <= 1'd1;
			main_sdram_bankmachine7_cmd_payload_is_cmd <= 1'd1;
			if ((~main_sdram_bankmachine7_refresh_req)) begin
				builder_bankmachine7_next_state <= 1'd0;
			end
		end
		3'd5: begin
			builder_bankmachine7_next_state <= 2'd3;
		end
		3'd6: begin
			builder_bankmachine7_next_state <= 1'd0;
		end
		default: begin
			if (main_sdram_bankmachine7_refresh_req) begin
				builder_bankmachine7_next_state <= 3'd4;
			end else begin
				if (main_sdram_bankmachine7_cmd_buffer_source_valid) begin
					if (main_sdram_bankmachine7_row_opened) begin
						if (main_sdram_bankmachine7_row_hit) begin
							main_sdram_bankmachine7_cmd_valid <= 1'd1;
							if (main_sdram_bankmachine7_cmd_buffer_source_payload_we) begin
								main_sdram_bankmachine7_req_wdata_ready <= main_sdram_bankmachine7_cmd_ready;
								main_sdram_bankmachine7_cmd_payload_is_write <= 1'd1;
								main_sdram_bankmachine7_cmd_payload_we <= 1'd1;
							end else begin
								main_sdram_bankmachine7_req_rdata_valid <= main_sdram_bankmachine7_cmd_ready;
								main_sdram_bankmachine7_cmd_payload_is_read <= 1'd1;
							end
							main_sdram_bankmachine7_cmd_payload_cas <= 1'd1;
							if ((main_sdram_bankmachine7_cmd_ready & main_sdram_bankmachine7_auto_precharge)) begin
								builder_bankmachine7_next_state <= 2'd2;
							end
						end else begin
							builder_bankmachine7_next_state <= 1'd1;
						end
					end else begin
						builder_bankmachine7_next_state <= 2'd3;
					end
				end
			end
		end
	endcase
end
assign main_sdram_trrdcon_valid = ((main_sdram_choose_cmd_cmd_valid & main_sdram_choose_cmd_cmd_ready) & ((main_sdram_choose_cmd_cmd_payload_ras & (~main_sdram_choose_cmd_cmd_payload_cas)) & (~main_sdram_choose_cmd_cmd_payload_we)));
assign main_sdram_tfawcon_valid = ((main_sdram_choose_cmd_cmd_valid & main_sdram_choose_cmd_cmd_ready) & ((main_sdram_choose_cmd_cmd_payload_ras & (~main_sdram_choose_cmd_cmd_payload_cas)) & (~main_sdram_choose_cmd_cmd_payload_we)));
assign main_sdram_ras_allowed = (main_sdram_trrdcon_ready & main_sdram_tfawcon_ready);
assign main_sdram_tccdcon_valid = ((main_sdram_choose_req_cmd_valid & main_sdram_choose_req_cmd_ready) & (main_sdram_choose_req_cmd_payload_is_write | main_sdram_choose_req_cmd_payload_is_read));
assign main_sdram_cas_allowed = main_sdram_tccdcon_ready;
assign main_sdram_twtrcon_valid = ((main_sdram_choose_req_cmd_valid & main_sdram_choose_req_cmd_ready) & main_sdram_choose_req_cmd_payload_is_write);
assign main_sdram_read_available = ((((((((main_sdram_bankmachine0_cmd_valid & main_sdram_bankmachine0_cmd_payload_is_read) | (main_sdram_bankmachine1_cmd_valid & main_sdram_bankmachine1_cmd_payload_is_read)) | (main_sdram_bankmachine2_cmd_valid & main_sdram_bankmachine2_cmd_payload_is_read)) | (main_sdram_bankmachine3_cmd_valid & main_sdram_bankmachine3_cmd_payload_is_read)) | (main_sdram_bankmachine4_cmd_valid & main_sdram_bankmachine4_cmd_payload_is_read)) | (main_sdram_bankmachine5_cmd_valid & main_sdram_bankmachine5_cmd_payload_is_read)) | (main_sdram_bankmachine6_cmd_valid & main_sdram_bankmachine6_cmd_payload_is_read)) | (main_sdram_bankmachine7_cmd_valid & main_sdram_bankmachine7_cmd_payload_is_read));
assign main_sdram_write_available = ((((((((main_sdram_bankmachine0_cmd_valid & main_sdram_bankmachine0_cmd_payload_is_write) | (main_sdram_bankmachine1_cmd_valid & main_sdram_bankmachine1_cmd_payload_is_write)) | (main_sdram_bankmachine2_cmd_valid & main_sdram_bankmachine2_cmd_payload_is_write)) | (main_sdram_bankmachine3_cmd_valid & main_sdram_bankmachine3_cmd_payload_is_write)) | (main_sdram_bankmachine4_cmd_valid & main_sdram_bankmachine4_cmd_payload_is_write)) | (main_sdram_bankmachine5_cmd_valid & main_sdram_bankmachine5_cmd_payload_is_write)) | (main_sdram_bankmachine6_cmd_valid & main_sdram_bankmachine6_cmd_payload_is_write)) | (main_sdram_bankmachine7_cmd_valid & main_sdram_bankmachine7_cmd_payload_is_write));
assign main_sdram_max_time0 = (main_sdram_time0 == 1'd0);
assign main_sdram_max_time1 = (main_sdram_time1 == 1'd0);
assign main_sdram_bankmachine0_refresh_req = main_sdram_cmd_valid;
assign main_sdram_bankmachine1_refresh_req = main_sdram_cmd_valid;
assign main_sdram_bankmachine2_refresh_req = main_sdram_cmd_valid;
assign main_sdram_bankmachine3_refresh_req = main_sdram_cmd_valid;
assign main_sdram_bankmachine4_refresh_req = main_sdram_cmd_valid;
assign main_sdram_bankmachine5_refresh_req = main_sdram_cmd_valid;
assign main_sdram_bankmachine6_refresh_req = main_sdram_cmd_valid;
assign main_sdram_bankmachine7_refresh_req = main_sdram_cmd_valid;
assign main_sdram_go_to_refresh = (((((((main_sdram_bankmachine0_refresh_gnt & main_sdram_bankmachine1_refresh_gnt) & main_sdram_bankmachine2_refresh_gnt) & main_sdram_bankmachine3_refresh_gnt) & main_sdram_bankmachine4_refresh_gnt) & main_sdram_bankmachine5_refresh_gnt) & main_sdram_bankmachine6_refresh_gnt) & main_sdram_bankmachine7_refresh_gnt);
assign main_sdram_interface_rdata = {main_sdram_dfi_p3_rddata, main_sdram_dfi_p2_rddata, main_sdram_dfi_p1_rddata, main_sdram_dfi_p0_rddata};
assign {main_sdram_dfi_p3_wrdata, main_sdram_dfi_p2_wrdata, main_sdram_dfi_p1_wrdata, main_sdram_dfi_p0_wrdata} = main_sdram_interface_wdata;
assign {main_sdram_dfi_p3_wrdata_mask, main_sdram_dfi_p2_wrdata_mask, main_sdram_dfi_p1_wrdata_mask, main_sdram_dfi_p0_wrdata_mask} = (~main_sdram_interface_wdata_we);
always @(*) begin
	main_sdram_choose_cmd_valids <= 8'd0;
	main_sdram_choose_cmd_valids[0] <= (main_sdram_bankmachine0_cmd_valid & (((main_sdram_bankmachine0_cmd_payload_is_cmd & main_sdram_choose_cmd_want_cmds) & ((~((main_sdram_bankmachine0_cmd_payload_ras & (~main_sdram_bankmachine0_cmd_payload_cas)) & (~main_sdram_bankmachine0_cmd_payload_we))) | main_sdram_choose_cmd_want_activates)) | ((main_sdram_bankmachine0_cmd_payload_is_read == main_sdram_choose_cmd_want_reads) & (main_sdram_bankmachine0_cmd_payload_is_write == main_sdram_choose_cmd_want_writes))));
	main_sdram_choose_cmd_valids[1] <= (main_sdram_bankmachine1_cmd_valid & (((main_sdram_bankmachine1_cmd_payload_is_cmd & main_sdram_choose_cmd_want_cmds) & ((~((main_sdram_bankmachine1_cmd_payload_ras & (~main_sdram_bankmachine1_cmd_payload_cas)) & (~main_sdram_bankmachine1_cmd_payload_we))) | main_sdram_choose_cmd_want_activates)) | ((main_sdram_bankmachine1_cmd_payload_is_read == main_sdram_choose_cmd_want_reads) & (main_sdram_bankmachine1_cmd_payload_is_write == main_sdram_choose_cmd_want_writes))));
	main_sdram_choose_cmd_valids[2] <= (main_sdram_bankmachine2_cmd_valid & (((main_sdram_bankmachine2_cmd_payload_is_cmd & main_sdram_choose_cmd_want_cmds) & ((~((main_sdram_bankmachine2_cmd_payload_ras & (~main_sdram_bankmachine2_cmd_payload_cas)) & (~main_sdram_bankmachine2_cmd_payload_we))) | main_sdram_choose_cmd_want_activates)) | ((main_sdram_bankmachine2_cmd_payload_is_read == main_sdram_choose_cmd_want_reads) & (main_sdram_bankmachine2_cmd_payload_is_write == main_sdram_choose_cmd_want_writes))));
	main_sdram_choose_cmd_valids[3] <= (main_sdram_bankmachine3_cmd_valid & (((main_sdram_bankmachine3_cmd_payload_is_cmd & main_sdram_choose_cmd_want_cmds) & ((~((main_sdram_bankmachine3_cmd_payload_ras & (~main_sdram_bankmachine3_cmd_payload_cas)) & (~main_sdram_bankmachine3_cmd_payload_we))) | main_sdram_choose_cmd_want_activates)) | ((main_sdram_bankmachine3_cmd_payload_is_read == main_sdram_choose_cmd_want_reads) & (main_sdram_bankmachine3_cmd_payload_is_write == main_sdram_choose_cmd_want_writes))));
	main_sdram_choose_cmd_valids[4] <= (main_sdram_bankmachine4_cmd_valid & (((main_sdram_bankmachine4_cmd_payload_is_cmd & main_sdram_choose_cmd_want_cmds) & ((~((main_sdram_bankmachine4_cmd_payload_ras & (~main_sdram_bankmachine4_cmd_payload_cas)) & (~main_sdram_bankmachine4_cmd_payload_we))) | main_sdram_choose_cmd_want_activates)) | ((main_sdram_bankmachine4_cmd_payload_is_read == main_sdram_choose_cmd_want_reads) & (main_sdram_bankmachine4_cmd_payload_is_write == main_sdram_choose_cmd_want_writes))));
	main_sdram_choose_cmd_valids[5] <= (main_sdram_bankmachine5_cmd_valid & (((main_sdram_bankmachine5_cmd_payload_is_cmd & main_sdram_choose_cmd_want_cmds) & ((~((main_sdram_bankmachine5_cmd_payload_ras & (~main_sdram_bankmachine5_cmd_payload_cas)) & (~main_sdram_bankmachine5_cmd_payload_we))) | main_sdram_choose_cmd_want_activates)) | ((main_sdram_bankmachine5_cmd_payload_is_read == main_sdram_choose_cmd_want_reads) & (main_sdram_bankmachine5_cmd_payload_is_write == main_sdram_choose_cmd_want_writes))));
	main_sdram_choose_cmd_valids[6] <= (main_sdram_bankmachine6_cmd_valid & (((main_sdram_bankmachine6_cmd_payload_is_cmd & main_sdram_choose_cmd_want_cmds) & ((~((main_sdram_bankmachine6_cmd_payload_ras & (~main_sdram_bankmachine6_cmd_payload_cas)) & (~main_sdram_bankmachine6_cmd_payload_we))) | main_sdram_choose_cmd_want_activates)) | ((main_sdram_bankmachine6_cmd_payload_is_read == main_sdram_choose_cmd_want_reads) & (main_sdram_bankmachine6_cmd_payload_is_write == main_sdram_choose_cmd_want_writes))));
	main_sdram_choose_cmd_valids[7] <= (main_sdram_bankmachine7_cmd_valid & (((main_sdram_bankmachine7_cmd_payload_is_cmd & main_sdram_choose_cmd_want_cmds) & ((~((main_sdram_bankmachine7_cmd_payload_ras & (~main_sdram_bankmachine7_cmd_payload_cas)) & (~main_sdram_bankmachine7_cmd_payload_we))) | main_sdram_choose_cmd_want_activates)) | ((main_sdram_bankmachine7_cmd_payload_is_read == main_sdram_choose_cmd_want_reads) & (main_sdram_bankmachine7_cmd_payload_is_write == main_sdram_choose_cmd_want_writes))));
end
assign main_sdram_choose_cmd_request = main_sdram_choose_cmd_valids;
assign main_sdram_choose_cmd_cmd_valid = builder_rhs_array_muxed0;
assign main_sdram_choose_cmd_cmd_payload_a = builder_rhs_array_muxed1;
assign main_sdram_choose_cmd_cmd_payload_ba = builder_rhs_array_muxed2;
assign main_sdram_choose_cmd_cmd_payload_is_read = builder_rhs_array_muxed3;
assign main_sdram_choose_cmd_cmd_payload_is_write = builder_rhs_array_muxed4;
assign main_sdram_choose_cmd_cmd_payload_is_cmd = builder_rhs_array_muxed5;
always @(*) begin
	main_sdram_choose_cmd_cmd_payload_cas <= 1'd0;
	if (main_sdram_choose_cmd_cmd_valid) begin
		main_sdram_choose_cmd_cmd_payload_cas <= builder_t_array_muxed0;
	end
end
always @(*) begin
	main_sdram_choose_cmd_cmd_payload_ras <= 1'd0;
	if (main_sdram_choose_cmd_cmd_valid) begin
		main_sdram_choose_cmd_cmd_payload_ras <= builder_t_array_muxed1;
	end
end
always @(*) begin
	main_sdram_choose_cmd_cmd_payload_we <= 1'd0;
	if (main_sdram_choose_cmd_cmd_valid) begin
		main_sdram_choose_cmd_cmd_payload_we <= builder_t_array_muxed2;
	end
end
assign main_sdram_choose_cmd_ce = (main_sdram_choose_cmd_cmd_ready | (~main_sdram_choose_cmd_cmd_valid));
always @(*) begin
	main_sdram_choose_req_valids <= 8'd0;
	main_sdram_choose_req_valids[0] <= (main_sdram_bankmachine0_cmd_valid & (((main_sdram_bankmachine0_cmd_payload_is_cmd & main_sdram_choose_req_want_cmds) & ((~((main_sdram_bankmachine0_cmd_payload_ras & (~main_sdram_bankmachine0_cmd_payload_cas)) & (~main_sdram_bankmachine0_cmd_payload_we))) | main_sdram_choose_req_want_activates)) | ((main_sdram_bankmachine0_cmd_payload_is_read == main_sdram_choose_req_want_reads) & (main_sdram_bankmachine0_cmd_payload_is_write == main_sdram_choose_req_want_writes))));
	main_sdram_choose_req_valids[1] <= (main_sdram_bankmachine1_cmd_valid & (((main_sdram_bankmachine1_cmd_payload_is_cmd & main_sdram_choose_req_want_cmds) & ((~((main_sdram_bankmachine1_cmd_payload_ras & (~main_sdram_bankmachine1_cmd_payload_cas)) & (~main_sdram_bankmachine1_cmd_payload_we))) | main_sdram_choose_req_want_activates)) | ((main_sdram_bankmachine1_cmd_payload_is_read == main_sdram_choose_req_want_reads) & (main_sdram_bankmachine1_cmd_payload_is_write == main_sdram_choose_req_want_writes))));
	main_sdram_choose_req_valids[2] <= (main_sdram_bankmachine2_cmd_valid & (((main_sdram_bankmachine2_cmd_payload_is_cmd & main_sdram_choose_req_want_cmds) & ((~((main_sdram_bankmachine2_cmd_payload_ras & (~main_sdram_bankmachine2_cmd_payload_cas)) & (~main_sdram_bankmachine2_cmd_payload_we))) | main_sdram_choose_req_want_activates)) | ((main_sdram_bankmachine2_cmd_payload_is_read == main_sdram_choose_req_want_reads) & (main_sdram_bankmachine2_cmd_payload_is_write == main_sdram_choose_req_want_writes))));
	main_sdram_choose_req_valids[3] <= (main_sdram_bankmachine3_cmd_valid & (((main_sdram_bankmachine3_cmd_payload_is_cmd & main_sdram_choose_req_want_cmds) & ((~((main_sdram_bankmachine3_cmd_payload_ras & (~main_sdram_bankmachine3_cmd_payload_cas)) & (~main_sdram_bankmachine3_cmd_payload_we))) | main_sdram_choose_req_want_activates)) | ((main_sdram_bankmachine3_cmd_payload_is_read == main_sdram_choose_req_want_reads) & (main_sdram_bankmachine3_cmd_payload_is_write == main_sdram_choose_req_want_writes))));
	main_sdram_choose_req_valids[4] <= (main_sdram_bankmachine4_cmd_valid & (((main_sdram_bankmachine4_cmd_payload_is_cmd & main_sdram_choose_req_want_cmds) & ((~((main_sdram_bankmachine4_cmd_payload_ras & (~main_sdram_bankmachine4_cmd_payload_cas)) & (~main_sdram_bankmachine4_cmd_payload_we))) | main_sdram_choose_req_want_activates)) | ((main_sdram_bankmachine4_cmd_payload_is_read == main_sdram_choose_req_want_reads) & (main_sdram_bankmachine4_cmd_payload_is_write == main_sdram_choose_req_want_writes))));
	main_sdram_choose_req_valids[5] <= (main_sdram_bankmachine5_cmd_valid & (((main_sdram_bankmachine5_cmd_payload_is_cmd & main_sdram_choose_req_want_cmds) & ((~((main_sdram_bankmachine5_cmd_payload_ras & (~main_sdram_bankmachine5_cmd_payload_cas)) & (~main_sdram_bankmachine5_cmd_payload_we))) | main_sdram_choose_req_want_activates)) | ((main_sdram_bankmachine5_cmd_payload_is_read == main_sdram_choose_req_want_reads) & (main_sdram_bankmachine5_cmd_payload_is_write == main_sdram_choose_req_want_writes))));
	main_sdram_choose_req_valids[6] <= (main_sdram_bankmachine6_cmd_valid & (((main_sdram_bankmachine6_cmd_payload_is_cmd & main_sdram_choose_req_want_cmds) & ((~((main_sdram_bankmachine6_cmd_payload_ras & (~main_sdram_bankmachine6_cmd_payload_cas)) & (~main_sdram_bankmachine6_cmd_payload_we))) | main_sdram_choose_req_want_activates)) | ((main_sdram_bankmachine6_cmd_payload_is_read == main_sdram_choose_req_want_reads) & (main_sdram_bankmachine6_cmd_payload_is_write == main_sdram_choose_req_want_writes))));
	main_sdram_choose_req_valids[7] <= (main_sdram_bankmachine7_cmd_valid & (((main_sdram_bankmachine7_cmd_payload_is_cmd & main_sdram_choose_req_want_cmds) & ((~((main_sdram_bankmachine7_cmd_payload_ras & (~main_sdram_bankmachine7_cmd_payload_cas)) & (~main_sdram_bankmachine7_cmd_payload_we))) | main_sdram_choose_req_want_activates)) | ((main_sdram_bankmachine7_cmd_payload_is_read == main_sdram_choose_req_want_reads) & (main_sdram_bankmachine7_cmd_payload_is_write == main_sdram_choose_req_want_writes))));
end
assign main_sdram_choose_req_request = main_sdram_choose_req_valids;
assign main_sdram_choose_req_cmd_valid = builder_rhs_array_muxed6;
assign main_sdram_choose_req_cmd_payload_a = builder_rhs_array_muxed7;
assign main_sdram_choose_req_cmd_payload_ba = builder_rhs_array_muxed8;
assign main_sdram_choose_req_cmd_payload_is_read = builder_rhs_array_muxed9;
assign main_sdram_choose_req_cmd_payload_is_write = builder_rhs_array_muxed10;
assign main_sdram_choose_req_cmd_payload_is_cmd = builder_rhs_array_muxed11;
always @(*) begin
	main_sdram_choose_req_cmd_payload_cas <= 1'd0;
	if (main_sdram_choose_req_cmd_valid) begin
		main_sdram_choose_req_cmd_payload_cas <= builder_t_array_muxed3;
	end
end
always @(*) begin
	main_sdram_choose_req_cmd_payload_ras <= 1'd0;
	if (main_sdram_choose_req_cmd_valid) begin
		main_sdram_choose_req_cmd_payload_ras <= builder_t_array_muxed4;
	end
end
always @(*) begin
	main_sdram_choose_req_cmd_payload_we <= 1'd0;
	if (main_sdram_choose_req_cmd_valid) begin
		main_sdram_choose_req_cmd_payload_we <= builder_t_array_muxed5;
	end
end
always @(*) begin
	main_sdram_bankmachine0_cmd_ready <= 1'd0;
	if (((main_sdram_choose_cmd_cmd_valid & main_sdram_choose_cmd_cmd_ready) & (main_sdram_choose_cmd_grant == 1'd0))) begin
		main_sdram_bankmachine0_cmd_ready <= 1'd1;
	end
	if (((main_sdram_choose_req_cmd_valid & main_sdram_choose_req_cmd_ready) & (main_sdram_choose_req_grant == 1'd0))) begin
		main_sdram_bankmachine0_cmd_ready <= 1'd1;
	end
end
always @(*) begin
	main_sdram_bankmachine1_cmd_ready <= 1'd0;
	if (((main_sdram_choose_cmd_cmd_valid & main_sdram_choose_cmd_cmd_ready) & (main_sdram_choose_cmd_grant == 1'd1))) begin
		main_sdram_bankmachine1_cmd_ready <= 1'd1;
	end
	if (((main_sdram_choose_req_cmd_valid & main_sdram_choose_req_cmd_ready) & (main_sdram_choose_req_grant == 1'd1))) begin
		main_sdram_bankmachine1_cmd_ready <= 1'd1;
	end
end
always @(*) begin
	main_sdram_bankmachine2_cmd_ready <= 1'd0;
	if (((main_sdram_choose_cmd_cmd_valid & main_sdram_choose_cmd_cmd_ready) & (main_sdram_choose_cmd_grant == 2'd2))) begin
		main_sdram_bankmachine2_cmd_ready <= 1'd1;
	end
	if (((main_sdram_choose_req_cmd_valid & main_sdram_choose_req_cmd_ready) & (main_sdram_choose_req_grant == 2'd2))) begin
		main_sdram_bankmachine2_cmd_ready <= 1'd1;
	end
end
always @(*) begin
	main_sdram_bankmachine3_cmd_ready <= 1'd0;
	if (((main_sdram_choose_cmd_cmd_valid & main_sdram_choose_cmd_cmd_ready) & (main_sdram_choose_cmd_grant == 2'd3))) begin
		main_sdram_bankmachine3_cmd_ready <= 1'd1;
	end
	if (((main_sdram_choose_req_cmd_valid & main_sdram_choose_req_cmd_ready) & (main_sdram_choose_req_grant == 2'd3))) begin
		main_sdram_bankmachine3_cmd_ready <= 1'd1;
	end
end
always @(*) begin
	main_sdram_bankmachine4_cmd_ready <= 1'd0;
	if (((main_sdram_choose_cmd_cmd_valid & main_sdram_choose_cmd_cmd_ready) & (main_sdram_choose_cmd_grant == 3'd4))) begin
		main_sdram_bankmachine4_cmd_ready <= 1'd1;
	end
	if (((main_sdram_choose_req_cmd_valid & main_sdram_choose_req_cmd_ready) & (main_sdram_choose_req_grant == 3'd4))) begin
		main_sdram_bankmachine4_cmd_ready <= 1'd1;
	end
end
always @(*) begin
	main_sdram_bankmachine5_cmd_ready <= 1'd0;
	if (((main_sdram_choose_cmd_cmd_valid & main_sdram_choose_cmd_cmd_ready) & (main_sdram_choose_cmd_grant == 3'd5))) begin
		main_sdram_bankmachine5_cmd_ready <= 1'd1;
	end
	if (((main_sdram_choose_req_cmd_valid & main_sdram_choose_req_cmd_ready) & (main_sdram_choose_req_grant == 3'd5))) begin
		main_sdram_bankmachine5_cmd_ready <= 1'd1;
	end
end
always @(*) begin
	main_sdram_bankmachine6_cmd_ready <= 1'd0;
	if (((main_sdram_choose_cmd_cmd_valid & main_sdram_choose_cmd_cmd_ready) & (main_sdram_choose_cmd_grant == 3'd6))) begin
		main_sdram_bankmachine6_cmd_ready <= 1'd1;
	end
	if (((main_sdram_choose_req_cmd_valid & main_sdram_choose_req_cmd_ready) & (main_sdram_choose_req_grant == 3'd6))) begin
		main_sdram_bankmachine6_cmd_ready <= 1'd1;
	end
end
always @(*) begin
	main_sdram_bankmachine7_cmd_ready <= 1'd0;
	if (((main_sdram_choose_cmd_cmd_valid & main_sdram_choose_cmd_cmd_ready) & (main_sdram_choose_cmd_grant == 3'd7))) begin
		main_sdram_bankmachine7_cmd_ready <= 1'd1;
	end
	if (((main_sdram_choose_req_cmd_valid & main_sdram_choose_req_cmd_ready) & (main_sdram_choose_req_grant == 3'd7))) begin
		main_sdram_bankmachine7_cmd_ready <= 1'd1;
	end
end
assign main_sdram_choose_req_ce = (main_sdram_choose_req_cmd_ready | (~main_sdram_choose_req_cmd_valid));
assign main_sdram_dfi_p0_reset_n = 1'd1;
assign main_sdram_dfi_p0_cke = {1{main_sdram_steerer0}};
assign main_sdram_dfi_p0_odt = {1{main_sdram_steerer1}};
assign main_sdram_dfi_p1_reset_n = 1'd1;
assign main_sdram_dfi_p1_cke = {1{main_sdram_steerer2}};
assign main_sdram_dfi_p1_odt = {1{main_sdram_steerer3}};
assign main_sdram_dfi_p2_reset_n = 1'd1;
assign main_sdram_dfi_p2_cke = {1{main_sdram_steerer4}};
assign main_sdram_dfi_p2_odt = {1{main_sdram_steerer5}};
assign main_sdram_dfi_p3_reset_n = 1'd1;
assign main_sdram_dfi_p3_cke = {1{main_sdram_steerer6}};
assign main_sdram_dfi_p3_odt = {1{main_sdram_steerer7}};
assign main_sdram_tfawcon_count = ((main_sdram_tfawcon_window[0] + main_sdram_tfawcon_window[1]) + main_sdram_tfawcon_window[2]);
always @(*) begin
	main_sdram_steerer_sel0 <= 2'd0;
	main_sdram_steerer_sel1 <= 2'd0;
	main_sdram_en0 <= 1'd0;
	main_sdram_steerer_sel2 <= 2'd0;
	main_sdram_choose_cmd_want_activates <= 1'd0;
	main_sdram_steerer_sel3 <= 2'd0;
	builder_multiplexer_next_state <= 4'd0;
	main_sdram_cmd_ready <= 1'd0;
	main_sdram_choose_cmd_cmd_ready <= 1'd0;
	main_sdram_choose_req_want_reads <= 1'd0;
	main_sdram_choose_req_want_writes <= 1'd0;
	main_sdram_en1 <= 1'd0;
	main_sdram_choose_req_cmd_ready <= 1'd0;
	builder_multiplexer_next_state <= builder_multiplexer_state;
	case (builder_multiplexer_state)
		1'd1: begin
			main_sdram_en1 <= 1'd1;
			main_sdram_choose_req_want_writes <= 1'd1;
			if (1'd0) begin
				main_sdram_choose_req_cmd_ready <= (main_sdram_cas_allowed & ((~((main_sdram_choose_req_cmd_payload_ras & (~main_sdram_choose_req_cmd_payload_cas)) & (~main_sdram_choose_req_cmd_payload_we))) | main_sdram_ras_allowed));
			end else begin
				main_sdram_choose_cmd_want_activates <= main_sdram_ras_allowed;
				main_sdram_choose_cmd_cmd_ready <= ((~((main_sdram_choose_cmd_cmd_payload_ras & (~main_sdram_choose_cmd_cmd_payload_cas)) & (~main_sdram_choose_cmd_cmd_payload_we))) | main_sdram_ras_allowed);
				main_sdram_choose_req_cmd_ready <= main_sdram_cas_allowed;
			end
			main_sdram_steerer_sel0 <= 1'd0;
			main_sdram_steerer_sel1 <= 1'd0;
			main_sdram_steerer_sel2 <= 1'd1;
			main_sdram_steerer_sel3 <= 2'd2;
			if (main_sdram_read_available) begin
				if (((~main_sdram_write_available) | main_sdram_max_time1)) begin
					builder_multiplexer_next_state <= 2'd3;
				end
			end
			if (main_sdram_go_to_refresh) begin
				builder_multiplexer_next_state <= 2'd2;
			end
		end
		2'd2: begin
			main_sdram_steerer_sel0 <= 2'd3;
			main_sdram_cmd_ready <= 1'd1;
			if (main_sdram_cmd_last) begin
				builder_multiplexer_next_state <= 1'd0;
			end
		end
		2'd3: begin
			if (main_sdram_twtrcon_ready) begin
				builder_multiplexer_next_state <= 1'd0;
			end
		end
		3'd4: begin
			builder_multiplexer_next_state <= 3'd5;
		end
		3'd5: begin
			builder_multiplexer_next_state <= 3'd6;
		end
		3'd6: begin
			builder_multiplexer_next_state <= 3'd7;
		end
		3'd7: begin
			builder_multiplexer_next_state <= 4'd8;
		end
		4'd8: begin
			builder_multiplexer_next_state <= 4'd9;
		end
		4'd9: begin
			builder_multiplexer_next_state <= 4'd10;
		end
		4'd10: begin
			builder_multiplexer_next_state <= 4'd11;
		end
		4'd11: begin
			builder_multiplexer_next_state <= 1'd1;
		end
		default: begin
			main_sdram_en0 <= 1'd1;
			main_sdram_choose_req_want_reads <= 1'd1;
			if (1'd0) begin
				main_sdram_choose_req_cmd_ready <= (main_sdram_cas_allowed & ((~((main_sdram_choose_req_cmd_payload_ras & (~main_sdram_choose_req_cmd_payload_cas)) & (~main_sdram_choose_req_cmd_payload_we))) | main_sdram_ras_allowed));
			end else begin
				main_sdram_choose_cmd_want_activates <= main_sdram_ras_allowed;
				main_sdram_choose_cmd_cmd_ready <= ((~((main_sdram_choose_cmd_cmd_payload_ras & (~main_sdram_choose_cmd_cmd_payload_cas)) & (~main_sdram_choose_cmd_cmd_payload_we))) | main_sdram_ras_allowed);
				main_sdram_choose_req_cmd_ready <= main_sdram_cas_allowed;
			end
			main_sdram_steerer_sel0 <= 1'd0;
			main_sdram_steerer_sel1 <= 1'd1;
			main_sdram_steerer_sel2 <= 2'd2;
			main_sdram_steerer_sel3 <= 1'd0;
			if (main_sdram_write_available) begin
				if (((~main_sdram_read_available) | main_sdram_max_time0)) begin
					builder_multiplexer_next_state <= 3'd4;
				end
			end
			if (main_sdram_go_to_refresh) begin
				builder_multiplexer_next_state <= 2'd2;
			end
		end
	endcase
end
assign builder_roundrobin0_request = {(((main_port_cmd_payload_addr[9:7] == 1'd0) & (~(((((((builder_locked0 | (main_sdram_interface_bank1_lock & (builder_roundrobin1_grant == 1'd0))) | (main_sdram_interface_bank2_lock & (builder_roundrobin2_grant == 1'd0))) | (main_sdram_interface_bank3_lock & (builder_roundrobin3_grant == 1'd0))) | (main_sdram_interface_bank4_lock & (builder_roundrobin4_grant == 1'd0))) | (main_sdram_interface_bank5_lock & (builder_roundrobin5_grant == 1'd0))) | (main_sdram_interface_bank6_lock & (builder_roundrobin6_grant == 1'd0))) | (main_sdram_interface_bank7_lock & (builder_roundrobin7_grant == 1'd0))))) & main_port_cmd_valid)};
assign builder_roundrobin0_ce = ((~main_sdram_interface_bank0_valid) & (~main_sdram_interface_bank0_lock));
assign main_sdram_interface_bank0_addr = builder_rhs_array_muxed12;
assign main_sdram_interface_bank0_we = builder_rhs_array_muxed13;
assign main_sdram_interface_bank0_valid = builder_rhs_array_muxed14;
assign builder_roundrobin1_request = {(((main_port_cmd_payload_addr[9:7] == 1'd1) & (~(((((((builder_locked1 | (main_sdram_interface_bank0_lock & (builder_roundrobin0_grant == 1'd0))) | (main_sdram_interface_bank2_lock & (builder_roundrobin2_grant == 1'd0))) | (main_sdram_interface_bank3_lock & (builder_roundrobin3_grant == 1'd0))) | (main_sdram_interface_bank4_lock & (builder_roundrobin4_grant == 1'd0))) | (main_sdram_interface_bank5_lock & (builder_roundrobin5_grant == 1'd0))) | (main_sdram_interface_bank6_lock & (builder_roundrobin6_grant == 1'd0))) | (main_sdram_interface_bank7_lock & (builder_roundrobin7_grant == 1'd0))))) & main_port_cmd_valid)};
assign builder_roundrobin1_ce = ((~main_sdram_interface_bank1_valid) & (~main_sdram_interface_bank1_lock));
assign main_sdram_interface_bank1_addr = builder_rhs_array_muxed15;
assign main_sdram_interface_bank1_we = builder_rhs_array_muxed16;
assign main_sdram_interface_bank1_valid = builder_rhs_array_muxed17;
assign builder_roundrobin2_request = {(((main_port_cmd_payload_addr[9:7] == 2'd2) & (~(((((((builder_locked2 | (main_sdram_interface_bank0_lock & (builder_roundrobin0_grant == 1'd0))) | (main_sdram_interface_bank1_lock & (builder_roundrobin1_grant == 1'd0))) | (main_sdram_interface_bank3_lock & (builder_roundrobin3_grant == 1'd0))) | (main_sdram_interface_bank4_lock & (builder_roundrobin4_grant == 1'd0))) | (main_sdram_interface_bank5_lock & (builder_roundrobin5_grant == 1'd0))) | (main_sdram_interface_bank6_lock & (builder_roundrobin6_grant == 1'd0))) | (main_sdram_interface_bank7_lock & (builder_roundrobin7_grant == 1'd0))))) & main_port_cmd_valid)};
assign builder_roundrobin2_ce = ((~main_sdram_interface_bank2_valid) & (~main_sdram_interface_bank2_lock));
assign main_sdram_interface_bank2_addr = builder_rhs_array_muxed18;
assign main_sdram_interface_bank2_we = builder_rhs_array_muxed19;
assign main_sdram_interface_bank2_valid = builder_rhs_array_muxed20;
assign builder_roundrobin3_request = {(((main_port_cmd_payload_addr[9:7] == 2'd3) & (~(((((((builder_locked3 | (main_sdram_interface_bank0_lock & (builder_roundrobin0_grant == 1'd0))) | (main_sdram_interface_bank1_lock & (builder_roundrobin1_grant == 1'd0))) | (main_sdram_interface_bank2_lock & (builder_roundrobin2_grant == 1'd0))) | (main_sdram_interface_bank4_lock & (builder_roundrobin4_grant == 1'd0))) | (main_sdram_interface_bank5_lock & (builder_roundrobin5_grant == 1'd0))) | (main_sdram_interface_bank6_lock & (builder_roundrobin6_grant == 1'd0))) | (main_sdram_interface_bank7_lock & (builder_roundrobin7_grant == 1'd0))))) & main_port_cmd_valid)};
assign builder_roundrobin3_ce = ((~main_sdram_interface_bank3_valid) & (~main_sdram_interface_bank3_lock));
assign main_sdram_interface_bank3_addr = builder_rhs_array_muxed21;
assign main_sdram_interface_bank3_we = builder_rhs_array_muxed22;
assign main_sdram_interface_bank3_valid = builder_rhs_array_muxed23;
assign builder_roundrobin4_request = {(((main_port_cmd_payload_addr[9:7] == 3'd4) & (~(((((((builder_locked4 | (main_sdram_interface_bank0_lock & (builder_roundrobin0_grant == 1'd0))) | (main_sdram_interface_bank1_lock & (builder_roundrobin1_grant == 1'd0))) | (main_sdram_interface_bank2_lock & (builder_roundrobin2_grant == 1'd0))) | (main_sdram_interface_bank3_lock & (builder_roundrobin3_grant == 1'd0))) | (main_sdram_interface_bank5_lock & (builder_roundrobin5_grant == 1'd0))) | (main_sdram_interface_bank6_lock & (builder_roundrobin6_grant == 1'd0))) | (main_sdram_interface_bank7_lock & (builder_roundrobin7_grant == 1'd0))))) & main_port_cmd_valid)};
assign builder_roundrobin4_ce = ((~main_sdram_interface_bank4_valid) & (~main_sdram_interface_bank4_lock));
assign main_sdram_interface_bank4_addr = builder_rhs_array_muxed24;
assign main_sdram_interface_bank4_we = builder_rhs_array_muxed25;
assign main_sdram_interface_bank4_valid = builder_rhs_array_muxed26;
assign builder_roundrobin5_request = {(((main_port_cmd_payload_addr[9:7] == 3'd5) & (~(((((((builder_locked5 | (main_sdram_interface_bank0_lock & (builder_roundrobin0_grant == 1'd0))) | (main_sdram_interface_bank1_lock & (builder_roundrobin1_grant == 1'd0))) | (main_sdram_interface_bank2_lock & (builder_roundrobin2_grant == 1'd0))) | (main_sdram_interface_bank3_lock & (builder_roundrobin3_grant == 1'd0))) | (main_sdram_interface_bank4_lock & (builder_roundrobin4_grant == 1'd0))) | (main_sdram_interface_bank6_lock & (builder_roundrobin6_grant == 1'd0))) | (main_sdram_interface_bank7_lock & (builder_roundrobin7_grant == 1'd0))))) & main_port_cmd_valid)};
assign builder_roundrobin5_ce = ((~main_sdram_interface_bank5_valid) & (~main_sdram_interface_bank5_lock));
assign main_sdram_interface_bank5_addr = builder_rhs_array_muxed27;
assign main_sdram_interface_bank5_we = builder_rhs_array_muxed28;
assign main_sdram_interface_bank5_valid = builder_rhs_array_muxed29;
assign builder_roundrobin6_request = {(((main_port_cmd_payload_addr[9:7] == 3'd6) & (~(((((((builder_locked6 | (main_sdram_interface_bank0_lock & (builder_roundrobin0_grant == 1'd0))) | (main_sdram_interface_bank1_lock & (builder_roundrobin1_grant == 1'd0))) | (main_sdram_interface_bank2_lock & (builder_roundrobin2_grant == 1'd0))) | (main_sdram_interface_bank3_lock & (builder_roundrobin3_grant == 1'd0))) | (main_sdram_interface_bank4_lock & (builder_roundrobin4_grant == 1'd0))) | (main_sdram_interface_bank5_lock & (builder_roundrobin5_grant == 1'd0))) | (main_sdram_interface_bank7_lock & (builder_roundrobin7_grant == 1'd0))))) & main_port_cmd_valid)};
assign builder_roundrobin6_ce = ((~main_sdram_interface_bank6_valid) & (~main_sdram_interface_bank6_lock));
assign main_sdram_interface_bank6_addr = builder_rhs_array_muxed30;
assign main_sdram_interface_bank6_we = builder_rhs_array_muxed31;
assign main_sdram_interface_bank6_valid = builder_rhs_array_muxed32;
assign builder_roundrobin7_request = {(((main_port_cmd_payload_addr[9:7] == 3'd7) & (~(((((((builder_locked7 | (main_sdram_interface_bank0_lock & (builder_roundrobin0_grant == 1'd0))) | (main_sdram_interface_bank1_lock & (builder_roundrobin1_grant == 1'd0))) | (main_sdram_interface_bank2_lock & (builder_roundrobin2_grant == 1'd0))) | (main_sdram_interface_bank3_lock & (builder_roundrobin3_grant == 1'd0))) | (main_sdram_interface_bank4_lock & (builder_roundrobin4_grant == 1'd0))) | (main_sdram_interface_bank5_lock & (builder_roundrobin5_grant == 1'd0))) | (main_sdram_interface_bank6_lock & (builder_roundrobin6_grant == 1'd0))))) & main_port_cmd_valid)};
assign builder_roundrobin7_ce = ((~main_sdram_interface_bank7_valid) & (~main_sdram_interface_bank7_lock));
assign main_sdram_interface_bank7_addr = builder_rhs_array_muxed33;
assign main_sdram_interface_bank7_we = builder_rhs_array_muxed34;
assign main_sdram_interface_bank7_valid = builder_rhs_array_muxed35;
assign main_port_cmd_ready = ((((((((1'd0 | (((builder_roundrobin0_grant == 1'd0) & ((main_port_cmd_payload_addr[9:7] == 1'd0) & (~(((((((builder_locked0 | (main_sdram_interface_bank1_lock & (builder_roundrobin1_grant == 1'd0))) | (main_sdram_interface_bank2_lock & (builder_roundrobin2_grant == 1'd0))) | (main_sdram_interface_bank3_lock & (builder_roundrobin3_grant == 1'd0))) | (main_sdram_interface_bank4_lock & (builder_roundrobin4_grant == 1'd0))) | (main_sdram_interface_bank5_lock & (builder_roundrobin5_grant == 1'd0))) | (main_sdram_interface_bank6_lock & (builder_roundrobin6_grant == 1'd0))) | (main_sdram_interface_bank7_lock & (builder_roundrobin7_grant == 1'd0)))))) & main_sdram_interface_bank0_ready)) | (((builder_roundrobin1_grant == 1'd0) & ((main_port_cmd_payload_addr[9:7] == 1'd1) & (~(((((((builder_locked1 | (main_sdram_interface_bank0_lock & (builder_roundrobin0_grant == 1'd0))) | (main_sdram_interface_bank2_lock & (builder_roundrobin2_grant == 1'd0))) | (main_sdram_interface_bank3_lock & (builder_roundrobin3_grant == 1'd0))) | (main_sdram_interface_bank4_lock & (builder_roundrobin4_grant == 1'd0))) | (main_sdram_interface_bank5_lock & (builder_roundrobin5_grant == 1'd0))) | (main_sdram_interface_bank6_lock & (builder_roundrobin6_grant == 1'd0))) | (main_sdram_interface_bank7_lock & (builder_roundrobin7_grant == 1'd0)))))) & main_sdram_interface_bank1_ready)) | (((builder_roundrobin2_grant == 1'd0) & ((main_port_cmd_payload_addr[9:7] == 2'd2) & (~(((((((builder_locked2 | (main_sdram_interface_bank0_lock & (builder_roundrobin0_grant == 1'd0))) | (main_sdram_interface_bank1_lock & (builder_roundrobin1_grant == 1'd0))) | (main_sdram_interface_bank3_lock & (builder_roundrobin3_grant == 1'd0))) | (main_sdram_interface_bank4_lock & (builder_roundrobin4_grant == 1'd0))) | (main_sdram_interface_bank5_lock & (builder_roundrobin5_grant == 1'd0))) | (main_sdram_interface_bank6_lock & (builder_roundrobin6_grant == 1'd0))) | (main_sdram_interface_bank7_lock & (builder_roundrobin7_grant == 1'd0)))))) & main_sdram_interface_bank2_ready)) | (((builder_roundrobin3_grant == 1'd0) & ((main_port_cmd_payload_addr[9:7] == 2'd3) & (~(((((((builder_locked3 | (main_sdram_interface_bank0_lock & (builder_roundrobin0_grant == 1'd0))) | (main_sdram_interface_bank1_lock & (builder_roundrobin1_grant == 1'd0))) | (main_sdram_interface_bank2_lock & (builder_roundrobin2_grant == 1'd0))) | (main_sdram_interface_bank4_lock & (builder_roundrobin4_grant == 1'd0))) | (main_sdram_interface_bank5_lock & (builder_roundrobin5_grant == 1'd0))) | (main_sdram_interface_bank6_lock & (builder_roundrobin6_grant == 1'd0))) | (main_sdram_interface_bank7_lock & (builder_roundrobin7_grant == 1'd0)))))) & main_sdram_interface_bank3_ready)) | (((builder_roundrobin4_grant == 1'd0) & ((main_port_cmd_payload_addr[9:7] == 3'd4) & (~(((((((builder_locked4 | (main_sdram_interface_bank0_lock & (builder_roundrobin0_grant == 1'd0))) | (main_sdram_interface_bank1_lock & (builder_roundrobin1_grant == 1'd0))) | (main_sdram_interface_bank2_lock & (builder_roundrobin2_grant == 1'd0))) | (main_sdram_interface_bank3_lock & (builder_roundrobin3_grant == 1'd0))) | (main_sdram_interface_bank5_lock & (builder_roundrobin5_grant == 1'd0))) | (main_sdram_interface_bank6_lock & (builder_roundrobin6_grant == 1'd0))) | (main_sdram_interface_bank7_lock & (builder_roundrobin7_grant == 1'd0)))))) & main_sdram_interface_bank4_ready)) | (((builder_roundrobin5_grant == 1'd0) & ((main_port_cmd_payload_addr[9:7] == 3'd5) & (~(((((((builder_locked5 | (main_sdram_interface_bank0_lock & (builder_roundrobin0_grant == 1'd0))) | (main_sdram_interface_bank1_lock & (builder_roundrobin1_grant == 1'd0))) | (main_sdram_interface_bank2_lock & (builder_roundrobin2_grant == 1'd0))) | (main_sdram_interface_bank3_lock & (builder_roundrobin3_grant == 1'd0))) | (main_sdram_interface_bank4_lock & (builder_roundrobin4_grant == 1'd0))) | (main_sdram_interface_bank6_lock & (builder_roundrobin6_grant == 1'd0))) | (main_sdram_interface_bank7_lock & (builder_roundrobin7_grant == 1'd0)))))) & main_sdram_interface_bank5_ready)) | (((builder_roundrobin6_grant == 1'd0) & ((main_port_cmd_payload_addr[9:7] == 3'd6) & (~(((((((builder_locked6 | (main_sdram_interface_bank0_lock & (builder_roundrobin0_grant == 1'd0))) | (main_sdram_interface_bank1_lock & (builder_roundrobin1_grant == 1'd0))) | (main_sdram_interface_bank2_lock & (builder_roundrobin2_grant == 1'd0))) | (main_sdram_interface_bank3_lock & (builder_roundrobin3_grant == 1'd0))) | (main_sdram_interface_bank4_lock & (builder_roundrobin4_grant == 1'd0))) | (main_sdram_interface_bank5_lock & (builder_roundrobin5_grant == 1'd0))) | (main_sdram_interface_bank7_lock & (builder_roundrobin7_grant == 1'd0)))))) & main_sdram_interface_bank6_ready)) | (((builder_roundrobin7_grant == 1'd0) & ((main_port_cmd_payload_addr[9:7] == 3'd7) & (~(((((((builder_locked7 | (main_sdram_interface_bank0_lock & (builder_roundrobin0_grant == 1'd0))) | (main_sdram_interface_bank1_lock & (builder_roundrobin1_grant == 1'd0))) | (main_sdram_interface_bank2_lock & (builder_roundrobin2_grant == 1'd0))) | (main_sdram_interface_bank3_lock & (builder_roundrobin3_grant == 1'd0))) | (main_sdram_interface_bank4_lock & (builder_roundrobin4_grant == 1'd0))) | (main_sdram_interface_bank5_lock & (builder_roundrobin5_grant == 1'd0))) | (main_sdram_interface_bank6_lock & (builder_roundrobin6_grant == 1'd0)))))) & main_sdram_interface_bank7_ready));
assign main_port_wdata_ready = builder_new_master_wdata_ready2;
assign main_port_rdata_valid = builder_new_master_rdata_valid9;
always @(*) begin
	main_sdram_interface_wdata <= 128'd0;
	main_sdram_interface_wdata_we <= 16'd0;
	case ({builder_new_master_wdata_ready2})
		1'd1: begin
			main_sdram_interface_wdata <= main_port_wdata_payload_data;
			main_sdram_interface_wdata_we <= main_port_wdata_payload_we;
		end
		default: begin
			main_sdram_interface_wdata <= 1'd0;
			main_sdram_interface_wdata_we <= 1'd0;
		end
	endcase
end
assign main_port_rdata_payload_data = main_sdram_interface_rdata;
assign builder_roundrobin0_grant = 1'd0;
assign builder_roundrobin1_grant = 1'd0;
assign builder_roundrobin2_grant = 1'd0;
assign builder_roundrobin3_grant = 1'd0;
assign builder_roundrobin4_grant = 1'd0;
assign builder_roundrobin5_grant = 1'd0;
assign builder_roundrobin6_grant = 1'd0;
assign builder_roundrobin7_grant = 1'd0;
assign main_data_port_adr = main_interface0_wb_sdram_adr[2];
always @(*) begin
	main_data_port_dat_w <= 128'd0;
	main_data_port_we <= 16'd0;
	if (main_write_from_slave) begin
		main_data_port_dat_w <= main_dat_r;
		main_data_port_we <= {16{1'd1}};
	end else begin
		main_data_port_dat_w <= {4{main_interface0_wb_sdram_dat_w}};
		if ((((main_interface0_wb_sdram_cyc & main_interface0_wb_sdram_stb) & main_interface0_wb_sdram_we) & main_interface0_wb_sdram_ack)) begin
			main_data_port_we <= {({4{(main_interface0_wb_sdram_adr[1:0] == 1'd0)}} & main_interface0_wb_sdram_sel), ({4{(main_interface0_wb_sdram_adr[1:0] == 1'd1)}} & main_interface0_wb_sdram_sel), ({4{(main_interface0_wb_sdram_adr[1:0] == 2'd2)}} & main_interface0_wb_sdram_sel), ({4{(main_interface0_wb_sdram_adr[1:0] == 2'd3)}} & main_interface0_wb_sdram_sel)};
		end
	end
end
assign main_dat_w = main_data_port_dat_r;
assign main_sel = 16'd65535;
always @(*) begin
	main_interface0_wb_sdram_dat_r <= 32'd0;
	case (main_adr_offset_r)
		1'd0: begin
			main_interface0_wb_sdram_dat_r <= main_data_port_dat_r[127:96];
		end
		1'd1: begin
			main_interface0_wb_sdram_dat_r <= main_data_port_dat_r[95:64];
		end
		2'd2: begin
			main_interface0_wb_sdram_dat_r <= main_data_port_dat_r[63:32];
		end
		default: begin
			main_interface0_wb_sdram_dat_r <= main_data_port_dat_r[31:0];
		end
	endcase
end
assign {main_tag_do_dirty, main_tag_do_tag} = main_tag_port_dat_r;
assign main_tag_port_dat_w = {main_tag_di_dirty, main_tag_di_tag};
assign main_tag_port_adr = main_interface0_wb_sdram_adr[2];
assign main_tag_di_tag = main_interface0_wb_sdram_adr[29:3];
assign main_adr = {main_tag_do_tag, main_interface0_wb_sdram_adr[2]};
always @(*) begin
	main_word_inc <= 1'd0;
	main_write_from_slave <= 1'd0;
	main_interface0_wb_sdram_ack <= 1'd0;
	main_cyc <= 1'd0;
	main_stb <= 1'd0;
	main_tag_port_we <= 1'd0;
	main_we <= 1'd0;
	builder_fullmemorywe_next_state <= 2'd0;
	main_tag_di_dirty <= 1'd0;
	main_word_clr <= 1'd0;
	builder_fullmemorywe_next_state <= builder_fullmemorywe_state;
	case (builder_fullmemorywe_state)
		1'd1: begin
			main_word_clr <= 1'd1;
			if ((main_tag_do_tag == main_interface0_wb_sdram_adr[29:3])) begin
				main_interface0_wb_sdram_ack <= 1'd1;
				if (main_interface0_wb_sdram_we) begin
					main_tag_di_dirty <= 1'd1;
					main_tag_port_we <= 1'd1;
				end
				builder_fullmemorywe_next_state <= 1'd0;
			end else begin
				if (main_tag_do_dirty) begin
					builder_fullmemorywe_next_state <= 2'd2;
				end else begin
					main_tag_port_we <= 1'd1;
					main_word_clr <= 1'd1;
					builder_fullmemorywe_next_state <= 2'd3;
				end
			end
		end
		2'd2: begin
			main_stb <= 1'd1;
			main_cyc <= 1'd1;
			main_we <= 1'd1;
			if (main_ack) begin
				main_word_inc <= 1'd1;
				if (1'd1) begin
					main_tag_port_we <= 1'd1;
					main_word_clr <= 1'd1;
					builder_fullmemorywe_next_state <= 2'd3;
				end
			end
		end
		2'd3: begin
			main_stb <= 1'd1;
			main_cyc <= 1'd1;
			main_we <= 1'd0;
			if (main_ack) begin
				main_write_from_slave <= 1'd1;
				main_word_inc <= 1'd1;
				if (1'd1) begin
					builder_fullmemorywe_next_state <= 1'd1;
				end else begin
					builder_fullmemorywe_next_state <= 2'd3;
				end
			end
		end
		default: begin
			if ((main_interface0_wb_sdram_cyc & main_interface0_wb_sdram_stb)) begin
				builder_fullmemorywe_next_state <= 1'd1;
			end
		end
	endcase
end
assign main_wdata_converter_sink_valid = ((main_cyc & main_stb) & main_we);
assign main_wdata_converter_sink_payload_data = main_dat_w;
assign main_wdata_converter_sink_payload_we = main_sel;
assign main_port_wdata_valid = main_wdata_converter_source_valid;
assign main_wdata_converter_source_ready = main_port_wdata_ready;
assign main_port_wdata_first = main_wdata_converter_source_first;
assign main_port_wdata_last = main_wdata_converter_source_last;
assign main_port_wdata_payload_data = main_wdata_converter_source_payload_data;
assign main_port_wdata_payload_we = main_wdata_converter_source_payload_we;
assign main_rdata_converter_sink_valid = main_port_rdata_valid;
assign main_port_rdata_ready = main_rdata_converter_sink_ready;
assign main_rdata_converter_sink_first = main_port_rdata_first;
assign main_rdata_converter_sink_last = main_port_rdata_last;
assign main_rdata_converter_sink_payload_data = main_port_rdata_payload_data;
assign main_rdata_converter_source_ready = 1'd1;
assign main_dat_r = main_rdata_converter_source_payload_data;
assign main_wdata_converter_converter_sink_valid = main_wdata_converter_sink_valid;
assign main_wdata_converter_converter_sink_first = main_wdata_converter_sink_first;
assign main_wdata_converter_converter_sink_last = main_wdata_converter_sink_last;
assign main_wdata_converter_sink_ready = main_wdata_converter_converter_sink_ready;
assign main_wdata_converter_converter_sink_payload_data = {main_wdata_converter_sink_payload_we, main_wdata_converter_sink_payload_data};
assign main_wdata_converter_source_valid = main_wdata_converter_source_source_valid;
assign main_wdata_converter_source_first = main_wdata_converter_source_source_first;
assign main_wdata_converter_source_last = main_wdata_converter_source_source_last;
assign main_wdata_converter_source_source_ready = main_wdata_converter_source_ready;
assign {main_wdata_converter_source_payload_we, main_wdata_converter_source_payload_data} = main_wdata_converter_source_source_payload_data;
assign main_wdata_converter_source_source_valid = main_wdata_converter_converter_source_valid;
assign main_wdata_converter_converter_source_ready = main_wdata_converter_source_source_ready;
assign main_wdata_converter_source_source_first = main_wdata_converter_converter_source_first;
assign main_wdata_converter_source_source_last = main_wdata_converter_converter_source_last;
assign main_wdata_converter_source_source_payload_data = main_wdata_converter_converter_source_payload_data;
assign main_wdata_converter_converter_source_valid = main_wdata_converter_converter_sink_valid;
assign main_wdata_converter_converter_sink_ready = main_wdata_converter_converter_source_ready;
assign main_wdata_converter_converter_source_first = main_wdata_converter_converter_sink_first;
assign main_wdata_converter_converter_source_last = main_wdata_converter_converter_sink_last;
assign main_wdata_converter_converter_source_payload_data = main_wdata_converter_converter_sink_payload_data;
assign main_wdata_converter_converter_source_payload_valid_token_count = 1'd1;
assign main_rdata_converter_converter_sink_valid = main_rdata_converter_sink_valid;
assign main_rdata_converter_converter_sink_first = main_rdata_converter_sink_first;
assign main_rdata_converter_converter_sink_last = main_rdata_converter_sink_last;
assign main_rdata_converter_sink_ready = main_rdata_converter_converter_sink_ready;
assign main_rdata_converter_converter_sink_payload_data = {main_rdata_converter_sink_payload_data};
assign main_rdata_converter_source_valid = main_rdata_converter_source_source_valid;
assign main_rdata_converter_source_first = main_rdata_converter_source_source_first;
assign main_rdata_converter_source_last = main_rdata_converter_source_source_last;
assign main_rdata_converter_source_source_ready = main_rdata_converter_source_ready;
assign {main_rdata_converter_source_payload_data} = main_rdata_converter_source_source_payload_data;
assign main_rdata_converter_source_source_valid = main_rdata_converter_converter_source_valid;
assign main_rdata_converter_converter_source_ready = main_rdata_converter_source_source_ready;
assign main_rdata_converter_source_source_first = main_rdata_converter_converter_source_first;
assign main_rdata_converter_source_source_last = main_rdata_converter_converter_source_last;
assign main_rdata_converter_source_source_payload_data = main_rdata_converter_converter_source_payload_data;
assign main_rdata_converter_converter_source_valid = main_rdata_converter_converter_sink_valid;
assign main_rdata_converter_converter_sink_ready = main_rdata_converter_converter_source_ready;
assign main_rdata_converter_converter_source_first = main_rdata_converter_converter_sink_first;
assign main_rdata_converter_converter_source_last = main_rdata_converter_converter_sink_last;
assign main_rdata_converter_converter_source_payload_data = main_rdata_converter_converter_sink_payload_data;
assign main_rdata_converter_converter_source_payload_valid_token_count = 1'd1;
always @(*) begin
	main_port_cmd_payload_addr <= 24'd0;
	main_count_next_value <= 1'd0;
	main_count_next_value_ce <= 1'd0;
	main_port_cmd_valid <= 1'd0;
	builder_litedramwishbone2native_next_state <= 2'd0;
	main_ack <= 1'd0;
	main_port_cmd_payload_we <= 1'd0;
	builder_litedramwishbone2native_next_state <= builder_litedramwishbone2native_state;
	case (builder_litedramwishbone2native_state)
		1'd1: begin
			if (main_wdata_converter_sink_ready) begin
				main_ack <= 1'd1;
				builder_litedramwishbone2native_next_state <= 1'd0;
			end
		end
		2'd2: begin
			if (main_rdata_converter_source_valid) begin
				main_ack <= 1'd1;
				builder_litedramwishbone2native_next_state <= 1'd0;
			end
		end
		default: begin
			main_port_cmd_valid <= (main_cyc & main_stb);
			main_port_cmd_payload_we <= main_we;
			main_port_cmd_payload_addr <= (((main_adr * 1'd1) + main_count) - 1'd0);
			if ((main_port_cmd_valid & main_port_cmd_ready)) begin
				main_count_next_value <= (main_count + 1'd1);
				main_count_next_value_ce <= 1'd1;
				if ((main_count == 1'd0)) begin
					main_count_next_value <= 1'd0;
					main_count_next_value_ce <= 1'd1;
					if (main_we) begin
						builder_litedramwishbone2native_next_state <= 1'd1;
					end else begin
						builder_litedramwishbone2native_next_state <= 2'd2;
					end
				end
			end
		end
	endcase
end
assign main_interface0_wb_sdram_adr = builder_rhs_array_muxed36;
assign main_interface0_wb_sdram_dat_w = builder_rhs_array_muxed37;
assign main_interface0_wb_sdram_sel = builder_rhs_array_muxed38;
assign main_interface0_wb_sdram_cyc = builder_rhs_array_muxed39;
assign main_interface0_wb_sdram_stb = builder_rhs_array_muxed40;
assign main_interface0_wb_sdram_we = builder_rhs_array_muxed41;
assign main_interface0_wb_sdram_cti = builder_rhs_array_muxed42;
assign main_interface0_wb_sdram_bte = builder_rhs_array_muxed43;
assign main_interface1_wb_sdram_dat_r = main_interface0_wb_sdram_dat_r;
assign main_interface1_wb_sdram_ack = (main_interface0_wb_sdram_ack & (builder_wb_sdram_con_grant == 1'd0));
assign main_interface1_wb_sdram_err = (main_interface0_wb_sdram_err & (builder_wb_sdram_con_grant == 1'd0));
assign builder_wb_sdram_con_request = {main_interface1_wb_sdram_cyc};
assign builder_wb_sdram_con_grant = 1'd0;
assign builder_basesoc_shared_adr = builder_rhs_array_muxed44;
assign builder_basesoc_shared_dat_w = builder_rhs_array_muxed45;
assign builder_basesoc_shared_sel = builder_rhs_array_muxed46;
assign builder_basesoc_shared_cyc = builder_rhs_array_muxed47;
assign builder_basesoc_shared_stb = builder_rhs_array_muxed48;
assign builder_basesoc_shared_we = builder_rhs_array_muxed49;
assign builder_basesoc_shared_cti = builder_rhs_array_muxed50;
assign builder_basesoc_shared_bte = builder_rhs_array_muxed51;
assign main_uart_wishbone_dat_r = builder_basesoc_shared_dat_r;
assign main_uart_wishbone_ack = (builder_basesoc_shared_ack & (builder_basesoc_grant == 1'd0));
assign main_uart_wishbone_err = (builder_basesoc_shared_err & (builder_basesoc_grant == 1'd0));
assign builder_basesoc_request = {main_uart_wishbone_cyc};
assign builder_basesoc_grant = 1'd0;
always @(*) begin
	builder_basesoc_slave_sel <= 3'd0;
	builder_basesoc_slave_sel[0] <= (builder_basesoc_shared_adr[28:10] == 13'd4096);
	builder_basesoc_slave_sel[1] <= (builder_basesoc_shared_adr[28:14] == 10'd512);
	builder_basesoc_slave_sel[2] <= (builder_basesoc_shared_adr[28:26] == 3'd4);
end
assign main_sram_bus_adr = builder_basesoc_shared_adr;
assign main_sram_bus_dat_w = builder_basesoc_shared_dat_w;
assign main_sram_bus_sel = builder_basesoc_shared_sel;
assign main_sram_bus_stb = builder_basesoc_shared_stb;
assign main_sram_bus_we = builder_basesoc_shared_we;
assign main_sram_bus_cti = builder_basesoc_shared_cti;
assign main_sram_bus_bte = builder_basesoc_shared_bte;
assign main_bus_wishbone_adr = builder_basesoc_shared_adr;
assign main_bus_wishbone_dat_w = builder_basesoc_shared_dat_w;
assign main_bus_wishbone_sel = builder_basesoc_shared_sel;
assign main_bus_wishbone_stb = builder_basesoc_shared_stb;
assign main_bus_wishbone_we = builder_basesoc_shared_we;
assign main_bus_wishbone_cti = builder_basesoc_shared_cti;
assign main_bus_wishbone_bte = builder_basesoc_shared_bte;
assign main_interface1_wb_sdram_adr = builder_basesoc_shared_adr;
assign main_interface1_wb_sdram_dat_w = builder_basesoc_shared_dat_w;
assign main_interface1_wb_sdram_sel = builder_basesoc_shared_sel;
assign main_interface1_wb_sdram_stb = builder_basesoc_shared_stb;
assign main_interface1_wb_sdram_we = builder_basesoc_shared_we;
assign main_interface1_wb_sdram_cti = builder_basesoc_shared_cti;
assign main_interface1_wb_sdram_bte = builder_basesoc_shared_bte;
assign main_sram_bus_cyc = (builder_basesoc_shared_cyc & builder_basesoc_slave_sel[0]);
assign main_bus_wishbone_cyc = (builder_basesoc_shared_cyc & builder_basesoc_slave_sel[1]);
assign main_interface1_wb_sdram_cyc = (builder_basesoc_shared_cyc & builder_basesoc_slave_sel[2]);
assign builder_basesoc_shared_err = ((main_sram_bus_err | main_bus_wishbone_err) | main_interface1_wb_sdram_err);
assign builder_basesoc_wait = ((builder_basesoc_shared_stb & builder_basesoc_shared_cyc) & (~builder_basesoc_shared_ack));
always @(*) begin
	builder_basesoc_shared_ack <= 1'd0;
	builder_basesoc_shared_dat_r <= 32'd0;
	builder_basesoc_error <= 1'd0;
	builder_basesoc_shared_ack <= ((main_sram_bus_ack | main_bus_wishbone_ack) | main_interface1_wb_sdram_ack);
	builder_basesoc_shared_dat_r <= ((({32{builder_basesoc_slave_sel_r[0]}} & main_sram_bus_dat_r) | ({32{builder_basesoc_slave_sel_r[1]}} & main_bus_wishbone_dat_r)) | ({32{builder_basesoc_slave_sel_r[2]}} & main_interface1_wb_sdram_dat_r));
	if (builder_basesoc_done) begin
		builder_basesoc_shared_dat_r <= 32'd4294967295;
		builder_basesoc_shared_ack <= 1'd1;
		builder_basesoc_error <= 1'd1;
	end
end
assign builder_basesoc_done = (builder_basesoc_count == 1'd0);
assign builder_basesoc_csrbankarray_csrbank0_sel = (builder_basesoc_csrbankarray_interface0_bank_bus_adr[13:9] == 1'd0);
assign builder_basesoc_csrbankarray_csrbank0_reset0_r = builder_basesoc_csrbankarray_interface0_bank_bus_dat_w[0];
assign builder_basesoc_csrbankarray_csrbank0_reset0_re = ((builder_basesoc_csrbankarray_csrbank0_sel & builder_basesoc_csrbankarray_interface0_bank_bus_we) & (builder_basesoc_csrbankarray_interface0_bank_bus_adr[3:0] == 1'd0));
assign builder_basesoc_csrbankarray_csrbank0_reset0_we = ((builder_basesoc_csrbankarray_csrbank0_sel & (~builder_basesoc_csrbankarray_interface0_bank_bus_we)) & (builder_basesoc_csrbankarray_interface0_bank_bus_adr[3:0] == 1'd0));
assign builder_basesoc_csrbankarray_csrbank0_scratch3_r = builder_basesoc_csrbankarray_interface0_bank_bus_dat_w[7:0];
assign builder_basesoc_csrbankarray_csrbank0_scratch3_re = ((builder_basesoc_csrbankarray_csrbank0_sel & builder_basesoc_csrbankarray_interface0_bank_bus_we) & (builder_basesoc_csrbankarray_interface0_bank_bus_adr[3:0] == 1'd1));
assign builder_basesoc_csrbankarray_csrbank0_scratch3_we = ((builder_basesoc_csrbankarray_csrbank0_sel & (~builder_basesoc_csrbankarray_interface0_bank_bus_we)) & (builder_basesoc_csrbankarray_interface0_bank_bus_adr[3:0] == 1'd1));
assign builder_basesoc_csrbankarray_csrbank0_scratch2_r = builder_basesoc_csrbankarray_interface0_bank_bus_dat_w[7:0];
assign builder_basesoc_csrbankarray_csrbank0_scratch2_re = ((builder_basesoc_csrbankarray_csrbank0_sel & builder_basesoc_csrbankarray_interface0_bank_bus_we) & (builder_basesoc_csrbankarray_interface0_bank_bus_adr[3:0] == 2'd2));
assign builder_basesoc_csrbankarray_csrbank0_scratch2_we = ((builder_basesoc_csrbankarray_csrbank0_sel & (~builder_basesoc_csrbankarray_interface0_bank_bus_we)) & (builder_basesoc_csrbankarray_interface0_bank_bus_adr[3:0] == 2'd2));
assign builder_basesoc_csrbankarray_csrbank0_scratch1_r = builder_basesoc_csrbankarray_interface0_bank_bus_dat_w[7:0];
assign builder_basesoc_csrbankarray_csrbank0_scratch1_re = ((builder_basesoc_csrbankarray_csrbank0_sel & builder_basesoc_csrbankarray_interface0_bank_bus_we) & (builder_basesoc_csrbankarray_interface0_bank_bus_adr[3:0] == 2'd3));
assign builder_basesoc_csrbankarray_csrbank0_scratch1_we = ((builder_basesoc_csrbankarray_csrbank0_sel & (~builder_basesoc_csrbankarray_interface0_bank_bus_we)) & (builder_basesoc_csrbankarray_interface0_bank_bus_adr[3:0] == 2'd3));
assign builder_basesoc_csrbankarray_csrbank0_scratch0_r = builder_basesoc_csrbankarray_interface0_bank_bus_dat_w[7:0];
assign builder_basesoc_csrbankarray_csrbank0_scratch0_re = ((builder_basesoc_csrbankarray_csrbank0_sel & builder_basesoc_csrbankarray_interface0_bank_bus_we) & (builder_basesoc_csrbankarray_interface0_bank_bus_adr[3:0] == 3'd4));
assign builder_basesoc_csrbankarray_csrbank0_scratch0_we = ((builder_basesoc_csrbankarray_csrbank0_sel & (~builder_basesoc_csrbankarray_interface0_bank_bus_we)) & (builder_basesoc_csrbankarray_interface0_bank_bus_adr[3:0] == 3'd4));
assign builder_basesoc_csrbankarray_csrbank0_bus_errors3_r = builder_basesoc_csrbankarray_interface0_bank_bus_dat_w[7:0];
assign builder_basesoc_csrbankarray_csrbank0_bus_errors3_re = ((builder_basesoc_csrbankarray_csrbank0_sel & builder_basesoc_csrbankarray_interface0_bank_bus_we) & (builder_basesoc_csrbankarray_interface0_bank_bus_adr[3:0] == 3'd5));
assign builder_basesoc_csrbankarray_csrbank0_bus_errors3_we = ((builder_basesoc_csrbankarray_csrbank0_sel & (~builder_basesoc_csrbankarray_interface0_bank_bus_we)) & (builder_basesoc_csrbankarray_interface0_bank_bus_adr[3:0] == 3'd5));
assign builder_basesoc_csrbankarray_csrbank0_bus_errors2_r = builder_basesoc_csrbankarray_interface0_bank_bus_dat_w[7:0];
assign builder_basesoc_csrbankarray_csrbank0_bus_errors2_re = ((builder_basesoc_csrbankarray_csrbank0_sel & builder_basesoc_csrbankarray_interface0_bank_bus_we) & (builder_basesoc_csrbankarray_interface0_bank_bus_adr[3:0] == 3'd6));
assign builder_basesoc_csrbankarray_csrbank0_bus_errors2_we = ((builder_basesoc_csrbankarray_csrbank0_sel & (~builder_basesoc_csrbankarray_interface0_bank_bus_we)) & (builder_basesoc_csrbankarray_interface0_bank_bus_adr[3:0] == 3'd6));
assign builder_basesoc_csrbankarray_csrbank0_bus_errors1_r = builder_basesoc_csrbankarray_interface0_bank_bus_dat_w[7:0];
assign builder_basesoc_csrbankarray_csrbank0_bus_errors1_re = ((builder_basesoc_csrbankarray_csrbank0_sel & builder_basesoc_csrbankarray_interface0_bank_bus_we) & (builder_basesoc_csrbankarray_interface0_bank_bus_adr[3:0] == 3'd7));
assign builder_basesoc_csrbankarray_csrbank0_bus_errors1_we = ((builder_basesoc_csrbankarray_csrbank0_sel & (~builder_basesoc_csrbankarray_interface0_bank_bus_we)) & (builder_basesoc_csrbankarray_interface0_bank_bus_adr[3:0] == 3'd7));
assign builder_basesoc_csrbankarray_csrbank0_bus_errors0_r = builder_basesoc_csrbankarray_interface0_bank_bus_dat_w[7:0];
assign builder_basesoc_csrbankarray_csrbank0_bus_errors0_re = ((builder_basesoc_csrbankarray_csrbank0_sel & builder_basesoc_csrbankarray_interface0_bank_bus_we) & (builder_basesoc_csrbankarray_interface0_bank_bus_adr[3:0] == 4'd8));
assign builder_basesoc_csrbankarray_csrbank0_bus_errors0_we = ((builder_basesoc_csrbankarray_csrbank0_sel & (~builder_basesoc_csrbankarray_interface0_bank_bus_we)) & (builder_basesoc_csrbankarray_interface0_bank_bus_adr[3:0] == 4'd8));
assign builder_basesoc_csrbankarray_csrbank0_reset0_w = main_ctrl_reset_storage;
assign builder_basesoc_csrbankarray_csrbank0_scratch3_w = main_ctrl_scratch_storage[31:24];
assign builder_basesoc_csrbankarray_csrbank0_scratch2_w = main_ctrl_scratch_storage[23:16];
assign builder_basesoc_csrbankarray_csrbank0_scratch1_w = main_ctrl_scratch_storage[15:8];
assign builder_basesoc_csrbankarray_csrbank0_scratch0_w = main_ctrl_scratch_storage[7:0];
assign builder_basesoc_csrbankarray_csrbank0_bus_errors3_w = main_ctrl_bus_errors_status[31:24];
assign builder_basesoc_csrbankarray_csrbank0_bus_errors2_w = main_ctrl_bus_errors_status[23:16];
assign builder_basesoc_csrbankarray_csrbank0_bus_errors1_w = main_ctrl_bus_errors_status[15:8];
assign builder_basesoc_csrbankarray_csrbank0_bus_errors0_w = main_ctrl_bus_errors_status[7:0];
assign main_ctrl_bus_errors_we = builder_basesoc_csrbankarray_csrbank0_bus_errors0_we;
assign builder_basesoc_csrbankarray_csrbank1_sel = (builder_basesoc_csrbankarray_interface1_bank_bus_adr[13:9] == 3'd5);
assign builder_basesoc_csrbankarray_csrbank1_half_sys8x_taps0_r = builder_basesoc_csrbankarray_interface1_bank_bus_dat_w[4:0];
assign builder_basesoc_csrbankarray_csrbank1_half_sys8x_taps0_re = ((builder_basesoc_csrbankarray_csrbank1_sel & builder_basesoc_csrbankarray_interface1_bank_bus_we) & (builder_basesoc_csrbankarray_interface1_bank_bus_adr[2:0] == 1'd0));
assign builder_basesoc_csrbankarray_csrbank1_half_sys8x_taps0_we = ((builder_basesoc_csrbankarray_csrbank1_sel & (~builder_basesoc_csrbankarray_interface1_bank_bus_we)) & (builder_basesoc_csrbankarray_interface1_bank_bus_adr[2:0] == 1'd0));
assign main_a7ddrphy_cdly_rst_r = builder_basesoc_csrbankarray_interface1_bank_bus_dat_w[0];
assign main_a7ddrphy_cdly_rst_re = ((builder_basesoc_csrbankarray_csrbank1_sel & builder_basesoc_csrbankarray_interface1_bank_bus_we) & (builder_basesoc_csrbankarray_interface1_bank_bus_adr[2:0] == 1'd1));
assign main_a7ddrphy_cdly_rst_we = ((builder_basesoc_csrbankarray_csrbank1_sel & (~builder_basesoc_csrbankarray_interface1_bank_bus_we)) & (builder_basesoc_csrbankarray_interface1_bank_bus_adr[2:0] == 1'd1));
assign main_a7ddrphy_cdly_inc_r = builder_basesoc_csrbankarray_interface1_bank_bus_dat_w[0];
assign main_a7ddrphy_cdly_inc_re = ((builder_basesoc_csrbankarray_csrbank1_sel & builder_basesoc_csrbankarray_interface1_bank_bus_we) & (builder_basesoc_csrbankarray_interface1_bank_bus_adr[2:0] == 2'd2));
assign main_a7ddrphy_cdly_inc_we = ((builder_basesoc_csrbankarray_csrbank1_sel & (~builder_basesoc_csrbankarray_interface1_bank_bus_we)) & (builder_basesoc_csrbankarray_interface1_bank_bus_adr[2:0] == 2'd2));
assign builder_basesoc_csrbankarray_csrbank1_dly_sel0_r = builder_basesoc_csrbankarray_interface1_bank_bus_dat_w[1:0];
assign builder_basesoc_csrbankarray_csrbank1_dly_sel0_re = ((builder_basesoc_csrbankarray_csrbank1_sel & builder_basesoc_csrbankarray_interface1_bank_bus_we) & (builder_basesoc_csrbankarray_interface1_bank_bus_adr[2:0] == 2'd3));
assign builder_basesoc_csrbankarray_csrbank1_dly_sel0_we = ((builder_basesoc_csrbankarray_csrbank1_sel & (~builder_basesoc_csrbankarray_interface1_bank_bus_we)) & (builder_basesoc_csrbankarray_interface1_bank_bus_adr[2:0] == 2'd3));
assign main_a7ddrphy_rdly_dq_rst_r = builder_basesoc_csrbankarray_interface1_bank_bus_dat_w[0];
assign main_a7ddrphy_rdly_dq_rst_re = ((builder_basesoc_csrbankarray_csrbank1_sel & builder_basesoc_csrbankarray_interface1_bank_bus_we) & (builder_basesoc_csrbankarray_interface1_bank_bus_adr[2:0] == 3'd4));
assign main_a7ddrphy_rdly_dq_rst_we = ((builder_basesoc_csrbankarray_csrbank1_sel & (~builder_basesoc_csrbankarray_interface1_bank_bus_we)) & (builder_basesoc_csrbankarray_interface1_bank_bus_adr[2:0] == 3'd4));
assign main_a7ddrphy_rdly_dq_inc_r = builder_basesoc_csrbankarray_interface1_bank_bus_dat_w[0];
assign main_a7ddrphy_rdly_dq_inc_re = ((builder_basesoc_csrbankarray_csrbank1_sel & builder_basesoc_csrbankarray_interface1_bank_bus_we) & (builder_basesoc_csrbankarray_interface1_bank_bus_adr[2:0] == 3'd5));
assign main_a7ddrphy_rdly_dq_inc_we = ((builder_basesoc_csrbankarray_csrbank1_sel & (~builder_basesoc_csrbankarray_interface1_bank_bus_we)) & (builder_basesoc_csrbankarray_interface1_bank_bus_adr[2:0] == 3'd5));
assign main_a7ddrphy_rdly_dq_bitslip_rst_r = builder_basesoc_csrbankarray_interface1_bank_bus_dat_w[0];
assign main_a7ddrphy_rdly_dq_bitslip_rst_re = ((builder_basesoc_csrbankarray_csrbank1_sel & builder_basesoc_csrbankarray_interface1_bank_bus_we) & (builder_basesoc_csrbankarray_interface1_bank_bus_adr[2:0] == 3'd6));
assign main_a7ddrphy_rdly_dq_bitslip_rst_we = ((builder_basesoc_csrbankarray_csrbank1_sel & (~builder_basesoc_csrbankarray_interface1_bank_bus_we)) & (builder_basesoc_csrbankarray_interface1_bank_bus_adr[2:0] == 3'd6));
assign main_a7ddrphy_rdly_dq_bitslip_r = builder_basesoc_csrbankarray_interface1_bank_bus_dat_w[0];
assign main_a7ddrphy_rdly_dq_bitslip_re = ((builder_basesoc_csrbankarray_csrbank1_sel & builder_basesoc_csrbankarray_interface1_bank_bus_we) & (builder_basesoc_csrbankarray_interface1_bank_bus_adr[2:0] == 3'd7));
assign main_a7ddrphy_rdly_dq_bitslip_we = ((builder_basesoc_csrbankarray_csrbank1_sel & (~builder_basesoc_csrbankarray_interface1_bank_bus_we)) & (builder_basesoc_csrbankarray_interface1_bank_bus_adr[2:0] == 3'd7));
assign builder_basesoc_csrbankarray_csrbank1_half_sys8x_taps0_w = main_a7ddrphy_half_sys8x_taps_storage[4:0];
assign builder_basesoc_csrbankarray_csrbank1_dly_sel0_w = main_a7ddrphy_dly_sel_storage[1:0];
assign builder_basesoc_csrbankarray_sel = (builder_basesoc_csrbankarray_sram_bus_adr[13:9] == 2'd3);
always @(*) begin
	builder_basesoc_csrbankarray_sram_bus_dat_r <= 8'd0;
	if (builder_basesoc_csrbankarray_sel_r) begin
		builder_basesoc_csrbankarray_sram_bus_dat_r <= builder_basesoc_csrbankarray_dat_r;
	end
end
assign builder_basesoc_csrbankarray_adr = builder_basesoc_csrbankarray_sram_bus_adr[6:0];
assign builder_basesoc_csrbankarray_csrbank2_sel = (builder_basesoc_csrbankarray_interface2_bank_bus_adr[13:9] == 4'd8);
assign builder_basesoc_csrbankarray_csrbank2_dfii_control0_r = builder_basesoc_csrbankarray_interface2_bank_bus_dat_w[3:0];
assign builder_basesoc_csrbankarray_csrbank2_dfii_control0_re = ((builder_basesoc_csrbankarray_csrbank2_sel & builder_basesoc_csrbankarray_interface2_bank_bus_we) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 1'd0));
assign builder_basesoc_csrbankarray_csrbank2_dfii_control0_we = ((builder_basesoc_csrbankarray_csrbank2_sel & (~builder_basesoc_csrbankarray_interface2_bank_bus_we)) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 1'd0));
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi0_command0_r = builder_basesoc_csrbankarray_interface2_bank_bus_dat_w[5:0];
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi0_command0_re = ((builder_basesoc_csrbankarray_csrbank2_sel & builder_basesoc_csrbankarray_interface2_bank_bus_we) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 1'd1));
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi0_command0_we = ((builder_basesoc_csrbankarray_csrbank2_sel & (~builder_basesoc_csrbankarray_interface2_bank_bus_we)) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 1'd1));
assign main_sdram_phaseinjector0_command_issue_r = builder_basesoc_csrbankarray_interface2_bank_bus_dat_w[0];
assign main_sdram_phaseinjector0_command_issue_re = ((builder_basesoc_csrbankarray_csrbank2_sel & builder_basesoc_csrbankarray_interface2_bank_bus_we) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 2'd2));
assign main_sdram_phaseinjector0_command_issue_we = ((builder_basesoc_csrbankarray_csrbank2_sel & (~builder_basesoc_csrbankarray_interface2_bank_bus_we)) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 2'd2));
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi0_address1_r = builder_basesoc_csrbankarray_interface2_bank_bus_dat_w[5:0];
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi0_address1_re = ((builder_basesoc_csrbankarray_csrbank2_sel & builder_basesoc_csrbankarray_interface2_bank_bus_we) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 2'd3));
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi0_address1_we = ((builder_basesoc_csrbankarray_csrbank2_sel & (~builder_basesoc_csrbankarray_interface2_bank_bus_we)) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 2'd3));
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi0_address0_r = builder_basesoc_csrbankarray_interface2_bank_bus_dat_w[7:0];
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi0_address0_re = ((builder_basesoc_csrbankarray_csrbank2_sel & builder_basesoc_csrbankarray_interface2_bank_bus_we) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 3'd4));
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi0_address0_we = ((builder_basesoc_csrbankarray_csrbank2_sel & (~builder_basesoc_csrbankarray_interface2_bank_bus_we)) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 3'd4));
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi0_baddress0_r = builder_basesoc_csrbankarray_interface2_bank_bus_dat_w[2:0];
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi0_baddress0_re = ((builder_basesoc_csrbankarray_csrbank2_sel & builder_basesoc_csrbankarray_interface2_bank_bus_we) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 3'd5));
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi0_baddress0_we = ((builder_basesoc_csrbankarray_csrbank2_sel & (~builder_basesoc_csrbankarray_interface2_bank_bus_we)) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 3'd5));
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi0_wrdata3_r = builder_basesoc_csrbankarray_interface2_bank_bus_dat_w[7:0];
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi0_wrdata3_re = ((builder_basesoc_csrbankarray_csrbank2_sel & builder_basesoc_csrbankarray_interface2_bank_bus_we) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 3'd6));
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi0_wrdata3_we = ((builder_basesoc_csrbankarray_csrbank2_sel & (~builder_basesoc_csrbankarray_interface2_bank_bus_we)) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 3'd6));
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi0_wrdata2_r = builder_basesoc_csrbankarray_interface2_bank_bus_dat_w[7:0];
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi0_wrdata2_re = ((builder_basesoc_csrbankarray_csrbank2_sel & builder_basesoc_csrbankarray_interface2_bank_bus_we) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 3'd7));
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi0_wrdata2_we = ((builder_basesoc_csrbankarray_csrbank2_sel & (~builder_basesoc_csrbankarray_interface2_bank_bus_we)) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 3'd7));
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi0_wrdata1_r = builder_basesoc_csrbankarray_interface2_bank_bus_dat_w[7:0];
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi0_wrdata1_re = ((builder_basesoc_csrbankarray_csrbank2_sel & builder_basesoc_csrbankarray_interface2_bank_bus_we) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 4'd8));
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi0_wrdata1_we = ((builder_basesoc_csrbankarray_csrbank2_sel & (~builder_basesoc_csrbankarray_interface2_bank_bus_we)) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 4'd8));
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi0_wrdata0_r = builder_basesoc_csrbankarray_interface2_bank_bus_dat_w[7:0];
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi0_wrdata0_re = ((builder_basesoc_csrbankarray_csrbank2_sel & builder_basesoc_csrbankarray_interface2_bank_bus_we) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 4'd9));
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi0_wrdata0_we = ((builder_basesoc_csrbankarray_csrbank2_sel & (~builder_basesoc_csrbankarray_interface2_bank_bus_we)) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 4'd9));
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi0_rddata3_r = builder_basesoc_csrbankarray_interface2_bank_bus_dat_w[7:0];
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi0_rddata3_re = ((builder_basesoc_csrbankarray_csrbank2_sel & builder_basesoc_csrbankarray_interface2_bank_bus_we) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 4'd10));
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi0_rddata3_we = ((builder_basesoc_csrbankarray_csrbank2_sel & (~builder_basesoc_csrbankarray_interface2_bank_bus_we)) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 4'd10));
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi0_rddata2_r = builder_basesoc_csrbankarray_interface2_bank_bus_dat_w[7:0];
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi0_rddata2_re = ((builder_basesoc_csrbankarray_csrbank2_sel & builder_basesoc_csrbankarray_interface2_bank_bus_we) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 4'd11));
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi0_rddata2_we = ((builder_basesoc_csrbankarray_csrbank2_sel & (~builder_basesoc_csrbankarray_interface2_bank_bus_we)) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 4'd11));
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi0_rddata1_r = builder_basesoc_csrbankarray_interface2_bank_bus_dat_w[7:0];
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi0_rddata1_re = ((builder_basesoc_csrbankarray_csrbank2_sel & builder_basesoc_csrbankarray_interface2_bank_bus_we) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 4'd12));
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi0_rddata1_we = ((builder_basesoc_csrbankarray_csrbank2_sel & (~builder_basesoc_csrbankarray_interface2_bank_bus_we)) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 4'd12));
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi0_rddata0_r = builder_basesoc_csrbankarray_interface2_bank_bus_dat_w[7:0];
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi0_rddata0_re = ((builder_basesoc_csrbankarray_csrbank2_sel & builder_basesoc_csrbankarray_interface2_bank_bus_we) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 4'd13));
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi0_rddata0_we = ((builder_basesoc_csrbankarray_csrbank2_sel & (~builder_basesoc_csrbankarray_interface2_bank_bus_we)) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 4'd13));
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi1_command0_r = builder_basesoc_csrbankarray_interface2_bank_bus_dat_w[5:0];
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi1_command0_re = ((builder_basesoc_csrbankarray_csrbank2_sel & builder_basesoc_csrbankarray_interface2_bank_bus_we) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 4'd14));
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi1_command0_we = ((builder_basesoc_csrbankarray_csrbank2_sel & (~builder_basesoc_csrbankarray_interface2_bank_bus_we)) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 4'd14));
assign main_sdram_phaseinjector1_command_issue_r = builder_basesoc_csrbankarray_interface2_bank_bus_dat_w[0];
assign main_sdram_phaseinjector1_command_issue_re = ((builder_basesoc_csrbankarray_csrbank2_sel & builder_basesoc_csrbankarray_interface2_bank_bus_we) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 4'd15));
assign main_sdram_phaseinjector1_command_issue_we = ((builder_basesoc_csrbankarray_csrbank2_sel & (~builder_basesoc_csrbankarray_interface2_bank_bus_we)) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 4'd15));
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi1_address1_r = builder_basesoc_csrbankarray_interface2_bank_bus_dat_w[5:0];
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi1_address1_re = ((builder_basesoc_csrbankarray_csrbank2_sel & builder_basesoc_csrbankarray_interface2_bank_bus_we) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 5'd16));
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi1_address1_we = ((builder_basesoc_csrbankarray_csrbank2_sel & (~builder_basesoc_csrbankarray_interface2_bank_bus_we)) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 5'd16));
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi1_address0_r = builder_basesoc_csrbankarray_interface2_bank_bus_dat_w[7:0];
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi1_address0_re = ((builder_basesoc_csrbankarray_csrbank2_sel & builder_basesoc_csrbankarray_interface2_bank_bus_we) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 5'd17));
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi1_address0_we = ((builder_basesoc_csrbankarray_csrbank2_sel & (~builder_basesoc_csrbankarray_interface2_bank_bus_we)) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 5'd17));
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi1_baddress0_r = builder_basesoc_csrbankarray_interface2_bank_bus_dat_w[2:0];
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi1_baddress0_re = ((builder_basesoc_csrbankarray_csrbank2_sel & builder_basesoc_csrbankarray_interface2_bank_bus_we) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 5'd18));
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi1_baddress0_we = ((builder_basesoc_csrbankarray_csrbank2_sel & (~builder_basesoc_csrbankarray_interface2_bank_bus_we)) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 5'd18));
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi1_wrdata3_r = builder_basesoc_csrbankarray_interface2_bank_bus_dat_w[7:0];
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi1_wrdata3_re = ((builder_basesoc_csrbankarray_csrbank2_sel & builder_basesoc_csrbankarray_interface2_bank_bus_we) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 5'd19));
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi1_wrdata3_we = ((builder_basesoc_csrbankarray_csrbank2_sel & (~builder_basesoc_csrbankarray_interface2_bank_bus_we)) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 5'd19));
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi1_wrdata2_r = builder_basesoc_csrbankarray_interface2_bank_bus_dat_w[7:0];
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi1_wrdata2_re = ((builder_basesoc_csrbankarray_csrbank2_sel & builder_basesoc_csrbankarray_interface2_bank_bus_we) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 5'd20));
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi1_wrdata2_we = ((builder_basesoc_csrbankarray_csrbank2_sel & (~builder_basesoc_csrbankarray_interface2_bank_bus_we)) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 5'd20));
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi1_wrdata1_r = builder_basesoc_csrbankarray_interface2_bank_bus_dat_w[7:0];
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi1_wrdata1_re = ((builder_basesoc_csrbankarray_csrbank2_sel & builder_basesoc_csrbankarray_interface2_bank_bus_we) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 5'd21));
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi1_wrdata1_we = ((builder_basesoc_csrbankarray_csrbank2_sel & (~builder_basesoc_csrbankarray_interface2_bank_bus_we)) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 5'd21));
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi1_wrdata0_r = builder_basesoc_csrbankarray_interface2_bank_bus_dat_w[7:0];
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi1_wrdata0_re = ((builder_basesoc_csrbankarray_csrbank2_sel & builder_basesoc_csrbankarray_interface2_bank_bus_we) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 5'd22));
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi1_wrdata0_we = ((builder_basesoc_csrbankarray_csrbank2_sel & (~builder_basesoc_csrbankarray_interface2_bank_bus_we)) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 5'd22));
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi1_rddata3_r = builder_basesoc_csrbankarray_interface2_bank_bus_dat_w[7:0];
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi1_rddata3_re = ((builder_basesoc_csrbankarray_csrbank2_sel & builder_basesoc_csrbankarray_interface2_bank_bus_we) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 5'd23));
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi1_rddata3_we = ((builder_basesoc_csrbankarray_csrbank2_sel & (~builder_basesoc_csrbankarray_interface2_bank_bus_we)) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 5'd23));
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi1_rddata2_r = builder_basesoc_csrbankarray_interface2_bank_bus_dat_w[7:0];
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi1_rddata2_re = ((builder_basesoc_csrbankarray_csrbank2_sel & builder_basesoc_csrbankarray_interface2_bank_bus_we) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 5'd24));
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi1_rddata2_we = ((builder_basesoc_csrbankarray_csrbank2_sel & (~builder_basesoc_csrbankarray_interface2_bank_bus_we)) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 5'd24));
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi1_rddata1_r = builder_basesoc_csrbankarray_interface2_bank_bus_dat_w[7:0];
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi1_rddata1_re = ((builder_basesoc_csrbankarray_csrbank2_sel & builder_basesoc_csrbankarray_interface2_bank_bus_we) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 5'd25));
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi1_rddata1_we = ((builder_basesoc_csrbankarray_csrbank2_sel & (~builder_basesoc_csrbankarray_interface2_bank_bus_we)) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 5'd25));
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi1_rddata0_r = builder_basesoc_csrbankarray_interface2_bank_bus_dat_w[7:0];
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi1_rddata0_re = ((builder_basesoc_csrbankarray_csrbank2_sel & builder_basesoc_csrbankarray_interface2_bank_bus_we) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 5'd26));
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi1_rddata0_we = ((builder_basesoc_csrbankarray_csrbank2_sel & (~builder_basesoc_csrbankarray_interface2_bank_bus_we)) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 5'd26));
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi2_command0_r = builder_basesoc_csrbankarray_interface2_bank_bus_dat_w[5:0];
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi2_command0_re = ((builder_basesoc_csrbankarray_csrbank2_sel & builder_basesoc_csrbankarray_interface2_bank_bus_we) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 5'd27));
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi2_command0_we = ((builder_basesoc_csrbankarray_csrbank2_sel & (~builder_basesoc_csrbankarray_interface2_bank_bus_we)) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 5'd27));
assign main_sdram_phaseinjector2_command_issue_r = builder_basesoc_csrbankarray_interface2_bank_bus_dat_w[0];
assign main_sdram_phaseinjector2_command_issue_re = ((builder_basesoc_csrbankarray_csrbank2_sel & builder_basesoc_csrbankarray_interface2_bank_bus_we) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 5'd28));
assign main_sdram_phaseinjector2_command_issue_we = ((builder_basesoc_csrbankarray_csrbank2_sel & (~builder_basesoc_csrbankarray_interface2_bank_bus_we)) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 5'd28));
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi2_address1_r = builder_basesoc_csrbankarray_interface2_bank_bus_dat_w[5:0];
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi2_address1_re = ((builder_basesoc_csrbankarray_csrbank2_sel & builder_basesoc_csrbankarray_interface2_bank_bus_we) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 5'd29));
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi2_address1_we = ((builder_basesoc_csrbankarray_csrbank2_sel & (~builder_basesoc_csrbankarray_interface2_bank_bus_we)) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 5'd29));
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi2_address0_r = builder_basesoc_csrbankarray_interface2_bank_bus_dat_w[7:0];
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi2_address0_re = ((builder_basesoc_csrbankarray_csrbank2_sel & builder_basesoc_csrbankarray_interface2_bank_bus_we) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 5'd30));
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi2_address0_we = ((builder_basesoc_csrbankarray_csrbank2_sel & (~builder_basesoc_csrbankarray_interface2_bank_bus_we)) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 5'd30));
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi2_baddress0_r = builder_basesoc_csrbankarray_interface2_bank_bus_dat_w[2:0];
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi2_baddress0_re = ((builder_basesoc_csrbankarray_csrbank2_sel & builder_basesoc_csrbankarray_interface2_bank_bus_we) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 5'd31));
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi2_baddress0_we = ((builder_basesoc_csrbankarray_csrbank2_sel & (~builder_basesoc_csrbankarray_interface2_bank_bus_we)) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 5'd31));
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi2_wrdata3_r = builder_basesoc_csrbankarray_interface2_bank_bus_dat_w[7:0];
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi2_wrdata3_re = ((builder_basesoc_csrbankarray_csrbank2_sel & builder_basesoc_csrbankarray_interface2_bank_bus_we) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 6'd32));
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi2_wrdata3_we = ((builder_basesoc_csrbankarray_csrbank2_sel & (~builder_basesoc_csrbankarray_interface2_bank_bus_we)) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 6'd32));
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi2_wrdata2_r = builder_basesoc_csrbankarray_interface2_bank_bus_dat_w[7:0];
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi2_wrdata2_re = ((builder_basesoc_csrbankarray_csrbank2_sel & builder_basesoc_csrbankarray_interface2_bank_bus_we) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 6'd33));
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi2_wrdata2_we = ((builder_basesoc_csrbankarray_csrbank2_sel & (~builder_basesoc_csrbankarray_interface2_bank_bus_we)) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 6'd33));
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi2_wrdata1_r = builder_basesoc_csrbankarray_interface2_bank_bus_dat_w[7:0];
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi2_wrdata1_re = ((builder_basesoc_csrbankarray_csrbank2_sel & builder_basesoc_csrbankarray_interface2_bank_bus_we) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 6'd34));
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi2_wrdata1_we = ((builder_basesoc_csrbankarray_csrbank2_sel & (~builder_basesoc_csrbankarray_interface2_bank_bus_we)) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 6'd34));
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi2_wrdata0_r = builder_basesoc_csrbankarray_interface2_bank_bus_dat_w[7:0];
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi2_wrdata0_re = ((builder_basesoc_csrbankarray_csrbank2_sel & builder_basesoc_csrbankarray_interface2_bank_bus_we) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 6'd35));
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi2_wrdata0_we = ((builder_basesoc_csrbankarray_csrbank2_sel & (~builder_basesoc_csrbankarray_interface2_bank_bus_we)) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 6'd35));
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi2_rddata3_r = builder_basesoc_csrbankarray_interface2_bank_bus_dat_w[7:0];
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi2_rddata3_re = ((builder_basesoc_csrbankarray_csrbank2_sel & builder_basesoc_csrbankarray_interface2_bank_bus_we) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 6'd36));
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi2_rddata3_we = ((builder_basesoc_csrbankarray_csrbank2_sel & (~builder_basesoc_csrbankarray_interface2_bank_bus_we)) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 6'd36));
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi2_rddata2_r = builder_basesoc_csrbankarray_interface2_bank_bus_dat_w[7:0];
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi2_rddata2_re = ((builder_basesoc_csrbankarray_csrbank2_sel & builder_basesoc_csrbankarray_interface2_bank_bus_we) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 6'd37));
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi2_rddata2_we = ((builder_basesoc_csrbankarray_csrbank2_sel & (~builder_basesoc_csrbankarray_interface2_bank_bus_we)) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 6'd37));
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi2_rddata1_r = builder_basesoc_csrbankarray_interface2_bank_bus_dat_w[7:0];
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi2_rddata1_re = ((builder_basesoc_csrbankarray_csrbank2_sel & builder_basesoc_csrbankarray_interface2_bank_bus_we) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 6'd38));
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi2_rddata1_we = ((builder_basesoc_csrbankarray_csrbank2_sel & (~builder_basesoc_csrbankarray_interface2_bank_bus_we)) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 6'd38));
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi2_rddata0_r = builder_basesoc_csrbankarray_interface2_bank_bus_dat_w[7:0];
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi2_rddata0_re = ((builder_basesoc_csrbankarray_csrbank2_sel & builder_basesoc_csrbankarray_interface2_bank_bus_we) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 6'd39));
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi2_rddata0_we = ((builder_basesoc_csrbankarray_csrbank2_sel & (~builder_basesoc_csrbankarray_interface2_bank_bus_we)) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 6'd39));
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi3_command0_r = builder_basesoc_csrbankarray_interface2_bank_bus_dat_w[5:0];
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi3_command0_re = ((builder_basesoc_csrbankarray_csrbank2_sel & builder_basesoc_csrbankarray_interface2_bank_bus_we) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 6'd40));
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi3_command0_we = ((builder_basesoc_csrbankarray_csrbank2_sel & (~builder_basesoc_csrbankarray_interface2_bank_bus_we)) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 6'd40));
assign main_sdram_phaseinjector3_command_issue_r = builder_basesoc_csrbankarray_interface2_bank_bus_dat_w[0];
assign main_sdram_phaseinjector3_command_issue_re = ((builder_basesoc_csrbankarray_csrbank2_sel & builder_basesoc_csrbankarray_interface2_bank_bus_we) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 6'd41));
assign main_sdram_phaseinjector3_command_issue_we = ((builder_basesoc_csrbankarray_csrbank2_sel & (~builder_basesoc_csrbankarray_interface2_bank_bus_we)) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 6'd41));
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi3_address1_r = builder_basesoc_csrbankarray_interface2_bank_bus_dat_w[5:0];
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi3_address1_re = ((builder_basesoc_csrbankarray_csrbank2_sel & builder_basesoc_csrbankarray_interface2_bank_bus_we) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 6'd42));
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi3_address1_we = ((builder_basesoc_csrbankarray_csrbank2_sel & (~builder_basesoc_csrbankarray_interface2_bank_bus_we)) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 6'd42));
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi3_address0_r = builder_basesoc_csrbankarray_interface2_bank_bus_dat_w[7:0];
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi3_address0_re = ((builder_basesoc_csrbankarray_csrbank2_sel & builder_basesoc_csrbankarray_interface2_bank_bus_we) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 6'd43));
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi3_address0_we = ((builder_basesoc_csrbankarray_csrbank2_sel & (~builder_basesoc_csrbankarray_interface2_bank_bus_we)) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 6'd43));
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi3_baddress0_r = builder_basesoc_csrbankarray_interface2_bank_bus_dat_w[2:0];
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi3_baddress0_re = ((builder_basesoc_csrbankarray_csrbank2_sel & builder_basesoc_csrbankarray_interface2_bank_bus_we) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 6'd44));
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi3_baddress0_we = ((builder_basesoc_csrbankarray_csrbank2_sel & (~builder_basesoc_csrbankarray_interface2_bank_bus_we)) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 6'd44));
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi3_wrdata3_r = builder_basesoc_csrbankarray_interface2_bank_bus_dat_w[7:0];
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi3_wrdata3_re = ((builder_basesoc_csrbankarray_csrbank2_sel & builder_basesoc_csrbankarray_interface2_bank_bus_we) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 6'd45));
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi3_wrdata3_we = ((builder_basesoc_csrbankarray_csrbank2_sel & (~builder_basesoc_csrbankarray_interface2_bank_bus_we)) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 6'd45));
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi3_wrdata2_r = builder_basesoc_csrbankarray_interface2_bank_bus_dat_w[7:0];
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi3_wrdata2_re = ((builder_basesoc_csrbankarray_csrbank2_sel & builder_basesoc_csrbankarray_interface2_bank_bus_we) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 6'd46));
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi3_wrdata2_we = ((builder_basesoc_csrbankarray_csrbank2_sel & (~builder_basesoc_csrbankarray_interface2_bank_bus_we)) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 6'd46));
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi3_wrdata1_r = builder_basesoc_csrbankarray_interface2_bank_bus_dat_w[7:0];
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi3_wrdata1_re = ((builder_basesoc_csrbankarray_csrbank2_sel & builder_basesoc_csrbankarray_interface2_bank_bus_we) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 6'd47));
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi3_wrdata1_we = ((builder_basesoc_csrbankarray_csrbank2_sel & (~builder_basesoc_csrbankarray_interface2_bank_bus_we)) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 6'd47));
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi3_wrdata0_r = builder_basesoc_csrbankarray_interface2_bank_bus_dat_w[7:0];
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi3_wrdata0_re = ((builder_basesoc_csrbankarray_csrbank2_sel & builder_basesoc_csrbankarray_interface2_bank_bus_we) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 6'd48));
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi3_wrdata0_we = ((builder_basesoc_csrbankarray_csrbank2_sel & (~builder_basesoc_csrbankarray_interface2_bank_bus_we)) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 6'd48));
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi3_rddata3_r = builder_basesoc_csrbankarray_interface2_bank_bus_dat_w[7:0];
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi3_rddata3_re = ((builder_basesoc_csrbankarray_csrbank2_sel & builder_basesoc_csrbankarray_interface2_bank_bus_we) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 6'd49));
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi3_rddata3_we = ((builder_basesoc_csrbankarray_csrbank2_sel & (~builder_basesoc_csrbankarray_interface2_bank_bus_we)) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 6'd49));
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi3_rddata2_r = builder_basesoc_csrbankarray_interface2_bank_bus_dat_w[7:0];
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi3_rddata2_re = ((builder_basesoc_csrbankarray_csrbank2_sel & builder_basesoc_csrbankarray_interface2_bank_bus_we) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 6'd50));
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi3_rddata2_we = ((builder_basesoc_csrbankarray_csrbank2_sel & (~builder_basesoc_csrbankarray_interface2_bank_bus_we)) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 6'd50));
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi3_rddata1_r = builder_basesoc_csrbankarray_interface2_bank_bus_dat_w[7:0];
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi3_rddata1_re = ((builder_basesoc_csrbankarray_csrbank2_sel & builder_basesoc_csrbankarray_interface2_bank_bus_we) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 6'd51));
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi3_rddata1_we = ((builder_basesoc_csrbankarray_csrbank2_sel & (~builder_basesoc_csrbankarray_interface2_bank_bus_we)) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 6'd51));
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi3_rddata0_r = builder_basesoc_csrbankarray_interface2_bank_bus_dat_w[7:0];
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi3_rddata0_re = ((builder_basesoc_csrbankarray_csrbank2_sel & builder_basesoc_csrbankarray_interface2_bank_bus_we) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 6'd52));
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi3_rddata0_we = ((builder_basesoc_csrbankarray_csrbank2_sel & (~builder_basesoc_csrbankarray_interface2_bank_bus_we)) & (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0] == 6'd52));
assign builder_basesoc_csrbankarray_csrbank2_dfii_control0_w = main_sdram_storage[3:0];
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi0_command0_w = main_sdram_phaseinjector0_command_storage[5:0];
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi0_address1_w = main_sdram_phaseinjector0_address_storage[13:8];
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi0_address0_w = main_sdram_phaseinjector0_address_storage[7:0];
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi0_baddress0_w = main_sdram_phaseinjector0_baddress_storage[2:0];
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi0_wrdata3_w = main_sdram_phaseinjector0_wrdata_storage[31:24];
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi0_wrdata2_w = main_sdram_phaseinjector0_wrdata_storage[23:16];
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi0_wrdata1_w = main_sdram_phaseinjector0_wrdata_storage[15:8];
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi0_wrdata0_w = main_sdram_phaseinjector0_wrdata_storage[7:0];
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi0_rddata3_w = main_sdram_phaseinjector0_status[31:24];
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi0_rddata2_w = main_sdram_phaseinjector0_status[23:16];
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi0_rddata1_w = main_sdram_phaseinjector0_status[15:8];
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi0_rddata0_w = main_sdram_phaseinjector0_status[7:0];
assign main_sdram_phaseinjector0_we = builder_basesoc_csrbankarray_csrbank2_dfii_pi0_rddata0_we;
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi1_command0_w = main_sdram_phaseinjector1_command_storage[5:0];
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi1_address1_w = main_sdram_phaseinjector1_address_storage[13:8];
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi1_address0_w = main_sdram_phaseinjector1_address_storage[7:0];
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi1_baddress0_w = main_sdram_phaseinjector1_baddress_storage[2:0];
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi1_wrdata3_w = main_sdram_phaseinjector1_wrdata_storage[31:24];
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi1_wrdata2_w = main_sdram_phaseinjector1_wrdata_storage[23:16];
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi1_wrdata1_w = main_sdram_phaseinjector1_wrdata_storage[15:8];
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi1_wrdata0_w = main_sdram_phaseinjector1_wrdata_storage[7:0];
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi1_rddata3_w = main_sdram_phaseinjector1_status[31:24];
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi1_rddata2_w = main_sdram_phaseinjector1_status[23:16];
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi1_rddata1_w = main_sdram_phaseinjector1_status[15:8];
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi1_rddata0_w = main_sdram_phaseinjector1_status[7:0];
assign main_sdram_phaseinjector1_we = builder_basesoc_csrbankarray_csrbank2_dfii_pi1_rddata0_we;
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi2_command0_w = main_sdram_phaseinjector2_command_storage[5:0];
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi2_address1_w = main_sdram_phaseinjector2_address_storage[13:8];
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi2_address0_w = main_sdram_phaseinjector2_address_storage[7:0];
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi2_baddress0_w = main_sdram_phaseinjector2_baddress_storage[2:0];
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi2_wrdata3_w = main_sdram_phaseinjector2_wrdata_storage[31:24];
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi2_wrdata2_w = main_sdram_phaseinjector2_wrdata_storage[23:16];
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi2_wrdata1_w = main_sdram_phaseinjector2_wrdata_storage[15:8];
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi2_wrdata0_w = main_sdram_phaseinjector2_wrdata_storage[7:0];
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi2_rddata3_w = main_sdram_phaseinjector2_status[31:24];
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi2_rddata2_w = main_sdram_phaseinjector2_status[23:16];
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi2_rddata1_w = main_sdram_phaseinjector2_status[15:8];
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi2_rddata0_w = main_sdram_phaseinjector2_status[7:0];
assign main_sdram_phaseinjector2_we = builder_basesoc_csrbankarray_csrbank2_dfii_pi2_rddata0_we;
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi3_command0_w = main_sdram_phaseinjector3_command_storage[5:0];
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi3_address1_w = main_sdram_phaseinjector3_address_storage[13:8];
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi3_address0_w = main_sdram_phaseinjector3_address_storage[7:0];
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi3_baddress0_w = main_sdram_phaseinjector3_baddress_storage[2:0];
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi3_wrdata3_w = main_sdram_phaseinjector3_wrdata_storage[31:24];
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi3_wrdata2_w = main_sdram_phaseinjector3_wrdata_storage[23:16];
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi3_wrdata1_w = main_sdram_phaseinjector3_wrdata_storage[15:8];
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi3_wrdata0_w = main_sdram_phaseinjector3_wrdata_storage[7:0];
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi3_rddata3_w = main_sdram_phaseinjector3_status[31:24];
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi3_rddata2_w = main_sdram_phaseinjector3_status[23:16];
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi3_rddata1_w = main_sdram_phaseinjector3_status[15:8];
assign builder_basesoc_csrbankarray_csrbank2_dfii_pi3_rddata0_w = main_sdram_phaseinjector3_status[7:0];
assign main_sdram_phaseinjector3_we = builder_basesoc_csrbankarray_csrbank2_dfii_pi3_rddata0_we;
assign builder_basesoc_csrbankarray_csrbank3_sel = (builder_basesoc_csrbankarray_interface3_bank_bus_adr[13:9] == 3'd4);
assign builder_basesoc_csrbankarray_csrbank3_load3_r = builder_basesoc_csrbankarray_interface3_bank_bus_dat_w[7:0];
assign builder_basesoc_csrbankarray_csrbank3_load3_re = ((builder_basesoc_csrbankarray_csrbank3_sel & builder_basesoc_csrbankarray_interface3_bank_bus_we) & (builder_basesoc_csrbankarray_interface3_bank_bus_adr[4:0] == 1'd0));
assign builder_basesoc_csrbankarray_csrbank3_load3_we = ((builder_basesoc_csrbankarray_csrbank3_sel & (~builder_basesoc_csrbankarray_interface3_bank_bus_we)) & (builder_basesoc_csrbankarray_interface3_bank_bus_adr[4:0] == 1'd0));
assign builder_basesoc_csrbankarray_csrbank3_load2_r = builder_basesoc_csrbankarray_interface3_bank_bus_dat_w[7:0];
assign builder_basesoc_csrbankarray_csrbank3_load2_re = ((builder_basesoc_csrbankarray_csrbank3_sel & builder_basesoc_csrbankarray_interface3_bank_bus_we) & (builder_basesoc_csrbankarray_interface3_bank_bus_adr[4:0] == 1'd1));
assign builder_basesoc_csrbankarray_csrbank3_load2_we = ((builder_basesoc_csrbankarray_csrbank3_sel & (~builder_basesoc_csrbankarray_interface3_bank_bus_we)) & (builder_basesoc_csrbankarray_interface3_bank_bus_adr[4:0] == 1'd1));
assign builder_basesoc_csrbankarray_csrbank3_load1_r = builder_basesoc_csrbankarray_interface3_bank_bus_dat_w[7:0];
assign builder_basesoc_csrbankarray_csrbank3_load1_re = ((builder_basesoc_csrbankarray_csrbank3_sel & builder_basesoc_csrbankarray_interface3_bank_bus_we) & (builder_basesoc_csrbankarray_interface3_bank_bus_adr[4:0] == 2'd2));
assign builder_basesoc_csrbankarray_csrbank3_load1_we = ((builder_basesoc_csrbankarray_csrbank3_sel & (~builder_basesoc_csrbankarray_interface3_bank_bus_we)) & (builder_basesoc_csrbankarray_interface3_bank_bus_adr[4:0] == 2'd2));
assign builder_basesoc_csrbankarray_csrbank3_load0_r = builder_basesoc_csrbankarray_interface3_bank_bus_dat_w[7:0];
assign builder_basesoc_csrbankarray_csrbank3_load0_re = ((builder_basesoc_csrbankarray_csrbank3_sel & builder_basesoc_csrbankarray_interface3_bank_bus_we) & (builder_basesoc_csrbankarray_interface3_bank_bus_adr[4:0] == 2'd3));
assign builder_basesoc_csrbankarray_csrbank3_load0_we = ((builder_basesoc_csrbankarray_csrbank3_sel & (~builder_basesoc_csrbankarray_interface3_bank_bus_we)) & (builder_basesoc_csrbankarray_interface3_bank_bus_adr[4:0] == 2'd3));
assign builder_basesoc_csrbankarray_csrbank3_reload3_r = builder_basesoc_csrbankarray_interface3_bank_bus_dat_w[7:0];
assign builder_basesoc_csrbankarray_csrbank3_reload3_re = ((builder_basesoc_csrbankarray_csrbank3_sel & builder_basesoc_csrbankarray_interface3_bank_bus_we) & (builder_basesoc_csrbankarray_interface3_bank_bus_adr[4:0] == 3'd4));
assign builder_basesoc_csrbankarray_csrbank3_reload3_we = ((builder_basesoc_csrbankarray_csrbank3_sel & (~builder_basesoc_csrbankarray_interface3_bank_bus_we)) & (builder_basesoc_csrbankarray_interface3_bank_bus_adr[4:0] == 3'd4));
assign builder_basesoc_csrbankarray_csrbank3_reload2_r = builder_basesoc_csrbankarray_interface3_bank_bus_dat_w[7:0];
assign builder_basesoc_csrbankarray_csrbank3_reload2_re = ((builder_basesoc_csrbankarray_csrbank3_sel & builder_basesoc_csrbankarray_interface3_bank_bus_we) & (builder_basesoc_csrbankarray_interface3_bank_bus_adr[4:0] == 3'd5));
assign builder_basesoc_csrbankarray_csrbank3_reload2_we = ((builder_basesoc_csrbankarray_csrbank3_sel & (~builder_basesoc_csrbankarray_interface3_bank_bus_we)) & (builder_basesoc_csrbankarray_interface3_bank_bus_adr[4:0] == 3'd5));
assign builder_basesoc_csrbankarray_csrbank3_reload1_r = builder_basesoc_csrbankarray_interface3_bank_bus_dat_w[7:0];
assign builder_basesoc_csrbankarray_csrbank3_reload1_re = ((builder_basesoc_csrbankarray_csrbank3_sel & builder_basesoc_csrbankarray_interface3_bank_bus_we) & (builder_basesoc_csrbankarray_interface3_bank_bus_adr[4:0] == 3'd6));
assign builder_basesoc_csrbankarray_csrbank3_reload1_we = ((builder_basesoc_csrbankarray_csrbank3_sel & (~builder_basesoc_csrbankarray_interface3_bank_bus_we)) & (builder_basesoc_csrbankarray_interface3_bank_bus_adr[4:0] == 3'd6));
assign builder_basesoc_csrbankarray_csrbank3_reload0_r = builder_basesoc_csrbankarray_interface3_bank_bus_dat_w[7:0];
assign builder_basesoc_csrbankarray_csrbank3_reload0_re = ((builder_basesoc_csrbankarray_csrbank3_sel & builder_basesoc_csrbankarray_interface3_bank_bus_we) & (builder_basesoc_csrbankarray_interface3_bank_bus_adr[4:0] == 3'd7));
assign builder_basesoc_csrbankarray_csrbank3_reload0_we = ((builder_basesoc_csrbankarray_csrbank3_sel & (~builder_basesoc_csrbankarray_interface3_bank_bus_we)) & (builder_basesoc_csrbankarray_interface3_bank_bus_adr[4:0] == 3'd7));
assign builder_basesoc_csrbankarray_csrbank3_en0_r = builder_basesoc_csrbankarray_interface3_bank_bus_dat_w[0];
assign builder_basesoc_csrbankarray_csrbank3_en0_re = ((builder_basesoc_csrbankarray_csrbank3_sel & builder_basesoc_csrbankarray_interface3_bank_bus_we) & (builder_basesoc_csrbankarray_interface3_bank_bus_adr[4:0] == 4'd8));
assign builder_basesoc_csrbankarray_csrbank3_en0_we = ((builder_basesoc_csrbankarray_csrbank3_sel & (~builder_basesoc_csrbankarray_interface3_bank_bus_we)) & (builder_basesoc_csrbankarray_interface3_bank_bus_adr[4:0] == 4'd8));
assign builder_basesoc_csrbankarray_csrbank3_update_value0_r = builder_basesoc_csrbankarray_interface3_bank_bus_dat_w[0];
assign builder_basesoc_csrbankarray_csrbank3_update_value0_re = ((builder_basesoc_csrbankarray_csrbank3_sel & builder_basesoc_csrbankarray_interface3_bank_bus_we) & (builder_basesoc_csrbankarray_interface3_bank_bus_adr[4:0] == 4'd9));
assign builder_basesoc_csrbankarray_csrbank3_update_value0_we = ((builder_basesoc_csrbankarray_csrbank3_sel & (~builder_basesoc_csrbankarray_interface3_bank_bus_we)) & (builder_basesoc_csrbankarray_interface3_bank_bus_adr[4:0] == 4'd9));
assign builder_basesoc_csrbankarray_csrbank3_value3_r = builder_basesoc_csrbankarray_interface3_bank_bus_dat_w[7:0];
assign builder_basesoc_csrbankarray_csrbank3_value3_re = ((builder_basesoc_csrbankarray_csrbank3_sel & builder_basesoc_csrbankarray_interface3_bank_bus_we) & (builder_basesoc_csrbankarray_interface3_bank_bus_adr[4:0] == 4'd10));
assign builder_basesoc_csrbankarray_csrbank3_value3_we = ((builder_basesoc_csrbankarray_csrbank3_sel & (~builder_basesoc_csrbankarray_interface3_bank_bus_we)) & (builder_basesoc_csrbankarray_interface3_bank_bus_adr[4:0] == 4'd10));
assign builder_basesoc_csrbankarray_csrbank3_value2_r = builder_basesoc_csrbankarray_interface3_bank_bus_dat_w[7:0];
assign builder_basesoc_csrbankarray_csrbank3_value2_re = ((builder_basesoc_csrbankarray_csrbank3_sel & builder_basesoc_csrbankarray_interface3_bank_bus_we) & (builder_basesoc_csrbankarray_interface3_bank_bus_adr[4:0] == 4'd11));
assign builder_basesoc_csrbankarray_csrbank3_value2_we = ((builder_basesoc_csrbankarray_csrbank3_sel & (~builder_basesoc_csrbankarray_interface3_bank_bus_we)) & (builder_basesoc_csrbankarray_interface3_bank_bus_adr[4:0] == 4'd11));
assign builder_basesoc_csrbankarray_csrbank3_value1_r = builder_basesoc_csrbankarray_interface3_bank_bus_dat_w[7:0];
assign builder_basesoc_csrbankarray_csrbank3_value1_re = ((builder_basesoc_csrbankarray_csrbank3_sel & builder_basesoc_csrbankarray_interface3_bank_bus_we) & (builder_basesoc_csrbankarray_interface3_bank_bus_adr[4:0] == 4'd12));
assign builder_basesoc_csrbankarray_csrbank3_value1_we = ((builder_basesoc_csrbankarray_csrbank3_sel & (~builder_basesoc_csrbankarray_interface3_bank_bus_we)) & (builder_basesoc_csrbankarray_interface3_bank_bus_adr[4:0] == 4'd12));
assign builder_basesoc_csrbankarray_csrbank3_value0_r = builder_basesoc_csrbankarray_interface3_bank_bus_dat_w[7:0];
assign builder_basesoc_csrbankarray_csrbank3_value0_re = ((builder_basesoc_csrbankarray_csrbank3_sel & builder_basesoc_csrbankarray_interface3_bank_bus_we) & (builder_basesoc_csrbankarray_interface3_bank_bus_adr[4:0] == 4'd13));
assign builder_basesoc_csrbankarray_csrbank3_value0_we = ((builder_basesoc_csrbankarray_csrbank3_sel & (~builder_basesoc_csrbankarray_interface3_bank_bus_we)) & (builder_basesoc_csrbankarray_interface3_bank_bus_adr[4:0] == 4'd13));
assign main_eventmanager_status_r = builder_basesoc_csrbankarray_interface3_bank_bus_dat_w[0];
assign main_eventmanager_status_re = ((builder_basesoc_csrbankarray_csrbank3_sel & builder_basesoc_csrbankarray_interface3_bank_bus_we) & (builder_basesoc_csrbankarray_interface3_bank_bus_adr[4:0] == 4'd14));
assign main_eventmanager_status_we = ((builder_basesoc_csrbankarray_csrbank3_sel & (~builder_basesoc_csrbankarray_interface3_bank_bus_we)) & (builder_basesoc_csrbankarray_interface3_bank_bus_adr[4:0] == 4'd14));
assign main_eventmanager_pending_r = builder_basesoc_csrbankarray_interface3_bank_bus_dat_w[0];
assign main_eventmanager_pending_re = ((builder_basesoc_csrbankarray_csrbank3_sel & builder_basesoc_csrbankarray_interface3_bank_bus_we) & (builder_basesoc_csrbankarray_interface3_bank_bus_adr[4:0] == 4'd15));
assign main_eventmanager_pending_we = ((builder_basesoc_csrbankarray_csrbank3_sel & (~builder_basesoc_csrbankarray_interface3_bank_bus_we)) & (builder_basesoc_csrbankarray_interface3_bank_bus_adr[4:0] == 4'd15));
assign builder_basesoc_csrbankarray_csrbank3_ev_enable0_r = builder_basesoc_csrbankarray_interface3_bank_bus_dat_w[0];
assign builder_basesoc_csrbankarray_csrbank3_ev_enable0_re = ((builder_basesoc_csrbankarray_csrbank3_sel & builder_basesoc_csrbankarray_interface3_bank_bus_we) & (builder_basesoc_csrbankarray_interface3_bank_bus_adr[4:0] == 5'd16));
assign builder_basesoc_csrbankarray_csrbank3_ev_enable0_we = ((builder_basesoc_csrbankarray_csrbank3_sel & (~builder_basesoc_csrbankarray_interface3_bank_bus_we)) & (builder_basesoc_csrbankarray_interface3_bank_bus_adr[4:0] == 5'd16));
assign builder_basesoc_csrbankarray_csrbank3_load3_w = main_load_storage[31:24];
assign builder_basesoc_csrbankarray_csrbank3_load2_w = main_load_storage[23:16];
assign builder_basesoc_csrbankarray_csrbank3_load1_w = main_load_storage[15:8];
assign builder_basesoc_csrbankarray_csrbank3_load0_w = main_load_storage[7:0];
assign builder_basesoc_csrbankarray_csrbank3_reload3_w = main_reload_storage[31:24];
assign builder_basesoc_csrbankarray_csrbank3_reload2_w = main_reload_storage[23:16];
assign builder_basesoc_csrbankarray_csrbank3_reload1_w = main_reload_storage[15:8];
assign builder_basesoc_csrbankarray_csrbank3_reload0_w = main_reload_storage[7:0];
assign builder_basesoc_csrbankarray_csrbank3_en0_w = main_en_storage;
assign builder_basesoc_csrbankarray_csrbank3_update_value0_w = main_update_value_storage;
assign builder_basesoc_csrbankarray_csrbank3_value3_w = main_value_status[31:24];
assign builder_basesoc_csrbankarray_csrbank3_value2_w = main_value_status[23:16];
assign builder_basesoc_csrbankarray_csrbank3_value1_w = main_value_status[15:8];
assign builder_basesoc_csrbankarray_csrbank3_value0_w = main_value_status[7:0];
assign main_value_we = builder_basesoc_csrbankarray_csrbank3_value0_we;
assign builder_basesoc_csrbankarray_csrbank3_ev_enable0_w = main_eventmanager_storage;
assign builder_basesoc_csrcon_adr = main_interface_adr;
assign builder_basesoc_csrcon_we = main_interface_we;
assign builder_basesoc_csrcon_dat_w = main_interface_dat_w;
assign main_interface_dat_r = builder_basesoc_csrcon_dat_r;
assign builder_basesoc_csrbankarray_interface0_bank_bus_adr = builder_basesoc_csrcon_adr;
assign builder_basesoc_csrbankarray_interface1_bank_bus_adr = builder_basesoc_csrcon_adr;
assign builder_basesoc_csrbankarray_interface2_bank_bus_adr = builder_basesoc_csrcon_adr;
assign builder_basesoc_csrbankarray_interface3_bank_bus_adr = builder_basesoc_csrcon_adr;
assign builder_basesoc_csrbankarray_sram_bus_adr = builder_basesoc_csrcon_adr;
assign builder_basesoc_csrbankarray_interface0_bank_bus_we = builder_basesoc_csrcon_we;
assign builder_basesoc_csrbankarray_interface1_bank_bus_we = builder_basesoc_csrcon_we;
assign builder_basesoc_csrbankarray_interface2_bank_bus_we = builder_basesoc_csrcon_we;
assign builder_basesoc_csrbankarray_interface3_bank_bus_we = builder_basesoc_csrcon_we;
assign builder_basesoc_csrbankarray_sram_bus_we = builder_basesoc_csrcon_we;
assign builder_basesoc_csrbankarray_interface0_bank_bus_dat_w = builder_basesoc_csrcon_dat_w;
assign builder_basesoc_csrbankarray_interface1_bank_bus_dat_w = builder_basesoc_csrcon_dat_w;
assign builder_basesoc_csrbankarray_interface2_bank_bus_dat_w = builder_basesoc_csrcon_dat_w;
assign builder_basesoc_csrbankarray_interface3_bank_bus_dat_w = builder_basesoc_csrcon_dat_w;
assign builder_basesoc_csrbankarray_sram_bus_dat_w = builder_basesoc_csrcon_dat_w;
assign builder_basesoc_csrcon_dat_r = ((((builder_basesoc_csrbankarray_interface0_bank_bus_dat_r | builder_basesoc_csrbankarray_interface1_bank_bus_dat_r) | builder_basesoc_csrbankarray_interface2_bank_bus_dat_r) | builder_basesoc_csrbankarray_interface3_bank_bus_dat_r) | builder_basesoc_csrbankarray_sram_bus_dat_r);
always @(*) begin
	builder_rhs_array_muxed0 <= 1'd0;
	case (main_sdram_choose_cmd_grant)
		1'd0: begin
			builder_rhs_array_muxed0 <= main_sdram_choose_cmd_valids[0];
		end
		1'd1: begin
			builder_rhs_array_muxed0 <= main_sdram_choose_cmd_valids[1];
		end
		2'd2: begin
			builder_rhs_array_muxed0 <= main_sdram_choose_cmd_valids[2];
		end
		2'd3: begin
			builder_rhs_array_muxed0 <= main_sdram_choose_cmd_valids[3];
		end
		3'd4: begin
			builder_rhs_array_muxed0 <= main_sdram_choose_cmd_valids[4];
		end
		3'd5: begin
			builder_rhs_array_muxed0 <= main_sdram_choose_cmd_valids[5];
		end
		3'd6: begin
			builder_rhs_array_muxed0 <= main_sdram_choose_cmd_valids[6];
		end
		default: begin
			builder_rhs_array_muxed0 <= main_sdram_choose_cmd_valids[7];
		end
	endcase
end
always @(*) begin
	builder_rhs_array_muxed1 <= 14'd0;
	case (main_sdram_choose_cmd_grant)
		1'd0: begin
			builder_rhs_array_muxed1 <= main_sdram_bankmachine0_cmd_payload_a;
		end
		1'd1: begin
			builder_rhs_array_muxed1 <= main_sdram_bankmachine1_cmd_payload_a;
		end
		2'd2: begin
			builder_rhs_array_muxed1 <= main_sdram_bankmachine2_cmd_payload_a;
		end
		2'd3: begin
			builder_rhs_array_muxed1 <= main_sdram_bankmachine3_cmd_payload_a;
		end
		3'd4: begin
			builder_rhs_array_muxed1 <= main_sdram_bankmachine4_cmd_payload_a;
		end
		3'd5: begin
			builder_rhs_array_muxed1 <= main_sdram_bankmachine5_cmd_payload_a;
		end
		3'd6: begin
			builder_rhs_array_muxed1 <= main_sdram_bankmachine6_cmd_payload_a;
		end
		default: begin
			builder_rhs_array_muxed1 <= main_sdram_bankmachine7_cmd_payload_a;
		end
	endcase
end
always @(*) begin
	builder_rhs_array_muxed2 <= 3'd0;
	case (main_sdram_choose_cmd_grant)
		1'd0: begin
			builder_rhs_array_muxed2 <= main_sdram_bankmachine0_cmd_payload_ba;
		end
		1'd1: begin
			builder_rhs_array_muxed2 <= main_sdram_bankmachine1_cmd_payload_ba;
		end
		2'd2: begin
			builder_rhs_array_muxed2 <= main_sdram_bankmachine2_cmd_payload_ba;
		end
		2'd3: begin
			builder_rhs_array_muxed2 <= main_sdram_bankmachine3_cmd_payload_ba;
		end
		3'd4: begin
			builder_rhs_array_muxed2 <= main_sdram_bankmachine4_cmd_payload_ba;
		end
		3'd5: begin
			builder_rhs_array_muxed2 <= main_sdram_bankmachine5_cmd_payload_ba;
		end
		3'd6: begin
			builder_rhs_array_muxed2 <= main_sdram_bankmachine6_cmd_payload_ba;
		end
		default: begin
			builder_rhs_array_muxed2 <= main_sdram_bankmachine7_cmd_payload_ba;
		end
	endcase
end
always @(*) begin
	builder_rhs_array_muxed3 <= 1'd0;
	case (main_sdram_choose_cmd_grant)
		1'd0: begin
			builder_rhs_array_muxed3 <= main_sdram_bankmachine0_cmd_payload_is_read;
		end
		1'd1: begin
			builder_rhs_array_muxed3 <= main_sdram_bankmachine1_cmd_payload_is_read;
		end
		2'd2: begin
			builder_rhs_array_muxed3 <= main_sdram_bankmachine2_cmd_payload_is_read;
		end
		2'd3: begin
			builder_rhs_array_muxed3 <= main_sdram_bankmachine3_cmd_payload_is_read;
		end
		3'd4: begin
			builder_rhs_array_muxed3 <= main_sdram_bankmachine4_cmd_payload_is_read;
		end
		3'd5: begin
			builder_rhs_array_muxed3 <= main_sdram_bankmachine5_cmd_payload_is_read;
		end
		3'd6: begin
			builder_rhs_array_muxed3 <= main_sdram_bankmachine6_cmd_payload_is_read;
		end
		default: begin
			builder_rhs_array_muxed3 <= main_sdram_bankmachine7_cmd_payload_is_read;
		end
	endcase
end
always @(*) begin
	builder_rhs_array_muxed4 <= 1'd0;
	case (main_sdram_choose_cmd_grant)
		1'd0: begin
			builder_rhs_array_muxed4 <= main_sdram_bankmachine0_cmd_payload_is_write;
		end
		1'd1: begin
			builder_rhs_array_muxed4 <= main_sdram_bankmachine1_cmd_payload_is_write;
		end
		2'd2: begin
			builder_rhs_array_muxed4 <= main_sdram_bankmachine2_cmd_payload_is_write;
		end
		2'd3: begin
			builder_rhs_array_muxed4 <= main_sdram_bankmachine3_cmd_payload_is_write;
		end
		3'd4: begin
			builder_rhs_array_muxed4 <= main_sdram_bankmachine4_cmd_payload_is_write;
		end
		3'd5: begin
			builder_rhs_array_muxed4 <= main_sdram_bankmachine5_cmd_payload_is_write;
		end
		3'd6: begin
			builder_rhs_array_muxed4 <= main_sdram_bankmachine6_cmd_payload_is_write;
		end
		default: begin
			builder_rhs_array_muxed4 <= main_sdram_bankmachine7_cmd_payload_is_write;
		end
	endcase
end
always @(*) begin
	builder_rhs_array_muxed5 <= 1'd0;
	case (main_sdram_choose_cmd_grant)
		1'd0: begin
			builder_rhs_array_muxed5 <= main_sdram_bankmachine0_cmd_payload_is_cmd;
		end
		1'd1: begin
			builder_rhs_array_muxed5 <= main_sdram_bankmachine1_cmd_payload_is_cmd;
		end
		2'd2: begin
			builder_rhs_array_muxed5 <= main_sdram_bankmachine2_cmd_payload_is_cmd;
		end
		2'd3: begin
			builder_rhs_array_muxed5 <= main_sdram_bankmachine3_cmd_payload_is_cmd;
		end
		3'd4: begin
			builder_rhs_array_muxed5 <= main_sdram_bankmachine4_cmd_payload_is_cmd;
		end
		3'd5: begin
			builder_rhs_array_muxed5 <= main_sdram_bankmachine5_cmd_payload_is_cmd;
		end
		3'd6: begin
			builder_rhs_array_muxed5 <= main_sdram_bankmachine6_cmd_payload_is_cmd;
		end
		default: begin
			builder_rhs_array_muxed5 <= main_sdram_bankmachine7_cmd_payload_is_cmd;
		end
	endcase
end
always @(*) begin
	builder_t_array_muxed0 <= 1'd0;
	case (main_sdram_choose_cmd_grant)
		1'd0: begin
			builder_t_array_muxed0 <= main_sdram_bankmachine0_cmd_payload_cas;
		end
		1'd1: begin
			builder_t_array_muxed0 <= main_sdram_bankmachine1_cmd_payload_cas;
		end
		2'd2: begin
			builder_t_array_muxed0 <= main_sdram_bankmachine2_cmd_payload_cas;
		end
		2'd3: begin
			builder_t_array_muxed0 <= main_sdram_bankmachine3_cmd_payload_cas;
		end
		3'd4: begin
			builder_t_array_muxed0 <= main_sdram_bankmachine4_cmd_payload_cas;
		end
		3'd5: begin
			builder_t_array_muxed0 <= main_sdram_bankmachine5_cmd_payload_cas;
		end
		3'd6: begin
			builder_t_array_muxed0 <= main_sdram_bankmachine6_cmd_payload_cas;
		end
		default: begin
			builder_t_array_muxed0 <= main_sdram_bankmachine7_cmd_payload_cas;
		end
	endcase
end
always @(*) begin
	builder_t_array_muxed1 <= 1'd0;
	case (main_sdram_choose_cmd_grant)
		1'd0: begin
			builder_t_array_muxed1 <= main_sdram_bankmachine0_cmd_payload_ras;
		end
		1'd1: begin
			builder_t_array_muxed1 <= main_sdram_bankmachine1_cmd_payload_ras;
		end
		2'd2: begin
			builder_t_array_muxed1 <= main_sdram_bankmachine2_cmd_payload_ras;
		end
		2'd3: begin
			builder_t_array_muxed1 <= main_sdram_bankmachine3_cmd_payload_ras;
		end
		3'd4: begin
			builder_t_array_muxed1 <= main_sdram_bankmachine4_cmd_payload_ras;
		end
		3'd5: begin
			builder_t_array_muxed1 <= main_sdram_bankmachine5_cmd_payload_ras;
		end
		3'd6: begin
			builder_t_array_muxed1 <= main_sdram_bankmachine6_cmd_payload_ras;
		end
		default: begin
			builder_t_array_muxed1 <= main_sdram_bankmachine7_cmd_payload_ras;
		end
	endcase
end
always @(*) begin
	builder_t_array_muxed2 <= 1'd0;
	case (main_sdram_choose_cmd_grant)
		1'd0: begin
			builder_t_array_muxed2 <= main_sdram_bankmachine0_cmd_payload_we;
		end
		1'd1: begin
			builder_t_array_muxed2 <= main_sdram_bankmachine1_cmd_payload_we;
		end
		2'd2: begin
			builder_t_array_muxed2 <= main_sdram_bankmachine2_cmd_payload_we;
		end
		2'd3: begin
			builder_t_array_muxed2 <= main_sdram_bankmachine3_cmd_payload_we;
		end
		3'd4: begin
			builder_t_array_muxed2 <= main_sdram_bankmachine4_cmd_payload_we;
		end
		3'd5: begin
			builder_t_array_muxed2 <= main_sdram_bankmachine5_cmd_payload_we;
		end
		3'd6: begin
			builder_t_array_muxed2 <= main_sdram_bankmachine6_cmd_payload_we;
		end
		default: begin
			builder_t_array_muxed2 <= main_sdram_bankmachine7_cmd_payload_we;
		end
	endcase
end
always @(*) begin
	builder_rhs_array_muxed6 <= 1'd0;
	case (main_sdram_choose_req_grant)
		1'd0: begin
			builder_rhs_array_muxed6 <= main_sdram_choose_req_valids[0];
		end
		1'd1: begin
			builder_rhs_array_muxed6 <= main_sdram_choose_req_valids[1];
		end
		2'd2: begin
			builder_rhs_array_muxed6 <= main_sdram_choose_req_valids[2];
		end
		2'd3: begin
			builder_rhs_array_muxed6 <= main_sdram_choose_req_valids[3];
		end
		3'd4: begin
			builder_rhs_array_muxed6 <= main_sdram_choose_req_valids[4];
		end
		3'd5: begin
			builder_rhs_array_muxed6 <= main_sdram_choose_req_valids[5];
		end
		3'd6: begin
			builder_rhs_array_muxed6 <= main_sdram_choose_req_valids[6];
		end
		default: begin
			builder_rhs_array_muxed6 <= main_sdram_choose_req_valids[7];
		end
	endcase
end
always @(*) begin
	builder_rhs_array_muxed7 <= 14'd0;
	case (main_sdram_choose_req_grant)
		1'd0: begin
			builder_rhs_array_muxed7 <= main_sdram_bankmachine0_cmd_payload_a;
		end
		1'd1: begin
			builder_rhs_array_muxed7 <= main_sdram_bankmachine1_cmd_payload_a;
		end
		2'd2: begin
			builder_rhs_array_muxed7 <= main_sdram_bankmachine2_cmd_payload_a;
		end
		2'd3: begin
			builder_rhs_array_muxed7 <= main_sdram_bankmachine3_cmd_payload_a;
		end
		3'd4: begin
			builder_rhs_array_muxed7 <= main_sdram_bankmachine4_cmd_payload_a;
		end
		3'd5: begin
			builder_rhs_array_muxed7 <= main_sdram_bankmachine5_cmd_payload_a;
		end
		3'd6: begin
			builder_rhs_array_muxed7 <= main_sdram_bankmachine6_cmd_payload_a;
		end
		default: begin
			builder_rhs_array_muxed7 <= main_sdram_bankmachine7_cmd_payload_a;
		end
	endcase
end
always @(*) begin
	builder_rhs_array_muxed8 <= 3'd0;
	case (main_sdram_choose_req_grant)
		1'd0: begin
			builder_rhs_array_muxed8 <= main_sdram_bankmachine0_cmd_payload_ba;
		end
		1'd1: begin
			builder_rhs_array_muxed8 <= main_sdram_bankmachine1_cmd_payload_ba;
		end
		2'd2: begin
			builder_rhs_array_muxed8 <= main_sdram_bankmachine2_cmd_payload_ba;
		end
		2'd3: begin
			builder_rhs_array_muxed8 <= main_sdram_bankmachine3_cmd_payload_ba;
		end
		3'd4: begin
			builder_rhs_array_muxed8 <= main_sdram_bankmachine4_cmd_payload_ba;
		end
		3'd5: begin
			builder_rhs_array_muxed8 <= main_sdram_bankmachine5_cmd_payload_ba;
		end
		3'd6: begin
			builder_rhs_array_muxed8 <= main_sdram_bankmachine6_cmd_payload_ba;
		end
		default: begin
			builder_rhs_array_muxed8 <= main_sdram_bankmachine7_cmd_payload_ba;
		end
	endcase
end
always @(*) begin
	builder_rhs_array_muxed9 <= 1'd0;
	case (main_sdram_choose_req_grant)
		1'd0: begin
			builder_rhs_array_muxed9 <= main_sdram_bankmachine0_cmd_payload_is_read;
		end
		1'd1: begin
			builder_rhs_array_muxed9 <= main_sdram_bankmachine1_cmd_payload_is_read;
		end
		2'd2: begin
			builder_rhs_array_muxed9 <= main_sdram_bankmachine2_cmd_payload_is_read;
		end
		2'd3: begin
			builder_rhs_array_muxed9 <= main_sdram_bankmachine3_cmd_payload_is_read;
		end
		3'd4: begin
			builder_rhs_array_muxed9 <= main_sdram_bankmachine4_cmd_payload_is_read;
		end
		3'd5: begin
			builder_rhs_array_muxed9 <= main_sdram_bankmachine5_cmd_payload_is_read;
		end
		3'd6: begin
			builder_rhs_array_muxed9 <= main_sdram_bankmachine6_cmd_payload_is_read;
		end
		default: begin
			builder_rhs_array_muxed9 <= main_sdram_bankmachine7_cmd_payload_is_read;
		end
	endcase
end
always @(*) begin
	builder_rhs_array_muxed10 <= 1'd0;
	case (main_sdram_choose_req_grant)
		1'd0: begin
			builder_rhs_array_muxed10 <= main_sdram_bankmachine0_cmd_payload_is_write;
		end
		1'd1: begin
			builder_rhs_array_muxed10 <= main_sdram_bankmachine1_cmd_payload_is_write;
		end
		2'd2: begin
			builder_rhs_array_muxed10 <= main_sdram_bankmachine2_cmd_payload_is_write;
		end
		2'd3: begin
			builder_rhs_array_muxed10 <= main_sdram_bankmachine3_cmd_payload_is_write;
		end
		3'd4: begin
			builder_rhs_array_muxed10 <= main_sdram_bankmachine4_cmd_payload_is_write;
		end
		3'd5: begin
			builder_rhs_array_muxed10 <= main_sdram_bankmachine5_cmd_payload_is_write;
		end
		3'd6: begin
			builder_rhs_array_muxed10 <= main_sdram_bankmachine6_cmd_payload_is_write;
		end
		default: begin
			builder_rhs_array_muxed10 <= main_sdram_bankmachine7_cmd_payload_is_write;
		end
	endcase
end
always @(*) begin
	builder_rhs_array_muxed11 <= 1'd0;
	case (main_sdram_choose_req_grant)
		1'd0: begin
			builder_rhs_array_muxed11 <= main_sdram_bankmachine0_cmd_payload_is_cmd;
		end
		1'd1: begin
			builder_rhs_array_muxed11 <= main_sdram_bankmachine1_cmd_payload_is_cmd;
		end
		2'd2: begin
			builder_rhs_array_muxed11 <= main_sdram_bankmachine2_cmd_payload_is_cmd;
		end
		2'd3: begin
			builder_rhs_array_muxed11 <= main_sdram_bankmachine3_cmd_payload_is_cmd;
		end
		3'd4: begin
			builder_rhs_array_muxed11 <= main_sdram_bankmachine4_cmd_payload_is_cmd;
		end
		3'd5: begin
			builder_rhs_array_muxed11 <= main_sdram_bankmachine5_cmd_payload_is_cmd;
		end
		3'd6: begin
			builder_rhs_array_muxed11 <= main_sdram_bankmachine6_cmd_payload_is_cmd;
		end
		default: begin
			builder_rhs_array_muxed11 <= main_sdram_bankmachine7_cmd_payload_is_cmd;
		end
	endcase
end
always @(*) begin
	builder_t_array_muxed3 <= 1'd0;
	case (main_sdram_choose_req_grant)
		1'd0: begin
			builder_t_array_muxed3 <= main_sdram_bankmachine0_cmd_payload_cas;
		end
		1'd1: begin
			builder_t_array_muxed3 <= main_sdram_bankmachine1_cmd_payload_cas;
		end
		2'd2: begin
			builder_t_array_muxed3 <= main_sdram_bankmachine2_cmd_payload_cas;
		end
		2'd3: begin
			builder_t_array_muxed3 <= main_sdram_bankmachine3_cmd_payload_cas;
		end
		3'd4: begin
			builder_t_array_muxed3 <= main_sdram_bankmachine4_cmd_payload_cas;
		end
		3'd5: begin
			builder_t_array_muxed3 <= main_sdram_bankmachine5_cmd_payload_cas;
		end
		3'd6: begin
			builder_t_array_muxed3 <= main_sdram_bankmachine6_cmd_payload_cas;
		end
		default: begin
			builder_t_array_muxed3 <= main_sdram_bankmachine7_cmd_payload_cas;
		end
	endcase
end
always @(*) begin
	builder_t_array_muxed4 <= 1'd0;
	case (main_sdram_choose_req_grant)
		1'd0: begin
			builder_t_array_muxed4 <= main_sdram_bankmachine0_cmd_payload_ras;
		end
		1'd1: begin
			builder_t_array_muxed4 <= main_sdram_bankmachine1_cmd_payload_ras;
		end
		2'd2: begin
			builder_t_array_muxed4 <= main_sdram_bankmachine2_cmd_payload_ras;
		end
		2'd3: begin
			builder_t_array_muxed4 <= main_sdram_bankmachine3_cmd_payload_ras;
		end
		3'd4: begin
			builder_t_array_muxed4 <= main_sdram_bankmachine4_cmd_payload_ras;
		end
		3'd5: begin
			builder_t_array_muxed4 <= main_sdram_bankmachine5_cmd_payload_ras;
		end
		3'd6: begin
			builder_t_array_muxed4 <= main_sdram_bankmachine6_cmd_payload_ras;
		end
		default: begin
			builder_t_array_muxed4 <= main_sdram_bankmachine7_cmd_payload_ras;
		end
	endcase
end
always @(*) begin
	builder_t_array_muxed5 <= 1'd0;
	case (main_sdram_choose_req_grant)
		1'd0: begin
			builder_t_array_muxed5 <= main_sdram_bankmachine0_cmd_payload_we;
		end
		1'd1: begin
			builder_t_array_muxed5 <= main_sdram_bankmachine1_cmd_payload_we;
		end
		2'd2: begin
			builder_t_array_muxed5 <= main_sdram_bankmachine2_cmd_payload_we;
		end
		2'd3: begin
			builder_t_array_muxed5 <= main_sdram_bankmachine3_cmd_payload_we;
		end
		3'd4: begin
			builder_t_array_muxed5 <= main_sdram_bankmachine4_cmd_payload_we;
		end
		3'd5: begin
			builder_t_array_muxed5 <= main_sdram_bankmachine5_cmd_payload_we;
		end
		3'd6: begin
			builder_t_array_muxed5 <= main_sdram_bankmachine6_cmd_payload_we;
		end
		default: begin
			builder_t_array_muxed5 <= main_sdram_bankmachine7_cmd_payload_we;
		end
	endcase
end
always @(*) begin
	builder_rhs_array_muxed12 <= 21'd0;
	case (builder_roundrobin0_grant)
		default: begin
			builder_rhs_array_muxed12 <= {main_port_cmd_payload_addr[23:10], main_port_cmd_payload_addr[6:0]};
		end
	endcase
end
always @(*) begin
	builder_rhs_array_muxed13 <= 1'd0;
	case (builder_roundrobin0_grant)
		default: begin
			builder_rhs_array_muxed13 <= main_port_cmd_payload_we;
		end
	endcase
end
always @(*) begin
	builder_rhs_array_muxed14 <= 1'd0;
	case (builder_roundrobin0_grant)
		default: begin
			builder_rhs_array_muxed14 <= (((main_port_cmd_payload_addr[9:7] == 1'd0) & (~(((((((builder_locked0 | (main_sdram_interface_bank1_lock & (builder_roundrobin1_grant == 1'd0))) | (main_sdram_interface_bank2_lock & (builder_roundrobin2_grant == 1'd0))) | (main_sdram_interface_bank3_lock & (builder_roundrobin3_grant == 1'd0))) | (main_sdram_interface_bank4_lock & (builder_roundrobin4_grant == 1'd0))) | (main_sdram_interface_bank5_lock & (builder_roundrobin5_grant == 1'd0))) | (main_sdram_interface_bank6_lock & (builder_roundrobin6_grant == 1'd0))) | (main_sdram_interface_bank7_lock & (builder_roundrobin7_grant == 1'd0))))) & main_port_cmd_valid);
		end
	endcase
end
always @(*) begin
	builder_rhs_array_muxed15 <= 21'd0;
	case (builder_roundrobin1_grant)
		default: begin
			builder_rhs_array_muxed15 <= {main_port_cmd_payload_addr[23:10], main_port_cmd_payload_addr[6:0]};
		end
	endcase
end
always @(*) begin
	builder_rhs_array_muxed16 <= 1'd0;
	case (builder_roundrobin1_grant)
		default: begin
			builder_rhs_array_muxed16 <= main_port_cmd_payload_we;
		end
	endcase
end
always @(*) begin
	builder_rhs_array_muxed17 <= 1'd0;
	case (builder_roundrobin1_grant)
		default: begin
			builder_rhs_array_muxed17 <= (((main_port_cmd_payload_addr[9:7] == 1'd1) & (~(((((((builder_locked1 | (main_sdram_interface_bank0_lock & (builder_roundrobin0_grant == 1'd0))) | (main_sdram_interface_bank2_lock & (builder_roundrobin2_grant == 1'd0))) | (main_sdram_interface_bank3_lock & (builder_roundrobin3_grant == 1'd0))) | (main_sdram_interface_bank4_lock & (builder_roundrobin4_grant == 1'd0))) | (main_sdram_interface_bank5_lock & (builder_roundrobin5_grant == 1'd0))) | (main_sdram_interface_bank6_lock & (builder_roundrobin6_grant == 1'd0))) | (main_sdram_interface_bank7_lock & (builder_roundrobin7_grant == 1'd0))))) & main_port_cmd_valid);
		end
	endcase
end
always @(*) begin
	builder_rhs_array_muxed18 <= 21'd0;
	case (builder_roundrobin2_grant)
		default: begin
			builder_rhs_array_muxed18 <= {main_port_cmd_payload_addr[23:10], main_port_cmd_payload_addr[6:0]};
		end
	endcase
end
always @(*) begin
	builder_rhs_array_muxed19 <= 1'd0;
	case (builder_roundrobin2_grant)
		default: begin
			builder_rhs_array_muxed19 <= main_port_cmd_payload_we;
		end
	endcase
end
always @(*) begin
	builder_rhs_array_muxed20 <= 1'd0;
	case (builder_roundrobin2_grant)
		default: begin
			builder_rhs_array_muxed20 <= (((main_port_cmd_payload_addr[9:7] == 2'd2) & (~(((((((builder_locked2 | (main_sdram_interface_bank0_lock & (builder_roundrobin0_grant == 1'd0))) | (main_sdram_interface_bank1_lock & (builder_roundrobin1_grant == 1'd0))) | (main_sdram_interface_bank3_lock & (builder_roundrobin3_grant == 1'd0))) | (main_sdram_interface_bank4_lock & (builder_roundrobin4_grant == 1'd0))) | (main_sdram_interface_bank5_lock & (builder_roundrobin5_grant == 1'd0))) | (main_sdram_interface_bank6_lock & (builder_roundrobin6_grant == 1'd0))) | (main_sdram_interface_bank7_lock & (builder_roundrobin7_grant == 1'd0))))) & main_port_cmd_valid);
		end
	endcase
end
always @(*) begin
	builder_rhs_array_muxed21 <= 21'd0;
	case (builder_roundrobin3_grant)
		default: begin
			builder_rhs_array_muxed21 <= {main_port_cmd_payload_addr[23:10], main_port_cmd_payload_addr[6:0]};
		end
	endcase
end
always @(*) begin
	builder_rhs_array_muxed22 <= 1'd0;
	case (builder_roundrobin3_grant)
		default: begin
			builder_rhs_array_muxed22 <= main_port_cmd_payload_we;
		end
	endcase
end
always @(*) begin
	builder_rhs_array_muxed23 <= 1'd0;
	case (builder_roundrobin3_grant)
		default: begin
			builder_rhs_array_muxed23 <= (((main_port_cmd_payload_addr[9:7] == 2'd3) & (~(((((((builder_locked3 | (main_sdram_interface_bank0_lock & (builder_roundrobin0_grant == 1'd0))) | (main_sdram_interface_bank1_lock & (builder_roundrobin1_grant == 1'd0))) | (main_sdram_interface_bank2_lock & (builder_roundrobin2_grant == 1'd0))) | (main_sdram_interface_bank4_lock & (builder_roundrobin4_grant == 1'd0))) | (main_sdram_interface_bank5_lock & (builder_roundrobin5_grant == 1'd0))) | (main_sdram_interface_bank6_lock & (builder_roundrobin6_grant == 1'd0))) | (main_sdram_interface_bank7_lock & (builder_roundrobin7_grant == 1'd0))))) & main_port_cmd_valid);
		end
	endcase
end
always @(*) begin
	builder_rhs_array_muxed24 <= 21'd0;
	case (builder_roundrobin4_grant)
		default: begin
			builder_rhs_array_muxed24 <= {main_port_cmd_payload_addr[23:10], main_port_cmd_payload_addr[6:0]};
		end
	endcase
end
always @(*) begin
	builder_rhs_array_muxed25 <= 1'd0;
	case (builder_roundrobin4_grant)
		default: begin
			builder_rhs_array_muxed25 <= main_port_cmd_payload_we;
		end
	endcase
end
always @(*) begin
	builder_rhs_array_muxed26 <= 1'd0;
	case (builder_roundrobin4_grant)
		default: begin
			builder_rhs_array_muxed26 <= (((main_port_cmd_payload_addr[9:7] == 3'd4) & (~(((((((builder_locked4 | (main_sdram_interface_bank0_lock & (builder_roundrobin0_grant == 1'd0))) | (main_sdram_interface_bank1_lock & (builder_roundrobin1_grant == 1'd0))) | (main_sdram_interface_bank2_lock & (builder_roundrobin2_grant == 1'd0))) | (main_sdram_interface_bank3_lock & (builder_roundrobin3_grant == 1'd0))) | (main_sdram_interface_bank5_lock & (builder_roundrobin5_grant == 1'd0))) | (main_sdram_interface_bank6_lock & (builder_roundrobin6_grant == 1'd0))) | (main_sdram_interface_bank7_lock & (builder_roundrobin7_grant == 1'd0))))) & main_port_cmd_valid);
		end
	endcase
end
always @(*) begin
	builder_rhs_array_muxed27 <= 21'd0;
	case (builder_roundrobin5_grant)
		default: begin
			builder_rhs_array_muxed27 <= {main_port_cmd_payload_addr[23:10], main_port_cmd_payload_addr[6:0]};
		end
	endcase
end
always @(*) begin
	builder_rhs_array_muxed28 <= 1'd0;
	case (builder_roundrobin5_grant)
		default: begin
			builder_rhs_array_muxed28 <= main_port_cmd_payload_we;
		end
	endcase
end
always @(*) begin
	builder_rhs_array_muxed29 <= 1'd0;
	case (builder_roundrobin5_grant)
		default: begin
			builder_rhs_array_muxed29 <= (((main_port_cmd_payload_addr[9:7] == 3'd5) & (~(((((((builder_locked5 | (main_sdram_interface_bank0_lock & (builder_roundrobin0_grant == 1'd0))) | (main_sdram_interface_bank1_lock & (builder_roundrobin1_grant == 1'd0))) | (main_sdram_interface_bank2_lock & (builder_roundrobin2_grant == 1'd0))) | (main_sdram_interface_bank3_lock & (builder_roundrobin3_grant == 1'd0))) | (main_sdram_interface_bank4_lock & (builder_roundrobin4_grant == 1'd0))) | (main_sdram_interface_bank6_lock & (builder_roundrobin6_grant == 1'd0))) | (main_sdram_interface_bank7_lock & (builder_roundrobin7_grant == 1'd0))))) & main_port_cmd_valid);
		end
	endcase
end
always @(*) begin
	builder_rhs_array_muxed30 <= 21'd0;
	case (builder_roundrobin6_grant)
		default: begin
			builder_rhs_array_muxed30 <= {main_port_cmd_payload_addr[23:10], main_port_cmd_payload_addr[6:0]};
		end
	endcase
end
always @(*) begin
	builder_rhs_array_muxed31 <= 1'd0;
	case (builder_roundrobin6_grant)
		default: begin
			builder_rhs_array_muxed31 <= main_port_cmd_payload_we;
		end
	endcase
end
always @(*) begin
	builder_rhs_array_muxed32 <= 1'd0;
	case (builder_roundrobin6_grant)
		default: begin
			builder_rhs_array_muxed32 <= (((main_port_cmd_payload_addr[9:7] == 3'd6) & (~(((((((builder_locked6 | (main_sdram_interface_bank0_lock & (builder_roundrobin0_grant == 1'd0))) | (main_sdram_interface_bank1_lock & (builder_roundrobin1_grant == 1'd0))) | (main_sdram_interface_bank2_lock & (builder_roundrobin2_grant == 1'd0))) | (main_sdram_interface_bank3_lock & (builder_roundrobin3_grant == 1'd0))) | (main_sdram_interface_bank4_lock & (builder_roundrobin4_grant == 1'd0))) | (main_sdram_interface_bank5_lock & (builder_roundrobin5_grant == 1'd0))) | (main_sdram_interface_bank7_lock & (builder_roundrobin7_grant == 1'd0))))) & main_port_cmd_valid);
		end
	endcase
end
always @(*) begin
	builder_rhs_array_muxed33 <= 21'd0;
	case (builder_roundrobin7_grant)
		default: begin
			builder_rhs_array_muxed33 <= {main_port_cmd_payload_addr[23:10], main_port_cmd_payload_addr[6:0]};
		end
	endcase
end
always @(*) begin
	builder_rhs_array_muxed34 <= 1'd0;
	case (builder_roundrobin7_grant)
		default: begin
			builder_rhs_array_muxed34 <= main_port_cmd_payload_we;
		end
	endcase
end
always @(*) begin
	builder_rhs_array_muxed35 <= 1'd0;
	case (builder_roundrobin7_grant)
		default: begin
			builder_rhs_array_muxed35 <= (((main_port_cmd_payload_addr[9:7] == 3'd7) & (~(((((((builder_locked7 | (main_sdram_interface_bank0_lock & (builder_roundrobin0_grant == 1'd0))) | (main_sdram_interface_bank1_lock & (builder_roundrobin1_grant == 1'd0))) | (main_sdram_interface_bank2_lock & (builder_roundrobin2_grant == 1'd0))) | (main_sdram_interface_bank3_lock & (builder_roundrobin3_grant == 1'd0))) | (main_sdram_interface_bank4_lock & (builder_roundrobin4_grant == 1'd0))) | (main_sdram_interface_bank5_lock & (builder_roundrobin5_grant == 1'd0))) | (main_sdram_interface_bank6_lock & (builder_roundrobin6_grant == 1'd0))))) & main_port_cmd_valid);
		end
	endcase
end
always @(*) begin
	builder_rhs_array_muxed36 <= 30'd0;
	case (builder_wb_sdram_con_grant)
		default: begin
			builder_rhs_array_muxed36 <= main_interface1_wb_sdram_adr;
		end
	endcase
end
always @(*) begin
	builder_rhs_array_muxed37 <= 32'd0;
	case (builder_wb_sdram_con_grant)
		default: begin
			builder_rhs_array_muxed37 <= main_interface1_wb_sdram_dat_w;
		end
	endcase
end
always @(*) begin
	builder_rhs_array_muxed38 <= 4'd0;
	case (builder_wb_sdram_con_grant)
		default: begin
			builder_rhs_array_muxed38 <= main_interface1_wb_sdram_sel;
		end
	endcase
end
always @(*) begin
	builder_rhs_array_muxed39 <= 1'd0;
	case (builder_wb_sdram_con_grant)
		default: begin
			builder_rhs_array_muxed39 <= main_interface1_wb_sdram_cyc;
		end
	endcase
end
always @(*) begin
	builder_rhs_array_muxed40 <= 1'd0;
	case (builder_wb_sdram_con_grant)
		default: begin
			builder_rhs_array_muxed40 <= main_interface1_wb_sdram_stb;
		end
	endcase
end
always @(*) begin
	builder_rhs_array_muxed41 <= 1'd0;
	case (builder_wb_sdram_con_grant)
		default: begin
			builder_rhs_array_muxed41 <= main_interface1_wb_sdram_we;
		end
	endcase
end
always @(*) begin
	builder_rhs_array_muxed42 <= 3'd0;
	case (builder_wb_sdram_con_grant)
		default: begin
			builder_rhs_array_muxed42 <= main_interface1_wb_sdram_cti;
		end
	endcase
end
always @(*) begin
	builder_rhs_array_muxed43 <= 2'd0;
	case (builder_wb_sdram_con_grant)
		default: begin
			builder_rhs_array_muxed43 <= main_interface1_wb_sdram_bte;
		end
	endcase
end
always @(*) begin
	builder_rhs_array_muxed44 <= 30'd0;
	case (builder_basesoc_grant)
		default: begin
			builder_rhs_array_muxed44 <= main_uart_wishbone_adr;
		end
	endcase
end
always @(*) begin
	builder_rhs_array_muxed45 <= 32'd0;
	case (builder_basesoc_grant)
		default: begin
			builder_rhs_array_muxed45 <= main_uart_wishbone_dat_w;
		end
	endcase
end
always @(*) begin
	builder_rhs_array_muxed46 <= 4'd0;
	case (builder_basesoc_grant)
		default: begin
			builder_rhs_array_muxed46 <= main_uart_wishbone_sel;
		end
	endcase
end
always @(*) begin
	builder_rhs_array_muxed47 <= 1'd0;
	case (builder_basesoc_grant)
		default: begin
			builder_rhs_array_muxed47 <= main_uart_wishbone_cyc;
		end
	endcase
end
always @(*) begin
	builder_rhs_array_muxed48 <= 1'd0;
	case (builder_basesoc_grant)
		default: begin
			builder_rhs_array_muxed48 <= main_uart_wishbone_stb;
		end
	endcase
end
always @(*) begin
	builder_rhs_array_muxed49 <= 1'd0;
	case (builder_basesoc_grant)
		default: begin
			builder_rhs_array_muxed49 <= main_uart_wishbone_we;
		end
	endcase
end
always @(*) begin
	builder_rhs_array_muxed50 <= 3'd0;
	case (builder_basesoc_grant)
		default: begin
			builder_rhs_array_muxed50 <= main_uart_wishbone_cti;
		end
	endcase
end
always @(*) begin
	builder_rhs_array_muxed51 <= 2'd0;
	case (builder_basesoc_grant)
		default: begin
			builder_rhs_array_muxed51 <= main_uart_wishbone_bte;
		end
	endcase
end
always @(*) begin
	builder_array_muxed0 <= 3'd0;
	case (main_sdram_steerer_sel0)
		1'd0: begin
			builder_array_muxed0 <= main_sdram_nop_ba[2:0];
		end
		1'd1: begin
			builder_array_muxed0 <= main_sdram_choose_cmd_cmd_payload_ba[2:0];
		end
		2'd2: begin
			builder_array_muxed0 <= main_sdram_choose_req_cmd_payload_ba[2:0];
		end
		default: begin
			builder_array_muxed0 <= main_sdram_cmd_payload_ba[2:0];
		end
	endcase
end
always @(*) begin
	builder_array_muxed1 <= 14'd0;
	case (main_sdram_steerer_sel0)
		1'd0: begin
			builder_array_muxed1 <= main_sdram_nop_a;
		end
		1'd1: begin
			builder_array_muxed1 <= main_sdram_choose_cmd_cmd_payload_a;
		end
		2'd2: begin
			builder_array_muxed1 <= main_sdram_choose_req_cmd_payload_a;
		end
		default: begin
			builder_array_muxed1 <= main_sdram_cmd_payload_a;
		end
	endcase
end
always @(*) begin
	builder_array_muxed2 <= 1'd0;
	case (main_sdram_steerer_sel0)
		1'd0: begin
			builder_array_muxed2 <= 1'd0;
		end
		1'd1: begin
			builder_array_muxed2 <= ((main_sdram_choose_cmd_cmd_valid & main_sdram_choose_cmd_cmd_ready) & main_sdram_choose_cmd_cmd_payload_cas);
		end
		2'd2: begin
			builder_array_muxed2 <= ((main_sdram_choose_req_cmd_valid & main_sdram_choose_req_cmd_ready) & main_sdram_choose_req_cmd_payload_cas);
		end
		default: begin
			builder_array_muxed2 <= ((main_sdram_cmd_valid & main_sdram_cmd_ready) & main_sdram_cmd_payload_cas);
		end
	endcase
end
always @(*) begin
	builder_array_muxed3 <= 1'd0;
	case (main_sdram_steerer_sel0)
		1'd0: begin
			builder_array_muxed3 <= 1'd0;
		end
		1'd1: begin
			builder_array_muxed3 <= ((main_sdram_choose_cmd_cmd_valid & main_sdram_choose_cmd_cmd_ready) & main_sdram_choose_cmd_cmd_payload_ras);
		end
		2'd2: begin
			builder_array_muxed3 <= ((main_sdram_choose_req_cmd_valid & main_sdram_choose_req_cmd_ready) & main_sdram_choose_req_cmd_payload_ras);
		end
		default: begin
			builder_array_muxed3 <= ((main_sdram_cmd_valid & main_sdram_cmd_ready) & main_sdram_cmd_payload_ras);
		end
	endcase
end
always @(*) begin
	builder_array_muxed4 <= 1'd0;
	case (main_sdram_steerer_sel0)
		1'd0: begin
			builder_array_muxed4 <= 1'd0;
		end
		1'd1: begin
			builder_array_muxed4 <= ((main_sdram_choose_cmd_cmd_valid & main_sdram_choose_cmd_cmd_ready) & main_sdram_choose_cmd_cmd_payload_we);
		end
		2'd2: begin
			builder_array_muxed4 <= ((main_sdram_choose_req_cmd_valid & main_sdram_choose_req_cmd_ready) & main_sdram_choose_req_cmd_payload_we);
		end
		default: begin
			builder_array_muxed4 <= ((main_sdram_cmd_valid & main_sdram_cmd_ready) & main_sdram_cmd_payload_we);
		end
	endcase
end
always @(*) begin
	builder_array_muxed5 <= 1'd0;
	case (main_sdram_steerer_sel0)
		1'd0: begin
			builder_array_muxed5 <= 1'd0;
		end
		1'd1: begin
			builder_array_muxed5 <= ((main_sdram_choose_cmd_cmd_valid & main_sdram_choose_cmd_cmd_ready) & main_sdram_choose_cmd_cmd_payload_is_read);
		end
		2'd2: begin
			builder_array_muxed5 <= ((main_sdram_choose_req_cmd_valid & main_sdram_choose_req_cmd_ready) & main_sdram_choose_req_cmd_payload_is_read);
		end
		default: begin
			builder_array_muxed5 <= ((main_sdram_cmd_valid & main_sdram_cmd_ready) & main_sdram_cmd_payload_is_read);
		end
	endcase
end
always @(*) begin
	builder_array_muxed6 <= 1'd0;
	case (main_sdram_steerer_sel0)
		1'd0: begin
			builder_array_muxed6 <= 1'd0;
		end
		1'd1: begin
			builder_array_muxed6 <= ((main_sdram_choose_cmd_cmd_valid & main_sdram_choose_cmd_cmd_ready) & main_sdram_choose_cmd_cmd_payload_is_write);
		end
		2'd2: begin
			builder_array_muxed6 <= ((main_sdram_choose_req_cmd_valid & main_sdram_choose_req_cmd_ready) & main_sdram_choose_req_cmd_payload_is_write);
		end
		default: begin
			builder_array_muxed6 <= ((main_sdram_cmd_valid & main_sdram_cmd_ready) & main_sdram_cmd_payload_is_write);
		end
	endcase
end
always @(*) begin
	builder_array_muxed7 <= 3'd0;
	case (main_sdram_steerer_sel1)
		1'd0: begin
			builder_array_muxed7 <= main_sdram_nop_ba[2:0];
		end
		1'd1: begin
			builder_array_muxed7 <= main_sdram_choose_cmd_cmd_payload_ba[2:0];
		end
		2'd2: begin
			builder_array_muxed7 <= main_sdram_choose_req_cmd_payload_ba[2:0];
		end
		default: begin
			builder_array_muxed7 <= main_sdram_cmd_payload_ba[2:0];
		end
	endcase
end
always @(*) begin
	builder_array_muxed8 <= 14'd0;
	case (main_sdram_steerer_sel1)
		1'd0: begin
			builder_array_muxed8 <= main_sdram_nop_a;
		end
		1'd1: begin
			builder_array_muxed8 <= main_sdram_choose_cmd_cmd_payload_a;
		end
		2'd2: begin
			builder_array_muxed8 <= main_sdram_choose_req_cmd_payload_a;
		end
		default: begin
			builder_array_muxed8 <= main_sdram_cmd_payload_a;
		end
	endcase
end
always @(*) begin
	builder_array_muxed9 <= 1'd0;
	case (main_sdram_steerer_sel1)
		1'd0: begin
			builder_array_muxed9 <= 1'd0;
		end
		1'd1: begin
			builder_array_muxed9 <= ((main_sdram_choose_cmd_cmd_valid & main_sdram_choose_cmd_cmd_ready) & main_sdram_choose_cmd_cmd_payload_cas);
		end
		2'd2: begin
			builder_array_muxed9 <= ((main_sdram_choose_req_cmd_valid & main_sdram_choose_req_cmd_ready) & main_sdram_choose_req_cmd_payload_cas);
		end
		default: begin
			builder_array_muxed9 <= ((main_sdram_cmd_valid & main_sdram_cmd_ready) & main_sdram_cmd_payload_cas);
		end
	endcase
end
always @(*) begin
	builder_array_muxed10 <= 1'd0;
	case (main_sdram_steerer_sel1)
		1'd0: begin
			builder_array_muxed10 <= 1'd0;
		end
		1'd1: begin
			builder_array_muxed10 <= ((main_sdram_choose_cmd_cmd_valid & main_sdram_choose_cmd_cmd_ready) & main_sdram_choose_cmd_cmd_payload_ras);
		end
		2'd2: begin
			builder_array_muxed10 <= ((main_sdram_choose_req_cmd_valid & main_sdram_choose_req_cmd_ready) & main_sdram_choose_req_cmd_payload_ras);
		end
		default: begin
			builder_array_muxed10 <= ((main_sdram_cmd_valid & main_sdram_cmd_ready) & main_sdram_cmd_payload_ras);
		end
	endcase
end
always @(*) begin
	builder_array_muxed11 <= 1'd0;
	case (main_sdram_steerer_sel1)
		1'd0: begin
			builder_array_muxed11 <= 1'd0;
		end
		1'd1: begin
			builder_array_muxed11 <= ((main_sdram_choose_cmd_cmd_valid & main_sdram_choose_cmd_cmd_ready) & main_sdram_choose_cmd_cmd_payload_we);
		end
		2'd2: begin
			builder_array_muxed11 <= ((main_sdram_choose_req_cmd_valid & main_sdram_choose_req_cmd_ready) & main_sdram_choose_req_cmd_payload_we);
		end
		default: begin
			builder_array_muxed11 <= ((main_sdram_cmd_valid & main_sdram_cmd_ready) & main_sdram_cmd_payload_we);
		end
	endcase
end
always @(*) begin
	builder_array_muxed12 <= 1'd0;
	case (main_sdram_steerer_sel1)
		1'd0: begin
			builder_array_muxed12 <= 1'd0;
		end
		1'd1: begin
			builder_array_muxed12 <= ((main_sdram_choose_cmd_cmd_valid & main_sdram_choose_cmd_cmd_ready) & main_sdram_choose_cmd_cmd_payload_is_read);
		end
		2'd2: begin
			builder_array_muxed12 <= ((main_sdram_choose_req_cmd_valid & main_sdram_choose_req_cmd_ready) & main_sdram_choose_req_cmd_payload_is_read);
		end
		default: begin
			builder_array_muxed12 <= ((main_sdram_cmd_valid & main_sdram_cmd_ready) & main_sdram_cmd_payload_is_read);
		end
	endcase
end
always @(*) begin
	builder_array_muxed13 <= 1'd0;
	case (main_sdram_steerer_sel1)
		1'd0: begin
			builder_array_muxed13 <= 1'd0;
		end
		1'd1: begin
			builder_array_muxed13 <= ((main_sdram_choose_cmd_cmd_valid & main_sdram_choose_cmd_cmd_ready) & main_sdram_choose_cmd_cmd_payload_is_write);
		end
		2'd2: begin
			builder_array_muxed13 <= ((main_sdram_choose_req_cmd_valid & main_sdram_choose_req_cmd_ready) & main_sdram_choose_req_cmd_payload_is_write);
		end
		default: begin
			builder_array_muxed13 <= ((main_sdram_cmd_valid & main_sdram_cmd_ready) & main_sdram_cmd_payload_is_write);
		end
	endcase
end
always @(*) begin
	builder_array_muxed14 <= 3'd0;
	case (main_sdram_steerer_sel2)
		1'd0: begin
			builder_array_muxed14 <= main_sdram_nop_ba[2:0];
		end
		1'd1: begin
			builder_array_muxed14 <= main_sdram_choose_cmd_cmd_payload_ba[2:0];
		end
		2'd2: begin
			builder_array_muxed14 <= main_sdram_choose_req_cmd_payload_ba[2:0];
		end
		default: begin
			builder_array_muxed14 <= main_sdram_cmd_payload_ba[2:0];
		end
	endcase
end
always @(*) begin
	builder_array_muxed15 <= 14'd0;
	case (main_sdram_steerer_sel2)
		1'd0: begin
			builder_array_muxed15 <= main_sdram_nop_a;
		end
		1'd1: begin
			builder_array_muxed15 <= main_sdram_choose_cmd_cmd_payload_a;
		end
		2'd2: begin
			builder_array_muxed15 <= main_sdram_choose_req_cmd_payload_a;
		end
		default: begin
			builder_array_muxed15 <= main_sdram_cmd_payload_a;
		end
	endcase
end
always @(*) begin
	builder_array_muxed16 <= 1'd0;
	case (main_sdram_steerer_sel2)
		1'd0: begin
			builder_array_muxed16 <= 1'd0;
		end
		1'd1: begin
			builder_array_muxed16 <= ((main_sdram_choose_cmd_cmd_valid & main_sdram_choose_cmd_cmd_ready) & main_sdram_choose_cmd_cmd_payload_cas);
		end
		2'd2: begin
			builder_array_muxed16 <= ((main_sdram_choose_req_cmd_valid & main_sdram_choose_req_cmd_ready) & main_sdram_choose_req_cmd_payload_cas);
		end
		default: begin
			builder_array_muxed16 <= ((main_sdram_cmd_valid & main_sdram_cmd_ready) & main_sdram_cmd_payload_cas);
		end
	endcase
end
always @(*) begin
	builder_array_muxed17 <= 1'd0;
	case (main_sdram_steerer_sel2)
		1'd0: begin
			builder_array_muxed17 <= 1'd0;
		end
		1'd1: begin
			builder_array_muxed17 <= ((main_sdram_choose_cmd_cmd_valid & main_sdram_choose_cmd_cmd_ready) & main_sdram_choose_cmd_cmd_payload_ras);
		end
		2'd2: begin
			builder_array_muxed17 <= ((main_sdram_choose_req_cmd_valid & main_sdram_choose_req_cmd_ready) & main_sdram_choose_req_cmd_payload_ras);
		end
		default: begin
			builder_array_muxed17 <= ((main_sdram_cmd_valid & main_sdram_cmd_ready) & main_sdram_cmd_payload_ras);
		end
	endcase
end
always @(*) begin
	builder_array_muxed18 <= 1'd0;
	case (main_sdram_steerer_sel2)
		1'd0: begin
			builder_array_muxed18 <= 1'd0;
		end
		1'd1: begin
			builder_array_muxed18 <= ((main_sdram_choose_cmd_cmd_valid & main_sdram_choose_cmd_cmd_ready) & main_sdram_choose_cmd_cmd_payload_we);
		end
		2'd2: begin
			builder_array_muxed18 <= ((main_sdram_choose_req_cmd_valid & main_sdram_choose_req_cmd_ready) & main_sdram_choose_req_cmd_payload_we);
		end
		default: begin
			builder_array_muxed18 <= ((main_sdram_cmd_valid & main_sdram_cmd_ready) & main_sdram_cmd_payload_we);
		end
	endcase
end
always @(*) begin
	builder_array_muxed19 <= 1'd0;
	case (main_sdram_steerer_sel2)
		1'd0: begin
			builder_array_muxed19 <= 1'd0;
		end
		1'd1: begin
			builder_array_muxed19 <= ((main_sdram_choose_cmd_cmd_valid & main_sdram_choose_cmd_cmd_ready) & main_sdram_choose_cmd_cmd_payload_is_read);
		end
		2'd2: begin
			builder_array_muxed19 <= ((main_sdram_choose_req_cmd_valid & main_sdram_choose_req_cmd_ready) & main_sdram_choose_req_cmd_payload_is_read);
		end
		default: begin
			builder_array_muxed19 <= ((main_sdram_cmd_valid & main_sdram_cmd_ready) & main_sdram_cmd_payload_is_read);
		end
	endcase
end
always @(*) begin
	builder_array_muxed20 <= 1'd0;
	case (main_sdram_steerer_sel2)
		1'd0: begin
			builder_array_muxed20 <= 1'd0;
		end
		1'd1: begin
			builder_array_muxed20 <= ((main_sdram_choose_cmd_cmd_valid & main_sdram_choose_cmd_cmd_ready) & main_sdram_choose_cmd_cmd_payload_is_write);
		end
		2'd2: begin
			builder_array_muxed20 <= ((main_sdram_choose_req_cmd_valid & main_sdram_choose_req_cmd_ready) & main_sdram_choose_req_cmd_payload_is_write);
		end
		default: begin
			builder_array_muxed20 <= ((main_sdram_cmd_valid & main_sdram_cmd_ready) & main_sdram_cmd_payload_is_write);
		end
	endcase
end
always @(*) begin
	builder_array_muxed21 <= 3'd0;
	case (main_sdram_steerer_sel3)
		1'd0: begin
			builder_array_muxed21 <= main_sdram_nop_ba[2:0];
		end
		1'd1: begin
			builder_array_muxed21 <= main_sdram_choose_cmd_cmd_payload_ba[2:0];
		end
		2'd2: begin
			builder_array_muxed21 <= main_sdram_choose_req_cmd_payload_ba[2:0];
		end
		default: begin
			builder_array_muxed21 <= main_sdram_cmd_payload_ba[2:0];
		end
	endcase
end
always @(*) begin
	builder_array_muxed22 <= 14'd0;
	case (main_sdram_steerer_sel3)
		1'd0: begin
			builder_array_muxed22 <= main_sdram_nop_a;
		end
		1'd1: begin
			builder_array_muxed22 <= main_sdram_choose_cmd_cmd_payload_a;
		end
		2'd2: begin
			builder_array_muxed22 <= main_sdram_choose_req_cmd_payload_a;
		end
		default: begin
			builder_array_muxed22 <= main_sdram_cmd_payload_a;
		end
	endcase
end
always @(*) begin
	builder_array_muxed23 <= 1'd0;
	case (main_sdram_steerer_sel3)
		1'd0: begin
			builder_array_muxed23 <= 1'd0;
		end
		1'd1: begin
			builder_array_muxed23 <= ((main_sdram_choose_cmd_cmd_valid & main_sdram_choose_cmd_cmd_ready) & main_sdram_choose_cmd_cmd_payload_cas);
		end
		2'd2: begin
			builder_array_muxed23 <= ((main_sdram_choose_req_cmd_valid & main_sdram_choose_req_cmd_ready) & main_sdram_choose_req_cmd_payload_cas);
		end
		default: begin
			builder_array_muxed23 <= ((main_sdram_cmd_valid & main_sdram_cmd_ready) & main_sdram_cmd_payload_cas);
		end
	endcase
end
always @(*) begin
	builder_array_muxed24 <= 1'd0;
	case (main_sdram_steerer_sel3)
		1'd0: begin
			builder_array_muxed24 <= 1'd0;
		end
		1'd1: begin
			builder_array_muxed24 <= ((main_sdram_choose_cmd_cmd_valid & main_sdram_choose_cmd_cmd_ready) & main_sdram_choose_cmd_cmd_payload_ras);
		end
		2'd2: begin
			builder_array_muxed24 <= ((main_sdram_choose_req_cmd_valid & main_sdram_choose_req_cmd_ready) & main_sdram_choose_req_cmd_payload_ras);
		end
		default: begin
			builder_array_muxed24 <= ((main_sdram_cmd_valid & main_sdram_cmd_ready) & main_sdram_cmd_payload_ras);
		end
	endcase
end
always @(*) begin
	builder_array_muxed25 <= 1'd0;
	case (main_sdram_steerer_sel3)
		1'd0: begin
			builder_array_muxed25 <= 1'd0;
		end
		1'd1: begin
			builder_array_muxed25 <= ((main_sdram_choose_cmd_cmd_valid & main_sdram_choose_cmd_cmd_ready) & main_sdram_choose_cmd_cmd_payload_we);
		end
		2'd2: begin
			builder_array_muxed25 <= ((main_sdram_choose_req_cmd_valid & main_sdram_choose_req_cmd_ready) & main_sdram_choose_req_cmd_payload_we);
		end
		default: begin
			builder_array_muxed25 <= ((main_sdram_cmd_valid & main_sdram_cmd_ready) & main_sdram_cmd_payload_we);
		end
	endcase
end
always @(*) begin
	builder_array_muxed26 <= 1'd0;
	case (main_sdram_steerer_sel3)
		1'd0: begin
			builder_array_muxed26 <= 1'd0;
		end
		1'd1: begin
			builder_array_muxed26 <= ((main_sdram_choose_cmd_cmd_valid & main_sdram_choose_cmd_cmd_ready) & main_sdram_choose_cmd_cmd_payload_is_read);
		end
		2'd2: begin
			builder_array_muxed26 <= ((main_sdram_choose_req_cmd_valid & main_sdram_choose_req_cmd_ready) & main_sdram_choose_req_cmd_payload_is_read);
		end
		default: begin
			builder_array_muxed26 <= ((main_sdram_cmd_valid & main_sdram_cmd_ready) & main_sdram_cmd_payload_is_read);
		end
	endcase
end
always @(*) begin
	builder_array_muxed27 <= 1'd0;
	case (main_sdram_steerer_sel3)
		1'd0: begin
			builder_array_muxed27 <= 1'd0;
		end
		1'd1: begin
			builder_array_muxed27 <= ((main_sdram_choose_cmd_cmd_valid & main_sdram_choose_cmd_cmd_ready) & main_sdram_choose_cmd_cmd_payload_is_write);
		end
		2'd2: begin
			builder_array_muxed27 <= ((main_sdram_choose_req_cmd_valid & main_sdram_choose_req_cmd_ready) & main_sdram_choose_req_cmd_payload_is_write);
		end
		default: begin
			builder_array_muxed27 <= ((main_sdram_cmd_valid & main_sdram_cmd_ready) & main_sdram_cmd_payload_is_write);
		end
	endcase
end
assign main_uart_rx = builder_regs1;
assign builder_xilinxasyncresetsynchronizerimpl0 = ((~main_locked) | main_reset);
assign builder_xilinxasyncresetsynchronizerimpl1 = ((~main_locked) | main_reset);
assign builder_xilinxasyncresetsynchronizerimpl2 = ((~main_locked) | main_reset);
assign builder_xilinxasyncresetsynchronizerimpl3 = ((~main_locked) | main_reset);
always @(posedge clk200_clk) begin
	if ((main_reset_counter != 1'd0)) begin
		main_reset_counter <= (main_reset_counter - 1'd1);
	end else begin
		main_ic_reset <= 1'd0;
	end
	if (clk200_rst) begin
		main_reset_counter <= 4'd15;
		main_ic_reset <= 1'd1;
	end
end
always @(posedge sys_clk) begin
	if ((main_ctrl_bus_errors != 32'd4294967295)) begin
		if (main_ctrl_bus_error) begin
			main_ctrl_bus_errors <= (main_ctrl_bus_errors + 1'd1);
		end
	end
	main_sram_bus_ack <= 1'd0;
	if (((main_sram_bus_cyc & main_sram_bus_stb) & (~main_sram_bus_ack))) begin
		main_sram_bus_ack <= 1'd1;
	end
	if (main_uart_byte_counter_reset) begin
		main_uart_byte_counter <= 1'd0;
	end else begin
		if (main_uart_byte_counter_ce) begin
			main_uart_byte_counter <= (main_uart_byte_counter + 1'd1);
		end
	end
	if (main_uart_word_counter_reset) begin
		main_uart_word_counter <= 1'd0;
	end else begin
		if (main_uart_word_counter_ce) begin
			main_uart_word_counter <= (main_uart_word_counter + 1'd1);
		end
	end
	if (main_uart_cmd_ce) begin
		main_uart_cmd <= main_uart_source_payload_data;
	end
	if (main_uart_length_ce) begin
		main_uart_length <= main_uart_source_payload_data;
	end
	if (main_uart_address_ce) begin
		main_uart_address <= {main_uart_address[23:0], main_uart_source_payload_data};
	end
	if (main_uart_rx_data_ce) begin
		main_uart_data <= {main_uart_data[23:0], main_uart_source_payload_data};
	end else begin
		if (main_uart_tx_data_ce) begin
			main_uart_data <= main_uart_wishbone_dat_r;
		end
	end
	main_uart_sink_ready <= 1'd0;
	if (((main_uart_sink_valid & (~main_uart_tx_busy)) & (~main_uart_sink_ready))) begin
		main_uart_tx_reg <= main_uart_sink_payload_data;
		main_uart_tx_bitcount <= 1'd0;
		main_uart_tx_busy <= 1'd1;
		serial_tx <= 1'd0;
	end else begin
		if ((main_uart_uart_clk_txen & main_uart_tx_busy)) begin
			main_uart_tx_bitcount <= (main_uart_tx_bitcount + 1'd1);
			if ((main_uart_tx_bitcount == 4'd8)) begin
				serial_tx <= 1'd1;
			end else begin
				if ((main_uart_tx_bitcount == 4'd9)) begin
					serial_tx <= 1'd1;
					main_uart_tx_busy <= 1'd0;
					main_uart_sink_ready <= 1'd1;
				end else begin
					serial_tx <= main_uart_tx_reg[0];
					main_uart_tx_reg <= {1'd0, main_uart_tx_reg[7:1]};
				end
			end
		end
	end
	if (main_uart_tx_busy) begin
		{main_uart_uart_clk_txen, main_uart_phase_accumulator_tx} <= (main_uart_phase_accumulator_tx + main_uart_storage);
	end else begin
		{main_uart_uart_clk_txen, main_uart_phase_accumulator_tx} <= 1'd0;
	end
	main_uart_source_valid <= 1'd0;
	main_uart_rx_r <= main_uart_rx;
	if ((~main_uart_rx_busy)) begin
		if (((~main_uart_rx) & main_uart_rx_r)) begin
			main_uart_rx_busy <= 1'd1;
			main_uart_rx_bitcount <= 1'd0;
		end
	end else begin
		if (main_uart_uart_clk_rxen) begin
			main_uart_rx_bitcount <= (main_uart_rx_bitcount + 1'd1);
			if ((main_uart_rx_bitcount == 1'd0)) begin
				if (main_uart_rx) begin
					main_uart_rx_busy <= 1'd0;
				end
			end else begin
				if ((main_uart_rx_bitcount == 4'd9)) begin
					main_uart_rx_busy <= 1'd0;
					if (main_uart_rx) begin
						main_uart_source_payload_data <= main_uart_rx_reg;
						main_uart_source_valid <= 1'd1;
					end
				end else begin
					main_uart_rx_reg <= {main_uart_rx, main_uart_rx_reg[7:1]};
				end
			end
		end
	end
	if (main_uart_rx_busy) begin
		{main_uart_uart_clk_rxen, main_uart_phase_accumulator_rx} <= (main_uart_phase_accumulator_rx + main_uart_storage);
	end else begin
		{main_uart_uart_clk_rxen, main_uart_phase_accumulator_rx} <= 32'd2147483648;
	end
	builder_uartwishbonebridge_state <= builder_uartwishbonebridge_next_state;
	if (main_uart_reset) begin
		builder_uartwishbonebridge_state <= 3'd0;
	end
	if (main_uart_wait) begin
		if ((~main_uart_done)) begin
			main_uart_count <= (main_uart_count - 1'd1);
		end
	end else begin
		main_uart_count <= 23'd5000000;
	end
	if (main_en_storage) begin
		if ((main_value == 1'd0)) begin
			main_value <= main_reload_storage;
		end else begin
			main_value <= (main_value - 1'd1);
		end
	end else begin
		main_value <= main_load_storage;
	end
	if (main_update_value_re) begin
		main_value_status <= main_value;
	end
	if (main_zero_clear) begin
		main_zero_pending <= 1'd0;
	end
	main_zero_old_trigger <= main_zero_trigger;
	if (((~main_zero_trigger) & main_zero_old_trigger)) begin
		main_zero_pending <= 1'd1;
	end
	builder_wb2csr_state <= builder_wb2csr_next_state;
	if (main_a7ddrphy_dly_sel_storage[0]) begin
		if (main_a7ddrphy_rdly_dq_bitslip_rst_re) begin
			main_a7ddrphy_bitslip0_value <= 1'd0;
		end else begin
			if (main_a7ddrphy_rdly_dq_bitslip_re) begin
				main_a7ddrphy_bitslip0_value <= (main_a7ddrphy_bitslip0_value + 1'd1);
			end
		end
	end
	if (main_a7ddrphy_dly_sel_storage[0]) begin
		if (main_a7ddrphy_rdly_dq_bitslip_rst_re) begin
			main_a7ddrphy_bitslip1_value <= 1'd0;
		end else begin
			if (main_a7ddrphy_rdly_dq_bitslip_re) begin
				main_a7ddrphy_bitslip1_value <= (main_a7ddrphy_bitslip1_value + 1'd1);
			end
		end
	end
	if (main_a7ddrphy_dly_sel_storage[0]) begin
		if (main_a7ddrphy_rdly_dq_bitslip_rst_re) begin
			main_a7ddrphy_bitslip2_value <= 1'd0;
		end else begin
			if (main_a7ddrphy_rdly_dq_bitslip_re) begin
				main_a7ddrphy_bitslip2_value <= (main_a7ddrphy_bitslip2_value + 1'd1);
			end
		end
	end
	if (main_a7ddrphy_dly_sel_storage[0]) begin
		if (main_a7ddrphy_rdly_dq_bitslip_rst_re) begin
			main_a7ddrphy_bitslip3_value <= 1'd0;
		end else begin
			if (main_a7ddrphy_rdly_dq_bitslip_re) begin
				main_a7ddrphy_bitslip3_value <= (main_a7ddrphy_bitslip3_value + 1'd1);
			end
		end
	end
	if (main_a7ddrphy_dly_sel_storage[0]) begin
		if (main_a7ddrphy_rdly_dq_bitslip_rst_re) begin
			main_a7ddrphy_bitslip4_value <= 1'd0;
		end else begin
			if (main_a7ddrphy_rdly_dq_bitslip_re) begin
				main_a7ddrphy_bitslip4_value <= (main_a7ddrphy_bitslip4_value + 1'd1);
			end
		end
	end
	if (main_a7ddrphy_dly_sel_storage[0]) begin
		if (main_a7ddrphy_rdly_dq_bitslip_rst_re) begin
			main_a7ddrphy_bitslip5_value <= 1'd0;
		end else begin
			if (main_a7ddrphy_rdly_dq_bitslip_re) begin
				main_a7ddrphy_bitslip5_value <= (main_a7ddrphy_bitslip5_value + 1'd1);
			end
		end
	end
	if (main_a7ddrphy_dly_sel_storage[0]) begin
		if (main_a7ddrphy_rdly_dq_bitslip_rst_re) begin
			main_a7ddrphy_bitslip6_value <= 1'd0;
		end else begin
			if (main_a7ddrphy_rdly_dq_bitslip_re) begin
				main_a7ddrphy_bitslip6_value <= (main_a7ddrphy_bitslip6_value + 1'd1);
			end
		end
	end
	if (main_a7ddrphy_dly_sel_storage[0]) begin
		if (main_a7ddrphy_rdly_dq_bitslip_rst_re) begin
			main_a7ddrphy_bitslip7_value <= 1'd0;
		end else begin
			if (main_a7ddrphy_rdly_dq_bitslip_re) begin
				main_a7ddrphy_bitslip7_value <= (main_a7ddrphy_bitslip7_value + 1'd1);
			end
		end
	end
	if (main_a7ddrphy_dly_sel_storage[1]) begin
		if (main_a7ddrphy_rdly_dq_bitslip_rst_re) begin
			main_a7ddrphy_bitslip8_value <= 1'd0;
		end else begin
			if (main_a7ddrphy_rdly_dq_bitslip_re) begin
				main_a7ddrphy_bitslip8_value <= (main_a7ddrphy_bitslip8_value + 1'd1);
			end
		end
	end
	if (main_a7ddrphy_dly_sel_storage[1]) begin
		if (main_a7ddrphy_rdly_dq_bitslip_rst_re) begin
			main_a7ddrphy_bitslip9_value <= 1'd0;
		end else begin
			if (main_a7ddrphy_rdly_dq_bitslip_re) begin
				main_a7ddrphy_bitslip9_value <= (main_a7ddrphy_bitslip9_value + 1'd1);
			end
		end
	end
	if (main_a7ddrphy_dly_sel_storage[1]) begin
		if (main_a7ddrphy_rdly_dq_bitslip_rst_re) begin
			main_a7ddrphy_bitslip10_value <= 1'd0;
		end else begin
			if (main_a7ddrphy_rdly_dq_bitslip_re) begin
				main_a7ddrphy_bitslip10_value <= (main_a7ddrphy_bitslip10_value + 1'd1);
			end
		end
	end
	if (main_a7ddrphy_dly_sel_storage[1]) begin
		if (main_a7ddrphy_rdly_dq_bitslip_rst_re) begin
			main_a7ddrphy_bitslip11_value <= 1'd0;
		end else begin
			if (main_a7ddrphy_rdly_dq_bitslip_re) begin
				main_a7ddrphy_bitslip11_value <= (main_a7ddrphy_bitslip11_value + 1'd1);
			end
		end
	end
	if (main_a7ddrphy_dly_sel_storage[1]) begin
		if (main_a7ddrphy_rdly_dq_bitslip_rst_re) begin
			main_a7ddrphy_bitslip12_value <= 1'd0;
		end else begin
			if (main_a7ddrphy_rdly_dq_bitslip_re) begin
				main_a7ddrphy_bitslip12_value <= (main_a7ddrphy_bitslip12_value + 1'd1);
			end
		end
	end
	if (main_a7ddrphy_dly_sel_storage[1]) begin
		if (main_a7ddrphy_rdly_dq_bitslip_rst_re) begin
			main_a7ddrphy_bitslip13_value <= 1'd0;
		end else begin
			if (main_a7ddrphy_rdly_dq_bitslip_re) begin
				main_a7ddrphy_bitslip13_value <= (main_a7ddrphy_bitslip13_value + 1'd1);
			end
		end
	end
	if (main_a7ddrphy_dly_sel_storage[1]) begin
		if (main_a7ddrphy_rdly_dq_bitslip_rst_re) begin
			main_a7ddrphy_bitslip14_value <= 1'd0;
		end else begin
			if (main_a7ddrphy_rdly_dq_bitslip_re) begin
				main_a7ddrphy_bitslip14_value <= (main_a7ddrphy_bitslip14_value + 1'd1);
			end
		end
	end
	if (main_a7ddrphy_dly_sel_storage[1]) begin
		if (main_a7ddrphy_rdly_dq_bitslip_rst_re) begin
			main_a7ddrphy_bitslip15_value <= 1'd0;
		end else begin
			if (main_a7ddrphy_rdly_dq_bitslip_re) begin
				main_a7ddrphy_bitslip15_value <= (main_a7ddrphy_bitslip15_value + 1'd1);
			end
		end
	end
	main_a7ddrphy_n_rddata_en0 <= main_a7ddrphy_dfi_p2_rddata_en;
	main_a7ddrphy_n_rddata_en1 <= main_a7ddrphy_n_rddata_en0;
	main_a7ddrphy_n_rddata_en2 <= main_a7ddrphy_n_rddata_en1;
	main_a7ddrphy_n_rddata_en3 <= main_a7ddrphy_n_rddata_en2;
	main_a7ddrphy_n_rddata_en4 <= main_a7ddrphy_n_rddata_en3;
	main_a7ddrphy_n_rddata_en5 <= main_a7ddrphy_n_rddata_en4;
	main_a7ddrphy_n_rddata_en6 <= main_a7ddrphy_n_rddata_en5;
	main_a7ddrphy_n_rddata_en7 <= main_a7ddrphy_n_rddata_en6;
	main_a7ddrphy_dfi_p0_rddata_valid <= main_a7ddrphy_n_rddata_en7;
	main_a7ddrphy_dfi_p1_rddata_valid <= main_a7ddrphy_n_rddata_en7;
	main_a7ddrphy_dfi_p2_rddata_valid <= main_a7ddrphy_n_rddata_en7;
	main_a7ddrphy_dfi_p3_rddata_valid <= main_a7ddrphy_n_rddata_en7;
	main_a7ddrphy_last_wrdata_en <= {main_a7ddrphy_last_wrdata_en[2:0], main_a7ddrphy_dfi_p3_wrdata_en};
	main_a7ddrphy_oe_dqs <= main_a7ddrphy_oe;
	main_a7ddrphy_oe_dq <= main_a7ddrphy_oe;
	main_a7ddrphy_bitslip0_r <= {main_a7ddrphy_bitslip0_i, main_a7ddrphy_bitslip0_r[15:8]};
	case (main_a7ddrphy_bitslip0_value)
		1'd0: begin
			main_a7ddrphy_bitslip0_o <= main_a7ddrphy_bitslip0_r[7:0];
		end
		1'd1: begin
			main_a7ddrphy_bitslip0_o <= main_a7ddrphy_bitslip0_r[8:1];
		end
		2'd2: begin
			main_a7ddrphy_bitslip0_o <= main_a7ddrphy_bitslip0_r[9:2];
		end
		2'd3: begin
			main_a7ddrphy_bitslip0_o <= main_a7ddrphy_bitslip0_r[10:3];
		end
		3'd4: begin
			main_a7ddrphy_bitslip0_o <= main_a7ddrphy_bitslip0_r[11:4];
		end
		3'd5: begin
			main_a7ddrphy_bitslip0_o <= main_a7ddrphy_bitslip0_r[12:5];
		end
		3'd6: begin
			main_a7ddrphy_bitslip0_o <= main_a7ddrphy_bitslip0_r[13:6];
		end
		3'd7: begin
			main_a7ddrphy_bitslip0_o <= main_a7ddrphy_bitslip0_r[14:7];
		end
	endcase
	main_a7ddrphy_bitslip1_r <= {main_a7ddrphy_bitslip1_i, main_a7ddrphy_bitslip1_r[15:8]};
	case (main_a7ddrphy_bitslip1_value)
		1'd0: begin
			main_a7ddrphy_bitslip1_o <= main_a7ddrphy_bitslip1_r[7:0];
		end
		1'd1: begin
			main_a7ddrphy_bitslip1_o <= main_a7ddrphy_bitslip1_r[8:1];
		end
		2'd2: begin
			main_a7ddrphy_bitslip1_o <= main_a7ddrphy_bitslip1_r[9:2];
		end
		2'd3: begin
			main_a7ddrphy_bitslip1_o <= main_a7ddrphy_bitslip1_r[10:3];
		end
		3'd4: begin
			main_a7ddrphy_bitslip1_o <= main_a7ddrphy_bitslip1_r[11:4];
		end
		3'd5: begin
			main_a7ddrphy_bitslip1_o <= main_a7ddrphy_bitslip1_r[12:5];
		end
		3'd6: begin
			main_a7ddrphy_bitslip1_o <= main_a7ddrphy_bitslip1_r[13:6];
		end
		3'd7: begin
			main_a7ddrphy_bitslip1_o <= main_a7ddrphy_bitslip1_r[14:7];
		end
	endcase
	main_a7ddrphy_bitslip2_r <= {main_a7ddrphy_bitslip2_i, main_a7ddrphy_bitslip2_r[15:8]};
	case (main_a7ddrphy_bitslip2_value)
		1'd0: begin
			main_a7ddrphy_bitslip2_o <= main_a7ddrphy_bitslip2_r[7:0];
		end
		1'd1: begin
			main_a7ddrphy_bitslip2_o <= main_a7ddrphy_bitslip2_r[8:1];
		end
		2'd2: begin
			main_a7ddrphy_bitslip2_o <= main_a7ddrphy_bitslip2_r[9:2];
		end
		2'd3: begin
			main_a7ddrphy_bitslip2_o <= main_a7ddrphy_bitslip2_r[10:3];
		end
		3'd4: begin
			main_a7ddrphy_bitslip2_o <= main_a7ddrphy_bitslip2_r[11:4];
		end
		3'd5: begin
			main_a7ddrphy_bitslip2_o <= main_a7ddrphy_bitslip2_r[12:5];
		end
		3'd6: begin
			main_a7ddrphy_bitslip2_o <= main_a7ddrphy_bitslip2_r[13:6];
		end
		3'd7: begin
			main_a7ddrphy_bitslip2_o <= main_a7ddrphy_bitslip2_r[14:7];
		end
	endcase
	main_a7ddrphy_bitslip3_r <= {main_a7ddrphy_bitslip3_i, main_a7ddrphy_bitslip3_r[15:8]};
	case (main_a7ddrphy_bitslip3_value)
		1'd0: begin
			main_a7ddrphy_bitslip3_o <= main_a7ddrphy_bitslip3_r[7:0];
		end
		1'd1: begin
			main_a7ddrphy_bitslip3_o <= main_a7ddrphy_bitslip3_r[8:1];
		end
		2'd2: begin
			main_a7ddrphy_bitslip3_o <= main_a7ddrphy_bitslip3_r[9:2];
		end
		2'd3: begin
			main_a7ddrphy_bitslip3_o <= main_a7ddrphy_bitslip3_r[10:3];
		end
		3'd4: begin
			main_a7ddrphy_bitslip3_o <= main_a7ddrphy_bitslip3_r[11:4];
		end
		3'd5: begin
			main_a7ddrphy_bitslip3_o <= main_a7ddrphy_bitslip3_r[12:5];
		end
		3'd6: begin
			main_a7ddrphy_bitslip3_o <= main_a7ddrphy_bitslip3_r[13:6];
		end
		3'd7: begin
			main_a7ddrphy_bitslip3_o <= main_a7ddrphy_bitslip3_r[14:7];
		end
	endcase
	main_a7ddrphy_bitslip4_r <= {main_a7ddrphy_bitslip4_i, main_a7ddrphy_bitslip4_r[15:8]};
	case (main_a7ddrphy_bitslip4_value)
		1'd0: begin
			main_a7ddrphy_bitslip4_o <= main_a7ddrphy_bitslip4_r[7:0];
		end
		1'd1: begin
			main_a7ddrphy_bitslip4_o <= main_a7ddrphy_bitslip4_r[8:1];
		end
		2'd2: begin
			main_a7ddrphy_bitslip4_o <= main_a7ddrphy_bitslip4_r[9:2];
		end
		2'd3: begin
			main_a7ddrphy_bitslip4_o <= main_a7ddrphy_bitslip4_r[10:3];
		end
		3'd4: begin
			main_a7ddrphy_bitslip4_o <= main_a7ddrphy_bitslip4_r[11:4];
		end
		3'd5: begin
			main_a7ddrphy_bitslip4_o <= main_a7ddrphy_bitslip4_r[12:5];
		end
		3'd6: begin
			main_a7ddrphy_bitslip4_o <= main_a7ddrphy_bitslip4_r[13:6];
		end
		3'd7: begin
			main_a7ddrphy_bitslip4_o <= main_a7ddrphy_bitslip4_r[14:7];
		end
	endcase
	main_a7ddrphy_bitslip5_r <= {main_a7ddrphy_bitslip5_i, main_a7ddrphy_bitslip5_r[15:8]};
	case (main_a7ddrphy_bitslip5_value)
		1'd0: begin
			main_a7ddrphy_bitslip5_o <= main_a7ddrphy_bitslip5_r[7:0];
		end
		1'd1: begin
			main_a7ddrphy_bitslip5_o <= main_a7ddrphy_bitslip5_r[8:1];
		end
		2'd2: begin
			main_a7ddrphy_bitslip5_o <= main_a7ddrphy_bitslip5_r[9:2];
		end
		2'd3: begin
			main_a7ddrphy_bitslip5_o <= main_a7ddrphy_bitslip5_r[10:3];
		end
		3'd4: begin
			main_a7ddrphy_bitslip5_o <= main_a7ddrphy_bitslip5_r[11:4];
		end
		3'd5: begin
			main_a7ddrphy_bitslip5_o <= main_a7ddrphy_bitslip5_r[12:5];
		end
		3'd6: begin
			main_a7ddrphy_bitslip5_o <= main_a7ddrphy_bitslip5_r[13:6];
		end
		3'd7: begin
			main_a7ddrphy_bitslip5_o <= main_a7ddrphy_bitslip5_r[14:7];
		end
	endcase
	main_a7ddrphy_bitslip6_r <= {main_a7ddrphy_bitslip6_i, main_a7ddrphy_bitslip6_r[15:8]};
	case (main_a7ddrphy_bitslip6_value)
		1'd0: begin
			main_a7ddrphy_bitslip6_o <= main_a7ddrphy_bitslip6_r[7:0];
		end
		1'd1: begin
			main_a7ddrphy_bitslip6_o <= main_a7ddrphy_bitslip6_r[8:1];
		end
		2'd2: begin
			main_a7ddrphy_bitslip6_o <= main_a7ddrphy_bitslip6_r[9:2];
		end
		2'd3: begin
			main_a7ddrphy_bitslip6_o <= main_a7ddrphy_bitslip6_r[10:3];
		end
		3'd4: begin
			main_a7ddrphy_bitslip6_o <= main_a7ddrphy_bitslip6_r[11:4];
		end
		3'd5: begin
			main_a7ddrphy_bitslip6_o <= main_a7ddrphy_bitslip6_r[12:5];
		end
		3'd6: begin
			main_a7ddrphy_bitslip6_o <= main_a7ddrphy_bitslip6_r[13:6];
		end
		3'd7: begin
			main_a7ddrphy_bitslip6_o <= main_a7ddrphy_bitslip6_r[14:7];
		end
	endcase
	main_a7ddrphy_bitslip7_r <= {main_a7ddrphy_bitslip7_i, main_a7ddrphy_bitslip7_r[15:8]};
	case (main_a7ddrphy_bitslip7_value)
		1'd0: begin
			main_a7ddrphy_bitslip7_o <= main_a7ddrphy_bitslip7_r[7:0];
		end
		1'd1: begin
			main_a7ddrphy_bitslip7_o <= main_a7ddrphy_bitslip7_r[8:1];
		end
		2'd2: begin
			main_a7ddrphy_bitslip7_o <= main_a7ddrphy_bitslip7_r[9:2];
		end
		2'd3: begin
			main_a7ddrphy_bitslip7_o <= main_a7ddrphy_bitslip7_r[10:3];
		end
		3'd4: begin
			main_a7ddrphy_bitslip7_o <= main_a7ddrphy_bitslip7_r[11:4];
		end
		3'd5: begin
			main_a7ddrphy_bitslip7_o <= main_a7ddrphy_bitslip7_r[12:5];
		end
		3'd6: begin
			main_a7ddrphy_bitslip7_o <= main_a7ddrphy_bitslip7_r[13:6];
		end
		3'd7: begin
			main_a7ddrphy_bitslip7_o <= main_a7ddrphy_bitslip7_r[14:7];
		end
	endcase
	main_a7ddrphy_bitslip8_r <= {main_a7ddrphy_bitslip8_i, main_a7ddrphy_bitslip8_r[15:8]};
	case (main_a7ddrphy_bitslip8_value)
		1'd0: begin
			main_a7ddrphy_bitslip8_o <= main_a7ddrphy_bitslip8_r[7:0];
		end
		1'd1: begin
			main_a7ddrphy_bitslip8_o <= main_a7ddrphy_bitslip8_r[8:1];
		end
		2'd2: begin
			main_a7ddrphy_bitslip8_o <= main_a7ddrphy_bitslip8_r[9:2];
		end
		2'd3: begin
			main_a7ddrphy_bitslip8_o <= main_a7ddrphy_bitslip8_r[10:3];
		end
		3'd4: begin
			main_a7ddrphy_bitslip8_o <= main_a7ddrphy_bitslip8_r[11:4];
		end
		3'd5: begin
			main_a7ddrphy_bitslip8_o <= main_a7ddrphy_bitslip8_r[12:5];
		end
		3'd6: begin
			main_a7ddrphy_bitslip8_o <= main_a7ddrphy_bitslip8_r[13:6];
		end
		3'd7: begin
			main_a7ddrphy_bitslip8_o <= main_a7ddrphy_bitslip8_r[14:7];
		end
	endcase
	main_a7ddrphy_bitslip9_r <= {main_a7ddrphy_bitslip9_i, main_a7ddrphy_bitslip9_r[15:8]};
	case (main_a7ddrphy_bitslip9_value)
		1'd0: begin
			main_a7ddrphy_bitslip9_o <= main_a7ddrphy_bitslip9_r[7:0];
		end
		1'd1: begin
			main_a7ddrphy_bitslip9_o <= main_a7ddrphy_bitslip9_r[8:1];
		end
		2'd2: begin
			main_a7ddrphy_bitslip9_o <= main_a7ddrphy_bitslip9_r[9:2];
		end
		2'd3: begin
			main_a7ddrphy_bitslip9_o <= main_a7ddrphy_bitslip9_r[10:3];
		end
		3'd4: begin
			main_a7ddrphy_bitslip9_o <= main_a7ddrphy_bitslip9_r[11:4];
		end
		3'd5: begin
			main_a7ddrphy_bitslip9_o <= main_a7ddrphy_bitslip9_r[12:5];
		end
		3'd6: begin
			main_a7ddrphy_bitslip9_o <= main_a7ddrphy_bitslip9_r[13:6];
		end
		3'd7: begin
			main_a7ddrphy_bitslip9_o <= main_a7ddrphy_bitslip9_r[14:7];
		end
	endcase
	main_a7ddrphy_bitslip10_r <= {main_a7ddrphy_bitslip10_i, main_a7ddrphy_bitslip10_r[15:8]};
	case (main_a7ddrphy_bitslip10_value)
		1'd0: begin
			main_a7ddrphy_bitslip10_o <= main_a7ddrphy_bitslip10_r[7:0];
		end
		1'd1: begin
			main_a7ddrphy_bitslip10_o <= main_a7ddrphy_bitslip10_r[8:1];
		end
		2'd2: begin
			main_a7ddrphy_bitslip10_o <= main_a7ddrphy_bitslip10_r[9:2];
		end
		2'd3: begin
			main_a7ddrphy_bitslip10_o <= main_a7ddrphy_bitslip10_r[10:3];
		end
		3'd4: begin
			main_a7ddrphy_bitslip10_o <= main_a7ddrphy_bitslip10_r[11:4];
		end
		3'd5: begin
			main_a7ddrphy_bitslip10_o <= main_a7ddrphy_bitslip10_r[12:5];
		end
		3'd6: begin
			main_a7ddrphy_bitslip10_o <= main_a7ddrphy_bitslip10_r[13:6];
		end
		3'd7: begin
			main_a7ddrphy_bitslip10_o <= main_a7ddrphy_bitslip10_r[14:7];
		end
	endcase
	main_a7ddrphy_bitslip11_r <= {main_a7ddrphy_bitslip11_i, main_a7ddrphy_bitslip11_r[15:8]};
	case (main_a7ddrphy_bitslip11_value)
		1'd0: begin
			main_a7ddrphy_bitslip11_o <= main_a7ddrphy_bitslip11_r[7:0];
		end
		1'd1: begin
			main_a7ddrphy_bitslip11_o <= main_a7ddrphy_bitslip11_r[8:1];
		end
		2'd2: begin
			main_a7ddrphy_bitslip11_o <= main_a7ddrphy_bitslip11_r[9:2];
		end
		2'd3: begin
			main_a7ddrphy_bitslip11_o <= main_a7ddrphy_bitslip11_r[10:3];
		end
		3'd4: begin
			main_a7ddrphy_bitslip11_o <= main_a7ddrphy_bitslip11_r[11:4];
		end
		3'd5: begin
			main_a7ddrphy_bitslip11_o <= main_a7ddrphy_bitslip11_r[12:5];
		end
		3'd6: begin
			main_a7ddrphy_bitslip11_o <= main_a7ddrphy_bitslip11_r[13:6];
		end
		3'd7: begin
			main_a7ddrphy_bitslip11_o <= main_a7ddrphy_bitslip11_r[14:7];
		end
	endcase
	main_a7ddrphy_bitslip12_r <= {main_a7ddrphy_bitslip12_i, main_a7ddrphy_bitslip12_r[15:8]};
	case (main_a7ddrphy_bitslip12_value)
		1'd0: begin
			main_a7ddrphy_bitslip12_o <= main_a7ddrphy_bitslip12_r[7:0];
		end
		1'd1: begin
			main_a7ddrphy_bitslip12_o <= main_a7ddrphy_bitslip12_r[8:1];
		end
		2'd2: begin
			main_a7ddrphy_bitslip12_o <= main_a7ddrphy_bitslip12_r[9:2];
		end
		2'd3: begin
			main_a7ddrphy_bitslip12_o <= main_a7ddrphy_bitslip12_r[10:3];
		end
		3'd4: begin
			main_a7ddrphy_bitslip12_o <= main_a7ddrphy_bitslip12_r[11:4];
		end
		3'd5: begin
			main_a7ddrphy_bitslip12_o <= main_a7ddrphy_bitslip12_r[12:5];
		end
		3'd6: begin
			main_a7ddrphy_bitslip12_o <= main_a7ddrphy_bitslip12_r[13:6];
		end
		3'd7: begin
			main_a7ddrphy_bitslip12_o <= main_a7ddrphy_bitslip12_r[14:7];
		end
	endcase
	main_a7ddrphy_bitslip13_r <= {main_a7ddrphy_bitslip13_i, main_a7ddrphy_bitslip13_r[15:8]};
	case (main_a7ddrphy_bitslip13_value)
		1'd0: begin
			main_a7ddrphy_bitslip13_o <= main_a7ddrphy_bitslip13_r[7:0];
		end
		1'd1: begin
			main_a7ddrphy_bitslip13_o <= main_a7ddrphy_bitslip13_r[8:1];
		end
		2'd2: begin
			main_a7ddrphy_bitslip13_o <= main_a7ddrphy_bitslip13_r[9:2];
		end
		2'd3: begin
			main_a7ddrphy_bitslip13_o <= main_a7ddrphy_bitslip13_r[10:3];
		end
		3'd4: begin
			main_a7ddrphy_bitslip13_o <= main_a7ddrphy_bitslip13_r[11:4];
		end
		3'd5: begin
			main_a7ddrphy_bitslip13_o <= main_a7ddrphy_bitslip13_r[12:5];
		end
		3'd6: begin
			main_a7ddrphy_bitslip13_o <= main_a7ddrphy_bitslip13_r[13:6];
		end
		3'd7: begin
			main_a7ddrphy_bitslip13_o <= main_a7ddrphy_bitslip13_r[14:7];
		end
	endcase
	main_a7ddrphy_bitslip14_r <= {main_a7ddrphy_bitslip14_i, main_a7ddrphy_bitslip14_r[15:8]};
	case (main_a7ddrphy_bitslip14_value)
		1'd0: begin
			main_a7ddrphy_bitslip14_o <= main_a7ddrphy_bitslip14_r[7:0];
		end
		1'd1: begin
			main_a7ddrphy_bitslip14_o <= main_a7ddrphy_bitslip14_r[8:1];
		end
		2'd2: begin
			main_a7ddrphy_bitslip14_o <= main_a7ddrphy_bitslip14_r[9:2];
		end
		2'd3: begin
			main_a7ddrphy_bitslip14_o <= main_a7ddrphy_bitslip14_r[10:3];
		end
		3'd4: begin
			main_a7ddrphy_bitslip14_o <= main_a7ddrphy_bitslip14_r[11:4];
		end
		3'd5: begin
			main_a7ddrphy_bitslip14_o <= main_a7ddrphy_bitslip14_r[12:5];
		end
		3'd6: begin
			main_a7ddrphy_bitslip14_o <= main_a7ddrphy_bitslip14_r[13:6];
		end
		3'd7: begin
			main_a7ddrphy_bitslip14_o <= main_a7ddrphy_bitslip14_r[14:7];
		end
	endcase
	main_a7ddrphy_bitslip15_r <= {main_a7ddrphy_bitslip15_i, main_a7ddrphy_bitslip15_r[15:8]};
	case (main_a7ddrphy_bitslip15_value)
		1'd0: begin
			main_a7ddrphy_bitslip15_o <= main_a7ddrphy_bitslip15_r[7:0];
		end
		1'd1: begin
			main_a7ddrphy_bitslip15_o <= main_a7ddrphy_bitslip15_r[8:1];
		end
		2'd2: begin
			main_a7ddrphy_bitslip15_o <= main_a7ddrphy_bitslip15_r[9:2];
		end
		2'd3: begin
			main_a7ddrphy_bitslip15_o <= main_a7ddrphy_bitslip15_r[10:3];
		end
		3'd4: begin
			main_a7ddrphy_bitslip15_o <= main_a7ddrphy_bitslip15_r[11:4];
		end
		3'd5: begin
			main_a7ddrphy_bitslip15_o <= main_a7ddrphy_bitslip15_r[12:5];
		end
		3'd6: begin
			main_a7ddrphy_bitslip15_o <= main_a7ddrphy_bitslip15_r[13:6];
		end
		3'd7: begin
			main_a7ddrphy_bitslip15_o <= main_a7ddrphy_bitslip15_r[14:7];
		end
	endcase
	if (main_sdram_inti_p0_rddata_valid) begin
		main_sdram_phaseinjector0_status <= main_sdram_inti_p0_rddata;
	end
	if (main_sdram_inti_p1_rddata_valid) begin
		main_sdram_phaseinjector1_status <= main_sdram_inti_p1_rddata;
	end
	if (main_sdram_inti_p2_rddata_valid) begin
		main_sdram_phaseinjector2_status <= main_sdram_inti_p2_rddata;
	end
	if (main_sdram_inti_p3_rddata_valid) begin
		main_sdram_phaseinjector3_status <= main_sdram_inti_p3_rddata;
	end
	if ((main_sdram_timer_wait & (~main_sdram_timer_done0))) begin
		main_sdram_timer_count1 <= (main_sdram_timer_count1 - 1'd1);
	end else begin
		main_sdram_timer_count1 <= 9'd390;
	end
	main_sdram_postponer_req_o <= 1'd0;
	if (main_sdram_postponer_req_i) begin
		main_sdram_postponer_count <= (main_sdram_postponer_count - 1'd1);
		if ((main_sdram_postponer_count == 1'd0)) begin
			main_sdram_postponer_count <= 1'd0;
			main_sdram_postponer_req_o <= 1'd1;
		end
	end
	if (main_sdram_sequencer_start0) begin
		main_sdram_sequencer_count <= 1'd0;
	end else begin
		if (main_sdram_sequencer_done1) begin
			if ((main_sdram_sequencer_count != 1'd0)) begin
				main_sdram_sequencer_count <= (main_sdram_sequencer_count - 1'd1);
			end
		end
	end
	main_sdram_cmd_payload_a <= 1'd0;
	main_sdram_cmd_payload_ba <= 1'd0;
	main_sdram_cmd_payload_cas <= 1'd0;
	main_sdram_cmd_payload_ras <= 1'd0;
	main_sdram_cmd_payload_we <= 1'd0;
	main_sdram_sequencer_done1 <= 1'd0;
	if ((main_sdram_sequencer_start1 & (main_sdram_sequencer_counter == 1'd0))) begin
		main_sdram_cmd_payload_a <= 11'd1024;
		main_sdram_cmd_payload_ba <= 1'd0;
		main_sdram_cmd_payload_cas <= 1'd0;
		main_sdram_cmd_payload_ras <= 1'd1;
		main_sdram_cmd_payload_we <= 1'd1;
	end
	if ((main_sdram_sequencer_counter == 2'd2)) begin
		main_sdram_cmd_payload_a <= 1'd0;
		main_sdram_cmd_payload_ba <= 1'd0;
		main_sdram_cmd_payload_cas <= 1'd1;
		main_sdram_cmd_payload_ras <= 1'd1;
		main_sdram_cmd_payload_we <= 1'd0;
	end
	if ((main_sdram_sequencer_counter == 6'd34)) begin
		main_sdram_cmd_payload_a <= 1'd0;
		main_sdram_cmd_payload_ba <= 1'd0;
		main_sdram_cmd_payload_cas <= 1'd0;
		main_sdram_cmd_payload_ras <= 1'd0;
		main_sdram_cmd_payload_we <= 1'd0;
		main_sdram_sequencer_done1 <= 1'd1;
	end
	if ((main_sdram_sequencer_counter == 6'd34)) begin
		main_sdram_sequencer_counter <= 1'd0;
	end else begin
		if ((main_sdram_sequencer_counter != 1'd0)) begin
			main_sdram_sequencer_counter <= (main_sdram_sequencer_counter + 1'd1);
		end else begin
			if (main_sdram_sequencer_start1) begin
				main_sdram_sequencer_counter <= 1'd1;
			end
		end
	end
	if ((main_sdram_zqcs_timer_wait & (~main_sdram_zqcs_timer_done0))) begin
		main_sdram_zqcs_timer_count1 <= (main_sdram_zqcs_timer_count1 - 1'd1);
	end else begin
		main_sdram_zqcs_timer_count1 <= 26'd49999999;
	end
	main_sdram_zqcs_executer_done <= 1'd0;
	if ((main_sdram_zqcs_executer_start & (main_sdram_zqcs_executer_counter == 1'd0))) begin
		main_sdram_cmd_payload_a <= 11'd1024;
		main_sdram_cmd_payload_ba <= 1'd0;
		main_sdram_cmd_payload_cas <= 1'd0;
		main_sdram_cmd_payload_ras <= 1'd1;
		main_sdram_cmd_payload_we <= 1'd1;
	end
	if ((main_sdram_zqcs_executer_counter == 2'd2)) begin
		main_sdram_cmd_payload_a <= 1'd0;
		main_sdram_cmd_payload_ba <= 1'd0;
		main_sdram_cmd_payload_cas <= 1'd0;
		main_sdram_cmd_payload_ras <= 1'd0;
		main_sdram_cmd_payload_we <= 1'd1;
	end
	if ((main_sdram_zqcs_executer_counter == 5'd18)) begin
		main_sdram_cmd_payload_a <= 1'd0;
		main_sdram_cmd_payload_ba <= 1'd0;
		main_sdram_cmd_payload_cas <= 1'd0;
		main_sdram_cmd_payload_ras <= 1'd0;
		main_sdram_cmd_payload_we <= 1'd0;
		main_sdram_zqcs_executer_done <= 1'd1;
	end
	if ((main_sdram_zqcs_executer_counter == 5'd18)) begin
		main_sdram_zqcs_executer_counter <= 1'd0;
	end else begin
		if ((main_sdram_zqcs_executer_counter != 1'd0)) begin
			main_sdram_zqcs_executer_counter <= (main_sdram_zqcs_executer_counter + 1'd1);
		end else begin
			if (main_sdram_zqcs_executer_start) begin
				main_sdram_zqcs_executer_counter <= 1'd1;
			end
		end
	end
	builder_refresher_state <= builder_refresher_next_state;
	if (main_sdram_bankmachine0_row_close) begin
		main_sdram_bankmachine0_row_opened <= 1'd0;
	end else begin
		if (main_sdram_bankmachine0_row_open) begin
			main_sdram_bankmachine0_row_opened <= 1'd1;
			main_sdram_bankmachine0_row <= main_sdram_bankmachine0_cmd_buffer_source_payload_addr[20:7];
		end
	end
	if (((main_sdram_bankmachine0_cmd_buffer_lookahead_syncfifo0_we & main_sdram_bankmachine0_cmd_buffer_lookahead_syncfifo0_writable) & (~main_sdram_bankmachine0_cmd_buffer_lookahead_replace))) begin
		main_sdram_bankmachine0_cmd_buffer_lookahead_produce <= (main_sdram_bankmachine0_cmd_buffer_lookahead_produce + 1'd1);
	end
	if (main_sdram_bankmachine0_cmd_buffer_lookahead_do_read) begin
		main_sdram_bankmachine0_cmd_buffer_lookahead_consume <= (main_sdram_bankmachine0_cmd_buffer_lookahead_consume + 1'd1);
	end
	if (((main_sdram_bankmachine0_cmd_buffer_lookahead_syncfifo0_we & main_sdram_bankmachine0_cmd_buffer_lookahead_syncfifo0_writable) & (~main_sdram_bankmachine0_cmd_buffer_lookahead_replace))) begin
		if ((~main_sdram_bankmachine0_cmd_buffer_lookahead_do_read)) begin
			main_sdram_bankmachine0_cmd_buffer_lookahead_level <= (main_sdram_bankmachine0_cmd_buffer_lookahead_level + 1'd1);
		end
	end else begin
		if (main_sdram_bankmachine0_cmd_buffer_lookahead_do_read) begin
			main_sdram_bankmachine0_cmd_buffer_lookahead_level <= (main_sdram_bankmachine0_cmd_buffer_lookahead_level - 1'd1);
		end
	end
	if (((~main_sdram_bankmachine0_cmd_buffer_source_valid) | main_sdram_bankmachine0_cmd_buffer_source_ready)) begin
		main_sdram_bankmachine0_cmd_buffer_source_valid <= main_sdram_bankmachine0_cmd_buffer_sink_valid;
		main_sdram_bankmachine0_cmd_buffer_source_first <= main_sdram_bankmachine0_cmd_buffer_sink_first;
		main_sdram_bankmachine0_cmd_buffer_source_last <= main_sdram_bankmachine0_cmd_buffer_sink_last;
		main_sdram_bankmachine0_cmd_buffer_source_payload_we <= main_sdram_bankmachine0_cmd_buffer_sink_payload_we;
		main_sdram_bankmachine0_cmd_buffer_source_payload_addr <= main_sdram_bankmachine0_cmd_buffer_sink_payload_addr;
	end
	if (main_sdram_bankmachine0_twtpcon_valid) begin
		main_sdram_bankmachine0_twtpcon_count <= 3'd4;
		if (1'd0) begin
			main_sdram_bankmachine0_twtpcon_ready <= 1'd1;
		end else begin
			main_sdram_bankmachine0_twtpcon_ready <= 1'd0;
		end
	end else begin
		if ((~main_sdram_bankmachine0_twtpcon_ready)) begin
			main_sdram_bankmachine0_twtpcon_count <= (main_sdram_bankmachine0_twtpcon_count - 1'd1);
			if ((main_sdram_bankmachine0_twtpcon_count == 1'd1)) begin
				main_sdram_bankmachine0_twtpcon_ready <= 1'd1;
			end
		end
	end
	if (main_sdram_bankmachine0_trccon_valid) begin
		main_sdram_bankmachine0_trccon_count <= 2'd3;
		if (1'd0) begin
			main_sdram_bankmachine0_trccon_ready <= 1'd1;
		end else begin
			main_sdram_bankmachine0_trccon_ready <= 1'd0;
		end
	end else begin
		if ((~main_sdram_bankmachine0_trccon_ready)) begin
			main_sdram_bankmachine0_trccon_count <= (main_sdram_bankmachine0_trccon_count - 1'd1);
			if ((main_sdram_bankmachine0_trccon_count == 1'd1)) begin
				main_sdram_bankmachine0_trccon_ready <= 1'd1;
			end
		end
	end
	if (main_sdram_bankmachine0_trascon_valid) begin
		main_sdram_bankmachine0_trascon_count <= 2'd2;
		if (1'd0) begin
			main_sdram_bankmachine0_trascon_ready <= 1'd1;
		end else begin
			main_sdram_bankmachine0_trascon_ready <= 1'd0;
		end
	end else begin
		if ((~main_sdram_bankmachine0_trascon_ready)) begin
			main_sdram_bankmachine0_trascon_count <= (main_sdram_bankmachine0_trascon_count - 1'd1);
			if ((main_sdram_bankmachine0_trascon_count == 1'd1)) begin
				main_sdram_bankmachine0_trascon_ready <= 1'd1;
			end
		end
	end
	builder_bankmachine0_state <= builder_bankmachine0_next_state;
	if (main_sdram_bankmachine1_row_close) begin
		main_sdram_bankmachine1_row_opened <= 1'd0;
	end else begin
		if (main_sdram_bankmachine1_row_open) begin
			main_sdram_bankmachine1_row_opened <= 1'd1;
			main_sdram_bankmachine1_row <= main_sdram_bankmachine1_cmd_buffer_source_payload_addr[20:7];
		end
	end
	if (((main_sdram_bankmachine1_cmd_buffer_lookahead_syncfifo1_we & main_sdram_bankmachine1_cmd_buffer_lookahead_syncfifo1_writable) & (~main_sdram_bankmachine1_cmd_buffer_lookahead_replace))) begin
		main_sdram_bankmachine1_cmd_buffer_lookahead_produce <= (main_sdram_bankmachine1_cmd_buffer_lookahead_produce + 1'd1);
	end
	if (main_sdram_bankmachine1_cmd_buffer_lookahead_do_read) begin
		main_sdram_bankmachine1_cmd_buffer_lookahead_consume <= (main_sdram_bankmachine1_cmd_buffer_lookahead_consume + 1'd1);
	end
	if (((main_sdram_bankmachine1_cmd_buffer_lookahead_syncfifo1_we & main_sdram_bankmachine1_cmd_buffer_lookahead_syncfifo1_writable) & (~main_sdram_bankmachine1_cmd_buffer_lookahead_replace))) begin
		if ((~main_sdram_bankmachine1_cmd_buffer_lookahead_do_read)) begin
			main_sdram_bankmachine1_cmd_buffer_lookahead_level <= (main_sdram_bankmachine1_cmd_buffer_lookahead_level + 1'd1);
		end
	end else begin
		if (main_sdram_bankmachine1_cmd_buffer_lookahead_do_read) begin
			main_sdram_bankmachine1_cmd_buffer_lookahead_level <= (main_sdram_bankmachine1_cmd_buffer_lookahead_level - 1'd1);
		end
	end
	if (((~main_sdram_bankmachine1_cmd_buffer_source_valid) | main_sdram_bankmachine1_cmd_buffer_source_ready)) begin
		main_sdram_bankmachine1_cmd_buffer_source_valid <= main_sdram_bankmachine1_cmd_buffer_sink_valid;
		main_sdram_bankmachine1_cmd_buffer_source_first <= main_sdram_bankmachine1_cmd_buffer_sink_first;
		main_sdram_bankmachine1_cmd_buffer_source_last <= main_sdram_bankmachine1_cmd_buffer_sink_last;
		main_sdram_bankmachine1_cmd_buffer_source_payload_we <= main_sdram_bankmachine1_cmd_buffer_sink_payload_we;
		main_sdram_bankmachine1_cmd_buffer_source_payload_addr <= main_sdram_bankmachine1_cmd_buffer_sink_payload_addr;
	end
	if (main_sdram_bankmachine1_twtpcon_valid) begin
		main_sdram_bankmachine1_twtpcon_count <= 3'd4;
		if (1'd0) begin
			main_sdram_bankmachine1_twtpcon_ready <= 1'd1;
		end else begin
			main_sdram_bankmachine1_twtpcon_ready <= 1'd0;
		end
	end else begin
		if ((~main_sdram_bankmachine1_twtpcon_ready)) begin
			main_sdram_bankmachine1_twtpcon_count <= (main_sdram_bankmachine1_twtpcon_count - 1'd1);
			if ((main_sdram_bankmachine1_twtpcon_count == 1'd1)) begin
				main_sdram_bankmachine1_twtpcon_ready <= 1'd1;
			end
		end
	end
	if (main_sdram_bankmachine1_trccon_valid) begin
		main_sdram_bankmachine1_trccon_count <= 2'd3;
		if (1'd0) begin
			main_sdram_bankmachine1_trccon_ready <= 1'd1;
		end else begin
			main_sdram_bankmachine1_trccon_ready <= 1'd0;
		end
	end else begin
		if ((~main_sdram_bankmachine1_trccon_ready)) begin
			main_sdram_bankmachine1_trccon_count <= (main_sdram_bankmachine1_trccon_count - 1'd1);
			if ((main_sdram_bankmachine1_trccon_count == 1'd1)) begin
				main_sdram_bankmachine1_trccon_ready <= 1'd1;
			end
		end
	end
	if (main_sdram_bankmachine1_trascon_valid) begin
		main_sdram_bankmachine1_trascon_count <= 2'd2;
		if (1'd0) begin
			main_sdram_bankmachine1_trascon_ready <= 1'd1;
		end else begin
			main_sdram_bankmachine1_trascon_ready <= 1'd0;
		end
	end else begin
		if ((~main_sdram_bankmachine1_trascon_ready)) begin
			main_sdram_bankmachine1_trascon_count <= (main_sdram_bankmachine1_trascon_count - 1'd1);
			if ((main_sdram_bankmachine1_trascon_count == 1'd1)) begin
				main_sdram_bankmachine1_trascon_ready <= 1'd1;
			end
		end
	end
	builder_bankmachine1_state <= builder_bankmachine1_next_state;
	if (main_sdram_bankmachine2_row_close) begin
		main_sdram_bankmachine2_row_opened <= 1'd0;
	end else begin
		if (main_sdram_bankmachine2_row_open) begin
			main_sdram_bankmachine2_row_opened <= 1'd1;
			main_sdram_bankmachine2_row <= main_sdram_bankmachine2_cmd_buffer_source_payload_addr[20:7];
		end
	end
	if (((main_sdram_bankmachine2_cmd_buffer_lookahead_syncfifo2_we & main_sdram_bankmachine2_cmd_buffer_lookahead_syncfifo2_writable) & (~main_sdram_bankmachine2_cmd_buffer_lookahead_replace))) begin
		main_sdram_bankmachine2_cmd_buffer_lookahead_produce <= (main_sdram_bankmachine2_cmd_buffer_lookahead_produce + 1'd1);
	end
	if (main_sdram_bankmachine2_cmd_buffer_lookahead_do_read) begin
		main_sdram_bankmachine2_cmd_buffer_lookahead_consume <= (main_sdram_bankmachine2_cmd_buffer_lookahead_consume + 1'd1);
	end
	if (((main_sdram_bankmachine2_cmd_buffer_lookahead_syncfifo2_we & main_sdram_bankmachine2_cmd_buffer_lookahead_syncfifo2_writable) & (~main_sdram_bankmachine2_cmd_buffer_lookahead_replace))) begin
		if ((~main_sdram_bankmachine2_cmd_buffer_lookahead_do_read)) begin
			main_sdram_bankmachine2_cmd_buffer_lookahead_level <= (main_sdram_bankmachine2_cmd_buffer_lookahead_level + 1'd1);
		end
	end else begin
		if (main_sdram_bankmachine2_cmd_buffer_lookahead_do_read) begin
			main_sdram_bankmachine2_cmd_buffer_lookahead_level <= (main_sdram_bankmachine2_cmd_buffer_lookahead_level - 1'd1);
		end
	end
	if (((~main_sdram_bankmachine2_cmd_buffer_source_valid) | main_sdram_bankmachine2_cmd_buffer_source_ready)) begin
		main_sdram_bankmachine2_cmd_buffer_source_valid <= main_sdram_bankmachine2_cmd_buffer_sink_valid;
		main_sdram_bankmachine2_cmd_buffer_source_first <= main_sdram_bankmachine2_cmd_buffer_sink_first;
		main_sdram_bankmachine2_cmd_buffer_source_last <= main_sdram_bankmachine2_cmd_buffer_sink_last;
		main_sdram_bankmachine2_cmd_buffer_source_payload_we <= main_sdram_bankmachine2_cmd_buffer_sink_payload_we;
		main_sdram_bankmachine2_cmd_buffer_source_payload_addr <= main_sdram_bankmachine2_cmd_buffer_sink_payload_addr;
	end
	if (main_sdram_bankmachine2_twtpcon_valid) begin
		main_sdram_bankmachine2_twtpcon_count <= 3'd4;
		if (1'd0) begin
			main_sdram_bankmachine2_twtpcon_ready <= 1'd1;
		end else begin
			main_sdram_bankmachine2_twtpcon_ready <= 1'd0;
		end
	end else begin
		if ((~main_sdram_bankmachine2_twtpcon_ready)) begin
			main_sdram_bankmachine2_twtpcon_count <= (main_sdram_bankmachine2_twtpcon_count - 1'd1);
			if ((main_sdram_bankmachine2_twtpcon_count == 1'd1)) begin
				main_sdram_bankmachine2_twtpcon_ready <= 1'd1;
			end
		end
	end
	if (main_sdram_bankmachine2_trccon_valid) begin
		main_sdram_bankmachine2_trccon_count <= 2'd3;
		if (1'd0) begin
			main_sdram_bankmachine2_trccon_ready <= 1'd1;
		end else begin
			main_sdram_bankmachine2_trccon_ready <= 1'd0;
		end
	end else begin
		if ((~main_sdram_bankmachine2_trccon_ready)) begin
			main_sdram_bankmachine2_trccon_count <= (main_sdram_bankmachine2_trccon_count - 1'd1);
			if ((main_sdram_bankmachine2_trccon_count == 1'd1)) begin
				main_sdram_bankmachine2_trccon_ready <= 1'd1;
			end
		end
	end
	if (main_sdram_bankmachine2_trascon_valid) begin
		main_sdram_bankmachine2_trascon_count <= 2'd2;
		if (1'd0) begin
			main_sdram_bankmachine2_trascon_ready <= 1'd1;
		end else begin
			main_sdram_bankmachine2_trascon_ready <= 1'd0;
		end
	end else begin
		if ((~main_sdram_bankmachine2_trascon_ready)) begin
			main_sdram_bankmachine2_trascon_count <= (main_sdram_bankmachine2_trascon_count - 1'd1);
			if ((main_sdram_bankmachine2_trascon_count == 1'd1)) begin
				main_sdram_bankmachine2_trascon_ready <= 1'd1;
			end
		end
	end
	builder_bankmachine2_state <= builder_bankmachine2_next_state;
	if (main_sdram_bankmachine3_row_close) begin
		main_sdram_bankmachine3_row_opened <= 1'd0;
	end else begin
		if (main_sdram_bankmachine3_row_open) begin
			main_sdram_bankmachine3_row_opened <= 1'd1;
			main_sdram_bankmachine3_row <= main_sdram_bankmachine3_cmd_buffer_source_payload_addr[20:7];
		end
	end
	if (((main_sdram_bankmachine3_cmd_buffer_lookahead_syncfifo3_we & main_sdram_bankmachine3_cmd_buffer_lookahead_syncfifo3_writable) & (~main_sdram_bankmachine3_cmd_buffer_lookahead_replace))) begin
		main_sdram_bankmachine3_cmd_buffer_lookahead_produce <= (main_sdram_bankmachine3_cmd_buffer_lookahead_produce + 1'd1);
	end
	if (main_sdram_bankmachine3_cmd_buffer_lookahead_do_read) begin
		main_sdram_bankmachine3_cmd_buffer_lookahead_consume <= (main_sdram_bankmachine3_cmd_buffer_lookahead_consume + 1'd1);
	end
	if (((main_sdram_bankmachine3_cmd_buffer_lookahead_syncfifo3_we & main_sdram_bankmachine3_cmd_buffer_lookahead_syncfifo3_writable) & (~main_sdram_bankmachine3_cmd_buffer_lookahead_replace))) begin
		if ((~main_sdram_bankmachine3_cmd_buffer_lookahead_do_read)) begin
			main_sdram_bankmachine3_cmd_buffer_lookahead_level <= (main_sdram_bankmachine3_cmd_buffer_lookahead_level + 1'd1);
		end
	end else begin
		if (main_sdram_bankmachine3_cmd_buffer_lookahead_do_read) begin
			main_sdram_bankmachine3_cmd_buffer_lookahead_level <= (main_sdram_bankmachine3_cmd_buffer_lookahead_level - 1'd1);
		end
	end
	if (((~main_sdram_bankmachine3_cmd_buffer_source_valid) | main_sdram_bankmachine3_cmd_buffer_source_ready)) begin
		main_sdram_bankmachine3_cmd_buffer_source_valid <= main_sdram_bankmachine3_cmd_buffer_sink_valid;
		main_sdram_bankmachine3_cmd_buffer_source_first <= main_sdram_bankmachine3_cmd_buffer_sink_first;
		main_sdram_bankmachine3_cmd_buffer_source_last <= main_sdram_bankmachine3_cmd_buffer_sink_last;
		main_sdram_bankmachine3_cmd_buffer_source_payload_we <= main_sdram_bankmachine3_cmd_buffer_sink_payload_we;
		main_sdram_bankmachine3_cmd_buffer_source_payload_addr <= main_sdram_bankmachine3_cmd_buffer_sink_payload_addr;
	end
	if (main_sdram_bankmachine3_twtpcon_valid) begin
		main_sdram_bankmachine3_twtpcon_count <= 3'd4;
		if (1'd0) begin
			main_sdram_bankmachine3_twtpcon_ready <= 1'd1;
		end else begin
			main_sdram_bankmachine3_twtpcon_ready <= 1'd0;
		end
	end else begin
		if ((~main_sdram_bankmachine3_twtpcon_ready)) begin
			main_sdram_bankmachine3_twtpcon_count <= (main_sdram_bankmachine3_twtpcon_count - 1'd1);
			if ((main_sdram_bankmachine3_twtpcon_count == 1'd1)) begin
				main_sdram_bankmachine3_twtpcon_ready <= 1'd1;
			end
		end
	end
	if (main_sdram_bankmachine3_trccon_valid) begin
		main_sdram_bankmachine3_trccon_count <= 2'd3;
		if (1'd0) begin
			main_sdram_bankmachine3_trccon_ready <= 1'd1;
		end else begin
			main_sdram_bankmachine3_trccon_ready <= 1'd0;
		end
	end else begin
		if ((~main_sdram_bankmachine3_trccon_ready)) begin
			main_sdram_bankmachine3_trccon_count <= (main_sdram_bankmachine3_trccon_count - 1'd1);
			if ((main_sdram_bankmachine3_trccon_count == 1'd1)) begin
				main_sdram_bankmachine3_trccon_ready <= 1'd1;
			end
		end
	end
	if (main_sdram_bankmachine3_trascon_valid) begin
		main_sdram_bankmachine3_trascon_count <= 2'd2;
		if (1'd0) begin
			main_sdram_bankmachine3_trascon_ready <= 1'd1;
		end else begin
			main_sdram_bankmachine3_trascon_ready <= 1'd0;
		end
	end else begin
		if ((~main_sdram_bankmachine3_trascon_ready)) begin
			main_sdram_bankmachine3_trascon_count <= (main_sdram_bankmachine3_trascon_count - 1'd1);
			if ((main_sdram_bankmachine3_trascon_count == 1'd1)) begin
				main_sdram_bankmachine3_trascon_ready <= 1'd1;
			end
		end
	end
	builder_bankmachine3_state <= builder_bankmachine3_next_state;
	if (main_sdram_bankmachine4_row_close) begin
		main_sdram_bankmachine4_row_opened <= 1'd0;
	end else begin
		if (main_sdram_bankmachine4_row_open) begin
			main_sdram_bankmachine4_row_opened <= 1'd1;
			main_sdram_bankmachine4_row <= main_sdram_bankmachine4_cmd_buffer_source_payload_addr[20:7];
		end
	end
	if (((main_sdram_bankmachine4_cmd_buffer_lookahead_syncfifo4_we & main_sdram_bankmachine4_cmd_buffer_lookahead_syncfifo4_writable) & (~main_sdram_bankmachine4_cmd_buffer_lookahead_replace))) begin
		main_sdram_bankmachine4_cmd_buffer_lookahead_produce <= (main_sdram_bankmachine4_cmd_buffer_lookahead_produce + 1'd1);
	end
	if (main_sdram_bankmachine4_cmd_buffer_lookahead_do_read) begin
		main_sdram_bankmachine4_cmd_buffer_lookahead_consume <= (main_sdram_bankmachine4_cmd_buffer_lookahead_consume + 1'd1);
	end
	if (((main_sdram_bankmachine4_cmd_buffer_lookahead_syncfifo4_we & main_sdram_bankmachine4_cmd_buffer_lookahead_syncfifo4_writable) & (~main_sdram_bankmachine4_cmd_buffer_lookahead_replace))) begin
		if ((~main_sdram_bankmachine4_cmd_buffer_lookahead_do_read)) begin
			main_sdram_bankmachine4_cmd_buffer_lookahead_level <= (main_sdram_bankmachine4_cmd_buffer_lookahead_level + 1'd1);
		end
	end else begin
		if (main_sdram_bankmachine4_cmd_buffer_lookahead_do_read) begin
			main_sdram_bankmachine4_cmd_buffer_lookahead_level <= (main_sdram_bankmachine4_cmd_buffer_lookahead_level - 1'd1);
		end
	end
	if (((~main_sdram_bankmachine4_cmd_buffer_source_valid) | main_sdram_bankmachine4_cmd_buffer_source_ready)) begin
		main_sdram_bankmachine4_cmd_buffer_source_valid <= main_sdram_bankmachine4_cmd_buffer_sink_valid;
		main_sdram_bankmachine4_cmd_buffer_source_first <= main_sdram_bankmachine4_cmd_buffer_sink_first;
		main_sdram_bankmachine4_cmd_buffer_source_last <= main_sdram_bankmachine4_cmd_buffer_sink_last;
		main_sdram_bankmachine4_cmd_buffer_source_payload_we <= main_sdram_bankmachine4_cmd_buffer_sink_payload_we;
		main_sdram_bankmachine4_cmd_buffer_source_payload_addr <= main_sdram_bankmachine4_cmd_buffer_sink_payload_addr;
	end
	if (main_sdram_bankmachine4_twtpcon_valid) begin
		main_sdram_bankmachine4_twtpcon_count <= 3'd4;
		if (1'd0) begin
			main_sdram_bankmachine4_twtpcon_ready <= 1'd1;
		end else begin
			main_sdram_bankmachine4_twtpcon_ready <= 1'd0;
		end
	end else begin
		if ((~main_sdram_bankmachine4_twtpcon_ready)) begin
			main_sdram_bankmachine4_twtpcon_count <= (main_sdram_bankmachine4_twtpcon_count - 1'd1);
			if ((main_sdram_bankmachine4_twtpcon_count == 1'd1)) begin
				main_sdram_bankmachine4_twtpcon_ready <= 1'd1;
			end
		end
	end
	if (main_sdram_bankmachine4_trccon_valid) begin
		main_sdram_bankmachine4_trccon_count <= 2'd3;
		if (1'd0) begin
			main_sdram_bankmachine4_trccon_ready <= 1'd1;
		end else begin
			main_sdram_bankmachine4_trccon_ready <= 1'd0;
		end
	end else begin
		if ((~main_sdram_bankmachine4_trccon_ready)) begin
			main_sdram_bankmachine4_trccon_count <= (main_sdram_bankmachine4_trccon_count - 1'd1);
			if ((main_sdram_bankmachine4_trccon_count == 1'd1)) begin
				main_sdram_bankmachine4_trccon_ready <= 1'd1;
			end
		end
	end
	if (main_sdram_bankmachine4_trascon_valid) begin
		main_sdram_bankmachine4_trascon_count <= 2'd2;
		if (1'd0) begin
			main_sdram_bankmachine4_trascon_ready <= 1'd1;
		end else begin
			main_sdram_bankmachine4_trascon_ready <= 1'd0;
		end
	end else begin
		if ((~main_sdram_bankmachine4_trascon_ready)) begin
			main_sdram_bankmachine4_trascon_count <= (main_sdram_bankmachine4_trascon_count - 1'd1);
			if ((main_sdram_bankmachine4_trascon_count == 1'd1)) begin
				main_sdram_bankmachine4_trascon_ready <= 1'd1;
			end
		end
	end
	builder_bankmachine4_state <= builder_bankmachine4_next_state;
	if (main_sdram_bankmachine5_row_close) begin
		main_sdram_bankmachine5_row_opened <= 1'd0;
	end else begin
		if (main_sdram_bankmachine5_row_open) begin
			main_sdram_bankmachine5_row_opened <= 1'd1;
			main_sdram_bankmachine5_row <= main_sdram_bankmachine5_cmd_buffer_source_payload_addr[20:7];
		end
	end
	if (((main_sdram_bankmachine5_cmd_buffer_lookahead_syncfifo5_we & main_sdram_bankmachine5_cmd_buffer_lookahead_syncfifo5_writable) & (~main_sdram_bankmachine5_cmd_buffer_lookahead_replace))) begin
		main_sdram_bankmachine5_cmd_buffer_lookahead_produce <= (main_sdram_bankmachine5_cmd_buffer_lookahead_produce + 1'd1);
	end
	if (main_sdram_bankmachine5_cmd_buffer_lookahead_do_read) begin
		main_sdram_bankmachine5_cmd_buffer_lookahead_consume <= (main_sdram_bankmachine5_cmd_buffer_lookahead_consume + 1'd1);
	end
	if (((main_sdram_bankmachine5_cmd_buffer_lookahead_syncfifo5_we & main_sdram_bankmachine5_cmd_buffer_lookahead_syncfifo5_writable) & (~main_sdram_bankmachine5_cmd_buffer_lookahead_replace))) begin
		if ((~main_sdram_bankmachine5_cmd_buffer_lookahead_do_read)) begin
			main_sdram_bankmachine5_cmd_buffer_lookahead_level <= (main_sdram_bankmachine5_cmd_buffer_lookahead_level + 1'd1);
		end
	end else begin
		if (main_sdram_bankmachine5_cmd_buffer_lookahead_do_read) begin
			main_sdram_bankmachine5_cmd_buffer_lookahead_level <= (main_sdram_bankmachine5_cmd_buffer_lookahead_level - 1'd1);
		end
	end
	if (((~main_sdram_bankmachine5_cmd_buffer_source_valid) | main_sdram_bankmachine5_cmd_buffer_source_ready)) begin
		main_sdram_bankmachine5_cmd_buffer_source_valid <= main_sdram_bankmachine5_cmd_buffer_sink_valid;
		main_sdram_bankmachine5_cmd_buffer_source_first <= main_sdram_bankmachine5_cmd_buffer_sink_first;
		main_sdram_bankmachine5_cmd_buffer_source_last <= main_sdram_bankmachine5_cmd_buffer_sink_last;
		main_sdram_bankmachine5_cmd_buffer_source_payload_we <= main_sdram_bankmachine5_cmd_buffer_sink_payload_we;
		main_sdram_bankmachine5_cmd_buffer_source_payload_addr <= main_sdram_bankmachine5_cmd_buffer_sink_payload_addr;
	end
	if (main_sdram_bankmachine5_twtpcon_valid) begin
		main_sdram_bankmachine5_twtpcon_count <= 3'd4;
		if (1'd0) begin
			main_sdram_bankmachine5_twtpcon_ready <= 1'd1;
		end else begin
			main_sdram_bankmachine5_twtpcon_ready <= 1'd0;
		end
	end else begin
		if ((~main_sdram_bankmachine5_twtpcon_ready)) begin
			main_sdram_bankmachine5_twtpcon_count <= (main_sdram_bankmachine5_twtpcon_count - 1'd1);
			if ((main_sdram_bankmachine5_twtpcon_count == 1'd1)) begin
				main_sdram_bankmachine5_twtpcon_ready <= 1'd1;
			end
		end
	end
	if (main_sdram_bankmachine5_trccon_valid) begin
		main_sdram_bankmachine5_trccon_count <= 2'd3;
		if (1'd0) begin
			main_sdram_bankmachine5_trccon_ready <= 1'd1;
		end else begin
			main_sdram_bankmachine5_trccon_ready <= 1'd0;
		end
	end else begin
		if ((~main_sdram_bankmachine5_trccon_ready)) begin
			main_sdram_bankmachine5_trccon_count <= (main_sdram_bankmachine5_trccon_count - 1'd1);
			if ((main_sdram_bankmachine5_trccon_count == 1'd1)) begin
				main_sdram_bankmachine5_trccon_ready <= 1'd1;
			end
		end
	end
	if (main_sdram_bankmachine5_trascon_valid) begin
		main_sdram_bankmachine5_trascon_count <= 2'd2;
		if (1'd0) begin
			main_sdram_bankmachine5_trascon_ready <= 1'd1;
		end else begin
			main_sdram_bankmachine5_trascon_ready <= 1'd0;
		end
	end else begin
		if ((~main_sdram_bankmachine5_trascon_ready)) begin
			main_sdram_bankmachine5_trascon_count <= (main_sdram_bankmachine5_trascon_count - 1'd1);
			if ((main_sdram_bankmachine5_trascon_count == 1'd1)) begin
				main_sdram_bankmachine5_trascon_ready <= 1'd1;
			end
		end
	end
	builder_bankmachine5_state <= builder_bankmachine5_next_state;
	if (main_sdram_bankmachine6_row_close) begin
		main_sdram_bankmachine6_row_opened <= 1'd0;
	end else begin
		if (main_sdram_bankmachine6_row_open) begin
			main_sdram_bankmachine6_row_opened <= 1'd1;
			main_sdram_bankmachine6_row <= main_sdram_bankmachine6_cmd_buffer_source_payload_addr[20:7];
		end
	end
	if (((main_sdram_bankmachine6_cmd_buffer_lookahead_syncfifo6_we & main_sdram_bankmachine6_cmd_buffer_lookahead_syncfifo6_writable) & (~main_sdram_bankmachine6_cmd_buffer_lookahead_replace))) begin
		main_sdram_bankmachine6_cmd_buffer_lookahead_produce <= (main_sdram_bankmachine6_cmd_buffer_lookahead_produce + 1'd1);
	end
	if (main_sdram_bankmachine6_cmd_buffer_lookahead_do_read) begin
		main_sdram_bankmachine6_cmd_buffer_lookahead_consume <= (main_sdram_bankmachine6_cmd_buffer_lookahead_consume + 1'd1);
	end
	if (((main_sdram_bankmachine6_cmd_buffer_lookahead_syncfifo6_we & main_sdram_bankmachine6_cmd_buffer_lookahead_syncfifo6_writable) & (~main_sdram_bankmachine6_cmd_buffer_lookahead_replace))) begin
		if ((~main_sdram_bankmachine6_cmd_buffer_lookahead_do_read)) begin
			main_sdram_bankmachine6_cmd_buffer_lookahead_level <= (main_sdram_bankmachine6_cmd_buffer_lookahead_level + 1'd1);
		end
	end else begin
		if (main_sdram_bankmachine6_cmd_buffer_lookahead_do_read) begin
			main_sdram_bankmachine6_cmd_buffer_lookahead_level <= (main_sdram_bankmachine6_cmd_buffer_lookahead_level - 1'd1);
		end
	end
	if (((~main_sdram_bankmachine6_cmd_buffer_source_valid) | main_sdram_bankmachine6_cmd_buffer_source_ready)) begin
		main_sdram_bankmachine6_cmd_buffer_source_valid <= main_sdram_bankmachine6_cmd_buffer_sink_valid;
		main_sdram_bankmachine6_cmd_buffer_source_first <= main_sdram_bankmachine6_cmd_buffer_sink_first;
		main_sdram_bankmachine6_cmd_buffer_source_last <= main_sdram_bankmachine6_cmd_buffer_sink_last;
		main_sdram_bankmachine6_cmd_buffer_source_payload_we <= main_sdram_bankmachine6_cmd_buffer_sink_payload_we;
		main_sdram_bankmachine6_cmd_buffer_source_payload_addr <= main_sdram_bankmachine6_cmd_buffer_sink_payload_addr;
	end
	if (main_sdram_bankmachine6_twtpcon_valid) begin
		main_sdram_bankmachine6_twtpcon_count <= 3'd4;
		if (1'd0) begin
			main_sdram_bankmachine6_twtpcon_ready <= 1'd1;
		end else begin
			main_sdram_bankmachine6_twtpcon_ready <= 1'd0;
		end
	end else begin
		if ((~main_sdram_bankmachine6_twtpcon_ready)) begin
			main_sdram_bankmachine6_twtpcon_count <= (main_sdram_bankmachine6_twtpcon_count - 1'd1);
			if ((main_sdram_bankmachine6_twtpcon_count == 1'd1)) begin
				main_sdram_bankmachine6_twtpcon_ready <= 1'd1;
			end
		end
	end
	if (main_sdram_bankmachine6_trccon_valid) begin
		main_sdram_bankmachine6_trccon_count <= 2'd3;
		if (1'd0) begin
			main_sdram_bankmachine6_trccon_ready <= 1'd1;
		end else begin
			main_sdram_bankmachine6_trccon_ready <= 1'd0;
		end
	end else begin
		if ((~main_sdram_bankmachine6_trccon_ready)) begin
			main_sdram_bankmachine6_trccon_count <= (main_sdram_bankmachine6_trccon_count - 1'd1);
			if ((main_sdram_bankmachine6_trccon_count == 1'd1)) begin
				main_sdram_bankmachine6_trccon_ready <= 1'd1;
			end
		end
	end
	if (main_sdram_bankmachine6_trascon_valid) begin
		main_sdram_bankmachine6_trascon_count <= 2'd2;
		if (1'd0) begin
			main_sdram_bankmachine6_trascon_ready <= 1'd1;
		end else begin
			main_sdram_bankmachine6_trascon_ready <= 1'd0;
		end
	end else begin
		if ((~main_sdram_bankmachine6_trascon_ready)) begin
			main_sdram_bankmachine6_trascon_count <= (main_sdram_bankmachine6_trascon_count - 1'd1);
			if ((main_sdram_bankmachine6_trascon_count == 1'd1)) begin
				main_sdram_bankmachine6_trascon_ready <= 1'd1;
			end
		end
	end
	builder_bankmachine6_state <= builder_bankmachine6_next_state;
	if (main_sdram_bankmachine7_row_close) begin
		main_sdram_bankmachine7_row_opened <= 1'd0;
	end else begin
		if (main_sdram_bankmachine7_row_open) begin
			main_sdram_bankmachine7_row_opened <= 1'd1;
			main_sdram_bankmachine7_row <= main_sdram_bankmachine7_cmd_buffer_source_payload_addr[20:7];
		end
	end
	if (((main_sdram_bankmachine7_cmd_buffer_lookahead_syncfifo7_we & main_sdram_bankmachine7_cmd_buffer_lookahead_syncfifo7_writable) & (~main_sdram_bankmachine7_cmd_buffer_lookahead_replace))) begin
		main_sdram_bankmachine7_cmd_buffer_lookahead_produce <= (main_sdram_bankmachine7_cmd_buffer_lookahead_produce + 1'd1);
	end
	if (main_sdram_bankmachine7_cmd_buffer_lookahead_do_read) begin
		main_sdram_bankmachine7_cmd_buffer_lookahead_consume <= (main_sdram_bankmachine7_cmd_buffer_lookahead_consume + 1'd1);
	end
	if (((main_sdram_bankmachine7_cmd_buffer_lookahead_syncfifo7_we & main_sdram_bankmachine7_cmd_buffer_lookahead_syncfifo7_writable) & (~main_sdram_bankmachine7_cmd_buffer_lookahead_replace))) begin
		if ((~main_sdram_bankmachine7_cmd_buffer_lookahead_do_read)) begin
			main_sdram_bankmachine7_cmd_buffer_lookahead_level <= (main_sdram_bankmachine7_cmd_buffer_lookahead_level + 1'd1);
		end
	end else begin
		if (main_sdram_bankmachine7_cmd_buffer_lookahead_do_read) begin
			main_sdram_bankmachine7_cmd_buffer_lookahead_level <= (main_sdram_bankmachine7_cmd_buffer_lookahead_level - 1'd1);
		end
	end
	if (((~main_sdram_bankmachine7_cmd_buffer_source_valid) | main_sdram_bankmachine7_cmd_buffer_source_ready)) begin
		main_sdram_bankmachine7_cmd_buffer_source_valid <= main_sdram_bankmachine7_cmd_buffer_sink_valid;
		main_sdram_bankmachine7_cmd_buffer_source_first <= main_sdram_bankmachine7_cmd_buffer_sink_first;
		main_sdram_bankmachine7_cmd_buffer_source_last <= main_sdram_bankmachine7_cmd_buffer_sink_last;
		main_sdram_bankmachine7_cmd_buffer_source_payload_we <= main_sdram_bankmachine7_cmd_buffer_sink_payload_we;
		main_sdram_bankmachine7_cmd_buffer_source_payload_addr <= main_sdram_bankmachine7_cmd_buffer_sink_payload_addr;
	end
	if (main_sdram_bankmachine7_twtpcon_valid) begin
		main_sdram_bankmachine7_twtpcon_count <= 3'd4;
		if (1'd0) begin
			main_sdram_bankmachine7_twtpcon_ready <= 1'd1;
		end else begin
			main_sdram_bankmachine7_twtpcon_ready <= 1'd0;
		end
	end else begin
		if ((~main_sdram_bankmachine7_twtpcon_ready)) begin
			main_sdram_bankmachine7_twtpcon_count <= (main_sdram_bankmachine7_twtpcon_count - 1'd1);
			if ((main_sdram_bankmachine7_twtpcon_count == 1'd1)) begin
				main_sdram_bankmachine7_twtpcon_ready <= 1'd1;
			end
		end
	end
	if (main_sdram_bankmachine7_trccon_valid) begin
		main_sdram_bankmachine7_trccon_count <= 2'd3;
		if (1'd0) begin
			main_sdram_bankmachine7_trccon_ready <= 1'd1;
		end else begin
			main_sdram_bankmachine7_trccon_ready <= 1'd0;
		end
	end else begin
		if ((~main_sdram_bankmachine7_trccon_ready)) begin
			main_sdram_bankmachine7_trccon_count <= (main_sdram_bankmachine7_trccon_count - 1'd1);
			if ((main_sdram_bankmachine7_trccon_count == 1'd1)) begin
				main_sdram_bankmachine7_trccon_ready <= 1'd1;
			end
		end
	end
	if (main_sdram_bankmachine7_trascon_valid) begin
		main_sdram_bankmachine7_trascon_count <= 2'd2;
		if (1'd0) begin
			main_sdram_bankmachine7_trascon_ready <= 1'd1;
		end else begin
			main_sdram_bankmachine7_trascon_ready <= 1'd0;
		end
	end else begin
		if ((~main_sdram_bankmachine7_trascon_ready)) begin
			main_sdram_bankmachine7_trascon_count <= (main_sdram_bankmachine7_trascon_count - 1'd1);
			if ((main_sdram_bankmachine7_trascon_count == 1'd1)) begin
				main_sdram_bankmachine7_trascon_ready <= 1'd1;
			end
		end
	end
	builder_bankmachine7_state <= builder_bankmachine7_next_state;
	if ((~main_sdram_en0)) begin
		main_sdram_time0 <= 5'd31;
	end else begin
		if ((~main_sdram_max_time0)) begin
			main_sdram_time0 <= (main_sdram_time0 - 1'd1);
		end
	end
	if ((~main_sdram_en1)) begin
		main_sdram_time1 <= 4'd15;
	end else begin
		if ((~main_sdram_max_time1)) begin
			main_sdram_time1 <= (main_sdram_time1 - 1'd1);
		end
	end
	if (main_sdram_choose_cmd_ce) begin
		case (main_sdram_choose_cmd_grant)
			1'd0: begin
				if (main_sdram_choose_cmd_request[1]) begin
					main_sdram_choose_cmd_grant <= 1'd1;
				end else begin
					if (main_sdram_choose_cmd_request[2]) begin
						main_sdram_choose_cmd_grant <= 2'd2;
					end else begin
						if (main_sdram_choose_cmd_request[3]) begin
							main_sdram_choose_cmd_grant <= 2'd3;
						end else begin
							if (main_sdram_choose_cmd_request[4]) begin
								main_sdram_choose_cmd_grant <= 3'd4;
							end else begin
								if (main_sdram_choose_cmd_request[5]) begin
									main_sdram_choose_cmd_grant <= 3'd5;
								end else begin
									if (main_sdram_choose_cmd_request[6]) begin
										main_sdram_choose_cmd_grant <= 3'd6;
									end else begin
										if (main_sdram_choose_cmd_request[7]) begin
											main_sdram_choose_cmd_grant <= 3'd7;
										end
									end
								end
							end
						end
					end
				end
			end
			1'd1: begin
				if (main_sdram_choose_cmd_request[2]) begin
					main_sdram_choose_cmd_grant <= 2'd2;
				end else begin
					if (main_sdram_choose_cmd_request[3]) begin
						main_sdram_choose_cmd_grant <= 2'd3;
					end else begin
						if (main_sdram_choose_cmd_request[4]) begin
							main_sdram_choose_cmd_grant <= 3'd4;
						end else begin
							if (main_sdram_choose_cmd_request[5]) begin
								main_sdram_choose_cmd_grant <= 3'd5;
							end else begin
								if (main_sdram_choose_cmd_request[6]) begin
									main_sdram_choose_cmd_grant <= 3'd6;
								end else begin
									if (main_sdram_choose_cmd_request[7]) begin
										main_sdram_choose_cmd_grant <= 3'd7;
									end else begin
										if (main_sdram_choose_cmd_request[0]) begin
											main_sdram_choose_cmd_grant <= 1'd0;
										end
									end
								end
							end
						end
					end
				end
			end
			2'd2: begin
				if (main_sdram_choose_cmd_request[3]) begin
					main_sdram_choose_cmd_grant <= 2'd3;
				end else begin
					if (main_sdram_choose_cmd_request[4]) begin
						main_sdram_choose_cmd_grant <= 3'd4;
					end else begin
						if (main_sdram_choose_cmd_request[5]) begin
							main_sdram_choose_cmd_grant <= 3'd5;
						end else begin
							if (main_sdram_choose_cmd_request[6]) begin
								main_sdram_choose_cmd_grant <= 3'd6;
							end else begin
								if (main_sdram_choose_cmd_request[7]) begin
									main_sdram_choose_cmd_grant <= 3'd7;
								end else begin
									if (main_sdram_choose_cmd_request[0]) begin
										main_sdram_choose_cmd_grant <= 1'd0;
									end else begin
										if (main_sdram_choose_cmd_request[1]) begin
											main_sdram_choose_cmd_grant <= 1'd1;
										end
									end
								end
							end
						end
					end
				end
			end
			2'd3: begin
				if (main_sdram_choose_cmd_request[4]) begin
					main_sdram_choose_cmd_grant <= 3'd4;
				end else begin
					if (main_sdram_choose_cmd_request[5]) begin
						main_sdram_choose_cmd_grant <= 3'd5;
					end else begin
						if (main_sdram_choose_cmd_request[6]) begin
							main_sdram_choose_cmd_grant <= 3'd6;
						end else begin
							if (main_sdram_choose_cmd_request[7]) begin
								main_sdram_choose_cmd_grant <= 3'd7;
							end else begin
								if (main_sdram_choose_cmd_request[0]) begin
									main_sdram_choose_cmd_grant <= 1'd0;
								end else begin
									if (main_sdram_choose_cmd_request[1]) begin
										main_sdram_choose_cmd_grant <= 1'd1;
									end else begin
										if (main_sdram_choose_cmd_request[2]) begin
											main_sdram_choose_cmd_grant <= 2'd2;
										end
									end
								end
							end
						end
					end
				end
			end
			3'd4: begin
				if (main_sdram_choose_cmd_request[5]) begin
					main_sdram_choose_cmd_grant <= 3'd5;
				end else begin
					if (main_sdram_choose_cmd_request[6]) begin
						main_sdram_choose_cmd_grant <= 3'd6;
					end else begin
						if (main_sdram_choose_cmd_request[7]) begin
							main_sdram_choose_cmd_grant <= 3'd7;
						end else begin
							if (main_sdram_choose_cmd_request[0]) begin
								main_sdram_choose_cmd_grant <= 1'd0;
							end else begin
								if (main_sdram_choose_cmd_request[1]) begin
									main_sdram_choose_cmd_grant <= 1'd1;
								end else begin
									if (main_sdram_choose_cmd_request[2]) begin
										main_sdram_choose_cmd_grant <= 2'd2;
									end else begin
										if (main_sdram_choose_cmd_request[3]) begin
											main_sdram_choose_cmd_grant <= 2'd3;
										end
									end
								end
							end
						end
					end
				end
			end
			3'd5: begin
				if (main_sdram_choose_cmd_request[6]) begin
					main_sdram_choose_cmd_grant <= 3'd6;
				end else begin
					if (main_sdram_choose_cmd_request[7]) begin
						main_sdram_choose_cmd_grant <= 3'd7;
					end else begin
						if (main_sdram_choose_cmd_request[0]) begin
							main_sdram_choose_cmd_grant <= 1'd0;
						end else begin
							if (main_sdram_choose_cmd_request[1]) begin
								main_sdram_choose_cmd_grant <= 1'd1;
							end else begin
								if (main_sdram_choose_cmd_request[2]) begin
									main_sdram_choose_cmd_grant <= 2'd2;
								end else begin
									if (main_sdram_choose_cmd_request[3]) begin
										main_sdram_choose_cmd_grant <= 2'd3;
									end else begin
										if (main_sdram_choose_cmd_request[4]) begin
											main_sdram_choose_cmd_grant <= 3'd4;
										end
									end
								end
							end
						end
					end
				end
			end
			3'd6: begin
				if (main_sdram_choose_cmd_request[7]) begin
					main_sdram_choose_cmd_grant <= 3'd7;
				end else begin
					if (main_sdram_choose_cmd_request[0]) begin
						main_sdram_choose_cmd_grant <= 1'd0;
					end else begin
						if (main_sdram_choose_cmd_request[1]) begin
							main_sdram_choose_cmd_grant <= 1'd1;
						end else begin
							if (main_sdram_choose_cmd_request[2]) begin
								main_sdram_choose_cmd_grant <= 2'd2;
							end else begin
								if (main_sdram_choose_cmd_request[3]) begin
									main_sdram_choose_cmd_grant <= 2'd3;
								end else begin
									if (main_sdram_choose_cmd_request[4]) begin
										main_sdram_choose_cmd_grant <= 3'd4;
									end else begin
										if (main_sdram_choose_cmd_request[5]) begin
											main_sdram_choose_cmd_grant <= 3'd5;
										end
									end
								end
							end
						end
					end
				end
			end
			3'd7: begin
				if (main_sdram_choose_cmd_request[0]) begin
					main_sdram_choose_cmd_grant <= 1'd0;
				end else begin
					if (main_sdram_choose_cmd_request[1]) begin
						main_sdram_choose_cmd_grant <= 1'd1;
					end else begin
						if (main_sdram_choose_cmd_request[2]) begin
							main_sdram_choose_cmd_grant <= 2'd2;
						end else begin
							if (main_sdram_choose_cmd_request[3]) begin
								main_sdram_choose_cmd_grant <= 2'd3;
							end else begin
								if (main_sdram_choose_cmd_request[4]) begin
									main_sdram_choose_cmd_grant <= 3'd4;
								end else begin
									if (main_sdram_choose_cmd_request[5]) begin
										main_sdram_choose_cmd_grant <= 3'd5;
									end else begin
										if (main_sdram_choose_cmd_request[6]) begin
											main_sdram_choose_cmd_grant <= 3'd6;
										end
									end
								end
							end
						end
					end
				end
			end
		endcase
	end
	if (main_sdram_choose_req_ce) begin
		case (main_sdram_choose_req_grant)
			1'd0: begin
				if (main_sdram_choose_req_request[1]) begin
					main_sdram_choose_req_grant <= 1'd1;
				end else begin
					if (main_sdram_choose_req_request[2]) begin
						main_sdram_choose_req_grant <= 2'd2;
					end else begin
						if (main_sdram_choose_req_request[3]) begin
							main_sdram_choose_req_grant <= 2'd3;
						end else begin
							if (main_sdram_choose_req_request[4]) begin
								main_sdram_choose_req_grant <= 3'd4;
							end else begin
								if (main_sdram_choose_req_request[5]) begin
									main_sdram_choose_req_grant <= 3'd5;
								end else begin
									if (main_sdram_choose_req_request[6]) begin
										main_sdram_choose_req_grant <= 3'd6;
									end else begin
										if (main_sdram_choose_req_request[7]) begin
											main_sdram_choose_req_grant <= 3'd7;
										end
									end
								end
							end
						end
					end
				end
			end
			1'd1: begin
				if (main_sdram_choose_req_request[2]) begin
					main_sdram_choose_req_grant <= 2'd2;
				end else begin
					if (main_sdram_choose_req_request[3]) begin
						main_sdram_choose_req_grant <= 2'd3;
					end else begin
						if (main_sdram_choose_req_request[4]) begin
							main_sdram_choose_req_grant <= 3'd4;
						end else begin
							if (main_sdram_choose_req_request[5]) begin
								main_sdram_choose_req_grant <= 3'd5;
							end else begin
								if (main_sdram_choose_req_request[6]) begin
									main_sdram_choose_req_grant <= 3'd6;
								end else begin
									if (main_sdram_choose_req_request[7]) begin
										main_sdram_choose_req_grant <= 3'd7;
									end else begin
										if (main_sdram_choose_req_request[0]) begin
											main_sdram_choose_req_grant <= 1'd0;
										end
									end
								end
							end
						end
					end
				end
			end
			2'd2: begin
				if (main_sdram_choose_req_request[3]) begin
					main_sdram_choose_req_grant <= 2'd3;
				end else begin
					if (main_sdram_choose_req_request[4]) begin
						main_sdram_choose_req_grant <= 3'd4;
					end else begin
						if (main_sdram_choose_req_request[5]) begin
							main_sdram_choose_req_grant <= 3'd5;
						end else begin
							if (main_sdram_choose_req_request[6]) begin
								main_sdram_choose_req_grant <= 3'd6;
							end else begin
								if (main_sdram_choose_req_request[7]) begin
									main_sdram_choose_req_grant <= 3'd7;
								end else begin
									if (main_sdram_choose_req_request[0]) begin
										main_sdram_choose_req_grant <= 1'd0;
									end else begin
										if (main_sdram_choose_req_request[1]) begin
											main_sdram_choose_req_grant <= 1'd1;
										end
									end
								end
							end
						end
					end
				end
			end
			2'd3: begin
				if (main_sdram_choose_req_request[4]) begin
					main_sdram_choose_req_grant <= 3'd4;
				end else begin
					if (main_sdram_choose_req_request[5]) begin
						main_sdram_choose_req_grant <= 3'd5;
					end else begin
						if (main_sdram_choose_req_request[6]) begin
							main_sdram_choose_req_grant <= 3'd6;
						end else begin
							if (main_sdram_choose_req_request[7]) begin
								main_sdram_choose_req_grant <= 3'd7;
							end else begin
								if (main_sdram_choose_req_request[0]) begin
									main_sdram_choose_req_grant <= 1'd0;
								end else begin
									if (main_sdram_choose_req_request[1]) begin
										main_sdram_choose_req_grant <= 1'd1;
									end else begin
										if (main_sdram_choose_req_request[2]) begin
											main_sdram_choose_req_grant <= 2'd2;
										end
									end
								end
							end
						end
					end
				end
			end
			3'd4: begin
				if (main_sdram_choose_req_request[5]) begin
					main_sdram_choose_req_grant <= 3'd5;
				end else begin
					if (main_sdram_choose_req_request[6]) begin
						main_sdram_choose_req_grant <= 3'd6;
					end else begin
						if (main_sdram_choose_req_request[7]) begin
							main_sdram_choose_req_grant <= 3'd7;
						end else begin
							if (main_sdram_choose_req_request[0]) begin
								main_sdram_choose_req_grant <= 1'd0;
							end else begin
								if (main_sdram_choose_req_request[1]) begin
									main_sdram_choose_req_grant <= 1'd1;
								end else begin
									if (main_sdram_choose_req_request[2]) begin
										main_sdram_choose_req_grant <= 2'd2;
									end else begin
										if (main_sdram_choose_req_request[3]) begin
											main_sdram_choose_req_grant <= 2'd3;
										end
									end
								end
							end
						end
					end
				end
			end
			3'd5: begin
				if (main_sdram_choose_req_request[6]) begin
					main_sdram_choose_req_grant <= 3'd6;
				end else begin
					if (main_sdram_choose_req_request[7]) begin
						main_sdram_choose_req_grant <= 3'd7;
					end else begin
						if (main_sdram_choose_req_request[0]) begin
							main_sdram_choose_req_grant <= 1'd0;
						end else begin
							if (main_sdram_choose_req_request[1]) begin
								main_sdram_choose_req_grant <= 1'd1;
							end else begin
								if (main_sdram_choose_req_request[2]) begin
									main_sdram_choose_req_grant <= 2'd2;
								end else begin
									if (main_sdram_choose_req_request[3]) begin
										main_sdram_choose_req_grant <= 2'd3;
									end else begin
										if (main_sdram_choose_req_request[4]) begin
											main_sdram_choose_req_grant <= 3'd4;
										end
									end
								end
							end
						end
					end
				end
			end
			3'd6: begin
				if (main_sdram_choose_req_request[7]) begin
					main_sdram_choose_req_grant <= 3'd7;
				end else begin
					if (main_sdram_choose_req_request[0]) begin
						main_sdram_choose_req_grant <= 1'd0;
					end else begin
						if (main_sdram_choose_req_request[1]) begin
							main_sdram_choose_req_grant <= 1'd1;
						end else begin
							if (main_sdram_choose_req_request[2]) begin
								main_sdram_choose_req_grant <= 2'd2;
							end else begin
								if (main_sdram_choose_req_request[3]) begin
									main_sdram_choose_req_grant <= 2'd3;
								end else begin
									if (main_sdram_choose_req_request[4]) begin
										main_sdram_choose_req_grant <= 3'd4;
									end else begin
										if (main_sdram_choose_req_request[5]) begin
											main_sdram_choose_req_grant <= 3'd5;
										end
									end
								end
							end
						end
					end
				end
			end
			3'd7: begin
				if (main_sdram_choose_req_request[0]) begin
					main_sdram_choose_req_grant <= 1'd0;
				end else begin
					if (main_sdram_choose_req_request[1]) begin
						main_sdram_choose_req_grant <= 1'd1;
					end else begin
						if (main_sdram_choose_req_request[2]) begin
							main_sdram_choose_req_grant <= 2'd2;
						end else begin
							if (main_sdram_choose_req_request[3]) begin
								main_sdram_choose_req_grant <= 2'd3;
							end else begin
								if (main_sdram_choose_req_request[4]) begin
									main_sdram_choose_req_grant <= 3'd4;
								end else begin
									if (main_sdram_choose_req_request[5]) begin
										main_sdram_choose_req_grant <= 3'd5;
									end else begin
										if (main_sdram_choose_req_request[6]) begin
											main_sdram_choose_req_grant <= 3'd6;
										end
									end
								end
							end
						end
					end
				end
			end
		endcase
	end
	main_sdram_dfi_p0_cs_n <= 1'd0;
	main_sdram_dfi_p0_bank <= builder_array_muxed0;
	main_sdram_dfi_p0_address <= builder_array_muxed1;
	main_sdram_dfi_p0_cas_n <= (~builder_array_muxed2);
	main_sdram_dfi_p0_ras_n <= (~builder_array_muxed3);
	main_sdram_dfi_p0_we_n <= (~builder_array_muxed4);
	main_sdram_dfi_p0_rddata_en <= builder_array_muxed5;
	main_sdram_dfi_p0_wrdata_en <= builder_array_muxed6;
	main_sdram_dfi_p1_cs_n <= 1'd0;
	main_sdram_dfi_p1_bank <= builder_array_muxed7;
	main_sdram_dfi_p1_address <= builder_array_muxed8;
	main_sdram_dfi_p1_cas_n <= (~builder_array_muxed9);
	main_sdram_dfi_p1_ras_n <= (~builder_array_muxed10);
	main_sdram_dfi_p1_we_n <= (~builder_array_muxed11);
	main_sdram_dfi_p1_rddata_en <= builder_array_muxed12;
	main_sdram_dfi_p1_wrdata_en <= builder_array_muxed13;
	main_sdram_dfi_p2_cs_n <= 1'd0;
	main_sdram_dfi_p2_bank <= builder_array_muxed14;
	main_sdram_dfi_p2_address <= builder_array_muxed15;
	main_sdram_dfi_p2_cas_n <= (~builder_array_muxed16);
	main_sdram_dfi_p2_ras_n <= (~builder_array_muxed17);
	main_sdram_dfi_p2_we_n <= (~builder_array_muxed18);
	main_sdram_dfi_p2_rddata_en <= builder_array_muxed19;
	main_sdram_dfi_p2_wrdata_en <= builder_array_muxed20;
	main_sdram_dfi_p3_cs_n <= 1'd0;
	main_sdram_dfi_p3_bank <= builder_array_muxed21;
	main_sdram_dfi_p3_address <= builder_array_muxed22;
	main_sdram_dfi_p3_cas_n <= (~builder_array_muxed23);
	main_sdram_dfi_p3_ras_n <= (~builder_array_muxed24);
	main_sdram_dfi_p3_we_n <= (~builder_array_muxed25);
	main_sdram_dfi_p3_rddata_en <= builder_array_muxed26;
	main_sdram_dfi_p3_wrdata_en <= builder_array_muxed27;
	if (main_sdram_trrdcon_valid) begin
		main_sdram_trrdcon_count <= 1'd1;
		if (1'd0) begin
			main_sdram_trrdcon_ready <= 1'd1;
		end else begin
			main_sdram_trrdcon_ready <= 1'd0;
		end
	end else begin
		if ((~main_sdram_trrdcon_ready)) begin
			main_sdram_trrdcon_count <= (main_sdram_trrdcon_count - 1'd1);
			if ((main_sdram_trrdcon_count == 1'd1)) begin
				main_sdram_trrdcon_ready <= 1'd1;
			end
		end
	end
	main_sdram_tfawcon_window <= {main_sdram_tfawcon_window, main_sdram_tfawcon_valid};
	if ((main_sdram_tfawcon_count < 3'd4)) begin
		if ((main_sdram_tfawcon_count == 2'd3)) begin
			main_sdram_tfawcon_ready <= (~main_sdram_tfawcon_valid);
		end else begin
			main_sdram_tfawcon_ready <= 1'd1;
		end
	end
	if (main_sdram_tccdcon_valid) begin
		main_sdram_tccdcon_count <= 1'd0;
		if (1'd1) begin
			main_sdram_tccdcon_ready <= 1'd1;
		end else begin
			main_sdram_tccdcon_ready <= 1'd0;
		end
	end else begin
		if ((~main_sdram_tccdcon_ready)) begin
			main_sdram_tccdcon_count <= (main_sdram_tccdcon_count - 1'd1);
			if ((main_sdram_tccdcon_count == 1'd1)) begin
				main_sdram_tccdcon_ready <= 1'd1;
			end
		end
	end
	if (main_sdram_twtrcon_valid) begin
		main_sdram_twtrcon_count <= 3'd4;
		if (1'd0) begin
			main_sdram_twtrcon_ready <= 1'd1;
		end else begin
			main_sdram_twtrcon_ready <= 1'd0;
		end
	end else begin
		if ((~main_sdram_twtrcon_ready)) begin
			main_sdram_twtrcon_count <= (main_sdram_twtrcon_count - 1'd1);
			if ((main_sdram_twtrcon_count == 1'd1)) begin
				main_sdram_twtrcon_ready <= 1'd1;
			end
		end
	end
	builder_multiplexer_state <= builder_multiplexer_next_state;
	if (((builder_roundrobin0_grant == 1'd0) & main_sdram_interface_bank0_rdata_valid)) begin
		builder_rbank <= 1'd0;
	end
	if (((builder_roundrobin0_grant == 1'd0) & main_sdram_interface_bank0_wdata_ready)) begin
		builder_wbank <= 1'd0;
	end
	if (((builder_roundrobin1_grant == 1'd0) & main_sdram_interface_bank1_rdata_valid)) begin
		builder_rbank <= 1'd1;
	end
	if (((builder_roundrobin1_grant == 1'd0) & main_sdram_interface_bank1_wdata_ready)) begin
		builder_wbank <= 1'd1;
	end
	if (((builder_roundrobin2_grant == 1'd0) & main_sdram_interface_bank2_rdata_valid)) begin
		builder_rbank <= 2'd2;
	end
	if (((builder_roundrobin2_grant == 1'd0) & main_sdram_interface_bank2_wdata_ready)) begin
		builder_wbank <= 2'd2;
	end
	if (((builder_roundrobin3_grant == 1'd0) & main_sdram_interface_bank3_rdata_valid)) begin
		builder_rbank <= 2'd3;
	end
	if (((builder_roundrobin3_grant == 1'd0) & main_sdram_interface_bank3_wdata_ready)) begin
		builder_wbank <= 2'd3;
	end
	if (((builder_roundrobin4_grant == 1'd0) & main_sdram_interface_bank4_rdata_valid)) begin
		builder_rbank <= 3'd4;
	end
	if (((builder_roundrobin4_grant == 1'd0) & main_sdram_interface_bank4_wdata_ready)) begin
		builder_wbank <= 3'd4;
	end
	if (((builder_roundrobin5_grant == 1'd0) & main_sdram_interface_bank5_rdata_valid)) begin
		builder_rbank <= 3'd5;
	end
	if (((builder_roundrobin5_grant == 1'd0) & main_sdram_interface_bank5_wdata_ready)) begin
		builder_wbank <= 3'd5;
	end
	if (((builder_roundrobin6_grant == 1'd0) & main_sdram_interface_bank6_rdata_valid)) begin
		builder_rbank <= 3'd6;
	end
	if (((builder_roundrobin6_grant == 1'd0) & main_sdram_interface_bank6_wdata_ready)) begin
		builder_wbank <= 3'd6;
	end
	if (((builder_roundrobin7_grant == 1'd0) & main_sdram_interface_bank7_rdata_valid)) begin
		builder_rbank <= 3'd7;
	end
	if (((builder_roundrobin7_grant == 1'd0) & main_sdram_interface_bank7_wdata_ready)) begin
		builder_wbank <= 3'd7;
	end
	builder_new_master_wdata_ready0 <= ((((((((1'd0 | ((builder_roundrobin0_grant == 1'd0) & main_sdram_interface_bank0_wdata_ready)) | ((builder_roundrobin1_grant == 1'd0) & main_sdram_interface_bank1_wdata_ready)) | ((builder_roundrobin2_grant == 1'd0) & main_sdram_interface_bank2_wdata_ready)) | ((builder_roundrobin3_grant == 1'd0) & main_sdram_interface_bank3_wdata_ready)) | ((builder_roundrobin4_grant == 1'd0) & main_sdram_interface_bank4_wdata_ready)) | ((builder_roundrobin5_grant == 1'd0) & main_sdram_interface_bank5_wdata_ready)) | ((builder_roundrobin6_grant == 1'd0) & main_sdram_interface_bank6_wdata_ready)) | ((builder_roundrobin7_grant == 1'd0) & main_sdram_interface_bank7_wdata_ready));
	builder_new_master_wdata_ready1 <= builder_new_master_wdata_ready0;
	builder_new_master_wdata_ready2 <= builder_new_master_wdata_ready1;
	builder_new_master_rdata_valid0 <= ((((((((1'd0 | ((builder_roundrobin0_grant == 1'd0) & main_sdram_interface_bank0_rdata_valid)) | ((builder_roundrobin1_grant == 1'd0) & main_sdram_interface_bank1_rdata_valid)) | ((builder_roundrobin2_grant == 1'd0) & main_sdram_interface_bank2_rdata_valid)) | ((builder_roundrobin3_grant == 1'd0) & main_sdram_interface_bank3_rdata_valid)) | ((builder_roundrobin4_grant == 1'd0) & main_sdram_interface_bank4_rdata_valid)) | ((builder_roundrobin5_grant == 1'd0) & main_sdram_interface_bank5_rdata_valid)) | ((builder_roundrobin6_grant == 1'd0) & main_sdram_interface_bank6_rdata_valid)) | ((builder_roundrobin7_grant == 1'd0) & main_sdram_interface_bank7_rdata_valid));
	builder_new_master_rdata_valid1 <= builder_new_master_rdata_valid0;
	builder_new_master_rdata_valid2 <= builder_new_master_rdata_valid1;
	builder_new_master_rdata_valid3 <= builder_new_master_rdata_valid2;
	builder_new_master_rdata_valid4 <= builder_new_master_rdata_valid3;
	builder_new_master_rdata_valid5 <= builder_new_master_rdata_valid4;
	builder_new_master_rdata_valid6 <= builder_new_master_rdata_valid5;
	builder_new_master_rdata_valid7 <= builder_new_master_rdata_valid6;
	builder_new_master_rdata_valid8 <= builder_new_master_rdata_valid7;
	builder_new_master_rdata_valid9 <= builder_new_master_rdata_valid8;
	main_adr_offset_r <= main_interface0_wb_sdram_adr[1:0];
	builder_fullmemorywe_state <= builder_fullmemorywe_next_state;
	builder_litedramwishbone2native_state <= builder_litedramwishbone2native_next_state;
	if (main_count_next_value_ce) begin
		main_count <= main_count_next_value;
	end
	builder_basesoc_slave_sel_r <= builder_basesoc_slave_sel;
	if (builder_basesoc_wait) begin
		if ((~builder_basesoc_done)) begin
			builder_basesoc_count <= (builder_basesoc_count - 1'd1);
		end
	end else begin
		builder_basesoc_count <= 20'd1000000;
	end
	builder_basesoc_csrbankarray_interface0_bank_bus_dat_r <= 1'd0;
	if (builder_basesoc_csrbankarray_csrbank0_sel) begin
		case (builder_basesoc_csrbankarray_interface0_bank_bus_adr[3:0])
			1'd0: begin
				builder_basesoc_csrbankarray_interface0_bank_bus_dat_r <= builder_basesoc_csrbankarray_csrbank0_reset0_w;
			end
			1'd1: begin
				builder_basesoc_csrbankarray_interface0_bank_bus_dat_r <= builder_basesoc_csrbankarray_csrbank0_scratch3_w;
			end
			2'd2: begin
				builder_basesoc_csrbankarray_interface0_bank_bus_dat_r <= builder_basesoc_csrbankarray_csrbank0_scratch2_w;
			end
			2'd3: begin
				builder_basesoc_csrbankarray_interface0_bank_bus_dat_r <= builder_basesoc_csrbankarray_csrbank0_scratch1_w;
			end
			3'd4: begin
				builder_basesoc_csrbankarray_interface0_bank_bus_dat_r <= builder_basesoc_csrbankarray_csrbank0_scratch0_w;
			end
			3'd5: begin
				builder_basesoc_csrbankarray_interface0_bank_bus_dat_r <= builder_basesoc_csrbankarray_csrbank0_bus_errors3_w;
			end
			3'd6: begin
				builder_basesoc_csrbankarray_interface0_bank_bus_dat_r <= builder_basesoc_csrbankarray_csrbank0_bus_errors2_w;
			end
			3'd7: begin
				builder_basesoc_csrbankarray_interface0_bank_bus_dat_r <= builder_basesoc_csrbankarray_csrbank0_bus_errors1_w;
			end
			4'd8: begin
				builder_basesoc_csrbankarray_interface0_bank_bus_dat_r <= builder_basesoc_csrbankarray_csrbank0_bus_errors0_w;
			end
		endcase
	end
	if (builder_basesoc_csrbankarray_csrbank0_reset0_re) begin
		main_ctrl_reset_storage <= builder_basesoc_csrbankarray_csrbank0_reset0_r;
	end
	main_ctrl_reset_re <= builder_basesoc_csrbankarray_csrbank0_reset0_re;
	if (builder_basesoc_csrbankarray_csrbank0_scratch3_re) begin
		main_ctrl_scratch_storage[31:24] <= builder_basesoc_csrbankarray_csrbank0_scratch3_r;
	end
	if (builder_basesoc_csrbankarray_csrbank0_scratch2_re) begin
		main_ctrl_scratch_storage[23:16] <= builder_basesoc_csrbankarray_csrbank0_scratch2_r;
	end
	if (builder_basesoc_csrbankarray_csrbank0_scratch1_re) begin
		main_ctrl_scratch_storage[15:8] <= builder_basesoc_csrbankarray_csrbank0_scratch1_r;
	end
	if (builder_basesoc_csrbankarray_csrbank0_scratch0_re) begin
		main_ctrl_scratch_storage[7:0] <= builder_basesoc_csrbankarray_csrbank0_scratch0_r;
	end
	main_ctrl_scratch_re <= builder_basesoc_csrbankarray_csrbank0_scratch0_re;
	builder_basesoc_csrbankarray_interface1_bank_bus_dat_r <= 1'd0;
	if (builder_basesoc_csrbankarray_csrbank1_sel) begin
		case (builder_basesoc_csrbankarray_interface1_bank_bus_adr[2:0])
			1'd0: begin
				builder_basesoc_csrbankarray_interface1_bank_bus_dat_r <= builder_basesoc_csrbankarray_csrbank1_half_sys8x_taps0_w;
			end
			1'd1: begin
				builder_basesoc_csrbankarray_interface1_bank_bus_dat_r <= main_a7ddrphy_cdly_rst_w;
			end
			2'd2: begin
				builder_basesoc_csrbankarray_interface1_bank_bus_dat_r <= main_a7ddrphy_cdly_inc_w;
			end
			2'd3: begin
				builder_basesoc_csrbankarray_interface1_bank_bus_dat_r <= builder_basesoc_csrbankarray_csrbank1_dly_sel0_w;
			end
			3'd4: begin
				builder_basesoc_csrbankarray_interface1_bank_bus_dat_r <= main_a7ddrphy_rdly_dq_rst_w;
			end
			3'd5: begin
				builder_basesoc_csrbankarray_interface1_bank_bus_dat_r <= main_a7ddrphy_rdly_dq_inc_w;
			end
			3'd6: begin
				builder_basesoc_csrbankarray_interface1_bank_bus_dat_r <= main_a7ddrphy_rdly_dq_bitslip_rst_w;
			end
			3'd7: begin
				builder_basesoc_csrbankarray_interface1_bank_bus_dat_r <= main_a7ddrphy_rdly_dq_bitslip_w;
			end
		endcase
	end
	if (builder_basesoc_csrbankarray_csrbank1_half_sys8x_taps0_re) begin
		main_a7ddrphy_half_sys8x_taps_storage[4:0] <= builder_basesoc_csrbankarray_csrbank1_half_sys8x_taps0_r;
	end
	main_a7ddrphy_half_sys8x_taps_re <= builder_basesoc_csrbankarray_csrbank1_half_sys8x_taps0_re;
	if (builder_basesoc_csrbankarray_csrbank1_dly_sel0_re) begin
		main_a7ddrphy_dly_sel_storage[1:0] <= builder_basesoc_csrbankarray_csrbank1_dly_sel0_r;
	end
	main_a7ddrphy_dly_sel_re <= builder_basesoc_csrbankarray_csrbank1_dly_sel0_re;
	builder_basesoc_csrbankarray_sel_r <= builder_basesoc_csrbankarray_sel;
	builder_basesoc_csrbankarray_interface2_bank_bus_dat_r <= 1'd0;
	if (builder_basesoc_csrbankarray_csrbank2_sel) begin
		case (builder_basesoc_csrbankarray_interface2_bank_bus_adr[5:0])
			1'd0: begin
				builder_basesoc_csrbankarray_interface2_bank_bus_dat_r <= builder_basesoc_csrbankarray_csrbank2_dfii_control0_w;
			end
			1'd1: begin
				builder_basesoc_csrbankarray_interface2_bank_bus_dat_r <= builder_basesoc_csrbankarray_csrbank2_dfii_pi0_command0_w;
			end
			2'd2: begin
				builder_basesoc_csrbankarray_interface2_bank_bus_dat_r <= main_sdram_phaseinjector0_command_issue_w;
			end
			2'd3: begin
				builder_basesoc_csrbankarray_interface2_bank_bus_dat_r <= builder_basesoc_csrbankarray_csrbank2_dfii_pi0_address1_w;
			end
			3'd4: begin
				builder_basesoc_csrbankarray_interface2_bank_bus_dat_r <= builder_basesoc_csrbankarray_csrbank2_dfii_pi0_address0_w;
			end
			3'd5: begin
				builder_basesoc_csrbankarray_interface2_bank_bus_dat_r <= builder_basesoc_csrbankarray_csrbank2_dfii_pi0_baddress0_w;
			end
			3'd6: begin
				builder_basesoc_csrbankarray_interface2_bank_bus_dat_r <= builder_basesoc_csrbankarray_csrbank2_dfii_pi0_wrdata3_w;
			end
			3'd7: begin
				builder_basesoc_csrbankarray_interface2_bank_bus_dat_r <= builder_basesoc_csrbankarray_csrbank2_dfii_pi0_wrdata2_w;
			end
			4'd8: begin
				builder_basesoc_csrbankarray_interface2_bank_bus_dat_r <= builder_basesoc_csrbankarray_csrbank2_dfii_pi0_wrdata1_w;
			end
			4'd9: begin
				builder_basesoc_csrbankarray_interface2_bank_bus_dat_r <= builder_basesoc_csrbankarray_csrbank2_dfii_pi0_wrdata0_w;
			end
			4'd10: begin
				builder_basesoc_csrbankarray_interface2_bank_bus_dat_r <= builder_basesoc_csrbankarray_csrbank2_dfii_pi0_rddata3_w;
			end
			4'd11: begin
				builder_basesoc_csrbankarray_interface2_bank_bus_dat_r <= builder_basesoc_csrbankarray_csrbank2_dfii_pi0_rddata2_w;
			end
			4'd12: begin
				builder_basesoc_csrbankarray_interface2_bank_bus_dat_r <= builder_basesoc_csrbankarray_csrbank2_dfii_pi0_rddata1_w;
			end
			4'd13: begin
				builder_basesoc_csrbankarray_interface2_bank_bus_dat_r <= builder_basesoc_csrbankarray_csrbank2_dfii_pi0_rddata0_w;
			end
			4'd14: begin
				builder_basesoc_csrbankarray_interface2_bank_bus_dat_r <= builder_basesoc_csrbankarray_csrbank2_dfii_pi1_command0_w;
			end
			4'd15: begin
				builder_basesoc_csrbankarray_interface2_bank_bus_dat_r <= main_sdram_phaseinjector1_command_issue_w;
			end
			5'd16: begin
				builder_basesoc_csrbankarray_interface2_bank_bus_dat_r <= builder_basesoc_csrbankarray_csrbank2_dfii_pi1_address1_w;
			end
			5'd17: begin
				builder_basesoc_csrbankarray_interface2_bank_bus_dat_r <= builder_basesoc_csrbankarray_csrbank2_dfii_pi1_address0_w;
			end
			5'd18: begin
				builder_basesoc_csrbankarray_interface2_bank_bus_dat_r <= builder_basesoc_csrbankarray_csrbank2_dfii_pi1_baddress0_w;
			end
			5'd19: begin
				builder_basesoc_csrbankarray_interface2_bank_bus_dat_r <= builder_basesoc_csrbankarray_csrbank2_dfii_pi1_wrdata3_w;
			end
			5'd20: begin
				builder_basesoc_csrbankarray_interface2_bank_bus_dat_r <= builder_basesoc_csrbankarray_csrbank2_dfii_pi1_wrdata2_w;
			end
			5'd21: begin
				builder_basesoc_csrbankarray_interface2_bank_bus_dat_r <= builder_basesoc_csrbankarray_csrbank2_dfii_pi1_wrdata1_w;
			end
			5'd22: begin
				builder_basesoc_csrbankarray_interface2_bank_bus_dat_r <= builder_basesoc_csrbankarray_csrbank2_dfii_pi1_wrdata0_w;
			end
			5'd23: begin
				builder_basesoc_csrbankarray_interface2_bank_bus_dat_r <= builder_basesoc_csrbankarray_csrbank2_dfii_pi1_rddata3_w;
			end
			5'd24: begin
				builder_basesoc_csrbankarray_interface2_bank_bus_dat_r <= builder_basesoc_csrbankarray_csrbank2_dfii_pi1_rddata2_w;
			end
			5'd25: begin
				builder_basesoc_csrbankarray_interface2_bank_bus_dat_r <= builder_basesoc_csrbankarray_csrbank2_dfii_pi1_rddata1_w;
			end
			5'd26: begin
				builder_basesoc_csrbankarray_interface2_bank_bus_dat_r <= builder_basesoc_csrbankarray_csrbank2_dfii_pi1_rddata0_w;
			end
			5'd27: begin
				builder_basesoc_csrbankarray_interface2_bank_bus_dat_r <= builder_basesoc_csrbankarray_csrbank2_dfii_pi2_command0_w;
			end
			5'd28: begin
				builder_basesoc_csrbankarray_interface2_bank_bus_dat_r <= main_sdram_phaseinjector2_command_issue_w;
			end
			5'd29: begin
				builder_basesoc_csrbankarray_interface2_bank_bus_dat_r <= builder_basesoc_csrbankarray_csrbank2_dfii_pi2_address1_w;
			end
			5'd30: begin
				builder_basesoc_csrbankarray_interface2_bank_bus_dat_r <= builder_basesoc_csrbankarray_csrbank2_dfii_pi2_address0_w;
			end
			5'd31: begin
				builder_basesoc_csrbankarray_interface2_bank_bus_dat_r <= builder_basesoc_csrbankarray_csrbank2_dfii_pi2_baddress0_w;
			end
			6'd32: begin
				builder_basesoc_csrbankarray_interface2_bank_bus_dat_r <= builder_basesoc_csrbankarray_csrbank2_dfii_pi2_wrdata3_w;
			end
			6'd33: begin
				builder_basesoc_csrbankarray_interface2_bank_bus_dat_r <= builder_basesoc_csrbankarray_csrbank2_dfii_pi2_wrdata2_w;
			end
			6'd34: begin
				builder_basesoc_csrbankarray_interface2_bank_bus_dat_r <= builder_basesoc_csrbankarray_csrbank2_dfii_pi2_wrdata1_w;
			end
			6'd35: begin
				builder_basesoc_csrbankarray_interface2_bank_bus_dat_r <= builder_basesoc_csrbankarray_csrbank2_dfii_pi2_wrdata0_w;
			end
			6'd36: begin
				builder_basesoc_csrbankarray_interface2_bank_bus_dat_r <= builder_basesoc_csrbankarray_csrbank2_dfii_pi2_rddata3_w;
			end
			6'd37: begin
				builder_basesoc_csrbankarray_interface2_bank_bus_dat_r <= builder_basesoc_csrbankarray_csrbank2_dfii_pi2_rddata2_w;
			end
			6'd38: begin
				builder_basesoc_csrbankarray_interface2_bank_bus_dat_r <= builder_basesoc_csrbankarray_csrbank2_dfii_pi2_rddata1_w;
			end
			6'd39: begin
				builder_basesoc_csrbankarray_interface2_bank_bus_dat_r <= builder_basesoc_csrbankarray_csrbank2_dfii_pi2_rddata0_w;
			end
			6'd40: begin
				builder_basesoc_csrbankarray_interface2_bank_bus_dat_r <= builder_basesoc_csrbankarray_csrbank2_dfii_pi3_command0_w;
			end
			6'd41: begin
				builder_basesoc_csrbankarray_interface2_bank_bus_dat_r <= main_sdram_phaseinjector3_command_issue_w;
			end
			6'd42: begin
				builder_basesoc_csrbankarray_interface2_bank_bus_dat_r <= builder_basesoc_csrbankarray_csrbank2_dfii_pi3_address1_w;
			end
			6'd43: begin
				builder_basesoc_csrbankarray_interface2_bank_bus_dat_r <= builder_basesoc_csrbankarray_csrbank2_dfii_pi3_address0_w;
			end
			6'd44: begin
				builder_basesoc_csrbankarray_interface2_bank_bus_dat_r <= builder_basesoc_csrbankarray_csrbank2_dfii_pi3_baddress0_w;
			end
			6'd45: begin
				builder_basesoc_csrbankarray_interface2_bank_bus_dat_r <= builder_basesoc_csrbankarray_csrbank2_dfii_pi3_wrdata3_w;
			end
			6'd46: begin
				builder_basesoc_csrbankarray_interface2_bank_bus_dat_r <= builder_basesoc_csrbankarray_csrbank2_dfii_pi3_wrdata2_w;
			end
			6'd47: begin
				builder_basesoc_csrbankarray_interface2_bank_bus_dat_r <= builder_basesoc_csrbankarray_csrbank2_dfii_pi3_wrdata1_w;
			end
			6'd48: begin
				builder_basesoc_csrbankarray_interface2_bank_bus_dat_r <= builder_basesoc_csrbankarray_csrbank2_dfii_pi3_wrdata0_w;
			end
			6'd49: begin
				builder_basesoc_csrbankarray_interface2_bank_bus_dat_r <= builder_basesoc_csrbankarray_csrbank2_dfii_pi3_rddata3_w;
			end
			6'd50: begin
				builder_basesoc_csrbankarray_interface2_bank_bus_dat_r <= builder_basesoc_csrbankarray_csrbank2_dfii_pi3_rddata2_w;
			end
			6'd51: begin
				builder_basesoc_csrbankarray_interface2_bank_bus_dat_r <= builder_basesoc_csrbankarray_csrbank2_dfii_pi3_rddata1_w;
			end
			6'd52: begin
				builder_basesoc_csrbankarray_interface2_bank_bus_dat_r <= builder_basesoc_csrbankarray_csrbank2_dfii_pi3_rddata0_w;
			end
		endcase
	end
	if (builder_basesoc_csrbankarray_csrbank2_dfii_control0_re) begin
		main_sdram_storage[3:0] <= builder_basesoc_csrbankarray_csrbank2_dfii_control0_r;
	end
	main_sdram_re <= builder_basesoc_csrbankarray_csrbank2_dfii_control0_re;
	if (builder_basesoc_csrbankarray_csrbank2_dfii_pi0_command0_re) begin
		main_sdram_phaseinjector0_command_storage[5:0] <= builder_basesoc_csrbankarray_csrbank2_dfii_pi0_command0_r;
	end
	main_sdram_phaseinjector0_command_re <= builder_basesoc_csrbankarray_csrbank2_dfii_pi0_command0_re;
	if (builder_basesoc_csrbankarray_csrbank2_dfii_pi0_address1_re) begin
		main_sdram_phaseinjector0_address_storage[13:8] <= builder_basesoc_csrbankarray_csrbank2_dfii_pi0_address1_r;
	end
	if (builder_basesoc_csrbankarray_csrbank2_dfii_pi0_address0_re) begin
		main_sdram_phaseinjector0_address_storage[7:0] <= builder_basesoc_csrbankarray_csrbank2_dfii_pi0_address0_r;
	end
	main_sdram_phaseinjector0_address_re <= builder_basesoc_csrbankarray_csrbank2_dfii_pi0_address0_re;
	if (builder_basesoc_csrbankarray_csrbank2_dfii_pi0_baddress0_re) begin
		main_sdram_phaseinjector0_baddress_storage[2:0] <= builder_basesoc_csrbankarray_csrbank2_dfii_pi0_baddress0_r;
	end
	main_sdram_phaseinjector0_baddress_re <= builder_basesoc_csrbankarray_csrbank2_dfii_pi0_baddress0_re;
	if (builder_basesoc_csrbankarray_csrbank2_dfii_pi0_wrdata3_re) begin
		main_sdram_phaseinjector0_wrdata_storage[31:24] <= builder_basesoc_csrbankarray_csrbank2_dfii_pi0_wrdata3_r;
	end
	if (builder_basesoc_csrbankarray_csrbank2_dfii_pi0_wrdata2_re) begin
		main_sdram_phaseinjector0_wrdata_storage[23:16] <= builder_basesoc_csrbankarray_csrbank2_dfii_pi0_wrdata2_r;
	end
	if (builder_basesoc_csrbankarray_csrbank2_dfii_pi0_wrdata1_re) begin
		main_sdram_phaseinjector0_wrdata_storage[15:8] <= builder_basesoc_csrbankarray_csrbank2_dfii_pi0_wrdata1_r;
	end
	if (builder_basesoc_csrbankarray_csrbank2_dfii_pi0_wrdata0_re) begin
		main_sdram_phaseinjector0_wrdata_storage[7:0] <= builder_basesoc_csrbankarray_csrbank2_dfii_pi0_wrdata0_r;
	end
	main_sdram_phaseinjector0_wrdata_re <= builder_basesoc_csrbankarray_csrbank2_dfii_pi0_wrdata0_re;
	if (builder_basesoc_csrbankarray_csrbank2_dfii_pi1_command0_re) begin
		main_sdram_phaseinjector1_command_storage[5:0] <= builder_basesoc_csrbankarray_csrbank2_dfii_pi1_command0_r;
	end
	main_sdram_phaseinjector1_command_re <= builder_basesoc_csrbankarray_csrbank2_dfii_pi1_command0_re;
	if (builder_basesoc_csrbankarray_csrbank2_dfii_pi1_address1_re) begin
		main_sdram_phaseinjector1_address_storage[13:8] <= builder_basesoc_csrbankarray_csrbank2_dfii_pi1_address1_r;
	end
	if (builder_basesoc_csrbankarray_csrbank2_dfii_pi1_address0_re) begin
		main_sdram_phaseinjector1_address_storage[7:0] <= builder_basesoc_csrbankarray_csrbank2_dfii_pi1_address0_r;
	end
	main_sdram_phaseinjector1_address_re <= builder_basesoc_csrbankarray_csrbank2_dfii_pi1_address0_re;
	if (builder_basesoc_csrbankarray_csrbank2_dfii_pi1_baddress0_re) begin
		main_sdram_phaseinjector1_baddress_storage[2:0] <= builder_basesoc_csrbankarray_csrbank2_dfii_pi1_baddress0_r;
	end
	main_sdram_phaseinjector1_baddress_re <= builder_basesoc_csrbankarray_csrbank2_dfii_pi1_baddress0_re;
	if (builder_basesoc_csrbankarray_csrbank2_dfii_pi1_wrdata3_re) begin
		main_sdram_phaseinjector1_wrdata_storage[31:24] <= builder_basesoc_csrbankarray_csrbank2_dfii_pi1_wrdata3_r;
	end
	if (builder_basesoc_csrbankarray_csrbank2_dfii_pi1_wrdata2_re) begin
		main_sdram_phaseinjector1_wrdata_storage[23:16] <= builder_basesoc_csrbankarray_csrbank2_dfii_pi1_wrdata2_r;
	end
	if (builder_basesoc_csrbankarray_csrbank2_dfii_pi1_wrdata1_re) begin
		main_sdram_phaseinjector1_wrdata_storage[15:8] <= builder_basesoc_csrbankarray_csrbank2_dfii_pi1_wrdata1_r;
	end
	if (builder_basesoc_csrbankarray_csrbank2_dfii_pi1_wrdata0_re) begin
		main_sdram_phaseinjector1_wrdata_storage[7:0] <= builder_basesoc_csrbankarray_csrbank2_dfii_pi1_wrdata0_r;
	end
	main_sdram_phaseinjector1_wrdata_re <= builder_basesoc_csrbankarray_csrbank2_dfii_pi1_wrdata0_re;
	if (builder_basesoc_csrbankarray_csrbank2_dfii_pi2_command0_re) begin
		main_sdram_phaseinjector2_command_storage[5:0] <= builder_basesoc_csrbankarray_csrbank2_dfii_pi2_command0_r;
	end
	main_sdram_phaseinjector2_command_re <= builder_basesoc_csrbankarray_csrbank2_dfii_pi2_command0_re;
	if (builder_basesoc_csrbankarray_csrbank2_dfii_pi2_address1_re) begin
		main_sdram_phaseinjector2_address_storage[13:8] <= builder_basesoc_csrbankarray_csrbank2_dfii_pi2_address1_r;
	end
	if (builder_basesoc_csrbankarray_csrbank2_dfii_pi2_address0_re) begin
		main_sdram_phaseinjector2_address_storage[7:0] <= builder_basesoc_csrbankarray_csrbank2_dfii_pi2_address0_r;
	end
	main_sdram_phaseinjector2_address_re <= builder_basesoc_csrbankarray_csrbank2_dfii_pi2_address0_re;
	if (builder_basesoc_csrbankarray_csrbank2_dfii_pi2_baddress0_re) begin
		main_sdram_phaseinjector2_baddress_storage[2:0] <= builder_basesoc_csrbankarray_csrbank2_dfii_pi2_baddress0_r;
	end
	main_sdram_phaseinjector2_baddress_re <= builder_basesoc_csrbankarray_csrbank2_dfii_pi2_baddress0_re;
	if (builder_basesoc_csrbankarray_csrbank2_dfii_pi2_wrdata3_re) begin
		main_sdram_phaseinjector2_wrdata_storage[31:24] <= builder_basesoc_csrbankarray_csrbank2_dfii_pi2_wrdata3_r;
	end
	if (builder_basesoc_csrbankarray_csrbank2_dfii_pi2_wrdata2_re) begin
		main_sdram_phaseinjector2_wrdata_storage[23:16] <= builder_basesoc_csrbankarray_csrbank2_dfii_pi2_wrdata2_r;
	end
	if (builder_basesoc_csrbankarray_csrbank2_dfii_pi2_wrdata1_re) begin
		main_sdram_phaseinjector2_wrdata_storage[15:8] <= builder_basesoc_csrbankarray_csrbank2_dfii_pi2_wrdata1_r;
	end
	if (builder_basesoc_csrbankarray_csrbank2_dfii_pi2_wrdata0_re) begin
		main_sdram_phaseinjector2_wrdata_storage[7:0] <= builder_basesoc_csrbankarray_csrbank2_dfii_pi2_wrdata0_r;
	end
	main_sdram_phaseinjector2_wrdata_re <= builder_basesoc_csrbankarray_csrbank2_dfii_pi2_wrdata0_re;
	if (builder_basesoc_csrbankarray_csrbank2_dfii_pi3_command0_re) begin
		main_sdram_phaseinjector3_command_storage[5:0] <= builder_basesoc_csrbankarray_csrbank2_dfii_pi3_command0_r;
	end
	main_sdram_phaseinjector3_command_re <= builder_basesoc_csrbankarray_csrbank2_dfii_pi3_command0_re;
	if (builder_basesoc_csrbankarray_csrbank2_dfii_pi3_address1_re) begin
		main_sdram_phaseinjector3_address_storage[13:8] <= builder_basesoc_csrbankarray_csrbank2_dfii_pi3_address1_r;
	end
	if (builder_basesoc_csrbankarray_csrbank2_dfii_pi3_address0_re) begin
		main_sdram_phaseinjector3_address_storage[7:0] <= builder_basesoc_csrbankarray_csrbank2_dfii_pi3_address0_r;
	end
	main_sdram_phaseinjector3_address_re <= builder_basesoc_csrbankarray_csrbank2_dfii_pi3_address0_re;
	if (builder_basesoc_csrbankarray_csrbank2_dfii_pi3_baddress0_re) begin
		main_sdram_phaseinjector3_baddress_storage[2:0] <= builder_basesoc_csrbankarray_csrbank2_dfii_pi3_baddress0_r;
	end
	main_sdram_phaseinjector3_baddress_re <= builder_basesoc_csrbankarray_csrbank2_dfii_pi3_baddress0_re;
	if (builder_basesoc_csrbankarray_csrbank2_dfii_pi3_wrdata3_re) begin
		main_sdram_phaseinjector3_wrdata_storage[31:24] <= builder_basesoc_csrbankarray_csrbank2_dfii_pi3_wrdata3_r;
	end
	if (builder_basesoc_csrbankarray_csrbank2_dfii_pi3_wrdata2_re) begin
		main_sdram_phaseinjector3_wrdata_storage[23:16] <= builder_basesoc_csrbankarray_csrbank2_dfii_pi3_wrdata2_r;
	end
	if (builder_basesoc_csrbankarray_csrbank2_dfii_pi3_wrdata1_re) begin
		main_sdram_phaseinjector3_wrdata_storage[15:8] <= builder_basesoc_csrbankarray_csrbank2_dfii_pi3_wrdata1_r;
	end
	if (builder_basesoc_csrbankarray_csrbank2_dfii_pi3_wrdata0_re) begin
		main_sdram_phaseinjector3_wrdata_storage[7:0] <= builder_basesoc_csrbankarray_csrbank2_dfii_pi3_wrdata0_r;
	end
	main_sdram_phaseinjector3_wrdata_re <= builder_basesoc_csrbankarray_csrbank2_dfii_pi3_wrdata0_re;
	builder_basesoc_csrbankarray_interface3_bank_bus_dat_r <= 1'd0;
	if (builder_basesoc_csrbankarray_csrbank3_sel) begin
		case (builder_basesoc_csrbankarray_interface3_bank_bus_adr[4:0])
			1'd0: begin
				builder_basesoc_csrbankarray_interface3_bank_bus_dat_r <= builder_basesoc_csrbankarray_csrbank3_load3_w;
			end
			1'd1: begin
				builder_basesoc_csrbankarray_interface3_bank_bus_dat_r <= builder_basesoc_csrbankarray_csrbank3_load2_w;
			end
			2'd2: begin
				builder_basesoc_csrbankarray_interface3_bank_bus_dat_r <= builder_basesoc_csrbankarray_csrbank3_load1_w;
			end
			2'd3: begin
				builder_basesoc_csrbankarray_interface3_bank_bus_dat_r <= builder_basesoc_csrbankarray_csrbank3_load0_w;
			end
			3'd4: begin
				builder_basesoc_csrbankarray_interface3_bank_bus_dat_r <= builder_basesoc_csrbankarray_csrbank3_reload3_w;
			end
			3'd5: begin
				builder_basesoc_csrbankarray_interface3_bank_bus_dat_r <= builder_basesoc_csrbankarray_csrbank3_reload2_w;
			end
			3'd6: begin
				builder_basesoc_csrbankarray_interface3_bank_bus_dat_r <= builder_basesoc_csrbankarray_csrbank3_reload1_w;
			end
			3'd7: begin
				builder_basesoc_csrbankarray_interface3_bank_bus_dat_r <= builder_basesoc_csrbankarray_csrbank3_reload0_w;
			end
			4'd8: begin
				builder_basesoc_csrbankarray_interface3_bank_bus_dat_r <= builder_basesoc_csrbankarray_csrbank3_en0_w;
			end
			4'd9: begin
				builder_basesoc_csrbankarray_interface3_bank_bus_dat_r <= builder_basesoc_csrbankarray_csrbank3_update_value0_w;
			end
			4'd10: begin
				builder_basesoc_csrbankarray_interface3_bank_bus_dat_r <= builder_basesoc_csrbankarray_csrbank3_value3_w;
			end
			4'd11: begin
				builder_basesoc_csrbankarray_interface3_bank_bus_dat_r <= builder_basesoc_csrbankarray_csrbank3_value2_w;
			end
			4'd12: begin
				builder_basesoc_csrbankarray_interface3_bank_bus_dat_r <= builder_basesoc_csrbankarray_csrbank3_value1_w;
			end
			4'd13: begin
				builder_basesoc_csrbankarray_interface3_bank_bus_dat_r <= builder_basesoc_csrbankarray_csrbank3_value0_w;
			end
			4'd14: begin
				builder_basesoc_csrbankarray_interface3_bank_bus_dat_r <= main_eventmanager_status_w;
			end
			4'd15: begin
				builder_basesoc_csrbankarray_interface3_bank_bus_dat_r <= main_eventmanager_pending_w;
			end
			5'd16: begin
				builder_basesoc_csrbankarray_interface3_bank_bus_dat_r <= builder_basesoc_csrbankarray_csrbank3_ev_enable0_w;
			end
		endcase
	end
	if (builder_basesoc_csrbankarray_csrbank3_load3_re) begin
		main_load_storage[31:24] <= builder_basesoc_csrbankarray_csrbank3_load3_r;
	end
	if (builder_basesoc_csrbankarray_csrbank3_load2_re) begin
		main_load_storage[23:16] <= builder_basesoc_csrbankarray_csrbank3_load2_r;
	end
	if (builder_basesoc_csrbankarray_csrbank3_load1_re) begin
		main_load_storage[15:8] <= builder_basesoc_csrbankarray_csrbank3_load1_r;
	end
	if (builder_basesoc_csrbankarray_csrbank3_load0_re) begin
		main_load_storage[7:0] <= builder_basesoc_csrbankarray_csrbank3_load0_r;
	end
	main_load_re <= builder_basesoc_csrbankarray_csrbank3_load0_re;
	if (builder_basesoc_csrbankarray_csrbank3_reload3_re) begin
		main_reload_storage[31:24] <= builder_basesoc_csrbankarray_csrbank3_reload3_r;
	end
	if (builder_basesoc_csrbankarray_csrbank3_reload2_re) begin
		main_reload_storage[23:16] <= builder_basesoc_csrbankarray_csrbank3_reload2_r;
	end
	if (builder_basesoc_csrbankarray_csrbank3_reload1_re) begin
		main_reload_storage[15:8] <= builder_basesoc_csrbankarray_csrbank3_reload1_r;
	end
	if (builder_basesoc_csrbankarray_csrbank3_reload0_re) begin
		main_reload_storage[7:0] <= builder_basesoc_csrbankarray_csrbank3_reload0_r;
	end
	main_reload_re <= builder_basesoc_csrbankarray_csrbank3_reload0_re;
	if (builder_basesoc_csrbankarray_csrbank3_en0_re) begin
		main_en_storage <= builder_basesoc_csrbankarray_csrbank3_en0_r;
	end
	main_en_re <= builder_basesoc_csrbankarray_csrbank3_en0_re;
	if (builder_basesoc_csrbankarray_csrbank3_update_value0_re) begin
		main_update_value_storage <= builder_basesoc_csrbankarray_csrbank3_update_value0_r;
	end
	main_update_value_re <= builder_basesoc_csrbankarray_csrbank3_update_value0_re;
	if (builder_basesoc_csrbankarray_csrbank3_ev_enable0_re) begin
		main_eventmanager_storage <= builder_basesoc_csrbankarray_csrbank3_ev_enable0_r;
	end
	main_eventmanager_re <= builder_basesoc_csrbankarray_csrbank3_ev_enable0_re;
	if (sys_rst) begin
		main_ctrl_reset_storage <= 1'd0;
		main_ctrl_reset_re <= 1'd0;
		main_ctrl_scratch_storage <= 32'd305419896;
		main_ctrl_scratch_re <= 1'd0;
		main_ctrl_bus_errors <= 32'd0;
		main_sram_bus_ack <= 1'd0;
		serial_tx <= 1'd1;
		main_uart_sink_ready <= 1'd0;
		main_uart_uart_clk_txen <= 1'd0;
		main_uart_phase_accumulator_tx <= 32'd0;
		main_uart_tx_reg <= 8'd0;
		main_uart_tx_bitcount <= 4'd0;
		main_uart_tx_busy <= 1'd0;
		main_uart_source_valid <= 1'd0;
		main_uart_source_payload_data <= 8'd0;
		main_uart_uart_clk_rxen <= 1'd0;
		main_uart_phase_accumulator_rx <= 32'd0;
		main_uart_rx_r <= 1'd0;
		main_uart_rx_reg <= 8'd0;
		main_uart_rx_bitcount <= 4'd0;
		main_uart_rx_busy <= 1'd0;
		main_uart_count <= 23'd5000000;
		main_load_storage <= 32'd0;
		main_load_re <= 1'd0;
		main_reload_storage <= 32'd0;
		main_reload_re <= 1'd0;
		main_en_storage <= 1'd0;
		main_en_re <= 1'd0;
		main_update_value_storage <= 1'd0;
		main_update_value_re <= 1'd0;
		main_value_status <= 32'd0;
		main_zero_pending <= 1'd0;
		main_zero_old_trigger <= 1'd0;
		main_eventmanager_storage <= 1'd0;
		main_eventmanager_re <= 1'd0;
		main_value <= 32'd0;
		main_a7ddrphy_half_sys8x_taps_storage <= 5'd16;
		main_a7ddrphy_half_sys8x_taps_re <= 1'd0;
		main_a7ddrphy_dly_sel_storage <= 2'd0;
		main_a7ddrphy_dly_sel_re <= 1'd0;
		main_a7ddrphy_dfi_p0_rddata_valid <= 1'd0;
		main_a7ddrphy_dfi_p1_rddata_valid <= 1'd0;
		main_a7ddrphy_dfi_p2_rddata_valid <= 1'd0;
		main_a7ddrphy_dfi_p3_rddata_valid <= 1'd0;
		main_a7ddrphy_oe_dqs <= 1'd0;
		main_a7ddrphy_oe_dq <= 1'd0;
		main_a7ddrphy_bitslip0_o <= 8'd0;
		main_a7ddrphy_bitslip0_value <= 3'd0;
		main_a7ddrphy_bitslip0_r <= 16'd0;
		main_a7ddrphy_bitslip1_o <= 8'd0;
		main_a7ddrphy_bitslip1_value <= 3'd0;
		main_a7ddrphy_bitslip1_r <= 16'd0;
		main_a7ddrphy_bitslip2_o <= 8'd0;
		main_a7ddrphy_bitslip2_value <= 3'd0;
		main_a7ddrphy_bitslip2_r <= 16'd0;
		main_a7ddrphy_bitslip3_o <= 8'd0;
		main_a7ddrphy_bitslip3_value <= 3'd0;
		main_a7ddrphy_bitslip3_r <= 16'd0;
		main_a7ddrphy_bitslip4_o <= 8'd0;
		main_a7ddrphy_bitslip4_value <= 3'd0;
		main_a7ddrphy_bitslip4_r <= 16'd0;
		main_a7ddrphy_bitslip5_o <= 8'd0;
		main_a7ddrphy_bitslip5_value <= 3'd0;
		main_a7ddrphy_bitslip5_r <= 16'd0;
		main_a7ddrphy_bitslip6_o <= 8'd0;
		main_a7ddrphy_bitslip6_value <= 3'd0;
		main_a7ddrphy_bitslip6_r <= 16'd0;
		main_a7ddrphy_bitslip7_o <= 8'd0;
		main_a7ddrphy_bitslip7_value <= 3'd0;
		main_a7ddrphy_bitslip7_r <= 16'd0;
		main_a7ddrphy_bitslip8_o <= 8'd0;
		main_a7ddrphy_bitslip8_value <= 3'd0;
		main_a7ddrphy_bitslip8_r <= 16'd0;
		main_a7ddrphy_bitslip9_o <= 8'd0;
		main_a7ddrphy_bitslip9_value <= 3'd0;
		main_a7ddrphy_bitslip9_r <= 16'd0;
		main_a7ddrphy_bitslip10_o <= 8'd0;
		main_a7ddrphy_bitslip10_value <= 3'd0;
		main_a7ddrphy_bitslip10_r <= 16'd0;
		main_a7ddrphy_bitslip11_o <= 8'd0;
		main_a7ddrphy_bitslip11_value <= 3'd0;
		main_a7ddrphy_bitslip11_r <= 16'd0;
		main_a7ddrphy_bitslip12_o <= 8'd0;
		main_a7ddrphy_bitslip12_value <= 3'd0;
		main_a7ddrphy_bitslip12_r <= 16'd0;
		main_a7ddrphy_bitslip13_o <= 8'd0;
		main_a7ddrphy_bitslip13_value <= 3'd0;
		main_a7ddrphy_bitslip13_r <= 16'd0;
		main_a7ddrphy_bitslip14_o <= 8'd0;
		main_a7ddrphy_bitslip14_value <= 3'd0;
		main_a7ddrphy_bitslip14_r <= 16'd0;
		main_a7ddrphy_bitslip15_o <= 8'd0;
		main_a7ddrphy_bitslip15_value <= 3'd0;
		main_a7ddrphy_bitslip15_r <= 16'd0;
		main_a7ddrphy_n_rddata_en0 <= 1'd0;
		main_a7ddrphy_n_rddata_en1 <= 1'd0;
		main_a7ddrphy_n_rddata_en2 <= 1'd0;
		main_a7ddrphy_n_rddata_en3 <= 1'd0;
		main_a7ddrphy_n_rddata_en4 <= 1'd0;
		main_a7ddrphy_n_rddata_en5 <= 1'd0;
		main_a7ddrphy_n_rddata_en6 <= 1'd0;
		main_a7ddrphy_n_rddata_en7 <= 1'd0;
		main_a7ddrphy_last_wrdata_en <= 4'd0;
		main_sdram_storage <= 4'd0;
		main_sdram_re <= 1'd0;
		main_sdram_phaseinjector0_command_storage <= 6'd0;
		main_sdram_phaseinjector0_command_re <= 1'd0;
		main_sdram_phaseinjector0_address_storage <= 14'd0;
		main_sdram_phaseinjector0_address_re <= 1'd0;
		main_sdram_phaseinjector0_baddress_storage <= 3'd0;
		main_sdram_phaseinjector0_baddress_re <= 1'd0;
		main_sdram_phaseinjector0_wrdata_storage <= 32'd0;
		main_sdram_phaseinjector0_wrdata_re <= 1'd0;
		main_sdram_phaseinjector0_status <= 32'd0;
		main_sdram_phaseinjector1_command_storage <= 6'd0;
		main_sdram_phaseinjector1_command_re <= 1'd0;
		main_sdram_phaseinjector1_address_storage <= 14'd0;
		main_sdram_phaseinjector1_address_re <= 1'd0;
		main_sdram_phaseinjector1_baddress_storage <= 3'd0;
		main_sdram_phaseinjector1_baddress_re <= 1'd0;
		main_sdram_phaseinjector1_wrdata_storage <= 32'd0;
		main_sdram_phaseinjector1_wrdata_re <= 1'd0;
		main_sdram_phaseinjector1_status <= 32'd0;
		main_sdram_phaseinjector2_command_storage <= 6'd0;
		main_sdram_phaseinjector2_command_re <= 1'd0;
		main_sdram_phaseinjector2_address_storage <= 14'd0;
		main_sdram_phaseinjector2_address_re <= 1'd0;
		main_sdram_phaseinjector2_baddress_storage <= 3'd0;
		main_sdram_phaseinjector2_baddress_re <= 1'd0;
		main_sdram_phaseinjector2_wrdata_storage <= 32'd0;
		main_sdram_phaseinjector2_wrdata_re <= 1'd0;
		main_sdram_phaseinjector2_status <= 32'd0;
		main_sdram_phaseinjector3_command_storage <= 6'd0;
		main_sdram_phaseinjector3_command_re <= 1'd0;
		main_sdram_phaseinjector3_address_storage <= 14'd0;
		main_sdram_phaseinjector3_address_re <= 1'd0;
		main_sdram_phaseinjector3_baddress_storage <= 3'd0;
		main_sdram_phaseinjector3_baddress_re <= 1'd0;
		main_sdram_phaseinjector3_wrdata_storage <= 32'd0;
		main_sdram_phaseinjector3_wrdata_re <= 1'd0;
		main_sdram_phaseinjector3_status <= 32'd0;
		main_sdram_dfi_p0_address <= 14'd0;
		main_sdram_dfi_p0_bank <= 3'd0;
		main_sdram_dfi_p0_cas_n <= 1'd1;
		main_sdram_dfi_p0_cs_n <= 1'd1;
		main_sdram_dfi_p0_ras_n <= 1'd1;
		main_sdram_dfi_p0_we_n <= 1'd1;
		main_sdram_dfi_p0_wrdata_en <= 1'd0;
		main_sdram_dfi_p0_rddata_en <= 1'd0;
		main_sdram_dfi_p1_address <= 14'd0;
		main_sdram_dfi_p1_bank <= 3'd0;
		main_sdram_dfi_p1_cas_n <= 1'd1;
		main_sdram_dfi_p1_cs_n <= 1'd1;
		main_sdram_dfi_p1_ras_n <= 1'd1;
		main_sdram_dfi_p1_we_n <= 1'd1;
		main_sdram_dfi_p1_wrdata_en <= 1'd0;
		main_sdram_dfi_p1_rddata_en <= 1'd0;
		main_sdram_dfi_p2_address <= 14'd0;
		main_sdram_dfi_p2_bank <= 3'd0;
		main_sdram_dfi_p2_cas_n <= 1'd1;
		main_sdram_dfi_p2_cs_n <= 1'd1;
		main_sdram_dfi_p2_ras_n <= 1'd1;
		main_sdram_dfi_p2_we_n <= 1'd1;
		main_sdram_dfi_p2_wrdata_en <= 1'd0;
		main_sdram_dfi_p2_rddata_en <= 1'd0;
		main_sdram_dfi_p3_address <= 14'd0;
		main_sdram_dfi_p3_bank <= 3'd0;
		main_sdram_dfi_p3_cas_n <= 1'd1;
		main_sdram_dfi_p3_cs_n <= 1'd1;
		main_sdram_dfi_p3_ras_n <= 1'd1;
		main_sdram_dfi_p3_we_n <= 1'd1;
		main_sdram_dfi_p3_wrdata_en <= 1'd0;
		main_sdram_dfi_p3_rddata_en <= 1'd0;
		main_sdram_cmd_payload_a <= 14'd0;
		main_sdram_cmd_payload_ba <= 3'd0;
		main_sdram_cmd_payload_cas <= 1'd0;
		main_sdram_cmd_payload_ras <= 1'd0;
		main_sdram_cmd_payload_we <= 1'd0;
		main_sdram_timer_count1 <= 9'd390;
		main_sdram_postponer_req_o <= 1'd0;
		main_sdram_postponer_count <= 1'd0;
		main_sdram_sequencer_done1 <= 1'd0;
		main_sdram_sequencer_counter <= 6'd0;
		main_sdram_sequencer_count <= 1'd0;
		main_sdram_zqcs_timer_count1 <= 26'd49999999;
		main_sdram_zqcs_executer_done <= 1'd0;
		main_sdram_zqcs_executer_counter <= 5'd0;
		main_sdram_bankmachine0_cmd_buffer_lookahead_level <= 4'd0;
		main_sdram_bankmachine0_cmd_buffer_lookahead_produce <= 3'd0;
		main_sdram_bankmachine0_cmd_buffer_lookahead_consume <= 3'd0;
		main_sdram_bankmachine0_cmd_buffer_source_valid <= 1'd0;
		main_sdram_bankmachine0_cmd_buffer_source_first <= 1'd0;
		main_sdram_bankmachine0_cmd_buffer_source_last <= 1'd0;
		main_sdram_bankmachine0_cmd_buffer_source_payload_we <= 1'd0;
		main_sdram_bankmachine0_cmd_buffer_source_payload_addr <= 21'd0;
		main_sdram_bankmachine0_row <= 14'd0;
		main_sdram_bankmachine0_row_opened <= 1'd0;
		main_sdram_bankmachine0_twtpcon_ready <= 1'd1;
		main_sdram_bankmachine0_twtpcon_count <= 3'd0;
		main_sdram_bankmachine0_trccon_ready <= 1'd1;
		main_sdram_bankmachine0_trccon_count <= 2'd0;
		main_sdram_bankmachine0_trascon_ready <= 1'd1;
		main_sdram_bankmachine0_trascon_count <= 2'd0;
		main_sdram_bankmachine1_cmd_buffer_lookahead_level <= 4'd0;
		main_sdram_bankmachine1_cmd_buffer_lookahead_produce <= 3'd0;
		main_sdram_bankmachine1_cmd_buffer_lookahead_consume <= 3'd0;
		main_sdram_bankmachine1_cmd_buffer_source_valid <= 1'd0;
		main_sdram_bankmachine1_cmd_buffer_source_first <= 1'd0;
		main_sdram_bankmachine1_cmd_buffer_source_last <= 1'd0;
		main_sdram_bankmachine1_cmd_buffer_source_payload_we <= 1'd0;
		main_sdram_bankmachine1_cmd_buffer_source_payload_addr <= 21'd0;
		main_sdram_bankmachine1_row <= 14'd0;
		main_sdram_bankmachine1_row_opened <= 1'd0;
		main_sdram_bankmachine1_twtpcon_ready <= 1'd1;
		main_sdram_bankmachine1_twtpcon_count <= 3'd0;
		main_sdram_bankmachine1_trccon_ready <= 1'd1;
		main_sdram_bankmachine1_trccon_count <= 2'd0;
		main_sdram_bankmachine1_trascon_ready <= 1'd1;
		main_sdram_bankmachine1_trascon_count <= 2'd0;
		main_sdram_bankmachine2_cmd_buffer_lookahead_level <= 4'd0;
		main_sdram_bankmachine2_cmd_buffer_lookahead_produce <= 3'd0;
		main_sdram_bankmachine2_cmd_buffer_lookahead_consume <= 3'd0;
		main_sdram_bankmachine2_cmd_buffer_source_valid <= 1'd0;
		main_sdram_bankmachine2_cmd_buffer_source_first <= 1'd0;
		main_sdram_bankmachine2_cmd_buffer_source_last <= 1'd0;
		main_sdram_bankmachine2_cmd_buffer_source_payload_we <= 1'd0;
		main_sdram_bankmachine2_cmd_buffer_source_payload_addr <= 21'd0;
		main_sdram_bankmachine2_row <= 14'd0;
		main_sdram_bankmachine2_row_opened <= 1'd0;
		main_sdram_bankmachine2_twtpcon_ready <= 1'd1;
		main_sdram_bankmachine2_twtpcon_count <= 3'd0;
		main_sdram_bankmachine2_trccon_ready <= 1'd1;
		main_sdram_bankmachine2_trccon_count <= 2'd0;
		main_sdram_bankmachine2_trascon_ready <= 1'd1;
		main_sdram_bankmachine2_trascon_count <= 2'd0;
		main_sdram_bankmachine3_cmd_buffer_lookahead_level <= 4'd0;
		main_sdram_bankmachine3_cmd_buffer_lookahead_produce <= 3'd0;
		main_sdram_bankmachine3_cmd_buffer_lookahead_consume <= 3'd0;
		main_sdram_bankmachine3_cmd_buffer_source_valid <= 1'd0;
		main_sdram_bankmachine3_cmd_buffer_source_first <= 1'd0;
		main_sdram_bankmachine3_cmd_buffer_source_last <= 1'd0;
		main_sdram_bankmachine3_cmd_buffer_source_payload_we <= 1'd0;
		main_sdram_bankmachine3_cmd_buffer_source_payload_addr <= 21'd0;
		main_sdram_bankmachine3_row <= 14'd0;
		main_sdram_bankmachine3_row_opened <= 1'd0;
		main_sdram_bankmachine3_twtpcon_ready <= 1'd1;
		main_sdram_bankmachine3_twtpcon_count <= 3'd0;
		main_sdram_bankmachine3_trccon_ready <= 1'd1;
		main_sdram_bankmachine3_trccon_count <= 2'd0;
		main_sdram_bankmachine3_trascon_ready <= 1'd1;
		main_sdram_bankmachine3_trascon_count <= 2'd0;
		main_sdram_bankmachine4_cmd_buffer_lookahead_level <= 4'd0;
		main_sdram_bankmachine4_cmd_buffer_lookahead_produce <= 3'd0;
		main_sdram_bankmachine4_cmd_buffer_lookahead_consume <= 3'd0;
		main_sdram_bankmachine4_cmd_buffer_source_valid <= 1'd0;
		main_sdram_bankmachine4_cmd_buffer_source_first <= 1'd0;
		main_sdram_bankmachine4_cmd_buffer_source_last <= 1'd0;
		main_sdram_bankmachine4_cmd_buffer_source_payload_we <= 1'd0;
		main_sdram_bankmachine4_cmd_buffer_source_payload_addr <= 21'd0;
		main_sdram_bankmachine4_row <= 14'd0;
		main_sdram_bankmachine4_row_opened <= 1'd0;
		main_sdram_bankmachine4_twtpcon_ready <= 1'd1;
		main_sdram_bankmachine4_twtpcon_count <= 3'd0;
		main_sdram_bankmachine4_trccon_ready <= 1'd1;
		main_sdram_bankmachine4_trccon_count <= 2'd0;
		main_sdram_bankmachine4_trascon_ready <= 1'd1;
		main_sdram_bankmachine4_trascon_count <= 2'd0;
		main_sdram_bankmachine5_cmd_buffer_lookahead_level <= 4'd0;
		main_sdram_bankmachine5_cmd_buffer_lookahead_produce <= 3'd0;
		main_sdram_bankmachine5_cmd_buffer_lookahead_consume <= 3'd0;
		main_sdram_bankmachine5_cmd_buffer_source_valid <= 1'd0;
		main_sdram_bankmachine5_cmd_buffer_source_first <= 1'd0;
		main_sdram_bankmachine5_cmd_buffer_source_last <= 1'd0;
		main_sdram_bankmachine5_cmd_buffer_source_payload_we <= 1'd0;
		main_sdram_bankmachine5_cmd_buffer_source_payload_addr <= 21'd0;
		main_sdram_bankmachine5_row <= 14'd0;
		main_sdram_bankmachine5_row_opened <= 1'd0;
		main_sdram_bankmachine5_twtpcon_ready <= 1'd1;
		main_sdram_bankmachine5_twtpcon_count <= 3'd0;
		main_sdram_bankmachine5_trccon_ready <= 1'd1;
		main_sdram_bankmachine5_trccon_count <= 2'd0;
		main_sdram_bankmachine5_trascon_ready <= 1'd1;
		main_sdram_bankmachine5_trascon_count <= 2'd0;
		main_sdram_bankmachine6_cmd_buffer_lookahead_level <= 4'd0;
		main_sdram_bankmachine6_cmd_buffer_lookahead_produce <= 3'd0;
		main_sdram_bankmachine6_cmd_buffer_lookahead_consume <= 3'd0;
		main_sdram_bankmachine6_cmd_buffer_source_valid <= 1'd0;
		main_sdram_bankmachine6_cmd_buffer_source_first <= 1'd0;
		main_sdram_bankmachine6_cmd_buffer_source_last <= 1'd0;
		main_sdram_bankmachine6_cmd_buffer_source_payload_we <= 1'd0;
		main_sdram_bankmachine6_cmd_buffer_source_payload_addr <= 21'd0;
		main_sdram_bankmachine6_row <= 14'd0;
		main_sdram_bankmachine6_row_opened <= 1'd0;
		main_sdram_bankmachine6_twtpcon_ready <= 1'd1;
		main_sdram_bankmachine6_twtpcon_count <= 3'd0;
		main_sdram_bankmachine6_trccon_ready <= 1'd1;
		main_sdram_bankmachine6_trccon_count <= 2'd0;
		main_sdram_bankmachine6_trascon_ready <= 1'd1;
		main_sdram_bankmachine6_trascon_count <= 2'd0;
		main_sdram_bankmachine7_cmd_buffer_lookahead_level <= 4'd0;
		main_sdram_bankmachine7_cmd_buffer_lookahead_produce <= 3'd0;
		main_sdram_bankmachine7_cmd_buffer_lookahead_consume <= 3'd0;
		main_sdram_bankmachine7_cmd_buffer_source_valid <= 1'd0;
		main_sdram_bankmachine7_cmd_buffer_source_first <= 1'd0;
		main_sdram_bankmachine7_cmd_buffer_source_last <= 1'd0;
		main_sdram_bankmachine7_cmd_buffer_source_payload_we <= 1'd0;
		main_sdram_bankmachine7_cmd_buffer_source_payload_addr <= 21'd0;
		main_sdram_bankmachine7_row <= 14'd0;
		main_sdram_bankmachine7_row_opened <= 1'd0;
		main_sdram_bankmachine7_twtpcon_ready <= 1'd1;
		main_sdram_bankmachine7_twtpcon_count <= 3'd0;
		main_sdram_bankmachine7_trccon_ready <= 1'd1;
		main_sdram_bankmachine7_trccon_count <= 2'd0;
		main_sdram_bankmachine7_trascon_ready <= 1'd1;
		main_sdram_bankmachine7_trascon_count <= 2'd0;
		main_sdram_choose_cmd_grant <= 3'd0;
		main_sdram_choose_req_grant <= 3'd0;
		main_sdram_trrdcon_ready <= 1'd1;
		main_sdram_trrdcon_count <= 1'd0;
		main_sdram_tfawcon_ready <= 1'd1;
		main_sdram_tfawcon_window <= 3'd0;
		main_sdram_tccdcon_ready <= 1'd1;
		main_sdram_tccdcon_count <= 1'd0;
		main_sdram_twtrcon_ready <= 1'd1;
		main_sdram_twtrcon_count <= 3'd0;
		main_sdram_time0 <= 5'd0;
		main_sdram_time1 <= 4'd0;
		main_adr_offset_r <= 2'd0;
		main_count <= 1'd0;
		builder_uartwishbonebridge_state <= 3'd0;
		builder_wb2csr_state <= 1'd0;
		builder_refresher_state <= 2'd0;
		builder_bankmachine0_state <= 3'd0;
		builder_bankmachine1_state <= 3'd0;
		builder_bankmachine2_state <= 3'd0;
		builder_bankmachine3_state <= 3'd0;
		builder_bankmachine4_state <= 3'd0;
		builder_bankmachine5_state <= 3'd0;
		builder_bankmachine6_state <= 3'd0;
		builder_bankmachine7_state <= 3'd0;
		builder_multiplexer_state <= 4'd0;
		builder_rbank <= 3'd0;
		builder_wbank <= 3'd0;
		builder_new_master_wdata_ready0 <= 1'd0;
		builder_new_master_wdata_ready1 <= 1'd0;
		builder_new_master_wdata_ready2 <= 1'd0;
		builder_new_master_rdata_valid0 <= 1'd0;
		builder_new_master_rdata_valid1 <= 1'd0;
		builder_new_master_rdata_valid2 <= 1'd0;
		builder_new_master_rdata_valid3 <= 1'd0;
		builder_new_master_rdata_valid4 <= 1'd0;
		builder_new_master_rdata_valid5 <= 1'd0;
		builder_new_master_rdata_valid6 <= 1'd0;
		builder_new_master_rdata_valid7 <= 1'd0;
		builder_new_master_rdata_valid8 <= 1'd0;
		builder_new_master_rdata_valid9 <= 1'd0;
		builder_fullmemorywe_state <= 2'd0;
		builder_litedramwishbone2native_state <= 2'd0;
		builder_basesoc_slave_sel_r <= 3'd0;
		builder_basesoc_count <= 20'd1000000;
		builder_basesoc_csrbankarray_interface0_bank_bus_dat_r <= 8'd0;
		builder_basesoc_csrbankarray_interface1_bank_bus_dat_r <= 8'd0;
		builder_basesoc_csrbankarray_sel_r <= 1'd0;
		builder_basesoc_csrbankarray_interface2_bank_bus_dat_r <= 8'd0;
		builder_basesoc_csrbankarray_interface3_bank_bus_dat_r <= 8'd0;
	end
	builder_regs0 <= serial_rx;
	builder_regs1 <= builder_regs0;
end
reg [31:0] mem[0:1023];
reg [9:0] memadr;
always @(posedge sys_clk) begin
	if (main_sram_we[0])
		mem[main_sram_adr][7:0] <= main_sram_dat_w[7:0];
	if (main_sram_we[1])
		mem[main_sram_adr][15:8] <= main_sram_dat_w[15:8];
	if (main_sram_we[2])
		mem[main_sram_adr][23:16] <= main_sram_dat_w[23:16];
	if (main_sram_we[3])
		mem[main_sram_adr][31:24] <= main_sram_dat_w[31:24];
	memadr <= main_sram_adr;
end
assign main_sram_dat_r = mem[memadr];
initial begin
	$readmemh("mem.init", mem);
end
reg [7:0] mem_1[0:73];
reg [6:0] memadr_1;
always @(posedge sys_clk) begin
	memadr_1 <= builder_basesoc_csrbankarray_adr;
end
assign builder_basesoc_csrbankarray_dat_r = mem_1[memadr_1];
initial begin
	$readmemh("mem_1.init", mem_1);
end
(* LOC="BUFGCTRL_X0Y16" *)
BUFG BUFG(
	.I(clk100),
	.O(main_pll_clkin)
);
(* LOC="BUFGCTRL_X0Y0" *)
BUFG BUFG_1(
	.I(main_clkout0),
	.O(main_clkout_buf0)
);
(* LOC="BUFGCTRL_X0Y1" *)
BUFG BUFG_2(
	.I(main_clkout1),
	.O(main_clkout_buf1)
);
(* LOC="BUFGCTRL_X0Y3" *)
BUFG BUFG_3(
	.I(main_clkout2),
	.O(main_clkout_buf2)
);
(* LOC="BUFGCTRL_X0Y2" *)
BUFG BUFG_4(
	.I(main_clkout3),
	.O(main_clkout_buf3)
);
(* LOC="BUFGCTRL_X0Y4" *)
BUFG BUFG_5(
	.I((~main_clkout_buf1)),
	.O(main_clkout_buf4)
);
(* LOC="IDELAYCTRL_X1Y0" *)
IDELAYCTRL IDELAYCTRL(
	.REFCLK(clk200_clk),
	.RST(main_ic_reset),
	.RDY(idelayctl_rdy)
);
wire tq;
OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(1'd0),
	.D2(1'd1),
	.D3(1'd0),
	.D4(1'd1),
	.D5(1'd0),
	.D6(1'd1),
	.D7(1'd0),
	.D8(1'd1),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(main_a7ddrphy_sd_clk_se_nodelay),
	.TQ(tq),
	.TCE(1'd1),
	.T1(1'b0)
);
OBUFTDS OBUFTDS_2(
	.I(main_a7ddrphy_sd_clk_se_nodelay),
	.O(ddram_clk_p),
	.OB(ddram_clk_n),
	.T(tq)
);
OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_1 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_a7ddrphy_dfi_p0_address[0]),
	.D2(main_a7ddrphy_dfi_p0_address[0]),
	.D3(main_a7ddrphy_dfi_p1_address[0]),
	.D4(main_a7ddrphy_dfi_p1_address[0]),
	.D5(main_a7ddrphy_dfi_p2_address[0]),
	.D6(main_a7ddrphy_dfi_p2_address[0]),
	.D7(main_a7ddrphy_dfi_p3_address[0]),
	.D8(main_a7ddrphy_dfi_p3_address[0]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a_iob[0])
);
OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_2 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_a7ddrphy_dfi_p0_address[1]),
	.D2(main_a7ddrphy_dfi_p0_address[1]),
	.D3(main_a7ddrphy_dfi_p1_address[1]),
	.D4(main_a7ddrphy_dfi_p1_address[1]),
	.D5(main_a7ddrphy_dfi_p2_address[1]),
	.D6(main_a7ddrphy_dfi_p2_address[1]),
	.D7(main_a7ddrphy_dfi_p3_address[1]),
	.D8(main_a7ddrphy_dfi_p3_address[1]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a_iob[1])
);
OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_3 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_a7ddrphy_dfi_p0_address[2]),
	.D2(main_a7ddrphy_dfi_p0_address[2]),
	.D3(main_a7ddrphy_dfi_p1_address[2]),
	.D4(main_a7ddrphy_dfi_p1_address[2]),
	.D5(main_a7ddrphy_dfi_p2_address[2]),
	.D6(main_a7ddrphy_dfi_p2_address[2]),
	.D7(main_a7ddrphy_dfi_p3_address[2]),
	.D8(main_a7ddrphy_dfi_p3_address[2]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a_iob[2])
);
OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_4 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_a7ddrphy_dfi_p0_address[3]),
	.D2(main_a7ddrphy_dfi_p0_address[3]),
	.D3(main_a7ddrphy_dfi_p1_address[3]),
	.D4(main_a7ddrphy_dfi_p1_address[3]),
	.D5(main_a7ddrphy_dfi_p2_address[3]),
	.D6(main_a7ddrphy_dfi_p2_address[3]),
	.D7(main_a7ddrphy_dfi_p3_address[3]),
	.D8(main_a7ddrphy_dfi_p3_address[3]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a_iob[3])
);
OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_5 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_a7ddrphy_dfi_p0_address[4]),
	.D2(main_a7ddrphy_dfi_p0_address[4]),
	.D3(main_a7ddrphy_dfi_p1_address[4]),
	.D4(main_a7ddrphy_dfi_p1_address[4]),
	.D5(main_a7ddrphy_dfi_p2_address[4]),
	.D6(main_a7ddrphy_dfi_p2_address[4]),
	.D7(main_a7ddrphy_dfi_p3_address[4]),
	.D8(main_a7ddrphy_dfi_p3_address[4]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a_iob[4])
);
OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_6 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_a7ddrphy_dfi_p0_address[5]),
	.D2(main_a7ddrphy_dfi_p0_address[5]),
	.D3(main_a7ddrphy_dfi_p1_address[5]),
	.D4(main_a7ddrphy_dfi_p1_address[5]),
	.D5(main_a7ddrphy_dfi_p2_address[5]),
	.D6(main_a7ddrphy_dfi_p2_address[5]),
	.D7(main_a7ddrphy_dfi_p3_address[5]),
	.D8(main_a7ddrphy_dfi_p3_address[5]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a_iob[5])
);
OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_7 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_a7ddrphy_dfi_p0_address[6]),
	.D2(main_a7ddrphy_dfi_p0_address[6]),
	.D3(main_a7ddrphy_dfi_p1_address[6]),
	.D4(main_a7ddrphy_dfi_p1_address[6]),
	.D5(main_a7ddrphy_dfi_p2_address[6]),
	.D6(main_a7ddrphy_dfi_p2_address[6]),
	.D7(main_a7ddrphy_dfi_p3_address[6]),
	.D8(main_a7ddrphy_dfi_p3_address[6]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a_iob[6])
);
OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_8 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_a7ddrphy_dfi_p0_address[7]),
	.D2(main_a7ddrphy_dfi_p0_address[7]),
	.D3(main_a7ddrphy_dfi_p1_address[7]),
	.D4(main_a7ddrphy_dfi_p1_address[7]),
	.D5(main_a7ddrphy_dfi_p2_address[7]),
	.D6(main_a7ddrphy_dfi_p2_address[7]),
	.D7(main_a7ddrphy_dfi_p3_address[7]),
	.D8(main_a7ddrphy_dfi_p3_address[7]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a_iob[7])
);
OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_9 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_a7ddrphy_dfi_p0_address[8]),
	.D2(main_a7ddrphy_dfi_p0_address[8]),
	.D3(main_a7ddrphy_dfi_p1_address[8]),
	.D4(main_a7ddrphy_dfi_p1_address[8]),
	.D5(main_a7ddrphy_dfi_p2_address[8]),
	.D6(main_a7ddrphy_dfi_p2_address[8]),
	.D7(main_a7ddrphy_dfi_p3_address[8]),
	.D8(main_a7ddrphy_dfi_p3_address[8]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a_iob[8])
);
OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_10 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_a7ddrphy_dfi_p0_address[9]),
	.D2(main_a7ddrphy_dfi_p0_address[9]),
	.D3(main_a7ddrphy_dfi_p1_address[9]),
	.D4(main_a7ddrphy_dfi_p1_address[9]),
	.D5(main_a7ddrphy_dfi_p2_address[9]),
	.D6(main_a7ddrphy_dfi_p2_address[9]),
	.D7(main_a7ddrphy_dfi_p3_address[9]),
	.D8(main_a7ddrphy_dfi_p3_address[9]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a_iob[9])
);
OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_11 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_a7ddrphy_dfi_p0_address[10]),
	.D2(main_a7ddrphy_dfi_p0_address[10]),
	.D3(main_a7ddrphy_dfi_p1_address[10]),
	.D4(main_a7ddrphy_dfi_p1_address[10]),
	.D5(main_a7ddrphy_dfi_p2_address[10]),
	.D6(main_a7ddrphy_dfi_p2_address[10]),
	.D7(main_a7ddrphy_dfi_p3_address[10]),
	.D8(main_a7ddrphy_dfi_p3_address[10]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a_iob[10])
);
OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_12 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_a7ddrphy_dfi_p0_address[11]),
	.D2(main_a7ddrphy_dfi_p0_address[11]),
	.D3(main_a7ddrphy_dfi_p1_address[11]),
	.D4(main_a7ddrphy_dfi_p1_address[11]),
	.D5(main_a7ddrphy_dfi_p2_address[11]),
	.D6(main_a7ddrphy_dfi_p2_address[11]),
	.D7(main_a7ddrphy_dfi_p3_address[11]),
	.D8(main_a7ddrphy_dfi_p3_address[11]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a_iob[11])
);
OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_13 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_a7ddrphy_dfi_p0_address[12]),
	.D2(main_a7ddrphy_dfi_p0_address[12]),
	.D3(main_a7ddrphy_dfi_p1_address[12]),
	.D4(main_a7ddrphy_dfi_p1_address[12]),
	.D5(main_a7ddrphy_dfi_p2_address[12]),
	.D6(main_a7ddrphy_dfi_p2_address[12]),
	.D7(main_a7ddrphy_dfi_p3_address[12]),
	.D8(main_a7ddrphy_dfi_p3_address[12]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a_iob[12])
);
OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_14 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_a7ddrphy_dfi_p0_address[13]),
	.D2(main_a7ddrphy_dfi_p0_address[13]),
	.D3(main_a7ddrphy_dfi_p1_address[13]),
	.D4(main_a7ddrphy_dfi_p1_address[13]),
	.D5(main_a7ddrphy_dfi_p2_address[13]),
	.D6(main_a7ddrphy_dfi_p2_address[13]),
	.D7(main_a7ddrphy_dfi_p3_address[13]),
	.D8(main_a7ddrphy_dfi_p3_address[13]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_a_iob[13])
);
OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_15 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_a7ddrphy_dfi_p0_bank[0]),
	.D2(main_a7ddrphy_dfi_p0_bank[0]),
	.D3(main_a7ddrphy_dfi_p1_bank[0]),
	.D4(main_a7ddrphy_dfi_p1_bank[0]),
	.D5(main_a7ddrphy_dfi_p2_bank[0]),
	.D6(main_a7ddrphy_dfi_p2_bank[0]),
	.D7(main_a7ddrphy_dfi_p3_bank[0]),
	.D8(main_a7ddrphy_dfi_p3_bank[0]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_ba_iob[0])
);
OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_16 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_a7ddrphy_dfi_p0_bank[1]),
	.D2(main_a7ddrphy_dfi_p0_bank[1]),
	.D3(main_a7ddrphy_dfi_p1_bank[1]),
	.D4(main_a7ddrphy_dfi_p1_bank[1]),
	.D5(main_a7ddrphy_dfi_p2_bank[1]),
	.D6(main_a7ddrphy_dfi_p2_bank[1]),
	.D7(main_a7ddrphy_dfi_p3_bank[1]),
	.D8(main_a7ddrphy_dfi_p3_bank[1]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_ba_iob[1])
);
OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_17 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_a7ddrphy_dfi_p0_bank[2]),
	.D2(main_a7ddrphy_dfi_p0_bank[2]),
	.D3(main_a7ddrphy_dfi_p1_bank[2]),
	.D4(main_a7ddrphy_dfi_p1_bank[2]),
	.D5(main_a7ddrphy_dfi_p2_bank[2]),
	.D6(main_a7ddrphy_dfi_p2_bank[2]),
	.D7(main_a7ddrphy_dfi_p3_bank[2]),
	.D8(main_a7ddrphy_dfi_p3_bank[2]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_ba_iob[2])
);
OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_18 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_a7ddrphy_dfi_p0_ras_n),
	.D2(main_a7ddrphy_dfi_p0_ras_n),
	.D3(main_a7ddrphy_dfi_p1_ras_n),
	.D4(main_a7ddrphy_dfi_p1_ras_n),
	.D5(main_a7ddrphy_dfi_p2_ras_n),
	.D6(main_a7ddrphy_dfi_p2_ras_n),
	.D7(main_a7ddrphy_dfi_p3_ras_n),
	.D8(main_a7ddrphy_dfi_p3_ras_n),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_ras_n_iob)
);
OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_19 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_a7ddrphy_dfi_p0_cas_n),
	.D2(main_a7ddrphy_dfi_p0_cas_n),
	.D3(main_a7ddrphy_dfi_p1_cas_n),
	.D4(main_a7ddrphy_dfi_p1_cas_n),
	.D5(main_a7ddrphy_dfi_p2_cas_n),
	.D6(main_a7ddrphy_dfi_p2_cas_n),
	.D7(main_a7ddrphy_dfi_p3_cas_n),
	.D8(main_a7ddrphy_dfi_p3_cas_n),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_cas_n_iob)
);
OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_20 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_a7ddrphy_dfi_p0_we_n),
	.D2(main_a7ddrphy_dfi_p0_we_n),
	.D3(main_a7ddrphy_dfi_p1_we_n),
	.D4(main_a7ddrphy_dfi_p1_we_n),
	.D5(main_a7ddrphy_dfi_p2_we_n),
	.D6(main_a7ddrphy_dfi_p2_we_n),
	.D7(main_a7ddrphy_dfi_p3_we_n),
	.D8(main_a7ddrphy_dfi_p3_we_n),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_we_n_iob)
);
OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_21 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_a7ddrphy_dfi_p0_cke),
	.D2(main_a7ddrphy_dfi_p0_cke),
	.D3(main_a7ddrphy_dfi_p1_cke),
	.D4(main_a7ddrphy_dfi_p1_cke),
	.D5(main_a7ddrphy_dfi_p2_cke),
	.D6(main_a7ddrphy_dfi_p2_cke),
	.D7(main_a7ddrphy_dfi_p3_cke),
	.D8(main_a7ddrphy_dfi_p3_cke),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_cke_iob)
);
OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_22 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_a7ddrphy_dfi_p0_odt),
	.D2(main_a7ddrphy_dfi_p0_odt),
	.D3(main_a7ddrphy_dfi_p1_odt),
	.D4(main_a7ddrphy_dfi_p1_odt),
	.D5(main_a7ddrphy_dfi_p2_odt),
	.D6(main_a7ddrphy_dfi_p2_odt),
	.D7(main_a7ddrphy_dfi_p3_odt),
	.D8(main_a7ddrphy_dfi_p3_odt),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_odt_iob)
);
OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_23 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_a7ddrphy_dfi_p0_reset_n),
	.D2(main_a7ddrphy_dfi_p0_reset_n),
	.D3(main_a7ddrphy_dfi_p1_reset_n),
	.D4(main_a7ddrphy_dfi_p1_reset_n),
	.D5(main_a7ddrphy_dfi_p2_reset_n),
	.D6(main_a7ddrphy_dfi_p2_reset_n),
	.D7(main_a7ddrphy_dfi_p3_reset_n),
	.D8(main_a7ddrphy_dfi_p3_reset_n),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_reset_n_iob)
);
OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_24 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_a7ddrphy_dfi_p0_cs_n),
	.D2(main_a7ddrphy_dfi_p0_cs_n),
	.D3(main_a7ddrphy_dfi_p1_cs_n),
	.D4(main_a7ddrphy_dfi_p1_cs_n),
	.D5(main_a7ddrphy_dfi_p2_cs_n),
	.D6(main_a7ddrphy_dfi_p2_cs_n),
	.D7(main_a7ddrphy_dfi_p3_cs_n),
	.D8(main_a7ddrphy_dfi_p3_cs_n),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_cs_n_iob)
);
OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_25 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_a7ddrphy_dfi_p0_wrdata_mask[0]),
	.D2(main_a7ddrphy_dfi_p0_wrdata_mask[2]),
	.D3(main_a7ddrphy_dfi_p1_wrdata_mask[0]),
	.D4(main_a7ddrphy_dfi_p1_wrdata_mask[2]),
	.D5(main_a7ddrphy_dfi_p2_wrdata_mask[0]),
	.D6(main_a7ddrphy_dfi_p2_wrdata_mask[2]),
	.D7(main_a7ddrphy_dfi_p3_wrdata_mask[0]),
	.D8(main_a7ddrphy_dfi_p3_wrdata_mask[2]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_dm_iob[0])
);
OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_26 (
	.CLK(sys4x_dqs_clk),
	.CLKDIV(sys_clk),
	.D1(main_a7ddrphy_dqs_serdes_pattern[0]),
	.D2(main_a7ddrphy_dqs_serdes_pattern[1]),
	.D3(main_a7ddrphy_dqs_serdes_pattern[2]),
	.D4(main_a7ddrphy_dqs_serdes_pattern[3]),
	.D5(main_a7ddrphy_dqs_serdes_pattern[4]),
	.D6(main_a7ddrphy_dqs_serdes_pattern[5]),
	.D7(main_a7ddrphy_dqs_serdes_pattern[6]),
	.D8(main_a7ddrphy_dqs_serdes_pattern[7]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_a7ddrphy_oe_dqs)),
	.TCE(1'd1),
	.OFB(main_a7ddrphy0),
	.OQ(main_a7ddrphy_dqs_nodelay0),
	.TQ(main_a7ddrphy_dqs_t0)
);
OBUFTDS OBUFTDS(
	.I(main_a7ddrphy_dqs_nodelay0),
	.T(main_a7ddrphy_dqs_t0),
	.O(ddram_dqs_p[0]),
	.OB(ddram_dqs_n[0])
);
OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_27 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_a7ddrphy_dfi_p0_wrdata_mask[1]),
	.D2(main_a7ddrphy_dfi_p0_wrdata_mask[3]),
	.D3(main_a7ddrphy_dfi_p1_wrdata_mask[1]),
	.D4(main_a7ddrphy_dfi_p1_wrdata_mask[3]),
	.D5(main_a7ddrphy_dfi_p2_wrdata_mask[1]),
	.D6(main_a7ddrphy_dfi_p2_wrdata_mask[3]),
	.D7(main_a7ddrphy_dfi_p3_wrdata_mask[1]),
	.D8(main_a7ddrphy_dfi_p3_wrdata_mask[3]),
	.OCE(1'd1),
	.RST(sys_rst),
	.OQ(ddram_dm_iob[1])
);
OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_28 (
	.CLK(sys4x_dqs_clk),
	.CLKDIV(sys_clk),
	.D1(main_a7ddrphy_dqs_serdes_pattern[0]),
	.D2(main_a7ddrphy_dqs_serdes_pattern[1]),
	.D3(main_a7ddrphy_dqs_serdes_pattern[2]),
	.D4(main_a7ddrphy_dqs_serdes_pattern[3]),
	.D5(main_a7ddrphy_dqs_serdes_pattern[4]),
	.D6(main_a7ddrphy_dqs_serdes_pattern[5]),
	.D7(main_a7ddrphy_dqs_serdes_pattern[6]),
	.D8(main_a7ddrphy_dqs_serdes_pattern[7]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_a7ddrphy_oe_dqs)),
	.TCE(1'd1),
	.OFB(main_a7ddrphy1),
	.OQ(main_a7ddrphy_dqs_nodelay1),
	.TQ(main_a7ddrphy_dqs_t1)
);
OBUFTDS OBUFTDS_1(
	.I(main_a7ddrphy_dqs_nodelay1),
	.T(main_a7ddrphy_dqs_t1),
	.O(ddram_dqs_p[1]),
	.OB(ddram_dqs_n[1])
);
OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_29 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_a7ddrphy_dfi_p0_wrdata[0]),
	.D2(main_a7ddrphy_dfi_p0_wrdata[16]),
	.D3(main_a7ddrphy_dfi_p1_wrdata[0]),
	.D4(main_a7ddrphy_dfi_p1_wrdata[16]),
	.D5(main_a7ddrphy_dfi_p2_wrdata[0]),
	.D6(main_a7ddrphy_dfi_p2_wrdata[16]),
	.D7(main_a7ddrphy_dfi_p3_wrdata[0]),
	.D8(main_a7ddrphy_dfi_p3_wrdata[16]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_a7ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_a7ddrphy_dq_o_nodelay0),
	.TQ(main_a7ddrphy_dq_t0)
);
ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2 (
	.BITSLIP(1'd0),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB(sys4x_clkb),
	.CLKDIV(sys_clk),
	.DDLY(main_a7ddrphy_dq_i_delayed0),
	.RST(sys_rst),
	.Q1(main_a7ddrphy_dq_i_data0[7]),
	.Q2(main_a7ddrphy_dq_i_data0[6]),
	.Q3(main_a7ddrphy_dq_i_data0[5]),
	.Q4(main_a7ddrphy_dq_i_data0[4]),
	.Q5(main_a7ddrphy_dq_i_data0[3]),
	.Q6(main_a7ddrphy_dq_i_data0[2]),
	.Q7(main_a7ddrphy_dq_i_data0[1]),
	.Q8(main_a7ddrphy_dq_i_data0[0])
);
IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2 (
	.C(sys_clk),
	.CE((main_a7ddrphy_dly_sel_storage[0] & main_a7ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_a7ddrphy_dq_i_nodelay0),
	.INC(1'd1),
	.LD((main_a7ddrphy_dly_sel_storage[0] & main_a7ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_a7ddrphy_dq_i_delayed0)
);
IOBUF IOBUF(
	.I(main_a7ddrphy_dq_o_nodelay0),
	.T(main_a7ddrphy_dq_t0),
	.IO(ddram_dq[0]),
	.O(main_a7ddrphy_dq_i_nodelay0)
);
OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_30 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_a7ddrphy_dfi_p0_wrdata[1]),
	.D2(main_a7ddrphy_dfi_p0_wrdata[17]),
	.D3(main_a7ddrphy_dfi_p1_wrdata[1]),
	.D4(main_a7ddrphy_dfi_p1_wrdata[17]),
	.D5(main_a7ddrphy_dfi_p2_wrdata[1]),
	.D6(main_a7ddrphy_dfi_p2_wrdata[17]),
	.D7(main_a7ddrphy_dfi_p3_wrdata[1]),
	.D8(main_a7ddrphy_dfi_p3_wrdata[17]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_a7ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_a7ddrphy_dq_o_nodelay1),
	.TQ(main_a7ddrphy_dq_t1)
);
ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_1 (
	.BITSLIP(1'd0),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB(sys4x_clkb),
	.CLKDIV(sys_clk),
	.DDLY(main_a7ddrphy_dq_i_delayed1),
	.RST(sys_rst),
	.Q1(main_a7ddrphy_dq_i_data1[7]),
	.Q2(main_a7ddrphy_dq_i_data1[6]),
	.Q3(main_a7ddrphy_dq_i_data1[5]),
	.Q4(main_a7ddrphy_dq_i_data1[4]),
	.Q5(main_a7ddrphy_dq_i_data1[3]),
	.Q6(main_a7ddrphy_dq_i_data1[2]),
	.Q7(main_a7ddrphy_dq_i_data1[1]),
	.Q8(main_a7ddrphy_dq_i_data1[0])
);
IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_1 (
	.C(sys_clk),
	.CE((main_a7ddrphy_dly_sel_storage[0] & main_a7ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_a7ddrphy_dq_i_nodelay1),
	.INC(1'd1),
	.LD((main_a7ddrphy_dly_sel_storage[0] & main_a7ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_a7ddrphy_dq_i_delayed1)
);
IOBUF IOBUF_1(
	.I(main_a7ddrphy_dq_o_nodelay1),
	.T(main_a7ddrphy_dq_t1),
	.IO(ddram_dq[1]),
	.O(main_a7ddrphy_dq_i_nodelay1)
);
OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_31 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_a7ddrphy_dfi_p0_wrdata[2]),
	.D2(main_a7ddrphy_dfi_p0_wrdata[18]),
	.D3(main_a7ddrphy_dfi_p1_wrdata[2]),
	.D4(main_a7ddrphy_dfi_p1_wrdata[18]),
	.D5(main_a7ddrphy_dfi_p2_wrdata[2]),
	.D6(main_a7ddrphy_dfi_p2_wrdata[18]),
	.D7(main_a7ddrphy_dfi_p3_wrdata[2]),
	.D8(main_a7ddrphy_dfi_p3_wrdata[18]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_a7ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_a7ddrphy_dq_o_nodelay2),
	.TQ(main_a7ddrphy_dq_t2)
);
ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_2 (
	.BITSLIP(1'd0),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB(sys4x_clkb),
	.CLKDIV(sys_clk),
	.DDLY(main_a7ddrphy_dq_i_delayed2),
	.RST(sys_rst),
	.Q1(main_a7ddrphy_dq_i_data2[7]),
	.Q2(main_a7ddrphy_dq_i_data2[6]),
	.Q3(main_a7ddrphy_dq_i_data2[5]),
	.Q4(main_a7ddrphy_dq_i_data2[4]),
	.Q5(main_a7ddrphy_dq_i_data2[3]),
	.Q6(main_a7ddrphy_dq_i_data2[2]),
	.Q7(main_a7ddrphy_dq_i_data2[1]),
	.Q8(main_a7ddrphy_dq_i_data2[0])
);
IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_2 (
	.C(sys_clk),
	.CE((main_a7ddrphy_dly_sel_storage[0] & main_a7ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_a7ddrphy_dq_i_nodelay2),
	.INC(1'd1),
	.LD((main_a7ddrphy_dly_sel_storage[0] & main_a7ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_a7ddrphy_dq_i_delayed2)
);
IOBUF IOBUF_2(
	.I(main_a7ddrphy_dq_o_nodelay2),
	.T(main_a7ddrphy_dq_t2),
	.IO(ddram_dq[2]),
	.O(main_a7ddrphy_dq_i_nodelay2)
);
OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_32 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_a7ddrphy_dfi_p0_wrdata[3]),
	.D2(main_a7ddrphy_dfi_p0_wrdata[19]),
	.D3(main_a7ddrphy_dfi_p1_wrdata[3]),
	.D4(main_a7ddrphy_dfi_p1_wrdata[19]),
	.D5(main_a7ddrphy_dfi_p2_wrdata[3]),
	.D6(main_a7ddrphy_dfi_p2_wrdata[19]),
	.D7(main_a7ddrphy_dfi_p3_wrdata[3]),
	.D8(main_a7ddrphy_dfi_p3_wrdata[19]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_a7ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_a7ddrphy_dq_o_nodelay3),
	.TQ(main_a7ddrphy_dq_t3)
);
ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_3 (
	.BITSLIP(1'd0),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB(sys4x_clkb),
	.CLKDIV(sys_clk),
	.DDLY(main_a7ddrphy_dq_i_delayed3),
	.RST(sys_rst),
	.Q1(main_a7ddrphy_dq_i_data3[7]),
	.Q2(main_a7ddrphy_dq_i_data3[6]),
	.Q3(main_a7ddrphy_dq_i_data3[5]),
	.Q4(main_a7ddrphy_dq_i_data3[4]),
	.Q5(main_a7ddrphy_dq_i_data3[3]),
	.Q6(main_a7ddrphy_dq_i_data3[2]),
	.Q7(main_a7ddrphy_dq_i_data3[1]),
	.Q8(main_a7ddrphy_dq_i_data3[0])
);
IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_3 (
	.C(sys_clk),
	.CE((main_a7ddrphy_dly_sel_storage[0] & main_a7ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_a7ddrphy_dq_i_nodelay3),
	.INC(1'd1),
	.LD((main_a7ddrphy_dly_sel_storage[0] & main_a7ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_a7ddrphy_dq_i_delayed3)
);
IOBUF IOBUF_3(
	.I(main_a7ddrphy_dq_o_nodelay3),
	.T(main_a7ddrphy_dq_t3),
	.IO(ddram_dq[3]),
	.O(main_a7ddrphy_dq_i_nodelay3)
);
OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_33 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_a7ddrphy_dfi_p0_wrdata[4]),
	.D2(main_a7ddrphy_dfi_p0_wrdata[20]),
	.D3(main_a7ddrphy_dfi_p1_wrdata[4]),
	.D4(main_a7ddrphy_dfi_p1_wrdata[20]),
	.D5(main_a7ddrphy_dfi_p2_wrdata[4]),
	.D6(main_a7ddrphy_dfi_p2_wrdata[20]),
	.D7(main_a7ddrphy_dfi_p3_wrdata[4]),
	.D8(main_a7ddrphy_dfi_p3_wrdata[20]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_a7ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_a7ddrphy_dq_o_nodelay4),
	.TQ(main_a7ddrphy_dq_t4)
);
ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_4 (
	.BITSLIP(1'd0),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB(sys4x_clkb),
	.CLKDIV(sys_clk),
	.DDLY(main_a7ddrphy_dq_i_delayed4),
	.RST(sys_rst),
	.Q1(main_a7ddrphy_dq_i_data4[7]),
	.Q2(main_a7ddrphy_dq_i_data4[6]),
	.Q3(main_a7ddrphy_dq_i_data4[5]),
	.Q4(main_a7ddrphy_dq_i_data4[4]),
	.Q5(main_a7ddrphy_dq_i_data4[3]),
	.Q6(main_a7ddrphy_dq_i_data4[2]),
	.Q7(main_a7ddrphy_dq_i_data4[1]),
	.Q8(main_a7ddrphy_dq_i_data4[0])
);
IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_4 (
	.C(sys_clk),
	.CE((main_a7ddrphy_dly_sel_storage[0] & main_a7ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_a7ddrphy_dq_i_nodelay4),
	.INC(1'd1),
	.LD((main_a7ddrphy_dly_sel_storage[0] & main_a7ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_a7ddrphy_dq_i_delayed4)
);
IOBUF IOBUF_4(
	.I(main_a7ddrphy_dq_o_nodelay4),
	.T(main_a7ddrphy_dq_t4),
	.IO(ddram_dq[4]),
	.O(main_a7ddrphy_dq_i_nodelay4)
);
OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_34 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_a7ddrphy_dfi_p0_wrdata[5]),
	.D2(main_a7ddrphy_dfi_p0_wrdata[21]),
	.D3(main_a7ddrphy_dfi_p1_wrdata[5]),
	.D4(main_a7ddrphy_dfi_p1_wrdata[21]),
	.D5(main_a7ddrphy_dfi_p2_wrdata[5]),
	.D6(main_a7ddrphy_dfi_p2_wrdata[21]),
	.D7(main_a7ddrphy_dfi_p3_wrdata[5]),
	.D8(main_a7ddrphy_dfi_p3_wrdata[21]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_a7ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_a7ddrphy_dq_o_nodelay5),
	.TQ(main_a7ddrphy_dq_t5)
);
ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_5 (
	.BITSLIP(1'd0),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB(sys4x_clkb),
	.CLKDIV(sys_clk),
	.DDLY(main_a7ddrphy_dq_i_delayed5),
	.RST(sys_rst),
	.Q1(main_a7ddrphy_dq_i_data5[7]),
	.Q2(main_a7ddrphy_dq_i_data5[6]),
	.Q3(main_a7ddrphy_dq_i_data5[5]),
	.Q4(main_a7ddrphy_dq_i_data5[4]),
	.Q5(main_a7ddrphy_dq_i_data5[3]),
	.Q6(main_a7ddrphy_dq_i_data5[2]),
	.Q7(main_a7ddrphy_dq_i_data5[1]),
	.Q8(main_a7ddrphy_dq_i_data5[0])
);
IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_5 (
	.C(sys_clk),
	.CE((main_a7ddrphy_dly_sel_storage[0] & main_a7ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_a7ddrphy_dq_i_nodelay5),
	.INC(1'd1),
	.LD((main_a7ddrphy_dly_sel_storage[0] & main_a7ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_a7ddrphy_dq_i_delayed5)
);
IOBUF IOBUF_5(
	.I(main_a7ddrphy_dq_o_nodelay5),
	.T(main_a7ddrphy_dq_t5),
	.IO(ddram_dq[5]),
	.O(main_a7ddrphy_dq_i_nodelay5)
);
OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_35 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_a7ddrphy_dfi_p0_wrdata[6]),
	.D2(main_a7ddrphy_dfi_p0_wrdata[22]),
	.D3(main_a7ddrphy_dfi_p1_wrdata[6]),
	.D4(main_a7ddrphy_dfi_p1_wrdata[22]),
	.D5(main_a7ddrphy_dfi_p2_wrdata[6]),
	.D6(main_a7ddrphy_dfi_p2_wrdata[22]),
	.D7(main_a7ddrphy_dfi_p3_wrdata[6]),
	.D8(main_a7ddrphy_dfi_p3_wrdata[22]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_a7ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_a7ddrphy_dq_o_nodelay6),
	.TQ(main_a7ddrphy_dq_t6)
);
ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_6 (
	.BITSLIP(1'd0),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB(sys4x_clkb),
	.CLKDIV(sys_clk),
	.DDLY(main_a7ddrphy_dq_i_delayed6),
	.RST(sys_rst),
	.Q1(main_a7ddrphy_dq_i_data6[7]),
	.Q2(main_a7ddrphy_dq_i_data6[6]),
	.Q3(main_a7ddrphy_dq_i_data6[5]),
	.Q4(main_a7ddrphy_dq_i_data6[4]),
	.Q5(main_a7ddrphy_dq_i_data6[3]),
	.Q6(main_a7ddrphy_dq_i_data6[2]),
	.Q7(main_a7ddrphy_dq_i_data6[1]),
	.Q8(main_a7ddrphy_dq_i_data6[0])
);
IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_6 (
	.C(sys_clk),
	.CE((main_a7ddrphy_dly_sel_storage[0] & main_a7ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_a7ddrphy_dq_i_nodelay6),
	.INC(1'd1),
	.LD((main_a7ddrphy_dly_sel_storage[0] & main_a7ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_a7ddrphy_dq_i_delayed6)
);
IOBUF IOBUF_6(
	.I(main_a7ddrphy_dq_o_nodelay6),
	.T(main_a7ddrphy_dq_t6),
	.IO(ddram_dq[6]),
	.O(main_a7ddrphy_dq_i_nodelay6)
);
OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_36 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_a7ddrphy_dfi_p0_wrdata[7]),
	.D2(main_a7ddrphy_dfi_p0_wrdata[23]),
	.D3(main_a7ddrphy_dfi_p1_wrdata[7]),
	.D4(main_a7ddrphy_dfi_p1_wrdata[23]),
	.D5(main_a7ddrphy_dfi_p2_wrdata[7]),
	.D6(main_a7ddrphy_dfi_p2_wrdata[23]),
	.D7(main_a7ddrphy_dfi_p3_wrdata[7]),
	.D8(main_a7ddrphy_dfi_p3_wrdata[23]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_a7ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_a7ddrphy_dq_o_nodelay7),
	.TQ(main_a7ddrphy_dq_t7)
);
ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_7 (
	.BITSLIP(1'd0),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB(sys4x_clkb),
	.CLKDIV(sys_clk),
	.DDLY(main_a7ddrphy_dq_i_delayed7),
	.RST(sys_rst),
	.Q1(main_a7ddrphy_dq_i_data7[7]),
	.Q2(main_a7ddrphy_dq_i_data7[6]),
	.Q3(main_a7ddrphy_dq_i_data7[5]),
	.Q4(main_a7ddrphy_dq_i_data7[4]),
	.Q5(main_a7ddrphy_dq_i_data7[3]),
	.Q6(main_a7ddrphy_dq_i_data7[2]),
	.Q7(main_a7ddrphy_dq_i_data7[1]),
	.Q8(main_a7ddrphy_dq_i_data7[0])
);
IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_7 (
	.C(sys_clk),
	.CE((main_a7ddrphy_dly_sel_storage[0] & main_a7ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_a7ddrphy_dq_i_nodelay7),
	.INC(1'd1),
	.LD((main_a7ddrphy_dly_sel_storage[0] & main_a7ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_a7ddrphy_dq_i_delayed7)
);
IOBUF IOBUF_7(
	.I(main_a7ddrphy_dq_o_nodelay7),
	.T(main_a7ddrphy_dq_t7),
	.IO(ddram_dq[7]),
	.O(main_a7ddrphy_dq_i_nodelay7)
);
OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_37 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_a7ddrphy_dfi_p0_wrdata[8]),
	.D2(main_a7ddrphy_dfi_p0_wrdata[24]),
	.D3(main_a7ddrphy_dfi_p1_wrdata[8]),
	.D4(main_a7ddrphy_dfi_p1_wrdata[24]),
	.D5(main_a7ddrphy_dfi_p2_wrdata[8]),
	.D6(main_a7ddrphy_dfi_p2_wrdata[24]),
	.D7(main_a7ddrphy_dfi_p3_wrdata[8]),
	.D8(main_a7ddrphy_dfi_p3_wrdata[24]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_a7ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_a7ddrphy_dq_o_nodelay8),
	.TQ(main_a7ddrphy_dq_t8)
);
ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_8 (
	.BITSLIP(1'd0),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB(sys4x_clkb),
	.CLKDIV(sys_clk),
	.DDLY(main_a7ddrphy_dq_i_delayed8),
	.RST(sys_rst),
	.Q1(main_a7ddrphy_dq_i_data8[7]),
	.Q2(main_a7ddrphy_dq_i_data8[6]),
	.Q3(main_a7ddrphy_dq_i_data8[5]),
	.Q4(main_a7ddrphy_dq_i_data8[4]),
	.Q5(main_a7ddrphy_dq_i_data8[3]),
	.Q6(main_a7ddrphy_dq_i_data8[2]),
	.Q7(main_a7ddrphy_dq_i_data8[1]),
	.Q8(main_a7ddrphy_dq_i_data8[0])
);
IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_8 (
	.C(sys_clk),
	.CE((main_a7ddrphy_dly_sel_storage[1] & main_a7ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_a7ddrphy_dq_i_nodelay8),
	.INC(1'd1),
	.LD((main_a7ddrphy_dly_sel_storage[1] & main_a7ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_a7ddrphy_dq_i_delayed8)
);
IOBUF IOBUF_8(
	.I(main_a7ddrphy_dq_o_nodelay8),
	.T(main_a7ddrphy_dq_t8),
	.IO(ddram_dq[8]),
	.O(main_a7ddrphy_dq_i_nodelay8)
);
OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_38 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_a7ddrphy_dfi_p0_wrdata[9]),
	.D2(main_a7ddrphy_dfi_p0_wrdata[25]),
	.D3(main_a7ddrphy_dfi_p1_wrdata[9]),
	.D4(main_a7ddrphy_dfi_p1_wrdata[25]),
	.D5(main_a7ddrphy_dfi_p2_wrdata[9]),
	.D6(main_a7ddrphy_dfi_p2_wrdata[25]),
	.D7(main_a7ddrphy_dfi_p3_wrdata[9]),
	.D8(main_a7ddrphy_dfi_p3_wrdata[25]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_a7ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_a7ddrphy_dq_o_nodelay9),
	.TQ(main_a7ddrphy_dq_t9)
);
ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_9 (
	.BITSLIP(1'd0),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB(sys4x_clkb),
	.CLKDIV(sys_clk),
	.DDLY(main_a7ddrphy_dq_i_delayed9),
	.RST(sys_rst),
	.Q1(main_a7ddrphy_dq_i_data9[7]),
	.Q2(main_a7ddrphy_dq_i_data9[6]),
	.Q3(main_a7ddrphy_dq_i_data9[5]),
	.Q4(main_a7ddrphy_dq_i_data9[4]),
	.Q5(main_a7ddrphy_dq_i_data9[3]),
	.Q6(main_a7ddrphy_dq_i_data9[2]),
	.Q7(main_a7ddrphy_dq_i_data9[1]),
	.Q8(main_a7ddrphy_dq_i_data9[0])
);
IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_9 (
	.C(sys_clk),
	.CE((main_a7ddrphy_dly_sel_storage[1] & main_a7ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_a7ddrphy_dq_i_nodelay9),
	.INC(1'd1),
	.LD((main_a7ddrphy_dly_sel_storage[1] & main_a7ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_a7ddrphy_dq_i_delayed9)
);
IOBUF IOBUF_9(
	.I(main_a7ddrphy_dq_o_nodelay9),
	.T(main_a7ddrphy_dq_t9),
	.IO(ddram_dq[9]),
	.O(main_a7ddrphy_dq_i_nodelay9)
);
OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_39 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_a7ddrphy_dfi_p0_wrdata[10]),
	.D2(main_a7ddrphy_dfi_p0_wrdata[26]),
	.D3(main_a7ddrphy_dfi_p1_wrdata[10]),
	.D4(main_a7ddrphy_dfi_p1_wrdata[26]),
	.D5(main_a7ddrphy_dfi_p2_wrdata[10]),
	.D6(main_a7ddrphy_dfi_p2_wrdata[26]),
	.D7(main_a7ddrphy_dfi_p3_wrdata[10]),
	.D8(main_a7ddrphy_dfi_p3_wrdata[26]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_a7ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_a7ddrphy_dq_o_nodelay10),
	.TQ(main_a7ddrphy_dq_t10)
);
ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_10 (
	.BITSLIP(1'd0),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB(sys4x_clkb),
	.CLKDIV(sys_clk),
	.DDLY(main_a7ddrphy_dq_i_delayed10),
	.RST(sys_rst),
	.Q1(main_a7ddrphy_dq_i_data10[7]),
	.Q2(main_a7ddrphy_dq_i_data10[6]),
	.Q3(main_a7ddrphy_dq_i_data10[5]),
	.Q4(main_a7ddrphy_dq_i_data10[4]),
	.Q5(main_a7ddrphy_dq_i_data10[3]),
	.Q6(main_a7ddrphy_dq_i_data10[2]),
	.Q7(main_a7ddrphy_dq_i_data10[1]),
	.Q8(main_a7ddrphy_dq_i_data10[0])
);
IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_10 (
	.C(sys_clk),
	.CE((main_a7ddrphy_dly_sel_storage[1] & main_a7ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_a7ddrphy_dq_i_nodelay10),
	.INC(1'd1),
	.LD((main_a7ddrphy_dly_sel_storage[1] & main_a7ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_a7ddrphy_dq_i_delayed10)
);
IOBUF IOBUF_10(
	.I(main_a7ddrphy_dq_o_nodelay10),
	.T(main_a7ddrphy_dq_t10),
	.IO(ddram_dq[10]),
	.O(main_a7ddrphy_dq_i_nodelay10)
);
OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_40 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_a7ddrphy_dfi_p0_wrdata[11]),
	.D2(main_a7ddrphy_dfi_p0_wrdata[27]),
	.D3(main_a7ddrphy_dfi_p1_wrdata[11]),
	.D4(main_a7ddrphy_dfi_p1_wrdata[27]),
	.D5(main_a7ddrphy_dfi_p2_wrdata[11]),
	.D6(main_a7ddrphy_dfi_p2_wrdata[27]),
	.D7(main_a7ddrphy_dfi_p3_wrdata[11]),
	.D8(main_a7ddrphy_dfi_p3_wrdata[27]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_a7ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_a7ddrphy_dq_o_nodelay11),
	.TQ(main_a7ddrphy_dq_t11)
);
ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_11 (
	.BITSLIP(1'd0),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB(sys4x_clkb),
	.CLKDIV(sys_clk),
	.DDLY(main_a7ddrphy_dq_i_delayed11),
	.RST(sys_rst),
	.Q1(main_a7ddrphy_dq_i_data11[7]),
	.Q2(main_a7ddrphy_dq_i_data11[6]),
	.Q3(main_a7ddrphy_dq_i_data11[5]),
	.Q4(main_a7ddrphy_dq_i_data11[4]),
	.Q5(main_a7ddrphy_dq_i_data11[3]),
	.Q6(main_a7ddrphy_dq_i_data11[2]),
	.Q7(main_a7ddrphy_dq_i_data11[1]),
	.Q8(main_a7ddrphy_dq_i_data11[0])
);
IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_11 (
	.C(sys_clk),
	.CE((main_a7ddrphy_dly_sel_storage[1] & main_a7ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_a7ddrphy_dq_i_nodelay11),
	.INC(1'd1),
	.LD((main_a7ddrphy_dly_sel_storage[1] & main_a7ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_a7ddrphy_dq_i_delayed11)
);
IOBUF IOBUF_11(
	.I(main_a7ddrphy_dq_o_nodelay11),
	.T(main_a7ddrphy_dq_t11),
	.IO(ddram_dq[11]),
	.O(main_a7ddrphy_dq_i_nodelay11)
);
OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_41 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_a7ddrphy_dfi_p0_wrdata[12]),
	.D2(main_a7ddrphy_dfi_p0_wrdata[28]),
	.D3(main_a7ddrphy_dfi_p1_wrdata[12]),
	.D4(main_a7ddrphy_dfi_p1_wrdata[28]),
	.D5(main_a7ddrphy_dfi_p2_wrdata[12]),
	.D6(main_a7ddrphy_dfi_p2_wrdata[28]),
	.D7(main_a7ddrphy_dfi_p3_wrdata[12]),
	.D8(main_a7ddrphy_dfi_p3_wrdata[28]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_a7ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_a7ddrphy_dq_o_nodelay12),
	.TQ(main_a7ddrphy_dq_t12)
);
ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_12 (
	.BITSLIP(1'd0),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB(sys4x_clkb),
	.CLKDIV(sys_clk),
	.DDLY(main_a7ddrphy_dq_i_delayed12),
	.RST(sys_rst),
	.Q1(main_a7ddrphy_dq_i_data12[7]),
	.Q2(main_a7ddrphy_dq_i_data12[6]),
	.Q3(main_a7ddrphy_dq_i_data12[5]),
	.Q4(main_a7ddrphy_dq_i_data12[4]),
	.Q5(main_a7ddrphy_dq_i_data12[3]),
	.Q6(main_a7ddrphy_dq_i_data12[2]),
	.Q7(main_a7ddrphy_dq_i_data12[1]),
	.Q8(main_a7ddrphy_dq_i_data12[0])
);
IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_12 (
	.C(sys_clk),
	.CE((main_a7ddrphy_dly_sel_storage[1] & main_a7ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_a7ddrphy_dq_i_nodelay12),
	.INC(1'd1),
	.LD((main_a7ddrphy_dly_sel_storage[1] & main_a7ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_a7ddrphy_dq_i_delayed12)
);
IOBUF IOBUF_12(
	.I(main_a7ddrphy_dq_o_nodelay12),
	.T(main_a7ddrphy_dq_t12),
	.IO(ddram_dq[12]),
	.O(main_a7ddrphy_dq_i_nodelay12)
);
OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_42 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_a7ddrphy_dfi_p0_wrdata[13]),
	.D2(main_a7ddrphy_dfi_p0_wrdata[29]),
	.D3(main_a7ddrphy_dfi_p1_wrdata[13]),
	.D4(main_a7ddrphy_dfi_p1_wrdata[29]),
	.D5(main_a7ddrphy_dfi_p2_wrdata[13]),
	.D6(main_a7ddrphy_dfi_p2_wrdata[29]),
	.D7(main_a7ddrphy_dfi_p3_wrdata[13]),
	.D8(main_a7ddrphy_dfi_p3_wrdata[29]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_a7ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_a7ddrphy_dq_o_nodelay13),
	.TQ(main_a7ddrphy_dq_t13)
);
ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_13 (
	.BITSLIP(1'd0),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB(sys4x_clkb),
	.CLKDIV(sys_clk),
	.DDLY(main_a7ddrphy_dq_i_delayed13),
	.RST(sys_rst),
	.Q1(main_a7ddrphy_dq_i_data13[7]),
	.Q2(main_a7ddrphy_dq_i_data13[6]),
	.Q3(main_a7ddrphy_dq_i_data13[5]),
	.Q4(main_a7ddrphy_dq_i_data13[4]),
	.Q5(main_a7ddrphy_dq_i_data13[3]),
	.Q6(main_a7ddrphy_dq_i_data13[2]),
	.Q7(main_a7ddrphy_dq_i_data13[1]),
	.Q8(main_a7ddrphy_dq_i_data13[0])
);
IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_13 (
	.C(sys_clk),
	.CE((main_a7ddrphy_dly_sel_storage[1] & main_a7ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_a7ddrphy_dq_i_nodelay13),
	.INC(1'd1),
	.LD((main_a7ddrphy_dly_sel_storage[1] & main_a7ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_a7ddrphy_dq_i_delayed13)
);
IOBUF IOBUF_13(
	.I(main_a7ddrphy_dq_o_nodelay13),
	.T(main_a7ddrphy_dq_t13),
	.IO(ddram_dq[13]),
	.O(main_a7ddrphy_dq_i_nodelay13)
);
OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_43 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_a7ddrphy_dfi_p0_wrdata[14]),
	.D2(main_a7ddrphy_dfi_p0_wrdata[30]),
	.D3(main_a7ddrphy_dfi_p1_wrdata[14]),
	.D4(main_a7ddrphy_dfi_p1_wrdata[30]),
	.D5(main_a7ddrphy_dfi_p2_wrdata[14]),
	.D6(main_a7ddrphy_dfi_p2_wrdata[30]),
	.D7(main_a7ddrphy_dfi_p3_wrdata[14]),
	.D8(main_a7ddrphy_dfi_p3_wrdata[30]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_a7ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_a7ddrphy_dq_o_nodelay14),
	.TQ(main_a7ddrphy_dq_t14)
);
ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_14 (
	.BITSLIP(1'd0),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB(sys4x_clkb),
	.CLKDIV(sys_clk),
	.DDLY(main_a7ddrphy_dq_i_delayed14),
	.RST(sys_rst),
	.Q1(main_a7ddrphy_dq_i_data14[7]),
	.Q2(main_a7ddrphy_dq_i_data14[6]),
	.Q3(main_a7ddrphy_dq_i_data14[5]),
	.Q4(main_a7ddrphy_dq_i_data14[4]),
	.Q5(main_a7ddrphy_dq_i_data14[3]),
	.Q6(main_a7ddrphy_dq_i_data14[2]),
	.Q7(main_a7ddrphy_dq_i_data14[1]),
	.Q8(main_a7ddrphy_dq_i_data14[0])
);
IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_14 (
	.C(sys_clk),
	.CE((main_a7ddrphy_dly_sel_storage[1] & main_a7ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_a7ddrphy_dq_i_nodelay14),
	.INC(1'd1),
	.LD((main_a7ddrphy_dly_sel_storage[1] & main_a7ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_a7ddrphy_dq_i_delayed14)
);
IOBUF IOBUF_14(
	.I(main_a7ddrphy_dq_o_nodelay14),
	.T(main_a7ddrphy_dq_t14),
	.IO(ddram_dq[14]),
	.O(main_a7ddrphy_dq_i_nodelay14)
);
OSERDESE2 #(
	.DATA_RATE_OQ("DDR"),
	.DATA_RATE_TQ("BUF"),
	.DATA_WIDTH(4'd8),
	.SERDES_MODE("MASTER"),
	.TRISTATE_WIDTH(1'd1)
) OSERDESE2_44 (
	.CLK(sys4x_clk),
	.CLKDIV(sys_clk),
	.D1(main_a7ddrphy_dfi_p0_wrdata[15]),
	.D2(main_a7ddrphy_dfi_p0_wrdata[31]),
	.D3(main_a7ddrphy_dfi_p1_wrdata[15]),
	.D4(main_a7ddrphy_dfi_p1_wrdata[31]),
	.D5(main_a7ddrphy_dfi_p2_wrdata[15]),
	.D6(main_a7ddrphy_dfi_p2_wrdata[31]),
	.D7(main_a7ddrphy_dfi_p3_wrdata[15]),
	.D8(main_a7ddrphy_dfi_p3_wrdata[31]),
	.OCE(1'd1),
	.RST(sys_rst),
	.T1((~main_a7ddrphy_oe_dq)),
	.TCE(1'd1),
	.OQ(main_a7ddrphy_dq_o_nodelay15),
	.TQ(main_a7ddrphy_dq_t15)
);
ISERDESE2 #(
	.DATA_RATE("DDR"),
	.DATA_WIDTH(4'd8),
	.INTERFACE_TYPE("NETWORKING"),
	.IOBDELAY("IFD"),
	.NUM_CE(1'd1),
	.SERDES_MODE("MASTER")
) ISERDESE2_15 (
	.BITSLIP(1'd0),
	.CE1(1'd1),
	.CLK(sys4x_clk),
	.CLKB(sys4x_clkb),
	.CLKDIV(sys_clk),
	.DDLY(main_a7ddrphy_dq_i_delayed15),
	.RST(sys_rst),
	.Q1(main_a7ddrphy_dq_i_data15[7]),
	.Q2(main_a7ddrphy_dq_i_data15[6]),
	.Q3(main_a7ddrphy_dq_i_data15[5]),
	.Q4(main_a7ddrphy_dq_i_data15[4]),
	.Q5(main_a7ddrphy_dq_i_data15[3]),
	.Q6(main_a7ddrphy_dq_i_data15[2]),
	.Q7(main_a7ddrphy_dq_i_data15[1]),
	.Q8(main_a7ddrphy_dq_i_data15[0])
);
IDELAYE2 #(
	.CINVCTRL_SEL("FALSE"),
	.DELAY_SRC("IDATAIN"),
	.HIGH_PERFORMANCE_MODE("TRUE"),
	.IDELAY_TYPE("VARIABLE"),
	.IDELAY_VALUE(1'd0),
	.PIPE_SEL("FALSE"),
	.REFCLK_FREQUENCY(200.0),
	.SIGNAL_PATTERN("DATA")
) IDELAYE2_15 (
	.C(sys_clk),
	.CE((main_a7ddrphy_dly_sel_storage[1] & main_a7ddrphy_rdly_dq_inc_re)),
	.IDATAIN(main_a7ddrphy_dq_i_nodelay15),
	.INC(1'd1),
	.LD((main_a7ddrphy_dly_sel_storage[1] & main_a7ddrphy_rdly_dq_rst_re)),
	.LDPIPEEN(1'd0),
	.DATAOUT(main_a7ddrphy_dq_i_delayed15)
);
IOBUF IOBUF_15(
	.I(main_a7ddrphy_dq_o_nodelay15),
	.T(main_a7ddrphy_dq_t15),
	.IO(ddram_dq[15]),
	.O(main_a7ddrphy_dq_i_nodelay15)
);
reg [23:0] storage[0:7];
reg [23:0] memdat;
always @(posedge sys_clk) begin
	if (main_sdram_bankmachine0_cmd_buffer_lookahead_wrport_we)
		storage[main_sdram_bankmachine0_cmd_buffer_lookahead_wrport_adr] <= main_sdram_bankmachine0_cmd_buffer_lookahead_wrport_dat_w;
	memdat <= storage[main_sdram_bankmachine0_cmd_buffer_lookahead_wrport_adr];
end
always @(posedge sys_clk) begin
end
assign main_sdram_bankmachine0_cmd_buffer_lookahead_wrport_dat_r = memdat;
assign main_sdram_bankmachine0_cmd_buffer_lookahead_rdport_dat_r = storage[main_sdram_bankmachine0_cmd_buffer_lookahead_rdport_adr];
reg [23:0] storage_1[0:7];
reg [23:0] memdat_1;
always @(posedge sys_clk) begin
	if (main_sdram_bankmachine1_cmd_buffer_lookahead_wrport_we)
		storage_1[main_sdram_bankmachine1_cmd_buffer_lookahead_wrport_adr] <= main_sdram_bankmachine1_cmd_buffer_lookahead_wrport_dat_w;
	memdat_1 <= storage_1[main_sdram_bankmachine1_cmd_buffer_lookahead_wrport_adr];
end
always @(posedge sys_clk) begin
end
assign main_sdram_bankmachine1_cmd_buffer_lookahead_wrport_dat_r = memdat_1;
assign main_sdram_bankmachine1_cmd_buffer_lookahead_rdport_dat_r = storage_1[main_sdram_bankmachine1_cmd_buffer_lookahead_rdport_adr];
reg [23:0] storage_2[0:7];
reg [23:0] memdat_2;
always @(posedge sys_clk) begin
	if (main_sdram_bankmachine2_cmd_buffer_lookahead_wrport_we)
		storage_2[main_sdram_bankmachine2_cmd_buffer_lookahead_wrport_adr] <= main_sdram_bankmachine2_cmd_buffer_lookahead_wrport_dat_w;
	memdat_2 <= storage_2[main_sdram_bankmachine2_cmd_buffer_lookahead_wrport_adr];
end
always @(posedge sys_clk) begin
end
assign main_sdram_bankmachine2_cmd_buffer_lookahead_wrport_dat_r = memdat_2;
assign main_sdram_bankmachine2_cmd_buffer_lookahead_rdport_dat_r = storage_2[main_sdram_bankmachine2_cmd_buffer_lookahead_rdport_adr];
reg [23:0] storage_3[0:7];
reg [23:0] memdat_3;
always @(posedge sys_clk) begin
	if (main_sdram_bankmachine3_cmd_buffer_lookahead_wrport_we)
		storage_3[main_sdram_bankmachine3_cmd_buffer_lookahead_wrport_adr] <= main_sdram_bankmachine3_cmd_buffer_lookahead_wrport_dat_w;
	memdat_3 <= storage_3[main_sdram_bankmachine3_cmd_buffer_lookahead_wrport_adr];
end
always @(posedge sys_clk) begin
end
assign main_sdram_bankmachine3_cmd_buffer_lookahead_wrport_dat_r = memdat_3;
assign main_sdram_bankmachine3_cmd_buffer_lookahead_rdport_dat_r = storage_3[main_sdram_bankmachine3_cmd_buffer_lookahead_rdport_adr];
reg [23:0] storage_4[0:7];
reg [23:0] memdat_4;
always @(posedge sys_clk) begin
	if (main_sdram_bankmachine4_cmd_buffer_lookahead_wrport_we)
		storage_4[main_sdram_bankmachine4_cmd_buffer_lookahead_wrport_adr] <= main_sdram_bankmachine4_cmd_buffer_lookahead_wrport_dat_w;
	memdat_4 <= storage_4[main_sdram_bankmachine4_cmd_buffer_lookahead_wrport_adr];
end
always @(posedge sys_clk) begin
end
assign main_sdram_bankmachine4_cmd_buffer_lookahead_wrport_dat_r = memdat_4;
assign main_sdram_bankmachine4_cmd_buffer_lookahead_rdport_dat_r = storage_4[main_sdram_bankmachine4_cmd_buffer_lookahead_rdport_adr];
reg [23:0] storage_5[0:7];
reg [23:0] memdat_5;
always @(posedge sys_clk) begin
	if (main_sdram_bankmachine5_cmd_buffer_lookahead_wrport_we)
		storage_5[main_sdram_bankmachine5_cmd_buffer_lookahead_wrport_adr] <= main_sdram_bankmachine5_cmd_buffer_lookahead_wrport_dat_w;
	memdat_5 <= storage_5[main_sdram_bankmachine5_cmd_buffer_lookahead_wrport_adr];
end
always @(posedge sys_clk) begin
end
assign main_sdram_bankmachine5_cmd_buffer_lookahead_wrport_dat_r = memdat_5;
assign main_sdram_bankmachine5_cmd_buffer_lookahead_rdport_dat_r = storage_5[main_sdram_bankmachine5_cmd_buffer_lookahead_rdport_adr];
reg [23:0] storage_6[0:7];
reg [23:0] memdat_6;
always @(posedge sys_clk) begin
	if (main_sdram_bankmachine6_cmd_buffer_lookahead_wrport_we)
		storage_6[main_sdram_bankmachine6_cmd_buffer_lookahead_wrport_adr] <= main_sdram_bankmachine6_cmd_buffer_lookahead_wrport_dat_w;
	memdat_6 <= storage_6[main_sdram_bankmachine6_cmd_buffer_lookahead_wrport_adr];
end
always @(posedge sys_clk) begin
end
assign main_sdram_bankmachine6_cmd_buffer_lookahead_wrport_dat_r = memdat_6;
assign main_sdram_bankmachine6_cmd_buffer_lookahead_rdport_dat_r = storage_6[main_sdram_bankmachine6_cmd_buffer_lookahead_rdport_adr];
reg [23:0] storage_7[0:7];
reg [23:0] memdat_7;
always @(posedge sys_clk) begin
	if (main_sdram_bankmachine7_cmd_buffer_lookahead_wrport_we)
		storage_7[main_sdram_bankmachine7_cmd_buffer_lookahead_wrport_adr] <= main_sdram_bankmachine7_cmd_buffer_lookahead_wrport_dat_w;
	memdat_7 <= storage_7[main_sdram_bankmachine7_cmd_buffer_lookahead_wrport_adr];
end
always @(posedge sys_clk) begin
end
assign main_sdram_bankmachine7_cmd_buffer_lookahead_wrport_dat_r = memdat_7;
assign main_sdram_bankmachine7_cmd_buffer_lookahead_rdport_dat_r = storage_7[main_sdram_bankmachine7_cmd_buffer_lookahead_rdport_adr];
reg [31:0] tag_mem[0:1];
reg [0:0] memadr_2;
always @(posedge sys_clk) begin
	if (main_tag_port_we)
		tag_mem[main_tag_port_adr] <= main_tag_port_dat_w;
	memadr_2 <= main_tag_port_adr;
end
assign main_tag_port_dat_r = tag_mem[memadr_2];
(* LOC="PLLE2_ADV_X1Y0" *)
PLLE2_ADV #(
	.CLKFBOUT_MULT(5'd16),
	.CLKIN1_PERIOD(10.0),
	.CLKOUT0_DIVIDE(6'd32),
	.CLKOUT0_PHASE(1'd0),
	.CLKOUT1_DIVIDE(4'd8),
	.CLKOUT1_PHASE(1'd0),
	.CLKOUT2_DIVIDE(4'd8),
	.CLKOUT2_PHASE(7'd90),
	.CLKOUT3_DIVIDE(4'd8),
	.CLKOUT3_PHASE(1'd0),
	.DIVCLK_DIVIDE(1'd1),
	.REF_JITTER1(0.01),
	.STARTUP_WAIT("FALSE")
) PLLE2_ADV (
	.CLKFBIN(builder_pll_fb),
	.CLKIN1(main_pll_clkin),
	.RST(main_reset),
	.CLKFBOUT(builder_pll_fb),
	.CLKOUT0(main_clkout0),
	.CLKOUT1(main_clkout1),
	.CLKOUT2(main_clkout2),
	.CLKOUT3(main_clkout3),
	.LOCKED(main_locked)
);
reg [7:0] data_mem_grain0[0:1];
reg [0:0] memadr_3;
always @(posedge sys_clk) begin
	if (main_data_port_we[0])
		data_mem_grain0[main_data_port_adr] <= main_data_port_dat_w[7:0];
	memadr_3 <= main_data_port_adr;
end
assign main_data_port_dat_r[7:0] = data_mem_grain0[memadr_3];
reg [7:0] data_mem_grain1[0:1];
reg [0:0] memadr_4;
always @(posedge sys_clk) begin
	if (main_data_port_we[1])
		data_mem_grain1[main_data_port_adr] <= main_data_port_dat_w[15:8];
	memadr_4 <= main_data_port_adr;
end
assign main_data_port_dat_r[15:8] = data_mem_grain1[memadr_4];
reg [7:0] data_mem_grain2[0:1];
reg [0:0] memadr_5;
always @(posedge sys_clk) begin
	if (main_data_port_we[2])
		data_mem_grain2[main_data_port_adr] <= main_data_port_dat_w[23:16];
	memadr_5 <= main_data_port_adr;
end
assign main_data_port_dat_r[23:16] = data_mem_grain2[memadr_5];
reg [7:0] data_mem_grain3[0:1];
reg [0:0] memadr_6;
always @(posedge sys_clk) begin
	if (main_data_port_we[3])
		data_mem_grain3[main_data_port_adr] <= main_data_port_dat_w[31:24];
	memadr_6 <= main_data_port_adr;
end
assign main_data_port_dat_r[31:24] = data_mem_grain3[memadr_6];
reg [7:0] data_mem_grain4[0:1];
reg [0:0] memadr_7;
always @(posedge sys_clk) begin
	if (main_data_port_we[4])
		data_mem_grain4[main_data_port_adr] <= main_data_port_dat_w[39:32];
	memadr_7 <= main_data_port_adr;
end
assign main_data_port_dat_r[39:32] = data_mem_grain4[memadr_7];
reg [7:0] data_mem_grain5[0:1];
reg [0:0] memadr_8;
always @(posedge sys_clk) begin
	if (main_data_port_we[5])
		data_mem_grain5[main_data_port_adr] <= main_data_port_dat_w[47:40];
	memadr_8 <= main_data_port_adr;
end
assign main_data_port_dat_r[47:40] = data_mem_grain5[memadr_8];
reg [7:0] data_mem_grain6[0:1];
reg [0:0] memadr_9;
always @(posedge sys_clk) begin
	if (main_data_port_we[6])
		data_mem_grain6[main_data_port_adr] <= main_data_port_dat_w[55:48];
	memadr_9 <= main_data_port_adr;
end
assign main_data_port_dat_r[55:48] = data_mem_grain6[memadr_9];
reg [7:0] data_mem_grain7[0:1];
reg [0:0] memadr_10;
always @(posedge sys_clk) begin
	if (main_data_port_we[7])
		data_mem_grain7[main_data_port_adr] <= main_data_port_dat_w[63:56];
	memadr_10 <= main_data_port_adr;
end
assign main_data_port_dat_r[63:56] = data_mem_grain7[memadr_10];
reg [7:0] data_mem_grain8[0:1];
reg [0:0] memadr_11;
always @(posedge sys_clk) begin
	if (main_data_port_we[8])
		data_mem_grain8[main_data_port_adr] <= main_data_port_dat_w[71:64];
	memadr_11 <= main_data_port_adr;
end
assign main_data_port_dat_r[71:64] = data_mem_grain8[memadr_11];
reg [7:0] data_mem_grain9[0:1];
reg [0:0] memadr_12;
always @(posedge sys_clk) begin
	if (main_data_port_we[9])
		data_mem_grain9[main_data_port_adr] <= main_data_port_dat_w[79:72];
	memadr_12 <= main_data_port_adr;
end
assign main_data_port_dat_r[79:72] = data_mem_grain9[memadr_12];
reg [7:0] data_mem_grain10[0:1];
reg [0:0] memadr_13;
always @(posedge sys_clk) begin
	if (main_data_port_we[10])
		data_mem_grain10[main_data_port_adr] <= main_data_port_dat_w[87:80];
	memadr_13 <= main_data_port_adr;
end
assign main_data_port_dat_r[87:80] = data_mem_grain10[memadr_13];
reg [7:0] data_mem_grain11[0:1];
reg [0:0] memadr_14;
always @(posedge sys_clk) begin
	if (main_data_port_we[11])
		data_mem_grain11[main_data_port_adr] <= main_data_port_dat_w[95:88];
	memadr_14 <= main_data_port_adr;
end
assign main_data_port_dat_r[95:88] = data_mem_grain11[memadr_14];
reg [7:0] data_mem_grain12[0:1];
reg [0:0] memadr_15;
always @(posedge sys_clk) begin
	if (main_data_port_we[12])
		data_mem_grain12[main_data_port_adr] <= main_data_port_dat_w[103:96];
	memadr_15 <= main_data_port_adr;
end
assign main_data_port_dat_r[103:96] = data_mem_grain12[memadr_15];
reg [7:0] data_mem_grain13[0:1];
reg [0:0] memadr_16;
always @(posedge sys_clk) begin
	if (main_data_port_we[13])
		data_mem_grain13[main_data_port_adr] <= main_data_port_dat_w[111:104];
	memadr_16 <= main_data_port_adr;
end
assign main_data_port_dat_r[111:104] = data_mem_grain13[memadr_16];
reg [7:0] data_mem_grain14[0:1];
reg [0:0] memadr_17;
always @(posedge sys_clk) begin
	if (main_data_port_we[14])
		data_mem_grain14[main_data_port_adr] <= main_data_port_dat_w[119:112];
	memadr_17 <= main_data_port_adr;
end
assign main_data_port_dat_r[119:112] = data_mem_grain14[memadr_17];
reg [7:0] data_mem_grain15[0:1];
reg [0:0] memadr_18;
always @(posedge sys_clk) begin
	if (main_data_port_we[15])
		data_mem_grain15[main_data_port_adr] <= main_data_port_dat_w[127:120];
	memadr_18 <= main_data_port_adr;
end
assign main_data_port_dat_r[127:120] = data_mem_grain15[memadr_18];
(* ars_ff1 = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE (
	.C(sys_clk),
	.CE(1'd1),
	.D(1'd0),
	.PRE(builder_xilinxasyncresetsynchronizerimpl0),
	.Q(builder_xilinxasyncresetsynchronizerimpl0_rst_meta)
);
(* ars_ff2 = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE_1 (
	.C(sys_clk),
	.CE(1'd1),
	.D(builder_xilinxasyncresetsynchronizerimpl0_rst_meta),
	.PRE(builder_xilinxasyncresetsynchronizerimpl0),
	.Q(sys_rst)
);
(* ars_ff1 = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE_2 (
	.C(sys4x_clk),
	.CE(1'd1),
	.D(1'd0),
	.PRE(builder_xilinxasyncresetsynchronizerimpl1),
	.Q(builder_xilinxasyncresetsynchronizerimpl1_rst_meta)
);
(* ars_ff2 = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE_3 (
	.C(sys4x_clk),
	.CE(1'd1),
	.D(builder_xilinxasyncresetsynchronizerimpl1_rst_meta),
	.PRE(builder_xilinxasyncresetsynchronizerimpl1),
	.Q(builder_xilinxasyncresetsynchronizerimpl1_expr)
);
(* ars_ff1 = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE_4 (
	.C(sys4x_dqs_clk),
	.CE(1'd1),
	.D(1'd0),
	.PRE(builder_xilinxasyncresetsynchronizerimpl2),
	.Q(builder_xilinxasyncresetsynchronizerimpl2_rst_meta)
);
(* ars_ff2 = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE_5 (
	.C(sys4x_dqs_clk),
	.CE(1'd1),
	.D(builder_xilinxasyncresetsynchronizerimpl2_rst_meta),
	.PRE(builder_xilinxasyncresetsynchronizerimpl2),
	.Q(builder_xilinxasyncresetsynchronizerimpl2_expr)
);
(* ars_ff1 = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE_6 (
	.C(clk200_clk),
	.CE(1'd1),
	.D(1'd0),
	.PRE(builder_xilinxasyncresetsynchronizerimpl3),
	.Q(builder_xilinxasyncresetsynchronizerimpl3_rst_meta)
);
(* ars_ff2 = "true", async_reg = "true" *) FDPE #(
	.INIT(1'd1)
) FDPE_7 (
	.C(clk200_clk),
	.CE(1'd1),
	.D(builder_xilinxasyncresetsynchronizerimpl3_rst_meta),
	.PRE(builder_xilinxasyncresetsynchronizerimpl3),
	.Q(clk200_rst)
);
endmodule