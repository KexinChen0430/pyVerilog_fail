module FE #(
`ifdef XIL_TIMING
  parameter LOC = "UNPLACED",
`endif
  parameter MODE = "TURBO_DECODE",
  parameter real PHYSICAL_UTILIZATION = 100.00,
  parameter SIM_DEVICE = "ULTRASCALE_PLUS",
  parameter STANDARD = "LTE",
  parameter real THROUGHPUT_UTILIZATION = 100.00
)(
  output [399:0] DEBUG_DOUT,
  output DEBUG_PHASE,
  output INTERRUPT,
  output [511:0] M_AXIS_DOUT_TDATA,
  output M_AXIS_DOUT_TLAST,
  output M_AXIS_DOUT_TVALID,
  output [31:0] M_AXIS_STATUS_TDATA,
  output M_AXIS_STATUS_TVALID,
  output [15:0] SPARE_OUT,
  output S_AXIS_CTRL_TREADY,
  output S_AXIS_DIN_TREADY,
  output S_AXIS_DIN_WORDS_TREADY,
  output S_AXIS_DOUT_WORDS_TREADY,
  output S_AXI_ARREADY,
  output S_AXI_AWREADY,
  output S_AXI_BVALID,
  output [31:0] S_AXI_RDATA,
  output S_AXI_RVALID,
  output S_AXI_WREADY,
  input CORE_CLK,
  input DEBUG_CLK_EN,
  input DEBUG_EN,
  input [3:0] DEBUG_SEL_IN,
  input M_AXIS_DOUT_ACLK,
  input M_AXIS_DOUT_TREADY,
  input M_AXIS_STATUS_ACLK,
  input M_AXIS_STATUS_TREADY,
  input RESET_N,
  input [15:0] SPARE_IN,
  input S_AXIS_CTRL_ACLK,
  input [31:0] S_AXIS_CTRL_TDATA,
  input S_AXIS_CTRL_TVALID,
  input S_AXIS_DIN_ACLK,
  input [511:0] S_AXIS_DIN_TDATA,
  input S_AXIS_DIN_TLAST,
  input S_AXIS_DIN_TVALID,
  input S_AXIS_DIN_WORDS_ACLK,
  input [31:0] S_AXIS_DIN_WORDS_TDATA,
  input S_AXIS_DIN_WORDS_TLAST,
  input S_AXIS_DIN_WORDS_TVALID,
  input S_AXIS_DOUT_WORDS_ACLK,
  input [31:0] S_AXIS_DOUT_WORDS_TDATA,
  input S_AXIS_DOUT_WORDS_TLAST,
  input S_AXIS_DOUT_WORDS_TVALID,
  input S_AXI_ACLK,
  input [17:0] S_AXI_ARADDR,
  input S_AXI_ARVALID,
  input [17:0] S_AXI_AWADDR,
  input S_AXI_AWVALID,
  input S_AXI_BREADY,
  input S_AXI_RREADY,
  input [31:0] S_AXI_WDATA,
  input S_AXI_WVALID
);
// define constants
  localparam MODULE_NAME = "FE";
  reg trig_attr;
// include dynamic registers - XILINX test only
`ifdef XIL_DR
  `include "FE_dr.v"
`else
  reg [96:1] MODE_REG = MODE;
  real PHYSICAL_UTILIZATION_REG = PHYSICAL_UTILIZATION;
  reg [152:1] SIM_DEVICE_REG = SIM_DEVICE;
  reg [48:1] STANDARD_REG = STANDARD;
  real THROUGHPUT_UTILIZATION_REG = THROUGHPUT_UTILIZATION;
`endif
`ifdef XIL_XECLIB
  wire [63:0] PHYSICAL_UTILIZATION_BIN;
  wire [63:0] THROUGHPUT_UTILIZATION_BIN;
`else
  reg [63:0] PHYSICAL_UTILIZATION_BIN;
  reg [63:0] THROUGHPUT_UTILIZATION_BIN;
`endif
`ifdef XIL_XECLIB
reg glblGSR = 1'b0;
`else
  tri0 glblGSR = glbl.GSR;
`endif
  wire CSSD_CLK_STOP_DONE_out;
  wire DEBUG_PHASE_out;
  wire INTERRUPT_out;
  wire MBIST_COMPSTAT_out;
  wire MBIST_TDO_out;
  wire M_AXIS_DOUT_TLAST_out;
  wire M_AXIS_DOUT_TVALID_out;
  wire M_AXIS_STATUS_TVALID_out;
  wire S_AXIS_CTRL_TREADY_out;
  wire S_AXIS_DIN_TREADY_out;
  wire S_AXIS_DIN_WORDS_TREADY_out;
  wire S_AXIS_DOUT_WORDS_TREADY_out;
  wire S_AXI_ARREADY_out;
  wire S_AXI_AWREADY_out;
  wire S_AXI_BVALID_out;
  wire S_AXI_RVALID_out;
  wire S_AXI_WREADY_out;
  wire [15:0] SPARE_OUT_out;
  wire [199:0] SCANOUT_out;
  wire [31:0] M_AXIS_STATUS_TDATA_out;
  wire [31:0] S_AXI_RDATA_out;
  wire [399:0] DEBUG_DOUT_out;
  wire [511:0] M_AXIS_DOUT_TDATA_out;
  wire [710:0] XIL_UNCONN_OUT_out;
  wire CORE_CLK_in;
  wire CSSD_RST_N_in;
  wire CTL_CSSD_EN_N_in;
  wire CTL_CSSD_SNGL_CHAIN_MD_N_in;
  wire DEBUG_CLK_EN_in;
  wire DEBUG_EN_in;
  wire DFTRAM_BYPASS_N_in;
  wire MBIST_TCK_in;
  wire MBIST_TDI_in;
  wire MBIST_TMS_in;
  wire MBIST_TRST_in;
  wire M_AXIS_DOUT_ACLK_in;
  wire M_AXIS_DOUT_TREADY_in;
  wire M_AXIS_STATUS_ACLK_in;
  wire M_AXIS_STATUS_TREADY_in;
  wire RESET_N_in;
  wire SCANENABLE_N_in;
  wire SCANMODE_N_in;
  wire SCAN_CLK_in;
  wire S_AXIS_CTRL_ACLK_in;
  wire S_AXIS_CTRL_TVALID_in;
  wire S_AXIS_DIN_ACLK_in;
  wire S_AXIS_DIN_TLAST_in;
  wire S_AXIS_DIN_TVALID_in;
  wire S_AXIS_DIN_WORDS_ACLK_in;
  wire S_AXIS_DIN_WORDS_TLAST_in;
  wire S_AXIS_DIN_WORDS_TVALID_in;
  wire S_AXIS_DOUT_WORDS_ACLK_in;
  wire S_AXIS_DOUT_WORDS_TLAST_in;
  wire S_AXIS_DOUT_WORDS_TVALID_in;
  wire S_AXI_ACLK_in;
  wire S_AXI_ARVALID_in;
  wire S_AXI_AWVALID_in;
  wire S_AXI_BREADY_in;
  wire S_AXI_RREADY_in;
  wire S_AXI_WVALID_in;
  wire TEST_MODE_PIN_CHAR_N_in;
  wire [15:0] CTL_CSSD_MRKR_START_INIT_in;
  wire [15:0] CTL_CSSD_MRKR_STOP_INIT_in;
  wire [15:0] SPARE_IN_in;
  wire [17:0] S_AXI_ARADDR_in;
  wire [17:0] S_AXI_AWADDR_in;
  wire [1861:0] XIL_UNCONN_IN_in;
  wire [199:0] SCANIN_in;
  wire [2:0] CTL_CSSD_ROOT_CLK_SEL_in;
  wire [31:0] S_AXIS_CTRL_TDATA_in;
  wire [31:0] S_AXIS_DIN_WORDS_TDATA_in;
  wire [31:0] S_AXIS_DOUT_WORDS_TDATA_in;
  wire [31:0] S_AXI_WDATA_in;
  wire [3:0] CSSD_CLK_STOP_EVENT_in;
  wire [3:0] DEBUG_SEL_IN_in;
  wire [469:0] XIL_UNCONN_CLK_in;
  wire [47:0] CTL_CSSD_STOP_COUNT_in;
  wire [511:0] S_AXIS_DIN_TDATA_in;
  wire [7:0] CTL_CSSD_ROOT_CLK_DIS_in;
`ifdef XIL_TIMING
  wire CORE_CLK_delay;
  wire DEBUG_EN_delay;
  wire M_AXIS_DOUT_ACLK_delay;
  wire M_AXIS_DOUT_TREADY_delay;
  wire M_AXIS_STATUS_ACLK_delay;
  wire M_AXIS_STATUS_TREADY_delay;
  wire S_AXIS_CTRL_ACLK_delay;
  wire S_AXIS_CTRL_TVALID_delay;
  wire S_AXIS_DIN_ACLK_delay;
  wire S_AXIS_DIN_TLAST_delay;
  wire S_AXIS_DIN_TVALID_delay;
  wire S_AXIS_DIN_WORDS_ACLK_delay;
  wire S_AXIS_DIN_WORDS_TLAST_delay;
  wire S_AXIS_DIN_WORDS_TVALID_delay;
  wire S_AXIS_DOUT_WORDS_ACLK_delay;
  wire S_AXIS_DOUT_WORDS_TLAST_delay;
  wire S_AXIS_DOUT_WORDS_TVALID_delay;
  wire S_AXI_ACLK_delay;
  wire S_AXI_ARVALID_delay;
  wire S_AXI_AWVALID_delay;
  wire S_AXI_BREADY_delay;
  wire S_AXI_RREADY_delay;
  wire S_AXI_WVALID_delay;
  wire [17:0] S_AXI_ARADDR_delay;
  wire [17:0] S_AXI_AWADDR_delay;
  wire [31:0] S_AXIS_CTRL_TDATA_delay;
  wire [31:0] S_AXIS_DIN_WORDS_TDATA_delay;
  wire [31:0] S_AXIS_DOUT_WORDS_TDATA_delay;
  wire [31:0] S_AXI_WDATA_delay;
  wire [511:0] S_AXIS_DIN_TDATA_delay;
`endif
  assign DEBUG_DOUT = DEBUG_DOUT_out;
  assign DEBUG_PHASE = DEBUG_PHASE_out;
  assign INTERRUPT = INTERRUPT_out;
  assign M_AXIS_DOUT_TDATA = M_AXIS_DOUT_TDATA_out;
  assign M_AXIS_DOUT_TLAST = M_AXIS_DOUT_TLAST_out;
  assign M_AXIS_DOUT_TVALID = M_AXIS_DOUT_TVALID_out;
  assign M_AXIS_STATUS_TDATA = M_AXIS_STATUS_TDATA_out;
  assign M_AXIS_STATUS_TVALID = M_AXIS_STATUS_TVALID_out;
  assign SPARE_OUT = SPARE_OUT_out;
  assign S_AXIS_CTRL_TREADY = S_AXIS_CTRL_TREADY_out;
  assign S_AXIS_DIN_TREADY = S_AXIS_DIN_TREADY_out;
  assign S_AXIS_DIN_WORDS_TREADY = S_AXIS_DIN_WORDS_TREADY_out;
  assign S_AXIS_DOUT_WORDS_TREADY = S_AXIS_DOUT_WORDS_TREADY_out;
  assign S_AXI_ARREADY = S_AXI_ARREADY_out;
  assign S_AXI_AWREADY = S_AXI_AWREADY_out;
  assign S_AXI_BVALID = S_AXI_BVALID_out;
  assign S_AXI_RDATA = S_AXI_RDATA_out;
  assign S_AXI_RVALID = S_AXI_RVALID_out;
  assign S_AXI_WREADY = S_AXI_WREADY_out;
`ifdef XIL_TIMING
  assign CORE_CLK_in = (CORE_CLK !== 1'bz) && CORE_CLK_delay; // rv 0
  assign DEBUG_EN_in = (DEBUG_EN === 1'bz) || DEBUG_EN_delay; // rv 1
  assign M_AXIS_DOUT_ACLK_in = (M_AXIS_DOUT_ACLK !== 1'bz) && M_AXIS_DOUT_ACLK_delay; // rv 0
  assign M_AXIS_DOUT_TREADY_in = (M_AXIS_DOUT_TREADY !== 1'bz) && M_AXIS_DOUT_TREADY_delay; // rv 0
  assign M_AXIS_STATUS_ACLK_in = (M_AXIS_STATUS_ACLK !== 1'bz) && M_AXIS_STATUS_ACLK_delay; // rv 0
  assign M_AXIS_STATUS_TREADY_in = (M_AXIS_STATUS_TREADY !== 1'bz) && M_AXIS_STATUS_TREADY_delay; // rv 0
  assign S_AXIS_CTRL_ACLK_in = (S_AXIS_CTRL_ACLK !== 1'bz) && S_AXIS_CTRL_ACLK_delay; // rv 0
  assign S_AXIS_CTRL_TDATA_in[0] = (S_AXIS_CTRL_TDATA[0] !== 1'bz) && S_AXIS_CTRL_TDATA_delay[0]; // rv 0
  assign S_AXIS_CTRL_TDATA_in[10] = (S_AXIS_CTRL_TDATA[10] !== 1'bz) && S_AXIS_CTRL_TDATA_delay[10]; // rv 0
  assign S_AXIS_CTRL_TDATA_in[11] = (S_AXIS_CTRL_TDATA[11] !== 1'bz) && S_AXIS_CTRL_TDATA_delay[11]; // rv 0
  assign S_AXIS_CTRL_TDATA_in[12] = (S_AXIS_CTRL_TDATA[12] !== 1'bz) && S_AXIS_CTRL_TDATA_delay[12]; // rv 0
  assign S_AXIS_CTRL_TDATA_in[13] = (S_AXIS_CTRL_TDATA[13] !== 1'bz) && S_AXIS_CTRL_TDATA_delay[13]; // rv 0
  assign S_AXIS_CTRL_TDATA_in[14] = (S_AXIS_CTRL_TDATA[14] !== 1'bz) && S_AXIS_CTRL_TDATA_delay[14]; // rv 0
  assign S_AXIS_CTRL_TDATA_in[15] = (S_AXIS_CTRL_TDATA[15] !== 1'bz) && S_AXIS_CTRL_TDATA_delay[15]; // rv 0
  assign S_AXIS_CTRL_TDATA_in[16] = (S_AXIS_CTRL_TDATA[16] !== 1'bz) && S_AXIS_CTRL_TDATA_delay[16]; // rv 0
  assign S_AXIS_CTRL_TDATA_in[17] = (S_AXIS_CTRL_TDATA[17] !== 1'bz) && S_AXIS_CTRL_TDATA_delay[17]; // rv 0
  assign S_AXIS_CTRL_TDATA_in[18] = (S_AXIS_CTRL_TDATA[18] !== 1'bz) && S_AXIS_CTRL_TDATA_delay[18]; // rv 0
  assign S_AXIS_CTRL_TDATA_in[19] = (S_AXIS_CTRL_TDATA[19] !== 1'bz) && S_AXIS_CTRL_TDATA_delay[19]; // rv 0
  assign S_AXIS_CTRL_TDATA_in[1] = (S_AXIS_CTRL_TDATA[1] !== 1'bz) && S_AXIS_CTRL_TDATA_delay[1]; // rv 0
  assign S_AXIS_CTRL_TDATA_in[20] = (S_AXIS_CTRL_TDATA[20] !== 1'bz) && S_AXIS_CTRL_TDATA_delay[20]; // rv 0
  assign S_AXIS_CTRL_TDATA_in[21] = (S_AXIS_CTRL_TDATA[21] !== 1'bz) && S_AXIS_CTRL_TDATA_delay[21]; // rv 0
  assign S_AXIS_CTRL_TDATA_in[22] = (S_AXIS_CTRL_TDATA[22] !== 1'bz) && S_AXIS_CTRL_TDATA_delay[22]; // rv 0
  assign S_AXIS_CTRL_TDATA_in[23] = (S_AXIS_CTRL_TDATA[23] !== 1'bz) && S_AXIS_CTRL_TDATA_delay[23]; // rv 0
  assign S_AXIS_CTRL_TDATA_in[24] = (S_AXIS_CTRL_TDATA[24] !== 1'bz) && S_AXIS_CTRL_TDATA_delay[24]; // rv 0
  assign S_AXIS_CTRL_TDATA_in[25] = (S_AXIS_CTRL_TDATA[25] !== 1'bz) && S_AXIS_CTRL_TDATA_delay[25]; // rv 0
  assign S_AXIS_CTRL_TDATA_in[26] = (S_AXIS_CTRL_TDATA[26] !== 1'bz) && S_AXIS_CTRL_TDATA_delay[26]; // rv 0
  assign S_AXIS_CTRL_TDATA_in[27] = (S_AXIS_CTRL_TDATA[27] !== 1'bz) && S_AXIS_CTRL_TDATA_delay[27]; // rv 0
  assign S_AXIS_CTRL_TDATA_in[28] = (S_AXIS_CTRL_TDATA[28] !== 1'bz) && S_AXIS_CTRL_TDATA_delay[28]; // rv 0
  assign S_AXIS_CTRL_TDATA_in[29] = (S_AXIS_CTRL_TDATA[29] !== 1'bz) && S_AXIS_CTRL_TDATA_delay[29]; // rv 0
  assign S_AXIS_CTRL_TDATA_in[2] = (S_AXIS_CTRL_TDATA[2] !== 1'bz) && S_AXIS_CTRL_TDATA_delay[2]; // rv 0
  assign S_AXIS_CTRL_TDATA_in[30] = (S_AXIS_CTRL_TDATA[30] !== 1'bz) && S_AXIS_CTRL_TDATA_delay[30]; // rv 0
  assign S_AXIS_CTRL_TDATA_in[31] = (S_AXIS_CTRL_TDATA[31] !== 1'bz) && S_AXIS_CTRL_TDATA_delay[31]; // rv 0
  assign S_AXIS_CTRL_TDATA_in[3] = (S_AXIS_CTRL_TDATA[3] !== 1'bz) && S_AXIS_CTRL_TDATA_delay[3]; // rv 0
  assign S_AXIS_CTRL_TDATA_in[4] = (S_AXIS_CTRL_TDATA[4] !== 1'bz) && S_AXIS_CTRL_TDATA_delay[4]; // rv 0
  assign S_AXIS_CTRL_TDATA_in[5] = (S_AXIS_CTRL_TDATA[5] !== 1'bz) && S_AXIS_CTRL_TDATA_delay[5]; // rv 0
  assign S_AXIS_CTRL_TDATA_in[6] = (S_AXIS_CTRL_TDATA[6] !== 1'bz) && S_AXIS_CTRL_TDATA_delay[6]; // rv 0
  assign S_AXIS_CTRL_TDATA_in[7] = (S_AXIS_CTRL_TDATA[7] !== 1'bz) && S_AXIS_CTRL_TDATA_delay[7]; // rv 0
  assign S_AXIS_CTRL_TDATA_in[8] = (S_AXIS_CTRL_TDATA[8] !== 1'bz) && S_AXIS_CTRL_TDATA_delay[8]; // rv 0
  assign S_AXIS_CTRL_TDATA_in[9] = (S_AXIS_CTRL_TDATA[9] !== 1'bz) && S_AXIS_CTRL_TDATA_delay[9]; // rv 0
  assign S_AXIS_CTRL_TVALID_in = (S_AXIS_CTRL_TVALID !== 1'bz) && S_AXIS_CTRL_TVALID_delay; // rv 0
  assign S_AXIS_DIN_ACLK_in = (S_AXIS_DIN_ACLK !== 1'bz) && S_AXIS_DIN_ACLK_delay; // rv 0
  assign S_AXIS_DIN_TDATA_in[0] = (S_AXIS_DIN_TDATA[0] !== 1'bz) && S_AXIS_DIN_TDATA_delay[0]; // rv 0
  assign S_AXIS_DIN_TDATA_in[100] = (S_AXIS_DIN_TDATA[100] !== 1'bz) && S_AXIS_DIN_TDATA_delay[100]; // rv 0
  assign S_AXIS_DIN_TDATA_in[101] = (S_AXIS_DIN_TDATA[101] !== 1'bz) && S_AXIS_DIN_TDATA_delay[101]; // rv 0
  assign S_AXIS_DIN_TDATA_in[102] = (S_AXIS_DIN_TDATA[102] !== 1'bz) && S_AXIS_DIN_TDATA_delay[102]; // rv 0
  assign S_AXIS_DIN_TDATA_in[103] = (S_AXIS_DIN_TDATA[103] !== 1'bz) && S_AXIS_DIN_TDATA_delay[103]; // rv 0
  assign S_AXIS_DIN_TDATA_in[104] = (S_AXIS_DIN_TDATA[104] !== 1'bz) && S_AXIS_DIN_TDATA_delay[104]; // rv 0
  assign S_AXIS_DIN_TDATA_in[105] = (S_AXIS_DIN_TDATA[105] !== 1'bz) && S_AXIS_DIN_TDATA_delay[105]; // rv 0
  assign S_AXIS_DIN_TDATA_in[106] = (S_AXIS_DIN_TDATA[106] !== 1'bz) && S_AXIS_DIN_TDATA_delay[106]; // rv 0
  assign S_AXIS_DIN_TDATA_in[107] = (S_AXIS_DIN_TDATA[107] !== 1'bz) && S_AXIS_DIN_TDATA_delay[107]; // rv 0
  assign S_AXIS_DIN_TDATA_in[108] = (S_AXIS_DIN_TDATA[108] !== 1'bz) && S_AXIS_DIN_TDATA_delay[108]; // rv 0
  assign S_AXIS_DIN_TDATA_in[109] = (S_AXIS_DIN_TDATA[109] !== 1'bz) && S_AXIS_DIN_TDATA_delay[109]; // rv 0
  assign S_AXIS_DIN_TDATA_in[10] = (S_AXIS_DIN_TDATA[10] !== 1'bz) && S_AXIS_DIN_TDATA_delay[10]; // rv 0
  assign S_AXIS_DIN_TDATA_in[110] = (S_AXIS_DIN_TDATA[110] !== 1'bz) && S_AXIS_DIN_TDATA_delay[110]; // rv 0
  assign S_AXIS_DIN_TDATA_in[111] = (S_AXIS_DIN_TDATA[111] !== 1'bz) && S_AXIS_DIN_TDATA_delay[111]; // rv 0
  assign S_AXIS_DIN_TDATA_in[112] = (S_AXIS_DIN_TDATA[112] !== 1'bz) && S_AXIS_DIN_TDATA_delay[112]; // rv 0
  assign S_AXIS_DIN_TDATA_in[113] = (S_AXIS_DIN_TDATA[113] !== 1'bz) && S_AXIS_DIN_TDATA_delay[113]; // rv 0
  assign S_AXIS_DIN_TDATA_in[114] = (S_AXIS_DIN_TDATA[114] !== 1'bz) && S_AXIS_DIN_TDATA_delay[114]; // rv 0
  assign S_AXIS_DIN_TDATA_in[115] = (S_AXIS_DIN_TDATA[115] !== 1'bz) && S_AXIS_DIN_TDATA_delay[115]; // rv 0
  assign S_AXIS_DIN_TDATA_in[116] = (S_AXIS_DIN_TDATA[116] !== 1'bz) && S_AXIS_DIN_TDATA_delay[116]; // rv 0
  assign S_AXIS_DIN_TDATA_in[117] = (S_AXIS_DIN_TDATA[117] !== 1'bz) && S_AXIS_DIN_TDATA_delay[117]; // rv 0
  assign S_AXIS_DIN_TDATA_in[118] = (S_AXIS_DIN_TDATA[118] !== 1'bz) && S_AXIS_DIN_TDATA_delay[118]; // rv 0
  assign S_AXIS_DIN_TDATA_in[119] = (S_AXIS_DIN_TDATA[119] !== 1'bz) && S_AXIS_DIN_TDATA_delay[119]; // rv 0
  assign S_AXIS_DIN_TDATA_in[11] = (S_AXIS_DIN_TDATA[11] !== 1'bz) && S_AXIS_DIN_TDATA_delay[11]; // rv 0
  assign S_AXIS_DIN_TDATA_in[120] = (S_AXIS_DIN_TDATA[120] !== 1'bz) && S_AXIS_DIN_TDATA_delay[120]; // rv 0
  assign S_AXIS_DIN_TDATA_in[121] = (S_AXIS_DIN_TDATA[121] !== 1'bz) && S_AXIS_DIN_TDATA_delay[121]; // rv 0
  assign S_AXIS_DIN_TDATA_in[122] = (S_AXIS_DIN_TDATA[122] !== 1'bz) && S_AXIS_DIN_TDATA_delay[122]; // rv 0
  assign S_AXIS_DIN_TDATA_in[123] = (S_AXIS_DIN_TDATA[123] !== 1'bz) && S_AXIS_DIN_TDATA_delay[123]; // rv 0
  assign S_AXIS_DIN_TDATA_in[124] = (S_AXIS_DIN_TDATA[124] !== 1'bz) && S_AXIS_DIN_TDATA_delay[124]; // rv 0
  assign S_AXIS_DIN_TDATA_in[125] = (S_AXIS_DIN_TDATA[125] !== 1'bz) && S_AXIS_DIN_TDATA_delay[125]; // rv 0
  assign S_AXIS_DIN_TDATA_in[126] = (S_AXIS_DIN_TDATA[126] !== 1'bz) && S_AXIS_DIN_TDATA_delay[126]; // rv 0
  assign S_AXIS_DIN_TDATA_in[127] = (S_AXIS_DIN_TDATA[127] !== 1'bz) && S_AXIS_DIN_TDATA_delay[127]; // rv 0
  assign S_AXIS_DIN_TDATA_in[128] = (S_AXIS_DIN_TDATA[128] !== 1'bz) && S_AXIS_DIN_TDATA_delay[128]; // rv 0
  assign S_AXIS_DIN_TDATA_in[129] = (S_AXIS_DIN_TDATA[129] !== 1'bz) && S_AXIS_DIN_TDATA_delay[129]; // rv 0
  assign S_AXIS_DIN_TDATA_in[12] = (S_AXIS_DIN_TDATA[12] !== 1'bz) && S_AXIS_DIN_TDATA_delay[12]; // rv 0
  assign S_AXIS_DIN_TDATA_in[130] = (S_AXIS_DIN_TDATA[130] !== 1'bz) && S_AXIS_DIN_TDATA_delay[130]; // rv 0
  assign S_AXIS_DIN_TDATA_in[131] = (S_AXIS_DIN_TDATA[131] !== 1'bz) && S_AXIS_DIN_TDATA_delay[131]; // rv 0
  assign S_AXIS_DIN_TDATA_in[132] = (S_AXIS_DIN_TDATA[132] !== 1'bz) && S_AXIS_DIN_TDATA_delay[132]; // rv 0
  assign S_AXIS_DIN_TDATA_in[133] = (S_AXIS_DIN_TDATA[133] !== 1'bz) && S_AXIS_DIN_TDATA_delay[133]; // rv 0
  assign S_AXIS_DIN_TDATA_in[134] = (S_AXIS_DIN_TDATA[134] !== 1'bz) && S_AXIS_DIN_TDATA_delay[134]; // rv 0
  assign S_AXIS_DIN_TDATA_in[135] = (S_AXIS_DIN_TDATA[135] !== 1'bz) && S_AXIS_DIN_TDATA_delay[135]; // rv 0
  assign S_AXIS_DIN_TDATA_in[136] = (S_AXIS_DIN_TDATA[136] !== 1'bz) && S_AXIS_DIN_TDATA_delay[136]; // rv 0
  assign S_AXIS_DIN_TDATA_in[137] = (S_AXIS_DIN_TDATA[137] !== 1'bz) && S_AXIS_DIN_TDATA_delay[137]; // rv 0
  assign S_AXIS_DIN_TDATA_in[138] = (S_AXIS_DIN_TDATA[138] !== 1'bz) && S_AXIS_DIN_TDATA_delay[138]; // rv 0
  assign S_AXIS_DIN_TDATA_in[139] = (S_AXIS_DIN_TDATA[139] !== 1'bz) && S_AXIS_DIN_TDATA_delay[139]; // rv 0
  assign S_AXIS_DIN_TDATA_in[13] = (S_AXIS_DIN_TDATA[13] !== 1'bz) && S_AXIS_DIN_TDATA_delay[13]; // rv 0
  assign S_AXIS_DIN_TDATA_in[140] = (S_AXIS_DIN_TDATA[140] !== 1'bz) && S_AXIS_DIN_TDATA_delay[140]; // rv 0
  assign S_AXIS_DIN_TDATA_in[141] = (S_AXIS_DIN_TDATA[141] !== 1'bz) && S_AXIS_DIN_TDATA_delay[141]; // rv 0
  assign S_AXIS_DIN_TDATA_in[142] = (S_AXIS_DIN_TDATA[142] !== 1'bz) && S_AXIS_DIN_TDATA_delay[142]; // rv 0
  assign S_AXIS_DIN_TDATA_in[143] = (S_AXIS_DIN_TDATA[143] !== 1'bz) && S_AXIS_DIN_TDATA_delay[143]; // rv 0
  assign S_AXIS_DIN_TDATA_in[144] = (S_AXIS_DIN_TDATA[144] !== 1'bz) && S_AXIS_DIN_TDATA_delay[144]; // rv 0
  assign S_AXIS_DIN_TDATA_in[145] = (S_AXIS_DIN_TDATA[145] !== 1'bz) && S_AXIS_DIN_TDATA_delay[145]; // rv 0
  assign S_AXIS_DIN_TDATA_in[146] = (S_AXIS_DIN_TDATA[146] !== 1'bz) && S_AXIS_DIN_TDATA_delay[146]; // rv 0
  assign S_AXIS_DIN_TDATA_in[147] = (S_AXIS_DIN_TDATA[147] !== 1'bz) && S_AXIS_DIN_TDATA_delay[147]; // rv 0
  assign S_AXIS_DIN_TDATA_in[148] = (S_AXIS_DIN_TDATA[148] !== 1'bz) && S_AXIS_DIN_TDATA_delay[148]; // rv 0
  assign S_AXIS_DIN_TDATA_in[149] = (S_AXIS_DIN_TDATA[149] !== 1'bz) && S_AXIS_DIN_TDATA_delay[149]; // rv 0
  assign S_AXIS_DIN_TDATA_in[14] = (S_AXIS_DIN_TDATA[14] !== 1'bz) && S_AXIS_DIN_TDATA_delay[14]; // rv 0
  assign S_AXIS_DIN_TDATA_in[150] = (S_AXIS_DIN_TDATA[150] !== 1'bz) && S_AXIS_DIN_TDATA_delay[150]; // rv 0
  assign S_AXIS_DIN_TDATA_in[151] = (S_AXIS_DIN_TDATA[151] !== 1'bz) && S_AXIS_DIN_TDATA_delay[151]; // rv 0
  assign S_AXIS_DIN_TDATA_in[152] = (S_AXIS_DIN_TDATA[152] !== 1'bz) && S_AXIS_DIN_TDATA_delay[152]; // rv 0
  assign S_AXIS_DIN_TDATA_in[153] = (S_AXIS_DIN_TDATA[153] !== 1'bz) && S_AXIS_DIN_TDATA_delay[153]; // rv 0
  assign S_AXIS_DIN_TDATA_in[154] = (S_AXIS_DIN_TDATA[154] !== 1'bz) && S_AXIS_DIN_TDATA_delay[154]; // rv 0
  assign S_AXIS_DIN_TDATA_in[155] = (S_AXIS_DIN_TDATA[155] !== 1'bz) && S_AXIS_DIN_TDATA_delay[155]; // rv 0
  assign S_AXIS_DIN_TDATA_in[156] = (S_AXIS_DIN_TDATA[156] !== 1'bz) && S_AXIS_DIN_TDATA_delay[156]; // rv 0
  assign S_AXIS_DIN_TDATA_in[157] = (S_AXIS_DIN_TDATA[157] !== 1'bz) && S_AXIS_DIN_TDATA_delay[157]; // rv 0
  assign S_AXIS_DIN_TDATA_in[158] = (S_AXIS_DIN_TDATA[158] !== 1'bz) && S_AXIS_DIN_TDATA_delay[158]; // rv 0
  assign S_AXIS_DIN_TDATA_in[159] = (S_AXIS_DIN_TDATA[159] !== 1'bz) && S_AXIS_DIN_TDATA_delay[159]; // rv 0
  assign S_AXIS_DIN_TDATA_in[15] = (S_AXIS_DIN_TDATA[15] !== 1'bz) && S_AXIS_DIN_TDATA_delay[15]; // rv 0
  assign S_AXIS_DIN_TDATA_in[160] = (S_AXIS_DIN_TDATA[160] !== 1'bz) && S_AXIS_DIN_TDATA_delay[160]; // rv 0
  assign S_AXIS_DIN_TDATA_in[161] = (S_AXIS_DIN_TDATA[161] !== 1'bz) && S_AXIS_DIN_TDATA_delay[161]; // rv 0
  assign S_AXIS_DIN_TDATA_in[162] = (S_AXIS_DIN_TDATA[162] !== 1'bz) && S_AXIS_DIN_TDATA_delay[162]; // rv 0
  assign S_AXIS_DIN_TDATA_in[163] = (S_AXIS_DIN_TDATA[163] !== 1'bz) && S_AXIS_DIN_TDATA_delay[163]; // rv 0
  assign S_AXIS_DIN_TDATA_in[164] = (S_AXIS_DIN_TDATA[164] !== 1'bz) && S_AXIS_DIN_TDATA_delay[164]; // rv 0
  assign S_AXIS_DIN_TDATA_in[165] = (S_AXIS_DIN_TDATA[165] !== 1'bz) && S_AXIS_DIN_TDATA_delay[165]; // rv 0
  assign S_AXIS_DIN_TDATA_in[166] = (S_AXIS_DIN_TDATA[166] !== 1'bz) && S_AXIS_DIN_TDATA_delay[166]; // rv 0
  assign S_AXIS_DIN_TDATA_in[167] = (S_AXIS_DIN_TDATA[167] !== 1'bz) && S_AXIS_DIN_TDATA_delay[167]; // rv 0
  assign S_AXIS_DIN_TDATA_in[168] = (S_AXIS_DIN_TDATA[168] !== 1'bz) && S_AXIS_DIN_TDATA_delay[168]; // rv 0
  assign S_AXIS_DIN_TDATA_in[169] = (S_AXIS_DIN_TDATA[169] !== 1'bz) && S_AXIS_DIN_TDATA_delay[169]; // rv 0
  assign S_AXIS_DIN_TDATA_in[16] = (S_AXIS_DIN_TDATA[16] !== 1'bz) && S_AXIS_DIN_TDATA_delay[16]; // rv 0
  assign S_AXIS_DIN_TDATA_in[170] = (S_AXIS_DIN_TDATA[170] !== 1'bz) && S_AXIS_DIN_TDATA_delay[170]; // rv 0
  assign S_AXIS_DIN_TDATA_in[171] = (S_AXIS_DIN_TDATA[171] !== 1'bz) && S_AXIS_DIN_TDATA_delay[171]; // rv 0
  assign S_AXIS_DIN_TDATA_in[172] = (S_AXIS_DIN_TDATA[172] !== 1'bz) && S_AXIS_DIN_TDATA_delay[172]; // rv 0
  assign S_AXIS_DIN_TDATA_in[173] = (S_AXIS_DIN_TDATA[173] !== 1'bz) && S_AXIS_DIN_TDATA_delay[173]; // rv 0
  assign S_AXIS_DIN_TDATA_in[174] = (S_AXIS_DIN_TDATA[174] !== 1'bz) && S_AXIS_DIN_TDATA_delay[174]; // rv 0
  assign S_AXIS_DIN_TDATA_in[175] = (S_AXIS_DIN_TDATA[175] !== 1'bz) && S_AXIS_DIN_TDATA_delay[175]; // rv 0
  assign S_AXIS_DIN_TDATA_in[176] = (S_AXIS_DIN_TDATA[176] !== 1'bz) && S_AXIS_DIN_TDATA_delay[176]; // rv 0
  assign S_AXIS_DIN_TDATA_in[177] = (S_AXIS_DIN_TDATA[177] !== 1'bz) && S_AXIS_DIN_TDATA_delay[177]; // rv 0
  assign S_AXIS_DIN_TDATA_in[178] = (S_AXIS_DIN_TDATA[178] !== 1'bz) && S_AXIS_DIN_TDATA_delay[178]; // rv 0
  assign S_AXIS_DIN_TDATA_in[179] = (S_AXIS_DIN_TDATA[179] !== 1'bz) && S_AXIS_DIN_TDATA_delay[179]; // rv 0
  assign S_AXIS_DIN_TDATA_in[17] = (S_AXIS_DIN_TDATA[17] !== 1'bz) && S_AXIS_DIN_TDATA_delay[17]; // rv 0
  assign S_AXIS_DIN_TDATA_in[180] = (S_AXIS_DIN_TDATA[180] !== 1'bz) && S_AXIS_DIN_TDATA_delay[180]; // rv 0
  assign S_AXIS_DIN_TDATA_in[181] = (S_AXIS_DIN_TDATA[181] !== 1'bz) && S_AXIS_DIN_TDATA_delay[181]; // rv 0
  assign S_AXIS_DIN_TDATA_in[182] = (S_AXIS_DIN_TDATA[182] !== 1'bz) && S_AXIS_DIN_TDATA_delay[182]; // rv 0
  assign S_AXIS_DIN_TDATA_in[183] = (S_AXIS_DIN_TDATA[183] !== 1'bz) && S_AXIS_DIN_TDATA_delay[183]; // rv 0
  assign S_AXIS_DIN_TDATA_in[184] = (S_AXIS_DIN_TDATA[184] !== 1'bz) && S_AXIS_DIN_TDATA_delay[184]; // rv 0
  assign S_AXIS_DIN_TDATA_in[185] = (S_AXIS_DIN_TDATA[185] !== 1'bz) && S_AXIS_DIN_TDATA_delay[185]; // rv 0
  assign S_AXIS_DIN_TDATA_in[186] = (S_AXIS_DIN_TDATA[186] !== 1'bz) && S_AXIS_DIN_TDATA_delay[186]; // rv 0
  assign S_AXIS_DIN_TDATA_in[187] = (S_AXIS_DIN_TDATA[187] !== 1'bz) && S_AXIS_DIN_TDATA_delay[187]; // rv 0
  assign S_AXIS_DIN_TDATA_in[188] = (S_AXIS_DIN_TDATA[188] !== 1'bz) && S_AXIS_DIN_TDATA_delay[188]; // rv 0
  assign S_AXIS_DIN_TDATA_in[189] = (S_AXIS_DIN_TDATA[189] !== 1'bz) && S_AXIS_DIN_TDATA_delay[189]; // rv 0
  assign S_AXIS_DIN_TDATA_in[18] = (S_AXIS_DIN_TDATA[18] !== 1'bz) && S_AXIS_DIN_TDATA_delay[18]; // rv 0
  assign S_AXIS_DIN_TDATA_in[190] = (S_AXIS_DIN_TDATA[190] !== 1'bz) && S_AXIS_DIN_TDATA_delay[190]; // rv 0
  assign S_AXIS_DIN_TDATA_in[191] = (S_AXIS_DIN_TDATA[191] !== 1'bz) && S_AXIS_DIN_TDATA_delay[191]; // rv 0
  assign S_AXIS_DIN_TDATA_in[192] = (S_AXIS_DIN_TDATA[192] !== 1'bz) && S_AXIS_DIN_TDATA_delay[192]; // rv 0
  assign S_AXIS_DIN_TDATA_in[193] = (S_AXIS_DIN_TDATA[193] !== 1'bz) && S_AXIS_DIN_TDATA_delay[193]; // rv 0
  assign S_AXIS_DIN_TDATA_in[194] = (S_AXIS_DIN_TDATA[194] !== 1'bz) && S_AXIS_DIN_TDATA_delay[194]; // rv 0
  assign S_AXIS_DIN_TDATA_in[195] = (S_AXIS_DIN_TDATA[195] !== 1'bz) && S_AXIS_DIN_TDATA_delay[195]; // rv 0
  assign S_AXIS_DIN_TDATA_in[196] = (S_AXIS_DIN_TDATA[196] !== 1'bz) && S_AXIS_DIN_TDATA_delay[196]; // rv 0
  assign S_AXIS_DIN_TDATA_in[197] = (S_AXIS_DIN_TDATA[197] !== 1'bz) && S_AXIS_DIN_TDATA_delay[197]; // rv 0
  assign S_AXIS_DIN_TDATA_in[198] = (S_AXIS_DIN_TDATA[198] !== 1'bz) && S_AXIS_DIN_TDATA_delay[198]; // rv 0
  assign S_AXIS_DIN_TDATA_in[199] = (S_AXIS_DIN_TDATA[199] !== 1'bz) && S_AXIS_DIN_TDATA_delay[199]; // rv 0
  assign S_AXIS_DIN_TDATA_in[19] = (S_AXIS_DIN_TDATA[19] !== 1'bz) && S_AXIS_DIN_TDATA_delay[19]; // rv 0
  assign S_AXIS_DIN_TDATA_in[1] = (S_AXIS_DIN_TDATA[1] !== 1'bz) && S_AXIS_DIN_TDATA_delay[1]; // rv 0
  assign S_AXIS_DIN_TDATA_in[200] = (S_AXIS_DIN_TDATA[200] !== 1'bz) && S_AXIS_DIN_TDATA_delay[200]; // rv 0
  assign S_AXIS_DIN_TDATA_in[201] = (S_AXIS_DIN_TDATA[201] !== 1'bz) && S_AXIS_DIN_TDATA_delay[201]; // rv 0
  assign S_AXIS_DIN_TDATA_in[202] = (S_AXIS_DIN_TDATA[202] !== 1'bz) && S_AXIS_DIN_TDATA_delay[202]; // rv 0
  assign S_AXIS_DIN_TDATA_in[203] = (S_AXIS_DIN_TDATA[203] !== 1'bz) && S_AXIS_DIN_TDATA_delay[203]; // rv 0
  assign S_AXIS_DIN_TDATA_in[204] = (S_AXIS_DIN_TDATA[204] !== 1'bz) && S_AXIS_DIN_TDATA_delay[204]; // rv 0
  assign S_AXIS_DIN_TDATA_in[205] = (S_AXIS_DIN_TDATA[205] !== 1'bz) && S_AXIS_DIN_TDATA_delay[205]; // rv 0
  assign S_AXIS_DIN_TDATA_in[206] = (S_AXIS_DIN_TDATA[206] !== 1'bz) && S_AXIS_DIN_TDATA_delay[206]; // rv 0
  assign S_AXIS_DIN_TDATA_in[207] = (S_AXIS_DIN_TDATA[207] !== 1'bz) && S_AXIS_DIN_TDATA_delay[207]; // rv 0
  assign S_AXIS_DIN_TDATA_in[208] = (S_AXIS_DIN_TDATA[208] !== 1'bz) && S_AXIS_DIN_TDATA_delay[208]; // rv 0
  assign S_AXIS_DIN_TDATA_in[209] = (S_AXIS_DIN_TDATA[209] !== 1'bz) && S_AXIS_DIN_TDATA_delay[209]; // rv 0
  assign S_AXIS_DIN_TDATA_in[20] = (S_AXIS_DIN_TDATA[20] !== 1'bz) && S_AXIS_DIN_TDATA_delay[20]; // rv 0
  assign S_AXIS_DIN_TDATA_in[210] = (S_AXIS_DIN_TDATA[210] !== 1'bz) && S_AXIS_DIN_TDATA_delay[210]; // rv 0
  assign S_AXIS_DIN_TDATA_in[211] = (S_AXIS_DIN_TDATA[211] !== 1'bz) && S_AXIS_DIN_TDATA_delay[211]; // rv 0
  assign S_AXIS_DIN_TDATA_in[212] = (S_AXIS_DIN_TDATA[212] !== 1'bz) && S_AXIS_DIN_TDATA_delay[212]; // rv 0
  assign S_AXIS_DIN_TDATA_in[213] = (S_AXIS_DIN_TDATA[213] !== 1'bz) && S_AXIS_DIN_TDATA_delay[213]; // rv 0
  assign S_AXIS_DIN_TDATA_in[214] = (S_AXIS_DIN_TDATA[214] !== 1'bz) && S_AXIS_DIN_TDATA_delay[214]; // rv 0
  assign S_AXIS_DIN_TDATA_in[215] = (S_AXIS_DIN_TDATA[215] !== 1'bz) && S_AXIS_DIN_TDATA_delay[215]; // rv 0
  assign S_AXIS_DIN_TDATA_in[216] = (S_AXIS_DIN_TDATA[216] !== 1'bz) && S_AXIS_DIN_TDATA_delay[216]; // rv 0
  assign S_AXIS_DIN_TDATA_in[217] = (S_AXIS_DIN_TDATA[217] !== 1'bz) && S_AXIS_DIN_TDATA_delay[217]; // rv 0
  assign S_AXIS_DIN_TDATA_in[218] = (S_AXIS_DIN_TDATA[218] !== 1'bz) && S_AXIS_DIN_TDATA_delay[218]; // rv 0
  assign S_AXIS_DIN_TDATA_in[219] = (S_AXIS_DIN_TDATA[219] !== 1'bz) && S_AXIS_DIN_TDATA_delay[219]; // rv 0
  assign S_AXIS_DIN_TDATA_in[21] = (S_AXIS_DIN_TDATA[21] !== 1'bz) && S_AXIS_DIN_TDATA_delay[21]; // rv 0
  assign S_AXIS_DIN_TDATA_in[220] = (S_AXIS_DIN_TDATA[220] !== 1'bz) && S_AXIS_DIN_TDATA_delay[220]; // rv 0
  assign S_AXIS_DIN_TDATA_in[221] = (S_AXIS_DIN_TDATA[221] !== 1'bz) && S_AXIS_DIN_TDATA_delay[221]; // rv 0
  assign S_AXIS_DIN_TDATA_in[222] = (S_AXIS_DIN_TDATA[222] !== 1'bz) && S_AXIS_DIN_TDATA_delay[222]; // rv 0
  assign S_AXIS_DIN_TDATA_in[223] = (S_AXIS_DIN_TDATA[223] !== 1'bz) && S_AXIS_DIN_TDATA_delay[223]; // rv 0
  assign S_AXIS_DIN_TDATA_in[224] = (S_AXIS_DIN_TDATA[224] !== 1'bz) && S_AXIS_DIN_TDATA_delay[224]; // rv 0
  assign S_AXIS_DIN_TDATA_in[225] = (S_AXIS_DIN_TDATA[225] !== 1'bz) && S_AXIS_DIN_TDATA_delay[225]; // rv 0
  assign S_AXIS_DIN_TDATA_in[226] = (S_AXIS_DIN_TDATA[226] !== 1'bz) && S_AXIS_DIN_TDATA_delay[226]; // rv 0
  assign S_AXIS_DIN_TDATA_in[227] = (S_AXIS_DIN_TDATA[227] !== 1'bz) && S_AXIS_DIN_TDATA_delay[227]; // rv 0
  assign S_AXIS_DIN_TDATA_in[228] = (S_AXIS_DIN_TDATA[228] !== 1'bz) && S_AXIS_DIN_TDATA_delay[228]; // rv 0
  assign S_AXIS_DIN_TDATA_in[229] = (S_AXIS_DIN_TDATA[229] !== 1'bz) && S_AXIS_DIN_TDATA_delay[229]; // rv 0
  assign S_AXIS_DIN_TDATA_in[22] = (S_AXIS_DIN_TDATA[22] !== 1'bz) && S_AXIS_DIN_TDATA_delay[22]; // rv 0
  assign S_AXIS_DIN_TDATA_in[230] = (S_AXIS_DIN_TDATA[230] !== 1'bz) && S_AXIS_DIN_TDATA_delay[230]; // rv 0
  assign S_AXIS_DIN_TDATA_in[231] = (S_AXIS_DIN_TDATA[231] !== 1'bz) && S_AXIS_DIN_TDATA_delay[231]; // rv 0
  assign S_AXIS_DIN_TDATA_in[232] = (S_AXIS_DIN_TDATA[232] !== 1'bz) && S_AXIS_DIN_TDATA_delay[232]; // rv 0
  assign S_AXIS_DIN_TDATA_in[233] = (S_AXIS_DIN_TDATA[233] !== 1'bz) && S_AXIS_DIN_TDATA_delay[233]; // rv 0
  assign S_AXIS_DIN_TDATA_in[234] = (S_AXIS_DIN_TDATA[234] !== 1'bz) && S_AXIS_DIN_TDATA_delay[234]; // rv 0
  assign S_AXIS_DIN_TDATA_in[235] = (S_AXIS_DIN_TDATA[235] !== 1'bz) && S_AXIS_DIN_TDATA_delay[235]; // rv 0
  assign S_AXIS_DIN_TDATA_in[236] = (S_AXIS_DIN_TDATA[236] !== 1'bz) && S_AXIS_DIN_TDATA_delay[236]; // rv 0
  assign S_AXIS_DIN_TDATA_in[237] = (S_AXIS_DIN_TDATA[237] !== 1'bz) && S_AXIS_DIN_TDATA_delay[237]; // rv 0
  assign S_AXIS_DIN_TDATA_in[238] = (S_AXIS_DIN_TDATA[238] !== 1'bz) && S_AXIS_DIN_TDATA_delay[238]; // rv 0
  assign S_AXIS_DIN_TDATA_in[239] = (S_AXIS_DIN_TDATA[239] !== 1'bz) && S_AXIS_DIN_TDATA_delay[239]; // rv 0
  assign S_AXIS_DIN_TDATA_in[23] = (S_AXIS_DIN_TDATA[23] !== 1'bz) && S_AXIS_DIN_TDATA_delay[23]; // rv 0
  assign S_AXIS_DIN_TDATA_in[240] = (S_AXIS_DIN_TDATA[240] !== 1'bz) && S_AXIS_DIN_TDATA_delay[240]; // rv 0
  assign S_AXIS_DIN_TDATA_in[241] = (S_AXIS_DIN_TDATA[241] !== 1'bz) && S_AXIS_DIN_TDATA_delay[241]; // rv 0
  assign S_AXIS_DIN_TDATA_in[242] = (S_AXIS_DIN_TDATA[242] !== 1'bz) && S_AXIS_DIN_TDATA_delay[242]; // rv 0
  assign S_AXIS_DIN_TDATA_in[243] = (S_AXIS_DIN_TDATA[243] !== 1'bz) && S_AXIS_DIN_TDATA_delay[243]; // rv 0
  assign S_AXIS_DIN_TDATA_in[244] = (S_AXIS_DIN_TDATA[244] !== 1'bz) && S_AXIS_DIN_TDATA_delay[244]; // rv 0
  assign S_AXIS_DIN_TDATA_in[245] = (S_AXIS_DIN_TDATA[245] !== 1'bz) && S_AXIS_DIN_TDATA_delay[245]; // rv 0
  assign S_AXIS_DIN_TDATA_in[246] = (S_AXIS_DIN_TDATA[246] !== 1'bz) && S_AXIS_DIN_TDATA_delay[246]; // rv 0
  assign S_AXIS_DIN_TDATA_in[247] = (S_AXIS_DIN_TDATA[247] !== 1'bz) && S_AXIS_DIN_TDATA_delay[247]; // rv 0
  assign S_AXIS_DIN_TDATA_in[248] = (S_AXIS_DIN_TDATA[248] !== 1'bz) && S_AXIS_DIN_TDATA_delay[248]; // rv 0
  assign S_AXIS_DIN_TDATA_in[249] = (S_AXIS_DIN_TDATA[249] !== 1'bz) && S_AXIS_DIN_TDATA_delay[249]; // rv 0
  assign S_AXIS_DIN_TDATA_in[24] = (S_AXIS_DIN_TDATA[24] !== 1'bz) && S_AXIS_DIN_TDATA_delay[24]; // rv 0
  assign S_AXIS_DIN_TDATA_in[250] = (S_AXIS_DIN_TDATA[250] !== 1'bz) && S_AXIS_DIN_TDATA_delay[250]; // rv 0
  assign S_AXIS_DIN_TDATA_in[251] = (S_AXIS_DIN_TDATA[251] !== 1'bz) && S_AXIS_DIN_TDATA_delay[251]; // rv 0
  assign S_AXIS_DIN_TDATA_in[252] = (S_AXIS_DIN_TDATA[252] !== 1'bz) && S_AXIS_DIN_TDATA_delay[252]; // rv 0
  assign S_AXIS_DIN_TDATA_in[253] = (S_AXIS_DIN_TDATA[253] !== 1'bz) && S_AXIS_DIN_TDATA_delay[253]; // rv 0
  assign S_AXIS_DIN_TDATA_in[254] = (S_AXIS_DIN_TDATA[254] !== 1'bz) && S_AXIS_DIN_TDATA_delay[254]; // rv 0
  assign S_AXIS_DIN_TDATA_in[255] = (S_AXIS_DIN_TDATA[255] !== 1'bz) && S_AXIS_DIN_TDATA_delay[255]; // rv 0
  assign S_AXIS_DIN_TDATA_in[256] = (S_AXIS_DIN_TDATA[256] !== 1'bz) && S_AXIS_DIN_TDATA_delay[256]; // rv 0
  assign S_AXIS_DIN_TDATA_in[257] = (S_AXIS_DIN_TDATA[257] !== 1'bz) && S_AXIS_DIN_TDATA_delay[257]; // rv 0
  assign S_AXIS_DIN_TDATA_in[258] = (S_AXIS_DIN_TDATA[258] !== 1'bz) && S_AXIS_DIN_TDATA_delay[258]; // rv 0
  assign S_AXIS_DIN_TDATA_in[259] = (S_AXIS_DIN_TDATA[259] !== 1'bz) && S_AXIS_DIN_TDATA_delay[259]; // rv 0
  assign S_AXIS_DIN_TDATA_in[25] = (S_AXIS_DIN_TDATA[25] !== 1'bz) && S_AXIS_DIN_TDATA_delay[25]; // rv 0
  assign S_AXIS_DIN_TDATA_in[260] = (S_AXIS_DIN_TDATA[260] !== 1'bz) && S_AXIS_DIN_TDATA_delay[260]; // rv 0
  assign S_AXIS_DIN_TDATA_in[261] = (S_AXIS_DIN_TDATA[261] !== 1'bz) && S_AXIS_DIN_TDATA_delay[261]; // rv 0
  assign S_AXIS_DIN_TDATA_in[262] = (S_AXIS_DIN_TDATA[262] !== 1'bz) && S_AXIS_DIN_TDATA_delay[262]; // rv 0
  assign S_AXIS_DIN_TDATA_in[263] = (S_AXIS_DIN_TDATA[263] !== 1'bz) && S_AXIS_DIN_TDATA_delay[263]; // rv 0
  assign S_AXIS_DIN_TDATA_in[264] = (S_AXIS_DIN_TDATA[264] !== 1'bz) && S_AXIS_DIN_TDATA_delay[264]; // rv 0
  assign S_AXIS_DIN_TDATA_in[265] = (S_AXIS_DIN_TDATA[265] !== 1'bz) && S_AXIS_DIN_TDATA_delay[265]; // rv 0
  assign S_AXIS_DIN_TDATA_in[266] = (S_AXIS_DIN_TDATA[266] !== 1'bz) && S_AXIS_DIN_TDATA_delay[266]; // rv 0
  assign S_AXIS_DIN_TDATA_in[267] = (S_AXIS_DIN_TDATA[267] !== 1'bz) && S_AXIS_DIN_TDATA_delay[267]; // rv 0
  assign S_AXIS_DIN_TDATA_in[268] = (S_AXIS_DIN_TDATA[268] !== 1'bz) && S_AXIS_DIN_TDATA_delay[268]; // rv 0
  assign S_AXIS_DIN_TDATA_in[269] = (S_AXIS_DIN_TDATA[269] !== 1'bz) && S_AXIS_DIN_TDATA_delay[269]; // rv 0
  assign S_AXIS_DIN_TDATA_in[26] = (S_AXIS_DIN_TDATA[26] !== 1'bz) && S_AXIS_DIN_TDATA_delay[26]; // rv 0
  assign S_AXIS_DIN_TDATA_in[270] = (S_AXIS_DIN_TDATA[270] !== 1'bz) && S_AXIS_DIN_TDATA_delay[270]; // rv 0
  assign S_AXIS_DIN_TDATA_in[271] = (S_AXIS_DIN_TDATA[271] !== 1'bz) && S_AXIS_DIN_TDATA_delay[271]; // rv 0
  assign S_AXIS_DIN_TDATA_in[272] = (S_AXIS_DIN_TDATA[272] !== 1'bz) && S_AXIS_DIN_TDATA_delay[272]; // rv 0
  assign S_AXIS_DIN_TDATA_in[273] = (S_AXIS_DIN_TDATA[273] !== 1'bz) && S_AXIS_DIN_TDATA_delay[273]; // rv 0
  assign S_AXIS_DIN_TDATA_in[274] = (S_AXIS_DIN_TDATA[274] !== 1'bz) && S_AXIS_DIN_TDATA_delay[274]; // rv 0
  assign S_AXIS_DIN_TDATA_in[275] = (S_AXIS_DIN_TDATA[275] !== 1'bz) && S_AXIS_DIN_TDATA_delay[275]; // rv 0
  assign S_AXIS_DIN_TDATA_in[276] = (S_AXIS_DIN_TDATA[276] !== 1'bz) && S_AXIS_DIN_TDATA_delay[276]; // rv 0
  assign S_AXIS_DIN_TDATA_in[277] = (S_AXIS_DIN_TDATA[277] !== 1'bz) && S_AXIS_DIN_TDATA_delay[277]; // rv 0
  assign S_AXIS_DIN_TDATA_in[278] = (S_AXIS_DIN_TDATA[278] !== 1'bz) && S_AXIS_DIN_TDATA_delay[278]; // rv 0
  assign S_AXIS_DIN_TDATA_in[279] = (S_AXIS_DIN_TDATA[279] !== 1'bz) && S_AXIS_DIN_TDATA_delay[279]; // rv 0
  assign S_AXIS_DIN_TDATA_in[27] = (S_AXIS_DIN_TDATA[27] !== 1'bz) && S_AXIS_DIN_TDATA_delay[27]; // rv 0
  assign S_AXIS_DIN_TDATA_in[280] = (S_AXIS_DIN_TDATA[280] !== 1'bz) && S_AXIS_DIN_TDATA_delay[280]; // rv 0
  assign S_AXIS_DIN_TDATA_in[281] = (S_AXIS_DIN_TDATA[281] !== 1'bz) && S_AXIS_DIN_TDATA_delay[281]; // rv 0
  assign S_AXIS_DIN_TDATA_in[282] = (S_AXIS_DIN_TDATA[282] !== 1'bz) && S_AXIS_DIN_TDATA_delay[282]; // rv 0
  assign S_AXIS_DIN_TDATA_in[283] = (S_AXIS_DIN_TDATA[283] !== 1'bz) && S_AXIS_DIN_TDATA_delay[283]; // rv 0
  assign S_AXIS_DIN_TDATA_in[284] = (S_AXIS_DIN_TDATA[284] !== 1'bz) && S_AXIS_DIN_TDATA_delay[284]; // rv 0
  assign S_AXIS_DIN_TDATA_in[285] = (S_AXIS_DIN_TDATA[285] !== 1'bz) && S_AXIS_DIN_TDATA_delay[285]; // rv 0
  assign S_AXIS_DIN_TDATA_in[286] = (S_AXIS_DIN_TDATA[286] !== 1'bz) && S_AXIS_DIN_TDATA_delay[286]; // rv 0
  assign S_AXIS_DIN_TDATA_in[287] = (S_AXIS_DIN_TDATA[287] !== 1'bz) && S_AXIS_DIN_TDATA_delay[287]; // rv 0
  assign S_AXIS_DIN_TDATA_in[288] = (S_AXIS_DIN_TDATA[288] !== 1'bz) && S_AXIS_DIN_TDATA_delay[288]; // rv 0
  assign S_AXIS_DIN_TDATA_in[289] = (S_AXIS_DIN_TDATA[289] !== 1'bz) && S_AXIS_DIN_TDATA_delay[289]; // rv 0
  assign S_AXIS_DIN_TDATA_in[28] = (S_AXIS_DIN_TDATA[28] !== 1'bz) && S_AXIS_DIN_TDATA_delay[28]; // rv 0
  assign S_AXIS_DIN_TDATA_in[290] = (S_AXIS_DIN_TDATA[290] !== 1'bz) && S_AXIS_DIN_TDATA_delay[290]; // rv 0
  assign S_AXIS_DIN_TDATA_in[291] = (S_AXIS_DIN_TDATA[291] !== 1'bz) && S_AXIS_DIN_TDATA_delay[291]; // rv 0
  assign S_AXIS_DIN_TDATA_in[292] = (S_AXIS_DIN_TDATA[292] !== 1'bz) && S_AXIS_DIN_TDATA_delay[292]; // rv 0
  assign S_AXIS_DIN_TDATA_in[293] = (S_AXIS_DIN_TDATA[293] !== 1'bz) && S_AXIS_DIN_TDATA_delay[293]; // rv 0
  assign S_AXIS_DIN_TDATA_in[294] = (S_AXIS_DIN_TDATA[294] !== 1'bz) && S_AXIS_DIN_TDATA_delay[294]; // rv 0
  assign S_AXIS_DIN_TDATA_in[295] = (S_AXIS_DIN_TDATA[295] !== 1'bz) && S_AXIS_DIN_TDATA_delay[295]; // rv 0
  assign S_AXIS_DIN_TDATA_in[296] = (S_AXIS_DIN_TDATA[296] !== 1'bz) && S_AXIS_DIN_TDATA_delay[296]; // rv 0
  assign S_AXIS_DIN_TDATA_in[297] = (S_AXIS_DIN_TDATA[297] !== 1'bz) && S_AXIS_DIN_TDATA_delay[297]; // rv 0
  assign S_AXIS_DIN_TDATA_in[298] = (S_AXIS_DIN_TDATA[298] !== 1'bz) && S_AXIS_DIN_TDATA_delay[298]; // rv 0
  assign S_AXIS_DIN_TDATA_in[299] = (S_AXIS_DIN_TDATA[299] !== 1'bz) && S_AXIS_DIN_TDATA_delay[299]; // rv 0
  assign S_AXIS_DIN_TDATA_in[29] = (S_AXIS_DIN_TDATA[29] !== 1'bz) && S_AXIS_DIN_TDATA_delay[29]; // rv 0
  assign S_AXIS_DIN_TDATA_in[2] = (S_AXIS_DIN_TDATA[2] !== 1'bz) && S_AXIS_DIN_TDATA_delay[2]; // rv 0
  assign S_AXIS_DIN_TDATA_in[300] = (S_AXIS_DIN_TDATA[300] !== 1'bz) && S_AXIS_DIN_TDATA_delay[300]; // rv 0
  assign S_AXIS_DIN_TDATA_in[301] = (S_AXIS_DIN_TDATA[301] !== 1'bz) && S_AXIS_DIN_TDATA_delay[301]; // rv 0
  assign S_AXIS_DIN_TDATA_in[302] = (S_AXIS_DIN_TDATA[302] !== 1'bz) && S_AXIS_DIN_TDATA_delay[302]; // rv 0
  assign S_AXIS_DIN_TDATA_in[303] = (S_AXIS_DIN_TDATA[303] !== 1'bz) && S_AXIS_DIN_TDATA_delay[303]; // rv 0
  assign S_AXIS_DIN_TDATA_in[304] = (S_AXIS_DIN_TDATA[304] !== 1'bz) && S_AXIS_DIN_TDATA_delay[304]; // rv 0
  assign S_AXIS_DIN_TDATA_in[305] = (S_AXIS_DIN_TDATA[305] !== 1'bz) && S_AXIS_DIN_TDATA_delay[305]; // rv 0
  assign S_AXIS_DIN_TDATA_in[306] = (S_AXIS_DIN_TDATA[306] !== 1'bz) && S_AXIS_DIN_TDATA_delay[306]; // rv 0
  assign S_AXIS_DIN_TDATA_in[307] = (S_AXIS_DIN_TDATA[307] !== 1'bz) && S_AXIS_DIN_TDATA_delay[307]; // rv 0
  assign S_AXIS_DIN_TDATA_in[308] = (S_AXIS_DIN_TDATA[308] !== 1'bz) && S_AXIS_DIN_TDATA_delay[308]; // rv 0
  assign S_AXIS_DIN_TDATA_in[309] = (S_AXIS_DIN_TDATA[309] !== 1'bz) && S_AXIS_DIN_TDATA_delay[309]; // rv 0
  assign S_AXIS_DIN_TDATA_in[30] = (S_AXIS_DIN_TDATA[30] !== 1'bz) && S_AXIS_DIN_TDATA_delay[30]; // rv 0
  assign S_AXIS_DIN_TDATA_in[310] = (S_AXIS_DIN_TDATA[310] !== 1'bz) && S_AXIS_DIN_TDATA_delay[310]; // rv 0
  assign S_AXIS_DIN_TDATA_in[311] = (S_AXIS_DIN_TDATA[311] !== 1'bz) && S_AXIS_DIN_TDATA_delay[311]; // rv 0
  assign S_AXIS_DIN_TDATA_in[312] = (S_AXIS_DIN_TDATA[312] !== 1'bz) && S_AXIS_DIN_TDATA_delay[312]; // rv 0
  assign S_AXIS_DIN_TDATA_in[313] = (S_AXIS_DIN_TDATA[313] !== 1'bz) && S_AXIS_DIN_TDATA_delay[313]; // rv 0
  assign S_AXIS_DIN_TDATA_in[314] = (S_AXIS_DIN_TDATA[314] !== 1'bz) && S_AXIS_DIN_TDATA_delay[314]; // rv 0
  assign S_AXIS_DIN_TDATA_in[315] = (S_AXIS_DIN_TDATA[315] !== 1'bz) && S_AXIS_DIN_TDATA_delay[315]; // rv 0
  assign S_AXIS_DIN_TDATA_in[316] = (S_AXIS_DIN_TDATA[316] !== 1'bz) && S_AXIS_DIN_TDATA_delay[316]; // rv 0
  assign S_AXIS_DIN_TDATA_in[317] = (S_AXIS_DIN_TDATA[317] !== 1'bz) && S_AXIS_DIN_TDATA_delay[317]; // rv 0
  assign S_AXIS_DIN_TDATA_in[318] = (S_AXIS_DIN_TDATA[318] !== 1'bz) && S_AXIS_DIN_TDATA_delay[318]; // rv 0
  assign S_AXIS_DIN_TDATA_in[319] = (S_AXIS_DIN_TDATA[319] !== 1'bz) && S_AXIS_DIN_TDATA_delay[319]; // rv 0
  assign S_AXIS_DIN_TDATA_in[31] = (S_AXIS_DIN_TDATA[31] !== 1'bz) && S_AXIS_DIN_TDATA_delay[31]; // rv 0
  assign S_AXIS_DIN_TDATA_in[320] = (S_AXIS_DIN_TDATA[320] !== 1'bz) && S_AXIS_DIN_TDATA_delay[320]; // rv 0
  assign S_AXIS_DIN_TDATA_in[321] = (S_AXIS_DIN_TDATA[321] !== 1'bz) && S_AXIS_DIN_TDATA_delay[321]; // rv 0
  assign S_AXIS_DIN_TDATA_in[322] = (S_AXIS_DIN_TDATA[322] !== 1'bz) && S_AXIS_DIN_TDATA_delay[322]; // rv 0
  assign S_AXIS_DIN_TDATA_in[323] = (S_AXIS_DIN_TDATA[323] !== 1'bz) && S_AXIS_DIN_TDATA_delay[323]; // rv 0
  assign S_AXIS_DIN_TDATA_in[324] = (S_AXIS_DIN_TDATA[324] !== 1'bz) && S_AXIS_DIN_TDATA_delay[324]; // rv 0
  assign S_AXIS_DIN_TDATA_in[325] = (S_AXIS_DIN_TDATA[325] !== 1'bz) && S_AXIS_DIN_TDATA_delay[325]; // rv 0
  assign S_AXIS_DIN_TDATA_in[326] = (S_AXIS_DIN_TDATA[326] !== 1'bz) && S_AXIS_DIN_TDATA_delay[326]; // rv 0
  assign S_AXIS_DIN_TDATA_in[327] = (S_AXIS_DIN_TDATA[327] !== 1'bz) && S_AXIS_DIN_TDATA_delay[327]; // rv 0
  assign S_AXIS_DIN_TDATA_in[328] = (S_AXIS_DIN_TDATA[328] !== 1'bz) && S_AXIS_DIN_TDATA_delay[328]; // rv 0
  assign S_AXIS_DIN_TDATA_in[329] = (S_AXIS_DIN_TDATA[329] !== 1'bz) && S_AXIS_DIN_TDATA_delay[329]; // rv 0
  assign S_AXIS_DIN_TDATA_in[32] = (S_AXIS_DIN_TDATA[32] !== 1'bz) && S_AXIS_DIN_TDATA_delay[32]; // rv 0
  assign S_AXIS_DIN_TDATA_in[330] = (S_AXIS_DIN_TDATA[330] !== 1'bz) && S_AXIS_DIN_TDATA_delay[330]; // rv 0
  assign S_AXIS_DIN_TDATA_in[331] = (S_AXIS_DIN_TDATA[331] !== 1'bz) && S_AXIS_DIN_TDATA_delay[331]; // rv 0
  assign S_AXIS_DIN_TDATA_in[332] = (S_AXIS_DIN_TDATA[332] !== 1'bz) && S_AXIS_DIN_TDATA_delay[332]; // rv 0
  assign S_AXIS_DIN_TDATA_in[333] = (S_AXIS_DIN_TDATA[333] !== 1'bz) && S_AXIS_DIN_TDATA_delay[333]; // rv 0
  assign S_AXIS_DIN_TDATA_in[334] = (S_AXIS_DIN_TDATA[334] !== 1'bz) && S_AXIS_DIN_TDATA_delay[334]; // rv 0
  assign S_AXIS_DIN_TDATA_in[335] = (S_AXIS_DIN_TDATA[335] !== 1'bz) && S_AXIS_DIN_TDATA_delay[335]; // rv 0
  assign S_AXIS_DIN_TDATA_in[336] = (S_AXIS_DIN_TDATA[336] !== 1'bz) && S_AXIS_DIN_TDATA_delay[336]; // rv 0
  assign S_AXIS_DIN_TDATA_in[337] = (S_AXIS_DIN_TDATA[337] !== 1'bz) && S_AXIS_DIN_TDATA_delay[337]; // rv 0
  assign S_AXIS_DIN_TDATA_in[338] = (S_AXIS_DIN_TDATA[338] !== 1'bz) && S_AXIS_DIN_TDATA_delay[338]; // rv 0
  assign S_AXIS_DIN_TDATA_in[339] = (S_AXIS_DIN_TDATA[339] !== 1'bz) && S_AXIS_DIN_TDATA_delay[339]; // rv 0
  assign S_AXIS_DIN_TDATA_in[33] = (S_AXIS_DIN_TDATA[33] !== 1'bz) && S_AXIS_DIN_TDATA_delay[33]; // rv 0
  assign S_AXIS_DIN_TDATA_in[340] = (S_AXIS_DIN_TDATA[340] !== 1'bz) && S_AXIS_DIN_TDATA_delay[340]; // rv 0
  assign S_AXIS_DIN_TDATA_in[341] = (S_AXIS_DIN_TDATA[341] !== 1'bz) && S_AXIS_DIN_TDATA_delay[341]; // rv 0
  assign S_AXIS_DIN_TDATA_in[342] = (S_AXIS_DIN_TDATA[342] !== 1'bz) && S_AXIS_DIN_TDATA_delay[342]; // rv 0
  assign S_AXIS_DIN_TDATA_in[343] = (S_AXIS_DIN_TDATA[343] !== 1'bz) && S_AXIS_DIN_TDATA_delay[343]; // rv 0
  assign S_AXIS_DIN_TDATA_in[344] = (S_AXIS_DIN_TDATA[344] !== 1'bz) && S_AXIS_DIN_TDATA_delay[344]; // rv 0
  assign S_AXIS_DIN_TDATA_in[345] = (S_AXIS_DIN_TDATA[345] !== 1'bz) && S_AXIS_DIN_TDATA_delay[345]; // rv 0
  assign S_AXIS_DIN_TDATA_in[346] = (S_AXIS_DIN_TDATA[346] !== 1'bz) && S_AXIS_DIN_TDATA_delay[346]; // rv 0
  assign S_AXIS_DIN_TDATA_in[347] = (S_AXIS_DIN_TDATA[347] !== 1'bz) && S_AXIS_DIN_TDATA_delay[347]; // rv 0
  assign S_AXIS_DIN_TDATA_in[348] = (S_AXIS_DIN_TDATA[348] !== 1'bz) && S_AXIS_DIN_TDATA_delay[348]; // rv 0
  assign S_AXIS_DIN_TDATA_in[349] = (S_AXIS_DIN_TDATA[349] !== 1'bz) && S_AXIS_DIN_TDATA_delay[349]; // rv 0
  assign S_AXIS_DIN_TDATA_in[34] = (S_AXIS_DIN_TDATA[34] !== 1'bz) && S_AXIS_DIN_TDATA_delay[34]; // rv 0
  assign S_AXIS_DIN_TDATA_in[350] = (S_AXIS_DIN_TDATA[350] !== 1'bz) && S_AXIS_DIN_TDATA_delay[350]; // rv 0
  assign S_AXIS_DIN_TDATA_in[351] = (S_AXIS_DIN_TDATA[351] !== 1'bz) && S_AXIS_DIN_TDATA_delay[351]; // rv 0
  assign S_AXIS_DIN_TDATA_in[352] = (S_AXIS_DIN_TDATA[352] !== 1'bz) && S_AXIS_DIN_TDATA_delay[352]; // rv 0
  assign S_AXIS_DIN_TDATA_in[353] = (S_AXIS_DIN_TDATA[353] !== 1'bz) && S_AXIS_DIN_TDATA_delay[353]; // rv 0
  assign S_AXIS_DIN_TDATA_in[354] = (S_AXIS_DIN_TDATA[354] !== 1'bz) && S_AXIS_DIN_TDATA_delay[354]; // rv 0
  assign S_AXIS_DIN_TDATA_in[355] = (S_AXIS_DIN_TDATA[355] !== 1'bz) && S_AXIS_DIN_TDATA_delay[355]; // rv 0
  assign S_AXIS_DIN_TDATA_in[356] = (S_AXIS_DIN_TDATA[356] !== 1'bz) && S_AXIS_DIN_TDATA_delay[356]; // rv 0
  assign S_AXIS_DIN_TDATA_in[357] = (S_AXIS_DIN_TDATA[357] !== 1'bz) && S_AXIS_DIN_TDATA_delay[357]; // rv 0
  assign S_AXIS_DIN_TDATA_in[358] = (S_AXIS_DIN_TDATA[358] !== 1'bz) && S_AXIS_DIN_TDATA_delay[358]; // rv 0
  assign S_AXIS_DIN_TDATA_in[359] = (S_AXIS_DIN_TDATA[359] !== 1'bz) && S_AXIS_DIN_TDATA_delay[359]; // rv 0
  assign S_AXIS_DIN_TDATA_in[35] = (S_AXIS_DIN_TDATA[35] !== 1'bz) && S_AXIS_DIN_TDATA_delay[35]; // rv 0
  assign S_AXIS_DIN_TDATA_in[360] = (S_AXIS_DIN_TDATA[360] !== 1'bz) && S_AXIS_DIN_TDATA_delay[360]; // rv 0
  assign S_AXIS_DIN_TDATA_in[361] = (S_AXIS_DIN_TDATA[361] !== 1'bz) && S_AXIS_DIN_TDATA_delay[361]; // rv 0
  assign S_AXIS_DIN_TDATA_in[362] = (S_AXIS_DIN_TDATA[362] !== 1'bz) && S_AXIS_DIN_TDATA_delay[362]; // rv 0
  assign S_AXIS_DIN_TDATA_in[363] = (S_AXIS_DIN_TDATA[363] !== 1'bz) && S_AXIS_DIN_TDATA_delay[363]; // rv 0
  assign S_AXIS_DIN_TDATA_in[364] = (S_AXIS_DIN_TDATA[364] !== 1'bz) && S_AXIS_DIN_TDATA_delay[364]; // rv 0
  assign S_AXIS_DIN_TDATA_in[365] = (S_AXIS_DIN_TDATA[365] !== 1'bz) && S_AXIS_DIN_TDATA_delay[365]; // rv 0
  assign S_AXIS_DIN_TDATA_in[366] = (S_AXIS_DIN_TDATA[366] !== 1'bz) && S_AXIS_DIN_TDATA_delay[366]; // rv 0
  assign S_AXIS_DIN_TDATA_in[367] = (S_AXIS_DIN_TDATA[367] !== 1'bz) && S_AXIS_DIN_TDATA_delay[367]; // rv 0
  assign S_AXIS_DIN_TDATA_in[368] = (S_AXIS_DIN_TDATA[368] !== 1'bz) && S_AXIS_DIN_TDATA_delay[368]; // rv 0
  assign S_AXIS_DIN_TDATA_in[369] = (S_AXIS_DIN_TDATA[369] !== 1'bz) && S_AXIS_DIN_TDATA_delay[369]; // rv 0
  assign S_AXIS_DIN_TDATA_in[36] = (S_AXIS_DIN_TDATA[36] !== 1'bz) && S_AXIS_DIN_TDATA_delay[36]; // rv 0
  assign S_AXIS_DIN_TDATA_in[370] = (S_AXIS_DIN_TDATA[370] !== 1'bz) && S_AXIS_DIN_TDATA_delay[370]; // rv 0
  assign S_AXIS_DIN_TDATA_in[371] = (S_AXIS_DIN_TDATA[371] !== 1'bz) && S_AXIS_DIN_TDATA_delay[371]; // rv 0
  assign S_AXIS_DIN_TDATA_in[372] = (S_AXIS_DIN_TDATA[372] !== 1'bz) && S_AXIS_DIN_TDATA_delay[372]; // rv 0
  assign S_AXIS_DIN_TDATA_in[373] = (S_AXIS_DIN_TDATA[373] !== 1'bz) && S_AXIS_DIN_TDATA_delay[373]; // rv 0
  assign S_AXIS_DIN_TDATA_in[374] = (S_AXIS_DIN_TDATA[374] !== 1'bz) && S_AXIS_DIN_TDATA_delay[374]; // rv 0
  assign S_AXIS_DIN_TDATA_in[375] = (S_AXIS_DIN_TDATA[375] !== 1'bz) && S_AXIS_DIN_TDATA_delay[375]; // rv 0
  assign S_AXIS_DIN_TDATA_in[376] = (S_AXIS_DIN_TDATA[376] !== 1'bz) && S_AXIS_DIN_TDATA_delay[376]; // rv 0
  assign S_AXIS_DIN_TDATA_in[377] = (S_AXIS_DIN_TDATA[377] !== 1'bz) && S_AXIS_DIN_TDATA_delay[377]; // rv 0
  assign S_AXIS_DIN_TDATA_in[378] = (S_AXIS_DIN_TDATA[378] !== 1'bz) && S_AXIS_DIN_TDATA_delay[378]; // rv 0
  assign S_AXIS_DIN_TDATA_in[379] = (S_AXIS_DIN_TDATA[379] !== 1'bz) && S_AXIS_DIN_TDATA_delay[379]; // rv 0
  assign S_AXIS_DIN_TDATA_in[37] = (S_AXIS_DIN_TDATA[37] !== 1'bz) && S_AXIS_DIN_TDATA_delay[37]; // rv 0
  assign S_AXIS_DIN_TDATA_in[380] = (S_AXIS_DIN_TDATA[380] !== 1'bz) && S_AXIS_DIN_TDATA_delay[380]; // rv 0
  assign S_AXIS_DIN_TDATA_in[381] = (S_AXIS_DIN_TDATA[381] !== 1'bz) && S_AXIS_DIN_TDATA_delay[381]; // rv 0
  assign S_AXIS_DIN_TDATA_in[382] = (S_AXIS_DIN_TDATA[382] !== 1'bz) && S_AXIS_DIN_TDATA_delay[382]; // rv 0
  assign S_AXIS_DIN_TDATA_in[383] = (S_AXIS_DIN_TDATA[383] !== 1'bz) && S_AXIS_DIN_TDATA_delay[383]; // rv 0
  assign S_AXIS_DIN_TDATA_in[384] = (S_AXIS_DIN_TDATA[384] !== 1'bz) && S_AXIS_DIN_TDATA_delay[384]; // rv 0
  assign S_AXIS_DIN_TDATA_in[385] = (S_AXIS_DIN_TDATA[385] !== 1'bz) && S_AXIS_DIN_TDATA_delay[385]; // rv 0
  assign S_AXIS_DIN_TDATA_in[386] = (S_AXIS_DIN_TDATA[386] !== 1'bz) && S_AXIS_DIN_TDATA_delay[386]; // rv 0
  assign S_AXIS_DIN_TDATA_in[387] = (S_AXIS_DIN_TDATA[387] !== 1'bz) && S_AXIS_DIN_TDATA_delay[387]; // rv 0
  assign S_AXIS_DIN_TDATA_in[388] = (S_AXIS_DIN_TDATA[388] !== 1'bz) && S_AXIS_DIN_TDATA_delay[388]; // rv 0
  assign S_AXIS_DIN_TDATA_in[389] = (S_AXIS_DIN_TDATA[389] !== 1'bz) && S_AXIS_DIN_TDATA_delay[389]; // rv 0
  assign S_AXIS_DIN_TDATA_in[38] = (S_AXIS_DIN_TDATA[38] !== 1'bz) && S_AXIS_DIN_TDATA_delay[38]; // rv 0
  assign S_AXIS_DIN_TDATA_in[390] = (S_AXIS_DIN_TDATA[390] !== 1'bz) && S_AXIS_DIN_TDATA_delay[390]; // rv 0
  assign S_AXIS_DIN_TDATA_in[391] = (S_AXIS_DIN_TDATA[391] !== 1'bz) && S_AXIS_DIN_TDATA_delay[391]; // rv 0
  assign S_AXIS_DIN_TDATA_in[392] = (S_AXIS_DIN_TDATA[392] !== 1'bz) && S_AXIS_DIN_TDATA_delay[392]; // rv 0
  assign S_AXIS_DIN_TDATA_in[393] = (S_AXIS_DIN_TDATA[393] !== 1'bz) && S_AXIS_DIN_TDATA_delay[393]; // rv 0
  assign S_AXIS_DIN_TDATA_in[394] = (S_AXIS_DIN_TDATA[394] !== 1'bz) && S_AXIS_DIN_TDATA_delay[394]; // rv 0
  assign S_AXIS_DIN_TDATA_in[395] = (S_AXIS_DIN_TDATA[395] !== 1'bz) && S_AXIS_DIN_TDATA_delay[395]; // rv 0
  assign S_AXIS_DIN_TDATA_in[396] = (S_AXIS_DIN_TDATA[396] !== 1'bz) && S_AXIS_DIN_TDATA_delay[396]; // rv 0
  assign S_AXIS_DIN_TDATA_in[397] = (S_AXIS_DIN_TDATA[397] !== 1'bz) && S_AXIS_DIN_TDATA_delay[397]; // rv 0
  assign S_AXIS_DIN_TDATA_in[398] = (S_AXIS_DIN_TDATA[398] !== 1'bz) && S_AXIS_DIN_TDATA_delay[398]; // rv 0
  assign S_AXIS_DIN_TDATA_in[399] = (S_AXIS_DIN_TDATA[399] !== 1'bz) && S_AXIS_DIN_TDATA_delay[399]; // rv 0
  assign S_AXIS_DIN_TDATA_in[39] = (S_AXIS_DIN_TDATA[39] !== 1'bz) && S_AXIS_DIN_TDATA_delay[39]; // rv 0
  assign S_AXIS_DIN_TDATA_in[3] = (S_AXIS_DIN_TDATA[3] !== 1'bz) && S_AXIS_DIN_TDATA_delay[3]; // rv 0
  assign S_AXIS_DIN_TDATA_in[400] = (S_AXIS_DIN_TDATA[400] !== 1'bz) && S_AXIS_DIN_TDATA_delay[400]; // rv 0
  assign S_AXIS_DIN_TDATA_in[401] = (S_AXIS_DIN_TDATA[401] !== 1'bz) && S_AXIS_DIN_TDATA_delay[401]; // rv 0
  assign S_AXIS_DIN_TDATA_in[402] = (S_AXIS_DIN_TDATA[402] !== 1'bz) && S_AXIS_DIN_TDATA_delay[402]; // rv 0
  assign S_AXIS_DIN_TDATA_in[403] = (S_AXIS_DIN_TDATA[403] !== 1'bz) && S_AXIS_DIN_TDATA_delay[403]; // rv 0
  assign S_AXIS_DIN_TDATA_in[404] = (S_AXIS_DIN_TDATA[404] !== 1'bz) && S_AXIS_DIN_TDATA_delay[404]; // rv 0
  assign S_AXIS_DIN_TDATA_in[405] = (S_AXIS_DIN_TDATA[405] !== 1'bz) && S_AXIS_DIN_TDATA_delay[405]; // rv 0
  assign S_AXIS_DIN_TDATA_in[406] = (S_AXIS_DIN_TDATA[406] !== 1'bz) && S_AXIS_DIN_TDATA_delay[406]; // rv 0
  assign S_AXIS_DIN_TDATA_in[407] = (S_AXIS_DIN_TDATA[407] !== 1'bz) && S_AXIS_DIN_TDATA_delay[407]; // rv 0
  assign S_AXIS_DIN_TDATA_in[408] = (S_AXIS_DIN_TDATA[408] !== 1'bz) && S_AXIS_DIN_TDATA_delay[408]; // rv 0
  assign S_AXIS_DIN_TDATA_in[409] = (S_AXIS_DIN_TDATA[409] !== 1'bz) && S_AXIS_DIN_TDATA_delay[409]; // rv 0
  assign S_AXIS_DIN_TDATA_in[40] = (S_AXIS_DIN_TDATA[40] !== 1'bz) && S_AXIS_DIN_TDATA_delay[40]; // rv 0
  assign S_AXIS_DIN_TDATA_in[410] = (S_AXIS_DIN_TDATA[410] !== 1'bz) && S_AXIS_DIN_TDATA_delay[410]; // rv 0
  assign S_AXIS_DIN_TDATA_in[411] = (S_AXIS_DIN_TDATA[411] !== 1'bz) && S_AXIS_DIN_TDATA_delay[411]; // rv 0
  assign S_AXIS_DIN_TDATA_in[412] = (S_AXIS_DIN_TDATA[412] !== 1'bz) && S_AXIS_DIN_TDATA_delay[412]; // rv 0
  assign S_AXIS_DIN_TDATA_in[413] = (S_AXIS_DIN_TDATA[413] !== 1'bz) && S_AXIS_DIN_TDATA_delay[413]; // rv 0
  assign S_AXIS_DIN_TDATA_in[414] = (S_AXIS_DIN_TDATA[414] !== 1'bz) && S_AXIS_DIN_TDATA_delay[414]; // rv 0
  assign S_AXIS_DIN_TDATA_in[415] = (S_AXIS_DIN_TDATA[415] !== 1'bz) && S_AXIS_DIN_TDATA_delay[415]; // rv 0
  assign S_AXIS_DIN_TDATA_in[416] = (S_AXIS_DIN_TDATA[416] !== 1'bz) && S_AXIS_DIN_TDATA_delay[416]; // rv 0
  assign S_AXIS_DIN_TDATA_in[417] = (S_AXIS_DIN_TDATA[417] !== 1'bz) && S_AXIS_DIN_TDATA_delay[417]; // rv 0
  assign S_AXIS_DIN_TDATA_in[418] = (S_AXIS_DIN_TDATA[418] !== 1'bz) && S_AXIS_DIN_TDATA_delay[418]; // rv 0
  assign S_AXIS_DIN_TDATA_in[419] = (S_AXIS_DIN_TDATA[419] !== 1'bz) && S_AXIS_DIN_TDATA_delay[419]; // rv 0
  assign S_AXIS_DIN_TDATA_in[41] = (S_AXIS_DIN_TDATA[41] !== 1'bz) && S_AXIS_DIN_TDATA_delay[41]; // rv 0
  assign S_AXIS_DIN_TDATA_in[420] = (S_AXIS_DIN_TDATA[420] !== 1'bz) && S_AXIS_DIN_TDATA_delay[420]; // rv 0
  assign S_AXIS_DIN_TDATA_in[421] = (S_AXIS_DIN_TDATA[421] !== 1'bz) && S_AXIS_DIN_TDATA_delay[421]; // rv 0
  assign S_AXIS_DIN_TDATA_in[422] = (S_AXIS_DIN_TDATA[422] !== 1'bz) && S_AXIS_DIN_TDATA_delay[422]; // rv 0
  assign S_AXIS_DIN_TDATA_in[423] = (S_AXIS_DIN_TDATA[423] !== 1'bz) && S_AXIS_DIN_TDATA_delay[423]; // rv 0
  assign S_AXIS_DIN_TDATA_in[424] = (S_AXIS_DIN_TDATA[424] !== 1'bz) && S_AXIS_DIN_TDATA_delay[424]; // rv 0
  assign S_AXIS_DIN_TDATA_in[425] = (S_AXIS_DIN_TDATA[425] !== 1'bz) && S_AXIS_DIN_TDATA_delay[425]; // rv 0
  assign S_AXIS_DIN_TDATA_in[426] = (S_AXIS_DIN_TDATA[426] !== 1'bz) && S_AXIS_DIN_TDATA_delay[426]; // rv 0
  assign S_AXIS_DIN_TDATA_in[427] = (S_AXIS_DIN_TDATA[427] !== 1'bz) && S_AXIS_DIN_TDATA_delay[427]; // rv 0
  assign S_AXIS_DIN_TDATA_in[428] = (S_AXIS_DIN_TDATA[428] !== 1'bz) && S_AXIS_DIN_TDATA_delay[428]; // rv 0
  assign S_AXIS_DIN_TDATA_in[429] = (S_AXIS_DIN_TDATA[429] !== 1'bz) && S_AXIS_DIN_TDATA_delay[429]; // rv 0
  assign S_AXIS_DIN_TDATA_in[42] = (S_AXIS_DIN_TDATA[42] !== 1'bz) && S_AXIS_DIN_TDATA_delay[42]; // rv 0
  assign S_AXIS_DIN_TDATA_in[430] = (S_AXIS_DIN_TDATA[430] !== 1'bz) && S_AXIS_DIN_TDATA_delay[430]; // rv 0
  assign S_AXIS_DIN_TDATA_in[431] = (S_AXIS_DIN_TDATA[431] !== 1'bz) && S_AXIS_DIN_TDATA_delay[431]; // rv 0
  assign S_AXIS_DIN_TDATA_in[432] = (S_AXIS_DIN_TDATA[432] !== 1'bz) && S_AXIS_DIN_TDATA_delay[432]; // rv 0
  assign S_AXIS_DIN_TDATA_in[433] = (S_AXIS_DIN_TDATA[433] !== 1'bz) && S_AXIS_DIN_TDATA_delay[433]; // rv 0
  assign S_AXIS_DIN_TDATA_in[434] = (S_AXIS_DIN_TDATA[434] !== 1'bz) && S_AXIS_DIN_TDATA_delay[434]; // rv 0
  assign S_AXIS_DIN_TDATA_in[435] = (S_AXIS_DIN_TDATA[435] !== 1'bz) && S_AXIS_DIN_TDATA_delay[435]; // rv 0
  assign S_AXIS_DIN_TDATA_in[436] = (S_AXIS_DIN_TDATA[436] !== 1'bz) && S_AXIS_DIN_TDATA_delay[436]; // rv 0
  assign S_AXIS_DIN_TDATA_in[437] = (S_AXIS_DIN_TDATA[437] !== 1'bz) && S_AXIS_DIN_TDATA_delay[437]; // rv 0
  assign S_AXIS_DIN_TDATA_in[438] = (S_AXIS_DIN_TDATA[438] !== 1'bz) && S_AXIS_DIN_TDATA_delay[438]; // rv 0
  assign S_AXIS_DIN_TDATA_in[439] = (S_AXIS_DIN_TDATA[439] !== 1'bz) && S_AXIS_DIN_TDATA_delay[439]; // rv 0
  assign S_AXIS_DIN_TDATA_in[43] = (S_AXIS_DIN_TDATA[43] !== 1'bz) && S_AXIS_DIN_TDATA_delay[43]; // rv 0
  assign S_AXIS_DIN_TDATA_in[440] = (S_AXIS_DIN_TDATA[440] !== 1'bz) && S_AXIS_DIN_TDATA_delay[440]; // rv 0
  assign S_AXIS_DIN_TDATA_in[441] = (S_AXIS_DIN_TDATA[441] !== 1'bz) && S_AXIS_DIN_TDATA_delay[441]; // rv 0
  assign S_AXIS_DIN_TDATA_in[442] = (S_AXIS_DIN_TDATA[442] !== 1'bz) && S_AXIS_DIN_TDATA_delay[442]; // rv 0
  assign S_AXIS_DIN_TDATA_in[443] = (S_AXIS_DIN_TDATA[443] !== 1'bz) && S_AXIS_DIN_TDATA_delay[443]; // rv 0
  assign S_AXIS_DIN_TDATA_in[444] = (S_AXIS_DIN_TDATA[444] !== 1'bz) && S_AXIS_DIN_TDATA_delay[444]; // rv 0
  assign S_AXIS_DIN_TDATA_in[445] = (S_AXIS_DIN_TDATA[445] !== 1'bz) && S_AXIS_DIN_TDATA_delay[445]; // rv 0
  assign S_AXIS_DIN_TDATA_in[446] = (S_AXIS_DIN_TDATA[446] !== 1'bz) && S_AXIS_DIN_TDATA_delay[446]; // rv 0
  assign S_AXIS_DIN_TDATA_in[447] = (S_AXIS_DIN_TDATA[447] !== 1'bz) && S_AXIS_DIN_TDATA_delay[447]; // rv 0
  assign S_AXIS_DIN_TDATA_in[448] = (S_AXIS_DIN_TDATA[448] !== 1'bz) && S_AXIS_DIN_TDATA_delay[448]; // rv 0
  assign S_AXIS_DIN_TDATA_in[449] = (S_AXIS_DIN_TDATA[449] !== 1'bz) && S_AXIS_DIN_TDATA_delay[449]; // rv 0
  assign S_AXIS_DIN_TDATA_in[44] = (S_AXIS_DIN_TDATA[44] !== 1'bz) && S_AXIS_DIN_TDATA_delay[44]; // rv 0
  assign S_AXIS_DIN_TDATA_in[450] = (S_AXIS_DIN_TDATA[450] !== 1'bz) && S_AXIS_DIN_TDATA_delay[450]; // rv 0
  assign S_AXIS_DIN_TDATA_in[451] = (S_AXIS_DIN_TDATA[451] !== 1'bz) && S_AXIS_DIN_TDATA_delay[451]; // rv 0
  assign S_AXIS_DIN_TDATA_in[452] = (S_AXIS_DIN_TDATA[452] !== 1'bz) && S_AXIS_DIN_TDATA_delay[452]; // rv 0
  assign S_AXIS_DIN_TDATA_in[453] = (S_AXIS_DIN_TDATA[453] !== 1'bz) && S_AXIS_DIN_TDATA_delay[453]; // rv 0
  assign S_AXIS_DIN_TDATA_in[454] = (S_AXIS_DIN_TDATA[454] !== 1'bz) && S_AXIS_DIN_TDATA_delay[454]; // rv 0
  assign S_AXIS_DIN_TDATA_in[455] = (S_AXIS_DIN_TDATA[455] !== 1'bz) && S_AXIS_DIN_TDATA_delay[455]; // rv 0
  assign S_AXIS_DIN_TDATA_in[456] = (S_AXIS_DIN_TDATA[456] !== 1'bz) && S_AXIS_DIN_TDATA_delay[456]; // rv 0
  assign S_AXIS_DIN_TDATA_in[457] = (S_AXIS_DIN_TDATA[457] !== 1'bz) && S_AXIS_DIN_TDATA_delay[457]; // rv 0
  assign S_AXIS_DIN_TDATA_in[458] = (S_AXIS_DIN_TDATA[458] !== 1'bz) && S_AXIS_DIN_TDATA_delay[458]; // rv 0
  assign S_AXIS_DIN_TDATA_in[459] = (S_AXIS_DIN_TDATA[459] !== 1'bz) && S_AXIS_DIN_TDATA_delay[459]; // rv 0
  assign S_AXIS_DIN_TDATA_in[45] = (S_AXIS_DIN_TDATA[45] !== 1'bz) && S_AXIS_DIN_TDATA_delay[45]; // rv 0
  assign S_AXIS_DIN_TDATA_in[460] = (S_AXIS_DIN_TDATA[460] !== 1'bz) && S_AXIS_DIN_TDATA_delay[460]; // rv 0
  assign S_AXIS_DIN_TDATA_in[461] = (S_AXIS_DIN_TDATA[461] !== 1'bz) && S_AXIS_DIN_TDATA_delay[461]; // rv 0
  assign S_AXIS_DIN_TDATA_in[462] = (S_AXIS_DIN_TDATA[462] !== 1'bz) && S_AXIS_DIN_TDATA_delay[462]; // rv 0
  assign S_AXIS_DIN_TDATA_in[463] = (S_AXIS_DIN_TDATA[463] !== 1'bz) && S_AXIS_DIN_TDATA_delay[463]; // rv 0
  assign S_AXIS_DIN_TDATA_in[464] = (S_AXIS_DIN_TDATA[464] !== 1'bz) && S_AXIS_DIN_TDATA_delay[464]; // rv 0
  assign S_AXIS_DIN_TDATA_in[465] = (S_AXIS_DIN_TDATA[465] !== 1'bz) && S_AXIS_DIN_TDATA_delay[465]; // rv 0
  assign S_AXIS_DIN_TDATA_in[466] = (S_AXIS_DIN_TDATA[466] !== 1'bz) && S_AXIS_DIN_TDATA_delay[466]; // rv 0
  assign S_AXIS_DIN_TDATA_in[467] = (S_AXIS_DIN_TDATA[467] !== 1'bz) && S_AXIS_DIN_TDATA_delay[467]; // rv 0
  assign S_AXIS_DIN_TDATA_in[468] = (S_AXIS_DIN_TDATA[468] !== 1'bz) && S_AXIS_DIN_TDATA_delay[468]; // rv 0
  assign S_AXIS_DIN_TDATA_in[469] = (S_AXIS_DIN_TDATA[469] !== 1'bz) && S_AXIS_DIN_TDATA_delay[469]; // rv 0
  assign S_AXIS_DIN_TDATA_in[46] = (S_AXIS_DIN_TDATA[46] !== 1'bz) && S_AXIS_DIN_TDATA_delay[46]; // rv 0
  assign S_AXIS_DIN_TDATA_in[470] = (S_AXIS_DIN_TDATA[470] !== 1'bz) && S_AXIS_DIN_TDATA_delay[470]; // rv 0
  assign S_AXIS_DIN_TDATA_in[471] = (S_AXIS_DIN_TDATA[471] !== 1'bz) && S_AXIS_DIN_TDATA_delay[471]; // rv 0
  assign S_AXIS_DIN_TDATA_in[472] = (S_AXIS_DIN_TDATA[472] !== 1'bz) && S_AXIS_DIN_TDATA_delay[472]; // rv 0
  assign S_AXIS_DIN_TDATA_in[473] = (S_AXIS_DIN_TDATA[473] !== 1'bz) && S_AXIS_DIN_TDATA_delay[473]; // rv 0
  assign S_AXIS_DIN_TDATA_in[474] = (S_AXIS_DIN_TDATA[474] !== 1'bz) && S_AXIS_DIN_TDATA_delay[474]; // rv 0
  assign S_AXIS_DIN_TDATA_in[475] = (S_AXIS_DIN_TDATA[475] !== 1'bz) && S_AXIS_DIN_TDATA_delay[475]; // rv 0
  assign S_AXIS_DIN_TDATA_in[476] = (S_AXIS_DIN_TDATA[476] !== 1'bz) && S_AXIS_DIN_TDATA_delay[476]; // rv 0
  assign S_AXIS_DIN_TDATA_in[477] = (S_AXIS_DIN_TDATA[477] !== 1'bz) && S_AXIS_DIN_TDATA_delay[477]; // rv 0
  assign S_AXIS_DIN_TDATA_in[478] = (S_AXIS_DIN_TDATA[478] !== 1'bz) && S_AXIS_DIN_TDATA_delay[478]; // rv 0
  assign S_AXIS_DIN_TDATA_in[479] = (S_AXIS_DIN_TDATA[479] !== 1'bz) && S_AXIS_DIN_TDATA_delay[479]; // rv 0
  assign S_AXIS_DIN_TDATA_in[47] = (S_AXIS_DIN_TDATA[47] !== 1'bz) && S_AXIS_DIN_TDATA_delay[47]; // rv 0
  assign S_AXIS_DIN_TDATA_in[480] = (S_AXIS_DIN_TDATA[480] !== 1'bz) && S_AXIS_DIN_TDATA_delay[480]; // rv 0
  assign S_AXIS_DIN_TDATA_in[481] = (S_AXIS_DIN_TDATA[481] !== 1'bz) && S_AXIS_DIN_TDATA_delay[481]; // rv 0
  assign S_AXIS_DIN_TDATA_in[482] = (S_AXIS_DIN_TDATA[482] !== 1'bz) && S_AXIS_DIN_TDATA_delay[482]; // rv 0
  assign S_AXIS_DIN_TDATA_in[483] = (S_AXIS_DIN_TDATA[483] !== 1'bz) && S_AXIS_DIN_TDATA_delay[483]; // rv 0
  assign S_AXIS_DIN_TDATA_in[484] = (S_AXIS_DIN_TDATA[484] !== 1'bz) && S_AXIS_DIN_TDATA_delay[484]; // rv 0
  assign S_AXIS_DIN_TDATA_in[485] = (S_AXIS_DIN_TDATA[485] !== 1'bz) && S_AXIS_DIN_TDATA_delay[485]; // rv 0
  assign S_AXIS_DIN_TDATA_in[486] = (S_AXIS_DIN_TDATA[486] !== 1'bz) && S_AXIS_DIN_TDATA_delay[486]; // rv 0
  assign S_AXIS_DIN_TDATA_in[487] = (S_AXIS_DIN_TDATA[487] !== 1'bz) && S_AXIS_DIN_TDATA_delay[487]; // rv 0
  assign S_AXIS_DIN_TDATA_in[488] = (S_AXIS_DIN_TDATA[488] !== 1'bz) && S_AXIS_DIN_TDATA_delay[488]; // rv 0
  assign S_AXIS_DIN_TDATA_in[489] = (S_AXIS_DIN_TDATA[489] !== 1'bz) && S_AXIS_DIN_TDATA_delay[489]; // rv 0
  assign S_AXIS_DIN_TDATA_in[48] = (S_AXIS_DIN_TDATA[48] !== 1'bz) && S_AXIS_DIN_TDATA_delay[48]; // rv 0
  assign S_AXIS_DIN_TDATA_in[490] = (S_AXIS_DIN_TDATA[490] !== 1'bz) && S_AXIS_DIN_TDATA_delay[490]; // rv 0
  assign S_AXIS_DIN_TDATA_in[491] = (S_AXIS_DIN_TDATA[491] !== 1'bz) && S_AXIS_DIN_TDATA_delay[491]; // rv 0
  assign S_AXIS_DIN_TDATA_in[492] = (S_AXIS_DIN_TDATA[492] !== 1'bz) && S_AXIS_DIN_TDATA_delay[492]; // rv 0
  assign S_AXIS_DIN_TDATA_in[493] = (S_AXIS_DIN_TDATA[493] !== 1'bz) && S_AXIS_DIN_TDATA_delay[493]; // rv 0
  assign S_AXIS_DIN_TDATA_in[494] = (S_AXIS_DIN_TDATA[494] !== 1'bz) && S_AXIS_DIN_TDATA_delay[494]; // rv 0
  assign S_AXIS_DIN_TDATA_in[495] = (S_AXIS_DIN_TDATA[495] !== 1'bz) && S_AXIS_DIN_TDATA_delay[495]; // rv 0
  assign S_AXIS_DIN_TDATA_in[496] = (S_AXIS_DIN_TDATA[496] !== 1'bz) && S_AXIS_DIN_TDATA_delay[496]; // rv 0
  assign S_AXIS_DIN_TDATA_in[497] = (S_AXIS_DIN_TDATA[497] !== 1'bz) && S_AXIS_DIN_TDATA_delay[497]; // rv 0
  assign S_AXIS_DIN_TDATA_in[498] = (S_AXIS_DIN_TDATA[498] !== 1'bz) && S_AXIS_DIN_TDATA_delay[498]; // rv 0
  assign S_AXIS_DIN_TDATA_in[499] = (S_AXIS_DIN_TDATA[499] !== 1'bz) && S_AXIS_DIN_TDATA_delay[499]; // rv 0
  assign S_AXIS_DIN_TDATA_in[49] = (S_AXIS_DIN_TDATA[49] !== 1'bz) && S_AXIS_DIN_TDATA_delay[49]; // rv 0
  assign S_AXIS_DIN_TDATA_in[4] = (S_AXIS_DIN_TDATA[4] !== 1'bz) && S_AXIS_DIN_TDATA_delay[4]; // rv 0
  assign S_AXIS_DIN_TDATA_in[500] = (S_AXIS_DIN_TDATA[500] !== 1'bz) && S_AXIS_DIN_TDATA_delay[500]; // rv 0
  assign S_AXIS_DIN_TDATA_in[501] = (S_AXIS_DIN_TDATA[501] !== 1'bz) && S_AXIS_DIN_TDATA_delay[501]; // rv 0
  assign S_AXIS_DIN_TDATA_in[502] = (S_AXIS_DIN_TDATA[502] !== 1'bz) && S_AXIS_DIN_TDATA_delay[502]; // rv 0
  assign S_AXIS_DIN_TDATA_in[503] = (S_AXIS_DIN_TDATA[503] !== 1'bz) && S_AXIS_DIN_TDATA_delay[503]; // rv 0
  assign S_AXIS_DIN_TDATA_in[504] = (S_AXIS_DIN_TDATA[504] !== 1'bz) && S_AXIS_DIN_TDATA_delay[504]; // rv 0
  assign S_AXIS_DIN_TDATA_in[505] = (S_AXIS_DIN_TDATA[505] !== 1'bz) && S_AXIS_DIN_TDATA_delay[505]; // rv 0
  assign S_AXIS_DIN_TDATA_in[506] = (S_AXIS_DIN_TDATA[506] !== 1'bz) && S_AXIS_DIN_TDATA_delay[506]; // rv 0
  assign S_AXIS_DIN_TDATA_in[507] = (S_AXIS_DIN_TDATA[507] !== 1'bz) && S_AXIS_DIN_TDATA_delay[507]; // rv 0
  assign S_AXIS_DIN_TDATA_in[508] = (S_AXIS_DIN_TDATA[508] !== 1'bz) && S_AXIS_DIN_TDATA_delay[508]; // rv 0
  assign S_AXIS_DIN_TDATA_in[509] = (S_AXIS_DIN_TDATA[509] !== 1'bz) && S_AXIS_DIN_TDATA_delay[509]; // rv 0
  assign S_AXIS_DIN_TDATA_in[50] = (S_AXIS_DIN_TDATA[50] !== 1'bz) && S_AXIS_DIN_TDATA_delay[50]; // rv 0
  assign S_AXIS_DIN_TDATA_in[510] = (S_AXIS_DIN_TDATA[510] !== 1'bz) && S_AXIS_DIN_TDATA_delay[510]; // rv 0
  assign S_AXIS_DIN_TDATA_in[511] = (S_AXIS_DIN_TDATA[511] !== 1'bz) && S_AXIS_DIN_TDATA_delay[511]; // rv 0
  assign S_AXIS_DIN_TDATA_in[51] = (S_AXIS_DIN_TDATA[51] !== 1'bz) && S_AXIS_DIN_TDATA_delay[51]; // rv 0
  assign S_AXIS_DIN_TDATA_in[52] = (S_AXIS_DIN_TDATA[52] !== 1'bz) && S_AXIS_DIN_TDATA_delay[52]; // rv 0
  assign S_AXIS_DIN_TDATA_in[53] = (S_AXIS_DIN_TDATA[53] !== 1'bz) && S_AXIS_DIN_TDATA_delay[53]; // rv 0
  assign S_AXIS_DIN_TDATA_in[54] = (S_AXIS_DIN_TDATA[54] !== 1'bz) && S_AXIS_DIN_TDATA_delay[54]; // rv 0
  assign S_AXIS_DIN_TDATA_in[55] = (S_AXIS_DIN_TDATA[55] !== 1'bz) && S_AXIS_DIN_TDATA_delay[55]; // rv 0
  assign S_AXIS_DIN_TDATA_in[56] = (S_AXIS_DIN_TDATA[56] !== 1'bz) && S_AXIS_DIN_TDATA_delay[56]; // rv 0
  assign S_AXIS_DIN_TDATA_in[57] = (S_AXIS_DIN_TDATA[57] !== 1'bz) && S_AXIS_DIN_TDATA_delay[57]; // rv 0
  assign S_AXIS_DIN_TDATA_in[58] = (S_AXIS_DIN_TDATA[58] !== 1'bz) && S_AXIS_DIN_TDATA_delay[58]; // rv 0
  assign S_AXIS_DIN_TDATA_in[59] = (S_AXIS_DIN_TDATA[59] !== 1'bz) && S_AXIS_DIN_TDATA_delay[59]; // rv 0
  assign S_AXIS_DIN_TDATA_in[5] = (S_AXIS_DIN_TDATA[5] !== 1'bz) && S_AXIS_DIN_TDATA_delay[5]; // rv 0
  assign S_AXIS_DIN_TDATA_in[60] = (S_AXIS_DIN_TDATA[60] !== 1'bz) && S_AXIS_DIN_TDATA_delay[60]; // rv 0
  assign S_AXIS_DIN_TDATA_in[61] = (S_AXIS_DIN_TDATA[61] !== 1'bz) && S_AXIS_DIN_TDATA_delay[61]; // rv 0
  assign S_AXIS_DIN_TDATA_in[62] = (S_AXIS_DIN_TDATA[62] !== 1'bz) && S_AXIS_DIN_TDATA_delay[62]; // rv 0
  assign S_AXIS_DIN_TDATA_in[63] = (S_AXIS_DIN_TDATA[63] !== 1'bz) && S_AXIS_DIN_TDATA_delay[63]; // rv 0
  assign S_AXIS_DIN_TDATA_in[64] = (S_AXIS_DIN_TDATA[64] !== 1'bz) && S_AXIS_DIN_TDATA_delay[64]; // rv 0
  assign S_AXIS_DIN_TDATA_in[65] = (S_AXIS_DIN_TDATA[65] !== 1'bz) && S_AXIS_DIN_TDATA_delay[65]; // rv 0
  assign S_AXIS_DIN_TDATA_in[66] = (S_AXIS_DIN_TDATA[66] !== 1'bz) && S_AXIS_DIN_TDATA_delay[66]; // rv 0
  assign S_AXIS_DIN_TDATA_in[67] = (S_AXIS_DIN_TDATA[67] !== 1'bz) && S_AXIS_DIN_TDATA_delay[67]; // rv 0
  assign S_AXIS_DIN_TDATA_in[68] = (S_AXIS_DIN_TDATA[68] !== 1'bz) && S_AXIS_DIN_TDATA_delay[68]; // rv 0
  assign S_AXIS_DIN_TDATA_in[69] = (S_AXIS_DIN_TDATA[69] !== 1'bz) && S_AXIS_DIN_TDATA_delay[69]; // rv 0
  assign S_AXIS_DIN_TDATA_in[6] = (S_AXIS_DIN_TDATA[6] !== 1'bz) && S_AXIS_DIN_TDATA_delay[6]; // rv 0
  assign S_AXIS_DIN_TDATA_in[70] = (S_AXIS_DIN_TDATA[70] !== 1'bz) && S_AXIS_DIN_TDATA_delay[70]; // rv 0
  assign S_AXIS_DIN_TDATA_in[71] = (S_AXIS_DIN_TDATA[71] !== 1'bz) && S_AXIS_DIN_TDATA_delay[71]; // rv 0
  assign S_AXIS_DIN_TDATA_in[72] = (S_AXIS_DIN_TDATA[72] !== 1'bz) && S_AXIS_DIN_TDATA_delay[72]; // rv 0
  assign S_AXIS_DIN_TDATA_in[73] = (S_AXIS_DIN_TDATA[73] !== 1'bz) && S_AXIS_DIN_TDATA_delay[73]; // rv 0
  assign S_AXIS_DIN_TDATA_in[74] = (S_AXIS_DIN_TDATA[74] !== 1'bz) && S_AXIS_DIN_TDATA_delay[74]; // rv 0
  assign S_AXIS_DIN_TDATA_in[75] = (S_AXIS_DIN_TDATA[75] !== 1'bz) && S_AXIS_DIN_TDATA_delay[75]; // rv 0
  assign S_AXIS_DIN_TDATA_in[76] = (S_AXIS_DIN_TDATA[76] !== 1'bz) && S_AXIS_DIN_TDATA_delay[76]; // rv 0
  assign S_AXIS_DIN_TDATA_in[77] = (S_AXIS_DIN_TDATA[77] !== 1'bz) && S_AXIS_DIN_TDATA_delay[77]; // rv 0
  assign S_AXIS_DIN_TDATA_in[78] = (S_AXIS_DIN_TDATA[78] !== 1'bz) && S_AXIS_DIN_TDATA_delay[78]; // rv 0
  assign S_AXIS_DIN_TDATA_in[79] = (S_AXIS_DIN_TDATA[79] !== 1'bz) && S_AXIS_DIN_TDATA_delay[79]; // rv 0
  assign S_AXIS_DIN_TDATA_in[7] = (S_AXIS_DIN_TDATA[7] !== 1'bz) && S_AXIS_DIN_TDATA_delay[7]; // rv 0
  assign S_AXIS_DIN_TDATA_in[80] = (S_AXIS_DIN_TDATA[80] !== 1'bz) && S_AXIS_DIN_TDATA_delay[80]; // rv 0
  assign S_AXIS_DIN_TDATA_in[81] = (S_AXIS_DIN_TDATA[81] !== 1'bz) && S_AXIS_DIN_TDATA_delay[81]; // rv 0
  assign S_AXIS_DIN_TDATA_in[82] = (S_AXIS_DIN_TDATA[82] !== 1'bz) && S_AXIS_DIN_TDATA_delay[82]; // rv 0
  assign S_AXIS_DIN_TDATA_in[83] = (S_AXIS_DIN_TDATA[83] !== 1'bz) && S_AXIS_DIN_TDATA_delay[83]; // rv 0
  assign S_AXIS_DIN_TDATA_in[84] = (S_AXIS_DIN_TDATA[84] !== 1'bz) && S_AXIS_DIN_TDATA_delay[84]; // rv 0
  assign S_AXIS_DIN_TDATA_in[85] = (S_AXIS_DIN_TDATA[85] !== 1'bz) && S_AXIS_DIN_TDATA_delay[85]; // rv 0
  assign S_AXIS_DIN_TDATA_in[86] = (S_AXIS_DIN_TDATA[86] !== 1'bz) && S_AXIS_DIN_TDATA_delay[86]; // rv 0
  assign S_AXIS_DIN_TDATA_in[87] = (S_AXIS_DIN_TDATA[87] !== 1'bz) && S_AXIS_DIN_TDATA_delay[87]; // rv 0
  assign S_AXIS_DIN_TDATA_in[88] = (S_AXIS_DIN_TDATA[88] !== 1'bz) && S_AXIS_DIN_TDATA_delay[88]; // rv 0
  assign S_AXIS_DIN_TDATA_in[89] = (S_AXIS_DIN_TDATA[89] !== 1'bz) && S_AXIS_DIN_TDATA_delay[89]; // rv 0
  assign S_AXIS_DIN_TDATA_in[8] = (S_AXIS_DIN_TDATA[8] !== 1'bz) && S_AXIS_DIN_TDATA_delay[8]; // rv 0
  assign S_AXIS_DIN_TDATA_in[90] = (S_AXIS_DIN_TDATA[90] !== 1'bz) && S_AXIS_DIN_TDATA_delay[90]; // rv 0
  assign S_AXIS_DIN_TDATA_in[91] = (S_AXIS_DIN_TDATA[91] !== 1'bz) && S_AXIS_DIN_TDATA_delay[91]; // rv 0
  assign S_AXIS_DIN_TDATA_in[92] = (S_AXIS_DIN_TDATA[92] !== 1'bz) && S_AXIS_DIN_TDATA_delay[92]; // rv 0
  assign S_AXIS_DIN_TDATA_in[93] = (S_AXIS_DIN_TDATA[93] !== 1'bz) && S_AXIS_DIN_TDATA_delay[93]; // rv 0
  assign S_AXIS_DIN_TDATA_in[94] = (S_AXIS_DIN_TDATA[94] !== 1'bz) && S_AXIS_DIN_TDATA_delay[94]; // rv 0
  assign S_AXIS_DIN_TDATA_in[95] = (S_AXIS_DIN_TDATA[95] !== 1'bz) && S_AXIS_DIN_TDATA_delay[95]; // rv 0
  assign S_AXIS_DIN_TDATA_in[96] = (S_AXIS_DIN_TDATA[96] !== 1'bz) && S_AXIS_DIN_TDATA_delay[96]; // rv 0
  assign S_AXIS_DIN_TDATA_in[97] = (S_AXIS_DIN_TDATA[97] !== 1'bz) && S_AXIS_DIN_TDATA_delay[97]; // rv 0
  assign S_AXIS_DIN_TDATA_in[98] = (S_AXIS_DIN_TDATA[98] !== 1'bz) && S_AXIS_DIN_TDATA_delay[98]; // rv 0
  assign S_AXIS_DIN_TDATA_in[99] = (S_AXIS_DIN_TDATA[99] !== 1'bz) && S_AXIS_DIN_TDATA_delay[99]; // rv 0
  assign S_AXIS_DIN_TDATA_in[9] = (S_AXIS_DIN_TDATA[9] !== 1'bz) && S_AXIS_DIN_TDATA_delay[9]; // rv 0
  assign S_AXIS_DIN_TLAST_in = (S_AXIS_DIN_TLAST !== 1'bz) && S_AXIS_DIN_TLAST_delay; // rv 0
  assign S_AXIS_DIN_TVALID_in = (S_AXIS_DIN_TVALID !== 1'bz) && S_AXIS_DIN_TVALID_delay; // rv 0
  assign S_AXIS_DIN_WORDS_ACLK_in = (S_AXIS_DIN_WORDS_ACLK !== 1'bz) && S_AXIS_DIN_WORDS_ACLK_delay; // rv 0
  assign S_AXIS_DIN_WORDS_TDATA_in[0] = (S_AXIS_DIN_WORDS_TDATA[0] !== 1'bz) && S_AXIS_DIN_WORDS_TDATA_delay[0]; // rv 0
  assign S_AXIS_DIN_WORDS_TDATA_in[10] = (S_AXIS_DIN_WORDS_TDATA[10] !== 1'bz) && S_AXIS_DIN_WORDS_TDATA_delay[10]; // rv 0
  assign S_AXIS_DIN_WORDS_TDATA_in[11] = (S_AXIS_DIN_WORDS_TDATA[11] !== 1'bz) && S_AXIS_DIN_WORDS_TDATA_delay[11]; // rv 0
  assign S_AXIS_DIN_WORDS_TDATA_in[12] = (S_AXIS_DIN_WORDS_TDATA[12] !== 1'bz) && S_AXIS_DIN_WORDS_TDATA_delay[12]; // rv 0
  assign S_AXIS_DIN_WORDS_TDATA_in[13] = (S_AXIS_DIN_WORDS_TDATA[13] !== 1'bz) && S_AXIS_DIN_WORDS_TDATA_delay[13]; // rv 0
  assign S_AXIS_DIN_WORDS_TDATA_in[14] = (S_AXIS_DIN_WORDS_TDATA[14] !== 1'bz) && S_AXIS_DIN_WORDS_TDATA_delay[14]; // rv 0
  assign S_AXIS_DIN_WORDS_TDATA_in[15] = (S_AXIS_DIN_WORDS_TDATA[15] !== 1'bz) && S_AXIS_DIN_WORDS_TDATA_delay[15]; // rv 0
  assign S_AXIS_DIN_WORDS_TDATA_in[16] = (S_AXIS_DIN_WORDS_TDATA[16] !== 1'bz) && S_AXIS_DIN_WORDS_TDATA_delay[16]; // rv 0
  assign S_AXIS_DIN_WORDS_TDATA_in[17] = (S_AXIS_DIN_WORDS_TDATA[17] !== 1'bz) && S_AXIS_DIN_WORDS_TDATA_delay[17]; // rv 0
  assign S_AXIS_DIN_WORDS_TDATA_in[18] = (S_AXIS_DIN_WORDS_TDATA[18] !== 1'bz) && S_AXIS_DIN_WORDS_TDATA_delay[18]; // rv 0
  assign S_AXIS_DIN_WORDS_TDATA_in[19] = (S_AXIS_DIN_WORDS_TDATA[19] !== 1'bz) && S_AXIS_DIN_WORDS_TDATA_delay[19]; // rv 0
  assign S_AXIS_DIN_WORDS_TDATA_in[1] = (S_AXIS_DIN_WORDS_TDATA[1] !== 1'bz) && S_AXIS_DIN_WORDS_TDATA_delay[1]; // rv 0
  assign S_AXIS_DIN_WORDS_TDATA_in[20] = (S_AXIS_DIN_WORDS_TDATA[20] !== 1'bz) && S_AXIS_DIN_WORDS_TDATA_delay[20]; // rv 0
  assign S_AXIS_DIN_WORDS_TDATA_in[21] = (S_AXIS_DIN_WORDS_TDATA[21] !== 1'bz) && S_AXIS_DIN_WORDS_TDATA_delay[21]; // rv 0
  assign S_AXIS_DIN_WORDS_TDATA_in[22] = (S_AXIS_DIN_WORDS_TDATA[22] !== 1'bz) && S_AXIS_DIN_WORDS_TDATA_delay[22]; // rv 0
  assign S_AXIS_DIN_WORDS_TDATA_in[23] = (S_AXIS_DIN_WORDS_TDATA[23] !== 1'bz) && S_AXIS_DIN_WORDS_TDATA_delay[23]; // rv 0
  assign S_AXIS_DIN_WORDS_TDATA_in[24] = (S_AXIS_DIN_WORDS_TDATA[24] !== 1'bz) && S_AXIS_DIN_WORDS_TDATA_delay[24]; // rv 0
  assign S_AXIS_DIN_WORDS_TDATA_in[25] = (S_AXIS_DIN_WORDS_TDATA[25] !== 1'bz) && S_AXIS_DIN_WORDS_TDATA_delay[25]; // rv 0
  assign S_AXIS_DIN_WORDS_TDATA_in[26] = (S_AXIS_DIN_WORDS_TDATA[26] !== 1'bz) && S_AXIS_DIN_WORDS_TDATA_delay[26]; // rv 0
  assign S_AXIS_DIN_WORDS_TDATA_in[27] = (S_AXIS_DIN_WORDS_TDATA[27] !== 1'bz) && S_AXIS_DIN_WORDS_TDATA_delay[27]; // rv 0
  assign S_AXIS_DIN_WORDS_TDATA_in[28] = (S_AXIS_DIN_WORDS_TDATA[28] !== 1'bz) && S_AXIS_DIN_WORDS_TDATA_delay[28]; // rv 0
  assign S_AXIS_DIN_WORDS_TDATA_in[29] = (S_AXIS_DIN_WORDS_TDATA[29] !== 1'bz) && S_AXIS_DIN_WORDS_TDATA_delay[29]; // rv 0
  assign S_AXIS_DIN_WORDS_TDATA_in[2] = (S_AXIS_DIN_WORDS_TDATA[2] !== 1'bz) && S_AXIS_DIN_WORDS_TDATA_delay[2]; // rv 0
  assign S_AXIS_DIN_WORDS_TDATA_in[30] = (S_AXIS_DIN_WORDS_TDATA[30] !== 1'bz) && S_AXIS_DIN_WORDS_TDATA_delay[30]; // rv 0
  assign S_AXIS_DIN_WORDS_TDATA_in[31] = (S_AXIS_DIN_WORDS_TDATA[31] !== 1'bz) && S_AXIS_DIN_WORDS_TDATA_delay[31]; // rv 0
  assign S_AXIS_DIN_WORDS_TDATA_in[3] = (S_AXIS_DIN_WORDS_TDATA[3] !== 1'bz) && S_AXIS_DIN_WORDS_TDATA_delay[3]; // rv 0
  assign S_AXIS_DIN_WORDS_TDATA_in[4] = (S_AXIS_DIN_WORDS_TDATA[4] !== 1'bz) && S_AXIS_DIN_WORDS_TDATA_delay[4]; // rv 0
  assign S_AXIS_DIN_WORDS_TDATA_in[5] = (S_AXIS_DIN_WORDS_TDATA[5] !== 1'bz) && S_AXIS_DIN_WORDS_TDATA_delay[5]; // rv 0
  assign S_AXIS_DIN_WORDS_TDATA_in[6] = (S_AXIS_DIN_WORDS_TDATA[6] !== 1'bz) && S_AXIS_DIN_WORDS_TDATA_delay[6]; // rv 0
  assign S_AXIS_DIN_WORDS_TDATA_in[7] = (S_AXIS_DIN_WORDS_TDATA[7] !== 1'bz) && S_AXIS_DIN_WORDS_TDATA_delay[7]; // rv 0
  assign S_AXIS_DIN_WORDS_TDATA_in[8] = (S_AXIS_DIN_WORDS_TDATA[8] !== 1'bz) && S_AXIS_DIN_WORDS_TDATA_delay[8]; // rv 0
  assign S_AXIS_DIN_WORDS_TDATA_in[9] = (S_AXIS_DIN_WORDS_TDATA[9] !== 1'bz) && S_AXIS_DIN_WORDS_TDATA_delay[9]; // rv 0
  assign S_AXIS_DIN_WORDS_TLAST_in = (S_AXIS_DIN_WORDS_TLAST !== 1'bz) && S_AXIS_DIN_WORDS_TLAST_delay; // rv 0
  assign S_AXIS_DIN_WORDS_TVALID_in = (S_AXIS_DIN_WORDS_TVALID !== 1'bz) && S_AXIS_DIN_WORDS_TVALID_delay; // rv 0
  assign S_AXIS_DOUT_WORDS_ACLK_in = (S_AXIS_DOUT_WORDS_ACLK !== 1'bz) && S_AXIS_DOUT_WORDS_ACLK_delay; // rv 0
  assign S_AXIS_DOUT_WORDS_TDATA_in[0] = (S_AXIS_DOUT_WORDS_TDATA[0] !== 1'bz) && S_AXIS_DOUT_WORDS_TDATA_delay[0]; // rv 0
  assign S_AXIS_DOUT_WORDS_TDATA_in[10] = (S_AXIS_DOUT_WORDS_TDATA[10] !== 1'bz) && S_AXIS_DOUT_WORDS_TDATA_delay[10]; // rv 0
  assign S_AXIS_DOUT_WORDS_TDATA_in[11] = (S_AXIS_DOUT_WORDS_TDATA[11] !== 1'bz) && S_AXIS_DOUT_WORDS_TDATA_delay[11]; // rv 0
  assign S_AXIS_DOUT_WORDS_TDATA_in[12] = (S_AXIS_DOUT_WORDS_TDATA[12] !== 1'bz) && S_AXIS_DOUT_WORDS_TDATA_delay[12]; // rv 0
  assign S_AXIS_DOUT_WORDS_TDATA_in[13] = (S_AXIS_DOUT_WORDS_TDATA[13] !== 1'bz) && S_AXIS_DOUT_WORDS_TDATA_delay[13]; // rv 0
  assign S_AXIS_DOUT_WORDS_TDATA_in[14] = (S_AXIS_DOUT_WORDS_TDATA[14] !== 1'bz) && S_AXIS_DOUT_WORDS_TDATA_delay[14]; // rv 0
  assign S_AXIS_DOUT_WORDS_TDATA_in[15] = (S_AXIS_DOUT_WORDS_TDATA[15] !== 1'bz) && S_AXIS_DOUT_WORDS_TDATA_delay[15]; // rv 0
  assign S_AXIS_DOUT_WORDS_TDATA_in[16] = (S_AXIS_DOUT_WORDS_TDATA[16] !== 1'bz) && S_AXIS_DOUT_WORDS_TDATA_delay[16]; // rv 0
  assign S_AXIS_DOUT_WORDS_TDATA_in[17] = (S_AXIS_DOUT_WORDS_TDATA[17] !== 1'bz) && S_AXIS_DOUT_WORDS_TDATA_delay[17]; // rv 0
  assign S_AXIS_DOUT_WORDS_TDATA_in[18] = (S_AXIS_DOUT_WORDS_TDATA[18] !== 1'bz) && S_AXIS_DOUT_WORDS_TDATA_delay[18]; // rv 0
  assign S_AXIS_DOUT_WORDS_TDATA_in[19] = (S_AXIS_DOUT_WORDS_TDATA[19] !== 1'bz) && S_AXIS_DOUT_WORDS_TDATA_delay[19]; // rv 0
  assign S_AXIS_DOUT_WORDS_TDATA_in[1] = (S_AXIS_DOUT_WORDS_TDATA[1] !== 1'bz) && S_AXIS_DOUT_WORDS_TDATA_delay[1]; // rv 0
  assign S_AXIS_DOUT_WORDS_TDATA_in[20] = (S_AXIS_DOUT_WORDS_TDATA[20] !== 1'bz) && S_AXIS_DOUT_WORDS_TDATA_delay[20]; // rv 0
  assign S_AXIS_DOUT_WORDS_TDATA_in[21] = (S_AXIS_DOUT_WORDS_TDATA[21] !== 1'bz) && S_AXIS_DOUT_WORDS_TDATA_delay[21]; // rv 0
  assign S_AXIS_DOUT_WORDS_TDATA_in[22] = (S_AXIS_DOUT_WORDS_TDATA[22] !== 1'bz) && S_AXIS_DOUT_WORDS_TDATA_delay[22]; // rv 0
  assign S_AXIS_DOUT_WORDS_TDATA_in[23] = (S_AXIS_DOUT_WORDS_TDATA[23] !== 1'bz) && S_AXIS_DOUT_WORDS_TDATA_delay[23]; // rv 0
  assign S_AXIS_DOUT_WORDS_TDATA_in[24] = (S_AXIS_DOUT_WORDS_TDATA[24] !== 1'bz) && S_AXIS_DOUT_WORDS_TDATA_delay[24]; // rv 0
  assign S_AXIS_DOUT_WORDS_TDATA_in[25] = (S_AXIS_DOUT_WORDS_TDATA[25] !== 1'bz) && S_AXIS_DOUT_WORDS_TDATA_delay[25]; // rv 0
  assign S_AXIS_DOUT_WORDS_TDATA_in[26] = (S_AXIS_DOUT_WORDS_TDATA[26] !== 1'bz) && S_AXIS_DOUT_WORDS_TDATA_delay[26]; // rv 0
  assign S_AXIS_DOUT_WORDS_TDATA_in[27] = (S_AXIS_DOUT_WORDS_TDATA[27] !== 1'bz) && S_AXIS_DOUT_WORDS_TDATA_delay[27]; // rv 0
  assign S_AXIS_DOUT_WORDS_TDATA_in[28] = (S_AXIS_DOUT_WORDS_TDATA[28] !== 1'bz) && S_AXIS_DOUT_WORDS_TDATA_delay[28]; // rv 0
  assign S_AXIS_DOUT_WORDS_TDATA_in[29] = (S_AXIS_DOUT_WORDS_TDATA[29] !== 1'bz) && S_AXIS_DOUT_WORDS_TDATA_delay[29]; // rv 0
  assign S_AXIS_DOUT_WORDS_TDATA_in[2] = (S_AXIS_DOUT_WORDS_TDATA[2] !== 1'bz) && S_AXIS_DOUT_WORDS_TDATA_delay[2]; // rv 0
  assign S_AXIS_DOUT_WORDS_TDATA_in[30] = (S_AXIS_DOUT_WORDS_TDATA[30] !== 1'bz) && S_AXIS_DOUT_WORDS_TDATA_delay[30]; // rv 0
  assign S_AXIS_DOUT_WORDS_TDATA_in[31] = (S_AXIS_DOUT_WORDS_TDATA[31] !== 1'bz) && S_AXIS_DOUT_WORDS_TDATA_delay[31]; // rv 0
  assign S_AXIS_DOUT_WORDS_TDATA_in[3] = (S_AXIS_DOUT_WORDS_TDATA[3] !== 1'bz) && S_AXIS_DOUT_WORDS_TDATA_delay[3]; // rv 0
  assign S_AXIS_DOUT_WORDS_TDATA_in[4] = (S_AXIS_DOUT_WORDS_TDATA[4] !== 1'bz) && S_AXIS_DOUT_WORDS_TDATA_delay[4]; // rv 0
  assign S_AXIS_DOUT_WORDS_TDATA_in[5] = (S_AXIS_DOUT_WORDS_TDATA[5] !== 1'bz) && S_AXIS_DOUT_WORDS_TDATA_delay[5]; // rv 0
  assign S_AXIS_DOUT_WORDS_TDATA_in[6] = (S_AXIS_DOUT_WORDS_TDATA[6] !== 1'bz) && S_AXIS_DOUT_WORDS_TDATA_delay[6]; // rv 0
  assign S_AXIS_DOUT_WORDS_TDATA_in[7] = (S_AXIS_DOUT_WORDS_TDATA[7] !== 1'bz) && S_AXIS_DOUT_WORDS_TDATA_delay[7]; // rv 0
  assign S_AXIS_DOUT_WORDS_TDATA_in[8] = (S_AXIS_DOUT_WORDS_TDATA[8] !== 1'bz) && S_AXIS_DOUT_WORDS_TDATA_delay[8]; // rv 0
  assign S_AXIS_DOUT_WORDS_TDATA_in[9] = (S_AXIS_DOUT_WORDS_TDATA[9] !== 1'bz) && S_AXIS_DOUT_WORDS_TDATA_delay[9]; // rv 0
  assign S_AXIS_DOUT_WORDS_TLAST_in = (S_AXIS_DOUT_WORDS_TLAST !== 1'bz) && S_AXIS_DOUT_WORDS_TLAST_delay; // rv 0
  assign S_AXIS_DOUT_WORDS_TVALID_in = (S_AXIS_DOUT_WORDS_TVALID !== 1'bz) && S_AXIS_DOUT_WORDS_TVALID_delay; // rv 0
  assign S_AXI_ACLK_in = (S_AXI_ACLK !== 1'bz) && S_AXI_ACLK_delay; // rv 0
  assign S_AXI_ARADDR_in[0] = (S_AXI_ARADDR[0] !== 1'bz) && S_AXI_ARADDR_delay[0]; // rv 0
  assign S_AXI_ARADDR_in[10] = (S_AXI_ARADDR[10] !== 1'bz) && S_AXI_ARADDR_delay[10]; // rv 0
  assign S_AXI_ARADDR_in[11] = (S_AXI_ARADDR[11] !== 1'bz) && S_AXI_ARADDR_delay[11]; // rv 0
  assign S_AXI_ARADDR_in[12] = (S_AXI_ARADDR[12] !== 1'bz) && S_AXI_ARADDR_delay[12]; // rv 0
  assign S_AXI_ARADDR_in[13] = (S_AXI_ARADDR[13] !== 1'bz) && S_AXI_ARADDR_delay[13]; // rv 0
  assign S_AXI_ARADDR_in[14] = (S_AXI_ARADDR[14] !== 1'bz) && S_AXI_ARADDR_delay[14]; // rv 0
  assign S_AXI_ARADDR_in[15] = (S_AXI_ARADDR[15] !== 1'bz) && S_AXI_ARADDR_delay[15]; // rv 0
  assign S_AXI_ARADDR_in[16] = (S_AXI_ARADDR[16] !== 1'bz) && S_AXI_ARADDR_delay[16]; // rv 0
  assign S_AXI_ARADDR_in[17] = (S_AXI_ARADDR[17] !== 1'bz) && S_AXI_ARADDR_delay[17]; // rv 0
  assign S_AXI_ARADDR_in[1] = (S_AXI_ARADDR[1] !== 1'bz) && S_AXI_ARADDR_delay[1]; // rv 0
  assign S_AXI_ARADDR_in[2] = (S_AXI_ARADDR[2] !== 1'bz) && S_AXI_ARADDR_delay[2]; // rv 0
  assign S_AXI_ARADDR_in[3] = (S_AXI_ARADDR[3] !== 1'bz) && S_AXI_ARADDR_delay[3]; // rv 0
  assign S_AXI_ARADDR_in[4] = (S_AXI_ARADDR[4] !== 1'bz) && S_AXI_ARADDR_delay[4]; // rv 0
  assign S_AXI_ARADDR_in[5] = (S_AXI_ARADDR[5] !== 1'bz) && S_AXI_ARADDR_delay[5]; // rv 0
  assign S_AXI_ARADDR_in[6] = (S_AXI_ARADDR[6] !== 1'bz) && S_AXI_ARADDR_delay[6]; // rv 0
  assign S_AXI_ARADDR_in[7] = (S_AXI_ARADDR[7] !== 1'bz) && S_AXI_ARADDR_delay[7]; // rv 0
  assign S_AXI_ARADDR_in[8] = (S_AXI_ARADDR[8] !== 1'bz) && S_AXI_ARADDR_delay[8]; // rv 0
  assign S_AXI_ARADDR_in[9] = (S_AXI_ARADDR[9] !== 1'bz) && S_AXI_ARADDR_delay[9]; // rv 0
  assign S_AXI_ARVALID_in = (S_AXI_ARVALID !== 1'bz) && S_AXI_ARVALID_delay; // rv 0
  assign S_AXI_AWADDR_in[0] = (S_AXI_AWADDR[0] !== 1'bz) && S_AXI_AWADDR_delay[0]; // rv 0
  assign S_AXI_AWADDR_in[10] = (S_AXI_AWADDR[10] !== 1'bz) && S_AXI_AWADDR_delay[10]; // rv 0
  assign S_AXI_AWADDR_in[11] = (S_AXI_AWADDR[11] !== 1'bz) && S_AXI_AWADDR_delay[11]; // rv 0
  assign S_AXI_AWADDR_in[12] = (S_AXI_AWADDR[12] !== 1'bz) && S_AXI_AWADDR_delay[12]; // rv 0
  assign S_AXI_AWADDR_in[13] = (S_AXI_AWADDR[13] !== 1'bz) && S_AXI_AWADDR_delay[13]; // rv 0
  assign S_AXI_AWADDR_in[14] = (S_AXI_AWADDR[14] !== 1'bz) && S_AXI_AWADDR_delay[14]; // rv 0
  assign S_AXI_AWADDR_in[15] = (S_AXI_AWADDR[15] !== 1'bz) && S_AXI_AWADDR_delay[15]; // rv 0
  assign S_AXI_AWADDR_in[16] = (S_AXI_AWADDR[16] !== 1'bz) && S_AXI_AWADDR_delay[16]; // rv 0
  assign S_AXI_AWADDR_in[17] = (S_AXI_AWADDR[17] !== 1'bz) && S_AXI_AWADDR_delay[17]; // rv 0
  assign S_AXI_AWADDR_in[1] = (S_AXI_AWADDR[1] !== 1'bz) && S_AXI_AWADDR_delay[1]; // rv 0
  assign S_AXI_AWADDR_in[2] = (S_AXI_AWADDR[2] !== 1'bz) && S_AXI_AWADDR_delay[2]; // rv 0
  assign S_AXI_AWADDR_in[3] = (S_AXI_AWADDR[3] !== 1'bz) && S_AXI_AWADDR_delay[3]; // rv 0
  assign S_AXI_AWADDR_in[4] = (S_AXI_AWADDR[4] !== 1'bz) && S_AXI_AWADDR_delay[4]; // rv 0
  assign S_AXI_AWADDR_in[5] = (S_AXI_AWADDR[5] !== 1'bz) && S_AXI_AWADDR_delay[5]; // rv 0
  assign S_AXI_AWADDR_in[6] = (S_AXI_AWADDR[6] !== 1'bz) && S_AXI_AWADDR_delay[6]; // rv 0
  assign S_AXI_AWADDR_in[7] = (S_AXI_AWADDR[7] !== 1'bz) && S_AXI_AWADDR_delay[7]; // rv 0
  assign S_AXI_AWADDR_in[8] = (S_AXI_AWADDR[8] !== 1'bz) && S_AXI_AWADDR_delay[8]; // rv 0
  assign S_AXI_AWADDR_in[9] = (S_AXI_AWADDR[9] !== 1'bz) && S_AXI_AWADDR_delay[9]; // rv 0
  assign S_AXI_AWVALID_in = (S_AXI_AWVALID !== 1'bz) && S_AXI_AWVALID_delay; // rv 0
  assign S_AXI_BREADY_in = (S_AXI_BREADY !== 1'bz) && S_AXI_BREADY_delay; // rv 0
  assign S_AXI_RREADY_in = (S_AXI_RREADY !== 1'bz) && S_AXI_RREADY_delay; // rv 0
  assign S_AXI_WDATA_in[0] = (S_AXI_WDATA[0] !== 1'bz) && S_AXI_WDATA_delay[0]; // rv 0
  assign S_AXI_WDATA_in[10] = (S_AXI_WDATA[10] !== 1'bz) && S_AXI_WDATA_delay[10]; // rv 0
  assign S_AXI_WDATA_in[11] = (S_AXI_WDATA[11] !== 1'bz) && S_AXI_WDATA_delay[11]; // rv 0
  assign S_AXI_WDATA_in[12] = (S_AXI_WDATA[12] !== 1'bz) && S_AXI_WDATA_delay[12]; // rv 0
  assign S_AXI_WDATA_in[13] = (S_AXI_WDATA[13] !== 1'bz) && S_AXI_WDATA_delay[13]; // rv 0
  assign S_AXI_WDATA_in[14] = (S_AXI_WDATA[14] !== 1'bz) && S_AXI_WDATA_delay[14]; // rv 0
  assign S_AXI_WDATA_in[15] = (S_AXI_WDATA[15] !== 1'bz) && S_AXI_WDATA_delay[15]; // rv 0
  assign S_AXI_WDATA_in[16] = (S_AXI_WDATA[16] !== 1'bz) && S_AXI_WDATA_delay[16]; // rv 0
  assign S_AXI_WDATA_in[17] = (S_AXI_WDATA[17] !== 1'bz) && S_AXI_WDATA_delay[17]; // rv 0
  assign S_AXI_WDATA_in[18] = (S_AXI_WDATA[18] !== 1'bz) && S_AXI_WDATA_delay[18]; // rv 0
  assign S_AXI_WDATA_in[19] = (S_AXI_WDATA[19] !== 1'bz) && S_AXI_WDATA_delay[19]; // rv 0
  assign S_AXI_WDATA_in[1] = (S_AXI_WDATA[1] !== 1'bz) && S_AXI_WDATA_delay[1]; // rv 0
  assign S_AXI_WDATA_in[20] = (S_AXI_WDATA[20] !== 1'bz) && S_AXI_WDATA_delay[20]; // rv 0
  assign S_AXI_WDATA_in[21] = (S_AXI_WDATA[21] !== 1'bz) && S_AXI_WDATA_delay[21]; // rv 0
  assign S_AXI_WDATA_in[22] = (S_AXI_WDATA[22] !== 1'bz) && S_AXI_WDATA_delay[22]; // rv 0
  assign S_AXI_WDATA_in[23] = (S_AXI_WDATA[23] !== 1'bz) && S_AXI_WDATA_delay[23]; // rv 0
  assign S_AXI_WDATA_in[24] = (S_AXI_WDATA[24] !== 1'bz) && S_AXI_WDATA_delay[24]; // rv 0
  assign S_AXI_WDATA_in[25] = (S_AXI_WDATA[25] !== 1'bz) && S_AXI_WDATA_delay[25]; // rv 0
  assign S_AXI_WDATA_in[26] = (S_AXI_WDATA[26] !== 1'bz) && S_AXI_WDATA_delay[26]; // rv 0
  assign S_AXI_WDATA_in[27] = (S_AXI_WDATA[27] !== 1'bz) && S_AXI_WDATA_delay[27]; // rv 0
  assign S_AXI_WDATA_in[28] = (S_AXI_WDATA[28] !== 1'bz) && S_AXI_WDATA_delay[28]; // rv 0
  assign S_AXI_WDATA_in[29] = (S_AXI_WDATA[29] !== 1'bz) && S_AXI_WDATA_delay[29]; // rv 0
  assign S_AXI_WDATA_in[2] = (S_AXI_WDATA[2] !== 1'bz) && S_AXI_WDATA_delay[2]; // rv 0
  assign S_AXI_WDATA_in[30] = (S_AXI_WDATA[30] !== 1'bz) && S_AXI_WDATA_delay[30]; // rv 0
  assign S_AXI_WDATA_in[31] = (S_AXI_WDATA[31] !== 1'bz) && S_AXI_WDATA_delay[31]; // rv 0
  assign S_AXI_WDATA_in[3] = (S_AXI_WDATA[3] !== 1'bz) && S_AXI_WDATA_delay[3]; // rv 0
  assign S_AXI_WDATA_in[4] = (S_AXI_WDATA[4] !== 1'bz) && S_AXI_WDATA_delay[4]; // rv 0
  assign S_AXI_WDATA_in[5] = (S_AXI_WDATA[5] !== 1'bz) && S_AXI_WDATA_delay[5]; // rv 0
  assign S_AXI_WDATA_in[6] = (S_AXI_WDATA[6] !== 1'bz) && S_AXI_WDATA_delay[6]; // rv 0
  assign S_AXI_WDATA_in[7] = (S_AXI_WDATA[7] !== 1'bz) && S_AXI_WDATA_delay[7]; // rv 0
  assign S_AXI_WDATA_in[8] = (S_AXI_WDATA[8] !== 1'bz) && S_AXI_WDATA_delay[8]; // rv 0
  assign S_AXI_WDATA_in[9] = (S_AXI_WDATA[9] !== 1'bz) && S_AXI_WDATA_delay[9]; // rv 0
  assign S_AXI_WVALID_in = (S_AXI_WVALID !== 1'bz) && S_AXI_WVALID_delay; // rv 0
`else
  assign CORE_CLK_in = (CORE_CLK !== 1'bz) && CORE_CLK; // rv 0
  assign DEBUG_EN_in = (DEBUG_EN === 1'bz) || DEBUG_EN; // rv 1
  assign M_AXIS_DOUT_ACLK_in = (M_AXIS_DOUT_ACLK !== 1'bz) && M_AXIS_DOUT_ACLK; // rv 0
  assign M_AXIS_DOUT_TREADY_in = (M_AXIS_DOUT_TREADY !== 1'bz) && M_AXIS_DOUT_TREADY; // rv 0
  assign M_AXIS_STATUS_ACLK_in = (M_AXIS_STATUS_ACLK !== 1'bz) && M_AXIS_STATUS_ACLK; // rv 0
  assign M_AXIS_STATUS_TREADY_in = (M_AXIS_STATUS_TREADY !== 1'bz) && M_AXIS_STATUS_TREADY; // rv 0
  assign S_AXIS_CTRL_ACLK_in = (S_AXIS_CTRL_ACLK !== 1'bz) && S_AXIS_CTRL_ACLK; // rv 0
  assign S_AXIS_CTRL_TDATA_in[0] = (S_AXIS_CTRL_TDATA[0] !== 1'bz) && S_AXIS_CTRL_TDATA[0]; // rv 0
  assign S_AXIS_CTRL_TDATA_in[10] = (S_AXIS_CTRL_TDATA[10] !== 1'bz) && S_AXIS_CTRL_TDATA[10]; // rv 0
  assign S_AXIS_CTRL_TDATA_in[11] = (S_AXIS_CTRL_TDATA[11] !== 1'bz) && S_AXIS_CTRL_TDATA[11]; // rv 0
  assign S_AXIS_CTRL_TDATA_in[12] = (S_AXIS_CTRL_TDATA[12] !== 1'bz) && S_AXIS_CTRL_TDATA[12]; // rv 0
  assign S_AXIS_CTRL_TDATA_in[13] = (S_AXIS_CTRL_TDATA[13] !== 1'bz) && S_AXIS_CTRL_TDATA[13]; // rv 0
  assign S_AXIS_CTRL_TDATA_in[14] = (S_AXIS_CTRL_TDATA[14] !== 1'bz) && S_AXIS_CTRL_TDATA[14]; // rv 0
  assign S_AXIS_CTRL_TDATA_in[15] = (S_AXIS_CTRL_TDATA[15] !== 1'bz) && S_AXIS_CTRL_TDATA[15]; // rv 0
  assign S_AXIS_CTRL_TDATA_in[16] = (S_AXIS_CTRL_TDATA[16] !== 1'bz) && S_AXIS_CTRL_TDATA[16]; // rv 0
  assign S_AXIS_CTRL_TDATA_in[17] = (S_AXIS_CTRL_TDATA[17] !== 1'bz) && S_AXIS_CTRL_TDATA[17]; // rv 0
  assign S_AXIS_CTRL_TDATA_in[18] = (S_AXIS_CTRL_TDATA[18] !== 1'bz) && S_AXIS_CTRL_TDATA[18]; // rv 0
  assign S_AXIS_CTRL_TDATA_in[19] = (S_AXIS_CTRL_TDATA[19] !== 1'bz) && S_AXIS_CTRL_TDATA[19]; // rv 0
  assign S_AXIS_CTRL_TDATA_in[1] = (S_AXIS_CTRL_TDATA[1] !== 1'bz) && S_AXIS_CTRL_TDATA[1]; // rv 0
  assign S_AXIS_CTRL_TDATA_in[20] = (S_AXIS_CTRL_TDATA[20] !== 1'bz) && S_AXIS_CTRL_TDATA[20]; // rv 0
  assign S_AXIS_CTRL_TDATA_in[21] = (S_AXIS_CTRL_TDATA[21] !== 1'bz) && S_AXIS_CTRL_TDATA[21]; // rv 0
  assign S_AXIS_CTRL_TDATA_in[22] = (S_AXIS_CTRL_TDATA[22] !== 1'bz) && S_AXIS_CTRL_TDATA[22]; // rv 0
  assign S_AXIS_CTRL_TDATA_in[23] = (S_AXIS_CTRL_TDATA[23] !== 1'bz) && S_AXIS_CTRL_TDATA[23]; // rv 0
  assign S_AXIS_CTRL_TDATA_in[24] = (S_AXIS_CTRL_TDATA[24] !== 1'bz) && S_AXIS_CTRL_TDATA[24]; // rv 0
  assign S_AXIS_CTRL_TDATA_in[25] = (S_AXIS_CTRL_TDATA[25] !== 1'bz) && S_AXIS_CTRL_TDATA[25]; // rv 0
  assign S_AXIS_CTRL_TDATA_in[26] = (S_AXIS_CTRL_TDATA[26] !== 1'bz) && S_AXIS_CTRL_TDATA[26]; // rv 0
  assign S_AXIS_CTRL_TDATA_in[27] = (S_AXIS_CTRL_TDATA[27] !== 1'bz) && S_AXIS_CTRL_TDATA[27]; // rv 0
  assign S_AXIS_CTRL_TDATA_in[28] = (S_AXIS_CTRL_TDATA[28] !== 1'bz) && S_AXIS_CTRL_TDATA[28]; // rv 0
  assign S_AXIS_CTRL_TDATA_in[29] = (S_AXIS_CTRL_TDATA[29] !== 1'bz) && S_AXIS_CTRL_TDATA[29]; // rv 0
  assign S_AXIS_CTRL_TDATA_in[2] = (S_AXIS_CTRL_TDATA[2] !== 1'bz) && S_AXIS_CTRL_TDATA[2]; // rv 0
  assign S_AXIS_CTRL_TDATA_in[30] = (S_AXIS_CTRL_TDATA[30] !== 1'bz) && S_AXIS_CTRL_TDATA[30]; // rv 0
  assign S_AXIS_CTRL_TDATA_in[31] = (S_AXIS_CTRL_TDATA[31] !== 1'bz) && S_AXIS_CTRL_TDATA[31]; // rv 0
  assign S_AXIS_CTRL_TDATA_in[3] = (S_AXIS_CTRL_TDATA[3] !== 1'bz) && S_AXIS_CTRL_TDATA[3]; // rv 0
  assign S_AXIS_CTRL_TDATA_in[4] = (S_AXIS_CTRL_TDATA[4] !== 1'bz) && S_AXIS_CTRL_TDATA[4]; // rv 0
  assign S_AXIS_CTRL_TDATA_in[5] = (S_AXIS_CTRL_TDATA[5] !== 1'bz) && S_AXIS_CTRL_TDATA[5]; // rv 0
  assign S_AXIS_CTRL_TDATA_in[6] = (S_AXIS_CTRL_TDATA[6] !== 1'bz) && S_AXIS_CTRL_TDATA[6]; // rv 0
  assign S_AXIS_CTRL_TDATA_in[7] = (S_AXIS_CTRL_TDATA[7] !== 1'bz) && S_AXIS_CTRL_TDATA[7]; // rv 0
  assign S_AXIS_CTRL_TDATA_in[8] = (S_AXIS_CTRL_TDATA[8] !== 1'bz) && S_AXIS_CTRL_TDATA[8]; // rv 0
  assign S_AXIS_CTRL_TDATA_in[9] = (S_AXIS_CTRL_TDATA[9] !== 1'bz) && S_AXIS_CTRL_TDATA[9]; // rv 0
  assign S_AXIS_CTRL_TVALID_in = (S_AXIS_CTRL_TVALID !== 1'bz) && S_AXIS_CTRL_TVALID; // rv 0
  assign S_AXIS_DIN_ACLK_in = (S_AXIS_DIN_ACLK !== 1'bz) && S_AXIS_DIN_ACLK; // rv 0
  assign S_AXIS_DIN_TDATA_in[0] = (S_AXIS_DIN_TDATA[0] !== 1'bz) && S_AXIS_DIN_TDATA[0]; // rv 0
  assign S_AXIS_DIN_TDATA_in[100] = (S_AXIS_DIN_TDATA[100] !== 1'bz) && S_AXIS_DIN_TDATA[100]; // rv 0
  assign S_AXIS_DIN_TDATA_in[101] = (S_AXIS_DIN_TDATA[101] !== 1'bz) && S_AXIS_DIN_TDATA[101]; // rv 0
  assign S_AXIS_DIN_TDATA_in[102] = (S_AXIS_DIN_TDATA[102] !== 1'bz) && S_AXIS_DIN_TDATA[102]; // rv 0
  assign S_AXIS_DIN_TDATA_in[103] = (S_AXIS_DIN_TDATA[103] !== 1'bz) && S_AXIS_DIN_TDATA[103]; // rv 0
  assign S_AXIS_DIN_TDATA_in[104] = (S_AXIS_DIN_TDATA[104] !== 1'bz) && S_AXIS_DIN_TDATA[104]; // rv 0
  assign S_AXIS_DIN_TDATA_in[105] = (S_AXIS_DIN_TDATA[105] !== 1'bz) && S_AXIS_DIN_TDATA[105]; // rv 0
  assign S_AXIS_DIN_TDATA_in[106] = (S_AXIS_DIN_TDATA[106] !== 1'bz) && S_AXIS_DIN_TDATA[106]; // rv 0
  assign S_AXIS_DIN_TDATA_in[107] = (S_AXIS_DIN_TDATA[107] !== 1'bz) && S_AXIS_DIN_TDATA[107]; // rv 0
  assign S_AXIS_DIN_TDATA_in[108] = (S_AXIS_DIN_TDATA[108] !== 1'bz) && S_AXIS_DIN_TDATA[108]; // rv 0
  assign S_AXIS_DIN_TDATA_in[109] = (S_AXIS_DIN_TDATA[109] !== 1'bz) && S_AXIS_DIN_TDATA[109]; // rv 0
  assign S_AXIS_DIN_TDATA_in[10] = (S_AXIS_DIN_TDATA[10] !== 1'bz) && S_AXIS_DIN_TDATA[10]; // rv 0
  assign S_AXIS_DIN_TDATA_in[110] = (S_AXIS_DIN_TDATA[110] !== 1'bz) && S_AXIS_DIN_TDATA[110]; // rv 0
  assign S_AXIS_DIN_TDATA_in[111] = (S_AXIS_DIN_TDATA[111] !== 1'bz) && S_AXIS_DIN_TDATA[111]; // rv 0
  assign S_AXIS_DIN_TDATA_in[112] = (S_AXIS_DIN_TDATA[112] !== 1'bz) && S_AXIS_DIN_TDATA[112]; // rv 0
  assign S_AXIS_DIN_TDATA_in[113] = (S_AXIS_DIN_TDATA[113] !== 1'bz) && S_AXIS_DIN_TDATA[113]; // rv 0
  assign S_AXIS_DIN_TDATA_in[114] = (S_AXIS_DIN_TDATA[114] !== 1'bz) && S_AXIS_DIN_TDATA[114]; // rv 0
  assign S_AXIS_DIN_TDATA_in[115] = (S_AXIS_DIN_TDATA[115] !== 1'bz) && S_AXIS_DIN_TDATA[115]; // rv 0
  assign S_AXIS_DIN_TDATA_in[116] = (S_AXIS_DIN_TDATA[116] !== 1'bz) && S_AXIS_DIN_TDATA[116]; // rv 0
  assign S_AXIS_DIN_TDATA_in[117] = (S_AXIS_DIN_TDATA[117] !== 1'bz) && S_AXIS_DIN_TDATA[117]; // rv 0
  assign S_AXIS_DIN_TDATA_in[118] = (S_AXIS_DIN_TDATA[118] !== 1'bz) && S_AXIS_DIN_TDATA[118]; // rv 0
  assign S_AXIS_DIN_TDATA_in[119] = (S_AXIS_DIN_TDATA[119] !== 1'bz) && S_AXIS_DIN_TDATA[119]; // rv 0
  assign S_AXIS_DIN_TDATA_in[11] = (S_AXIS_DIN_TDATA[11] !== 1'bz) && S_AXIS_DIN_TDATA[11]; // rv 0
  assign S_AXIS_DIN_TDATA_in[120] = (S_AXIS_DIN_TDATA[120] !== 1'bz) && S_AXIS_DIN_TDATA[120]; // rv 0
  assign S_AXIS_DIN_TDATA_in[121] = (S_AXIS_DIN_TDATA[121] !== 1'bz) && S_AXIS_DIN_TDATA[121]; // rv 0
  assign S_AXIS_DIN_TDATA_in[122] = (S_AXIS_DIN_TDATA[122] !== 1'bz) && S_AXIS_DIN_TDATA[122]; // rv 0
  assign S_AXIS_DIN_TDATA_in[123] = (S_AXIS_DIN_TDATA[123] !== 1'bz) && S_AXIS_DIN_TDATA[123]; // rv 0
  assign S_AXIS_DIN_TDATA_in[124] = (S_AXIS_DIN_TDATA[124] !== 1'bz) && S_AXIS_DIN_TDATA[124]; // rv 0
  assign S_AXIS_DIN_TDATA_in[125] = (S_AXIS_DIN_TDATA[125] !== 1'bz) && S_AXIS_DIN_TDATA[125]; // rv 0
  assign S_AXIS_DIN_TDATA_in[126] = (S_AXIS_DIN_TDATA[126] !== 1'bz) && S_AXIS_DIN_TDATA[126]; // rv 0
  assign S_AXIS_DIN_TDATA_in[127] = (S_AXIS_DIN_TDATA[127] !== 1'bz) && S_AXIS_DIN_TDATA[127]; // rv 0
  assign S_AXIS_DIN_TDATA_in[128] = (S_AXIS_DIN_TDATA[128] !== 1'bz) && S_AXIS_DIN_TDATA[128]; // rv 0
  assign S_AXIS_DIN_TDATA_in[129] = (S_AXIS_DIN_TDATA[129] !== 1'bz) && S_AXIS_DIN_TDATA[129]; // rv 0
  assign S_AXIS_DIN_TDATA_in[12] = (S_AXIS_DIN_TDATA[12] !== 1'bz) && S_AXIS_DIN_TDATA[12]; // rv 0
  assign S_AXIS_DIN_TDATA_in[130] = (S_AXIS_DIN_TDATA[130] !== 1'bz) && S_AXIS_DIN_TDATA[130]; // rv 0
  assign S_AXIS_DIN_TDATA_in[131] = (S_AXIS_DIN_TDATA[131] !== 1'bz) && S_AXIS_DIN_TDATA[131]; // rv 0
  assign S_AXIS_DIN_TDATA_in[132] = (S_AXIS_DIN_TDATA[132] !== 1'bz) && S_AXIS_DIN_TDATA[132]; // rv 0
  assign S_AXIS_DIN_TDATA_in[133] = (S_AXIS_DIN_TDATA[133] !== 1'bz) && S_AXIS_DIN_TDATA[133]; // rv 0
  assign S_AXIS_DIN_TDATA_in[134] = (S_AXIS_DIN_TDATA[134] !== 1'bz) && S_AXIS_DIN_TDATA[134]; // rv 0
  assign S_AXIS_DIN_TDATA_in[135] = (S_AXIS_DIN_TDATA[135] !== 1'bz) && S_AXIS_DIN_TDATA[135]; // rv 0
  assign S_AXIS_DIN_TDATA_in[136] = (S_AXIS_DIN_TDATA[136] !== 1'bz) && S_AXIS_DIN_TDATA[136]; // rv 0
  assign S_AXIS_DIN_TDATA_in[137] = (S_AXIS_DIN_TDATA[137] !== 1'bz) && S_AXIS_DIN_TDATA[137]; // rv 0
  assign S_AXIS_DIN_TDATA_in[138] = (S_AXIS_DIN_TDATA[138] !== 1'bz) && S_AXIS_DIN_TDATA[138]; // rv 0
  assign S_AXIS_DIN_TDATA_in[139] = (S_AXIS_DIN_TDATA[139] !== 1'bz) && S_AXIS_DIN_TDATA[139]; // rv 0
  assign S_AXIS_DIN_TDATA_in[13] = (S_AXIS_DIN_TDATA[13] !== 1'bz) && S_AXIS_DIN_TDATA[13]; // rv 0
  assign S_AXIS_DIN_TDATA_in[140] = (S_AXIS_DIN_TDATA[140] !== 1'bz) && S_AXIS_DIN_TDATA[140]; // rv 0
  assign S_AXIS_DIN_TDATA_in[141] = (S_AXIS_DIN_TDATA[141] !== 1'bz) && S_AXIS_DIN_TDATA[141]; // rv 0
  assign S_AXIS_DIN_TDATA_in[142] = (S_AXIS_DIN_TDATA[142] !== 1'bz) && S_AXIS_DIN_TDATA[142]; // rv 0
  assign S_AXIS_DIN_TDATA_in[143] = (S_AXIS_DIN_TDATA[143] !== 1'bz) && S_AXIS_DIN_TDATA[143]; // rv 0
  assign S_AXIS_DIN_TDATA_in[144] = (S_AXIS_DIN_TDATA[144] !== 1'bz) && S_AXIS_DIN_TDATA[144]; // rv 0
  assign S_AXIS_DIN_TDATA_in[145] = (S_AXIS_DIN_TDATA[145] !== 1'bz) && S_AXIS_DIN_TDATA[145]; // rv 0
  assign S_AXIS_DIN_TDATA_in[146] = (S_AXIS_DIN_TDATA[146] !== 1'bz) && S_AXIS_DIN_TDATA[146]; // rv 0
  assign S_AXIS_DIN_TDATA_in[147] = (S_AXIS_DIN_TDATA[147] !== 1'bz) && S_AXIS_DIN_TDATA[147]; // rv 0
  assign S_AXIS_DIN_TDATA_in[148] = (S_AXIS_DIN_TDATA[148] !== 1'bz) && S_AXIS_DIN_TDATA[148]; // rv 0
  assign S_AXIS_DIN_TDATA_in[149] = (S_AXIS_DIN_TDATA[149] !== 1'bz) && S_AXIS_DIN_TDATA[149]; // rv 0
  assign S_AXIS_DIN_TDATA_in[14] = (S_AXIS_DIN_TDATA[14] !== 1'bz) && S_AXIS_DIN_TDATA[14]; // rv 0
  assign S_AXIS_DIN_TDATA_in[150] = (S_AXIS_DIN_TDATA[150] !== 1'bz) && S_AXIS_DIN_TDATA[150]; // rv 0
  assign S_AXIS_DIN_TDATA_in[151] = (S_AXIS_DIN_TDATA[151] !== 1'bz) && S_AXIS_DIN_TDATA[151]; // rv 0
  assign S_AXIS_DIN_TDATA_in[152] = (S_AXIS_DIN_TDATA[152] !== 1'bz) && S_AXIS_DIN_TDATA[152]; // rv 0
  assign S_AXIS_DIN_TDATA_in[153] = (S_AXIS_DIN_TDATA[153] !== 1'bz) && S_AXIS_DIN_TDATA[153]; // rv 0
  assign S_AXIS_DIN_TDATA_in[154] = (S_AXIS_DIN_TDATA[154] !== 1'bz) && S_AXIS_DIN_TDATA[154]; // rv 0
  assign S_AXIS_DIN_TDATA_in[155] = (S_AXIS_DIN_TDATA[155] !== 1'bz) && S_AXIS_DIN_TDATA[155]; // rv 0
  assign S_AXIS_DIN_TDATA_in[156] = (S_AXIS_DIN_TDATA[156] !== 1'bz) && S_AXIS_DIN_TDATA[156]; // rv 0
  assign S_AXIS_DIN_TDATA_in[157] = (S_AXIS_DIN_TDATA[157] !== 1'bz) && S_AXIS_DIN_TDATA[157]; // rv 0
  assign S_AXIS_DIN_TDATA_in[158] = (S_AXIS_DIN_TDATA[158] !== 1'bz) && S_AXIS_DIN_TDATA[158]; // rv 0
  assign S_AXIS_DIN_TDATA_in[159] = (S_AXIS_DIN_TDATA[159] !== 1'bz) && S_AXIS_DIN_TDATA[159]; // rv 0
  assign S_AXIS_DIN_TDATA_in[15] = (S_AXIS_DIN_TDATA[15] !== 1'bz) && S_AXIS_DIN_TDATA[15]; // rv 0
  assign S_AXIS_DIN_TDATA_in[160] = (S_AXIS_DIN_TDATA[160] !== 1'bz) && S_AXIS_DIN_TDATA[160]; // rv 0
  assign S_AXIS_DIN_TDATA_in[161] = (S_AXIS_DIN_TDATA[161] !== 1'bz) && S_AXIS_DIN_TDATA[161]; // rv 0
  assign S_AXIS_DIN_TDATA_in[162] = (S_AXIS_DIN_TDATA[162] !== 1'bz) && S_AXIS_DIN_TDATA[162]; // rv 0
  assign S_AXIS_DIN_TDATA_in[163] = (S_AXIS_DIN_TDATA[163] !== 1'bz) && S_AXIS_DIN_TDATA[163]; // rv 0
  assign S_AXIS_DIN_TDATA_in[164] = (S_AXIS_DIN_TDATA[164] !== 1'bz) && S_AXIS_DIN_TDATA[164]; // rv 0
  assign S_AXIS_DIN_TDATA_in[165] = (S_AXIS_DIN_TDATA[165] !== 1'bz) && S_AXIS_DIN_TDATA[165]; // rv 0
  assign S_AXIS_DIN_TDATA_in[166] = (S_AXIS_DIN_TDATA[166] !== 1'bz) && S_AXIS_DIN_TDATA[166]; // rv 0
  assign S_AXIS_DIN_TDATA_in[167] = (S_AXIS_DIN_TDATA[167] !== 1'bz) && S_AXIS_DIN_TDATA[167]; // rv 0
  assign S_AXIS_DIN_TDATA_in[168] = (S_AXIS_DIN_TDATA[168] !== 1'bz) && S_AXIS_DIN_TDATA[168]; // rv 0
  assign S_AXIS_DIN_TDATA_in[169] = (S_AXIS_DIN_TDATA[169] !== 1'bz) && S_AXIS_DIN_TDATA[169]; // rv 0
  assign S_AXIS_DIN_TDATA_in[16] = (S_AXIS_DIN_TDATA[16] !== 1'bz) && S_AXIS_DIN_TDATA[16]; // rv 0
  assign S_AXIS_DIN_TDATA_in[170] = (S_AXIS_DIN_TDATA[170] !== 1'bz) && S_AXIS_DIN_TDATA[170]; // rv 0
  assign S_AXIS_DIN_TDATA_in[171] = (S_AXIS_DIN_TDATA[171] !== 1'bz) && S_AXIS_DIN_TDATA[171]; // rv 0
  assign S_AXIS_DIN_TDATA_in[172] = (S_AXIS_DIN_TDATA[172] !== 1'bz) && S_AXIS_DIN_TDATA[172]; // rv 0
  assign S_AXIS_DIN_TDATA_in[173] = (S_AXIS_DIN_TDATA[173] !== 1'bz) && S_AXIS_DIN_TDATA[173]; // rv 0
  assign S_AXIS_DIN_TDATA_in[174] = (S_AXIS_DIN_TDATA[174] !== 1'bz) && S_AXIS_DIN_TDATA[174]; // rv 0
  assign S_AXIS_DIN_TDATA_in[175] = (S_AXIS_DIN_TDATA[175] !== 1'bz) && S_AXIS_DIN_TDATA[175]; // rv 0
  assign S_AXIS_DIN_TDATA_in[176] = (S_AXIS_DIN_TDATA[176] !== 1'bz) && S_AXIS_DIN_TDATA[176]; // rv 0
  assign S_AXIS_DIN_TDATA_in[177] = (S_AXIS_DIN_TDATA[177] !== 1'bz) && S_AXIS_DIN_TDATA[177]; // rv 0
  assign S_AXIS_DIN_TDATA_in[178] = (S_AXIS_DIN_TDATA[178] !== 1'bz) && S_AXIS_DIN_TDATA[178]; // rv 0
  assign S_AXIS_DIN_TDATA_in[179] = (S_AXIS_DIN_TDATA[179] !== 1'bz) && S_AXIS_DIN_TDATA[179]; // rv 0
  assign S_AXIS_DIN_TDATA_in[17] = (S_AXIS_DIN_TDATA[17] !== 1'bz) && S_AXIS_DIN_TDATA[17]; // rv 0
  assign S_AXIS_DIN_TDATA_in[180] = (S_AXIS_DIN_TDATA[180] !== 1'bz) && S_AXIS_DIN_TDATA[180]; // rv 0
  assign S_AXIS_DIN_TDATA_in[181] = (S_AXIS_DIN_TDATA[181] !== 1'bz) && S_AXIS_DIN_TDATA[181]; // rv 0
  assign S_AXIS_DIN_TDATA_in[182] = (S_AXIS_DIN_TDATA[182] !== 1'bz) && S_AXIS_DIN_TDATA[182]; // rv 0
  assign S_AXIS_DIN_TDATA_in[183] = (S_AXIS_DIN_TDATA[183] !== 1'bz) && S_AXIS_DIN_TDATA[183]; // rv 0
  assign S_AXIS_DIN_TDATA_in[184] = (S_AXIS_DIN_TDATA[184] !== 1'bz) && S_AXIS_DIN_TDATA[184]; // rv 0
  assign S_AXIS_DIN_TDATA_in[185] = (S_AXIS_DIN_TDATA[185] !== 1'bz) && S_AXIS_DIN_TDATA[185]; // rv 0
  assign S_AXIS_DIN_TDATA_in[186] = (S_AXIS_DIN_TDATA[186] !== 1'bz) && S_AXIS_DIN_TDATA[186]; // rv 0
  assign S_AXIS_DIN_TDATA_in[187] = (S_AXIS_DIN_TDATA[187] !== 1'bz) && S_AXIS_DIN_TDATA[187]; // rv 0
  assign S_AXIS_DIN_TDATA_in[188] = (S_AXIS_DIN_TDATA[188] !== 1'bz) && S_AXIS_DIN_TDATA[188]; // rv 0
  assign S_AXIS_DIN_TDATA_in[189] = (S_AXIS_DIN_TDATA[189] !== 1'bz) && S_AXIS_DIN_TDATA[189]; // rv 0
  assign S_AXIS_DIN_TDATA_in[18] = (S_AXIS_DIN_TDATA[18] !== 1'bz) && S_AXIS_DIN_TDATA[18]; // rv 0
  assign S_AXIS_DIN_TDATA_in[190] = (S_AXIS_DIN_TDATA[190] !== 1'bz) && S_AXIS_DIN_TDATA[190]; // rv 0
  assign S_AXIS_DIN_TDATA_in[191] = (S_AXIS_DIN_TDATA[191] !== 1'bz) && S_AXIS_DIN_TDATA[191]; // rv 0
  assign S_AXIS_DIN_TDATA_in[192] = (S_AXIS_DIN_TDATA[192] !== 1'bz) && S_AXIS_DIN_TDATA[192]; // rv 0
  assign S_AXIS_DIN_TDATA_in[193] = (S_AXIS_DIN_TDATA[193] !== 1'bz) && S_AXIS_DIN_TDATA[193]; // rv 0
  assign S_AXIS_DIN_TDATA_in[194] = (S_AXIS_DIN_TDATA[194] !== 1'bz) && S_AXIS_DIN_TDATA[194]; // rv 0
  assign S_AXIS_DIN_TDATA_in[195] = (S_AXIS_DIN_TDATA[195] !== 1'bz) && S_AXIS_DIN_TDATA[195]; // rv 0
  assign S_AXIS_DIN_TDATA_in[196] = (S_AXIS_DIN_TDATA[196] !== 1'bz) && S_AXIS_DIN_TDATA[196]; // rv 0
  assign S_AXIS_DIN_TDATA_in[197] = (S_AXIS_DIN_TDATA[197] !== 1'bz) && S_AXIS_DIN_TDATA[197]; // rv 0
  assign S_AXIS_DIN_TDATA_in[198] = (S_AXIS_DIN_TDATA[198] !== 1'bz) && S_AXIS_DIN_TDATA[198]; // rv 0
  assign S_AXIS_DIN_TDATA_in[199] = (S_AXIS_DIN_TDATA[199] !== 1'bz) && S_AXIS_DIN_TDATA[199]; // rv 0
  assign S_AXIS_DIN_TDATA_in[19] = (S_AXIS_DIN_TDATA[19] !== 1'bz) && S_AXIS_DIN_TDATA[19]; // rv 0
  assign S_AXIS_DIN_TDATA_in[1] = (S_AXIS_DIN_TDATA[1] !== 1'bz) && S_AXIS_DIN_TDATA[1]; // rv 0
  assign S_AXIS_DIN_TDATA_in[200] = (S_AXIS_DIN_TDATA[200] !== 1'bz) && S_AXIS_DIN_TDATA[200]; // rv 0
  assign S_AXIS_DIN_TDATA_in[201] = (S_AXIS_DIN_TDATA[201] !== 1'bz) && S_AXIS_DIN_TDATA[201]; // rv 0
  assign S_AXIS_DIN_TDATA_in[202] = (S_AXIS_DIN_TDATA[202] !== 1'bz) && S_AXIS_DIN_TDATA[202]; // rv 0
  assign S_AXIS_DIN_TDATA_in[203] = (S_AXIS_DIN_TDATA[203] !== 1'bz) && S_AXIS_DIN_TDATA[203]; // rv 0
  assign S_AXIS_DIN_TDATA_in[204] = (S_AXIS_DIN_TDATA[204] !== 1'bz) && S_AXIS_DIN_TDATA[204]; // rv 0
  assign S_AXIS_DIN_TDATA_in[205] = (S_AXIS_DIN_TDATA[205] !== 1'bz) && S_AXIS_DIN_TDATA[205]; // rv 0
  assign S_AXIS_DIN_TDATA_in[206] = (S_AXIS_DIN_TDATA[206] !== 1'bz) && S_AXIS_DIN_TDATA[206]; // rv 0
  assign S_AXIS_DIN_TDATA_in[207] = (S_AXIS_DIN_TDATA[207] !== 1'bz) && S_AXIS_DIN_TDATA[207]; // rv 0
  assign S_AXIS_DIN_TDATA_in[208] = (S_AXIS_DIN_TDATA[208] !== 1'bz) && S_AXIS_DIN_TDATA[208]; // rv 0
  assign S_AXIS_DIN_TDATA_in[209] = (S_AXIS_DIN_TDATA[209] !== 1'bz) && S_AXIS_DIN_TDATA[209]; // rv 0
  assign S_AXIS_DIN_TDATA_in[20] = (S_AXIS_DIN_TDATA[20] !== 1'bz) && S_AXIS_DIN_TDATA[20]; // rv 0
  assign S_AXIS_DIN_TDATA_in[210] = (S_AXIS_DIN_TDATA[210] !== 1'bz) && S_AXIS_DIN_TDATA[210]; // rv 0
  assign S_AXIS_DIN_TDATA_in[211] = (S_AXIS_DIN_TDATA[211] !== 1'bz) && S_AXIS_DIN_TDATA[211]; // rv 0
  assign S_AXIS_DIN_TDATA_in[212] = (S_AXIS_DIN_TDATA[212] !== 1'bz) && S_AXIS_DIN_TDATA[212]; // rv 0
  assign S_AXIS_DIN_TDATA_in[213] = (S_AXIS_DIN_TDATA[213] !== 1'bz) && S_AXIS_DIN_TDATA[213]; // rv 0
  assign S_AXIS_DIN_TDATA_in[214] = (S_AXIS_DIN_TDATA[214] !== 1'bz) && S_AXIS_DIN_TDATA[214]; // rv 0
  assign S_AXIS_DIN_TDATA_in[215] = (S_AXIS_DIN_TDATA[215] !== 1'bz) && S_AXIS_DIN_TDATA[215]; // rv 0
  assign S_AXIS_DIN_TDATA_in[216] = (S_AXIS_DIN_TDATA[216] !== 1'bz) && S_AXIS_DIN_TDATA[216]; // rv 0
  assign S_AXIS_DIN_TDATA_in[217] = (S_AXIS_DIN_TDATA[217] !== 1'bz) && S_AXIS_DIN_TDATA[217]; // rv 0
  assign S_AXIS_DIN_TDATA_in[218] = (S_AXIS_DIN_TDATA[218] !== 1'bz) && S_AXIS_DIN_TDATA[218]; // rv 0
  assign S_AXIS_DIN_TDATA_in[219] = (S_AXIS_DIN_TDATA[219] !== 1'bz) && S_AXIS_DIN_TDATA[219]; // rv 0
  assign S_AXIS_DIN_TDATA_in[21] = (S_AXIS_DIN_TDATA[21] !== 1'bz) && S_AXIS_DIN_TDATA[21]; // rv 0
  assign S_AXIS_DIN_TDATA_in[220] = (S_AXIS_DIN_TDATA[220] !== 1'bz) && S_AXIS_DIN_TDATA[220]; // rv 0
  assign S_AXIS_DIN_TDATA_in[221] = (S_AXIS_DIN_TDATA[221] !== 1'bz) && S_AXIS_DIN_TDATA[221]; // rv 0
  assign S_AXIS_DIN_TDATA_in[222] = (S_AXIS_DIN_TDATA[222] !== 1'bz) && S_AXIS_DIN_TDATA[222]; // rv 0
  assign S_AXIS_DIN_TDATA_in[223] = (S_AXIS_DIN_TDATA[223] !== 1'bz) && S_AXIS_DIN_TDATA[223]; // rv 0
  assign S_AXIS_DIN_TDATA_in[224] = (S_AXIS_DIN_TDATA[224] !== 1'bz) && S_AXIS_DIN_TDATA[224]; // rv 0
  assign S_AXIS_DIN_TDATA_in[225] = (S_AXIS_DIN_TDATA[225] !== 1'bz) && S_AXIS_DIN_TDATA[225]; // rv 0
  assign S_AXIS_DIN_TDATA_in[226] = (S_AXIS_DIN_TDATA[226] !== 1'bz) && S_AXIS_DIN_TDATA[226]; // rv 0
  assign S_AXIS_DIN_TDATA_in[227] = (S_AXIS_DIN_TDATA[227] !== 1'bz) && S_AXIS_DIN_TDATA[227]; // rv 0
  assign S_AXIS_DIN_TDATA_in[228] = (S_AXIS_DIN_TDATA[228] !== 1'bz) && S_AXIS_DIN_TDATA[228]; // rv 0
  assign S_AXIS_DIN_TDATA_in[229] = (S_AXIS_DIN_TDATA[229] !== 1'bz) && S_AXIS_DIN_TDATA[229]; // rv 0
  assign S_AXIS_DIN_TDATA_in[22] = (S_AXIS_DIN_TDATA[22] !== 1'bz) && S_AXIS_DIN_TDATA[22]; // rv 0
  assign S_AXIS_DIN_TDATA_in[230] = (S_AXIS_DIN_TDATA[230] !== 1'bz) && S_AXIS_DIN_TDATA[230]; // rv 0
  assign S_AXIS_DIN_TDATA_in[231] = (S_AXIS_DIN_TDATA[231] !== 1'bz) && S_AXIS_DIN_TDATA[231]; // rv 0
  assign S_AXIS_DIN_TDATA_in[232] = (S_AXIS_DIN_TDATA[232] !== 1'bz) && S_AXIS_DIN_TDATA[232]; // rv 0
  assign S_AXIS_DIN_TDATA_in[233] = (S_AXIS_DIN_TDATA[233] !== 1'bz) && S_AXIS_DIN_TDATA[233]; // rv 0
  assign S_AXIS_DIN_TDATA_in[234] = (S_AXIS_DIN_TDATA[234] !== 1'bz) && S_AXIS_DIN_TDATA[234]; // rv 0
  assign S_AXIS_DIN_TDATA_in[235] = (S_AXIS_DIN_TDATA[235] !== 1'bz) && S_AXIS_DIN_TDATA[235]; // rv 0
  assign S_AXIS_DIN_TDATA_in[236] = (S_AXIS_DIN_TDATA[236] !== 1'bz) && S_AXIS_DIN_TDATA[236]; // rv 0
  assign S_AXIS_DIN_TDATA_in[237] = (S_AXIS_DIN_TDATA[237] !== 1'bz) && S_AXIS_DIN_TDATA[237]; // rv 0
  assign S_AXIS_DIN_TDATA_in[238] = (S_AXIS_DIN_TDATA[238] !== 1'bz) && S_AXIS_DIN_TDATA[238]; // rv 0
  assign S_AXIS_DIN_TDATA_in[239] = (S_AXIS_DIN_TDATA[239] !== 1'bz) && S_AXIS_DIN_TDATA[239]; // rv 0
  assign S_AXIS_DIN_TDATA_in[23] = (S_AXIS_DIN_TDATA[23] !== 1'bz) && S_AXIS_DIN_TDATA[23]; // rv 0
  assign S_AXIS_DIN_TDATA_in[240] = (S_AXIS_DIN_TDATA[240] !== 1'bz) && S_AXIS_DIN_TDATA[240]; // rv 0
  assign S_AXIS_DIN_TDATA_in[241] = (S_AXIS_DIN_TDATA[241] !== 1'bz) && S_AXIS_DIN_TDATA[241]; // rv 0
  assign S_AXIS_DIN_TDATA_in[242] = (S_AXIS_DIN_TDATA[242] !== 1'bz) && S_AXIS_DIN_TDATA[242]; // rv 0
  assign S_AXIS_DIN_TDATA_in[243] = (S_AXIS_DIN_TDATA[243] !== 1'bz) && S_AXIS_DIN_TDATA[243]; // rv 0
  assign S_AXIS_DIN_TDATA_in[244] = (S_AXIS_DIN_TDATA[244] !== 1'bz) && S_AXIS_DIN_TDATA[244]; // rv 0
  assign S_AXIS_DIN_TDATA_in[245] = (S_AXIS_DIN_TDATA[245] !== 1'bz) && S_AXIS_DIN_TDATA[245]; // rv 0
  assign S_AXIS_DIN_TDATA_in[246] = (S_AXIS_DIN_TDATA[246] !== 1'bz) && S_AXIS_DIN_TDATA[246]; // rv 0
  assign S_AXIS_DIN_TDATA_in[247] = (S_AXIS_DIN_TDATA[247] !== 1'bz) && S_AXIS_DIN_TDATA[247]; // rv 0
  assign S_AXIS_DIN_TDATA_in[248] = (S_AXIS_DIN_TDATA[248] !== 1'bz) && S_AXIS_DIN_TDATA[248]; // rv 0
  assign S_AXIS_DIN_TDATA_in[249] = (S_AXIS_DIN_TDATA[249] !== 1'bz) && S_AXIS_DIN_TDATA[249]; // rv 0
  assign S_AXIS_DIN_TDATA_in[24] = (S_AXIS_DIN_TDATA[24] !== 1'bz) && S_AXIS_DIN_TDATA[24]; // rv 0
  assign S_AXIS_DIN_TDATA_in[250] = (S_AXIS_DIN_TDATA[250] !== 1'bz) && S_AXIS_DIN_TDATA[250]; // rv 0
  assign S_AXIS_DIN_TDATA_in[251] = (S_AXIS_DIN_TDATA[251] !== 1'bz) && S_AXIS_DIN_TDATA[251]; // rv 0
  assign S_AXIS_DIN_TDATA_in[252] = (S_AXIS_DIN_TDATA[252] !== 1'bz) && S_AXIS_DIN_TDATA[252]; // rv 0
  assign S_AXIS_DIN_TDATA_in[253] = (S_AXIS_DIN_TDATA[253] !== 1'bz) && S_AXIS_DIN_TDATA[253]; // rv 0
  assign S_AXIS_DIN_TDATA_in[254] = (S_AXIS_DIN_TDATA[254] !== 1'bz) && S_AXIS_DIN_TDATA[254]; // rv 0
  assign S_AXIS_DIN_TDATA_in[255] = (S_AXIS_DIN_TDATA[255] !== 1'bz) && S_AXIS_DIN_TDATA[255]; // rv 0
  assign S_AXIS_DIN_TDATA_in[256] = (S_AXIS_DIN_TDATA[256] !== 1'bz) && S_AXIS_DIN_TDATA[256]; // rv 0
  assign S_AXIS_DIN_TDATA_in[257] = (S_AXIS_DIN_TDATA[257] !== 1'bz) && S_AXIS_DIN_TDATA[257]; // rv 0
  assign S_AXIS_DIN_TDATA_in[258] = (S_AXIS_DIN_TDATA[258] !== 1'bz) && S_AXIS_DIN_TDATA[258]; // rv 0
  assign S_AXIS_DIN_TDATA_in[259] = (S_AXIS_DIN_TDATA[259] !== 1'bz) && S_AXIS_DIN_TDATA[259]; // rv 0
  assign S_AXIS_DIN_TDATA_in[25] = (S_AXIS_DIN_TDATA[25] !== 1'bz) && S_AXIS_DIN_TDATA[25]; // rv 0
  assign S_AXIS_DIN_TDATA_in[260] = (S_AXIS_DIN_TDATA[260] !== 1'bz) && S_AXIS_DIN_TDATA[260]; // rv 0
  assign S_AXIS_DIN_TDATA_in[261] = (S_AXIS_DIN_TDATA[261] !== 1'bz) && S_AXIS_DIN_TDATA[261]; // rv 0
  assign S_AXIS_DIN_TDATA_in[262] = (S_AXIS_DIN_TDATA[262] !== 1'bz) && S_AXIS_DIN_TDATA[262]; // rv 0
  assign S_AXIS_DIN_TDATA_in[263] = (S_AXIS_DIN_TDATA[263] !== 1'bz) && S_AXIS_DIN_TDATA[263]; // rv 0
  assign S_AXIS_DIN_TDATA_in[264] = (S_AXIS_DIN_TDATA[264] !== 1'bz) && S_AXIS_DIN_TDATA[264]; // rv 0
  assign S_AXIS_DIN_TDATA_in[265] = (S_AXIS_DIN_TDATA[265] !== 1'bz) && S_AXIS_DIN_TDATA[265]; // rv 0
  assign S_AXIS_DIN_TDATA_in[266] = (S_AXIS_DIN_TDATA[266] !== 1'bz) && S_AXIS_DIN_TDATA[266]; // rv 0
  assign S_AXIS_DIN_TDATA_in[267] = (S_AXIS_DIN_TDATA[267] !== 1'bz) && S_AXIS_DIN_TDATA[267]; // rv 0
  assign S_AXIS_DIN_TDATA_in[268] = (S_AXIS_DIN_TDATA[268] !== 1'bz) && S_AXIS_DIN_TDATA[268]; // rv 0
  assign S_AXIS_DIN_TDATA_in[269] = (S_AXIS_DIN_TDATA[269] !== 1'bz) && S_AXIS_DIN_TDATA[269]; // rv 0
  assign S_AXIS_DIN_TDATA_in[26] = (S_AXIS_DIN_TDATA[26] !== 1'bz) && S_AXIS_DIN_TDATA[26]; // rv 0
  assign S_AXIS_DIN_TDATA_in[270] = (S_AXIS_DIN_TDATA[270] !== 1'bz) && S_AXIS_DIN_TDATA[270]; // rv 0
  assign S_AXIS_DIN_TDATA_in[271] = (S_AXIS_DIN_TDATA[271] !== 1'bz) && S_AXIS_DIN_TDATA[271]; // rv 0
  assign S_AXIS_DIN_TDATA_in[272] = (S_AXIS_DIN_TDATA[272] !== 1'bz) && S_AXIS_DIN_TDATA[272]; // rv 0
  assign S_AXIS_DIN_TDATA_in[273] = (S_AXIS_DIN_TDATA[273] !== 1'bz) && S_AXIS_DIN_TDATA[273]; // rv 0
  assign S_AXIS_DIN_TDATA_in[274] = (S_AXIS_DIN_TDATA[274] !== 1'bz) && S_AXIS_DIN_TDATA[274]; // rv 0
  assign S_AXIS_DIN_TDATA_in[275] = (S_AXIS_DIN_TDATA[275] !== 1'bz) && S_AXIS_DIN_TDATA[275]; // rv 0
  assign S_AXIS_DIN_TDATA_in[276] = (S_AXIS_DIN_TDATA[276] !== 1'bz) && S_AXIS_DIN_TDATA[276]; // rv 0
  assign S_AXIS_DIN_TDATA_in[277] = (S_AXIS_DIN_TDATA[277] !== 1'bz) && S_AXIS_DIN_TDATA[277]; // rv 0
  assign S_AXIS_DIN_TDATA_in[278] = (S_AXIS_DIN_TDATA[278] !== 1'bz) && S_AXIS_DIN_TDATA[278]; // rv 0
  assign S_AXIS_DIN_TDATA_in[279] = (S_AXIS_DIN_TDATA[279] !== 1'bz) && S_AXIS_DIN_TDATA[279]; // rv 0
  assign S_AXIS_DIN_TDATA_in[27] = (S_AXIS_DIN_TDATA[27] !== 1'bz) && S_AXIS_DIN_TDATA[27]; // rv 0
  assign S_AXIS_DIN_TDATA_in[280] = (S_AXIS_DIN_TDATA[280] !== 1'bz) && S_AXIS_DIN_TDATA[280]; // rv 0
  assign S_AXIS_DIN_TDATA_in[281] = (S_AXIS_DIN_TDATA[281] !== 1'bz) && S_AXIS_DIN_TDATA[281]; // rv 0
  assign S_AXIS_DIN_TDATA_in[282] = (S_AXIS_DIN_TDATA[282] !== 1'bz) && S_AXIS_DIN_TDATA[282]; // rv 0
  assign S_AXIS_DIN_TDATA_in[283] = (S_AXIS_DIN_TDATA[283] !== 1'bz) && S_AXIS_DIN_TDATA[283]; // rv 0
  assign S_AXIS_DIN_TDATA_in[284] = (S_AXIS_DIN_TDATA[284] !== 1'bz) && S_AXIS_DIN_TDATA[284]; // rv 0
  assign S_AXIS_DIN_TDATA_in[285] = (S_AXIS_DIN_TDATA[285] !== 1'bz) && S_AXIS_DIN_TDATA[285]; // rv 0
  assign S_AXIS_DIN_TDATA_in[286] = (S_AXIS_DIN_TDATA[286] !== 1'bz) && S_AXIS_DIN_TDATA[286]; // rv 0
  assign S_AXIS_DIN_TDATA_in[287] = (S_AXIS_DIN_TDATA[287] !== 1'bz) && S_AXIS_DIN_TDATA[287]; // rv 0
  assign S_AXIS_DIN_TDATA_in[288] = (S_AXIS_DIN_TDATA[288] !== 1'bz) && S_AXIS_DIN_TDATA[288]; // rv 0
  assign S_AXIS_DIN_TDATA_in[289] = (S_AXIS_DIN_TDATA[289] !== 1'bz) && S_AXIS_DIN_TDATA[289]; // rv 0
  assign S_AXIS_DIN_TDATA_in[28] = (S_AXIS_DIN_TDATA[28] !== 1'bz) && S_AXIS_DIN_TDATA[28]; // rv 0
  assign S_AXIS_DIN_TDATA_in[290] = (S_AXIS_DIN_TDATA[290] !== 1'bz) && S_AXIS_DIN_TDATA[290]; // rv 0
  assign S_AXIS_DIN_TDATA_in[291] = (S_AXIS_DIN_TDATA[291] !== 1'bz) && S_AXIS_DIN_TDATA[291]; // rv 0
  assign S_AXIS_DIN_TDATA_in[292] = (S_AXIS_DIN_TDATA[292] !== 1'bz) && S_AXIS_DIN_TDATA[292]; // rv 0
  assign S_AXIS_DIN_TDATA_in[293] = (S_AXIS_DIN_TDATA[293] !== 1'bz) && S_AXIS_DIN_TDATA[293]; // rv 0
  assign S_AXIS_DIN_TDATA_in[294] = (S_AXIS_DIN_TDATA[294] !== 1'bz) && S_AXIS_DIN_TDATA[294]; // rv 0
  assign S_AXIS_DIN_TDATA_in[295] = (S_AXIS_DIN_TDATA[295] !== 1'bz) && S_AXIS_DIN_TDATA[295]; // rv 0
  assign S_AXIS_DIN_TDATA_in[296] = (S_AXIS_DIN_TDATA[296] !== 1'bz) && S_AXIS_DIN_TDATA[296]; // rv 0
  assign S_AXIS_DIN_TDATA_in[297] = (S_AXIS_DIN_TDATA[297] !== 1'bz) && S_AXIS_DIN_TDATA[297]; // rv 0
  assign S_AXIS_DIN_TDATA_in[298] = (S_AXIS_DIN_TDATA[298] !== 1'bz) && S_AXIS_DIN_TDATA[298]; // rv 0
  assign S_AXIS_DIN_TDATA_in[299] = (S_AXIS_DIN_TDATA[299] !== 1'bz) && S_AXIS_DIN_TDATA[299]; // rv 0
  assign S_AXIS_DIN_TDATA_in[29] = (S_AXIS_DIN_TDATA[29] !== 1'bz) && S_AXIS_DIN_TDATA[29]; // rv 0
  assign S_AXIS_DIN_TDATA_in[2] = (S_AXIS_DIN_TDATA[2] !== 1'bz) && S_AXIS_DIN_TDATA[2]; // rv 0
  assign S_AXIS_DIN_TDATA_in[300] = (S_AXIS_DIN_TDATA[300] !== 1'bz) && S_AXIS_DIN_TDATA[300]; // rv 0
  assign S_AXIS_DIN_TDATA_in[301] = (S_AXIS_DIN_TDATA[301] !== 1'bz) && S_AXIS_DIN_TDATA[301]; // rv 0
  assign S_AXIS_DIN_TDATA_in[302] = (S_AXIS_DIN_TDATA[302] !== 1'bz) && S_AXIS_DIN_TDATA[302]; // rv 0
  assign S_AXIS_DIN_TDATA_in[303] = (S_AXIS_DIN_TDATA[303] !== 1'bz) && S_AXIS_DIN_TDATA[303]; // rv 0
  assign S_AXIS_DIN_TDATA_in[304] = (S_AXIS_DIN_TDATA[304] !== 1'bz) && S_AXIS_DIN_TDATA[304]; // rv 0
  assign S_AXIS_DIN_TDATA_in[305] = (S_AXIS_DIN_TDATA[305] !== 1'bz) && S_AXIS_DIN_TDATA[305]; // rv 0
  assign S_AXIS_DIN_TDATA_in[306] = (S_AXIS_DIN_TDATA[306] !== 1'bz) && S_AXIS_DIN_TDATA[306]; // rv 0
  assign S_AXIS_DIN_TDATA_in[307] = (S_AXIS_DIN_TDATA[307] !== 1'bz) && S_AXIS_DIN_TDATA[307]; // rv 0
  assign S_AXIS_DIN_TDATA_in[308] = (S_AXIS_DIN_TDATA[308] !== 1'bz) && S_AXIS_DIN_TDATA[308]; // rv 0
  assign S_AXIS_DIN_TDATA_in[309] = (S_AXIS_DIN_TDATA[309] !== 1'bz) && S_AXIS_DIN_TDATA[309]; // rv 0
  assign S_AXIS_DIN_TDATA_in[30] = (S_AXIS_DIN_TDATA[30] !== 1'bz) && S_AXIS_DIN_TDATA[30]; // rv 0
  assign S_AXIS_DIN_TDATA_in[310] = (S_AXIS_DIN_TDATA[310] !== 1'bz) && S_AXIS_DIN_TDATA[310]; // rv 0
  assign S_AXIS_DIN_TDATA_in[311] = (S_AXIS_DIN_TDATA[311] !== 1'bz) && S_AXIS_DIN_TDATA[311]; // rv 0
  assign S_AXIS_DIN_TDATA_in[312] = (S_AXIS_DIN_TDATA[312] !== 1'bz) && S_AXIS_DIN_TDATA[312]; // rv 0
  assign S_AXIS_DIN_TDATA_in[313] = (S_AXIS_DIN_TDATA[313] !== 1'bz) && S_AXIS_DIN_TDATA[313]; // rv 0
  assign S_AXIS_DIN_TDATA_in[314] = (S_AXIS_DIN_TDATA[314] !== 1'bz) && S_AXIS_DIN_TDATA[314]; // rv 0
  assign S_AXIS_DIN_TDATA_in[315] = (S_AXIS_DIN_TDATA[315] !== 1'bz) && S_AXIS_DIN_TDATA[315]; // rv 0
  assign S_AXIS_DIN_TDATA_in[316] = (S_AXIS_DIN_TDATA[316] !== 1'bz) && S_AXIS_DIN_TDATA[316]; // rv 0
  assign S_AXIS_DIN_TDATA_in[317] = (S_AXIS_DIN_TDATA[317] !== 1'bz) && S_AXIS_DIN_TDATA[317]; // rv 0
  assign S_AXIS_DIN_TDATA_in[318] = (S_AXIS_DIN_TDATA[318] !== 1'bz) && S_AXIS_DIN_TDATA[318]; // rv 0
  assign S_AXIS_DIN_TDATA_in[319] = (S_AXIS_DIN_TDATA[319] !== 1'bz) && S_AXIS_DIN_TDATA[319]; // rv 0
  assign S_AXIS_DIN_TDATA_in[31] = (S_AXIS_DIN_TDATA[31] !== 1'bz) && S_AXIS_DIN_TDATA[31]; // rv 0
  assign S_AXIS_DIN_TDATA_in[320] = (S_AXIS_DIN_TDATA[320] !== 1'bz) && S_AXIS_DIN_TDATA[320]; // rv 0
  assign S_AXIS_DIN_TDATA_in[321] = (S_AXIS_DIN_TDATA[321] !== 1'bz) && S_AXIS_DIN_TDATA[321]; // rv 0
  assign S_AXIS_DIN_TDATA_in[322] = (S_AXIS_DIN_TDATA[322] !== 1'bz) && S_AXIS_DIN_TDATA[322]; // rv 0
  assign S_AXIS_DIN_TDATA_in[323] = (S_AXIS_DIN_TDATA[323] !== 1'bz) && S_AXIS_DIN_TDATA[323]; // rv 0
  assign S_AXIS_DIN_TDATA_in[324] = (S_AXIS_DIN_TDATA[324] !== 1'bz) && S_AXIS_DIN_TDATA[324]; // rv 0
  assign S_AXIS_DIN_TDATA_in[325] = (S_AXIS_DIN_TDATA[325] !== 1'bz) && S_AXIS_DIN_TDATA[325]; // rv 0
  assign S_AXIS_DIN_TDATA_in[326] = (S_AXIS_DIN_TDATA[326] !== 1'bz) && S_AXIS_DIN_TDATA[326]; // rv 0
  assign S_AXIS_DIN_TDATA_in[327] = (S_AXIS_DIN_TDATA[327] !== 1'bz) && S_AXIS_DIN_TDATA[327]; // rv 0
  assign S_AXIS_DIN_TDATA_in[328] = (S_AXIS_DIN_TDATA[328] !== 1'bz) && S_AXIS_DIN_TDATA[328]; // rv 0
  assign S_AXIS_DIN_TDATA_in[329] = (S_AXIS_DIN_TDATA[329] !== 1'bz) && S_AXIS_DIN_TDATA[329]; // rv 0
  assign S_AXIS_DIN_TDATA_in[32] = (S_AXIS_DIN_TDATA[32] !== 1'bz) && S_AXIS_DIN_TDATA[32]; // rv 0
  assign S_AXIS_DIN_TDATA_in[330] = (S_AXIS_DIN_TDATA[330] !== 1'bz) && S_AXIS_DIN_TDATA[330]; // rv 0
  assign S_AXIS_DIN_TDATA_in[331] = (S_AXIS_DIN_TDATA[331] !== 1'bz) && S_AXIS_DIN_TDATA[331]; // rv 0
  assign S_AXIS_DIN_TDATA_in[332] = (S_AXIS_DIN_TDATA[332] !== 1'bz) && S_AXIS_DIN_TDATA[332]; // rv 0
  assign S_AXIS_DIN_TDATA_in[333] = (S_AXIS_DIN_TDATA[333] !== 1'bz) && S_AXIS_DIN_TDATA[333]; // rv 0
  assign S_AXIS_DIN_TDATA_in[334] = (S_AXIS_DIN_TDATA[334] !== 1'bz) && S_AXIS_DIN_TDATA[334]; // rv 0
  assign S_AXIS_DIN_TDATA_in[335] = (S_AXIS_DIN_TDATA[335] !== 1'bz) && S_AXIS_DIN_TDATA[335]; // rv 0
  assign S_AXIS_DIN_TDATA_in[336] = (S_AXIS_DIN_TDATA[336] !== 1'bz) && S_AXIS_DIN_TDATA[336]; // rv 0
  assign S_AXIS_DIN_TDATA_in[337] = (S_AXIS_DIN_TDATA[337] !== 1'bz) && S_AXIS_DIN_TDATA[337]; // rv 0
  assign S_AXIS_DIN_TDATA_in[338] = (S_AXIS_DIN_TDATA[338] !== 1'bz) && S_AXIS_DIN_TDATA[338]; // rv 0
  assign S_AXIS_DIN_TDATA_in[339] = (S_AXIS_DIN_TDATA[339] !== 1'bz) && S_AXIS_DIN_TDATA[339]; // rv 0
  assign S_AXIS_DIN_TDATA_in[33] = (S_AXIS_DIN_TDATA[33] !== 1'bz) && S_AXIS_DIN_TDATA[33]; // rv 0
  assign S_AXIS_DIN_TDATA_in[340] = (S_AXIS_DIN_TDATA[340] !== 1'bz) && S_AXIS_DIN_TDATA[340]; // rv 0
  assign S_AXIS_DIN_TDATA_in[341] = (S_AXIS_DIN_TDATA[341] !== 1'bz) && S_AXIS_DIN_TDATA[341]; // rv 0
  assign S_AXIS_DIN_TDATA_in[342] = (S_AXIS_DIN_TDATA[342] !== 1'bz) && S_AXIS_DIN_TDATA[342]; // rv 0
  assign S_AXIS_DIN_TDATA_in[343] = (S_AXIS_DIN_TDATA[343] !== 1'bz) && S_AXIS_DIN_TDATA[343]; // rv 0
  assign S_AXIS_DIN_TDATA_in[344] = (S_AXIS_DIN_TDATA[344] !== 1'bz) && S_AXIS_DIN_TDATA[344]; // rv 0
  assign S_AXIS_DIN_TDATA_in[345] = (S_AXIS_DIN_TDATA[345] !== 1'bz) && S_AXIS_DIN_TDATA[345]; // rv 0
  assign S_AXIS_DIN_TDATA_in[346] = (S_AXIS_DIN_TDATA[346] !== 1'bz) && S_AXIS_DIN_TDATA[346]; // rv 0
  assign S_AXIS_DIN_TDATA_in[347] = (S_AXIS_DIN_TDATA[347] !== 1'bz) && S_AXIS_DIN_TDATA[347]; // rv 0
  assign S_AXIS_DIN_TDATA_in[348] = (S_AXIS_DIN_TDATA[348] !== 1'bz) && S_AXIS_DIN_TDATA[348]; // rv 0
  assign S_AXIS_DIN_TDATA_in[349] = (S_AXIS_DIN_TDATA[349] !== 1'bz) && S_AXIS_DIN_TDATA[349]; // rv 0
  assign S_AXIS_DIN_TDATA_in[34] = (S_AXIS_DIN_TDATA[34] !== 1'bz) && S_AXIS_DIN_TDATA[34]; // rv 0
  assign S_AXIS_DIN_TDATA_in[350] = (S_AXIS_DIN_TDATA[350] !== 1'bz) && S_AXIS_DIN_TDATA[350]; // rv 0
  assign S_AXIS_DIN_TDATA_in[351] = (S_AXIS_DIN_TDATA[351] !== 1'bz) && S_AXIS_DIN_TDATA[351]; // rv 0
  assign S_AXIS_DIN_TDATA_in[352] = (S_AXIS_DIN_TDATA[352] !== 1'bz) && S_AXIS_DIN_TDATA[352]; // rv 0
  assign S_AXIS_DIN_TDATA_in[353] = (S_AXIS_DIN_TDATA[353] !== 1'bz) && S_AXIS_DIN_TDATA[353]; // rv 0
  assign S_AXIS_DIN_TDATA_in[354] = (S_AXIS_DIN_TDATA[354] !== 1'bz) && S_AXIS_DIN_TDATA[354]; // rv 0
  assign S_AXIS_DIN_TDATA_in[355] = (S_AXIS_DIN_TDATA[355] !== 1'bz) && S_AXIS_DIN_TDATA[355]; // rv 0
  assign S_AXIS_DIN_TDATA_in[356] = (S_AXIS_DIN_TDATA[356] !== 1'bz) && S_AXIS_DIN_TDATA[356]; // rv 0
  assign S_AXIS_DIN_TDATA_in[357] = (S_AXIS_DIN_TDATA[357] !== 1'bz) && S_AXIS_DIN_TDATA[357]; // rv 0
  assign S_AXIS_DIN_TDATA_in[358] = (S_AXIS_DIN_TDATA[358] !== 1'bz) && S_AXIS_DIN_TDATA[358]; // rv 0
  assign S_AXIS_DIN_TDATA_in[359] = (S_AXIS_DIN_TDATA[359] !== 1'bz) && S_AXIS_DIN_TDATA[359]; // rv 0
  assign S_AXIS_DIN_TDATA_in[35] = (S_AXIS_DIN_TDATA[35] !== 1'bz) && S_AXIS_DIN_TDATA[35]; // rv 0
  assign S_AXIS_DIN_TDATA_in[360] = (S_AXIS_DIN_TDATA[360] !== 1'bz) && S_AXIS_DIN_TDATA[360]; // rv 0
  assign S_AXIS_DIN_TDATA_in[361] = (S_AXIS_DIN_TDATA[361] !== 1'bz) && S_AXIS_DIN_TDATA[361]; // rv 0
  assign S_AXIS_DIN_TDATA_in[362] = (S_AXIS_DIN_TDATA[362] !== 1'bz) && S_AXIS_DIN_TDATA[362]; // rv 0
  assign S_AXIS_DIN_TDATA_in[363] = (S_AXIS_DIN_TDATA[363] !== 1'bz) && S_AXIS_DIN_TDATA[363]; // rv 0
  assign S_AXIS_DIN_TDATA_in[364] = (S_AXIS_DIN_TDATA[364] !== 1'bz) && S_AXIS_DIN_TDATA[364]; // rv 0
  assign S_AXIS_DIN_TDATA_in[365] = (S_AXIS_DIN_TDATA[365] !== 1'bz) && S_AXIS_DIN_TDATA[365]; // rv 0
  assign S_AXIS_DIN_TDATA_in[366] = (S_AXIS_DIN_TDATA[366] !== 1'bz) && S_AXIS_DIN_TDATA[366]; // rv 0
  assign S_AXIS_DIN_TDATA_in[367] = (S_AXIS_DIN_TDATA[367] !== 1'bz) && S_AXIS_DIN_TDATA[367]; // rv 0
  assign S_AXIS_DIN_TDATA_in[368] = (S_AXIS_DIN_TDATA[368] !== 1'bz) && S_AXIS_DIN_TDATA[368]; // rv 0
  assign S_AXIS_DIN_TDATA_in[369] = (S_AXIS_DIN_TDATA[369] !== 1'bz) && S_AXIS_DIN_TDATA[369]; // rv 0
  assign S_AXIS_DIN_TDATA_in[36] = (S_AXIS_DIN_TDATA[36] !== 1'bz) && S_AXIS_DIN_TDATA[36]; // rv 0
  assign S_AXIS_DIN_TDATA_in[370] = (S_AXIS_DIN_TDATA[370] !== 1'bz) && S_AXIS_DIN_TDATA[370]; // rv 0
  assign S_AXIS_DIN_TDATA_in[371] = (S_AXIS_DIN_TDATA[371] !== 1'bz) && S_AXIS_DIN_TDATA[371]; // rv 0
  assign S_AXIS_DIN_TDATA_in[372] = (S_AXIS_DIN_TDATA[372] !== 1'bz) && S_AXIS_DIN_TDATA[372]; // rv 0
  assign S_AXIS_DIN_TDATA_in[373] = (S_AXIS_DIN_TDATA[373] !== 1'bz) && S_AXIS_DIN_TDATA[373]; // rv 0
  assign S_AXIS_DIN_TDATA_in[374] = (S_AXIS_DIN_TDATA[374] !== 1'bz) && S_AXIS_DIN_TDATA[374]; // rv 0
  assign S_AXIS_DIN_TDATA_in[375] = (S_AXIS_DIN_TDATA[375] !== 1'bz) && S_AXIS_DIN_TDATA[375]; // rv 0
  assign S_AXIS_DIN_TDATA_in[376] = (S_AXIS_DIN_TDATA[376] !== 1'bz) && S_AXIS_DIN_TDATA[376]; // rv 0
  assign S_AXIS_DIN_TDATA_in[377] = (S_AXIS_DIN_TDATA[377] !== 1'bz) && S_AXIS_DIN_TDATA[377]; // rv 0
  assign S_AXIS_DIN_TDATA_in[378] = (S_AXIS_DIN_TDATA[378] !== 1'bz) && S_AXIS_DIN_TDATA[378]; // rv 0
  assign S_AXIS_DIN_TDATA_in[379] = (S_AXIS_DIN_TDATA[379] !== 1'bz) && S_AXIS_DIN_TDATA[379]; // rv 0
  assign S_AXIS_DIN_TDATA_in[37] = (S_AXIS_DIN_TDATA[37] !== 1'bz) && S_AXIS_DIN_TDATA[37]; // rv 0
  assign S_AXIS_DIN_TDATA_in[380] = (S_AXIS_DIN_TDATA[380] !== 1'bz) && S_AXIS_DIN_TDATA[380]; // rv 0
  assign S_AXIS_DIN_TDATA_in[381] = (S_AXIS_DIN_TDATA[381] !== 1'bz) && S_AXIS_DIN_TDATA[381]; // rv 0
  assign S_AXIS_DIN_TDATA_in[382] = (S_AXIS_DIN_TDATA[382] !== 1'bz) && S_AXIS_DIN_TDATA[382]; // rv 0
  assign S_AXIS_DIN_TDATA_in[383] = (S_AXIS_DIN_TDATA[383] !== 1'bz) && S_AXIS_DIN_TDATA[383]; // rv 0
  assign S_AXIS_DIN_TDATA_in[384] = (S_AXIS_DIN_TDATA[384] !== 1'bz) && S_AXIS_DIN_TDATA[384]; // rv 0
  assign S_AXIS_DIN_TDATA_in[385] = (S_AXIS_DIN_TDATA[385] !== 1'bz) && S_AXIS_DIN_TDATA[385]; // rv 0
  assign S_AXIS_DIN_TDATA_in[386] = (S_AXIS_DIN_TDATA[386] !== 1'bz) && S_AXIS_DIN_TDATA[386]; // rv 0
  assign S_AXIS_DIN_TDATA_in[387] = (S_AXIS_DIN_TDATA[387] !== 1'bz) && S_AXIS_DIN_TDATA[387]; // rv 0
  assign S_AXIS_DIN_TDATA_in[388] = (S_AXIS_DIN_TDATA[388] !== 1'bz) && S_AXIS_DIN_TDATA[388]; // rv 0
  assign S_AXIS_DIN_TDATA_in[389] = (S_AXIS_DIN_TDATA[389] !== 1'bz) && S_AXIS_DIN_TDATA[389]; // rv 0
  assign S_AXIS_DIN_TDATA_in[38] = (S_AXIS_DIN_TDATA[38] !== 1'bz) && S_AXIS_DIN_TDATA[38]; // rv 0
  assign S_AXIS_DIN_TDATA_in[390] = (S_AXIS_DIN_TDATA[390] !== 1'bz) && S_AXIS_DIN_TDATA[390]; // rv 0
  assign S_AXIS_DIN_TDATA_in[391] = (S_AXIS_DIN_TDATA[391] !== 1'bz) && S_AXIS_DIN_TDATA[391]; // rv 0
  assign S_AXIS_DIN_TDATA_in[392] = (S_AXIS_DIN_TDATA[392] !== 1'bz) && S_AXIS_DIN_TDATA[392]; // rv 0
  assign S_AXIS_DIN_TDATA_in[393] = (S_AXIS_DIN_TDATA[393] !== 1'bz) && S_AXIS_DIN_TDATA[393]; // rv 0
  assign S_AXIS_DIN_TDATA_in[394] = (S_AXIS_DIN_TDATA[394] !== 1'bz) && S_AXIS_DIN_TDATA[394]; // rv 0
  assign S_AXIS_DIN_TDATA_in[395] = (S_AXIS_DIN_TDATA[395] !== 1'bz) && S_AXIS_DIN_TDATA[395]; // rv 0
  assign S_AXIS_DIN_TDATA_in[396] = (S_AXIS_DIN_TDATA[396] !== 1'bz) && S_AXIS_DIN_TDATA[396]; // rv 0
  assign S_AXIS_DIN_TDATA_in[397] = (S_AXIS_DIN_TDATA[397] !== 1'bz) && S_AXIS_DIN_TDATA[397]; // rv 0
  assign S_AXIS_DIN_TDATA_in[398] = (S_AXIS_DIN_TDATA[398] !== 1'bz) && S_AXIS_DIN_TDATA[398]; // rv 0
  assign S_AXIS_DIN_TDATA_in[399] = (S_AXIS_DIN_TDATA[399] !== 1'bz) && S_AXIS_DIN_TDATA[399]; // rv 0
  assign S_AXIS_DIN_TDATA_in[39] = (S_AXIS_DIN_TDATA[39] !== 1'bz) && S_AXIS_DIN_TDATA[39]; // rv 0
  assign S_AXIS_DIN_TDATA_in[3] = (S_AXIS_DIN_TDATA[3] !== 1'bz) && S_AXIS_DIN_TDATA[3]; // rv 0
  assign S_AXIS_DIN_TDATA_in[400] = (S_AXIS_DIN_TDATA[400] !== 1'bz) && S_AXIS_DIN_TDATA[400]; // rv 0
  assign S_AXIS_DIN_TDATA_in[401] = (S_AXIS_DIN_TDATA[401] !== 1'bz) && S_AXIS_DIN_TDATA[401]; // rv 0
  assign S_AXIS_DIN_TDATA_in[402] = (S_AXIS_DIN_TDATA[402] !== 1'bz) && S_AXIS_DIN_TDATA[402]; // rv 0
  assign S_AXIS_DIN_TDATA_in[403] = (S_AXIS_DIN_TDATA[403] !== 1'bz) && S_AXIS_DIN_TDATA[403]; // rv 0
  assign S_AXIS_DIN_TDATA_in[404] = (S_AXIS_DIN_TDATA[404] !== 1'bz) && S_AXIS_DIN_TDATA[404]; // rv 0
  assign S_AXIS_DIN_TDATA_in[405] = (S_AXIS_DIN_TDATA[405] !== 1'bz) && S_AXIS_DIN_TDATA[405]; // rv 0
  assign S_AXIS_DIN_TDATA_in[406] = (S_AXIS_DIN_TDATA[406] !== 1'bz) && S_AXIS_DIN_TDATA[406]; // rv 0
  assign S_AXIS_DIN_TDATA_in[407] = (S_AXIS_DIN_TDATA[407] !== 1'bz) && S_AXIS_DIN_TDATA[407]; // rv 0
  assign S_AXIS_DIN_TDATA_in[408] = (S_AXIS_DIN_TDATA[408] !== 1'bz) && S_AXIS_DIN_TDATA[408]; // rv 0
  assign S_AXIS_DIN_TDATA_in[409] = (S_AXIS_DIN_TDATA[409] !== 1'bz) && S_AXIS_DIN_TDATA[409]; // rv 0
  assign S_AXIS_DIN_TDATA_in[40] = (S_AXIS_DIN_TDATA[40] !== 1'bz) && S_AXIS_DIN_TDATA[40]; // rv 0
  assign S_AXIS_DIN_TDATA_in[410] = (S_AXIS_DIN_TDATA[410] !== 1'bz) && S_AXIS_DIN_TDATA[410]; // rv 0
  assign S_AXIS_DIN_TDATA_in[411] = (S_AXIS_DIN_TDATA[411] !== 1'bz) && S_AXIS_DIN_TDATA[411]; // rv 0
  assign S_AXIS_DIN_TDATA_in[412] = (S_AXIS_DIN_TDATA[412] !== 1'bz) && S_AXIS_DIN_TDATA[412]; // rv 0
  assign S_AXIS_DIN_TDATA_in[413] = (S_AXIS_DIN_TDATA[413] !== 1'bz) && S_AXIS_DIN_TDATA[413]; // rv 0
  assign S_AXIS_DIN_TDATA_in[414] = (S_AXIS_DIN_TDATA[414] !== 1'bz) && S_AXIS_DIN_TDATA[414]; // rv 0
  assign S_AXIS_DIN_TDATA_in[415] = (S_AXIS_DIN_TDATA[415] !== 1'bz) && S_AXIS_DIN_TDATA[415]; // rv 0
  assign S_AXIS_DIN_TDATA_in[416] = (S_AXIS_DIN_TDATA[416] !== 1'bz) && S_AXIS_DIN_TDATA[416]; // rv 0
  assign S_AXIS_DIN_TDATA_in[417] = (S_AXIS_DIN_TDATA[417] !== 1'bz) && S_AXIS_DIN_TDATA[417]; // rv 0
  assign S_AXIS_DIN_TDATA_in[418] = (S_AXIS_DIN_TDATA[418] !== 1'bz) && S_AXIS_DIN_TDATA[418]; // rv 0
  assign S_AXIS_DIN_TDATA_in[419] = (S_AXIS_DIN_TDATA[419] !== 1'bz) && S_AXIS_DIN_TDATA[419]; // rv 0
  assign S_AXIS_DIN_TDATA_in[41] = (S_AXIS_DIN_TDATA[41] !== 1'bz) && S_AXIS_DIN_TDATA[41]; // rv 0
  assign S_AXIS_DIN_TDATA_in[420] = (S_AXIS_DIN_TDATA[420] !== 1'bz) && S_AXIS_DIN_TDATA[420]; // rv 0
  assign S_AXIS_DIN_TDATA_in[421] = (S_AXIS_DIN_TDATA[421] !== 1'bz) && S_AXIS_DIN_TDATA[421]; // rv 0
  assign S_AXIS_DIN_TDATA_in[422] = (S_AXIS_DIN_TDATA[422] !== 1'bz) && S_AXIS_DIN_TDATA[422]; // rv 0
  assign S_AXIS_DIN_TDATA_in[423] = (S_AXIS_DIN_TDATA[423] !== 1'bz) && S_AXIS_DIN_TDATA[423]; // rv 0
  assign S_AXIS_DIN_TDATA_in[424] = (S_AXIS_DIN_TDATA[424] !== 1'bz) && S_AXIS_DIN_TDATA[424]; // rv 0
  assign S_AXIS_DIN_TDATA_in[425] = (S_AXIS_DIN_TDATA[425] !== 1'bz) && S_AXIS_DIN_TDATA[425]; // rv 0
  assign S_AXIS_DIN_TDATA_in[426] = (S_AXIS_DIN_TDATA[426] !== 1'bz) && S_AXIS_DIN_TDATA[426]; // rv 0
  assign S_AXIS_DIN_TDATA_in[427] = (S_AXIS_DIN_TDATA[427] !== 1'bz) && S_AXIS_DIN_TDATA[427]; // rv 0
  assign S_AXIS_DIN_TDATA_in[428] = (S_AXIS_DIN_TDATA[428] !== 1'bz) && S_AXIS_DIN_TDATA[428]; // rv 0
  assign S_AXIS_DIN_TDATA_in[429] = (S_AXIS_DIN_TDATA[429] !== 1'bz) && S_AXIS_DIN_TDATA[429]; // rv 0
  assign S_AXIS_DIN_TDATA_in[42] = (S_AXIS_DIN_TDATA[42] !== 1'bz) && S_AXIS_DIN_TDATA[42]; // rv 0
  assign S_AXIS_DIN_TDATA_in[430] = (S_AXIS_DIN_TDATA[430] !== 1'bz) && S_AXIS_DIN_TDATA[430]; // rv 0
  assign S_AXIS_DIN_TDATA_in[431] = (S_AXIS_DIN_TDATA[431] !== 1'bz) && S_AXIS_DIN_TDATA[431]; // rv 0
  assign S_AXIS_DIN_TDATA_in[432] = (S_AXIS_DIN_TDATA[432] !== 1'bz) && S_AXIS_DIN_TDATA[432]; // rv 0
  assign S_AXIS_DIN_TDATA_in[433] = (S_AXIS_DIN_TDATA[433] !== 1'bz) && S_AXIS_DIN_TDATA[433]; // rv 0
  assign S_AXIS_DIN_TDATA_in[434] = (S_AXIS_DIN_TDATA[434] !== 1'bz) && S_AXIS_DIN_TDATA[434]; // rv 0
  assign S_AXIS_DIN_TDATA_in[435] = (S_AXIS_DIN_TDATA[435] !== 1'bz) && S_AXIS_DIN_TDATA[435]; // rv 0
  assign S_AXIS_DIN_TDATA_in[436] = (S_AXIS_DIN_TDATA[436] !== 1'bz) && S_AXIS_DIN_TDATA[436]; // rv 0
  assign S_AXIS_DIN_TDATA_in[437] = (S_AXIS_DIN_TDATA[437] !== 1'bz) && S_AXIS_DIN_TDATA[437]; // rv 0
  assign S_AXIS_DIN_TDATA_in[438] = (S_AXIS_DIN_TDATA[438] !== 1'bz) && S_AXIS_DIN_TDATA[438]; // rv 0
  assign S_AXIS_DIN_TDATA_in[439] = (S_AXIS_DIN_TDATA[439] !== 1'bz) && S_AXIS_DIN_TDATA[439]; // rv 0
  assign S_AXIS_DIN_TDATA_in[43] = (S_AXIS_DIN_TDATA[43] !== 1'bz) && S_AXIS_DIN_TDATA[43]; // rv 0
  assign S_AXIS_DIN_TDATA_in[440] = (S_AXIS_DIN_TDATA[440] !== 1'bz) && S_AXIS_DIN_TDATA[440]; // rv 0
  assign S_AXIS_DIN_TDATA_in[441] = (S_AXIS_DIN_TDATA[441] !== 1'bz) && S_AXIS_DIN_TDATA[441]; // rv 0
  assign S_AXIS_DIN_TDATA_in[442] = (S_AXIS_DIN_TDATA[442] !== 1'bz) && S_AXIS_DIN_TDATA[442]; // rv 0
  assign S_AXIS_DIN_TDATA_in[443] = (S_AXIS_DIN_TDATA[443] !== 1'bz) && S_AXIS_DIN_TDATA[443]; // rv 0
  assign S_AXIS_DIN_TDATA_in[444] = (S_AXIS_DIN_TDATA[444] !== 1'bz) && S_AXIS_DIN_TDATA[444]; // rv 0
  assign S_AXIS_DIN_TDATA_in[445] = (S_AXIS_DIN_TDATA[445] !== 1'bz) && S_AXIS_DIN_TDATA[445]; // rv 0
  assign S_AXIS_DIN_TDATA_in[446] = (S_AXIS_DIN_TDATA[446] !== 1'bz) && S_AXIS_DIN_TDATA[446]; // rv 0
  assign S_AXIS_DIN_TDATA_in[447] = (S_AXIS_DIN_TDATA[447] !== 1'bz) && S_AXIS_DIN_TDATA[447]; // rv 0
  assign S_AXIS_DIN_TDATA_in[448] = (S_AXIS_DIN_TDATA[448] !== 1'bz) && S_AXIS_DIN_TDATA[448]; // rv 0
  assign S_AXIS_DIN_TDATA_in[449] = (S_AXIS_DIN_TDATA[449] !== 1'bz) && S_AXIS_DIN_TDATA[449]; // rv 0
  assign S_AXIS_DIN_TDATA_in[44] = (S_AXIS_DIN_TDATA[44] !== 1'bz) && S_AXIS_DIN_TDATA[44]; // rv 0
  assign S_AXIS_DIN_TDATA_in[450] = (S_AXIS_DIN_TDATA[450] !== 1'bz) && S_AXIS_DIN_TDATA[450]; // rv 0
  assign S_AXIS_DIN_TDATA_in[451] = (S_AXIS_DIN_TDATA[451] !== 1'bz) && S_AXIS_DIN_TDATA[451]; // rv 0
  assign S_AXIS_DIN_TDATA_in[452] = (S_AXIS_DIN_TDATA[452] !== 1'bz) && S_AXIS_DIN_TDATA[452]; // rv 0
  assign S_AXIS_DIN_TDATA_in[453] = (S_AXIS_DIN_TDATA[453] !== 1'bz) && S_AXIS_DIN_TDATA[453]; // rv 0
  assign S_AXIS_DIN_TDATA_in[454] = (S_AXIS_DIN_TDATA[454] !== 1'bz) && S_AXIS_DIN_TDATA[454]; // rv 0
  assign S_AXIS_DIN_TDATA_in[455] = (S_AXIS_DIN_TDATA[455] !== 1'bz) && S_AXIS_DIN_TDATA[455]; // rv 0
  assign S_AXIS_DIN_TDATA_in[456] = (S_AXIS_DIN_TDATA[456] !== 1'bz) && S_AXIS_DIN_TDATA[456]; // rv 0
  assign S_AXIS_DIN_TDATA_in[457] = (S_AXIS_DIN_TDATA[457] !== 1'bz) && S_AXIS_DIN_TDATA[457]; // rv 0
  assign S_AXIS_DIN_TDATA_in[458] = (S_AXIS_DIN_TDATA[458] !== 1'bz) && S_AXIS_DIN_TDATA[458]; // rv 0
  assign S_AXIS_DIN_TDATA_in[459] = (S_AXIS_DIN_TDATA[459] !== 1'bz) && S_AXIS_DIN_TDATA[459]; // rv 0
  assign S_AXIS_DIN_TDATA_in[45] = (S_AXIS_DIN_TDATA[45] !== 1'bz) && S_AXIS_DIN_TDATA[45]; // rv 0
  assign S_AXIS_DIN_TDATA_in[460] = (S_AXIS_DIN_TDATA[460] !== 1'bz) && S_AXIS_DIN_TDATA[460]; // rv 0
  assign S_AXIS_DIN_TDATA_in[461] = (S_AXIS_DIN_TDATA[461] !== 1'bz) && S_AXIS_DIN_TDATA[461]; // rv 0
  assign S_AXIS_DIN_TDATA_in[462] = (S_AXIS_DIN_TDATA[462] !== 1'bz) && S_AXIS_DIN_TDATA[462]; // rv 0
  assign S_AXIS_DIN_TDATA_in[463] = (S_AXIS_DIN_TDATA[463] !== 1'bz) && S_AXIS_DIN_TDATA[463]; // rv 0
  assign S_AXIS_DIN_TDATA_in[464] = (S_AXIS_DIN_TDATA[464] !== 1'bz) && S_AXIS_DIN_TDATA[464]; // rv 0
  assign S_AXIS_DIN_TDATA_in[465] = (S_AXIS_DIN_TDATA[465] !== 1'bz) && S_AXIS_DIN_TDATA[465]; // rv 0
  assign S_AXIS_DIN_TDATA_in[466] = (S_AXIS_DIN_TDATA[466] !== 1'bz) && S_AXIS_DIN_TDATA[466]; // rv 0
  assign S_AXIS_DIN_TDATA_in[467] = (S_AXIS_DIN_TDATA[467] !== 1'bz) && S_AXIS_DIN_TDATA[467]; // rv 0
  assign S_AXIS_DIN_TDATA_in[468] = (S_AXIS_DIN_TDATA[468] !== 1'bz) && S_AXIS_DIN_TDATA[468]; // rv 0
  assign S_AXIS_DIN_TDATA_in[469] = (S_AXIS_DIN_TDATA[469] !== 1'bz) && S_AXIS_DIN_TDATA[469]; // rv 0
  assign S_AXIS_DIN_TDATA_in[46] = (S_AXIS_DIN_TDATA[46] !== 1'bz) && S_AXIS_DIN_TDATA[46]; // rv 0
  assign S_AXIS_DIN_TDATA_in[470] = (S_AXIS_DIN_TDATA[470] !== 1'bz) && S_AXIS_DIN_TDATA[470]; // rv 0
  assign S_AXIS_DIN_TDATA_in[471] = (S_AXIS_DIN_TDATA[471] !== 1'bz) && S_AXIS_DIN_TDATA[471]; // rv 0
  assign S_AXIS_DIN_TDATA_in[472] = (S_AXIS_DIN_TDATA[472] !== 1'bz) && S_AXIS_DIN_TDATA[472]; // rv 0
  assign S_AXIS_DIN_TDATA_in[473] = (S_AXIS_DIN_TDATA[473] !== 1'bz) && S_AXIS_DIN_TDATA[473]; // rv 0
  assign S_AXIS_DIN_TDATA_in[474] = (S_AXIS_DIN_TDATA[474] !== 1'bz) && S_AXIS_DIN_TDATA[474]; // rv 0
  assign S_AXIS_DIN_TDATA_in[475] = (S_AXIS_DIN_TDATA[475] !== 1'bz) && S_AXIS_DIN_TDATA[475]; // rv 0
  assign S_AXIS_DIN_TDATA_in[476] = (S_AXIS_DIN_TDATA[476] !== 1'bz) && S_AXIS_DIN_TDATA[476]; // rv 0
  assign S_AXIS_DIN_TDATA_in[477] = (S_AXIS_DIN_TDATA[477] !== 1'bz) && S_AXIS_DIN_TDATA[477]; // rv 0
  assign S_AXIS_DIN_TDATA_in[478] = (S_AXIS_DIN_TDATA[478] !== 1'bz) && S_AXIS_DIN_TDATA[478]; // rv 0
  assign S_AXIS_DIN_TDATA_in[479] = (S_AXIS_DIN_TDATA[479] !== 1'bz) && S_AXIS_DIN_TDATA[479]; // rv 0
  assign S_AXIS_DIN_TDATA_in[47] = (S_AXIS_DIN_TDATA[47] !== 1'bz) && S_AXIS_DIN_TDATA[47]; // rv 0
  assign S_AXIS_DIN_TDATA_in[480] = (S_AXIS_DIN_TDATA[480] !== 1'bz) && S_AXIS_DIN_TDATA[480]; // rv 0
  assign S_AXIS_DIN_TDATA_in[481] = (S_AXIS_DIN_TDATA[481] !== 1'bz) && S_AXIS_DIN_TDATA[481]; // rv 0
  assign S_AXIS_DIN_TDATA_in[482] = (S_AXIS_DIN_TDATA[482] !== 1'bz) && S_AXIS_DIN_TDATA[482]; // rv 0
  assign S_AXIS_DIN_TDATA_in[483] = (S_AXIS_DIN_TDATA[483] !== 1'bz) && S_AXIS_DIN_TDATA[483]; // rv 0
  assign S_AXIS_DIN_TDATA_in[484] = (S_AXIS_DIN_TDATA[484] !== 1'bz) && S_AXIS_DIN_TDATA[484]; // rv 0
  assign S_AXIS_DIN_TDATA_in[485] = (S_AXIS_DIN_TDATA[485] !== 1'bz) && S_AXIS_DIN_TDATA[485]; // rv 0
  assign S_AXIS_DIN_TDATA_in[486] = (S_AXIS_DIN_TDATA[486] !== 1'bz) && S_AXIS_DIN_TDATA[486]; // rv 0
  assign S_AXIS_DIN_TDATA_in[487] = (S_AXIS_DIN_TDATA[487] !== 1'bz) && S_AXIS_DIN_TDATA[487]; // rv 0
  assign S_AXIS_DIN_TDATA_in[488] = (S_AXIS_DIN_TDATA[488] !== 1'bz) && S_AXIS_DIN_TDATA[488]; // rv 0
  assign S_AXIS_DIN_TDATA_in[489] = (S_AXIS_DIN_TDATA[489] !== 1'bz) && S_AXIS_DIN_TDATA[489]; // rv 0
  assign S_AXIS_DIN_TDATA_in[48] = (S_AXIS_DIN_TDATA[48] !== 1'bz) && S_AXIS_DIN_TDATA[48]; // rv 0
  assign S_AXIS_DIN_TDATA_in[490] = (S_AXIS_DIN_TDATA[490] !== 1'bz) && S_AXIS_DIN_TDATA[490]; // rv 0
  assign S_AXIS_DIN_TDATA_in[491] = (S_AXIS_DIN_TDATA[491] !== 1'bz) && S_AXIS_DIN_TDATA[491]; // rv 0
  assign S_AXIS_DIN_TDATA_in[492] = (S_AXIS_DIN_TDATA[492] !== 1'bz) && S_AXIS_DIN_TDATA[492]; // rv 0
  assign S_AXIS_DIN_TDATA_in[493] = (S_AXIS_DIN_TDATA[493] !== 1'bz) && S_AXIS_DIN_TDATA[493]; // rv 0
  assign S_AXIS_DIN_TDATA_in[494] = (S_AXIS_DIN_TDATA[494] !== 1'bz) && S_AXIS_DIN_TDATA[494]; // rv 0
  assign S_AXIS_DIN_TDATA_in[495] = (S_AXIS_DIN_TDATA[495] !== 1'bz) && S_AXIS_DIN_TDATA[495]; // rv 0
  assign S_AXIS_DIN_TDATA_in[496] = (S_AXIS_DIN_TDATA[496] !== 1'bz) && S_AXIS_DIN_TDATA[496]; // rv 0
  assign S_AXIS_DIN_TDATA_in[497] = (S_AXIS_DIN_TDATA[497] !== 1'bz) && S_AXIS_DIN_TDATA[497]; // rv 0
  assign S_AXIS_DIN_TDATA_in[498] = (S_AXIS_DIN_TDATA[498] !== 1'bz) && S_AXIS_DIN_TDATA[498]; // rv 0
  assign S_AXIS_DIN_TDATA_in[499] = (S_AXIS_DIN_TDATA[499] !== 1'bz) && S_AXIS_DIN_TDATA[499]; // rv 0
  assign S_AXIS_DIN_TDATA_in[49] = (S_AXIS_DIN_TDATA[49] !== 1'bz) && S_AXIS_DIN_TDATA[49]; // rv 0
  assign S_AXIS_DIN_TDATA_in[4] = (S_AXIS_DIN_TDATA[4] !== 1'bz) && S_AXIS_DIN_TDATA[4]; // rv 0
  assign S_AXIS_DIN_TDATA_in[500] = (S_AXIS_DIN_TDATA[500] !== 1'bz) && S_AXIS_DIN_TDATA[500]; // rv 0
  assign S_AXIS_DIN_TDATA_in[501] = (S_AXIS_DIN_TDATA[501] !== 1'bz) && S_AXIS_DIN_TDATA[501]; // rv 0
  assign S_AXIS_DIN_TDATA_in[502] = (S_AXIS_DIN_TDATA[502] !== 1'bz) && S_AXIS_DIN_TDATA[502]; // rv 0
  assign S_AXIS_DIN_TDATA_in[503] = (S_AXIS_DIN_TDATA[503] !== 1'bz) && S_AXIS_DIN_TDATA[503]; // rv 0
  assign S_AXIS_DIN_TDATA_in[504] = (S_AXIS_DIN_TDATA[504] !== 1'bz) && S_AXIS_DIN_TDATA[504]; // rv 0
  assign S_AXIS_DIN_TDATA_in[505] = (S_AXIS_DIN_TDATA[505] !== 1'bz) && S_AXIS_DIN_TDATA[505]; // rv 0
  assign S_AXIS_DIN_TDATA_in[506] = (S_AXIS_DIN_TDATA[506] !== 1'bz) && S_AXIS_DIN_TDATA[506]; // rv 0
  assign S_AXIS_DIN_TDATA_in[507] = (S_AXIS_DIN_TDATA[507] !== 1'bz) && S_AXIS_DIN_TDATA[507]; // rv 0
  assign S_AXIS_DIN_TDATA_in[508] = (S_AXIS_DIN_TDATA[508] !== 1'bz) && S_AXIS_DIN_TDATA[508]; // rv 0
  assign S_AXIS_DIN_TDATA_in[509] = (S_AXIS_DIN_TDATA[509] !== 1'bz) && S_AXIS_DIN_TDATA[509]; // rv 0
  assign S_AXIS_DIN_TDATA_in[50] = (S_AXIS_DIN_TDATA[50] !== 1'bz) && S_AXIS_DIN_TDATA[50]; // rv 0
  assign S_AXIS_DIN_TDATA_in[510] = (S_AXIS_DIN_TDATA[510] !== 1'bz) && S_AXIS_DIN_TDATA[510]; // rv 0
  assign S_AXIS_DIN_TDATA_in[511] = (S_AXIS_DIN_TDATA[511] !== 1'bz) && S_AXIS_DIN_TDATA[511]; // rv 0
  assign S_AXIS_DIN_TDATA_in[51] = (S_AXIS_DIN_TDATA[51] !== 1'bz) && S_AXIS_DIN_TDATA[51]; // rv 0
  assign S_AXIS_DIN_TDATA_in[52] = (S_AXIS_DIN_TDATA[52] !== 1'bz) && S_AXIS_DIN_TDATA[52]; // rv 0
  assign S_AXIS_DIN_TDATA_in[53] = (S_AXIS_DIN_TDATA[53] !== 1'bz) && S_AXIS_DIN_TDATA[53]; // rv 0
  assign S_AXIS_DIN_TDATA_in[54] = (S_AXIS_DIN_TDATA[54] !== 1'bz) && S_AXIS_DIN_TDATA[54]; // rv 0
  assign S_AXIS_DIN_TDATA_in[55] = (S_AXIS_DIN_TDATA[55] !== 1'bz) && S_AXIS_DIN_TDATA[55]; // rv 0
  assign S_AXIS_DIN_TDATA_in[56] = (S_AXIS_DIN_TDATA[56] !== 1'bz) && S_AXIS_DIN_TDATA[56]; // rv 0
  assign S_AXIS_DIN_TDATA_in[57] = (S_AXIS_DIN_TDATA[57] !== 1'bz) && S_AXIS_DIN_TDATA[57]; // rv 0
  assign S_AXIS_DIN_TDATA_in[58] = (S_AXIS_DIN_TDATA[58] !== 1'bz) && S_AXIS_DIN_TDATA[58]; // rv 0
  assign S_AXIS_DIN_TDATA_in[59] = (S_AXIS_DIN_TDATA[59] !== 1'bz) && S_AXIS_DIN_TDATA[59]; // rv 0
  assign S_AXIS_DIN_TDATA_in[5] = (S_AXIS_DIN_TDATA[5] !== 1'bz) && S_AXIS_DIN_TDATA[5]; // rv 0
  assign S_AXIS_DIN_TDATA_in[60] = (S_AXIS_DIN_TDATA[60] !== 1'bz) && S_AXIS_DIN_TDATA[60]; // rv 0
  assign S_AXIS_DIN_TDATA_in[61] = (S_AXIS_DIN_TDATA[61] !== 1'bz) && S_AXIS_DIN_TDATA[61]; // rv 0
  assign S_AXIS_DIN_TDATA_in[62] = (S_AXIS_DIN_TDATA[62] !== 1'bz) && S_AXIS_DIN_TDATA[62]; // rv 0
  assign S_AXIS_DIN_TDATA_in[63] = (S_AXIS_DIN_TDATA[63] !== 1'bz) && S_AXIS_DIN_TDATA[63]; // rv 0
  assign S_AXIS_DIN_TDATA_in[64] = (S_AXIS_DIN_TDATA[64] !== 1'bz) && S_AXIS_DIN_TDATA[64]; // rv 0
  assign S_AXIS_DIN_TDATA_in[65] = (S_AXIS_DIN_TDATA[65] !== 1'bz) && S_AXIS_DIN_TDATA[65]; // rv 0
  assign S_AXIS_DIN_TDATA_in[66] = (S_AXIS_DIN_TDATA[66] !== 1'bz) && S_AXIS_DIN_TDATA[66]; // rv 0
  assign S_AXIS_DIN_TDATA_in[67] = (S_AXIS_DIN_TDATA[67] !== 1'bz) && S_AXIS_DIN_TDATA[67]; // rv 0
  assign S_AXIS_DIN_TDATA_in[68] = (S_AXIS_DIN_TDATA[68] !== 1'bz) && S_AXIS_DIN_TDATA[68]; // rv 0
  assign S_AXIS_DIN_TDATA_in[69] = (S_AXIS_DIN_TDATA[69] !== 1'bz) && S_AXIS_DIN_TDATA[69]; // rv 0
  assign S_AXIS_DIN_TDATA_in[6] = (S_AXIS_DIN_TDATA[6] !== 1'bz) && S_AXIS_DIN_TDATA[6]; // rv 0
  assign S_AXIS_DIN_TDATA_in[70] = (S_AXIS_DIN_TDATA[70] !== 1'bz) && S_AXIS_DIN_TDATA[70]; // rv 0
  assign S_AXIS_DIN_TDATA_in[71] = (S_AXIS_DIN_TDATA[71] !== 1'bz) && S_AXIS_DIN_TDATA[71]; // rv 0
  assign S_AXIS_DIN_TDATA_in[72] = (S_AXIS_DIN_TDATA[72] !== 1'bz) && S_AXIS_DIN_TDATA[72]; // rv 0
  assign S_AXIS_DIN_TDATA_in[73] = (S_AXIS_DIN_TDATA[73] !== 1'bz) && S_AXIS_DIN_TDATA[73]; // rv 0
  assign S_AXIS_DIN_TDATA_in[74] = (S_AXIS_DIN_TDATA[74] !== 1'bz) && S_AXIS_DIN_TDATA[74]; // rv 0
  assign S_AXIS_DIN_TDATA_in[75] = (S_AXIS_DIN_TDATA[75] !== 1'bz) && S_AXIS_DIN_TDATA[75]; // rv 0
  assign S_AXIS_DIN_TDATA_in[76] = (S_AXIS_DIN_TDATA[76] !== 1'bz) && S_AXIS_DIN_TDATA[76]; // rv 0
  assign S_AXIS_DIN_TDATA_in[77] = (S_AXIS_DIN_TDATA[77] !== 1'bz) && S_AXIS_DIN_TDATA[77]; // rv 0
  assign S_AXIS_DIN_TDATA_in[78] = (S_AXIS_DIN_TDATA[78] !== 1'bz) && S_AXIS_DIN_TDATA[78]; // rv 0
  assign S_AXIS_DIN_TDATA_in[79] = (S_AXIS_DIN_TDATA[79] !== 1'bz) && S_AXIS_DIN_TDATA[79]; // rv 0
  assign S_AXIS_DIN_TDATA_in[7] = (S_AXIS_DIN_TDATA[7] !== 1'bz) && S_AXIS_DIN_TDATA[7]; // rv 0
  assign S_AXIS_DIN_TDATA_in[80] = (S_AXIS_DIN_TDATA[80] !== 1'bz) && S_AXIS_DIN_TDATA[80]; // rv 0
  assign S_AXIS_DIN_TDATA_in[81] = (S_AXIS_DIN_TDATA[81] !== 1'bz) && S_AXIS_DIN_TDATA[81]; // rv 0
  assign S_AXIS_DIN_TDATA_in[82] = (S_AXIS_DIN_TDATA[82] !== 1'bz) && S_AXIS_DIN_TDATA[82]; // rv 0
  assign S_AXIS_DIN_TDATA_in[83] = (S_AXIS_DIN_TDATA[83] !== 1'bz) && S_AXIS_DIN_TDATA[83]; // rv 0
  assign S_AXIS_DIN_TDATA_in[84] = (S_AXIS_DIN_TDATA[84] !== 1'bz) && S_AXIS_DIN_TDATA[84]; // rv 0
  assign S_AXIS_DIN_TDATA_in[85] = (S_AXIS_DIN_TDATA[85] !== 1'bz) && S_AXIS_DIN_TDATA[85]; // rv 0
  assign S_AXIS_DIN_TDATA_in[86] = (S_AXIS_DIN_TDATA[86] !== 1'bz) && S_AXIS_DIN_TDATA[86]; // rv 0
  assign S_AXIS_DIN_TDATA_in[87] = (S_AXIS_DIN_TDATA[87] !== 1'bz) && S_AXIS_DIN_TDATA[87]; // rv 0
  assign S_AXIS_DIN_TDATA_in[88] = (S_AXIS_DIN_TDATA[88] !== 1'bz) && S_AXIS_DIN_TDATA[88]; // rv 0
  assign S_AXIS_DIN_TDATA_in[89] = (S_AXIS_DIN_TDATA[89] !== 1'bz) && S_AXIS_DIN_TDATA[89]; // rv 0
  assign S_AXIS_DIN_TDATA_in[8] = (S_AXIS_DIN_TDATA[8] !== 1'bz) && S_AXIS_DIN_TDATA[8]; // rv 0
  assign S_AXIS_DIN_TDATA_in[90] = (S_AXIS_DIN_TDATA[90] !== 1'bz) && S_AXIS_DIN_TDATA[90]; // rv 0
  assign S_AXIS_DIN_TDATA_in[91] = (S_AXIS_DIN_TDATA[91] !== 1'bz) && S_AXIS_DIN_TDATA[91]; // rv 0
  assign S_AXIS_DIN_TDATA_in[92] = (S_AXIS_DIN_TDATA[92] !== 1'bz) && S_AXIS_DIN_TDATA[92]; // rv 0
  assign S_AXIS_DIN_TDATA_in[93] = (S_AXIS_DIN_TDATA[93] !== 1'bz) && S_AXIS_DIN_TDATA[93]; // rv 0
  assign S_AXIS_DIN_TDATA_in[94] = (S_AXIS_DIN_TDATA[94] !== 1'bz) && S_AXIS_DIN_TDATA[94]; // rv 0
  assign S_AXIS_DIN_TDATA_in[95] = (S_AXIS_DIN_TDATA[95] !== 1'bz) && S_AXIS_DIN_TDATA[95]; // rv 0
  assign S_AXIS_DIN_TDATA_in[96] = (S_AXIS_DIN_TDATA[96] !== 1'bz) && S_AXIS_DIN_TDATA[96]; // rv 0
  assign S_AXIS_DIN_TDATA_in[97] = (S_AXIS_DIN_TDATA[97] !== 1'bz) && S_AXIS_DIN_TDATA[97]; // rv 0
  assign S_AXIS_DIN_TDATA_in[98] = (S_AXIS_DIN_TDATA[98] !== 1'bz) && S_AXIS_DIN_TDATA[98]; // rv 0
  assign S_AXIS_DIN_TDATA_in[99] = (S_AXIS_DIN_TDATA[99] !== 1'bz) && S_AXIS_DIN_TDATA[99]; // rv 0
  assign S_AXIS_DIN_TDATA_in[9] = (S_AXIS_DIN_TDATA[9] !== 1'bz) && S_AXIS_DIN_TDATA[9]; // rv 0
  assign S_AXIS_DIN_TLAST_in = (S_AXIS_DIN_TLAST !== 1'bz) && S_AXIS_DIN_TLAST; // rv 0
  assign S_AXIS_DIN_TVALID_in = (S_AXIS_DIN_TVALID !== 1'bz) && S_AXIS_DIN_TVALID; // rv 0
  assign S_AXIS_DIN_WORDS_ACLK_in = (S_AXIS_DIN_WORDS_ACLK !== 1'bz) && S_AXIS_DIN_WORDS_ACLK; // rv 0
  assign S_AXIS_DIN_WORDS_TDATA_in[0] = (S_AXIS_DIN_WORDS_TDATA[0] !== 1'bz) && S_AXIS_DIN_WORDS_TDATA[0]; // rv 0
  assign S_AXIS_DIN_WORDS_TDATA_in[10] = (S_AXIS_DIN_WORDS_TDATA[10] !== 1'bz) && S_AXIS_DIN_WORDS_TDATA[10]; // rv 0
  assign S_AXIS_DIN_WORDS_TDATA_in[11] = (S_AXIS_DIN_WORDS_TDATA[11] !== 1'bz) && S_AXIS_DIN_WORDS_TDATA[11]; // rv 0
  assign S_AXIS_DIN_WORDS_TDATA_in[12] = (S_AXIS_DIN_WORDS_TDATA[12] !== 1'bz) && S_AXIS_DIN_WORDS_TDATA[12]; // rv 0
  assign S_AXIS_DIN_WORDS_TDATA_in[13] = (S_AXIS_DIN_WORDS_TDATA[13] !== 1'bz) && S_AXIS_DIN_WORDS_TDATA[13]; // rv 0
  assign S_AXIS_DIN_WORDS_TDATA_in[14] = (S_AXIS_DIN_WORDS_TDATA[14] !== 1'bz) && S_AXIS_DIN_WORDS_TDATA[14]; // rv 0
  assign S_AXIS_DIN_WORDS_TDATA_in[15] = (S_AXIS_DIN_WORDS_TDATA[15] !== 1'bz) && S_AXIS_DIN_WORDS_TDATA[15]; // rv 0
  assign S_AXIS_DIN_WORDS_TDATA_in[16] = (S_AXIS_DIN_WORDS_TDATA[16] !== 1'bz) && S_AXIS_DIN_WORDS_TDATA[16]; // rv 0
  assign S_AXIS_DIN_WORDS_TDATA_in[17] = (S_AXIS_DIN_WORDS_TDATA[17] !== 1'bz) && S_AXIS_DIN_WORDS_TDATA[17]; // rv 0
  assign S_AXIS_DIN_WORDS_TDATA_in[18] = (S_AXIS_DIN_WORDS_TDATA[18] !== 1'bz) && S_AXIS_DIN_WORDS_TDATA[18]; // rv 0
  assign S_AXIS_DIN_WORDS_TDATA_in[19] = (S_AXIS_DIN_WORDS_TDATA[19] !== 1'bz) && S_AXIS_DIN_WORDS_TDATA[19]; // rv 0
  assign S_AXIS_DIN_WORDS_TDATA_in[1] = (S_AXIS_DIN_WORDS_TDATA[1] !== 1'bz) && S_AXIS_DIN_WORDS_TDATA[1]; // rv 0
  assign S_AXIS_DIN_WORDS_TDATA_in[20] = (S_AXIS_DIN_WORDS_TDATA[20] !== 1'bz) && S_AXIS_DIN_WORDS_TDATA[20]; // rv 0
  assign S_AXIS_DIN_WORDS_TDATA_in[21] = (S_AXIS_DIN_WORDS_TDATA[21] !== 1'bz) && S_AXIS_DIN_WORDS_TDATA[21]; // rv 0
  assign S_AXIS_DIN_WORDS_TDATA_in[22] = (S_AXIS_DIN_WORDS_TDATA[22] !== 1'bz) && S_AXIS_DIN_WORDS_TDATA[22]; // rv 0
  assign S_AXIS_DIN_WORDS_TDATA_in[23] = (S_AXIS_DIN_WORDS_TDATA[23] !== 1'bz) && S_AXIS_DIN_WORDS_TDATA[23]; // rv 0
  assign S_AXIS_DIN_WORDS_TDATA_in[24] = (S_AXIS_DIN_WORDS_TDATA[24] !== 1'bz) && S_AXIS_DIN_WORDS_TDATA[24]; // rv 0
  assign S_AXIS_DIN_WORDS_TDATA_in[25] = (S_AXIS_DIN_WORDS_TDATA[25] !== 1'bz) && S_AXIS_DIN_WORDS_TDATA[25]; // rv 0
  assign S_AXIS_DIN_WORDS_TDATA_in[26] = (S_AXIS_DIN_WORDS_TDATA[26] !== 1'bz) && S_AXIS_DIN_WORDS_TDATA[26]; // rv 0
  assign S_AXIS_DIN_WORDS_TDATA_in[27] = (S_AXIS_DIN_WORDS_TDATA[27] !== 1'bz) && S_AXIS_DIN_WORDS_TDATA[27]; // rv 0
  assign S_AXIS_DIN_WORDS_TDATA_in[28] = (S_AXIS_DIN_WORDS_TDATA[28] !== 1'bz) && S_AXIS_DIN_WORDS_TDATA[28]; // rv 0
  assign S_AXIS_DIN_WORDS_TDATA_in[29] = (S_AXIS_DIN_WORDS_TDATA[29] !== 1'bz) && S_AXIS_DIN_WORDS_TDATA[29]; // rv 0
  assign S_AXIS_DIN_WORDS_TDATA_in[2] = (S_AXIS_DIN_WORDS_TDATA[2] !== 1'bz) && S_AXIS_DIN_WORDS_TDATA[2]; // rv 0
  assign S_AXIS_DIN_WORDS_TDATA_in[30] = (S_AXIS_DIN_WORDS_TDATA[30] !== 1'bz) && S_AXIS_DIN_WORDS_TDATA[30]; // rv 0
  assign S_AXIS_DIN_WORDS_TDATA_in[31] = (S_AXIS_DIN_WORDS_TDATA[31] !== 1'bz) && S_AXIS_DIN_WORDS_TDATA[31]; // rv 0
  assign S_AXIS_DIN_WORDS_TDATA_in[3] = (S_AXIS_DIN_WORDS_TDATA[3] !== 1'bz) && S_AXIS_DIN_WORDS_TDATA[3]; // rv 0
  assign S_AXIS_DIN_WORDS_TDATA_in[4] = (S_AXIS_DIN_WORDS_TDATA[4] !== 1'bz) && S_AXIS_DIN_WORDS_TDATA[4]; // rv 0
  assign S_AXIS_DIN_WORDS_TDATA_in[5] = (S_AXIS_DIN_WORDS_TDATA[5] !== 1'bz) && S_AXIS_DIN_WORDS_TDATA[5]; // rv 0
  assign S_AXIS_DIN_WORDS_TDATA_in[6] = (S_AXIS_DIN_WORDS_TDATA[6] !== 1'bz) && S_AXIS_DIN_WORDS_TDATA[6]; // rv 0
  assign S_AXIS_DIN_WORDS_TDATA_in[7] = (S_AXIS_DIN_WORDS_TDATA[7] !== 1'bz) && S_AXIS_DIN_WORDS_TDATA[7]; // rv 0
  assign S_AXIS_DIN_WORDS_TDATA_in[8] = (S_AXIS_DIN_WORDS_TDATA[8] !== 1'bz) && S_AXIS_DIN_WORDS_TDATA[8]; // rv 0
  assign S_AXIS_DIN_WORDS_TDATA_in[9] = (S_AXIS_DIN_WORDS_TDATA[9] !== 1'bz) && S_AXIS_DIN_WORDS_TDATA[9]; // rv 0
  assign S_AXIS_DIN_WORDS_TLAST_in = (S_AXIS_DIN_WORDS_TLAST !== 1'bz) && S_AXIS_DIN_WORDS_TLAST; // rv 0
  assign S_AXIS_DIN_WORDS_TVALID_in = (S_AXIS_DIN_WORDS_TVALID !== 1'bz) && S_AXIS_DIN_WORDS_TVALID; // rv 0
  assign S_AXIS_DOUT_WORDS_ACLK_in = (S_AXIS_DOUT_WORDS_ACLK !== 1'bz) && S_AXIS_DOUT_WORDS_ACLK; // rv 0
  assign S_AXIS_DOUT_WORDS_TDATA_in[0] = (S_AXIS_DOUT_WORDS_TDATA[0] !== 1'bz) && S_AXIS_DOUT_WORDS_TDATA[0]; // rv 0
  assign S_AXIS_DOUT_WORDS_TDATA_in[10] = (S_AXIS_DOUT_WORDS_TDATA[10] !== 1'bz) && S_AXIS_DOUT_WORDS_TDATA[10]; // rv 0
  assign S_AXIS_DOUT_WORDS_TDATA_in[11] = (S_AXIS_DOUT_WORDS_TDATA[11] !== 1'bz) && S_AXIS_DOUT_WORDS_TDATA[11]; // rv 0
  assign S_AXIS_DOUT_WORDS_TDATA_in[12] = (S_AXIS_DOUT_WORDS_TDATA[12] !== 1'bz) && S_AXIS_DOUT_WORDS_TDATA[12]; // rv 0
  assign S_AXIS_DOUT_WORDS_TDATA_in[13] = (S_AXIS_DOUT_WORDS_TDATA[13] !== 1'bz) && S_AXIS_DOUT_WORDS_TDATA[13]; // rv 0
  assign S_AXIS_DOUT_WORDS_TDATA_in[14] = (S_AXIS_DOUT_WORDS_TDATA[14] !== 1'bz) && S_AXIS_DOUT_WORDS_TDATA[14]; // rv 0
  assign S_AXIS_DOUT_WORDS_TDATA_in[15] = (S_AXIS_DOUT_WORDS_TDATA[15] !== 1'bz) && S_AXIS_DOUT_WORDS_TDATA[15]; // rv 0
  assign S_AXIS_DOUT_WORDS_TDATA_in[16] = (S_AXIS_DOUT_WORDS_TDATA[16] !== 1'bz) && S_AXIS_DOUT_WORDS_TDATA[16]; // rv 0
  assign S_AXIS_DOUT_WORDS_TDATA_in[17] = (S_AXIS_DOUT_WORDS_TDATA[17] !== 1'bz) && S_AXIS_DOUT_WORDS_TDATA[17]; // rv 0
  assign S_AXIS_DOUT_WORDS_TDATA_in[18] = (S_AXIS_DOUT_WORDS_TDATA[18] !== 1'bz) && S_AXIS_DOUT_WORDS_TDATA[18]; // rv 0
  assign S_AXIS_DOUT_WORDS_TDATA_in[19] = (S_AXIS_DOUT_WORDS_TDATA[19] !== 1'bz) && S_AXIS_DOUT_WORDS_TDATA[19]; // rv 0
  assign S_AXIS_DOUT_WORDS_TDATA_in[1] = (S_AXIS_DOUT_WORDS_TDATA[1] !== 1'bz) && S_AXIS_DOUT_WORDS_TDATA[1]; // rv 0
  assign S_AXIS_DOUT_WORDS_TDATA_in[20] = (S_AXIS_DOUT_WORDS_TDATA[20] !== 1'bz) && S_AXIS_DOUT_WORDS_TDATA[20]; // rv 0
  assign S_AXIS_DOUT_WORDS_TDATA_in[21] = (S_AXIS_DOUT_WORDS_TDATA[21] !== 1'bz) && S_AXIS_DOUT_WORDS_TDATA[21]; // rv 0
  assign S_AXIS_DOUT_WORDS_TDATA_in[22] = (S_AXIS_DOUT_WORDS_TDATA[22] !== 1'bz) && S_AXIS_DOUT_WORDS_TDATA[22]; // rv 0
  assign S_AXIS_DOUT_WORDS_TDATA_in[23] = (S_AXIS_DOUT_WORDS_TDATA[23] !== 1'bz) && S_AXIS_DOUT_WORDS_TDATA[23]; // rv 0
  assign S_AXIS_DOUT_WORDS_TDATA_in[24] = (S_AXIS_DOUT_WORDS_TDATA[24] !== 1'bz) && S_AXIS_DOUT_WORDS_TDATA[24]; // rv 0
  assign S_AXIS_DOUT_WORDS_TDATA_in[25] = (S_AXIS_DOUT_WORDS_TDATA[25] !== 1'bz) && S_AXIS_DOUT_WORDS_TDATA[25]; // rv 0
  assign S_AXIS_DOUT_WORDS_TDATA_in[26] = (S_AXIS_DOUT_WORDS_TDATA[26] !== 1'bz) && S_AXIS_DOUT_WORDS_TDATA[26]; // rv 0
  assign S_AXIS_DOUT_WORDS_TDATA_in[27] = (S_AXIS_DOUT_WORDS_TDATA[27] !== 1'bz) && S_AXIS_DOUT_WORDS_TDATA[27]; // rv 0
  assign S_AXIS_DOUT_WORDS_TDATA_in[28] = (S_AXIS_DOUT_WORDS_TDATA[28] !== 1'bz) && S_AXIS_DOUT_WORDS_TDATA[28]; // rv 0
  assign S_AXIS_DOUT_WORDS_TDATA_in[29] = (S_AXIS_DOUT_WORDS_TDATA[29] !== 1'bz) && S_AXIS_DOUT_WORDS_TDATA[29]; // rv 0
  assign S_AXIS_DOUT_WORDS_TDATA_in[2] = (S_AXIS_DOUT_WORDS_TDATA[2] !== 1'bz) && S_AXIS_DOUT_WORDS_TDATA[2]; // rv 0
  assign S_AXIS_DOUT_WORDS_TDATA_in[30] = (S_AXIS_DOUT_WORDS_TDATA[30] !== 1'bz) && S_AXIS_DOUT_WORDS_TDATA[30]; // rv 0
  assign S_AXIS_DOUT_WORDS_TDATA_in[31] = (S_AXIS_DOUT_WORDS_TDATA[31] !== 1'bz) && S_AXIS_DOUT_WORDS_TDATA[31]; // rv 0
  assign S_AXIS_DOUT_WORDS_TDATA_in[3] = (S_AXIS_DOUT_WORDS_TDATA[3] !== 1'bz) && S_AXIS_DOUT_WORDS_TDATA[3]; // rv 0
  assign S_AXIS_DOUT_WORDS_TDATA_in[4] = (S_AXIS_DOUT_WORDS_TDATA[4] !== 1'bz) && S_AXIS_DOUT_WORDS_TDATA[4]; // rv 0
  assign S_AXIS_DOUT_WORDS_TDATA_in[5] = (S_AXIS_DOUT_WORDS_TDATA[5] !== 1'bz) && S_AXIS_DOUT_WORDS_TDATA[5]; // rv 0
  assign S_AXIS_DOUT_WORDS_TDATA_in[6] = (S_AXIS_DOUT_WORDS_TDATA[6] !== 1'bz) && S_AXIS_DOUT_WORDS_TDATA[6]; // rv 0
  assign S_AXIS_DOUT_WORDS_TDATA_in[7] = (S_AXIS_DOUT_WORDS_TDATA[7] !== 1'bz) && S_AXIS_DOUT_WORDS_TDATA[7]; // rv 0
  assign S_AXIS_DOUT_WORDS_TDATA_in[8] = (S_AXIS_DOUT_WORDS_TDATA[8] !== 1'bz) && S_AXIS_DOUT_WORDS_TDATA[8]; // rv 0
  assign S_AXIS_DOUT_WORDS_TDATA_in[9] = (S_AXIS_DOUT_WORDS_TDATA[9] !== 1'bz) && S_AXIS_DOUT_WORDS_TDATA[9]; // rv 0
  assign S_AXIS_DOUT_WORDS_TLAST_in = (S_AXIS_DOUT_WORDS_TLAST !== 1'bz) && S_AXIS_DOUT_WORDS_TLAST; // rv 0
  assign S_AXIS_DOUT_WORDS_TVALID_in = (S_AXIS_DOUT_WORDS_TVALID !== 1'bz) && S_AXIS_DOUT_WORDS_TVALID; // rv 0
  assign S_AXI_ACLK_in = (S_AXI_ACLK !== 1'bz) && S_AXI_ACLK; // rv 0
  assign S_AXI_ARADDR_in[0] = (S_AXI_ARADDR[0] !== 1'bz) && S_AXI_ARADDR[0]; // rv 0
  assign S_AXI_ARADDR_in[10] = (S_AXI_ARADDR[10] !== 1'bz) && S_AXI_ARADDR[10]; // rv 0
  assign S_AXI_ARADDR_in[11] = (S_AXI_ARADDR[11] !== 1'bz) && S_AXI_ARADDR[11]; // rv 0
  assign S_AXI_ARADDR_in[12] = (S_AXI_ARADDR[12] !== 1'bz) && S_AXI_ARADDR[12]; // rv 0
  assign S_AXI_ARADDR_in[13] = (S_AXI_ARADDR[13] !== 1'bz) && S_AXI_ARADDR[13]; // rv 0
  assign S_AXI_ARADDR_in[14] = (S_AXI_ARADDR[14] !== 1'bz) && S_AXI_ARADDR[14]; // rv 0
  assign S_AXI_ARADDR_in[15] = (S_AXI_ARADDR[15] !== 1'bz) && S_AXI_ARADDR[15]; // rv 0
  assign S_AXI_ARADDR_in[16] = (S_AXI_ARADDR[16] !== 1'bz) && S_AXI_ARADDR[16]; // rv 0
  assign S_AXI_ARADDR_in[17] = (S_AXI_ARADDR[17] !== 1'bz) && S_AXI_ARADDR[17]; // rv 0
  assign S_AXI_ARADDR_in[1] = (S_AXI_ARADDR[1] !== 1'bz) && S_AXI_ARADDR[1]; // rv 0
  assign S_AXI_ARADDR_in[2] = (S_AXI_ARADDR[2] !== 1'bz) && S_AXI_ARADDR[2]; // rv 0
  assign S_AXI_ARADDR_in[3] = (S_AXI_ARADDR[3] !== 1'bz) && S_AXI_ARADDR[3]; // rv 0
  assign S_AXI_ARADDR_in[4] = (S_AXI_ARADDR[4] !== 1'bz) && S_AXI_ARADDR[4]; // rv 0
  assign S_AXI_ARADDR_in[5] = (S_AXI_ARADDR[5] !== 1'bz) && S_AXI_ARADDR[5]; // rv 0
  assign S_AXI_ARADDR_in[6] = (S_AXI_ARADDR[6] !== 1'bz) && S_AXI_ARADDR[6]; // rv 0
  assign S_AXI_ARADDR_in[7] = (S_AXI_ARADDR[7] !== 1'bz) && S_AXI_ARADDR[7]; // rv 0
  assign S_AXI_ARADDR_in[8] = (S_AXI_ARADDR[8] !== 1'bz) && S_AXI_ARADDR[8]; // rv 0
  assign S_AXI_ARADDR_in[9] = (S_AXI_ARADDR[9] !== 1'bz) && S_AXI_ARADDR[9]; // rv 0
  assign S_AXI_ARVALID_in = (S_AXI_ARVALID !== 1'bz) && S_AXI_ARVALID; // rv 0
  assign S_AXI_AWADDR_in[0] = (S_AXI_AWADDR[0] !== 1'bz) && S_AXI_AWADDR[0]; // rv 0
  assign S_AXI_AWADDR_in[10] = (S_AXI_AWADDR[10] !== 1'bz) && S_AXI_AWADDR[10]; // rv 0
  assign S_AXI_AWADDR_in[11] = (S_AXI_AWADDR[11] !== 1'bz) && S_AXI_AWADDR[11]; // rv 0
  assign S_AXI_AWADDR_in[12] = (S_AXI_AWADDR[12] !== 1'bz) && S_AXI_AWADDR[12]; // rv 0
  assign S_AXI_AWADDR_in[13] = (S_AXI_AWADDR[13] !== 1'bz) && S_AXI_AWADDR[13]; // rv 0
  assign S_AXI_AWADDR_in[14] = (S_AXI_AWADDR[14] !== 1'bz) && S_AXI_AWADDR[14]; // rv 0
  assign S_AXI_AWADDR_in[15] = (S_AXI_AWADDR[15] !== 1'bz) && S_AXI_AWADDR[15]; // rv 0
  assign S_AXI_AWADDR_in[16] = (S_AXI_AWADDR[16] !== 1'bz) && S_AXI_AWADDR[16]; // rv 0
  assign S_AXI_AWADDR_in[17] = (S_AXI_AWADDR[17] !== 1'bz) && S_AXI_AWADDR[17]; // rv 0
  assign S_AXI_AWADDR_in[1] = (S_AXI_AWADDR[1] !== 1'bz) && S_AXI_AWADDR[1]; // rv 0
  assign S_AXI_AWADDR_in[2] = (S_AXI_AWADDR[2] !== 1'bz) && S_AXI_AWADDR[2]; // rv 0
  assign S_AXI_AWADDR_in[3] = (S_AXI_AWADDR[3] !== 1'bz) && S_AXI_AWADDR[3]; // rv 0
  assign S_AXI_AWADDR_in[4] = (S_AXI_AWADDR[4] !== 1'bz) && S_AXI_AWADDR[4]; // rv 0
  assign S_AXI_AWADDR_in[5] = (S_AXI_AWADDR[5] !== 1'bz) && S_AXI_AWADDR[5]; // rv 0
  assign S_AXI_AWADDR_in[6] = (S_AXI_AWADDR[6] !== 1'bz) && S_AXI_AWADDR[6]; // rv 0
  assign S_AXI_AWADDR_in[7] = (S_AXI_AWADDR[7] !== 1'bz) && S_AXI_AWADDR[7]; // rv 0
  assign S_AXI_AWADDR_in[8] = (S_AXI_AWADDR[8] !== 1'bz) && S_AXI_AWADDR[8]; // rv 0
  assign S_AXI_AWADDR_in[9] = (S_AXI_AWADDR[9] !== 1'bz) && S_AXI_AWADDR[9]; // rv 0
  assign S_AXI_AWVALID_in = (S_AXI_AWVALID !== 1'bz) && S_AXI_AWVALID; // rv 0
  assign S_AXI_BREADY_in = (S_AXI_BREADY !== 1'bz) && S_AXI_BREADY; // rv 0
  assign S_AXI_RREADY_in = (S_AXI_RREADY !== 1'bz) && S_AXI_RREADY; // rv 0
  assign S_AXI_WDATA_in[0] = (S_AXI_WDATA[0] !== 1'bz) && S_AXI_WDATA[0]; // rv 0
  assign S_AXI_WDATA_in[10] = (S_AXI_WDATA[10] !== 1'bz) && S_AXI_WDATA[10]; // rv 0
  assign S_AXI_WDATA_in[11] = (S_AXI_WDATA[11] !== 1'bz) && S_AXI_WDATA[11]; // rv 0
  assign S_AXI_WDATA_in[12] = (S_AXI_WDATA[12] !== 1'bz) && S_AXI_WDATA[12]; // rv 0
  assign S_AXI_WDATA_in[13] = (S_AXI_WDATA[13] !== 1'bz) && S_AXI_WDATA[13]; // rv 0
  assign S_AXI_WDATA_in[14] = (S_AXI_WDATA[14] !== 1'bz) && S_AXI_WDATA[14]; // rv 0
  assign S_AXI_WDATA_in[15] = (S_AXI_WDATA[15] !== 1'bz) && S_AXI_WDATA[15]; // rv 0
  assign S_AXI_WDATA_in[16] = (S_AXI_WDATA[16] !== 1'bz) && S_AXI_WDATA[16]; // rv 0
  assign S_AXI_WDATA_in[17] = (S_AXI_WDATA[17] !== 1'bz) && S_AXI_WDATA[17]; // rv 0
  assign S_AXI_WDATA_in[18] = (S_AXI_WDATA[18] !== 1'bz) && S_AXI_WDATA[18]; // rv 0
  assign S_AXI_WDATA_in[19] = (S_AXI_WDATA[19] !== 1'bz) && S_AXI_WDATA[19]; // rv 0
  assign S_AXI_WDATA_in[1] = (S_AXI_WDATA[1] !== 1'bz) && S_AXI_WDATA[1]; // rv 0
  assign S_AXI_WDATA_in[20] = (S_AXI_WDATA[20] !== 1'bz) && S_AXI_WDATA[20]; // rv 0
  assign S_AXI_WDATA_in[21] = (S_AXI_WDATA[21] !== 1'bz) && S_AXI_WDATA[21]; // rv 0
  assign S_AXI_WDATA_in[22] = (S_AXI_WDATA[22] !== 1'bz) && S_AXI_WDATA[22]; // rv 0
  assign S_AXI_WDATA_in[23] = (S_AXI_WDATA[23] !== 1'bz) && S_AXI_WDATA[23]; // rv 0
  assign S_AXI_WDATA_in[24] = (S_AXI_WDATA[24] !== 1'bz) && S_AXI_WDATA[24]; // rv 0
  assign S_AXI_WDATA_in[25] = (S_AXI_WDATA[25] !== 1'bz) && S_AXI_WDATA[25]; // rv 0
  assign S_AXI_WDATA_in[26] = (S_AXI_WDATA[26] !== 1'bz) && S_AXI_WDATA[26]; // rv 0
  assign S_AXI_WDATA_in[27] = (S_AXI_WDATA[27] !== 1'bz) && S_AXI_WDATA[27]; // rv 0
  assign S_AXI_WDATA_in[28] = (S_AXI_WDATA[28] !== 1'bz) && S_AXI_WDATA[28]; // rv 0
  assign S_AXI_WDATA_in[29] = (S_AXI_WDATA[29] !== 1'bz) && S_AXI_WDATA[29]; // rv 0
  assign S_AXI_WDATA_in[2] = (S_AXI_WDATA[2] !== 1'bz) && S_AXI_WDATA[2]; // rv 0
  assign S_AXI_WDATA_in[30] = (S_AXI_WDATA[30] !== 1'bz) && S_AXI_WDATA[30]; // rv 0
  assign S_AXI_WDATA_in[31] = (S_AXI_WDATA[31] !== 1'bz) && S_AXI_WDATA[31]; // rv 0
  assign S_AXI_WDATA_in[3] = (S_AXI_WDATA[3] !== 1'bz) && S_AXI_WDATA[3]; // rv 0
  assign S_AXI_WDATA_in[4] = (S_AXI_WDATA[4] !== 1'bz) && S_AXI_WDATA[4]; // rv 0
  assign S_AXI_WDATA_in[5] = (S_AXI_WDATA[5] !== 1'bz) && S_AXI_WDATA[5]; // rv 0
  assign S_AXI_WDATA_in[6] = (S_AXI_WDATA[6] !== 1'bz) && S_AXI_WDATA[6]; // rv 0
  assign S_AXI_WDATA_in[7] = (S_AXI_WDATA[7] !== 1'bz) && S_AXI_WDATA[7]; // rv 0
  assign S_AXI_WDATA_in[8] = (S_AXI_WDATA[8] !== 1'bz) && S_AXI_WDATA[8]; // rv 0
  assign S_AXI_WDATA_in[9] = (S_AXI_WDATA[9] !== 1'bz) && S_AXI_WDATA[9]; // rv 0
  assign S_AXI_WVALID_in = (S_AXI_WVALID !== 1'bz) && S_AXI_WVALID; // rv 0
`endif
  assign DEBUG_CLK_EN_in = (DEBUG_CLK_EN !== 1'bz) && DEBUG_CLK_EN; // rv 0
  assign DEBUG_SEL_IN_in[0] = (DEBUG_SEL_IN[0] !== 1'bz) && DEBUG_SEL_IN[0]; // rv 0
  assign DEBUG_SEL_IN_in[1] = (DEBUG_SEL_IN[1] !== 1'bz) && DEBUG_SEL_IN[1]; // rv 0
  assign DEBUG_SEL_IN_in[2] = (DEBUG_SEL_IN[2] !== 1'bz) && DEBUG_SEL_IN[2]; // rv 0
  assign DEBUG_SEL_IN_in[3] = (DEBUG_SEL_IN[3] !== 1'bz) && DEBUG_SEL_IN[3]; // rv 0
  assign RESET_N_in = (RESET_N === 1'bz) || RESET_N; // rv 1
  assign SPARE_IN_in[0] = (SPARE_IN[0] !== 1'bz) && SPARE_IN[0]; // rv 0
  assign SPARE_IN_in[10] = (SPARE_IN[10] !== 1'bz) && SPARE_IN[10]; // rv 0
  assign SPARE_IN_in[11] = (SPARE_IN[11] !== 1'bz) && SPARE_IN[11]; // rv 0
  assign SPARE_IN_in[12] = (SPARE_IN[12] !== 1'bz) && SPARE_IN[12]; // rv 0
  assign SPARE_IN_in[13] = (SPARE_IN[13] !== 1'bz) && SPARE_IN[13]; // rv 0
  assign SPARE_IN_in[14] = (SPARE_IN[14] !== 1'bz) && SPARE_IN[14]; // rv 0
  assign SPARE_IN_in[15] = (SPARE_IN[15] !== 1'bz) && SPARE_IN[15]; // rv 0
  assign SPARE_IN_in[1] = (SPARE_IN[1] !== 1'bz) && SPARE_IN[1]; // rv 0
  assign SPARE_IN_in[2] = (SPARE_IN[2] !== 1'bz) && SPARE_IN[2]; // rv 0
  assign SPARE_IN_in[3] = (SPARE_IN[3] !== 1'bz) && SPARE_IN[3]; // rv 0
  assign SPARE_IN_in[4] = (SPARE_IN[4] !== 1'bz) && SPARE_IN[4]; // rv 0
  assign SPARE_IN_in[5] = (SPARE_IN[5] !== 1'bz) && SPARE_IN[5]; // rv 0
  assign SPARE_IN_in[6] = (SPARE_IN[6] !== 1'bz) && SPARE_IN[6]; // rv 0
  assign SPARE_IN_in[7] = (SPARE_IN[7] !== 1'bz) && SPARE_IN[7]; // rv 0
  assign SPARE_IN_in[8] = (SPARE_IN[8] !== 1'bz) && SPARE_IN[8]; // rv 0
  assign SPARE_IN_in[9] = (SPARE_IN[9] !== 1'bz) && SPARE_IN[9]; // rv 0
`ifndef XIL_XECLIB
  reg attr_test;
  reg attr_err;
  initial begin
  trig_attr = 1'b0;
  `ifdef XIL_ATTR_TEST
    attr_test = 1'b1;
  `else
    attr_test = 1'b0;
  `endif
    attr_err = 1'b0;
    #1;
    trig_attr = ~trig_attr;
  end
`endif
`ifdef XIL_XECLIB
  assign PHYSICAL_UTILIZATION_BIN = PHYSICAL_UTILIZATION_REG * 1000;
  assign THROUGHPUT_UTILIZATION_BIN = THROUGHPUT_UTILIZATION_REG * 1000;
`else
  always @ (trig_attr) begin
  #1;
  PHYSICAL_UTILIZATION_BIN = PHYSICAL_UTILIZATION_REG * 1000;
  THROUGHPUT_UTILIZATION_BIN = THROUGHPUT_UTILIZATION_REG * 1000;
  end
`endif
`ifndef XIL_XECLIB
always @ (trig_attr) begin
  #1;
  if ((attr_test == 1'b1) ||
        ((MODE_REG != "TURBO_DECODE") &&
         (MODE_REG != "LDPC_DECODE") &&
         (MODE_REG != "LDPC_ENCODE"))) begin
      $display("Error: [Unisim %s-101] MODE attribute is set to %s.  Legal values for this attribute are TURBO_DECODE, LDPC_DECODE or LDPC_ENCODE. Instance: %m", MODULE_NAME, MODE_REG);
    attr_err = 1'b1;
  end
  if ((attr_test == 1'b1) ||
        (PHYSICAL_UTILIZATION_REG < 0.00 || PHYSICAL_UTILIZATION_REG > 100.00)) begin
      $display("Error: [Unisim %s-102] PHYSICAL_UTILIZATION attribute is set to %f.  Legal values for this attribute are 0.00 to 100.00. Instance: %m", MODULE_NAME, PHYSICAL_UTILIZATION_REG);
    attr_err = 1'b1;
  end
  if ((attr_test == 1'b1) ||
      ((SIM_DEVICE_REG != "ULTRASCALE_PLUS") &&
       (SIM_DEVICE_REG != "ULTRASCALE_PLUS_ES1") &&
       (SIM_DEVICE_REG != "ULTRASCALE_PLUS_ES2"))) begin
    $display("Error: [Unisim %s-103] SIM_DEVICE attribute is set to %s.  Legal values for this attribute are ULTRASCALE_PLUS, ULTRASCALE_PLUS_ES1 or ULTRASCALE_PLUS_ES2. Instance: %m", MODULE_NAME, SIM_DEVICE_REG);
    attr_err = 1'b1;
  end
  if ((attr_test == 1'b1) ||
        ((STANDARD_REG != "LTE") &&
         (STANDARD_REG != "5G") &&
         (STANDARD_REG != "CUSTOM") &&
         (STANDARD_REG != "DOCSIS") &&
         (STANDARD_REG != "WIFI"))) begin
      $display("Error: [Unisim %s-104] STANDARD attribute is set to %s.  Legal values for this attribute are LTE, 5G, CUSTOM, DOCSIS or WIFI. Instance: %m", MODULE_NAME, STANDARD_REG);
      attr_err = 1'b1;
    end
    if ((attr_test == 1'b1) ||
        (THROUGHPUT_UTILIZATION_REG < 0.00 || THROUGHPUT_UTILIZATION_REG > 100.00)) begin
      $display("Error: [Unisim %s-105] THROUGHPUT_UTILIZATION attribute is set to %f.  Legal values for this attribute are 0.00 to 100.00. Instance: %m", MODULE_NAME, THROUGHPUT_UTILIZATION_REG);
    attr_err = 1'b1;
  end
  if (attr_err == 1'b1) #1 $finish;
end
`endif
assign MBIST_TCK_in = 1'b1; // tie off
assign SCAN_CLK_in = 1'b1; // tie off
assign XIL_UNCONN_CLK_in = 470'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111; // tie off
assign CSSD_CLK_STOP_EVENT_in = 4'b1111; // tie off
assign CSSD_RST_N_in = 1'b1; // tie off
assign CTL_CSSD_EN_N_in = 1'b1; // tie off
assign CTL_CSSD_MRKR_START_INIT_in = 16'b1111111111111111; // tie off
assign CTL_CSSD_MRKR_STOP_INIT_in = 16'b1111111111111111; // tie off
assign CTL_CSSD_ROOT_CLK_DIS_in = 8'b11111111; // tie off
assign CTL_CSSD_ROOT_CLK_SEL_in = 3'b111; // tie off
assign CTL_CSSD_SNGL_CHAIN_MD_N_in = 1'b1; // tie off
assign CTL_CSSD_STOP_COUNT_in = 48'b111111111111111111111111111111111111111111111111; // tie off
assign DFTRAM_BYPASS_N_in = 1'b1; // tie off
assign MBIST_TDI_in = 1'b1; // tie off
assign MBIST_TMS_in = 1'b1; // tie off
assign MBIST_TRST_in = 1'b1; // tie off
assign SCANENABLE_N_in = 1'b1; // tie off
assign SCANIN_in = 200'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111; // tie off
assign SCANMODE_N_in = 1'b1; // tie off
assign TEST_MODE_PIN_CHAR_N_in = 1'b1; // tie off
assign XIL_UNCONN_IN_in = 1862'b11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111; // tie off
SIP_FE SIP_FE_INST (
.CSSD_CLK_STOP_DONE (CSSD_CLK_STOP_DONE_out),
.DEBUG_DOUT (DEBUG_DOUT_out),
.DEBUG_PHASE (DEBUG_PHASE_out),
.INTERRUPT (INTERRUPT_out),
.MBIST_COMPSTAT (MBIST_COMPSTAT_out),
.MBIST_TDO (MBIST_TDO_out),
.M_AXIS_DOUT_TDATA (M_AXIS_DOUT_TDATA_out),
.M_AXIS_DOUT_TLAST (M_AXIS_DOUT_TLAST_out),
.M_AXIS_DOUT_TVALID (M_AXIS_DOUT_TVALID_out),
.M_AXIS_STATUS_TDATA (M_AXIS_STATUS_TDATA_out),
.M_AXIS_STATUS_TVALID (M_AXIS_STATUS_TVALID_out),
.SCANOUT (SCANOUT_out),
.SPARE_OUT (SPARE_OUT_out),
.S_AXIS_CTRL_TREADY (S_AXIS_CTRL_TREADY_out),
.S_AXIS_DIN_TREADY (S_AXIS_DIN_TREADY_out),
.S_AXIS_DIN_WORDS_TREADY (S_AXIS_DIN_WORDS_TREADY_out),
.S_AXIS_DOUT_WORDS_TREADY (S_AXIS_DOUT_WORDS_TREADY_out),
.S_AXI_ARREADY (S_AXI_ARREADY_out),
.S_AXI_AWREADY (S_AXI_AWREADY_out),
.S_AXI_BVALID (S_AXI_BVALID_out),
.S_AXI_RDATA (S_AXI_RDATA_out),
.S_AXI_RVALID (S_AXI_RVALID_out),
.S_AXI_WREADY (S_AXI_WREADY_out),
.XIL_UNCONN_OUT (XIL_UNCONN_OUT_out),
.CORE_CLK (CORE_CLK_in),
.CSSD_CLK_STOP_EVENT (CSSD_CLK_STOP_EVENT_in),
.CSSD_RST_N (CSSD_RST_N_in),
.CTL_CSSD_EN_N (CTL_CSSD_EN_N_in),
.CTL_CSSD_MRKR_START_INIT (CTL_CSSD_MRKR_START_INIT_in),
.CTL_CSSD_MRKR_STOP_INIT (CTL_CSSD_MRKR_STOP_INIT_in),
.CTL_CSSD_ROOT_CLK_DIS (CTL_CSSD_ROOT_CLK_DIS_in),
.CTL_CSSD_ROOT_CLK_SEL (CTL_CSSD_ROOT_CLK_SEL_in),
.CTL_CSSD_SNGL_CHAIN_MD_N (CTL_CSSD_SNGL_CHAIN_MD_N_in),
.CTL_CSSD_STOP_COUNT (CTL_CSSD_STOP_COUNT_in),
.DEBUG_CLK_EN (DEBUG_CLK_EN_in),
.DEBUG_EN (DEBUG_EN_in),
.DEBUG_SEL_IN (DEBUG_SEL_IN_in),
.DFTRAM_BYPASS_N (DFTRAM_BYPASS_N_in),
.MBIST_TCK (MBIST_TCK_in),
.MBIST_TDI (MBIST_TDI_in),
.MBIST_TMS (MBIST_TMS_in),
.MBIST_TRST (MBIST_TRST_in),
.M_AXIS_DOUT_ACLK (M_AXIS_DOUT_ACLK_in),
.M_AXIS_DOUT_TREADY (M_AXIS_DOUT_TREADY_in),
.M_AXIS_STATUS_ACLK (M_AXIS_STATUS_ACLK_in),
.M_AXIS_STATUS_TREADY (M_AXIS_STATUS_TREADY_in),
.RESET_N (RESET_N_in),
.SCANENABLE_N (SCANENABLE_N_in),
.SCANIN (SCANIN_in),
.SCANMODE_N (SCANMODE_N_in),
.SCAN_CLK (SCAN_CLK_in),
.SPARE_IN (SPARE_IN_in),
.S_AXIS_CTRL_ACLK (S_AXIS_CTRL_ACLK_in),
.S_AXIS_CTRL_TDATA (S_AXIS_CTRL_TDATA_in),
.S_AXIS_CTRL_TVALID (S_AXIS_CTRL_TVALID_in),
.S_AXIS_DIN_ACLK (S_AXIS_DIN_ACLK_in),
.S_AXIS_DIN_TDATA (S_AXIS_DIN_TDATA_in),
.S_AXIS_DIN_TLAST (S_AXIS_DIN_TLAST_in),
.S_AXIS_DIN_TVALID (S_AXIS_DIN_TVALID_in),
.S_AXIS_DIN_WORDS_ACLK (S_AXIS_DIN_WORDS_ACLK_in),
.S_AXIS_DIN_WORDS_TDATA (S_AXIS_DIN_WORDS_TDATA_in),
.S_AXIS_DIN_WORDS_TLAST (S_AXIS_DIN_WORDS_TLAST_in),
.S_AXIS_DIN_WORDS_TVALID (S_AXIS_DIN_WORDS_TVALID_in),
.S_AXIS_DOUT_WORDS_ACLK (S_AXIS_DOUT_WORDS_ACLK_in),
.S_AXIS_DOUT_WORDS_TDATA (S_AXIS_DOUT_WORDS_TDATA_in),
.S_AXIS_DOUT_WORDS_TLAST (S_AXIS_DOUT_WORDS_TLAST_in),
.S_AXIS_DOUT_WORDS_TVALID (S_AXIS_DOUT_WORDS_TVALID_in),
.S_AXI_ACLK (S_AXI_ACLK_in),
.S_AXI_ARADDR (S_AXI_ARADDR_in),
.S_AXI_ARVALID (S_AXI_ARVALID_in),
.S_AXI_AWADDR (S_AXI_AWADDR_in),
.S_AXI_AWVALID (S_AXI_AWVALID_in),
.S_AXI_BREADY (S_AXI_BREADY_in),
.S_AXI_RREADY (S_AXI_RREADY_in),
.S_AXI_WDATA (S_AXI_WDATA_in),
.S_AXI_WVALID (S_AXI_WVALID_in),
.TEST_MODE_PIN_CHAR_N (TEST_MODE_PIN_CHAR_N_in),
.XIL_UNCONN_CLK (XIL_UNCONN_CLK_in),
.XIL_UNCONN_IN (XIL_UNCONN_IN_in),
.GSR (glblGSR)
);
`ifdef XIL_TIMING
  reg notifier;
`endif
`ifndef XIL_XECLIB
  specify
    (CORE_CLK => DEBUG_DOUT[0]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[100]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[101]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[102]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[103]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[104]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[105]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[106]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[107]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[108]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[109]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[10]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[110]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[111]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[112]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[113]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[114]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[115]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[116]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[117]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[118]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[119]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[11]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[120]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[121]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[122]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[123]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[124]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[125]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[126]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[127]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[128]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[129]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[12]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[130]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[131]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[132]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[133]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[134]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[135]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[136]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[137]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[138]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[139]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[13]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[140]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[141]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[142]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[143]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[144]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[145]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[146]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[147]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[148]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[149]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[14]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[150]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[151]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[152]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[153]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[154]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[155]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[156]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[157]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[158]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[159]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[15]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[160]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[161]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[162]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[163]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[164]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[165]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[166]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[167]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[168]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[169]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[16]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[170]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[171]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[172]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[173]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[174]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[175]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[176]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[177]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[178]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[179]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[17]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[180]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[181]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[182]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[183]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[184]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[185]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[186]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[187]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[188]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[189]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[18]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[190]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[191]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[192]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[193]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[194]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[195]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[196]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[197]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[198]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[199]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[19]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[1]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[200]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[201]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[202]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[203]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[204]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[205]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[206]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[207]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[208]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[209]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[20]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[210]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[211]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[212]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[213]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[214]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[215]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[216]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[217]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[218]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[219]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[21]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[220]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[221]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[222]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[223]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[224]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[225]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[226]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[227]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[228]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[229]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[22]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[230]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[231]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[232]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[233]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[234]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[235]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[236]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[237]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[238]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[239]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[23]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[240]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[241]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[242]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[243]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[244]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[245]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[246]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[247]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[248]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[249]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[24]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[250]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[251]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[252]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[253]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[254]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[255]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[256]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[257]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[258]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[259]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[25]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[260]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[261]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[262]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[263]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[264]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[265]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[266]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[267]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[268]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[269]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[26]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[270]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[271]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[272]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[273]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[274]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[275]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[276]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[277]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[278]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[279]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[27]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[280]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[281]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[282]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[283]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[284]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[285]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[286]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[287]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[288]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[289]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[28]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[290]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[291]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[292]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[293]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[294]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[295]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[296]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[297]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[298]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[299]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[29]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[2]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[300]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[301]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[302]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[303]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[304]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[305]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[306]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[307]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[308]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[309]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[30]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[310]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[311]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[312]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[313]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[314]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[315]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[316]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[317]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[318]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[319]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[31]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[320]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[321]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[322]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[323]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[324]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[325]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[326]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[327]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[328]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[329]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[32]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[330]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[331]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[332]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[333]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[334]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[335]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[336]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[337]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[338]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[339]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[33]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[340]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[341]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[342]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[343]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[344]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[345]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[346]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[347]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[348]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[349]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[34]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[350]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[351]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[352]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[353]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[354]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[355]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[356]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[357]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[358]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[359]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[35]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[360]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[361]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[362]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[363]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[364]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[365]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[366]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[367]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[368]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[369]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[36]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[370]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[371]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[372]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[373]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[374]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[375]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[376]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[377]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[378]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[379]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[37]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[380]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[381]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[382]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[383]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[384]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[385]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[386]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[387]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[388]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[389]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[38]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[390]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[391]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[392]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[393]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[394]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[395]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[396]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[397]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[398]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[399]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[39]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[3]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[40]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[41]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[42]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[43]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[44]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[45]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[46]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[47]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[48]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[49]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[4]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[50]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[51]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[52]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[53]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[54]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[55]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[56]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[57]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[58]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[59]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[5]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[60]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[61]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[62]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[63]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[64]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[65]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[66]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[67]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[68]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[69]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[6]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[70]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[71]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[72]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[73]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[74]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[75]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[76]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[77]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[78]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[79]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[7]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[80]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[81]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[82]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[83]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[84]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[85]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[86]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[87]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[88]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[89]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[8]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[90]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[91]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[92]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[93]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[94]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[95]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[96]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[97]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[98]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[99]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_DOUT[9]) = (100:100:100, 100:100:100);
    (CORE_CLK => DEBUG_PHASE) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[0]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[100]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[101]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[102]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[103]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[104]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[105]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[106]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[107]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[108]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[109]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[10]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[110]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[111]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[112]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[113]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[114]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[115]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[116]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[117]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[118]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[119]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[11]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[120]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[121]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[122]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[123]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[124]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[125]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[126]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[127]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[128]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[129]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[12]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[130]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[131]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[132]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[133]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[134]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[135]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[136]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[137]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[138]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[139]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[13]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[140]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[141]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[142]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[143]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[144]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[145]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[146]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[147]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[148]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[149]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[14]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[150]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[151]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[152]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[153]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[154]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[155]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[156]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[157]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[158]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[159]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[15]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[160]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[161]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[162]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[163]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[164]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[165]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[166]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[167]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[168]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[169]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[16]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[170]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[171]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[172]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[173]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[174]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[175]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[176]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[177]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[178]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[179]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[17]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[180]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[181]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[182]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[183]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[184]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[185]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[186]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[187]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[188]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[189]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[18]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[190]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[191]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[192]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[193]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[194]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[195]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[196]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[197]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[198]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[199]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[19]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[1]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[200]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[201]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[202]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[203]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[204]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[205]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[206]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[207]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[208]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[209]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[20]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[210]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[211]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[212]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[213]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[214]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[215]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[216]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[217]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[218]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[219]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[21]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[220]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[221]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[222]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[223]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[224]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[225]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[226]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[227]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[228]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[229]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[22]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[230]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[231]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[232]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[233]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[234]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[235]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[236]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[237]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[238]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[239]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[23]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[240]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[241]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[242]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[243]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[244]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[245]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[246]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[247]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[248]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[249]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[24]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[250]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[251]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[252]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[253]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[254]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[255]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[256]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[257]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[258]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[259]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[25]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[260]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[261]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[262]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[263]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[264]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[265]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[266]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[267]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[268]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[269]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[26]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[270]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[271]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[272]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[273]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[274]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[275]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[276]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[277]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[278]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[279]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[27]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[280]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[281]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[282]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[283]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[284]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[285]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[286]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[287]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[288]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[289]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[28]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[290]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[291]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[292]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[293]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[294]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[295]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[296]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[297]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[298]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[299]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[29]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[2]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[300]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[301]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[302]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[303]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[304]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[305]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[306]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[307]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[308]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[309]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[30]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[310]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[311]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[312]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[313]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[314]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[315]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[316]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[317]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[318]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[319]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[31]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[320]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[321]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[322]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[323]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[324]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[325]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[326]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[327]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[328]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[329]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[32]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[330]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[331]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[332]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[333]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[334]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[335]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[336]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[337]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[338]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[339]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[33]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[340]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[341]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[342]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[343]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[344]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[345]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[346]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[347]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[348]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[349]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[34]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[350]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[351]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[352]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[353]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[354]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[355]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[356]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[357]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[358]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[359]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[35]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[360]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[361]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[362]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[363]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[364]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[365]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[366]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[367]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[368]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[369]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[36]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[370]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[371]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[372]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[373]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[374]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[375]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[376]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[377]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[378]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[379]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[37]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[380]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[381]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[382]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[383]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[384]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[385]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[386]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[387]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[388]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[389]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[38]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[390]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[391]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[392]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[393]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[394]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[395]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[396]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[397]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[398]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[399]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[39]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[3]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[400]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[401]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[402]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[403]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[404]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[405]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[406]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[407]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[408]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[409]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[40]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[410]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[411]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[412]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[413]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[414]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[415]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[416]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[417]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[418]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[419]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[41]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[420]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[421]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[422]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[423]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[424]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[425]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[426]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[427]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[428]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[429]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[42]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[430]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[431]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[432]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[433]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[434]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[435]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[436]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[437]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[438]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[439]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[43]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[440]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[441]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[442]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[443]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[444]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[445]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[446]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[447]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[448]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[449]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[44]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[450]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[451]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[452]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[453]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[454]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[455]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[456]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[457]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[458]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[459]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[45]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[460]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[461]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[462]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[463]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[464]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[465]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[466]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[467]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[468]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[469]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[46]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[470]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[471]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[472]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[473]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[474]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[475]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[476]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[477]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[478]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[479]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[47]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[480]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[481]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[482]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[483]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[484]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[485]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[486]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[487]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[488]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[489]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[48]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[490]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[491]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[492]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[493]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[494]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[495]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[496]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[497]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[498]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[499]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[49]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[4]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[500]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[501]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[502]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[503]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[504]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[505]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[506]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[507]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[508]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[509]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[50]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[510]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[511]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[51]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[52]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[53]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[54]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[55]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[56]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[57]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[58]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[59]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[5]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[60]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[61]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[62]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[63]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[64]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[65]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[66]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[67]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[68]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[69]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[6]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[70]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[71]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[72]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[73]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[74]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[75]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[76]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[77]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[78]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[79]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[7]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[80]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[81]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[82]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[83]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[84]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[85]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[86]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[87]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[88]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[89]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[8]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[90]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[91]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[92]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[93]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[94]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[95]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[96]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[97]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[98]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[99]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TDATA[9]) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TLAST) = (100:100:100, 100:100:100);
    (M_AXIS_DOUT_ACLK => M_AXIS_DOUT_TVALID) = (100:100:100, 100:100:100);
    (M_AXIS_STATUS_ACLK => M_AXIS_STATUS_TDATA[0]) = (100:100:100, 100:100:100);
    (M_AXIS_STATUS_ACLK => M_AXIS_STATUS_TDATA[10]) = (100:100:100, 100:100:100);
    (M_AXIS_STATUS_ACLK => M_AXIS_STATUS_TDATA[11]) = (100:100:100, 100:100:100);
    (M_AXIS_STATUS_ACLK => M_AXIS_STATUS_TDATA[12]) = (100:100:100, 100:100:100);
    (M_AXIS_STATUS_ACLK => M_AXIS_STATUS_TDATA[13]) = (100:100:100, 100:100:100);
    (M_AXIS_STATUS_ACLK => M_AXIS_STATUS_TDATA[14]) = (100:100:100, 100:100:100);
    (M_AXIS_STATUS_ACLK => M_AXIS_STATUS_TDATA[15]) = (100:100:100, 100:100:100);
    (M_AXIS_STATUS_ACLK => M_AXIS_STATUS_TDATA[16]) = (100:100:100, 100:100:100);
    (M_AXIS_STATUS_ACLK => M_AXIS_STATUS_TDATA[17]) = (100:100:100, 100:100:100);
    (M_AXIS_STATUS_ACLK => M_AXIS_STATUS_TDATA[18]) = (100:100:100, 100:100:100);
    (M_AXIS_STATUS_ACLK => M_AXIS_STATUS_TDATA[19]) = (100:100:100, 100:100:100);
    (M_AXIS_STATUS_ACLK => M_AXIS_STATUS_TDATA[1]) = (100:100:100, 100:100:100);
    (M_AXIS_STATUS_ACLK => M_AXIS_STATUS_TDATA[20]) = (100:100:100, 100:100:100);
    (M_AXIS_STATUS_ACLK => M_AXIS_STATUS_TDATA[21]) = (100:100:100, 100:100:100);
    (M_AXIS_STATUS_ACLK => M_AXIS_STATUS_TDATA[22]) = (100:100:100, 100:100:100);
    (M_AXIS_STATUS_ACLK => M_AXIS_STATUS_TDATA[23]) = (100:100:100, 100:100:100);
    (M_AXIS_STATUS_ACLK => M_AXIS_STATUS_TDATA[24]) = (100:100:100, 100:100:100);
    (M_AXIS_STATUS_ACLK => M_AXIS_STATUS_TDATA[25]) = (100:100:100, 100:100:100);
    (M_AXIS_STATUS_ACLK => M_AXIS_STATUS_TDATA[26]) = (100:100:100, 100:100:100);
    (M_AXIS_STATUS_ACLK => M_AXIS_STATUS_TDATA[27]) = (100:100:100, 100:100:100);
    (M_AXIS_STATUS_ACLK => M_AXIS_STATUS_TDATA[28]) = (100:100:100, 100:100:100);
    (M_AXIS_STATUS_ACLK => M_AXIS_STATUS_TDATA[29]) = (100:100:100, 100:100:100);
    (M_AXIS_STATUS_ACLK => M_AXIS_STATUS_TDATA[2]) = (100:100:100, 100:100:100);
    (M_AXIS_STATUS_ACLK => M_AXIS_STATUS_TDATA[30]) = (100:100:100, 100:100:100);
    (M_AXIS_STATUS_ACLK => M_AXIS_STATUS_TDATA[31]) = (100:100:100, 100:100:100);
    (M_AXIS_STATUS_ACLK => M_AXIS_STATUS_TDATA[3]) = (100:100:100, 100:100:100);
    (M_AXIS_STATUS_ACLK => M_AXIS_STATUS_TDATA[4]) = (100:100:100, 100:100:100);
    (M_AXIS_STATUS_ACLK => M_AXIS_STATUS_TDATA[5]) = (100:100:100, 100:100:100);
    (M_AXIS_STATUS_ACLK => M_AXIS_STATUS_TDATA[6]) = (100:100:100, 100:100:100);
    (M_AXIS_STATUS_ACLK => M_AXIS_STATUS_TDATA[7]) = (100:100:100, 100:100:100);
    (M_AXIS_STATUS_ACLK => M_AXIS_STATUS_TDATA[8]) = (100:100:100, 100:100:100);
    (M_AXIS_STATUS_ACLK => M_AXIS_STATUS_TDATA[9]) = (100:100:100, 100:100:100);
    (M_AXIS_STATUS_ACLK => M_AXIS_STATUS_TVALID) = (100:100:100, 100:100:100);
    (S_AXIS_CTRL_ACLK => S_AXIS_CTRL_TREADY) = (100:100:100, 100:100:100);
    (S_AXIS_DIN_ACLK => S_AXIS_DIN_TREADY) = (100:100:100, 100:100:100);
    (S_AXIS_DIN_WORDS_ACLK => S_AXIS_DIN_WORDS_TREADY) = (100:100:100, 100:100:100);
    (S_AXIS_DOUT_WORDS_ACLK => S_AXIS_DOUT_WORDS_TREADY) = (100:100:100, 100:100:100);
    (S_AXI_ACLK => INTERRUPT) = (100:100:100, 100:100:100);
    (S_AXI_ACLK => S_AXI_ARREADY) = (100:100:100, 100:100:100);
    (S_AXI_ACLK => S_AXI_AWREADY) = (100:100:100, 100:100:100);
    (S_AXI_ACLK => S_AXI_BVALID) = (100:100:100, 100:100:100);
    (S_AXI_ACLK => S_AXI_RDATA[0]) = (100:100:100, 100:100:100);
    (S_AXI_ACLK => S_AXI_RDATA[10]) = (100:100:100, 100:100:100);
    (S_AXI_ACLK => S_AXI_RDATA[11]) = (100:100:100, 100:100:100);
    (S_AXI_ACLK => S_AXI_RDATA[12]) = (100:100:100, 100:100:100);
    (S_AXI_ACLK => S_AXI_RDATA[13]) = (100:100:100, 100:100:100);
    (S_AXI_ACLK => S_AXI_RDATA[14]) = (100:100:100, 100:100:100);
    (S_AXI_ACLK => S_AXI_RDATA[15]) = (100:100:100, 100:100:100);
    (S_AXI_ACLK => S_AXI_RDATA[16]) = (100:100:100, 100:100:100);
    (S_AXI_ACLK => S_AXI_RDATA[17]) = (100:100:100, 100:100:100);
    (S_AXI_ACLK => S_AXI_RDATA[18]) = (100:100:100, 100:100:100);
    (S_AXI_ACLK => S_AXI_RDATA[19]) = (100:100:100, 100:100:100);
    (S_AXI_ACLK => S_AXI_RDATA[1]) = (100:100:100, 100:100:100);
    (S_AXI_ACLK => S_AXI_RDATA[20]) = (100:100:100, 100:100:100);
    (S_AXI_ACLK => S_AXI_RDATA[21]) = (100:100:100, 100:100:100);
    (S_AXI_ACLK => S_AXI_RDATA[22]) = (100:100:100, 100:100:100);
    (S_AXI_ACLK => S_AXI_RDATA[23]) = (100:100:100, 100:100:100);
    (S_AXI_ACLK => S_AXI_RDATA[24]) = (100:100:100, 100:100:100);
    (S_AXI_ACLK => S_AXI_RDATA[25]) = (100:100:100, 100:100:100);
    (S_AXI_ACLK => S_AXI_RDATA[26]) = (100:100:100, 100:100:100);
    (S_AXI_ACLK => S_AXI_RDATA[27]) = (100:100:100, 100:100:100);
    (S_AXI_ACLK => S_AXI_RDATA[28]) = (100:100:100, 100:100:100);
    (S_AXI_ACLK => S_AXI_RDATA[29]) = (100:100:100, 100:100:100);
    (S_AXI_ACLK => S_AXI_RDATA[2]) = (100:100:100, 100:100:100);
    (S_AXI_ACLK => S_AXI_RDATA[30]) = (100:100:100, 100:100:100);
    (S_AXI_ACLK => S_AXI_RDATA[31]) = (100:100:100, 100:100:100);
    (S_AXI_ACLK => S_AXI_RDATA[3]) = (100:100:100, 100:100:100);
    (S_AXI_ACLK => S_AXI_RDATA[4]) = (100:100:100, 100:100:100);
    (S_AXI_ACLK => S_AXI_RDATA[5]) = (100:100:100, 100:100:100);
    (S_AXI_ACLK => S_AXI_RDATA[6]) = (100:100:100, 100:100:100);
    (S_AXI_ACLK => S_AXI_RDATA[7]) = (100:100:100, 100:100:100);
    (S_AXI_ACLK => S_AXI_RDATA[8]) = (100:100:100, 100:100:100);
    (S_AXI_ACLK => S_AXI_RDATA[9]) = (100:100:100, 100:100:100);
    (S_AXI_ACLK => S_AXI_RVALID) = (100:100:100, 100:100:100);
    (S_AXI_ACLK => S_AXI_WREADY) = (100:100:100, 100:100:100);
`ifdef XIL_TIMING
    $period (negedge CORE_CLK, 0:0:0, notifier);
    $period (negedge M_AXIS_DOUT_ACLK, 0:0:0, notifier);
    $period (negedge M_AXIS_STATUS_ACLK, 0:0:0, notifier);
    $period (negedge S_AXIS_CTRL_ACLK, 0:0:0, notifier);
    $period (negedge S_AXIS_DIN_ACLK, 0:0:0, notifier);
    $period (negedge S_AXIS_DIN_WORDS_ACLK, 0:0:0, notifier);
    $period (negedge S_AXIS_DOUT_WORDS_ACLK, 0:0:0, notifier);
    $period (negedge S_AXI_ACLK, 0:0:0, notifier);
    $period (posedge CORE_CLK, 0:0:0, notifier);
    $period (posedge M_AXIS_DOUT_ACLK, 0:0:0, notifier);
    $period (posedge M_AXIS_STATUS_ACLK, 0:0:0, notifier);
    $period (posedge S_AXIS_CTRL_ACLK, 0:0:0, notifier);
    $period (posedge S_AXIS_DIN_ACLK, 0:0:0, notifier);
    $period (posedge S_AXIS_DIN_WORDS_ACLK, 0:0:0, notifier);
    $period (posedge S_AXIS_DOUT_WORDS_ACLK, 0:0:0, notifier);
    $period (posedge S_AXI_ACLK, 0:0:0, notifier);
    $setuphold (posedge CORE_CLK, negedge DEBUG_EN, 0:0:0, 0:0:0, notifier, , , CORE_CLK_delay, DEBUG_EN_delay);
    $setuphold (posedge CORE_CLK, posedge DEBUG_EN, 0:0:0, 0:0:0, notifier, , , CORE_CLK_delay, DEBUG_EN_delay);
    $setuphold (posedge M_AXIS_DOUT_ACLK, negedge M_AXIS_DOUT_TREADY, 0:0:0, 0:0:0, notifier, , , M_AXIS_DOUT_ACLK_delay, M_AXIS_DOUT_TREADY_delay);
    $setuphold (posedge M_AXIS_DOUT_ACLK, posedge M_AXIS_DOUT_TREADY, 0:0:0, 0:0:0, notifier, , , M_AXIS_DOUT_ACLK_delay, M_AXIS_DOUT_TREADY_delay);
    $setuphold (posedge M_AXIS_STATUS_ACLK, negedge M_AXIS_STATUS_TREADY, 0:0:0, 0:0:0, notifier, , , M_AXIS_STATUS_ACLK_delay, M_AXIS_STATUS_TREADY_delay);
    $setuphold (posedge M_AXIS_STATUS_ACLK, posedge M_AXIS_STATUS_TREADY, 0:0:0, 0:0:0, notifier, , , M_AXIS_STATUS_ACLK_delay, M_AXIS_STATUS_TREADY_delay);
    $setuphold (posedge S_AXIS_CTRL_ACLK, negedge S_AXIS_CTRL_TDATA[0], 0:0:0, 0:0:0, notifier, , , S_AXIS_CTRL_ACLK_delay, S_AXIS_CTRL_TDATA_delay[0]);
    $setuphold (posedge S_AXIS_CTRL_ACLK, negedge S_AXIS_CTRL_TDATA[10], 0:0:0, 0:0:0, notifier, , , S_AXIS_CTRL_ACLK_delay, S_AXIS_CTRL_TDATA_delay[10]);
    $setuphold (posedge S_AXIS_CTRL_ACLK, negedge S_AXIS_CTRL_TDATA[11], 0:0:0, 0:0:0, notifier, , , S_AXIS_CTRL_ACLK_delay, S_AXIS_CTRL_TDATA_delay[11]);
    $setuphold (posedge S_AXIS_CTRL_ACLK, negedge S_AXIS_CTRL_TDATA[12], 0:0:0, 0:0:0, notifier, , , S_AXIS_CTRL_ACLK_delay, S_AXIS_CTRL_TDATA_delay[12]);
    $setuphold (posedge S_AXIS_CTRL_ACLK, negedge S_AXIS_CTRL_TDATA[13], 0:0:0, 0:0:0, notifier, , , S_AXIS_CTRL_ACLK_delay, S_AXIS_CTRL_TDATA_delay[13]);
    $setuphold (posedge S_AXIS_CTRL_ACLK, negedge S_AXIS_CTRL_TDATA[14], 0:0:0, 0:0:0, notifier, , , S_AXIS_CTRL_ACLK_delay, S_AXIS_CTRL_TDATA_delay[14]);
    $setuphold (posedge S_AXIS_CTRL_ACLK, negedge S_AXIS_CTRL_TDATA[15], 0:0:0, 0:0:0, notifier, , , S_AXIS_CTRL_ACLK_delay, S_AXIS_CTRL_TDATA_delay[15]);
    $setuphold (posedge S_AXIS_CTRL_ACLK, negedge S_AXIS_CTRL_TDATA[16], 0:0:0, 0:0:0, notifier, , , S_AXIS_CTRL_ACLK_delay, S_AXIS_CTRL_TDATA_delay[16]);
    $setuphold (posedge S_AXIS_CTRL_ACLK, negedge S_AXIS_CTRL_TDATA[17], 0:0:0, 0:0:0, notifier, , , S_AXIS_CTRL_ACLK_delay, S_AXIS_CTRL_TDATA_delay[17]);
    $setuphold (posedge S_AXIS_CTRL_ACLK, negedge S_AXIS_CTRL_TDATA[18], 0:0:0, 0:0:0, notifier, , , S_AXIS_CTRL_ACLK_delay, S_AXIS_CTRL_TDATA_delay[18]);
    $setuphold (posedge S_AXIS_CTRL_ACLK, negedge S_AXIS_CTRL_TDATA[19], 0:0:0, 0:0:0, notifier, , , S_AXIS_CTRL_ACLK_delay, S_AXIS_CTRL_TDATA_delay[19]);
    $setuphold (posedge S_AXIS_CTRL_ACLK, negedge S_AXIS_CTRL_TDATA[1], 0:0:0, 0:0:0, notifier, , , S_AXIS_CTRL_ACLK_delay, S_AXIS_CTRL_TDATA_delay[1]);
    $setuphold (posedge S_AXIS_CTRL_ACLK, negedge S_AXIS_CTRL_TDATA[20], 0:0:0, 0:0:0, notifier, , , S_AXIS_CTRL_ACLK_delay, S_AXIS_CTRL_TDATA_delay[20]);
    $setuphold (posedge S_AXIS_CTRL_ACLK, negedge S_AXIS_CTRL_TDATA[21], 0:0:0, 0:0:0, notifier, , , S_AXIS_CTRL_ACLK_delay, S_AXIS_CTRL_TDATA_delay[21]);
    $setuphold (posedge S_AXIS_CTRL_ACLK, negedge S_AXIS_CTRL_TDATA[22], 0:0:0, 0:0:0, notifier, , , S_AXIS_CTRL_ACLK_delay, S_AXIS_CTRL_TDATA_delay[22]);
    $setuphold (posedge S_AXIS_CTRL_ACLK, negedge S_AXIS_CTRL_TDATA[23], 0:0:0, 0:0:0, notifier, , , S_AXIS_CTRL_ACLK_delay, S_AXIS_CTRL_TDATA_delay[23]);
    $setuphold (posedge S_AXIS_CTRL_ACLK, negedge S_AXIS_CTRL_TDATA[24], 0:0:0, 0:0:0, notifier, , , S_AXIS_CTRL_ACLK_delay, S_AXIS_CTRL_TDATA_delay[24]);
    $setuphold (posedge S_AXIS_CTRL_ACLK, negedge S_AXIS_CTRL_TDATA[25], 0:0:0, 0:0:0, notifier, , , S_AXIS_CTRL_ACLK_delay, S_AXIS_CTRL_TDATA_delay[25]);
    $setuphold (posedge S_AXIS_CTRL_ACLK, negedge S_AXIS_CTRL_TDATA[26], 0:0:0, 0:0:0, notifier, , , S_AXIS_CTRL_ACLK_delay, S_AXIS_CTRL_TDATA_delay[26]);
    $setuphold (posedge S_AXIS_CTRL_ACLK, negedge S_AXIS_CTRL_TDATA[27], 0:0:0, 0:0:0, notifier, , , S_AXIS_CTRL_ACLK_delay, S_AXIS_CTRL_TDATA_delay[27]);
    $setuphold (posedge S_AXIS_CTRL_ACLK, negedge S_AXIS_CTRL_TDATA[28], 0:0:0, 0:0:0, notifier, , , S_AXIS_CTRL_ACLK_delay, S_AXIS_CTRL_TDATA_delay[28]);
    $setuphold (posedge S_AXIS_CTRL_ACLK, negedge S_AXIS_CTRL_TDATA[29], 0:0:0, 0:0:0, notifier, , , S_AXIS_CTRL_ACLK_delay, S_AXIS_CTRL_TDATA_delay[29]);
    $setuphold (posedge S_AXIS_CTRL_ACLK, negedge S_AXIS_CTRL_TDATA[2], 0:0:0, 0:0:0, notifier, , , S_AXIS_CTRL_ACLK_delay, S_AXIS_CTRL_TDATA_delay[2]);
    $setuphold (posedge S_AXIS_CTRL_ACLK, negedge S_AXIS_CTRL_TDATA[30], 0:0:0, 0:0:0, notifier, , , S_AXIS_CTRL_ACLK_delay, S_AXIS_CTRL_TDATA_delay[30]);
    $setuphold (posedge S_AXIS_CTRL_ACLK, negedge S_AXIS_CTRL_TDATA[31], 0:0:0, 0:0:0, notifier, , , S_AXIS_CTRL_ACLK_delay, S_AXIS_CTRL_TDATA_delay[31]);
    $setuphold (posedge S_AXIS_CTRL_ACLK, negedge S_AXIS_CTRL_TDATA[3], 0:0:0, 0:0:0, notifier, , , S_AXIS_CTRL_ACLK_delay, S_AXIS_CTRL_TDATA_delay[3]);
    $setuphold (posedge S_AXIS_CTRL_ACLK, negedge S_AXIS_CTRL_TDATA[4], 0:0:0, 0:0:0, notifier, , , S_AXIS_CTRL_ACLK_delay, S_AXIS_CTRL_TDATA_delay[4]);
    $setuphold (posedge S_AXIS_CTRL_ACLK, negedge S_AXIS_CTRL_TDATA[5], 0:0:0, 0:0:0, notifier, , , S_AXIS_CTRL_ACLK_delay, S_AXIS_CTRL_TDATA_delay[5]);
    $setuphold (posedge S_AXIS_CTRL_ACLK, negedge S_AXIS_CTRL_TDATA[6], 0:0:0, 0:0:0, notifier, , , S_AXIS_CTRL_ACLK_delay, S_AXIS_CTRL_TDATA_delay[6]);
    $setuphold (posedge S_AXIS_CTRL_ACLK, negedge S_AXIS_CTRL_TDATA[7], 0:0:0, 0:0:0, notifier, , , S_AXIS_CTRL_ACLK_delay, S_AXIS_CTRL_TDATA_delay[7]);
    $setuphold (posedge S_AXIS_CTRL_ACLK, negedge S_AXIS_CTRL_TDATA[8], 0:0:0, 0:0:0, notifier, , , S_AXIS_CTRL_ACLK_delay, S_AXIS_CTRL_TDATA_delay[8]);
    $setuphold (posedge S_AXIS_CTRL_ACLK, negedge S_AXIS_CTRL_TDATA[9], 0:0:0, 0:0:0, notifier, , , S_AXIS_CTRL_ACLK_delay, S_AXIS_CTRL_TDATA_delay[9]);
    $setuphold (posedge S_AXIS_CTRL_ACLK, negedge S_AXIS_CTRL_TVALID, 0:0:0, 0:0:0, notifier, , , S_AXIS_CTRL_ACLK_delay, S_AXIS_CTRL_TVALID_delay);
    $setuphold (posedge S_AXIS_CTRL_ACLK, posedge S_AXIS_CTRL_TDATA[0], 0:0:0, 0:0:0, notifier, , , S_AXIS_CTRL_ACLK_delay, S_AXIS_CTRL_TDATA_delay[0]);
    $setuphold (posedge S_AXIS_CTRL_ACLK, posedge S_AXIS_CTRL_TDATA[10], 0:0:0, 0:0:0, notifier, , , S_AXIS_CTRL_ACLK_delay, S_AXIS_CTRL_TDATA_delay[10]);
    $setuphold (posedge S_AXIS_CTRL_ACLK, posedge S_AXIS_CTRL_TDATA[11], 0:0:0, 0:0:0, notifier, , , S_AXIS_CTRL_ACLK_delay, S_AXIS_CTRL_TDATA_delay[11]);
    $setuphold (posedge S_AXIS_CTRL_ACLK, posedge S_AXIS_CTRL_TDATA[12], 0:0:0, 0:0:0, notifier, , , S_AXIS_CTRL_ACLK_delay, S_AXIS_CTRL_TDATA_delay[12]);
    $setuphold (posedge S_AXIS_CTRL_ACLK, posedge S_AXIS_CTRL_TDATA[13], 0:0:0, 0:0:0, notifier, , , S_AXIS_CTRL_ACLK_delay, S_AXIS_CTRL_TDATA_delay[13]);
    $setuphold (posedge S_AXIS_CTRL_ACLK, posedge S_AXIS_CTRL_TDATA[14], 0:0:0, 0:0:0, notifier, , , S_AXIS_CTRL_ACLK_delay, S_AXIS_CTRL_TDATA_delay[14]);
    $setuphold (posedge S_AXIS_CTRL_ACLK, posedge S_AXIS_CTRL_TDATA[15], 0:0:0, 0:0:0, notifier, , , S_AXIS_CTRL_ACLK_delay, S_AXIS_CTRL_TDATA_delay[15]);
    $setuphold (posedge S_AXIS_CTRL_ACLK, posedge S_AXIS_CTRL_TDATA[16], 0:0:0, 0:0:0, notifier, , , S_AXIS_CTRL_ACLK_delay, S_AXIS_CTRL_TDATA_delay[16]);
    $setuphold (posedge S_AXIS_CTRL_ACLK, posedge S_AXIS_CTRL_TDATA[17], 0:0:0, 0:0:0, notifier, , , S_AXIS_CTRL_ACLK_delay, S_AXIS_CTRL_TDATA_delay[17]);
    $setuphold (posedge S_AXIS_CTRL_ACLK, posedge S_AXIS_CTRL_TDATA[18], 0:0:0, 0:0:0, notifier, , , S_AXIS_CTRL_ACLK_delay, S_AXIS_CTRL_TDATA_delay[18]);
    $setuphold (posedge S_AXIS_CTRL_ACLK, posedge S_AXIS_CTRL_TDATA[19], 0:0:0, 0:0:0, notifier, , , S_AXIS_CTRL_ACLK_delay, S_AXIS_CTRL_TDATA_delay[19]);
    $setuphold (posedge S_AXIS_CTRL_ACLK, posedge S_AXIS_CTRL_TDATA[1], 0:0:0, 0:0:0, notifier, , , S_AXIS_CTRL_ACLK_delay, S_AXIS_CTRL_TDATA_delay[1]);
    $setuphold (posedge S_AXIS_CTRL_ACLK, posedge S_AXIS_CTRL_TDATA[20], 0:0:0, 0:0:0, notifier, , , S_AXIS_CTRL_ACLK_delay, S_AXIS_CTRL_TDATA_delay[20]);
    $setuphold (posedge S_AXIS_CTRL_ACLK, posedge S_AXIS_CTRL_TDATA[21], 0:0:0, 0:0:0, notifier, , , S_AXIS_CTRL_ACLK_delay, S_AXIS_CTRL_TDATA_delay[21]);
    $setuphold (posedge S_AXIS_CTRL_ACLK, posedge S_AXIS_CTRL_TDATA[22], 0:0:0, 0:0:0, notifier, , , S_AXIS_CTRL_ACLK_delay, S_AXIS_CTRL_TDATA_delay[22]);
    $setuphold (posedge S_AXIS_CTRL_ACLK, posedge S_AXIS_CTRL_TDATA[23], 0:0:0, 0:0:0, notifier, , , S_AXIS_CTRL_ACLK_delay, S_AXIS_CTRL_TDATA_delay[23]);
    $setuphold (posedge S_AXIS_CTRL_ACLK, posedge S_AXIS_CTRL_TDATA[24], 0:0:0, 0:0:0, notifier, , , S_AXIS_CTRL_ACLK_delay, S_AXIS_CTRL_TDATA_delay[24]);
    $setuphold (posedge S_AXIS_CTRL_ACLK, posedge S_AXIS_CTRL_TDATA[25], 0:0:0, 0:0:0, notifier, , , S_AXIS_CTRL_ACLK_delay, S_AXIS_CTRL_TDATA_delay[25]);
    $setuphold (posedge S_AXIS_CTRL_ACLK, posedge S_AXIS_CTRL_TDATA[26], 0:0:0, 0:0:0, notifier, , , S_AXIS_CTRL_ACLK_delay, S_AXIS_CTRL_TDATA_delay[26]);
    $setuphold (posedge S_AXIS_CTRL_ACLK, posedge S_AXIS_CTRL_TDATA[27], 0:0:0, 0:0:0, notifier, , , S_AXIS_CTRL_ACLK_delay, S_AXIS_CTRL_TDATA_delay[27]);
    $setuphold (posedge S_AXIS_CTRL_ACLK, posedge S_AXIS_CTRL_TDATA[28], 0:0:0, 0:0:0, notifier, , , S_AXIS_CTRL_ACLK_delay, S_AXIS_CTRL_TDATA_delay[28]);
    $setuphold (posedge S_AXIS_CTRL_ACLK, posedge S_AXIS_CTRL_TDATA[29], 0:0:0, 0:0:0, notifier, , , S_AXIS_CTRL_ACLK_delay, S_AXIS_CTRL_TDATA_delay[29]);
    $setuphold (posedge S_AXIS_CTRL_ACLK, posedge S_AXIS_CTRL_TDATA[2], 0:0:0, 0:0:0, notifier, , , S_AXIS_CTRL_ACLK_delay, S_AXIS_CTRL_TDATA_delay[2]);
    $setuphold (posedge S_AXIS_CTRL_ACLK, posedge S_AXIS_CTRL_TDATA[30], 0:0:0, 0:0:0, notifier, , , S_AXIS_CTRL_ACLK_delay, S_AXIS_CTRL_TDATA_delay[30]);
    $setuphold (posedge S_AXIS_CTRL_ACLK, posedge S_AXIS_CTRL_TDATA[31], 0:0:0, 0:0:0, notifier, , , S_AXIS_CTRL_ACLK_delay, S_AXIS_CTRL_TDATA_delay[31]);
    $setuphold (posedge S_AXIS_CTRL_ACLK, posedge S_AXIS_CTRL_TDATA[3], 0:0:0, 0:0:0, notifier, , , S_AXIS_CTRL_ACLK_delay, S_AXIS_CTRL_TDATA_delay[3]);
    $setuphold (posedge S_AXIS_CTRL_ACLK, posedge S_AXIS_CTRL_TDATA[4], 0:0:0, 0:0:0, notifier, , , S_AXIS_CTRL_ACLK_delay, S_AXIS_CTRL_TDATA_delay[4]);
    $setuphold (posedge S_AXIS_CTRL_ACLK, posedge S_AXIS_CTRL_TDATA[5], 0:0:0, 0:0:0, notifier, , , S_AXIS_CTRL_ACLK_delay, S_AXIS_CTRL_TDATA_delay[5]);
    $setuphold (posedge S_AXIS_CTRL_ACLK, posedge S_AXIS_CTRL_TDATA[6], 0:0:0, 0:0:0, notifier, , , S_AXIS_CTRL_ACLK_delay, S_AXIS_CTRL_TDATA_delay[6]);
    $setuphold (posedge S_AXIS_CTRL_ACLK, posedge S_AXIS_CTRL_TDATA[7], 0:0:0, 0:0:0, notifier, , , S_AXIS_CTRL_ACLK_delay, S_AXIS_CTRL_TDATA_delay[7]);
    $setuphold (posedge S_AXIS_CTRL_ACLK, posedge S_AXIS_CTRL_TDATA[8], 0:0:0, 0:0:0, notifier, , , S_AXIS_CTRL_ACLK_delay, S_AXIS_CTRL_TDATA_delay[8]);
    $setuphold (posedge S_AXIS_CTRL_ACLK, posedge S_AXIS_CTRL_TDATA[9], 0:0:0, 0:0:0, notifier, , , S_AXIS_CTRL_ACLK_delay, S_AXIS_CTRL_TDATA_delay[9]);
    $setuphold (posedge S_AXIS_CTRL_ACLK, posedge S_AXIS_CTRL_TVALID, 0:0:0, 0:0:0, notifier, , , S_AXIS_CTRL_ACLK_delay, S_AXIS_CTRL_TVALID_delay);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[0], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[0]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[100], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[100]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[101], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[101]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[102], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[102]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[103], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[103]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[104], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[104]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[105], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[105]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[106], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[106]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[107], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[107]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[108], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[108]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[109], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[109]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[10], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[10]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[110], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[110]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[111], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[111]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[112], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[112]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[113], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[113]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[114], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[114]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[115], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[115]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[116], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[116]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[117], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[117]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[118], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[118]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[119], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[119]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[11], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[11]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[120], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[120]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[121], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[121]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[122], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[122]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[123], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[123]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[124], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[124]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[125], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[125]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[126], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[126]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[127], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[127]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[128], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[128]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[129], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[129]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[12], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[12]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[130], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[130]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[131], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[131]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[132], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[132]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[133], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[133]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[134], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[134]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[135], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[135]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[136], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[136]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[137], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[137]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[138], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[138]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[139], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[139]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[13], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[13]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[140], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[140]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[141], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[141]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[142], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[142]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[143], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[143]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[144], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[144]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[145], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[145]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[146], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[146]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[147], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[147]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[148], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[148]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[149], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[149]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[14], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[14]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[150], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[150]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[151], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[151]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[152], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[152]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[153], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[153]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[154], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[154]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[155], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[155]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[156], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[156]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[157], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[157]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[158], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[158]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[159], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[159]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[15], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[15]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[160], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[160]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[161], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[161]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[162], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[162]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[163], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[163]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[164], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[164]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[165], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[165]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[166], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[166]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[167], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[167]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[168], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[168]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[169], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[169]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[16], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[16]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[170], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[170]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[171], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[171]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[172], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[172]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[173], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[173]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[174], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[174]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[175], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[175]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[176], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[176]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[177], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[177]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[178], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[178]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[179], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[179]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[17], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[17]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[180], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[180]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[181], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[181]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[182], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[182]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[183], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[183]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[184], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[184]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[185], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[185]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[186], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[186]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[187], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[187]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[188], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[188]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[189], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[189]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[18], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[18]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[190], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[190]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[191], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[191]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[192], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[192]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[193], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[193]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[194], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[194]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[195], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[195]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[196], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[196]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[197], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[197]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[198], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[198]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[199], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[199]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[19], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[19]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[1], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[1]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[200], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[200]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[201], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[201]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[202], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[202]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[203], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[203]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[204], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[204]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[205], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[205]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[206], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[206]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[207], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[207]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[208], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[208]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[209], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[209]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[20], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[20]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[210], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[210]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[211], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[211]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[212], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[212]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[213], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[213]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[214], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[214]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[215], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[215]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[216], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[216]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[217], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[217]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[218], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[218]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[219], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[219]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[21], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[21]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[220], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[220]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[221], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[221]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[222], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[222]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[223], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[223]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[224], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[224]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[225], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[225]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[226], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[226]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[227], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[227]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[228], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[228]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[229], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[229]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[22], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[22]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[230], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[230]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[231], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[231]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[232], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[232]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[233], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[233]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[234], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[234]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[235], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[235]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[236], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[236]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[237], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[237]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[238], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[238]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[239], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[239]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[23], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[23]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[240], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[240]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[241], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[241]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[242], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[242]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[243], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[243]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[244], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[244]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[245], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[245]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[246], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[246]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[247], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[247]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[248], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[248]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[249], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[249]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[24], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[24]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[250], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[250]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[251], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[251]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[252], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[252]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[253], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[253]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[254], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[254]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[255], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[255]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[256], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[256]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[257], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[257]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[258], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[258]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[259], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[259]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[25], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[25]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[260], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[260]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[261], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[261]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[262], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[262]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[263], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[263]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[264], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[264]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[265], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[265]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[266], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[266]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[267], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[267]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[268], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[268]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[269], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[269]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[26], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[26]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[270], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[270]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[271], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[271]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[272], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[272]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[273], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[273]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[274], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[274]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[275], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[275]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[276], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[276]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[277], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[277]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[278], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[278]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[279], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[279]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[27], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[27]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[280], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[280]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[281], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[281]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[282], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[282]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[283], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[283]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[284], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[284]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[285], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[285]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[286], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[286]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[287], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[287]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[288], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[288]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[289], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[289]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[28], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[28]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[290], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[290]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[291], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[291]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[292], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[292]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[293], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[293]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[294], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[294]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[295], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[295]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[296], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[296]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[297], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[297]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[298], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[298]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[299], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[299]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[29], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[29]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[2], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[2]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[300], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[300]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[301], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[301]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[302], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[302]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[303], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[303]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[304], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[304]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[305], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[305]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[306], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[306]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[307], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[307]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[308], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[308]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[309], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[309]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[30], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[30]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[310], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[310]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[311], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[311]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[312], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[312]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[313], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[313]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[314], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[314]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[315], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[315]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[316], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[316]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[317], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[317]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[318], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[318]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[319], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[319]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[31], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[31]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[320], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[320]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[321], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[321]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[322], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[322]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[323], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[323]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[324], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[324]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[325], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[325]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[326], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[326]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[327], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[327]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[328], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[328]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[329], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[329]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[32], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[32]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[330], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[330]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[331], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[331]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[332], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[332]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[333], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[333]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[334], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[334]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[335], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[335]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[336], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[336]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[337], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[337]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[338], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[338]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[339], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[339]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[33], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[33]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[340], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[340]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[341], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[341]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[342], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[342]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[343], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[343]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[344], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[344]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[345], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[345]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[346], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[346]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[347], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[347]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[348], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[348]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[349], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[349]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[34], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[34]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[350], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[350]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[351], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[351]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[352], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[352]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[353], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[353]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[354], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[354]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[355], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[355]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[356], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[356]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[357], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[357]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[358], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[358]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[359], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[359]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[35], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[35]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[360], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[360]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[361], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[361]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[362], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[362]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[363], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[363]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[364], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[364]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[365], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[365]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[366], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[366]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[367], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[367]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[368], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[368]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[369], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[369]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[36], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[36]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[370], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[370]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[371], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[371]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[372], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[372]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[373], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[373]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[374], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[374]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[375], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[375]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[376], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[376]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[377], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[377]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[378], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[378]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[379], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[379]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[37], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[37]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[380], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[380]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[381], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[381]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[382], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[382]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[383], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[383]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[384], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[384]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[385], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[385]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[386], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[386]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[387], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[387]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[388], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[388]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[389], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[389]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[38], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[38]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[390], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[390]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[391], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[391]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[392], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[392]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[393], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[393]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[394], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[394]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[395], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[395]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[396], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[396]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[397], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[397]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[398], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[398]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[399], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[399]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[39], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[39]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[3], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[3]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[400], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[400]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[401], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[401]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[402], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[402]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[403], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[403]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[404], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[404]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[405], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[405]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[406], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[406]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[407], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[407]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[408], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[408]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[409], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[409]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[40], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[40]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[410], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[410]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[411], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[411]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[412], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[412]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[413], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[413]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[414], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[414]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[415], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[415]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[416], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[416]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[417], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[417]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[418], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[418]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[419], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[419]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[41], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[41]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[420], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[420]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[421], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[421]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[422], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[422]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[423], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[423]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[424], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[424]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[425], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[425]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[426], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[426]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[427], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[427]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[428], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[428]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[429], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[429]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[42], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[42]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[430], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[430]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[431], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[431]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[432], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[432]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[433], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[433]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[434], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[434]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[435], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[435]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[436], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[436]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[437], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[437]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[438], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[438]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[439], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[439]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[43], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[43]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[440], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[440]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[441], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[441]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[442], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[442]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[443], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[443]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[444], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[444]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[445], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[445]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[446], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[446]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[447], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[447]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[448], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[448]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[449], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[449]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[44], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[44]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[450], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[450]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[451], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[451]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[452], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[452]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[453], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[453]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[454], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[454]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[455], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[455]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[456], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[456]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[457], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[457]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[458], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[458]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[459], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[459]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[45], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[45]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[460], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[460]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[461], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[461]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[462], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[462]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[463], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[463]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[464], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[464]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[465], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[465]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[466], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[466]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[467], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[467]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[468], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[468]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[469], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[469]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[46], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[46]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[470], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[470]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[471], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[471]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[472], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[472]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[473], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[473]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[474], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[474]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[475], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[475]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[476], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[476]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[477], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[477]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[478], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[478]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[479], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[479]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[47], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[47]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[480], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[480]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[481], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[481]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[482], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[482]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[483], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[483]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[484], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[484]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[485], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[485]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[486], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[486]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[487], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[487]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[488], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[488]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[489], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[489]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[48], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[48]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[490], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[490]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[491], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[491]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[492], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[492]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[493], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[493]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[494], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[494]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[495], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[495]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[496], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[496]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[497], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[497]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[498], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[498]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[499], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[499]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[49], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[49]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[4], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[4]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[500], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[500]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[501], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[501]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[502], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[502]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[503], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[503]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[504], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[504]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[505], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[505]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[506], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[506]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[507], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[507]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[508], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[508]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[509], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[509]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[50], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[50]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[510], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[510]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[511], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[511]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[51], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[51]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[52], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[52]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[53], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[53]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[54], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[54]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[55], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[55]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[56], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[56]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[57], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[57]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[58], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[58]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[59], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[59]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[5], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[5]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[60], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[60]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[61], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[61]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[62], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[62]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[63], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[63]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[64], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[64]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[65], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[65]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[66], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[66]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[67], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[67]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[68], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[68]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[69], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[69]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[6], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[6]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[70], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[70]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[71], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[71]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[72], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[72]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[73], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[73]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[74], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[74]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[75], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[75]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[76], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[76]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[77], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[77]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[78], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[78]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[79], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[79]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[7], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[7]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[80], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[80]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[81], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[81]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[82], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[82]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[83], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[83]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[84], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[84]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[85], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[85]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[86], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[86]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[87], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[87]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[88], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[88]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[89], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[89]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[8], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[8]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[90], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[90]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[91], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[91]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[92], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[92]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[93], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[93]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[94], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[94]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[95], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[95]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[96], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[96]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[97], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[97]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[98], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[98]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[99], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[99]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TDATA[9], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[9]);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TLAST, 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TLAST_delay);
    $setuphold (posedge S_AXIS_DIN_ACLK, negedge S_AXIS_DIN_TVALID, 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TVALID_delay);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[0], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[0]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[100], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[100]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[101], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[101]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[102], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[102]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[103], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[103]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[104], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[104]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[105], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[105]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[106], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[106]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[107], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[107]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[108], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[108]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[109], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[109]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[10], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[10]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[110], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[110]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[111], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[111]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[112], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[112]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[113], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[113]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[114], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[114]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[115], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[115]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[116], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[116]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[117], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[117]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[118], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[118]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[119], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[119]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[11], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[11]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[120], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[120]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[121], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[121]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[122], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[122]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[123], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[123]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[124], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[124]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[125], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[125]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[126], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[126]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[127], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[127]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[128], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[128]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[129], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[129]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[12], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[12]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[130], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[130]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[131], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[131]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[132], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[132]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[133], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[133]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[134], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[134]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[135], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[135]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[136], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[136]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[137], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[137]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[138], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[138]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[139], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[139]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[13], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[13]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[140], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[140]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[141], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[141]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[142], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[142]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[143], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[143]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[144], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[144]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[145], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[145]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[146], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[146]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[147], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[147]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[148], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[148]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[149], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[149]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[14], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[14]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[150], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[150]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[151], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[151]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[152], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[152]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[153], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[153]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[154], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[154]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[155], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[155]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[156], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[156]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[157], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[157]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[158], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[158]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[159], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[159]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[15], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[15]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[160], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[160]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[161], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[161]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[162], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[162]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[163], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[163]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[164], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[164]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[165], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[165]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[166], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[166]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[167], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[167]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[168], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[168]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[169], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[169]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[16], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[16]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[170], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[170]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[171], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[171]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[172], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[172]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[173], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[173]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[174], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[174]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[175], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[175]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[176], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[176]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[177], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[177]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[178], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[178]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[179], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[179]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[17], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[17]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[180], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[180]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[181], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[181]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[182], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[182]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[183], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[183]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[184], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[184]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[185], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[185]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[186], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[186]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[187], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[187]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[188], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[188]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[189], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[189]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[18], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[18]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[190], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[190]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[191], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[191]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[192], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[192]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[193], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[193]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[194], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[194]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[195], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[195]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[196], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[196]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[197], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[197]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[198], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[198]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[199], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[199]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[19], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[19]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[1], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[1]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[200], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[200]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[201], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[201]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[202], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[202]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[203], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[203]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[204], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[204]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[205], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[205]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[206], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[206]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[207], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[207]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[208], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[208]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[209], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[209]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[20], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[20]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[210], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[210]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[211], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[211]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[212], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[212]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[213], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[213]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[214], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[214]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[215], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[215]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[216], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[216]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[217], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[217]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[218], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[218]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[219], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[219]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[21], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[21]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[220], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[220]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[221], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[221]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[222], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[222]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[223], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[223]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[224], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[224]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[225], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[225]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[226], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[226]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[227], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[227]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[228], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[228]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[229], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[229]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[22], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[22]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[230], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[230]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[231], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[231]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[232], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[232]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[233], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[233]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[234], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[234]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[235], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[235]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[236], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[236]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[237], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[237]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[238], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[238]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[239], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[239]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[23], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[23]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[240], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[240]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[241], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[241]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[242], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[242]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[243], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[243]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[244], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[244]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[245], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[245]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[246], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[246]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[247], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[247]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[248], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[248]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[249], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[249]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[24], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[24]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[250], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[250]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[251], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[251]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[252], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[252]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[253], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[253]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[254], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[254]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[255], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[255]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[256], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[256]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[257], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[257]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[258], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[258]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[259], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[259]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[25], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[25]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[260], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[260]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[261], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[261]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[262], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[262]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[263], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[263]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[264], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[264]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[265], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[265]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[266], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[266]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[267], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[267]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[268], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[268]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[269], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[269]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[26], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[26]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[270], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[270]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[271], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[271]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[272], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[272]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[273], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[273]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[274], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[274]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[275], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[275]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[276], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[276]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[277], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[277]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[278], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[278]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[279], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[279]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[27], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[27]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[280], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[280]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[281], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[281]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[282], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[282]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[283], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[283]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[284], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[284]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[285], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[285]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[286], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[286]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[287], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[287]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[288], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[288]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[289], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[289]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[28], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[28]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[290], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[290]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[291], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[291]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[292], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[292]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[293], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[293]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[294], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[294]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[295], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[295]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[296], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[296]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[297], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[297]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[298], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[298]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[299], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[299]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[29], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[29]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[2], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[2]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[300], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[300]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[301], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[301]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[302], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[302]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[303], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[303]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[304], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[304]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[305], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[305]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[306], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[306]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[307], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[307]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[308], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[308]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[309], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[309]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[30], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[30]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[310], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[310]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[311], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[311]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[312], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[312]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[313], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[313]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[314], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[314]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[315], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[315]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[316], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[316]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[317], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[317]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[318], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[318]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[319], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[319]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[31], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[31]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[320], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[320]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[321], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[321]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[322], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[322]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[323], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[323]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[324], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[324]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[325], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[325]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[326], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[326]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[327], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[327]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[328], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[328]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[329], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[329]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[32], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[32]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[330], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[330]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[331], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[331]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[332], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[332]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[333], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[333]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[334], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[334]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[335], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[335]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[336], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[336]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[337], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[337]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[338], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[338]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[339], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[339]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[33], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[33]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[340], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[340]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[341], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[341]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[342], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[342]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[343], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[343]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[344], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[344]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[345], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[345]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[346], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[346]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[347], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[347]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[348], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[348]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[349], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[349]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[34], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[34]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[350], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[350]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[351], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[351]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[352], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[352]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[353], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[353]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[354], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[354]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[355], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[355]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[356], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[356]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[357], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[357]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[358], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[358]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[359], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[359]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[35], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[35]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[360], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[360]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[361], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[361]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[362], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[362]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[363], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[363]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[364], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[364]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[365], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[365]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[366], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[366]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[367], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[367]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[368], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[368]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[369], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[369]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[36], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[36]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[370], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[370]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[371], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[371]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[372], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[372]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[373], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[373]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[374], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[374]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[375], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[375]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[376], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[376]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[377], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[377]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[378], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[378]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[379], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[379]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[37], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[37]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[380], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[380]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[381], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[381]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[382], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[382]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[383], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[383]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[384], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[384]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[385], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[385]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[386], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[386]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[387], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[387]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[388], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[388]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[389], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[389]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[38], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[38]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[390], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[390]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[391], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[391]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[392], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[392]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[393], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[393]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[394], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[394]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[395], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[395]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[396], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[396]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[397], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[397]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[398], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[398]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[399], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[399]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[39], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[39]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[3], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[3]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[400], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[400]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[401], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[401]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[402], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[402]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[403], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[403]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[404], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[404]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[405], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[405]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[406], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[406]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[407], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[407]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[408], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[408]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[409], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[409]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[40], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[40]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[410], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[410]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[411], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[411]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[412], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[412]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[413], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[413]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[414], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[414]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[415], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[415]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[416], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[416]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[417], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[417]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[418], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[418]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[419], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[419]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[41], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[41]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[420], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[420]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[421], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[421]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[422], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[422]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[423], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[423]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[424], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[424]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[425], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[425]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[426], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[426]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[427], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[427]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[428], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[428]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[429], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[429]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[42], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[42]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[430], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[430]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[431], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[431]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[432], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[432]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[433], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[433]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[434], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[434]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[435], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[435]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[436], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[436]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[437], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[437]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[438], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[438]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[439], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[439]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[43], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[43]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[440], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[440]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[441], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[441]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[442], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[442]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[443], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[443]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[444], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[444]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[445], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[445]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[446], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[446]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[447], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[447]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[448], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[448]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[449], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[449]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[44], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[44]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[450], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[450]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[451], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[451]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[452], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[452]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[453], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[453]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[454], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[454]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[455], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[455]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[456], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[456]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[457], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[457]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[458], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[458]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[459], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[459]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[45], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[45]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[460], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[460]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[461], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[461]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[462], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[462]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[463], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[463]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[464], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[464]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[465], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[465]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[466], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[466]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[467], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[467]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[468], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[468]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[469], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[469]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[46], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[46]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[470], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[470]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[471], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[471]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[472], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[472]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[473], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[473]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[474], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[474]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[475], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[475]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[476], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[476]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[477], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[477]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[478], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[478]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[479], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[479]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[47], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[47]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[480], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[480]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[481], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[481]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[482], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[482]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[483], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[483]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[484], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[484]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[485], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[485]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[486], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[486]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[487], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[487]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[488], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[488]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[489], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[489]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[48], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[48]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[490], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[490]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[491], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[491]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[492], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[492]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[493], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[493]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[494], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[494]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[495], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[495]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[496], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[496]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[497], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[497]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[498], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[498]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[499], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[499]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[49], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[49]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[4], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[4]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[500], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[500]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[501], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[501]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[502], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[502]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[503], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[503]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[504], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[504]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[505], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[505]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[506], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[506]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[507], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[507]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[508], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[508]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[509], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[509]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[50], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[50]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[510], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[510]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[511], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[511]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[51], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[51]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[52], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[52]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[53], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[53]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[54], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[54]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[55], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[55]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[56], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[56]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[57], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[57]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[58], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[58]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[59], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[59]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[5], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[5]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[60], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[60]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[61], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[61]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[62], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[62]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[63], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[63]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[64], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[64]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[65], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[65]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[66], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[66]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[67], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[67]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[68], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[68]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[69], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[69]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[6], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[6]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[70], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[70]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[71], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[71]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[72], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[72]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[73], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[73]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[74], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[74]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[75], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[75]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[76], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[76]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[77], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[77]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[78], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[78]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[79], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[79]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[7], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[7]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[80], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[80]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[81], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[81]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[82], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[82]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[83], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[83]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[84], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[84]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[85], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[85]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[86], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[86]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[87], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[87]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[88], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[88]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[89], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[89]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[8], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[8]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[90], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[90]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[91], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[91]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[92], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[92]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[93], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[93]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[94], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[94]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[95], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[95]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[96], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[96]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[97], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[97]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[98], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[98]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[99], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[99]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TDATA[9], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TDATA_delay[9]);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TLAST, 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TLAST_delay);
    $setuphold (posedge S_AXIS_DIN_ACLK, posedge S_AXIS_DIN_TVALID, 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_ACLK_delay, S_AXIS_DIN_TVALID_delay);
    $setuphold (posedge S_AXIS_DIN_WORDS_ACLK, negedge S_AXIS_DIN_WORDS_TDATA[0], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_WORDS_ACLK_delay, S_AXIS_DIN_WORDS_TDATA_delay[0]);
    $setuphold (posedge S_AXIS_DIN_WORDS_ACLK, negedge S_AXIS_DIN_WORDS_TDATA[10], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_WORDS_ACLK_delay, S_AXIS_DIN_WORDS_TDATA_delay[10]);
    $setuphold (posedge S_AXIS_DIN_WORDS_ACLK, negedge S_AXIS_DIN_WORDS_TDATA[11], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_WORDS_ACLK_delay, S_AXIS_DIN_WORDS_TDATA_delay[11]);
    $setuphold (posedge S_AXIS_DIN_WORDS_ACLK, negedge S_AXIS_DIN_WORDS_TDATA[12], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_WORDS_ACLK_delay, S_AXIS_DIN_WORDS_TDATA_delay[12]);
    $setuphold (posedge S_AXIS_DIN_WORDS_ACLK, negedge S_AXIS_DIN_WORDS_TDATA[16], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_WORDS_ACLK_delay, S_AXIS_DIN_WORDS_TDATA_delay[16]);
    $setuphold (posedge S_AXIS_DIN_WORDS_ACLK, negedge S_AXIS_DIN_WORDS_TDATA[17], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_WORDS_ACLK_delay, S_AXIS_DIN_WORDS_TDATA_delay[17]);
    $setuphold (posedge S_AXIS_DIN_WORDS_ACLK, negedge S_AXIS_DIN_WORDS_TDATA[18], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_WORDS_ACLK_delay, S_AXIS_DIN_WORDS_TDATA_delay[18]);
    $setuphold (posedge S_AXIS_DIN_WORDS_ACLK, negedge S_AXIS_DIN_WORDS_TDATA[19], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_WORDS_ACLK_delay, S_AXIS_DIN_WORDS_TDATA_delay[19]);
    $setuphold (posedge S_AXIS_DIN_WORDS_ACLK, negedge S_AXIS_DIN_WORDS_TDATA[1], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_WORDS_ACLK_delay, S_AXIS_DIN_WORDS_TDATA_delay[1]);
    $setuphold (posedge S_AXIS_DIN_WORDS_ACLK, negedge S_AXIS_DIN_WORDS_TDATA[20], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_WORDS_ACLK_delay, S_AXIS_DIN_WORDS_TDATA_delay[20]);
    $setuphold (posedge S_AXIS_DIN_WORDS_ACLK, negedge S_AXIS_DIN_WORDS_TDATA[24], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_WORDS_ACLK_delay, S_AXIS_DIN_WORDS_TDATA_delay[24]);
    $setuphold (posedge S_AXIS_DIN_WORDS_ACLK, negedge S_AXIS_DIN_WORDS_TDATA[25], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_WORDS_ACLK_delay, S_AXIS_DIN_WORDS_TDATA_delay[25]);
    $setuphold (posedge S_AXIS_DIN_WORDS_ACLK, negedge S_AXIS_DIN_WORDS_TDATA[26], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_WORDS_ACLK_delay, S_AXIS_DIN_WORDS_TDATA_delay[26]);
    $setuphold (posedge S_AXIS_DIN_WORDS_ACLK, negedge S_AXIS_DIN_WORDS_TDATA[27], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_WORDS_ACLK_delay, S_AXIS_DIN_WORDS_TDATA_delay[27]);
    $setuphold (posedge S_AXIS_DIN_WORDS_ACLK, negedge S_AXIS_DIN_WORDS_TDATA[28], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_WORDS_ACLK_delay, S_AXIS_DIN_WORDS_TDATA_delay[28]);
    $setuphold (posedge S_AXIS_DIN_WORDS_ACLK, negedge S_AXIS_DIN_WORDS_TDATA[2], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_WORDS_ACLK_delay, S_AXIS_DIN_WORDS_TDATA_delay[2]);
    $setuphold (posedge S_AXIS_DIN_WORDS_ACLK, negedge S_AXIS_DIN_WORDS_TDATA[3], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_WORDS_ACLK_delay, S_AXIS_DIN_WORDS_TDATA_delay[3]);
    $setuphold (posedge S_AXIS_DIN_WORDS_ACLK, negedge S_AXIS_DIN_WORDS_TDATA[4], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_WORDS_ACLK_delay, S_AXIS_DIN_WORDS_TDATA_delay[4]);
    $setuphold (posedge S_AXIS_DIN_WORDS_ACLK, negedge S_AXIS_DIN_WORDS_TDATA[8], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_WORDS_ACLK_delay, S_AXIS_DIN_WORDS_TDATA_delay[8]);
    $setuphold (posedge S_AXIS_DIN_WORDS_ACLK, negedge S_AXIS_DIN_WORDS_TDATA[9], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_WORDS_ACLK_delay, S_AXIS_DIN_WORDS_TDATA_delay[9]);
    $setuphold (posedge S_AXIS_DIN_WORDS_ACLK, negedge S_AXIS_DIN_WORDS_TLAST, 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_WORDS_ACLK_delay, S_AXIS_DIN_WORDS_TLAST_delay);
    $setuphold (posedge S_AXIS_DIN_WORDS_ACLK, negedge S_AXIS_DIN_WORDS_TVALID, 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_WORDS_ACLK_delay, S_AXIS_DIN_WORDS_TVALID_delay);
    $setuphold (posedge S_AXIS_DIN_WORDS_ACLK, posedge S_AXIS_DIN_WORDS_TDATA[0], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_WORDS_ACLK_delay, S_AXIS_DIN_WORDS_TDATA_delay[0]);
    $setuphold (posedge S_AXIS_DIN_WORDS_ACLK, posedge S_AXIS_DIN_WORDS_TDATA[10], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_WORDS_ACLK_delay, S_AXIS_DIN_WORDS_TDATA_delay[10]);
    $setuphold (posedge S_AXIS_DIN_WORDS_ACLK, posedge S_AXIS_DIN_WORDS_TDATA[11], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_WORDS_ACLK_delay, S_AXIS_DIN_WORDS_TDATA_delay[11]);
    $setuphold (posedge S_AXIS_DIN_WORDS_ACLK, posedge S_AXIS_DIN_WORDS_TDATA[12], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_WORDS_ACLK_delay, S_AXIS_DIN_WORDS_TDATA_delay[12]);
    $setuphold (posedge S_AXIS_DIN_WORDS_ACLK, posedge S_AXIS_DIN_WORDS_TDATA[16], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_WORDS_ACLK_delay, S_AXIS_DIN_WORDS_TDATA_delay[16]);
    $setuphold (posedge S_AXIS_DIN_WORDS_ACLK, posedge S_AXIS_DIN_WORDS_TDATA[17], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_WORDS_ACLK_delay, S_AXIS_DIN_WORDS_TDATA_delay[17]);
    $setuphold (posedge S_AXIS_DIN_WORDS_ACLK, posedge S_AXIS_DIN_WORDS_TDATA[18], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_WORDS_ACLK_delay, S_AXIS_DIN_WORDS_TDATA_delay[18]);
    $setuphold (posedge S_AXIS_DIN_WORDS_ACLK, posedge S_AXIS_DIN_WORDS_TDATA[19], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_WORDS_ACLK_delay, S_AXIS_DIN_WORDS_TDATA_delay[19]);
    $setuphold (posedge S_AXIS_DIN_WORDS_ACLK, posedge S_AXIS_DIN_WORDS_TDATA[1], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_WORDS_ACLK_delay, S_AXIS_DIN_WORDS_TDATA_delay[1]);
    $setuphold (posedge S_AXIS_DIN_WORDS_ACLK, posedge S_AXIS_DIN_WORDS_TDATA[20], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_WORDS_ACLK_delay, S_AXIS_DIN_WORDS_TDATA_delay[20]);
    $setuphold (posedge S_AXIS_DIN_WORDS_ACLK, posedge S_AXIS_DIN_WORDS_TDATA[24], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_WORDS_ACLK_delay, S_AXIS_DIN_WORDS_TDATA_delay[24]);
    $setuphold (posedge S_AXIS_DIN_WORDS_ACLK, posedge S_AXIS_DIN_WORDS_TDATA[25], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_WORDS_ACLK_delay, S_AXIS_DIN_WORDS_TDATA_delay[25]);
    $setuphold (posedge S_AXIS_DIN_WORDS_ACLK, posedge S_AXIS_DIN_WORDS_TDATA[26], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_WORDS_ACLK_delay, S_AXIS_DIN_WORDS_TDATA_delay[26]);
    $setuphold (posedge S_AXIS_DIN_WORDS_ACLK, posedge S_AXIS_DIN_WORDS_TDATA[27], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_WORDS_ACLK_delay, S_AXIS_DIN_WORDS_TDATA_delay[27]);
    $setuphold (posedge S_AXIS_DIN_WORDS_ACLK, posedge S_AXIS_DIN_WORDS_TDATA[28], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_WORDS_ACLK_delay, S_AXIS_DIN_WORDS_TDATA_delay[28]);
    $setuphold (posedge S_AXIS_DIN_WORDS_ACLK, posedge S_AXIS_DIN_WORDS_TDATA[2], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_WORDS_ACLK_delay, S_AXIS_DIN_WORDS_TDATA_delay[2]);
    $setuphold (posedge S_AXIS_DIN_WORDS_ACLK, posedge S_AXIS_DIN_WORDS_TDATA[3], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_WORDS_ACLK_delay, S_AXIS_DIN_WORDS_TDATA_delay[3]);
    $setuphold (posedge S_AXIS_DIN_WORDS_ACLK, posedge S_AXIS_DIN_WORDS_TDATA[4], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_WORDS_ACLK_delay, S_AXIS_DIN_WORDS_TDATA_delay[4]);
    $setuphold (posedge S_AXIS_DIN_WORDS_ACLK, posedge S_AXIS_DIN_WORDS_TDATA[8], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_WORDS_ACLK_delay, S_AXIS_DIN_WORDS_TDATA_delay[8]);
    $setuphold (posedge S_AXIS_DIN_WORDS_ACLK, posedge S_AXIS_DIN_WORDS_TDATA[9], 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_WORDS_ACLK_delay, S_AXIS_DIN_WORDS_TDATA_delay[9]);
    $setuphold (posedge S_AXIS_DIN_WORDS_ACLK, posedge S_AXIS_DIN_WORDS_TLAST, 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_WORDS_ACLK_delay, S_AXIS_DIN_WORDS_TLAST_delay);
    $setuphold (posedge S_AXIS_DIN_WORDS_ACLK, posedge S_AXIS_DIN_WORDS_TVALID, 0:0:0, 0:0:0, notifier, , , S_AXIS_DIN_WORDS_ACLK_delay, S_AXIS_DIN_WORDS_TVALID_delay);
    $setuphold (posedge S_AXIS_DOUT_WORDS_ACLK, negedge S_AXIS_DOUT_WORDS_TDATA[0], 0:0:0, 0:0:0, notifier, , , S_AXIS_DOUT_WORDS_ACLK_delay, S_AXIS_DOUT_WORDS_TDATA_delay[0]);
    $setuphold (posedge S_AXIS_DOUT_WORDS_ACLK, negedge S_AXIS_DOUT_WORDS_TDATA[10], 0:0:0, 0:0:0, notifier, , , S_AXIS_DOUT_WORDS_ACLK_delay, S_AXIS_DOUT_WORDS_TDATA_delay[10]);
    $setuphold (posedge S_AXIS_DOUT_WORDS_ACLK, negedge S_AXIS_DOUT_WORDS_TDATA[11], 0:0:0, 0:0:0, notifier, , , S_AXIS_DOUT_WORDS_ACLK_delay, S_AXIS_DOUT_WORDS_TDATA_delay[11]);
    $setuphold (posedge S_AXIS_DOUT_WORDS_ACLK, negedge S_AXIS_DOUT_WORDS_TDATA[12], 0:0:0, 0:0:0, notifier, , , S_AXIS_DOUT_WORDS_ACLK_delay, S_AXIS_DOUT_WORDS_TDATA_delay[12]);
    $setuphold (posedge S_AXIS_DOUT_WORDS_ACLK, negedge S_AXIS_DOUT_WORDS_TDATA[16], 0:0:0, 0:0:0, notifier, , , S_AXIS_DOUT_WORDS_ACLK_delay, S_AXIS_DOUT_WORDS_TDATA_delay[16]);
    $setuphold (posedge S_AXIS_DOUT_WORDS_ACLK, negedge S_AXIS_DOUT_WORDS_TDATA[17], 0:0:0, 0:0:0, notifier, , , S_AXIS_DOUT_WORDS_ACLK_delay, S_AXIS_DOUT_WORDS_TDATA_delay[17]);
    $setuphold (posedge S_AXIS_DOUT_WORDS_ACLK, negedge S_AXIS_DOUT_WORDS_TDATA[18], 0:0:0, 0:0:0, notifier, , , S_AXIS_DOUT_WORDS_ACLK_delay, S_AXIS_DOUT_WORDS_TDATA_delay[18]);
    $setuphold (posedge S_AXIS_DOUT_WORDS_ACLK, negedge S_AXIS_DOUT_WORDS_TDATA[19], 0:0:0, 0:0:0, notifier, , , S_AXIS_DOUT_WORDS_ACLK_delay, S_AXIS_DOUT_WORDS_TDATA_delay[19]);
    $setuphold (posedge S_AXIS_DOUT_WORDS_ACLK, negedge S_AXIS_DOUT_WORDS_TDATA[1], 0:0:0, 0:0:0, notifier, , , S_AXIS_DOUT_WORDS_ACLK_delay, S_AXIS_DOUT_WORDS_TDATA_delay[1]);
    $setuphold (posedge S_AXIS_DOUT_WORDS_ACLK, negedge S_AXIS_DOUT_WORDS_TDATA[20], 0:0:0, 0:0:0, notifier, , , S_AXIS_DOUT_WORDS_ACLK_delay, S_AXIS_DOUT_WORDS_TDATA_delay[20]);
    $setuphold (posedge S_AXIS_DOUT_WORDS_ACLK, negedge S_AXIS_DOUT_WORDS_TDATA[24], 0:0:0, 0:0:0, notifier, , , S_AXIS_DOUT_WORDS_ACLK_delay, S_AXIS_DOUT_WORDS_TDATA_delay[24]);
    $setuphold (posedge S_AXIS_DOUT_WORDS_ACLK, negedge S_AXIS_DOUT_WORDS_TDATA[25], 0:0:0, 0:0:0, notifier, , , S_AXIS_DOUT_WORDS_ACLK_delay, S_AXIS_DOUT_WORDS_TDATA_delay[25]);
    $setuphold (posedge S_AXIS_DOUT_WORDS_ACLK, negedge S_AXIS_DOUT_WORDS_TDATA[26], 0:0:0, 0:0:0, notifier, , , S_AXIS_DOUT_WORDS_ACLK_delay, S_AXIS_DOUT_WORDS_TDATA_delay[26]);
    $setuphold (posedge S_AXIS_DOUT_WORDS_ACLK, negedge S_AXIS_DOUT_WORDS_TDATA[27], 0:0:0, 0:0:0, notifier, , , S_AXIS_DOUT_WORDS_ACLK_delay, S_AXIS_DOUT_WORDS_TDATA_delay[27]);
    $setuphold (posedge S_AXIS_DOUT_WORDS_ACLK, negedge S_AXIS_DOUT_WORDS_TDATA[28], 0:0:0, 0:0:0, notifier, , , S_AXIS_DOUT_WORDS_ACLK_delay, S_AXIS_DOUT_WORDS_TDATA_delay[28]);
    $setuphold (posedge S_AXIS_DOUT_WORDS_ACLK, negedge S_AXIS_DOUT_WORDS_TDATA[2], 0:0:0, 0:0:0, notifier, , , S_AXIS_DOUT_WORDS_ACLK_delay, S_AXIS_DOUT_WORDS_TDATA_delay[2]);
    $setuphold (posedge S_AXIS_DOUT_WORDS_ACLK, negedge S_AXIS_DOUT_WORDS_TDATA[3], 0:0:0, 0:0:0, notifier, , , S_AXIS_DOUT_WORDS_ACLK_delay, S_AXIS_DOUT_WORDS_TDATA_delay[3]);
    $setuphold (posedge S_AXIS_DOUT_WORDS_ACLK, negedge S_AXIS_DOUT_WORDS_TDATA[4], 0:0:0, 0:0:0, notifier, , , S_AXIS_DOUT_WORDS_ACLK_delay, S_AXIS_DOUT_WORDS_TDATA_delay[4]);
    $setuphold (posedge S_AXIS_DOUT_WORDS_ACLK, negedge S_AXIS_DOUT_WORDS_TDATA[8], 0:0:0, 0:0:0, notifier, , , S_AXIS_DOUT_WORDS_ACLK_delay, S_AXIS_DOUT_WORDS_TDATA_delay[8]);
    $setuphold (posedge S_AXIS_DOUT_WORDS_ACLK, negedge S_AXIS_DOUT_WORDS_TDATA[9], 0:0:0, 0:0:0, notifier, , , S_AXIS_DOUT_WORDS_ACLK_delay, S_AXIS_DOUT_WORDS_TDATA_delay[9]);
    $setuphold (posedge S_AXIS_DOUT_WORDS_ACLK, negedge S_AXIS_DOUT_WORDS_TLAST, 0:0:0, 0:0:0, notifier, , , S_AXIS_DOUT_WORDS_ACLK_delay, S_AXIS_DOUT_WORDS_TLAST_delay);
    $setuphold (posedge S_AXIS_DOUT_WORDS_ACLK, negedge S_AXIS_DOUT_WORDS_TVALID, 0:0:0, 0:0:0, notifier, , , S_AXIS_DOUT_WORDS_ACLK_delay, S_AXIS_DOUT_WORDS_TVALID_delay);
    $setuphold (posedge S_AXIS_DOUT_WORDS_ACLK, posedge S_AXIS_DOUT_WORDS_TDATA[0], 0:0:0, 0:0:0, notifier, , , S_AXIS_DOUT_WORDS_ACLK_delay, S_AXIS_DOUT_WORDS_TDATA_delay[0]);
    $setuphold (posedge S_AXIS_DOUT_WORDS_ACLK, posedge S_AXIS_DOUT_WORDS_TDATA[10], 0:0:0, 0:0:0, notifier, , , S_AXIS_DOUT_WORDS_ACLK_delay, S_AXIS_DOUT_WORDS_TDATA_delay[10]);
    $setuphold (posedge S_AXIS_DOUT_WORDS_ACLK, posedge S_AXIS_DOUT_WORDS_TDATA[11], 0:0:0, 0:0:0, notifier, , , S_AXIS_DOUT_WORDS_ACLK_delay, S_AXIS_DOUT_WORDS_TDATA_delay[11]);
    $setuphold (posedge S_AXIS_DOUT_WORDS_ACLK, posedge S_AXIS_DOUT_WORDS_TDATA[12], 0:0:0, 0:0:0, notifier, , , S_AXIS_DOUT_WORDS_ACLK_delay, S_AXIS_DOUT_WORDS_TDATA_delay[12]);
    $setuphold (posedge S_AXIS_DOUT_WORDS_ACLK, posedge S_AXIS_DOUT_WORDS_TDATA[16], 0:0:0, 0:0:0, notifier, , , S_AXIS_DOUT_WORDS_ACLK_delay, S_AXIS_DOUT_WORDS_TDATA_delay[16]);
    $setuphold (posedge S_AXIS_DOUT_WORDS_ACLK, posedge S_AXIS_DOUT_WORDS_TDATA[17], 0:0:0, 0:0:0, notifier, , , S_AXIS_DOUT_WORDS_ACLK_delay, S_AXIS_DOUT_WORDS_TDATA_delay[17]);
    $setuphold (posedge S_AXIS_DOUT_WORDS_ACLK, posedge S_AXIS_DOUT_WORDS_TDATA[18], 0:0:0, 0:0:0, notifier, , , S_AXIS_DOUT_WORDS_ACLK_delay, S_AXIS_DOUT_WORDS_TDATA_delay[18]);
    $setuphold (posedge S_AXIS_DOUT_WORDS_ACLK, posedge S_AXIS_DOUT_WORDS_TDATA[19], 0:0:0, 0:0:0, notifier, , , S_AXIS_DOUT_WORDS_ACLK_delay, S_AXIS_DOUT_WORDS_TDATA_delay[19]);
    $setuphold (posedge S_AXIS_DOUT_WORDS_ACLK, posedge S_AXIS_DOUT_WORDS_TDATA[1], 0:0:0, 0:0:0, notifier, , , S_AXIS_DOUT_WORDS_ACLK_delay, S_AXIS_DOUT_WORDS_TDATA_delay[1]);
    $setuphold (posedge S_AXIS_DOUT_WORDS_ACLK, posedge S_AXIS_DOUT_WORDS_TDATA[20], 0:0:0, 0:0:0, notifier, , , S_AXIS_DOUT_WORDS_ACLK_delay, S_AXIS_DOUT_WORDS_TDATA_delay[20]);
    $setuphold (posedge S_AXIS_DOUT_WORDS_ACLK, posedge S_AXIS_DOUT_WORDS_TDATA[24], 0:0:0, 0:0:0, notifier, , , S_AXIS_DOUT_WORDS_ACLK_delay, S_AXIS_DOUT_WORDS_TDATA_delay[24]);
    $setuphold (posedge S_AXIS_DOUT_WORDS_ACLK, posedge S_AXIS_DOUT_WORDS_TDATA[25], 0:0:0, 0:0:0, notifier, , , S_AXIS_DOUT_WORDS_ACLK_delay, S_AXIS_DOUT_WORDS_TDATA_delay[25]);
    $setuphold (posedge S_AXIS_DOUT_WORDS_ACLK, posedge S_AXIS_DOUT_WORDS_TDATA[26], 0:0:0, 0:0:0, notifier, , , S_AXIS_DOUT_WORDS_ACLK_delay, S_AXIS_DOUT_WORDS_TDATA_delay[26]);
    $setuphold (posedge S_AXIS_DOUT_WORDS_ACLK, posedge S_AXIS_DOUT_WORDS_TDATA[27], 0:0:0, 0:0:0, notifier, , , S_AXIS_DOUT_WORDS_ACLK_delay, S_AXIS_DOUT_WORDS_TDATA_delay[27]);
    $setuphold (posedge S_AXIS_DOUT_WORDS_ACLK, posedge S_AXIS_DOUT_WORDS_TDATA[28], 0:0:0, 0:0:0, notifier, , , S_AXIS_DOUT_WORDS_ACLK_delay, S_AXIS_DOUT_WORDS_TDATA_delay[28]);
    $setuphold (posedge S_AXIS_DOUT_WORDS_ACLK, posedge S_AXIS_DOUT_WORDS_TDATA[2], 0:0:0, 0:0:0, notifier, , , S_AXIS_DOUT_WORDS_ACLK_delay, S_AXIS_DOUT_WORDS_TDATA_delay[2]);
    $setuphold (posedge S_AXIS_DOUT_WORDS_ACLK, posedge S_AXIS_DOUT_WORDS_TDATA[3], 0:0:0, 0:0:0, notifier, , , S_AXIS_DOUT_WORDS_ACLK_delay, S_AXIS_DOUT_WORDS_TDATA_delay[3]);
    $setuphold (posedge S_AXIS_DOUT_WORDS_ACLK, posedge S_AXIS_DOUT_WORDS_TDATA[4], 0:0:0, 0:0:0, notifier, , , S_AXIS_DOUT_WORDS_ACLK_delay, S_AXIS_DOUT_WORDS_TDATA_delay[4]);
    $setuphold (posedge S_AXIS_DOUT_WORDS_ACLK, posedge S_AXIS_DOUT_WORDS_TDATA[8], 0:0:0, 0:0:0, notifier, , , S_AXIS_DOUT_WORDS_ACLK_delay, S_AXIS_DOUT_WORDS_TDATA_delay[8]);
    $setuphold (posedge S_AXIS_DOUT_WORDS_ACLK, posedge S_AXIS_DOUT_WORDS_TDATA[9], 0:0:0, 0:0:0, notifier, , , S_AXIS_DOUT_WORDS_ACLK_delay, S_AXIS_DOUT_WORDS_TDATA_delay[9]);
    $setuphold (posedge S_AXIS_DOUT_WORDS_ACLK, posedge S_AXIS_DOUT_WORDS_TLAST, 0:0:0, 0:0:0, notifier, , , S_AXIS_DOUT_WORDS_ACLK_delay, S_AXIS_DOUT_WORDS_TLAST_delay);
    $setuphold (posedge S_AXIS_DOUT_WORDS_ACLK, posedge S_AXIS_DOUT_WORDS_TVALID, 0:0:0, 0:0:0, notifier, , , S_AXIS_DOUT_WORDS_ACLK_delay, S_AXIS_DOUT_WORDS_TVALID_delay);
    $setuphold (posedge S_AXI_ACLK, negedge S_AXI_ARADDR[10], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_ARADDR_delay[10]);
    $setuphold (posedge S_AXI_ACLK, negedge S_AXI_ARADDR[11], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_ARADDR_delay[11]);
    $setuphold (posedge S_AXI_ACLK, negedge S_AXI_ARADDR[12], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_ARADDR_delay[12]);
    $setuphold (posedge S_AXI_ACLK, negedge S_AXI_ARADDR[13], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_ARADDR_delay[13]);
    $setuphold (posedge S_AXI_ACLK, negedge S_AXI_ARADDR[14], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_ARADDR_delay[14]);
    $setuphold (posedge S_AXI_ACLK, negedge S_AXI_ARADDR[15], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_ARADDR_delay[15]);
    $setuphold (posedge S_AXI_ACLK, negedge S_AXI_ARADDR[16], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_ARADDR_delay[16]);
    $setuphold (posedge S_AXI_ACLK, negedge S_AXI_ARADDR[17], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_ARADDR_delay[17]);
    $setuphold (posedge S_AXI_ACLK, negedge S_AXI_ARADDR[2], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_ARADDR_delay[2]);
    $setuphold (posedge S_AXI_ACLK, negedge S_AXI_ARADDR[3], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_ARADDR_delay[3]);
    $setuphold (posedge S_AXI_ACLK, negedge S_AXI_ARADDR[4], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_ARADDR_delay[4]);
    $setuphold (posedge S_AXI_ACLK, negedge S_AXI_ARADDR[5], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_ARADDR_delay[5]);
    $setuphold (posedge S_AXI_ACLK, negedge S_AXI_ARADDR[6], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_ARADDR_delay[6]);
    $setuphold (posedge S_AXI_ACLK, negedge S_AXI_ARADDR[7], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_ARADDR_delay[7]);
    $setuphold (posedge S_AXI_ACLK, negedge S_AXI_ARADDR[8], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_ARADDR_delay[8]);
    $setuphold (posedge S_AXI_ACLK, negedge S_AXI_ARADDR[9], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_ARADDR_delay[9]);
    $setuphold (posedge S_AXI_ACLK, negedge S_AXI_ARVALID, 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_ARVALID_delay);
    $setuphold (posedge S_AXI_ACLK, negedge S_AXI_AWADDR[10], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_AWADDR_delay[10]);
    $setuphold (posedge S_AXI_ACLK, negedge S_AXI_AWADDR[11], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_AWADDR_delay[11]);
    $setuphold (posedge S_AXI_ACLK, negedge S_AXI_AWADDR[12], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_AWADDR_delay[12]);
    $setuphold (posedge S_AXI_ACLK, negedge S_AXI_AWADDR[13], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_AWADDR_delay[13]);
    $setuphold (posedge S_AXI_ACLK, negedge S_AXI_AWADDR[14], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_AWADDR_delay[14]);
    $setuphold (posedge S_AXI_ACLK, negedge S_AXI_AWADDR[15], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_AWADDR_delay[15]);
    $setuphold (posedge S_AXI_ACLK, negedge S_AXI_AWADDR[16], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_AWADDR_delay[16]);
    $setuphold (posedge S_AXI_ACLK, negedge S_AXI_AWADDR[17], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_AWADDR_delay[17]);
    $setuphold (posedge S_AXI_ACLK, negedge S_AXI_AWADDR[2], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_AWADDR_delay[2]);
    $setuphold (posedge S_AXI_ACLK, negedge S_AXI_AWADDR[3], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_AWADDR_delay[3]);
    $setuphold (posedge S_AXI_ACLK, negedge S_AXI_AWADDR[4], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_AWADDR_delay[4]);
    $setuphold (posedge S_AXI_ACLK, negedge S_AXI_AWADDR[5], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_AWADDR_delay[5]);
    $setuphold (posedge S_AXI_ACLK, negedge S_AXI_AWADDR[6], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_AWADDR_delay[6]);
    $setuphold (posedge S_AXI_ACLK, negedge S_AXI_AWADDR[7], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_AWADDR_delay[7]);
    $setuphold (posedge S_AXI_ACLK, negedge S_AXI_AWADDR[8], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_AWADDR_delay[8]);
    $setuphold (posedge S_AXI_ACLK, negedge S_AXI_AWADDR[9], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_AWADDR_delay[9]);
    $setuphold (posedge S_AXI_ACLK, negedge S_AXI_AWVALID, 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_AWVALID_delay);
    $setuphold (posedge S_AXI_ACLK, negedge S_AXI_BREADY, 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_BREADY_delay);
    $setuphold (posedge S_AXI_ACLK, negedge S_AXI_RREADY, 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_RREADY_delay);
    $setuphold (posedge S_AXI_ACLK, negedge S_AXI_WDATA[0], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_WDATA_delay[0]);
    $setuphold (posedge S_AXI_ACLK, negedge S_AXI_WDATA[10], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_WDATA_delay[10]);
    $setuphold (posedge S_AXI_ACLK, negedge S_AXI_WDATA[11], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_WDATA_delay[11]);
    $setuphold (posedge S_AXI_ACLK, negedge S_AXI_WDATA[12], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_WDATA_delay[12]);
    $setuphold (posedge S_AXI_ACLK, negedge S_AXI_WDATA[13], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_WDATA_delay[13]);
    $setuphold (posedge S_AXI_ACLK, negedge S_AXI_WDATA[14], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_WDATA_delay[14]);
    $setuphold (posedge S_AXI_ACLK, negedge S_AXI_WDATA[15], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_WDATA_delay[15]);
    $setuphold (posedge S_AXI_ACLK, negedge S_AXI_WDATA[16], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_WDATA_delay[16]);
    $setuphold (posedge S_AXI_ACLK, negedge S_AXI_WDATA[17], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_WDATA_delay[17]);
    $setuphold (posedge S_AXI_ACLK, negedge S_AXI_WDATA[18], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_WDATA_delay[18]);
    $setuphold (posedge S_AXI_ACLK, negedge S_AXI_WDATA[19], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_WDATA_delay[19]);
    $setuphold (posedge S_AXI_ACLK, negedge S_AXI_WDATA[1], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_WDATA_delay[1]);
    $setuphold (posedge S_AXI_ACLK, negedge S_AXI_WDATA[20], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_WDATA_delay[20]);
    $setuphold (posedge S_AXI_ACLK, negedge S_AXI_WDATA[21], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_WDATA_delay[21]);
    $setuphold (posedge S_AXI_ACLK, negedge S_AXI_WDATA[22], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_WDATA_delay[22]);
    $setuphold (posedge S_AXI_ACLK, negedge S_AXI_WDATA[23], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_WDATA_delay[23]);
    $setuphold (posedge S_AXI_ACLK, negedge S_AXI_WDATA[24], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_WDATA_delay[24]);
    $setuphold (posedge S_AXI_ACLK, negedge S_AXI_WDATA[25], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_WDATA_delay[25]);
    $setuphold (posedge S_AXI_ACLK, negedge S_AXI_WDATA[26], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_WDATA_delay[26]);
    $setuphold (posedge S_AXI_ACLK, negedge S_AXI_WDATA[27], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_WDATA_delay[27]);
    $setuphold (posedge S_AXI_ACLK, negedge S_AXI_WDATA[28], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_WDATA_delay[28]);
    $setuphold (posedge S_AXI_ACLK, negedge S_AXI_WDATA[29], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_WDATA_delay[29]);
    $setuphold (posedge S_AXI_ACLK, negedge S_AXI_WDATA[2], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_WDATA_delay[2]);
    $setuphold (posedge S_AXI_ACLK, negedge S_AXI_WDATA[30], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_WDATA_delay[30]);
    $setuphold (posedge S_AXI_ACLK, negedge S_AXI_WDATA[31], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_WDATA_delay[31]);
    $setuphold (posedge S_AXI_ACLK, negedge S_AXI_WDATA[3], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_WDATA_delay[3]);
    $setuphold (posedge S_AXI_ACLK, negedge S_AXI_WDATA[4], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_WDATA_delay[4]);
    $setuphold (posedge S_AXI_ACLK, negedge S_AXI_WDATA[5], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_WDATA_delay[5]);
    $setuphold (posedge S_AXI_ACLK, negedge S_AXI_WDATA[6], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_WDATA_delay[6]);
    $setuphold (posedge S_AXI_ACLK, negedge S_AXI_WDATA[7], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_WDATA_delay[7]);
    $setuphold (posedge S_AXI_ACLK, negedge S_AXI_WDATA[8], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_WDATA_delay[8]);
    $setuphold (posedge S_AXI_ACLK, negedge S_AXI_WDATA[9], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_WDATA_delay[9]);
    $setuphold (posedge S_AXI_ACLK, negedge S_AXI_WVALID, 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_WVALID_delay);
    $setuphold (posedge S_AXI_ACLK, posedge S_AXI_ARADDR[10], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_ARADDR_delay[10]);
    $setuphold (posedge S_AXI_ACLK, posedge S_AXI_ARADDR[11], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_ARADDR_delay[11]);
    $setuphold (posedge S_AXI_ACLK, posedge S_AXI_ARADDR[12], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_ARADDR_delay[12]);
    $setuphold (posedge S_AXI_ACLK, posedge S_AXI_ARADDR[13], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_ARADDR_delay[13]);
    $setuphold (posedge S_AXI_ACLK, posedge S_AXI_ARADDR[14], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_ARADDR_delay[14]);
    $setuphold (posedge S_AXI_ACLK, posedge S_AXI_ARADDR[15], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_ARADDR_delay[15]);
    $setuphold (posedge S_AXI_ACLK, posedge S_AXI_ARADDR[16], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_ARADDR_delay[16]);
    $setuphold (posedge S_AXI_ACLK, posedge S_AXI_ARADDR[17], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_ARADDR_delay[17]);
    $setuphold (posedge S_AXI_ACLK, posedge S_AXI_ARADDR[2], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_ARADDR_delay[2]);
    $setuphold (posedge S_AXI_ACLK, posedge S_AXI_ARADDR[3], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_ARADDR_delay[3]);
    $setuphold (posedge S_AXI_ACLK, posedge S_AXI_ARADDR[4], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_ARADDR_delay[4]);
    $setuphold (posedge S_AXI_ACLK, posedge S_AXI_ARADDR[5], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_ARADDR_delay[5]);
    $setuphold (posedge S_AXI_ACLK, posedge S_AXI_ARADDR[6], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_ARADDR_delay[6]);
    $setuphold (posedge S_AXI_ACLK, posedge S_AXI_ARADDR[7], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_ARADDR_delay[7]);
    $setuphold (posedge S_AXI_ACLK, posedge S_AXI_ARADDR[8], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_ARADDR_delay[8]);
    $setuphold (posedge S_AXI_ACLK, posedge S_AXI_ARADDR[9], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_ARADDR_delay[9]);
    $setuphold (posedge S_AXI_ACLK, posedge S_AXI_ARVALID, 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_ARVALID_delay);
    $setuphold (posedge S_AXI_ACLK, posedge S_AXI_AWADDR[10], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_AWADDR_delay[10]);
    $setuphold (posedge S_AXI_ACLK, posedge S_AXI_AWADDR[11], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_AWADDR_delay[11]);
    $setuphold (posedge S_AXI_ACLK, posedge S_AXI_AWADDR[12], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_AWADDR_delay[12]);
    $setuphold (posedge S_AXI_ACLK, posedge S_AXI_AWADDR[13], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_AWADDR_delay[13]);
    $setuphold (posedge S_AXI_ACLK, posedge S_AXI_AWADDR[14], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_AWADDR_delay[14]);
    $setuphold (posedge S_AXI_ACLK, posedge S_AXI_AWADDR[15], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_AWADDR_delay[15]);
    $setuphold (posedge S_AXI_ACLK, posedge S_AXI_AWADDR[16], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_AWADDR_delay[16]);
    $setuphold (posedge S_AXI_ACLK, posedge S_AXI_AWADDR[17], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_AWADDR_delay[17]);
    $setuphold (posedge S_AXI_ACLK, posedge S_AXI_AWADDR[2], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_AWADDR_delay[2]);
    $setuphold (posedge S_AXI_ACLK, posedge S_AXI_AWADDR[3], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_AWADDR_delay[3]);
    $setuphold (posedge S_AXI_ACLK, posedge S_AXI_AWADDR[4], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_AWADDR_delay[4]);
    $setuphold (posedge S_AXI_ACLK, posedge S_AXI_AWADDR[5], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_AWADDR_delay[5]);
    $setuphold (posedge S_AXI_ACLK, posedge S_AXI_AWADDR[6], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_AWADDR_delay[6]);
    $setuphold (posedge S_AXI_ACLK, posedge S_AXI_AWADDR[7], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_AWADDR_delay[7]);
    $setuphold (posedge S_AXI_ACLK, posedge S_AXI_AWADDR[8], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_AWADDR_delay[8]);
    $setuphold (posedge S_AXI_ACLK, posedge S_AXI_AWADDR[9], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_AWADDR_delay[9]);
    $setuphold (posedge S_AXI_ACLK, posedge S_AXI_AWVALID, 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_AWVALID_delay);
    $setuphold (posedge S_AXI_ACLK, posedge S_AXI_BREADY, 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_BREADY_delay);
    $setuphold (posedge S_AXI_ACLK, posedge S_AXI_RREADY, 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_RREADY_delay);
    $setuphold (posedge S_AXI_ACLK, posedge S_AXI_WDATA[0], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_WDATA_delay[0]);
    $setuphold (posedge S_AXI_ACLK, posedge S_AXI_WDATA[10], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_WDATA_delay[10]);
    $setuphold (posedge S_AXI_ACLK, posedge S_AXI_WDATA[11], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_WDATA_delay[11]);
    $setuphold (posedge S_AXI_ACLK, posedge S_AXI_WDATA[12], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_WDATA_delay[12]);
    $setuphold (posedge S_AXI_ACLK, posedge S_AXI_WDATA[13], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_WDATA_delay[13]);
    $setuphold (posedge S_AXI_ACLK, posedge S_AXI_WDATA[14], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_WDATA_delay[14]);
    $setuphold (posedge S_AXI_ACLK, posedge S_AXI_WDATA[15], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_WDATA_delay[15]);
    $setuphold (posedge S_AXI_ACLK, posedge S_AXI_WDATA[16], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_WDATA_delay[16]);
    $setuphold (posedge S_AXI_ACLK, posedge S_AXI_WDATA[17], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_WDATA_delay[17]);
    $setuphold (posedge S_AXI_ACLK, posedge S_AXI_WDATA[18], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_WDATA_delay[18]);
    $setuphold (posedge S_AXI_ACLK, posedge S_AXI_WDATA[19], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_WDATA_delay[19]);
    $setuphold (posedge S_AXI_ACLK, posedge S_AXI_WDATA[1], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_WDATA_delay[1]);
    $setuphold (posedge S_AXI_ACLK, posedge S_AXI_WDATA[20], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_WDATA_delay[20]);
    $setuphold (posedge S_AXI_ACLK, posedge S_AXI_WDATA[21], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_WDATA_delay[21]);
    $setuphold (posedge S_AXI_ACLK, posedge S_AXI_WDATA[22], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_WDATA_delay[22]);
    $setuphold (posedge S_AXI_ACLK, posedge S_AXI_WDATA[23], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_WDATA_delay[23]);
    $setuphold (posedge S_AXI_ACLK, posedge S_AXI_WDATA[24], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_WDATA_delay[24]);
    $setuphold (posedge S_AXI_ACLK, posedge S_AXI_WDATA[25], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_WDATA_delay[25]);
    $setuphold (posedge S_AXI_ACLK, posedge S_AXI_WDATA[26], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_WDATA_delay[26]);
    $setuphold (posedge S_AXI_ACLK, posedge S_AXI_WDATA[27], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_WDATA_delay[27]);
    $setuphold (posedge S_AXI_ACLK, posedge S_AXI_WDATA[28], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_WDATA_delay[28]);
    $setuphold (posedge S_AXI_ACLK, posedge S_AXI_WDATA[29], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_WDATA_delay[29]);
    $setuphold (posedge S_AXI_ACLK, posedge S_AXI_WDATA[2], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_WDATA_delay[2]);
    $setuphold (posedge S_AXI_ACLK, posedge S_AXI_WDATA[30], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_WDATA_delay[30]);
    $setuphold (posedge S_AXI_ACLK, posedge S_AXI_WDATA[31], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_WDATA_delay[31]);
    $setuphold (posedge S_AXI_ACLK, posedge S_AXI_WDATA[3], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_WDATA_delay[3]);
    $setuphold (posedge S_AXI_ACLK, posedge S_AXI_WDATA[4], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_WDATA_delay[4]);
    $setuphold (posedge S_AXI_ACLK, posedge S_AXI_WDATA[5], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_WDATA_delay[5]);
    $setuphold (posedge S_AXI_ACLK, posedge S_AXI_WDATA[6], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_WDATA_delay[6]);
    $setuphold (posedge S_AXI_ACLK, posedge S_AXI_WDATA[7], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_WDATA_delay[7]);
    $setuphold (posedge S_AXI_ACLK, posedge S_AXI_WDATA[8], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_WDATA_delay[8]);
    $setuphold (posedge S_AXI_ACLK, posedge S_AXI_WDATA[9], 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_WDATA_delay[9]);
    $setuphold (posedge S_AXI_ACLK, posedge S_AXI_WVALID, 0:0:0, 0:0:0, notifier, , , S_AXI_ACLK_delay, S_AXI_WVALID_delay);
    $width (negedge CORE_CLK, 0:0:0, 0, notifier);
    $width (negedge M_AXIS_DOUT_ACLK, 0:0:0, 0, notifier);
    $width (negedge M_AXIS_STATUS_ACLK, 0:0:0, 0, notifier);
    $width (negedge S_AXIS_CTRL_ACLK, 0:0:0, 0, notifier);
    $width (negedge S_AXIS_DIN_ACLK, 0:0:0, 0, notifier);
    $width (negedge S_AXIS_DIN_WORDS_ACLK, 0:0:0, 0, notifier);
    $width (negedge S_AXIS_DOUT_WORDS_ACLK, 0:0:0, 0, notifier);
    $width (negedge S_AXI_ACLK, 0:0:0, 0, notifier);
    $width (posedge CORE_CLK, 0:0:0, 0, notifier);
    $width (posedge M_AXIS_DOUT_ACLK, 0:0:0, 0, notifier);
    $width (posedge M_AXIS_STATUS_ACLK, 0:0:0, 0, notifier);
    $width (posedge S_AXIS_CTRL_ACLK, 0:0:0, 0, notifier);
    $width (posedge S_AXIS_DIN_ACLK, 0:0:0, 0, notifier);
    $width (posedge S_AXIS_DIN_WORDS_ACLK, 0:0:0, 0, notifier);
    $width (posedge S_AXIS_DOUT_WORDS_ACLK, 0:0:0, 0, notifier);
    $width (posedge S_AXI_ACLK, 0:0:0, 0, notifier);
`endif
    specparam PATHPULSE$ = 0;
  endspecify
`endif
endmodule