module sim;
  // VCD Dump
  //initial begin
  //  $dumpfile("run.vcd");
  //  $dumpvars;
  //end
  // Generate Clock
  reg clk = 1'b0;
  always #5 clk = ~clk;
  // MulDiv Unit
  reg   [1:0] verbose;
  reg   [2:0] src_msg_fn;
  reg  [31:0] nmults;
  reg  [31:0] src_msg_a;
  reg  [31:0] src_msg_b;
  reg         src_val = 1'b0;
  wire        src_rdy;
  //wire [63:0] sink_msg;
  wire [31:0] sink_msg;
  wire        sink_val;
  wire        sink_rdy = 1'b1; // Always ready to accept result
  wire        muldivreq_go  = src_val  && src_rdy;
  wire        muldivresp_go = sink_val && sink_rdy;
  reg reset = 1'b1;
  imuldiv_IntMulVariable imul
  (
    .clk                (clk),
    .reset              (reset),
    .mulreq_msg_a       (src_msg_a),
    .mulreq_msg_b       (src_msg_b),
    .mulreq_val         (src_val),
    .mulreq_rdy         (src_rdy),
    .mulresp_msg_result (sink_msg),
    .mulresp_val        (sink_val),
    .mulresp_rdy        (sink_rdy)
  );
  // Test Vectors
  integer idx;
  reg [31:0] in0[999:0];
  reg [31:0] in1[999:0];
  reg [31:0] out[999:0];
  initial begin
    idx = 0;
    in0[  0]=32'h67f34f6d; in1[  0]=32'h24c617a0; out[  0]=32'h96826f20;
    in0[  1]=32'hb5d9ed18; in1[  1]=32'h7eb389c5; out[  1]=32'h285d4b78;
    in0[  2]=32'h5786f1db; in1[  2]=32'h435acae1; out[  2]=32'hc06f5f7b;
    in0[  3]=32'h70047e7d; in1[  3]=32'hff3e1308; out[  3]=32'hfacd3ae8;
    in0[  4]=32'h5530cbf5; in1[  4]=32'hc4984d96; out[  4]=32'h4568328e;
    in0[  5]=32'h34147951; in1[  5]=32'hf65b9385; out[  5]=32'hc6178a15;
    in0[  6]=32'h75174485; in1[  6]=32'h2920e6bc; out[  6]=32'hc245cfac;
    in0[  7]=32'h26171439; in1[  7]=32'h8c871861; out[  7]=32'h6eb30199;
    in0[  8]=32'h117cb918; in1[  8]=32'h2c809d62; out[  8]=32'hdb429330;
    in0[  9]=32'h4164f86c; in1[  9]=32'h7995f109; out[  9]=32'hfd4667cc;
    in0[ 10]=32'hf2c40f62; in1[ 10]=32'h897e310f; out[ 10]=32'hc4aaa8be;
    in0[ 11]=32'h610082d8; in1[ 11]=32'hb6fdc399; out[ 11]=32'h3c70bb18;
    in0[ 12]=32'hfdb3bc12; in1[ 12]=32'hbb9dd55e; out[ 12]=32'h3084089c;
    in0[ 13]=32'h1da3dd7e; in1[ 13]=32'h89ec653a; out[ 13]=32'hfbaae48c;
    in0[ 14]=32'hcc0d8e74; in1[ 14]=32'h9b30bcb3; out[ 14]=32'h93d7cb1c;
    in0[ 15]=32'ha37d20a5; in1[ 15]=32'hf5de555a; out[ 15]=32'h3dea4302;
    in0[ 16]=32'h892ea376; in1[ 16]=32'had1c78fd; out[ 16]=32'h0e9edb9e;
    in0[ 17]=32'he1d01c91; in1[ 17]=32'h3793ff36; out[ 17]=32'h7c9d7596;
    in0[ 18]=32'he5867c11; in1[ 18]=32'ha0e0ee12; out[ 18]=32'h59ac8732;
    in0[ 19]=32'hd119415a; in1[ 19]=32'h906fa0b0; out[ 19]=32'h803b2de0;
    in0[ 20]=32'ha52d20c0; in1[ 20]=32'hb70ab4a1; out[ 20]=32'h23e898c0;
    in0[ 21]=32'h988bebd1; in1[ 21]=32'h7365b610; out[ 21]=32'heeda5310;
    in0[ 22]=32'hf5412b23; in1[ 22]=32'hdbf52a72; out[ 22]=32'h2197f396;
    in0[ 23]=32'he16f4ef6; in1[ 23]=32'h761bd7f5; out[ 23]=32'hf2c92b6e;
    in0[ 24]=32'h7b85eeb6; in1[ 24]=32'hac28c326; out[ 24]=32'hef261104;
    in0[ 25]=32'h3be0f2e1; in1[ 25]=32'hfcf48677; out[ 25]=32'h8f26ac97;
    in0[ 26]=32'h85ec31ac; in1[ 26]=32'h5a4dd21e; out[ 26]=32'hdb28ea28;
    in0[ 27]=32'h47d041ec; in1[ 27]=32'h74df3ccc; out[ 27]=32'h65fbd810;
    in0[ 28]=32'h4048c934; in1[ 28]=32'h49827b21; out[ 28]=32'h4275ebb4;
    in0[ 29]=32'h49469987; in1[ 29]=32'hd87f15d7; out[ 29]=32'h66dc0361;
    in0[ 30]=32'hc981f522; in1[ 30]=32'h8ac94675; out[ 30]=32'h6d1e548a;
    in0[ 31]=32'h093a1e26; in1[ 31]=32'hd677487d; out[ 31]=32'ha185688e;
    in0[ 32]=32'haf27aab1; in1[ 32]=32'h931b1789; out[ 32]=32'hf03b3fb9;
    in0[ 33]=32'he4981875; in1[ 33]=32'h004ae4cf; out[ 33]=32'h5e95fa9b;
    in0[ 34]=32'hbbea7acf; in1[ 34]=32'hb32d6451; out[ 34]=32'h608cb77f;
    in0[ 35]=32'hc3a0da02; in1[ 35]=32'hf99ff344; out[ 35]=32'hfee7ce88;
    in0[ 36]=32'h4c9d8ecb; in1[ 36]=32'hfa56f325; out[ 36]=32'hd7825457;
    in0[ 37]=32'hec8d9cc4; in1[ 37]=32'hb1c15a91; out[ 37]=32'h7916b304;
    in0[ 38]=32'he9400bcb; in1[ 38]=32'hcefa10a8; out[ 38]=32'hf1026d38;
    in0[ 39]=32'h8482ecc4; in1[ 39]=32'h0d4ebc72; out[ 39]=32'h3fe55f48;
    in0[ 40]=32'h0a15e96b; in1[ 40]=32'h203af540; out[ 40]=32'hc01bc1c0;
    in0[ 41]=32'ha4653582; in1[ 41]=32'hdae36b48; out[ 41]=32'hb01a6290;
    in0[ 42]=32'h08b9ea64; in1[ 42]=32'h5b8f48cc; out[ 42]=32'hb7eee7b0;
    in0[ 43]=32'h419c1ce8; in1[ 43]=32'ha69a4650; out[ 43]=32'h04407880;
    in0[ 44]=32'h575e10f4; in1[ 44]=32'habc8117a; out[ 44]=32'h1c944848;
    in0[ 45]=32'h75c41c0d; in1[ 45]=32'h596944c7; out[ 45]=32'ha93a421b;
    in0[ 46]=32'hec0ffb99; in1[ 46]=32'h1db25718; out[ 46]=32'hd5629558;
    in0[ 47]=32'h6064f66a; in1[ 47]=32'hca550c64; out[ 47]=32'hd82f3968;
    in0[ 48]=32'h10754117; in1[ 48]=32'hcaec691b; out[ 48]=32'hfb444c6d;
    in0[ 49]=32'h74cadc3d; in1[ 49]=32'h8db4a155; out[ 49]=32'hcfc17d41;
    in0[ 50]=32'h371d921d; in1[ 50]=32'h3d616d79; out[ 50]=32'hea2d68b5;
    in0[ 51]=32'h6e841170; in1[ 51]=32'he57ead4b; out[ 51]=32'h6599cbd0;
    in0[ 52]=32'h6464ffd4; in1[ 52]=32'h692633d0; out[ 52]=32'h9e7f1840;
    in0[ 53]=32'h0f2356e6; in1[ 53]=32'h592afec1; out[ 53]=32'hb198b766;
    in0[ 54]=32'h9c7f213a; in1[ 54]=32'hd10fabf3; out[ 54]=32'hc444480e;
    in0[ 55]=32'hb45d0921; in1[ 55]=32'h67f680ec; out[ 55]=32'hd70aea6c;
    in0[ 56]=32'h6331711a; in1[ 56]=32'hd89f5d10; out[ 56]=32'h585383a0;
    in0[ 57]=32'h2dae0b84; in1[ 57]=32'h436b815b; out[ 57]=32'h4cd79bec;
    in0[ 58]=32'hcefbd30f; in1[ 58]=32'hf8c9e39f; out[ 58]=32'h19556351;
    in0[ 59]=32'h432d54cc; in1[ 59]=32'hfb5e1791; out[ 59]=32'h46335b8c;
    in0[ 60]=32'h7249d9b7; in1[ 60]=32'he6ae8883; out[ 60]=32'h1bd5a0a5;
    in0[ 61]=32'hd1a06415; in1[ 61]=32'hc530a942; out[ 61]=32'hda5baa6a;
    in0[ 62]=32'h1f6e422d; in1[ 62]=32'h08fc6c4e; out[ 62]=32'ha3cf25b6;
    in0[ 63]=32'h91896038; in1[ 63]=32'hb107b9a4; out[ 63]=32'hdc121be0;
    in0[ 64]=32'h3f79e4fd; in1[ 64]=32'h1534b813; out[ 64]=32'h9705d6c7;
    in0[ 65]=32'hee3ac762; in1[ 65]=32'h0385a7d9; out[ 65]=32'h03cdf012;
    in0[ 66]=32'h0baffde4; in1[ 66]=32'h55d6f147; out[ 66]=32'hdc6b0e3c;
    in0[ 67]=32'h6ad2a566; in1[ 67]=32'hc9b12c54; out[ 67]=32'hb311cd78;
    in0[ 68]=32'ha518fa06; in1[ 68]=32'hea8216c2; out[ 68]=32'hb575fc8c;
    in0[ 69]=32'h5e87c367; in1[ 69]=32'h79fdd610; out[ 69]=32'h319f5070;
    in0[ 70]=32'h7e3a298b; in1[ 70]=32'h66d0b415; out[ 70]=32'h62eb2467;
    in0[ 71]=32'h50d7d8ed; in1[ 71]=32'h84485084; out[ 71]=32'h59bdea34;
    in0[ 72]=32'h453530fc; in1[ 72]=32'h24c557ea; out[ 72]=32'h78306a58;
    in0[ 73]=32'h829e2190; in1[ 73]=32'hff9f7faf; out[ 73]=32'h052f6170;
    in0[ 74]=32'h38a8b121; in1[ 74]=32'hc5506a3a; out[ 74]=32'h6edfcb7a;
    in0[ 75]=32'hed137b52; in1[ 75]=32'h2f30695a; out[ 75]=32'h83cdfcd4;
    in0[ 76]=32'ha524c9bd; in1[ 76]=32'h4fd2fae2; out[ 76]=32'h8786aada;
    in0[ 77]=32'he3ef9ace; in1[ 77]=32'h6e2ee860; out[ 77]=32'hf328bd40;
    in0[ 78]=32'hbe1a989b; in1[ 78]=32'h908efb5e; out[ 78]=32'hb75e01ea;
    in0[ 79]=32'h83f1d8dd; in1[ 79]=32'h01cfe0f4; out[ 79]=32'h97f712a4;
    in0[ 80]=32'hbb9a2450; in1[ 80]=32'h482efb5b; out[ 80]=32'hd7c55870;
    in0[ 81]=32'he6c0a9d6; in1[ 81]=32'h8b0481f7; out[ 81]=32'h92d0b37a;
    in0[ 82]=32'h3562690a; in1[ 82]=32'h032471f1; out[ 82]=32'h956a4c6a;
    in0[ 83]=32'hd0ff2e60; in1[ 83]=32'heff8f177; out[ 83]=32'hee46eea0;
    in0[ 84]=32'hb4b16f6e; in1[ 84]=32'h12442bcf; out[ 84]=32'h3e6893f2;
    in0[ 85]=32'h1c6ffba1; in1[ 85]=32'h713c6b02; out[ 85]=32'h11c84242;
    in0[ 86]=32'h657c6487; in1[ 86]=32'h7fc1e97e; out[ 86]=32'hed7f5972;
    in0[ 87]=32'h611488f2; in1[ 87]=32'he8948161; out[ 87]=32'h9db1d5b2;
    in0[ 88]=32'h0b2dc798; in1[ 88]=32'h2efbd35e; out[ 88]=32'hd85991d0;
    in0[ 89]=32'h976b00b2; in1[ 89]=32'hffa8326b; out[ 89]=32'hf2ac0e66;
    in0[ 90]=32'h88a725b6; in1[ 90]=32'h1912dbf3; out[ 90]=32'h20b77dc2;
    in0[ 91]=32'hcf4bb68f; in1[ 91]=32'h085b63b0; out[ 91]=32'h287bcf50;
    in0[ 92]=32'h1965d1cb; in1[ 92]=32'h819cb1cb; out[ 92]=32'hac7eb6f9;
    in0[ 93]=32'hc0ff188b; in1[ 93]=32'h0e04a247; out[ 93]=32'hf073c48d;
    in0[ 94]=32'h7ea2e156; in1[ 94]=32'hb133fdca; out[ 94]=32'h3f59cbdc;
    in0[ 95]=32'h7c5433dd; in1[ 95]=32'h9880bdc7; out[ 95]=32'hf63e79cb;
    in0[ 96]=32'h4c04c579; in1[ 96]=32'h8c835b5e; out[ 96]=32'hd4dd856e;
    in0[ 97]=32'hbc7af287; in1[ 97]=32'hf25842a4; out[ 97]=32'h6db22c7c;
    in0[ 98]=32'he5bb2796; in1[ 98]=32'hd67b3899; out[ 98]=32'ha69578a6;
    in0[ 99]=32'h3b3f1b45; in1[ 99]=32'hf0591df6; out[ 99]=32'h3fb8054e;
    in0[100]=32'hef6965de; in1[100]=32'hcc392eac; out[100]=32'h618c5528;
    in0[101]=32'h75db7464; in1[101]=32'hde732e12; out[101]=32'hb9442708;
    in0[102]=32'h3ceb3472; in1[102]=32'h7da99e66; out[102]=32'hb957416c;
    in0[103]=32'h8b95d7fb; in1[103]=32'h4d749456; out[103]=32'he1efaa52;
    in0[104]=32'hb884bbf4; in1[104]=32'h43967e77; out[104]=32'h172d766c;
    in0[105]=32'hee9c1a25; in1[105]=32'h434b6b99; out[105]=32'h3210171d;
    in0[106]=32'h4dac2709; in1[106]=32'h17ce8672; out[106]=32'heb561802;
    in0[107]=32'h3605bc3e; in1[107]=32'h701fb675; out[107]=32'haff51c56;
    in0[108]=32'h93f73d6f; in1[108]=32'h2119bc20; out[108]=32'h5edc31e0;
    in0[109]=32'he418c577; in1[109]=32'h81e9baec; out[109]=32'hf69d7fb4;
    in0[110]=32'h490bf0e3; in1[110]=32'h768b1f88; out[110]=32'hadc47598;
    in0[111]=32'h0b0f0343; in1[111]=32'h10a2d939; out[111]=32'h708184eb;
    in0[112]=32'hd5bafb2f; in1[112]=32'h777d0f74; out[112]=32'h4c64924c;
    in0[113]=32'h64825c2a; in1[113]=32'hec544896; out[113]=32'h8415d09c;
    in0[114]=32'h6e3b29ea; in1[114]=32'h4fb87322; out[114]=32'h8ddfaf14;
    in0[115]=32'h450c98d8; in1[115]=32'h07b2b48b; out[115]=32'h877edd48;
    in0[116]=32'hbe4d28de; in1[116]=32'hfbe99445; out[116]=32'hc27a5bd6;
    in0[117]=32'ha38665e6; in1[117]=32'hd2b26222; out[117]=32'hb0c7948c;
    in0[118]=32'hfff19cc1; in1[118]=32'h1f642cfa; out[118]=32'h1348407a;
    in0[119]=32'h1ea06a92; in1[119]=32'h8cf6caa4; out[119]=32'h73277988;
    in0[120]=32'hab045171; in1[120]=32'hcd50ae58; out[120]=32'ha926ccd8;
    in0[121]=32'hb24505ff; in1[121]=32'hc5a5bec7; out[121]=32'he675eb39;
    in0[122]=32'h48b02005; in1[122]=32'hd4f6ac00; out[122]=32'h3e515c00;
    in0[123]=32'hf8480a15; in1[123]=32'h7c525722; out[123]=32'hdbb879ca;
    in0[124]=32'h510984e2; in1[124]=32'hba1d8d46; out[124]=32'ha864cfcc;
    in0[125]=32'h824683ac; in1[125]=32'hde34f160; out[125]=32'h23564c80;
    in0[126]=32'h6d95ea79; in1[126]=32'h459b1b4d; out[126]=32'h5a154965;
    in0[127]=32'h4d6c5b12; in1[127]=32'h9f2d863a; out[127]=32'h72620e14;
    in0[128]=32'h2ef0f552; in1[128]=32'h9113c4a5; out[128]=32'h6436e5da;
    in0[129]=32'hc86138ac; in1[129]=32'he1fd5a8b; out[129]=32'h28b23d64;
    in0[130]=32'h705b3dfc; in1[130]=32'hd96c9081; out[130]=32'hb327fbfc;
    in0[131]=32'he3a1b6bb; in1[131]=32'h2e3872a1; out[131]=32'hbefb319b;
    in0[132]=32'h11e5bd1b; in1[132]=32'hea07e059; out[132]=32'h18135e63;
    in0[133]=32'h2104ead6; in1[133]=32'h74824168; out[133]=32'he24bbcf0;
    in0[134]=32'h2a405c7f; in1[134]=32'h5fdbde20; out[134]=32'h59e6b1e0;
    in0[135]=32'hf70431db; in1[135]=32'h1a70d446; out[135]=32'h123efde2;
    in0[136]=32'h620bae7f; in1[136]=32'h845a8375; out[136]=32'h9e47bd0b;
    in0[137]=32'hb3068fc5; in1[137]=32'h6e31c02c; out[137]=32'hdba975dc;
    in0[138]=32'h7a50dbb8; in1[138]=32'he0670e3a; out[138]=32'h895dd7b0;
    in0[139]=32'h8b58ae0c; in1[139]=32'h15e1c4e2; out[139]=32'hde16d698;
    in0[140]=32'hc9105594; in1[140]=32'hf3ab2e40; out[140]=32'hd951fd00;
    in0[141]=32'hb87b5f8e; in1[141]=32'hb0b053ce; out[141]=32'hc4e1ee44;
    in0[142]=32'h36353408; in1[142]=32'hb9d1350a; out[142]=32'h6461b050;
    in0[143]=32'h19f612af; in1[143]=32'hc8d4c354; out[143]=32'h25e56e6c;
    in0[144]=32'h6da5ea7e; in1[144]=32'h2b6316d8; out[144]=32'h9edeae50;
    in0[145]=32'h24273c49; in1[145]=32'hb9a5cb6c; out[145]=32'hf96851cc;
    in0[146]=32'h284209d1; in1[146]=32'h15aa7a66; out[146]=32'h2cc78346;
    in0[147]=32'h2cfced3c; in1[147]=32'h6957d6a3; out[147]=32'h4ebf3534;
    in0[148]=32'ha92c257a; in1[148]=32'hf1f072ac; out[148]=32'h4eb981f8;
    in0[149]=32'h59fd3ff7; in1[149]=32'h72a961c1; out[149]=32'h0538d037;
    in0[150]=32'h885be472; in1[150]=32'hb547ebbb; out[150]=32'heb728546;
    in0[151]=32'h0c766ef7; in1[151]=32'h4073156d; out[151]=32'h9e7c822b;
    in0[152]=32'h0a79a0b1; in1[152]=32'hac32059e; out[152]=32'h25c6a23e;
    in0[153]=32'h58cec29e; in1[153]=32'h5a436932; out[153]=32'ha18ed0dc;
    in0[154]=32'h29ea5695; in1[154]=32'he56aace8; out[154]=32'h913c9308;
    in0[155]=32'he66e0225; in1[155]=32'h532fed3c; out[155]=32'h3d8fc1ac;
    in0[156]=32'h8f8d88cc; in1[156]=32'h919679d7; out[156]=32'h290e4f54;
    in0[157]=32'h38df8e47; in1[157]=32'h1f0c945f; out[157]=32'h9d8ad859;
    in0[158]=32'hbc4b3ab7; in1[158]=32'h5a52e8dd; out[158]=32'hdec587fb;
    in0[159]=32'h085b46c2; in1[159]=32'hdd8f4894; out[159]=32'h81097828;
    in0[160]=32'hefd70ecc; in1[160]=32'h869adb8e; out[160]=32'hb1aab928;
    in0[161]=32'h75c13e5c; in1[161]=32'h17546ddf; out[161]=32'h95127e24;
    in0[162]=32'hbcef8505; in1[162]=32'h0971bccd; out[162]=32'h15b23101;
    in0[163]=32'h91c64a6e; in1[163]=32'h77e35119; out[163]=32'h1b7412be;
    in0[164]=32'h802486ca; in1[164]=32'hc2080107; out[164]=32'hefd67986;
    in0[165]=32'ha84c5fda; in1[165]=32'hbd7afe58; out[165]=32'h413f3ef0;
    in0[166]=32'hdb171d57; in1[166]=32'hc68f1932; out[166]=32'hb9fa39fe;
    in0[167]=32'h75c16123; in1[167]=32'h40ea150b; out[167]=32'h76450b81;
    in0[168]=32'hc1e1b5cc; in1[168]=32'h592df361; out[168]=32'h96f2864c;
    in0[169]=32'hfb00829b; in1[169]=32'h8572e7b4; out[169]=32'ha23bb1fc;
    in0[170]=32'hef3ae1c5; in1[170]=32'h9c06943c; out[170]=32'h72f0ce2c;
    in0[171]=32'h52feee10; in1[171]=32'h09683863; out[171]=32'h23299030;
    in0[172]=32'h5d3d1fd9; in1[172]=32'hff2b58b6; out[172]=32'hccda3c46;
    in0[173]=32'h9223c2ac; in1[173]=32'hd92da212; out[173]=32'hebf08818;
    in0[174]=32'h5a95f71f; in1[174]=32'hdf61f1d2; out[174]=32'h2067e66e;
    in0[175]=32'hd7a387b5; in1[175]=32'he268fd80; out[175]=32'h5a69bb80;
    in0[176]=32'h5e3e30a0; in1[176]=32'hf32a25c1; out[176]=32'he429c8a0;
    in0[177]=32'h193d9671; in1[177]=32'ha8502aad; out[177]=32'h549d345d;
    in0[178]=32'h5d7ec9f5; in1[178]=32'hd3cffcc3; out[178]=32'h427c019f;
    in0[179]=32'h335ad266; in1[179]=32'h37f1b415; out[179]=32'h0e68fa5e;
    in0[180]=32'h6ef9f02e; in1[180]=32'h4bfee527; out[180]=32'h4390bd02;
    in0[181]=32'h7dd02a51; in1[181]=32'hdfc72649; out[181]=32'h3a9b1719;
    in0[182]=32'hc5e0d16b; in1[182]=32'hd50e4f5e; out[182]=32'h8406ea4a;
    in0[183]=32'h6c7722dc; in1[183]=32'hcfb3c156; out[183]=32'h852191e8;
    in0[184]=32'h5a9e2e9e; in1[184]=32'hd5fb12f4; out[184]=32'ha8f58a98;
    in0[185]=32'h47bb68fb; in1[185]=32'h3ee2cc52; out[185]=32'hc945a466;
    in0[186]=32'h712ba121; in1[186]=32'h3661d998; out[186]=32'h30fda498;
    in0[187]=32'he74a85f7; in1[187]=32'h42064cdb; out[187]=32'hce4fee4d;
    in0[188]=32'h0d358178; in1[188]=32'he398216f; out[188]=32'he7239b08;
    in0[189]=32'h4f019ae7; in1[189]=32'h1301b1cf; out[189]=32'hbe4cf7c9;
    in0[190]=32'h9475aae5; in1[190]=32'h2137e41e; out[190]=32'h6e30fad6;
    in0[191]=32'h3a97727d; in1[191]=32'h9432ab85; out[191]=32'h3a91f9f1;
    in0[192]=32'h5b2245b2; in1[192]=32'h619774ac; out[192]=32'h50997b98;
    in0[193]=32'hed2c2809; in1[193]=32'hd488d86a; out[193]=32'h2ed82bba;
    in0[194]=32'hfbc2ee41; in1[194]=32'hd764c9c5; out[194]=32'h72766105;
    in0[195]=32'h7e1418fb; in1[195]=32'h84d5236d; out[195]=32'ha2cff3df;
    in0[196]=32'ha0cff57e; in1[196]=32'h7c1b5264; out[196]=32'h5a284138;
    in0[197]=32'h8b40e8d4; in1[197]=32'h2c89813d; out[197]=32'hed3e4e84;
    in0[198]=32'ha45f7fbe; in1[198]=32'h1d6583b0; out[198]=32'hcbfc0ca0;
    in0[199]=32'hdafd79b9; in1[199]=32'h9d0f20d7; out[199]=32'h30ef5a5f;
    in0[200]=32'hc5c0be81; in1[200]=32'hcf1215ea; out[200]=32'h45e0b6ea;
    in0[201]=32'h9346d97a; in1[201]=32'hcb8cf452; out[201]=32'h60b1f114;
    in0[202]=32'h166e124d; in1[202]=32'h49fb3fb4; out[202]=32'hc264d124;
    in0[203]=32'h3553c7d9; in1[203]=32'h9ce0c010; out[203]=32'h44ff3d90;
    in0[204]=32'h9bb30307; in1[204]=32'h08aa175e; out[204]=32'h7ba6bd92;
    in0[205]=32'h5deb4426; in1[205]=32'h39b68ba7; out[205]=32'heb7e16ca;
    in0[206]=32'h4744250b; in1[206]=32'h9e9219ab; out[206]=32'h2c68d159;
    in0[207]=32'ha9d355c2; in1[207]=32'h0ddcb0ed; out[207]=32'h1053c49a;
    in0[208]=32'h001a1c66; in1[208]=32'h9de73758; out[208]=32'hd31dad10;
    in0[209]=32'hc8a2d971; in1[209]=32'h46444aef; out[209]=32'h0ae7aa7f;
    in0[210]=32'h13d7bea0; in1[210]=32'h4d28230a; out[210]=32'h2e7d5240;
    in0[211]=32'hd5415afc; in1[211]=32'h82dcf376; out[211]=32'h7e0d2428;
    in0[212]=32'hd8bc8ce0; in1[212]=32'h0b3f3b10; out[212]=32'h4b606e00;
    in0[213]=32'h05f84252; in1[213]=32'h40bc9890; out[213]=32'hf73dfe20;
    in0[214]=32'hfc644a3a; in1[214]=32'hd195f70e; out[214]=32'h1edc052c;
    in0[215]=32'he894a00d; in1[215]=32'h799595bd; out[215]=32'h8372ba99;
    in0[216]=32'h71b0cf67; in1[216]=32'h6f9f6364; out[216]=32'h433ed93c;
    in0[217]=32'h37e55cb4; in1[217]=32'hab0612f8; out[217]=32'haeee7660;
    in0[218]=32'hd3fce285; in1[218]=32'he652436a; out[218]=32'h02989a12;
    in0[219]=32'hb0a1907a; in1[219]=32'h9b7c35b3; out[219]=32'hccf9474e;
    in0[220]=32'hb501460b; in1[220]=32'h276b709e; out[220]=32'h39070aca;
    in0[221]=32'hf258edba; in1[221]=32'he7e5eb82; out[221]=32'h30c47674;
    in0[222]=32'h04836a14; in1[222]=32'h470cc4d9; out[222]=32'hf58c3af4;
    in0[223]=32'h5a3380b3; in1[223]=32'hbcb021b3; out[223]=32'ha4aa1029;
    in0[224]=32'ha99556be; in1[224]=32'he1f6840c; out[224]=32'h4c4e08e8;
    in0[225]=32'he2ab629d; in1[225]=32'ha56dddd6; out[225]=32'h9d3ef83e;
    in0[226]=32'h742114f4; in1[226]=32'h87e84d8c; out[226]=32'h1e84d970;
    in0[227]=32'h062133cb; in1[227]=32'h605c3d31; out[227]=32'hd2a648db;
    in0[228]=32'h253163d7; in1[228]=32'h265cf808; out[228]=32'hcd8766b8;
    in0[229]=32'hc714ae5c; in1[229]=32'h1de35fd3; out[229]=32'hca53d9d4;
    in0[230]=32'h6d6deaba; in1[230]=32'h4574eae8; out[230]=32'h2272bc90;
    in0[231]=32'ha4e12a2f; in1[231]=32'h969453c8; out[231]=32'hbdc231b8;
    in0[232]=32'h9ecef5ed; in1[232]=32'h9e40bd89; out[232]=32'h899194d5;
    in0[233]=32'h0c88088c; in1[233]=32'h26cb1b1a; out[233]=32'h2dbba238;
    in0[234]=32'h0301a7f4; in1[234]=32'he4831e32; out[234]=32'h09dd65a8;
    in0[235]=32'hb4d1df26; in1[235]=32'h5e78ab10; out[235]=32'h0afc5460;
    in0[236]=32'h07aa454b; in1[236]=32'hc0045727; out[236]=32'h5da90b6d;
    in0[237]=32'h87cf6cdc; in1[237]=32'ha1fcbf84; out[237]=32'h4dbc4570;
    in0[238]=32'hb88e2c54; in1[238]=32'h01906ab6; out[238]=32'h56ae4bb8;
    in0[239]=32'hc9c74a91; in1[239]=32'hed0abd5a; out[239]=32'h38c743fa;
    in0[240]=32'h205b6f69; in1[240]=32'h6db1c399; out[240]=32'hb91b90c1;
    in0[241]=32'h9fdb295c; in1[241]=32'h8a17a800; out[241]=32'h22686000;
    in0[242]=32'h49f8456b; in1[242]=32'hf747f782; out[242]=32'h98ba7d56;
    in0[243]=32'ha77cbdb4; in1[243]=32'hefbc6e2c; out[243]=32'hbf23f2f0;
    in0[244]=32'h3f6b9639; in1[244]=32'hac7d6c79; out[244]=32'h030f0cf1;
    in0[245]=32'h0e36d935; in1[245]=32'hc3a7585f; out[245]=32'h3197d2ab;
    in0[246]=32'h4dcfbc10; in1[246]=32'h6c46ce0e; out[246]=32'h971128e0;
    in0[247]=32'hf964d8ec; in1[247]=32'hb28129af; out[247]=32'h099a1554;
    in0[248]=32'hab1cce1c; in1[248]=32'h88a2ee89; out[248]=32'ha7c054fc;
    in0[249]=32'h266b218d; in1[249]=32'h5a394ff2; out[249]=32'h6b053a4a;
    in0[250]=32'h32270ce5; in1[250]=32'h0a0cef9f; out[250]=32'h2806cd3b;
    in0[251]=32'h26664bc3; in1[251]=32'h5001d320; out[251]=32'h58fe3160;
    in0[252]=32'h23a3f25d; in1[252]=32'hbd775ef6; out[252]=32'hc4c40b5e;
    in0[253]=32'hfe0d1219; in1[253]=32'hef7313c3; out[253]=32'hf487a40b;
    in0[254]=32'hc6bae0ce; in1[254]=32'h4a37eff6; out[254]=32'h47b657f4;
    in0[255]=32'hf14eb26f; in1[255]=32'h54fa7895; out[255]=32'h02d7e29b;
    in0[256]=32'ha7779e11; in1[256]=32'hd7d1c505; out[256]=32'ha4da2b55;
    in0[257]=32'h487286a7; in1[257]=32'h783de1f0; out[257]=32'hf1820390;
    in0[258]=32'h6d0a23ba; in1[258]=32'h7faa616a; out[258]=32'hfd404504;
    in0[259]=32'h8508150c; in1[259]=32'h24a4c40a; out[259]=32'h8e1e0278;
    in0[260]=32'h434541b1; in1[260]=32'h6a265a0a; out[260]=32'h0412caea;
    in0[261]=32'hc7bb828e; in1[261]=32'hdccae8cf; out[261]=32'h7afb40d2;
    in0[262]=32'h383379f5; in1[262]=32'h04975ccc; out[262]=32'h0c5c3b3c;
    in0[263]=32'h4f7a11db; in1[263]=32'hcab990ff; out[263]=32'h89e5f925;
    in0[264]=32'h683ffeb4; in1[264]=32'hb1e2531b; out[264]=32'h0d3c38fc;
    in0[265]=32'h830492cb; in1[265]=32'h2409d01c; out[265]=32'hc0e7fe34;
    in0[266]=32'h2ed4e2c0; in1[266]=32'h0910246b; out[266]=32'h6eddc640;
    in0[267]=32'h05cce361; in1[267]=32'hf7c2072b; out[267]=32'h7a23d84b;
    in0[268]=32'h6b0d8e18; in1[268]=32'h76ebeec4; out[268]=32'h10831a60;
    in0[269]=32'h309edc08; in1[269]=32'hc4e2319e; out[269]=32'hc93954f0;
    in0[270]=32'h62885fbc; in1[270]=32'he67c3b35; out[270]=32'h1b5c25ec;
    in0[271]=32'h9c0d22e9; in1[271]=32'h9f23050e; out[271]=32'h474175be;
    in0[272]=32'h1091462e; in1[272]=32'hb676cb3d; out[272]=32'h327832f6;
    in0[273]=32'hc28b4b48; in1[273]=32'h764876ee; out[273]=32'h6e732cf0;
    in0[274]=32'h91c732e4; in1[274]=32'hf26df08b; out[274]=32'h19f261cc;
    in0[275]=32'h686f510b; in1[275]=32'h202c24b9; out[275]=32'h6dbb1cf3;
    in0[276]=32'h307c7801; in1[276]=32'h534cc6a4; out[276]=32'h47d9a6a4;
    in0[277]=32'hf050d7d6; in1[277]=32'h1e936a7b; out[277]=32'hf4184fd2;
    in0[278]=32'h860d3200; in1[278]=32'h51debf7b; out[278]=32'h9ca50600;
    in0[279]=32'h7683c0f8; in1[279]=32'h2c10b734; out[279]=32'hf1347a60;
    in0[280]=32'h8791b65a; in1[280]=32'h656cfa9a; out[280]=32'h49b39624;
    in0[281]=32'h59dd85c8; in1[281]=32'h51b9a59a; out[281]=32'hcc046250;
    in0[282]=32'h8c20197f; in1[282]=32'h51dceda3; out[282]=32'h082ecedd;
    in0[283]=32'hbaf7c487; in1[283]=32'h2dde9bc0; out[283]=32'h65e32240;
    in0[284]=32'h32887e2d; in1[284]=32'hb1c0d168; out[284]=32'hb535ff48;
    in0[285]=32'h68fe2a8f; in1[285]=32'h689f0f2b; out[285]=32'h0e008705;
    in0[286]=32'h868ccca9; in1[286]=32'h2944e26a; out[286]=32'h70ddeffa;
    in0[287]=32'hc745aba5; in1[287]=32'h12e5d12b; out[287]=32'h7e6e89b7;
    in0[288]=32'h4669f0bd; in1[288]=32'hf07de8bf; out[288]=32'h477ee503;
    in0[289]=32'h44ef4adf; in1[289]=32'h4735c1c8; out[289]=32'h9b8f9d38;
    in0[290]=32'h7d4faa6e; in1[290]=32'he51ccc78; out[290]=32'h432f8b90;
    in0[291]=32'h65186931; in1[291]=32'h9901ee55; out[291]=32'hf5177b45;
    in0[292]=32'hb52815f6; in1[292]=32'h3a4c714e; out[292]=32'h24f046f4;
    in0[293]=32'hed8f3e7d; in1[293]=32'he69dc5e3; out[293]=32'h81c399d7;
    in0[294]=32'h2e78dfb1; in1[294]=32'h82c02c5e; out[294]=32'h7d948efe;
    in0[295]=32'h03396cd0; in1[295]=32'haf9c1966; out[295]=32'h6341aae0;
    in0[296]=32'h1d7ec22f; in1[296]=32'h18e5279f; out[296]=32'hbd5ac431;
    in0[297]=32'h9e3299bd; in1[297]=32'h9922b25f; out[297]=32'h43c67723;
    in0[298]=32'hec01bdfa; in1[298]=32'he76557d9; out[298]=32'h2eabfeea;
    in0[299]=32'h313c30b1; in1[299]=32'h52cd2e9a; out[299]=32'h1eb2187a;
    in0[300]=32'h4929e525; in1[300]=32'h87b996a9; out[300]=32'hf3a8f36d;
    in0[301]=32'h21ba358e; in1[301]=32'h5dc1ca81; out[301]=32'he325088e;
    in0[302]=32'hcd39e881; in1[302]=32'h0bc71b25; out[302]=32'h0c2b35a5;
    in0[303]=32'h7bdb4c17; in1[303]=32'hc179439e; out[303]=32'h2421fb32;
    in0[304]=32'hbe1f82ea; in1[304]=32'h20c67732; out[304]=32'h48fe57b4;
    in0[305]=32'hd23a4e6f; in1[305]=32'h2b647012; out[305]=32'h92c613ce;
    in0[306]=32'hbdd7052b; in1[306]=32'h55483457; out[306]=32'hec377d9d;
    in0[307]=32'hceef2e5a; in1[307]=32'h36571fd8; out[307]=32'h4d0201f0;
    in0[308]=32'ha542c9a4; in1[308]=32'h0fe359e3; out[308]=32'h2abed06c;
    in0[309]=32'h22ea522a; in1[309]=32'h7ca89e7e; out[309]=32'h119a5cac;
    in0[310]=32'h09969daf; in1[310]=32'hd4954bf3; out[310]=32'hed04f21d;
    in0[311]=32'h3e2e3058; in1[311]=32'h10644993; out[311]=32'h42aeda88;
    in0[312]=32'h04c28347; in1[312]=32'h47b7fa8c; out[312]=32'h175420d4;
    in0[313]=32'h844a8205; in1[313]=32'hafde939e; out[313]=32'h99fb1e16;
    in0[314]=32'h3e9d095d; in1[314]=32'h51befdc6; out[314]=32'hffbc26ee;
    in0[315]=32'h9edbab39; in1[315]=32'hd8719469; out[315]=32'hd33f2e61;
    in0[316]=32'he307c937; in1[316]=32'hdb5ee340; out[316]=32'h989012c0;
    in0[317]=32'hfe15712a; in1[317]=32'h3de33ef7; out[317]=32'hb2565b86;
    in0[318]=32'h1a1cb012; in1[318]=32'h90eca548; out[318]=32'h46251f10;
    in0[319]=32'h1f17cff4; in1[319]=32'h6dbd01e4; out[319]=32'h34292950;
    in0[320]=32'h105bc55a; in1[320]=32'hffd76e1e; out[320]=32'hbe23cc8c;
    in0[321]=32'hfb093a3e; in1[321]=32'he2662482; out[321]=32'hb7944b7c;
    in0[322]=32'h059e15a3; in1[322]=32'h29931c55; out[322]=32'haf74031f;
    in0[323]=32'h3ae8e1c4; in1[323]=32'h85202c97; out[323]=32'hd2aada9c;
    in0[324]=32'hbc19e2a4; in1[324]=32'h57c1cfe5; out[324]=32'hcb0e58b4;
    in0[325]=32'ha981aa5a; in1[325]=32'h10aa07d5; out[325]=32'h544f32e2;
    in0[326]=32'hdb7f68b3; in1[326]=32'hc20a33aa; out[326]=32'he1752fde;
    in0[327]=32'h23a84380; in1[327]=32'h3a25422c; out[327]=32'h43d29a00;
    in0[328]=32'h5e94cd95; in1[328]=32'h3c88d1b7; out[328]=32'h3b5d9a83;
    in0[329]=32'h40593305; in1[329]=32'hed9922f7; out[329]=32'h0dd3e3d3;
    in0[330]=32'heacfa854; in1[330]=32'h74c78ae0; out[330]=32'h4fbc9180;
    in0[331]=32'he09aafbc; in1[331]=32'hbd1335d5; out[331]=32'hbe0a236c;
    in0[332]=32'hb583bc7f; in1[332]=32'h4b1b9eef; out[332]=32'hdab85c91;
    in0[333]=32'h72f2be80; in1[333]=32'h9bc8c686; out[333]=32'h3e66b700;
    in0[334]=32'h02a33ce1; in1[334]=32'hea5f2fde; out[334]=32'h833b1a1e;
    in0[335]=32'h73586a52; in1[335]=32'h9aa9a950; out[335]=32'hedf35ba0;
    in0[336]=32'ha71510b7; in1[336]=32'h3d67fcbf; out[336]=32'hb9cc9c89;
    in0[337]=32'h78846532; in1[337]=32'h3d37b4a6; out[337]=32'he4bec66c;
    in0[338]=32'h87317543; in1[338]=32'he87b2fdb; out[338]=32'hcb079d51;
    in0[339]=32'h7faf79cf; in1[339]=32'h52e1678c; out[339]=32'hcae7e634;
    in0[340]=32'h918d4bad; in1[340]=32'hcf193505; out[340]=32'h5f524b61;
    in0[341]=32'hbec49725; in1[341]=32'h38014301; out[341]=32'he1784625;
    in0[342]=32'hcba2d5c6; in1[342]=32'h677b98a2; out[342]=32'hec1ad74c;
    in0[343]=32'he0d8f342; in1[343]=32'he3ec2b50; out[343]=32'h7b801aa0;
    in0[344]=32'h09a26145; in1[344]=32'h1a40571f; out[344]=32'hacf83a5b;
    in0[345]=32'h398ad762; in1[345]=32'h4d3e963c; out[345]=32'h7a79e6f8;
    in0[346]=32'h5a7b1fb8; in1[346]=32'h54da3cf4; out[346]=32'h7b795b60;
    in0[347]=32'hf59f933f; in1[347]=32'hef3df99e; out[347]=32'hb5b827e2;
    in0[348]=32'h47f452fa; in1[348]=32'h72270452; out[348]=32'hd5a47c14;
    in0[349]=32'h382e7b64; in1[349]=32'h8ca6f02f; out[349]=32'h970e675c;
    in0[350]=32'h5977e140; in1[350]=32'h45216187; out[350]=32'he3d108c0;
    in0[351]=32'hce4b4aab; in1[351]=32'hf0100490; out[351]=32'h3234ac30;
    in0[352]=32'h4ab70502; in1[352]=32'h1edbb5db; out[352]=32'hd5d1b2b6;
    in0[353]=32'hc1b9756e; in1[353]=32'h04d51d64; out[353]=32'h1b4554f8;
    in0[354]=32'h0f5bd55b; in1[354]=32'hd1a139eb; out[354]=32'h05091d89;
    in0[355]=32'h5292538b; in1[355]=32'h787f45e7; out[355]=32'h8c82d96d;
    in0[356]=32'h073509d8; in1[356]=32'hcc982bbf; out[356]=32'h4179a028;
    in0[357]=32'ha38a7dd3; in1[357]=32'h7c9977d0; out[357]=32'ha81e5070;
    in0[358]=32'he3ce3ed3; in1[358]=32'h90970998; out[358]=32'h411fb848;
    in0[359]=32'hf3eac30a; in1[359]=32'hacc60367; out[359]=32'h75799706;
    in0[360]=32'hdb03760a; in1[360]=32'h02e54338; out[360]=32'h7b987030;
    in0[361]=32'h97278147; in1[361]=32'he8c4f906; out[361]=32'h4a0716aa;
    in0[362]=32'h10655e95; in1[362]=32'h1fe5e0d2; out[362]=32'hcc32f63a;
    in0[363]=32'hf8e70168; in1[363]=32'h5f6eae1f; out[363]=32'h599ddb98;
    in0[364]=32'hf3441422; in1[364]=32'h6f510056; out[364]=32'hd5a0c36c;
    in0[365]=32'h844c484f; in1[365]=32'hf563c8c0; out[365]=32'h6340f340;
    in0[366]=32'he067ec5b; in1[366]=32'h3cdff143; out[366]=32'hc7f986d1;
    in0[367]=32'h69e7963d; in1[367]=32'h7fb283a7; out[367]=32'h515e38cb;
    in0[368]=32'h8503508c; in1[368]=32'h07bccccc; out[368]=32'h9da3bf90;
    in0[369]=32'hbfef7179; in1[369]=32'h13fd890d; out[369]=32'h02778425;
    in0[370]=32'hc26b607f; in1[370]=32'h5cf54b56; out[370]=32'hc2e29faa;
    in0[371]=32'hfd20103d; in1[371]=32'h02e206a5; out[371]=32'hb5e5e551;
    in0[372]=32'h8c17bc54; in1[372]=32'hfb1a5315; out[372]=32'hac89aee4;
    in0[373]=32'hd87e0a47; in1[373]=32'hd061f51c; out[373]=32'he28612c4;
    in0[374]=32'h0de756f3; in1[374]=32'hc8405ee0; out[374]=32'hb1194ea0;
    in0[375]=32'h9d308733; in1[375]=32'h42171331; out[375]=32'hfbe7a9c3;
    in0[376]=32'h2236b91b; in1[376]=32'hcb664cee; out[376]=32'h37961b1a;
    in0[377]=32'hc4643707; in1[377]=32'he183b560; out[377]=32'hd01195a0;
    in0[378]=32'h50eb5fee; in1[378]=32'hb51c65dd; out[378]=32'h7c12b676;
    in0[379]=32'h4424567b; in1[379]=32'h81fc7dd5; out[379]=32'h8c8a0357;
    in0[380]=32'h4772bdcb; in1[380]=32'h9e13308b; out[380]=32'haef41d39;
    in0[381]=32'hc651ba43; in1[381]=32'h5224d51d; out[381]=32'h1ea7d897;
    in0[382]=32'h784e9df5; in1[382]=32'hbca44184; out[382]=32'h1b98a754;
    in0[383]=32'haa3f78c6; in1[383]=32'h170c1fdf; out[383]=32'h70322e7a;
    in0[384]=32'hdfdb7a1a; in1[384]=32'hdf6fe8a9; out[384]=32'h45d12b2a;
    in0[385]=32'h689e6563; in1[385]=32'hf1615f30; out[385]=32'h02d5bf90;
    in0[386]=32'hd98a8701; in1[386]=32'hc150d721; out[386]=32'h538d3e21;
    in0[387]=32'he8ac8645; in1[387]=32'he459d68b; out[387]=32'hafe79577;
    in0[388]=32'he5275a4c; in1[388]=32'h274b64f8; out[388]=32'h65a929a0;
    in0[389]=32'hc887f403; in1[389]=32'hbcb6ed2b; out[389]=32'h39dec381;
    in0[390]=32'h262c77d7; in1[390]=32'h9b83b13d; out[390]=32'h5779353b;
    in0[391]=32'hbe39e2a6; in1[391]=32'h6d4d84fe; out[391]=32'h703a78b4;
    in0[392]=32'hfd4b62bf; in1[392]=32'h63da7958; out[392]=32'ha73c38a8;
    in0[393]=32'h31eb0ed8; in1[393]=32'hdd14ee95; out[393]=32'h367c73b8;
    in0[394]=32'h314032d7; in1[394]=32'h89d32311; out[394]=32'h026bc547;
    in0[395]=32'h293052f3; in1[395]=32'haddf4d11; out[395]=32'hbdd59923;
    in0[396]=32'h4c833be5; in1[396]=32'h09ddd75c; out[396]=32'h7827d94c;
    in0[397]=32'h235a5d6c; in1[397]=32'h39aca3af; out[397]=32'h84d1a0d4;
    in0[398]=32'h911e32a6; in1[398]=32'h8ea73717; out[398]=32'ha4e236ea;
    in0[399]=32'he05082e8; in1[399]=32'he5253ed5; out[399]=32'h96391b08;
    in0[400]=32'h804eff2c; in1[400]=32'h41e9ccfe; out[400]=32'hacc43da8;
    in0[401]=32'h9ea72601; in1[401]=32'h09dba185; out[401]=32'h17985f85;
    in0[402]=32'ha23e06cb; in1[402]=32'hc1ca0660; out[402]=32'hb2994e20;
    in0[403]=32'had826f8d; in1[403]=32'he4f1f77b; out[403]=32'hcf09a3bf;
    in0[404]=32'h64d61f05; in1[404]=32'h863a0036; out[404]=32'hea4c8b0e;
    in0[405]=32'h4c4fbfdc; in1[405]=32'h871225c2; out[405]=32'hdca230b8;
    in0[406]=32'h66cd4776; in1[406]=32'hd1e1a1b7; out[406]=32'hbb654b5a;
    in0[407]=32'h2375dcf3; in1[407]=32'hb3ae9815; out[407]=32'hfa0567ef;
    in0[408]=32'h2fff94b5; in1[408]=32'h4ff79261; out[408]=32'h48499295;
    in0[409]=32'h82da5afe; in1[409]=32'h61151514; out[409]=32'hd75bf1d8;
    in0[410]=32'h177a273d; in1[410]=32'h10d532c3; out[410]=32'h3376cd77;
    in0[411]=32'h09995287; in1[411]=32'h44e45613; out[411]=32'h94567a05;
    in0[412]=32'hcb34d9a0; in1[412]=32'h3c3d6423; out[412]=32'hc85c40e0;
    in0[413]=32'h1268632d; in1[413]=32'hf12c0a70; out[413]=32'h8a4725b0;
    in0[414]=32'h76401fd9; in1[414]=32'hd1f42c0b; out[414]=32'h9e0eaa53;
    in0[415]=32'hc05114ce; in1[415]=32'ha170c28f; out[415]=32'h872ebb12;
    in0[416]=32'h0494598b; in1[416]=32'hf554b1bc; out[416]=32'h5776dd14;
    in0[417]=32'hb6d04f2d; in1[417]=32'h1c3e6562; out[417]=32'h43e1103a;
    in0[418]=32'h4bb2c190; in1[418]=32'h7766ca7b; out[418]=32'h7afea030;
    in0[419]=32'hbb7eb320; in1[419]=32'hda5b814f; out[419]=32'ha0bc66e0;
    in0[420]=32'h8f023613; in1[420]=32'h5a55bad7; out[420]=32'h587437f5;
    in0[421]=32'h284c2a9e; in1[421]=32'h6fbb8289; out[421]=32'he1d10a8e;
    in0[422]=32'h860ba2cf; in1[422]=32'ha6ca3ff2; out[422]=32'h4566d8ae;
    in0[423]=32'hcdc95e87; in1[423]=32'h61c93b9f; out[423]=32'h97d9d2d9;
    in0[424]=32'h540a20e4; in1[424]=32'hd91cd541; out[424]=32'ha0e00de4;
    in0[425]=32'ha65feeac; in1[425]=32'h46780927; out[425]=32'ha0a16834;
    in0[426]=32'h7155396b; in1[426]=32'hbdb9af06; out[426]=32'h67927d82;
    in0[427]=32'h86e5b808; in1[427]=32'h16ff4c33; out[427]=32'h125e0998;
    in0[428]=32'hb08aa190; in1[428]=32'h567f53b1; out[428]=32'h88ab6490;
    in0[429]=32'h56cfa254; in1[429]=32'h3822c24d; out[429]=32'h649f7b44;
    in0[430]=32'hda1b2555; in1[430]=32'ha6e633e3; out[430]=32'h76e0095f;
    in0[431]=32'h68ab91e8; in1[431]=32'h29232139; out[431]=32'h86ba64a8;
    in0[432]=32'hf68f4ddb; in1[432]=32'hcb28e872; out[432]=32'h7d972386;
    in0[433]=32'h80cf194b; in1[433]=32'h7179939e; out[433]=32'h7acaad4a;
    in0[434]=32'h5422ba61; in1[434]=32'hc93d6242; out[434]=32'h8e6a2f02;
    in0[435]=32'hf21be95d; in1[435]=32'h72317b0e; out[435]=32'hbb737216;
    in0[436]=32'h4842eef8; in1[436]=32'h4c05c0c6; out[436]=32'h61d6d3d0;
    in0[437]=32'hc97c8d0f; in1[437]=32'h4e4a2df7; out[437]=32'ha44dbc79;
    in0[438]=32'h302dcc6e; in1[438]=32'hed4e7e2d; out[438]=32'h222f1356;
    in0[439]=32'h206fb5fa; in1[439]=32'h4dcae4df; out[439]=32'h88a62cc6;
    in0[440]=32'h87e9cd9c; in1[440]=32'h4f148f6c; out[440]=32'h24ace1d0;
    in0[441]=32'h4adfca26; in1[441]=32'h15d6152d; out[441]=32'h9eafa6ae;
    in0[442]=32'hdf201a3d; in1[442]=32'hbc1d2eb3; out[442]=32'h8d124ea7;
    in0[443]=32'h4ee10118; in1[443]=32'h32f33004; out[443]=32'h25808460;
    in0[444]=32'hb6b40dd1; in1[444]=32'h0bff6268; out[444]=32'he49e9ee8;
    in0[445]=32'h14f9899a; in1[445]=32'h7b8edb59; out[445]=32'h14e3948a;
    in0[446]=32'heb3347b1; in1[446]=32'h6a582040; out[446]=32'h24a00c40;
    in0[447]=32'habab26f8; in1[447]=32'h07b60af7; out[447]=32'hcdf84948;
    in0[448]=32'h352ba96f; in1[448]=32'h446c5805; out[448]=32'h02ec772b;
    in0[449]=32'h704cea88; in1[449]=32'h2cf7157c; out[449]=32'h5db6c1e0;
    in0[450]=32'h499b6d22; in1[450]=32'h0dcc5865; out[450]=32'h28edbe6a;
    in0[451]=32'h36a88abf; in1[451]=32'h4eea4439; out[451]=32'hf4f7a087;
    in0[452]=32'h1395da31; in1[452]=32'hc248d001; out[452]=32'h54a5aa31;
    in0[453]=32'h0ecaa2e7; in1[453]=32'hf8c80ad1; out[453]=32'h0a440497;
    in0[454]=32'h71d790f0; in1[454]=32'h8aafdf0c; out[454]=32'h916bdb40;
    in0[455]=32'hea22c667; in1[455]=32'h65efd9c6; out[455]=32'h6e3bc2aa;
    in0[456]=32'h85c46717; in1[456]=32'h1c950314; out[456]=32'h44f052cc;
    in0[457]=32'h26b1ecc5; in1[457]=32'h6cb2f76d; out[457]=32'he22de2e1;
    in0[458]=32'hba2b3b2c; in1[458]=32'hdcd50e4f; out[458]=32'hdc2faa94;
    in0[459]=32'hc5fddfc2; in1[459]=32'h44fec335; out[459]=32'he97c192a;
    in0[460]=32'h5ab76cfb; in1[460]=32'ha0db97e9; out[460]=32'hdcf33d73;
    in0[461]=32'hb6752a70; in1[461]=32'ha1739668; out[461]=32'h46c6dd80;
    in0[462]=32'h349d7305; in1[462]=32'h37bfaf4a; out[462]=32'hbadeaa72;
    in0[463]=32'hc333e1bd; in1[463]=32'h45eb971c; out[463]=32'h1d522bac;
    in0[464]=32'h3ac73949; in1[464]=32'ha3343292; out[464]=32'h8ca2eda2;
    in0[465]=32'h777ee05c; in1[465]=32'h9098a488; out[465]=32'hb9c220e0;
    in0[466]=32'h63bdcff6; in1[466]=32'hf2c4623f; out[466]=32'hf9aa598a;
    in0[467]=32'h8796d48d; in1[467]=32'hf97c012a; out[467]=32'heedf6c22;
    in0[468]=32'h7bb98415; in1[468]=32'h724aba9e; out[468]=32'hae88c6f6;
    in0[469]=32'h891dc838; in1[469]=32'h4621c8b5; out[469]=32'h55b24f98;
    in0[470]=32'h5b7f7e4e; in1[470]=32'h3cf85d6f; out[470]=32'ha0ba19d2;
    in0[471]=32'h98db9ea5; in1[471]=32'h53f0dca5; out[471]=32'h7b930c59;
    in0[472]=32'h2dafcd38; in1[472]=32'h621dee9f; out[472]=32'h805285c8;
    in0[473]=32'h02fda827; in1[473]=32'hf93d4fdc; out[473]=32'hd92b8a84;
    in0[474]=32'hccd04b7a; in1[474]=32'h8bbe0522; out[474]=32'h87af6834;
    in0[475]=32'h61c20952; in1[475]=32'h6d9bb2bb; out[475]=32'he1ddd2e6;
    in0[476]=32'h371926a4; in1[476]=32'h18f0a985; out[476]=32'hd4535734;
    in0[477]=32'hda36a2f8; in1[477]=32'h7a927ea6; out[477]=32'h8513bcd0;
    in0[478]=32'h5c1013f0; in1[478]=32'h853f4ed8; out[478]=32'h2bb3f280;
    in0[479]=32'had1b0674; in1[479]=32'h1e3f3f39; out[479]=32'h6026fbd4;
    in0[480]=32'hb58a7c06; in1[480]=32'h799b3188; out[480]=32'he0f10930;
    in0[481]=32'h56c235d2; in1[481]=32'h0cea1d88; out[481]=32'h21396190;
    in0[482]=32'h25bbb347; in1[482]=32'hb2155ac4; out[482]=32'hf38f385c;
    in0[483]=32'h83d0ae04; in1[483]=32'h1f51d507; out[483]=32'hc6c2161c;
    in0[484]=32'ha90fa26e; in1[484]=32'hf27b24fd; out[484]=32'h4e24feb6;
    in0[485]=32'h85a919b2; in1[485]=32'h7f5db65d; out[485]=32'h6a5ce1aa;
    in0[486]=32'h6b920915; in1[486]=32'h3601d3cb; out[486]=32'h215e82a7;
    in0[487]=32'hc05ec16d; in1[487]=32'h4d0c8d02; out[487]=32'h8b628bda;
    in0[488]=32'h00242b86; in1[488]=32'h28d8cd5d; out[488]=32'had0e1dae;
    in0[489]=32'heb173b4f; in1[489]=32'h06dbdd7f; out[489]=32'h454e9f31;
    in0[490]=32'h9655f377; in1[490]=32'h7a8376e6; out[490]=32'hfb5696ea;
    in0[491]=32'h5b4cae40; in1[491]=32'h19682e80; out[491]=32'h77a6a000;
    in0[492]=32'hd1108034; in1[492]=32'h6a811e3e; out[492]=32'hb3392498;
    in0[493]=32'h17be06f3; in1[493]=32'h059f4211; out[493]=32'ha1561c23;
    in0[494]=32'hd161b06a; in1[494]=32'h0e55840d; out[494]=32'h601e9d62;
    in0[495]=32'hebb047e5; in1[495]=32'hc351738e; out[495]=32'h1a88c006;
    in0[496]=32'h919c1779; in1[496]=32'h468a4bcd; out[496]=32'h12193ee5;
    in0[497]=32'hb33b88a3; in1[497]=32'h1ce82a35; out[497]=32'h877607bf;
    in0[498]=32'h94c75b34; in1[498]=32'hacaaa1af; out[498]=32'h952b0c8c;
    in0[499]=32'hbff5cfed; in1[499]=32'hb7706b7e; out[499]=32'h9b9465a6;
    in0[500]=32'h89ff8ef9; in1[500]=32'h05d853ec; out[500]=32'h920a888c;
    in0[501]=32'h1fc79367; in1[501]=32'h87a66236; out[501]=32'h005085ba;
    in0[502]=32'h9927705e; in1[502]=32'h38d4162a; out[502]=32'h21f8836c;
    in0[503]=32'h07e72040; in1[503]=32'h9a5f9952; out[503]=32'h220e9480;
    in0[504]=32'h7cb50803; in1[504]=32'h50ffc714; out[504]=32'h625bf53c;
    in0[505]=32'h8c8b46f1; in1[505]=32'hbc9b8979; out[505]=32'he6b680e9;
    in0[506]=32'h6ecd8416; in1[506]=32'ha750bce8; out[506]=32'hf81fdbf0;
    in0[507]=32'h26c011c5; in1[507]=32'hfe40b9d4; out[507]=32'hcb261424;
    in0[508]=32'h61f851bd; in1[508]=32'hcc74ce70; out[508]=32'h540dd8b0;
    in0[509]=32'h5969dc0c; in1[509]=32'h7d1feeb3; out[509]=32'h710c0464;
    in0[510]=32'h9afe52a4; in1[510]=32'h801528f2; out[510]=32'h08c7bf08;
    in0[511]=32'h596e2d01; in1[511]=32'heb0559b5; out[511]=32'h54902ab5;
    in0[512]=32'hfa03b872; in1[512]=32'h5ee2c65c; out[512]=32'h6aa274f8;
    in0[513]=32'h65eae2fc; in1[513]=32'hf5a727a0; out[513]=32'hb9c64180;
    in0[514]=32'haa962b3c; in1[514]=32'h81435276; out[514]=32'h47c525a8;
    in0[515]=32'hb6286f44; in1[515]=32'hd4739e93; out[515]=32'hd96fdc0c;
    in0[516]=32'h58f8eae9; in1[516]=32'h925f6c51; out[516]=32'h38539fb9;
    in0[517]=32'h30cc3af1; in1[517]=32'h74ded52a; out[517]=32'h3f8a308a;
    in0[518]=32'hf6dfd1b0; in1[518]=32'hdfffd3bf; out[518]=32'hd9218250;
    in0[519]=32'hb2731da8; in1[519]=32'h1f3750a0; out[519]=32'h384f0900;
    in0[520]=32'h2a15c3a5; in1[520]=32'h5b6e2c4b; out[520]=32'hc9e6ad57;
    in0[521]=32'h25eba5cb; in1[521]=32'hfed480f9; out[521]=32'h6b35c273;
    in0[522]=32'hfcf372a9; in1[522]=32'hc3d99169; out[522]=32'h900cc051;
    in0[523]=32'h3355b468; in1[523]=32'h14ffc7fb; out[523]=32'hc7dcb9f8;
    in0[524]=32'hd657194e; in1[524]=32'hfcd3eb6e; out[524]=32'hb0f17984;
    in0[525]=32'h7b33e115; in1[525]=32'h16ba7f29; out[525]=32'hcf3a775d;
    in0[526]=32'hfed76553; in1[526]=32'h4aad8b6f; out[526]=32'hea7ffffd;
    in0[527]=32'h8ea179fd; in1[527]=32'h02f53ab6; out[527]=32'hb5910bde;
    in0[528]=32'hb562e909; in1[528]=32'h3ed2309a; out[528]=32'h0093df6a;
    in0[529]=32'hea1fc4a5; in1[529]=32'h455fb3c6; out[529]=32'hbd4c769e;
    in0[530]=32'h6bd38a89; in1[530]=32'h5f9dd850; out[530]=32'hfc03e2d0;
    in0[531]=32'h3eb364ab; in1[531]=32'hed83bd79; out[531]=32'he69dd3d3;
    in0[532]=32'h423ed877; in1[532]=32'h57b6f1f0; out[532]=32'h9a4cf690;
    in0[533]=32'h713913b1; in1[533]=32'h4be69ec1; out[533]=32'h22351671;
    in0[534]=32'hd461bb54; in1[534]=32'ha829ae18; out[534]=32'h76f0a7e0;
    in0[535]=32'h7b219ec1; in1[535]=32'ha8472222; out[535]=32'h8113b7a2;
    in0[536]=32'h8b0fd506; in1[536]=32'hdedfdbaf; out[536]=32'h5f48c11a;
    in0[537]=32'hbc65b0c9; in1[537]=32'h35197ac0; out[537]=32'ha32560c0;
    in0[538]=32'he00858c4; in1[538]=32'hdcc57312; out[538]=32'h3f4a49c8;
    in0[539]=32'h1ffc98a0; in1[539]=32'hd366c955; out[539]=32'ha2744d20;
    in0[540]=32'ha900400b; in1[540]=32'hbd96d03d; out[540]=32'h1e8a329f;
    in0[541]=32'h20150d4a; in1[541]=32'h1193e1e1; out[541]=32'h3eacb80a;
    in0[542]=32'h9aee50d7; in1[542]=32'h4822b24c; out[542]=32'he7837dd4;
    in0[543]=32'hab02ba00; in1[543]=32'hee969349; out[543]=32'h50950a00;
    in0[544]=32'h02ecab3e; in1[544]=32'h2635c3b6; out[544]=32'h0287f814;
    in0[545]=32'hb46883dc; in1[545]=32'h534f4f75; out[545]=32'hb959278c;
    in0[546]=32'h497cceb1; in1[546]=32'h26369698; out[546]=32'ha28c6f18;
    in0[547]=32'h7419250a; in1[547]=32'h8d9e1d0c; out[547]=32'ha88bde78;
    in0[548]=32'h53e951ad; in1[548]=32'hbfe3e969; out[548]=32'h456ff4f5;
    in0[549]=32'hd3e7e1d5; in1[549]=32'h69b2f158; out[549]=32'h86692638;
    in0[550]=32'ha9adb447; in1[550]=32'h54003bc8; out[550]=32'he4413478;
    in0[551]=32'h3f520473; in1[551]=32'h3d254083; out[551]=32'hf3b406d9;
    in0[552]=32'h2303edc4; in1[552]=32'haf905811; out[552]=32'h673e2a04;
    in0[553]=32'h2acb1125; in1[553]=32'he0a557e4; out[553]=32'h8c87d7f4;
    in0[554]=32'hd51195e6; in1[554]=32'h3da9aa0b; out[554]=32'h98222ce2;
    in0[555]=32'hfabcb732; in1[555]=32'h74028e64; out[555]=32'hb5b94b88;
    in0[556]=32'hf332a118; in1[556]=32'h4d47bac1; out[556]=32'h07dee318;
    in0[557]=32'h7f4fa284; in1[557]=32'h1d098de9; out[557]=32'h66a19e24;
    in0[558]=32'h1d03d1b0; in1[558]=32'hbb5d4118; out[558]=32'h6d895880;
    in0[559]=32'hcdb562c0; in1[559]=32'hbaca3103; out[559]=32'h8c86e840;
    in0[560]=32'h25ec4393; in1[560]=32'hae307454; out[560]=32'h15b4c83c;
    in0[561]=32'hfd2bb67d; in1[561]=32'h3cea30cc; out[561]=32'h0b4edb9c;
    in0[562]=32'h874150af; in1[562]=32'h6ae97300; out[562]=32'h3c859d00;
    in0[563]=32'h7d7a33d5; in1[563]=32'h492a8a69; out[563]=32'h9502145d;
    in0[564]=32'hd02c2ba7; in1[564]=32'h2fa112d4; out[564]=32'h9cace44c;
    in0[565]=32'ha403a2d5; in1[565]=32'h34733e55; out[565]=32'hc053a6b9;
    in0[566]=32'h8d39b22e; in1[566]=32'h6b7d02c2; out[566]=32'hb39362dc;
    in0[567]=32'hd17ed76f; in1[567]=32'h40efbdd9; out[567]=32'h1a329017;
    in0[568]=32'h592b57c9; in1[568]=32'h10d1d169; out[568]=32'h308b1a71;
    in0[569]=32'hef4a481a; in1[569]=32'h080cdf17; out[569]=32'h65b32056;
    in0[570]=32'h01bb0ea7; in1[570]=32'hdcc150c9; out[570]=32'h6059b11f;
    in0[571]=32'h2a2d02f8; in1[571]=32'hf6737d51; out[571]=32'hf8190878;
    in0[572]=32'h7456a02b; in1[572]=32'hdc65f8fb; out[572]=32'h210fb229;
    in0[573]=32'h029b7ea6; in1[573]=32'h0f857fb2; out[573]=32'h7a30696c;
    in0[574]=32'hb4bf93c8; in1[574]=32'h7118978f; out[574]=32'h19ee84b8;
    in0[575]=32'h3097015d; in1[575]=32'h6e17d021; out[575]=32'h09edbcfd;
    in0[576]=32'had591abc; in1[576]=32'hc9a69bde; out[576]=32'h385d0308;
    in0[577]=32'h2d0d6180; in1[577]=32'h71e29d49; out[577]=32'ha09c4d80;
    in0[578]=32'hc2f96071; in1[578]=32'h7baec102; out[578]=32'h5f75f1e2;
    in0[579]=32'h799e088a; in1[579]=32'h3bb3f07a; out[579]=32'he3cf71c4;
    in0[580]=32'hf732dfbf; in1[580]=32'h376699fb; out[580]=32'hf5b48745;
    in0[581]=32'h3dd97323; in1[581]=32'he67130a7; out[581]=32'h62e3abd5;
    in0[582]=32'h89225c2f; in1[582]=32'hf30295eb; out[582]=32'h378ffa25;
    in0[583]=32'h17028136; in1[583]=32'hb3ccd87b; out[583]=32'he441a4f2;
    in0[584]=32'hb82753b2; in1[584]=32'hdeb3c49f; out[584]=32'h5df7438e;
    in0[585]=32'h4d9096b8; in1[585]=32'h47de1f97; out[585]=32'hfe192e88;
    in0[586]=32'hc724b7d6; in1[586]=32'h7ff733f3; out[586]=32'he1f42222;
    in0[587]=32'h0231ac72; in1[587]=32'h719d6f45; out[587]=32'h3512e8ba;
    in0[588]=32'ha7492361; in1[588]=32'hff0eccee; out[588]=32'h5c7e302e;
    in0[589]=32'h5bdbead0; in1[589]=32'h2bc6e750; out[589]=32'hb27b1100;
    in0[590]=32'h97493a77; in1[590]=32'h5612b597; out[590]=32'h18e59f31;
    in0[591]=32'hd8c36f47; in1[591]=32'ha3ec09ce; out[591]=32'h16a10a22;
    in0[592]=32'h224acbbb; in1[592]=32'h13c381bb; out[592]=32'hcdbd0c99;
    in0[593]=32'h912feb62; in1[593]=32'h76af5ba0; out[593]=32'hda9cf340;
    in0[594]=32'h85e9bd5d; in1[594]=32'h7210866a; out[594]=32'h0bb71682;
    in0[595]=32'hfabdcbbf; in1[595]=32'h2a5ffa74; out[595]=32'he8d9d88c;
    in0[596]=32'h82c768ab; in1[596]=32'h8ab12274; out[596]=32'h4a7d237c;
    in0[597]=32'h3dcf547d; in1[597]=32'h3dafe7e0; out[597]=32'hb519b860;
    in0[598]=32'ha0250a6f; in1[598]=32'hed3bbedf; out[598]=32'h289778b1;
    in0[599]=32'hea55bca3; in1[599]=32'h568f7f3e; out[599]=32'h6a658c7a;
    in0[600]=32'h87fb9dc1; in1[600]=32'h30123066; out[600]=32'ha3670ae6;
    in0[601]=32'hefe1d3b0; in1[601]=32'h53b6d309; out[601]=32'h1f8a8130;
    in0[602]=32'h56587563; in1[602]=32'h0ac2ca74; out[602]=32'hbfbb4edc;
    in0[603]=32'h8b235b6f; in1[603]=32'hac12258c; out[603]=32'h355b0bb4;
    in0[604]=32'h05886c3e; in1[604]=32'hfb375146; out[604]=32'hb8df36f4;
    in0[605]=32'h876f7539; in1[605]=32'h3b5798c0; out[605]=32'hba90c2c0;
    in0[606]=32'h3ae3c831; in1[606]=32'h11d05d42; out[606]=32'hd74369a2;
    in0[607]=32'hca9571c8; in1[607]=32'h9810d340; out[607]=32'haea44a00;
    in0[608]=32'h4974dfa0; in1[608]=32'h242f8fe2; out[608]=32'hb077cb40;
    in0[609]=32'hd1f68af5; in1[609]=32'h4c3dd4d5; out[609]=32'hb59581d9;
    in0[610]=32'h1234876e; in1[610]=32'h6fd23c2c; out[610]=32'h3b010ee8;
    in0[611]=32'hcbebc633; in1[611]=32'h46815271; out[611]=32'h5a41d283;
    in0[612]=32'h81fd0bb0; in1[612]=32'hbc61436a; out[612]=32'hba85e6e0;
    in0[613]=32'h8ee65edd; in1[613]=32'hf0473ebd; out[613]=32'hca588f29;
    in0[614]=32'h5d6057d0; in1[614]=32'hcc357ca4; out[614]=32'h6a510140;
    in0[615]=32'h1f3d4dab; in1[615]=32'h8b9bd016; out[615]=32'h5de89cb2;
    in0[616]=32'h22941b26; in1[616]=32'hc62018c2; out[616]=32'hdf8822cc;
    in0[617]=32'haac3dfab; in1[617]=32'h9376ac38; out[617]=32'h3ef1d168;
    in0[618]=32'hfd607cd8; in1[618]=32'h4117ff5b; out[618]=32'h3d0f88c8;
    in0[619]=32'h5b4c6de2; in1[619]=32'h56c53038; out[619]=32'hc83c6970;
    in0[620]=32'hd9a5ae02; in1[620]=32'hc1d8b01a; out[620]=32'h56250c34;
    in0[621]=32'h55a72bae; in1[621]=32'ha61fc92b; out[621]=32'hc271f43a;
    in0[622]=32'hc7c38beb; in1[622]=32'hf406edf0; out[622]=32'h935dbb50;
    in0[623]=32'ha8750abb; in1[623]=32'hf7c0694e; out[623]=32'hce4ff7fa;
    in0[624]=32'h9d40d9c4; in1[624]=32'h90d13696; out[624]=32'hdaf2f0d8;
    in0[625]=32'hd448b4e8; in1[625]=32'haef03704; out[625]=32'h3980aba0;
    in0[626]=32'h157d6dc3; in1[626]=32'h0461d998; out[626]=32'hb76676c8;
    in0[627]=32'h27c72fd0; in1[627]=32'hfaea5bbb; out[627]=32'hb09edcf0;
    in0[628]=32'haf1da01c; in1[628]=32'hbc4f693f; out[628]=32'h3799e2e4;
    in0[629]=32'h40ecf94e; in1[629]=32'hfb7579db; out[629]=32'hf73523ba;
    in0[630]=32'hcea7c3c8; in1[630]=32'hff742f61; out[630]=32'h0922e6c8;
    in0[631]=32'h95432aee; in1[631]=32'hc25239a6; out[631]=32'hda58d454;
    in0[632]=32'hf82443be; in1[632]=32'h4442a039; out[632]=32'hd965d54e;
    in0[633]=32'h75d3408a; in1[633]=32'h7120507b; out[633]=32'h9beb224e;
    in0[634]=32'h62083c5c; in1[634]=32'h8ccf7ac0; out[634]=32'h91551d00;
    in0[635]=32'h07c9240a; in1[635]=32'he61749ec; out[635]=32'hc19a1338;
    in0[636]=32'h3fe90226; in1[636]=32'hc6073f6e; out[636]=32'h40b04654;
    in0[637]=32'h825c6e19; in1[637]=32'h8beb9bb3; out[637]=32'hc13d1e7b;
    in0[638]=32'hc201a99d; in1[638]=32'h56942350; out[638]=32'ha7797810;
    in0[639]=32'h8fd51d04; in1[639]=32'h4bf23fb7; out[639]=32'hdd43b9dc;
    in0[640]=32'h96e4844a; in1[640]=32'h01b150c5; out[640]=32'h485aecf2;
    in0[641]=32'h2d57626e; in1[641]=32'h6a6eb968; out[641]=32'h68e57ab0;
    in0[642]=32'h096a8dc8; in1[642]=32'h169c0b08; out[642]=32'h754c0640;
    in0[643]=32'h7e7aeffd; in1[643]=32'h88224367; out[643]=32'h57dfc5cb;
    in0[644]=32'h80cd4236; in1[644]=32'hb37920f4; out[644]=32'h796fdb78;
    in0[645]=32'hdd4d04e4; in1[645]=32'h6d085209; out[645]=32'hae663404;
    in0[646]=32'h72ec3ec0; in1[646]=32'h15eb8379; out[646]=32'h9005e8c0;
    in0[647]=32'h8ea6c2fc; in1[647]=32'h14341276; out[647]=32'hc5c39828;
    in0[648]=32'he2025ba8; in1[648]=32'h1b5995a9; out[648]=32'h284f49e8;
    in0[649]=32'he97bc552; in1[649]=32'hdee3413d; out[649]=32'h234dd68a;
    in0[650]=32'h6906e47a; in1[650]=32'h53018a4e; out[650]=32'h29bd612c;
    in0[651]=32'h973e9bf7; in1[651]=32'hb306187b; out[651]=32'he67e17ad;
    in0[652]=32'h7bc417c5; in1[652]=32'h8e641f54; out[652]=32'hea2ca7a4;
    in0[653]=32'h369aedd7; in1[653]=32'h54b20920; out[653]=32'h313849e0;
    in0[654]=32'h8eeba447; in1[654]=32'h587e2c11; out[654]=32'h40d41cb7;
    in0[655]=32'h4c56b073; in1[655]=32'h83755923; out[655]=32'h10c11ab9;
    in0[656]=32'h00136160; in1[656]=32'h11ae7a11; out[656]=32'hccf13760;
    in0[657]=32'h0402862c; in1[657]=32'headccba9; out[657]=32'h2bdf770c;
    in0[658]=32'h8be5b7d3; in1[658]=32'hafafef8f; out[658]=32'h822cabdd;
    in0[659]=32'h7e6db5b4; in1[659]=32'h29d9c9f5; out[659]=32'hfc3d3944;
    in0[660]=32'h72e81c44; in1[660]=32'h3106e68c; out[660]=32'h0dec8d30;
    in0[661]=32'h65e95c4b; in1[661]=32'hf10d887d; out[661]=32'h06c8e89f;
    in0[662]=32'h427c12db; in1[662]=32'ha728f4f1; out[662]=32'ha7fe7c2b;
    in0[663]=32'h7b24fac1; in1[663]=32'h155c1eb8; out[663]=32'hca52d8b8;
    in0[664]=32'he62ff57c; in1[664]=32'h68b743da; out[664]=32'h6dba7f98;
    in0[665]=32'h1d8e8137; in1[665]=32'h97a9775d; out[665]=32'hb92481fb;
    in0[666]=32'hd6e7073a; in1[666]=32'h46b25771; out[666]=32'h41c2e69a;
    in0[667]=32'hb7f302aa; in1[667]=32'h682eedd5; out[667]=32'h91349972;
    in0[668]=32'hf4d85e7d; in1[668]=32'h3774d316; out[668]=32'h0c1d25be;
    in0[669]=32'h4ac2ccb4; in1[669]=32'h73c38095; out[669]=32'hb2d724c4;
    in0[670]=32'h18412b6f; in1[670]=32'h4c1d46d6; out[670]=32'hf7eda8ca;
    in0[671]=32'hebda608e; in1[671]=32'he31266f4; out[671]=32'h82989b58;
    in0[672]=32'hc00901b3; in1[672]=32'h7081a590; out[672]=32'hfe5c53b0;
    in0[673]=32'h666afa58; in1[673]=32'hbf353f2b; out[673]=32'h03cbb4c8;
    in0[674]=32'h15cb6357; in1[674]=32'h0b98c51c; out[674]=32'h9e58d084;
    in0[675]=32'hf5fd2041; in1[675]=32'hc1b1c680; out[675]=32'h13736680;
    in0[676]=32'hc6c5c409; in1[676]=32'h85461587; out[676]=32'h52d51dbf;
    in0[677]=32'h5040e891; in1[677]=32'h8f07df1b; out[677]=32'h5c65d64b;
    in0[678]=32'hb4a99fca; in1[678]=32'hb390472a; out[678]=32'hcec53d24;
    in0[679]=32'hd34375eb; in1[679]=32'h2bd60958; out[679]=32'h09c7cbc8;
    in0[680]=32'ha24a4f77; in1[680]=32'h752f7ea0; out[680]=32'hfb673c60;
    in0[681]=32'h52ea42cd; in1[681]=32'h0c2e0c6e; out[681]=32'h38a05016;
    in0[682]=32'h87722f16; in1[682]=32'he14b9ba6; out[682]=32'h17feda44;
    in0[683]=32'h14f8199c; in1[683]=32'h5a666afe; out[683]=32'h94ec00c8;
    in0[684]=32'h7d3021cc; in1[684]=32'hcd21a278; out[684]=32'hdb3eefa0;
    in0[685]=32'h71f6fb9d; in1[685]=32'h8c619d0d; out[685]=32'h74570ff9;
    in0[686]=32'h8eebf651; in1[686]=32'h32d358b2; out[686]=32'h53801c52;
    in0[687]=32'h5b00fe01; in1[687]=32'h568dc61f; out[687]=32'h0620881f;
    in0[688]=32'h2e270509; in1[688]=32'hcd077e90; out[688]=32'h82ac4310;
    in0[689]=32'h4774fb11; in1[689]=32'hf8b59e18; out[689]=32'he0f10798;
    in0[690]=32'h0fb27a6c; in1[690]=32'h0ca73923; out[690]=32'hcf1cc8c4;
    in0[691]=32'h3682c016; in1[691]=32'h0d60f88c; out[691]=32'h9fd65c08;
    in0[692]=32'h6f2a83e8; in1[692]=32'h9409c561; out[692]=32'h99c582e8;
    in0[693]=32'h7df19d31; in1[693]=32'h37011b1e; out[693]=32'h621596be;
    in0[694]=32'h5ea794ab; in1[694]=32'h8f4a8691; out[694]=32'hd32ab6db;
    in0[695]=32'h43100787; in1[695]=32'hf96809ae; out[695]=32'h8300dcc2;
    in0[696]=32'h77c01544; in1[696]=32'h4ac54aba; out[696]=32'h8d091b68;
    in0[697]=32'h49e8b394; in1[697]=32'hc0be3494; out[697]=32'h46d9e190;
    in0[698]=32'h844caad1; in1[698]=32'h8945c43f; out[698]=32'h24fb0d6f;
    in0[699]=32'he72c42fe; in1[699]=32'h11b4cdf5; out[699]=32'ha7998316;
    in0[700]=32'h917a0541; in1[700]=32'h6e2012a4; out[700]=32'h5ca9efa4;
    in0[701]=32'hf97bbefd; in1[701]=32'h105a8443; out[701]=32'h0ecf7037;
    in0[702]=32'h019c0f4c; in1[702]=32'h4def12a0; out[702]=32'h1e90e780;
    in0[703]=32'h8ef2a455; in1[703]=32'hd86aa729; out[703]=32'hf141c49d;
    in0[704]=32'h57a6a204; in1[704]=32'h2548d392; out[704]=32'h79b1b248;
    in0[705]=32'hff59eb92; in1[705]=32'haa09a630; out[705]=32'h6bbed760;
    in0[706]=32'hbbb1abdb; in1[706]=32'h35bf1565; out[706]=32'h2f96c467;
    in0[707]=32'h27f61653; in1[707]=32'h6abc4caf; out[707]=32'h22cde6bd;
    in0[708]=32'h8eeacd2f; in1[708]=32'h3e6d227e; out[708]=32'h45d43b22;
    in0[709]=32'h0653ce53; in1[709]=32'h8c906eb8; out[709]=32'h0193f5a8;
    in0[710]=32'h4f9f9aba; in1[710]=32'he837410f; out[710]=32'hfe994ae6;
    in0[711]=32'h7c966fa1; in1[711]=32'hec3b7766; out[711]=32'hb7ef5126;
    in0[712]=32'h862ac559; in1[712]=32'h00c4dd91; out[712]=32'h02bb9c69;
    in0[713]=32'hc26a33f9; in1[713]=32'h12e86478; out[713]=32'h39bda0b8;
    in0[714]=32'h661865df; in1[714]=32'hd9dd4d21; out[714]=32'h784c34bf;
    in0[715]=32'h3a70efaa; in1[715]=32'hca1f1c5e; out[715]=32'hf944986c;
    in0[716]=32'h2a8bc4ba; in1[716]=32'hb7bcf1cd; out[716]=32'h14b7a2f2;
    in0[717]=32'h10a60431; in1[717]=32'h56527b18; out[717]=32'h2145ef98;
    in0[718]=32'h6547c7e7; in1[718]=32'h34b4772e; out[718]=32'h0b3e4c82;
    in0[719]=32'h5fa4ece7; in1[719]=32'h740f6a04; out[719]=32'h5634599c;
    in0[720]=32'h90bc5c64; in1[720]=32'h31ab5289; out[720]=32'ha5317984;
    in0[721]=32'hd2b11a5f; in1[721]=32'h948a6dee; out[721]=32'h6c16f752;
    in0[722]=32'hf66a76d6; in1[722]=32'h29e420f5; out[722]=32'h3f567ace;
    in0[723]=32'h6e9f031f; in1[723]=32'ha75dd3c8; out[723]=32'hd70ffd38;
    in0[724]=32'h379cf2ce; in1[724]=32'h209eb256; out[724]=32'h6ab0cd34;
    in0[725]=32'h3ae6592f; in1[725]=32'hd0c40792; out[725]=32'h5bcb25ce;
    in0[726]=32'h3671fe35; in1[726]=32'h7d4d2807; out[726]=32'ha3c73b73;
    in0[727]=32'h6e8f629d; in1[727]=32'h47721cad; out[727]=32'hda98d019;
    in0[728]=32'h425527f6; in1[728]=32'h251e188c; out[728]=32'h7f24ea88;
    in0[729]=32'haefe5814; in1[729]=32'ha3ff5562; out[729]=32'he8885ba8;
    in0[730]=32'h5b6c52a8; in1[730]=32'he64d321c; out[730]=32'hf485da60;
    in0[731]=32'h0255bf54; in1[731]=32'h9cc835af; out[731]=32'h02da2e6c;
    in0[732]=32'h77708c8b; in1[732]=32'hea9e5ef5; out[732]=32'h6e1b8b07;
    in0[733]=32'hfae1fe5e; in1[733]=32'h22f8e542; out[733]=32'hbdddaa3c;
    in0[734]=32'hb5c7f26b; in1[734]=32'h626325c5; out[734]=32'h7e480357;
    in0[735]=32'hfb39148c; in1[735]=32'hf4cb47e8; out[735]=32'h3b7172e0;
    in0[736]=32'h7b94f843; in1[736]=32'h5553c887; out[736]=32'h4a3c4355;
    in0[737]=32'h7fd29a19; in1[737]=32'hdf534038; out[737]=32'h59b2f578;
    in0[738]=32'h8620dda4; in1[738]=32'h0169e6e5; out[738]=32'h0ecb9bb4;
    in0[739]=32'h285806fc; in1[739]=32'h610c8a7c; out[739]=32'hce373a10;
    in0[740]=32'hbe333c61; in1[740]=32'h42ed5a6c; out[740]=32'h28a492ec;
    in0[741]=32'hded9ac0e; in1[741]=32'hd8d5ef7d; out[741]=32'hff9014d6;
    in0[742]=32'h73c7d1ca; in1[742]=32'hc7b921b4; out[742]=32'hcb848c08;
    in0[743]=32'he1d7ad49; in1[743]=32'hbddb8f99; out[743]=32'h962557a1;
    in0[744]=32'h74a9793a; in1[744]=32'hb9752fb1; out[744]=32'h17f0771a;
    in0[745]=32'h220ff634; in1[745]=32'h37b8d725; out[745]=32'h75744184;
    in0[746]=32'hea79cbec; in1[746]=32'h9df0c356; out[746]=32'h747f4548;
    in0[747]=32'h896762fc; in1[747]=32'hdafa21ff; out[747]=32'h73d61504;
    in0[748]=32'he869d9a0; in1[748]=32'h416a4f22; out[748]=32'h44774740;
    in0[749]=32'hc6f401cf; in1[749]=32'h3c353c5d; out[749]=32'h5aec2c33;
    in0[750]=32'h3be1843a; in1[750]=32'hd0408184; out[750]=32'hb26967e8;
    in0[751]=32'h6d4e0539; in1[751]=32'h50a8b9a0; out[751]=32'heff174a0;
    in0[752]=32'h84b97e74; in1[752]=32'h9abeb48e; out[752]=32'hade5b458;
    in0[753]=32'h6f18a5ec; in1[753]=32'he3291fd3; out[753]=32'h64345584;
    in0[754]=32'h70a80ccf; in1[754]=32'h300874d4; out[754]=32'ha770676c;
    in0[755]=32'h70e7b0ca; in1[755]=32'h691c8a80; out[755]=32'h893d4900;
    in0[756]=32'h03754d8e; in1[756]=32'h99172ce4; out[756]=32'h138f7a78;
    in0[757]=32'hb00070aa; in1[757]=32'hec60dfa8; out[757]=32'hda2e0590;
    in0[758]=32'hb0882116; in1[758]=32'he26d92d5; out[758]=32'h0680134e;
    in0[759]=32'h50b2120e; in1[759]=32'habc4e180; out[759]=32'h079f5500;
    in0[760]=32'h797ed0d9; in1[760]=32'he6666469; out[760]=32'h8b0e6d01;
    in0[761]=32'h01c7c842; in1[761]=32'h926f1856; out[761]=32'hcc81762c;
    in0[762]=32'h8edef358; in1[762]=32'h4b249b5c; out[762]=32'h55d5bba0;
    in0[763]=32'h7673a8a9; in1[763]=32'hc771a080; out[763]=32'h54d6f480;
    in0[764]=32'h4852a3fb; in1[764]=32'h7371ddc2; out[764]=32'h48faf336;
    in0[765]=32'h5846b456; in1[765]=32'h3a31aa36; out[765]=32'h93212624;
    in0[766]=32'hafaa67d4; in1[766]=32'h4b5f9bc8; out[766]=32'h0daa79a0;
    in0[767]=32'h0dbfef5c; in1[767]=32'hb3716244; out[767]=32'h1c38cc70;
    in0[768]=32'h6cda3af6; in1[768]=32'h08a0ce5c; out[768]=32'h439f2468;
    in0[769]=32'h0442d79f; in1[769]=32'h1366fa20; out[769]=32'h854639e0;
    in0[770]=32'hd34713a5; in1[770]=32'h16047b31; out[770]=32'h139f0995;
    in0[771]=32'hceb1e054; in1[771]=32'h70b6c0e3; out[771]=32'hebb0ea7c;
    in0[772]=32'hf4a4cd59; in1[772]=32'hc0e499f2; out[772]=32'h65c84f22;
    in0[773]=32'h9f05d316; in1[773]=32'ha88caebc; out[773]=32'h9dc7f828;
    in0[774]=32'h28e105fe; in1[774]=32'h2c7d6c34; out[774]=32'hd1425f98;
    in0[775]=32'hd784f726; in1[775]=32'h93817d07; out[775]=32'h2d76500a;
    in0[776]=32'h4c214b9e; in1[776]=32'hfa577085; out[776]=32'h1d136916;
    in0[777]=32'hbaef164a; in1[777]=32'h37bebb5d; out[777]=32'hff0f26e2;
    in0[778]=32'ha19a251b; in1[778]=32'hd4fc42a5; out[778]=32'hc87ee067;
    in0[779]=32'hb7f3695f; in1[779]=32'h1d28c52f; out[779]=32'h4f9e7371;
    in0[780]=32'he62456e2; in1[780]=32'hc372bdee; out[780]=32'ha091a01c;
    in0[781]=32'h037c942e; in1[781]=32'h1a85f375; out[781]=32'h807d6306;
    in0[782]=32'hb8527030; in1[782]=32'h9018c157; out[782]=32'h4f185050;
    in0[783]=32'hd2cfd45d; in1[783]=32'hcc3ae070; out[783]=32'h4dd048b0;
    in0[784]=32'ha6901834; in1[784]=32'h13c7e1c8; out[784]=32'h72449ca0;
    in0[785]=32'hfdb87188; in1[785]=32'h48d5a74c; out[785]=32'h5af96c60;
    in0[786]=32'he7e70713; in1[786]=32'h494afa79; out[786]=32'haf98e5fb;
    in0[787]=32'ha05cc6de; in1[787]=32'h4fe9e5e2; out[787]=32'h11da25fc;
    in0[788]=32'hc5a510d0; in1[788]=32'h0e60adee; out[788]=32'hf9d23160;
    in0[789]=32'hd32f17b7; in1[789]=32'h7b52eb64; out[789]=32'h3ec8407c;
    in0[790]=32'h9bbb131c; in1[790]=32'hf73f47b2; out[790]=32'he2440d78;
    in0[791]=32'hfc428160; in1[791]=32'h98cd9b51; out[791]=32'haf400f60;
    in0[792]=32'h3d363a31; in1[792]=32'h7a504f4a; out[792]=32'hf6f1f12a;
    in0[793]=32'he74cb373; in1[793]=32'h09e893f0; out[793]=32'h8e2b44d0;
    in0[794]=32'he411903b; in1[794]=32'hf10f0ba0; out[794]=32'h4aa1ade0;
    in0[795]=32'h19cc3dbd; in1[795]=32'ha2e74acf; out[795]=32'h35898dd3;
    in0[796]=32'hb379882b; in1[796]=32'hacebbba7; out[796]=32'hbe383d0d;
    in0[797]=32'h42035c62; in1[797]=32'h72b030af; out[797]=32'he8fe86fe;
    in0[798]=32'hf0869abf; in1[798]=32'h6a8b433e; out[798]=32'h96ce7742;
    in0[799]=32'h2f808a99; in1[799]=32'h4cc5586a; out[799]=32'hee9afb5a;
    in0[800]=32'h22e37496; in1[800]=32'h9b910e76; out[800]=32'h602df124;
    in0[801]=32'hf14018ee; in1[801]=32'h2398e799; out[801]=32'h5d1da83e;
    in0[802]=32'h87c6b61a; in1[802]=32'h7a4194d3; out[802]=32'h6aa91f6e;
    in0[803]=32'h5e922448; in1[803]=32'hb3216d0f; out[803]=32'hc94ac838;
    in0[804]=32'hcef689b5; in1[804]=32'h0f9adbd6; out[804]=32'h5bc6f44e;
    in0[805]=32'h2b6f3a06; in1[805]=32'h9808c945; out[805]=32'h69b9599e;
    in0[806]=32'haad8fd6f; in1[806]=32'h9b44f677; out[806]=32'h74e27899;
    in0[807]=32'h07cbd38d; in1[807]=32'hb9e8e3bb; out[807]=32'h0b418eff;
    in0[808]=32'hee8d1192; in1[808]=32'h06c8b07e; out[808]=32'h8b9305dc;
    in0[809]=32'h9331da71; in1[809]=32'h0e33cc67; out[809]=32'ha5a3ef77;
    in0[810]=32'h48fc6a82; in1[810]=32'hd7c0a2b4; out[810]=32'h1c612768;
    in0[811]=32'hb040f69f; in1[811]=32'h45a9eb6f; out[811]=32'hb885e3f1;
    in0[812]=32'hdfae8626; in1[812]=32'h40eb4e2c; out[812]=32'h43c0a288;
    in0[813]=32'h590b54c7; in1[813]=32'h2ca8f127; out[813]=32'h12214151;
    in0[814]=32'hbbd5e2c3; in1[814]=32'hf95b758a; out[814]=32'h48405c1e;
    in0[815]=32'hb59400e7; in1[815]=32'h5dd78643; out[815]=32'hab362675;
    in0[816]=32'he61f8fb6; in1[816]=32'ha58877da; out[816]=32'h495dfafc;
    in0[817]=32'hd148953a; in1[817]=32'he73c2677; out[817]=32'h5e7bf9f6;
    in0[818]=32'h22713626; in1[818]=32'hd5516982; out[818]=32'hacb9154c;
    in0[819]=32'h0db9b7b2; in1[819]=32'ha079bc61; out[819]=32'ha9675272;
    in0[820]=32'had6c96cb; in1[820]=32'hace39dd6; out[820]=32'hab418cb2;
    in0[821]=32'h01347f50; in1[821]=32'h48612c2f; out[821]=32'hfbd51fb0;
    in0[822]=32'h6f03624d; in1[822]=32'h12fcd0ff; out[822]=32'h82097ab3;
    in0[823]=32'h42b2dd3b; in1[823]=32'h52b02b2d; out[823]=32'hc329cc5f;
    in0[824]=32'h4e994709; in1[824]=32'hb5f33af9; out[824]=32'hf7b921c1;
    in0[825]=32'h96d0a1fd; in1[825]=32'h46ff7537; out[825]=32'h49de6e5b;
    in0[826]=32'h56ea80f4; in1[826]=32'h465718a2; out[826]=32'h87687a68;
    in0[827]=32'h600688d9; in1[827]=32'h76315ed2; out[827]=32'h6324f002;
    in0[828]=32'hdb339f89; in1[828]=32'h02f0f4e9; out[828]=32'h587ac7b1;
    in0[829]=32'h031fd187; in1[829]=32'he343d99c; out[829]=32'h6b541d44;
    in0[830]=32'h34793c57; in1[830]=32'h79465db3; out[830]=32'h5a7acbd5;
    in0[831]=32'h63bf7a71; in1[831]=32'h16b9e6f6; out[831]=32'h13aa2e96;
    in0[832]=32'h469dfdfd; in1[832]=32'hacdb76b0; out[832]=32'ha3203bf0;
    in0[833]=32'hf59925a7; in1[833]=32'he81e5206; out[833]=32'h91385fea;
    in0[834]=32'had739049; in1[834]=32'hf2cea905; out[834]=32'hca40026d;
    in0[835]=32'h36efae1b; in1[835]=32'h64495a45; out[835]=32'h43826b47;
    in0[836]=32'h238258df; in1[836]=32'h249f7b37; out[836]=32'hd0353ce9;
    in0[837]=32'h1cc4ba42; in1[837]=32'hfe959706; out[837]=32'h9ae34b8c;
    in0[838]=32'h0fe91ce1; in1[838]=32'h52151a39; out[838]=32'ha84b4819;
    in0[839]=32'h30e9bd88; in1[839]=32'h66a69821; out[839]=32'h2cda2e88;
    in0[840]=32'ha7a45ee9; in1[840]=32'h422d160a; out[840]=32'h6d88bb1a;
    in0[841]=32'h1ea2eeee; in1[841]=32'ha9582e4f; out[841]=32'hfb067f72;
    in0[842]=32'h9357886d; in1[842]=32'hdcae50e6; out[842]=32'h215ca1ee;
    in0[843]=32'h993c3957; in1[843]=32'hf5bccb34; out[843]=32'h4097a2ac;
    in0[844]=32'hb5c4c627; in1[844]=32'h5e72e629; out[844]=32'h75e8c63f;
    in0[845]=32'hdd4e0948; in1[845]=32'ha45f4f98; out[845]=32'h0ceabac0;
    in0[846]=32'hd57ff30e; in1[846]=32'h35ce6e8b; out[846]=32'h622cfc9a;
    in0[847]=32'hba754df0; in1[847]=32'h5e18b749; out[847]=32'h74a9c970;
    in0[848]=32'h002c110f; in1[848]=32'h3575c2cb; out[848]=32'h6eb9e4e5;
    in0[849]=32'h42f1ec67; in1[849]=32'h301725e2; out[849]=32'h9dfe95ee;
    in0[850]=32'h8570223f; in1[850]=32'he2ab824d; out[850]=32'h92334af3;
    in0[851]=32'hb08dab1a; in1[851]=32'h6982262b; out[851]=32'h3c65995e;
    in0[852]=32'h1ce61f60; in1[852]=32'hb635f9e9; out[852]=32'he0d6ee60;
    in0[853]=32'h6166676b; in1[853]=32'h80c4ee72; out[853]=32'h41ab87a6;
    in0[854]=32'h60a9faf9; in1[854]=32'hf7b24cd7; out[854]=32'h6565b31f;
    in0[855]=32'hf7fc5bd8; in1[855]=32'hddf61c0c; out[855]=32'hf36fee20;
    in0[856]=32'h8280d70b; in1[856]=32'h62676aa4; out[856]=32'haf01510c;
    in0[857]=32'hbc571b36; in1[857]=32'hee5ce41a; out[857]=32'hb07cdb7c;
    in0[858]=32'h4debbae5; in1[858]=32'ha3344c1d; out[858]=32'h94b427f1;
    in0[859]=32'h6673942b; in1[859]=32'h0cd9b768; out[859]=32'hda51ee78;
    in0[860]=32'h929de9ff; in1[860]=32'h7ba8e6b8; out[860]=32'h56134948;
    in0[861]=32'h48e72bc9; in1[861]=32'h02c25c75; out[861]=32'h25b53edd;
    in0[862]=32'h5c969b37; in1[862]=32'h9a758feb; out[862]=32'h2517347d;
    in0[863]=32'h2b4973bf; in1[863]=32'hecfc9fec; out[863]=32'h8a9e5514;
    in0[864]=32'haa214d5f; in1[864]=32'h22c10bd5; out[864]=32'heea7750b;
    in0[865]=32'hfac69c8b; in1[865]=32'h8a85d7f4; out[865]=32'h14fcf17c;
    in0[866]=32'hbb6d593f; in1[866]=32'hb4333fd7; out[866]=32'h655974e9;
    in0[867]=32'h201bdf98; in1[867]=32'hdc6dcd01; out[867]=32'h45e09798;
    in0[868]=32'hd9dbb1ae; in1[868]=32'he7fa7b47; out[868]=32'h8038e142;
    in0[869]=32'he83f9c2c; in1[869]=32'h861bcd00; out[869]=32'h70b33c00;
    in0[870]=32'hdfe7ab14; in1[870]=32'h72a00316; out[870]=32'hc969efb8;
    in0[871]=32'h18b9f119; in1[871]=32'h2d2995e1; out[871]=32'hf6c173f9;
    in0[872]=32'h290de2a2; in1[872]=32'h1168f552; out[872]=32'h4427a1e4;
    in0[873]=32'h6540deed; in1[873]=32'ha0a6bace; out[873]=32'h49d994b6;
    in0[874]=32'hd9c933dc; in1[874]=32'h9d47677e; out[874]=32'h72e90a48;
    in0[875]=32'hafd53f92; in1[875]=32'h9cb6a46a; out[875]=32'h94d1da74;
    in0[876]=32'h9b95ff41; in1[876]=32'h9624304a; out[876]=32'h145bf8ca;
    in0[877]=32'h0f9690d2; in1[877]=32'h978b2515; out[877]=32'h8a4e3b3a;
    in0[878]=32'h024e4482; in1[878]=32'ha711e8a6; out[878]=32'hc7783c4c;
    in0[879]=32'h5ab0c19e; in1[879]=32'h4194d5c3; out[879]=32'h3313f15a;
    in0[880]=32'hf10559e8; in1[880]=32'h7982f9e4; out[880]=32'h2d06baa0;
    in0[881]=32'hb4bace11; in1[881]=32'h120867fe; out[881]=32'h1cc94bde;
    in0[882]=32'ha1192886; in1[882]=32'hef88349c; out[882]=32'he8bfe9a8;
    in0[883]=32'hd3da0c6b; in1[883]=32'hdb6fa8a9; out[883]=32'hde7d6aa3;
    in0[884]=32'ha542a42c; in1[884]=32'hc744f219; out[884]=32'hf263a04c;
    in0[885]=32'h27b54b1d; in1[885]=32'h8d45f01c; out[885]=32'h8610672c;
    in0[886]=32'h8c6ca4b1; in1[886]=32'h6fb43912; out[886]=32'h9bc2fd72;
    in0[887]=32'h3838a3ae; in1[887]=32'h2ad7068b; out[887]=32'hddb8f37a;
    in0[888]=32'h6361d786; in1[888]=32'hd057b4a4; out[888]=32'h94c249d8;
    in0[889]=32'h52f576e6; in1[889]=32'h70df5d01; out[889]=32'hb18104e6;
    in0[890]=32'h425e7c2a; in1[890]=32'hbfbe4942; out[890]=32'h8aeffcd4;
    in0[891]=32'h32ae06a3; in1[891]=32'h6ffb74d0; out[891]=32'h37384070;
    in0[892]=32'h1f9299de; in1[892]=32'h9d3beba6; out[892]=32'ha8788ff4;
    in0[893]=32'he00034af; in1[893]=32'h60e869f0; out[893]=32'h74652b10;
    in0[894]=32'he46090cc; in1[894]=32'h5eca7b95; out[894]=32'h7abe4abc;
    in0[895]=32'h6df504dc; in1[895]=32'h10549105; out[895]=32'h45b9b44c;
    in0[896]=32'hea69b44c; in1[896]=32'h44cfc6da; out[896]=32'h58ea50b8;
    in0[897]=32'hd998f2cf; in1[897]=32'ha331e107; out[897]=32'ha73592a9;
    in0[898]=32'h8dee83c7; in1[898]=32'h9db08e22; out[898]=32'hca95e26e;
    in0[899]=32'he90b1d77; in1[899]=32'h4f042daf; out[899]=32'h71a30f59;
    in0[900]=32'h2d3808e7; in1[900]=32'h875ee752; out[900]=32'h21cd4afe;
    in0[901]=32'h512b991e; in1[901]=32'hd1601039; out[901]=32'hb586f7ae;
    in0[902]=32'h52555c7b; in1[902]=32'hb7645560; out[902]=32'h44c38520;
    in0[903]=32'h9b87db2b; in1[903]=32'hff276316; out[903]=32'h1ffb76b2;
    in0[904]=32'h4b6a1102; in1[904]=32'h82d5f871; out[904]=32'h34f571e2;
    in0[905]=32'hee9fc019; in1[905]=32'h0f7587f5; out[905]=32'hdf9d06ed;
    in0[906]=32'h03d5e1ce; in1[906]=32'hf4584465; out[906]=32'h4a2cce46;
    in0[907]=32'h4e13a879; in1[907]=32'h1dc77e41; out[907]=32'h2af854b9;
    in0[908]=32'hd6c35404; in1[908]=32'h5b962024; out[908]=32'h44505090;
    in0[909]=32'h449712a2; in1[909]=32'h2185b14f; out[909]=32'h2eaac1fe;
    in0[910]=32'h620027dc; in1[910]=32'hd82f8e03; out[910]=32'h2d807f94;
    in0[911]=32'h5b87389b; in1[911]=32'he02dfe04; out[911]=32'h2b85ac6c;
    in0[912]=32'hff7b67e8; in1[912]=32'h03c02cd4; out[912]=32'h6e0dec20;
    in0[913]=32'h7922eb46; in1[913]=32'h0afab1f0; out[913]=32'h33c3f7a0;
    in0[914]=32'h830ef7de; in1[914]=32'hf587d3eb; out[914]=32'hd11b82ca;
    in0[915]=32'h3d7cad14; in1[915]=32'h0224d4d1; out[915]=32'hf0eddd54;
    in0[916]=32'h400214f0; in1[916]=32'h7ffc383a; out[916]=32'ha14d3e60;
    in0[917]=32'h9cea8cc1; in1[917]=32'h5be30a05; out[917]=32'ha43749c5;
    in0[918]=32'h65c3d702; in1[918]=32'h5b8cf6e4; out[918]=32'h1e1f69c8;
    in0[919]=32'h586e040f; in1[919]=32'he0cc912a; out[919]=32'h2e4d2976;
    in0[920]=32'h0adceb49; in1[920]=32'hae1858fd; out[920]=32'h5a0d9f25;
    in0[921]=32'h44fbed33; in1[921]=32'h41b15987; out[921]=32'he993d0e5;
    in0[922]=32'ha1361dfb; in1[922]=32'h9fc369fb; out[922]=32'hfd8c5819;
    in0[923]=32'hedddf017; in1[923]=32'hf52bc1b9; out[923]=32'h8e40d79f;
    in0[924]=32'h6b2ac1d8; in1[924]=32'hbedaa861; out[924]=32'h0c5932d8;
    in0[925]=32'ha2538568; in1[925]=32'h89011976; out[925]=32'h27eea5f0;
    in0[926]=32'hb38b2c97; in1[926]=32'h22d1d502; out[926]=32'ha876fc2e;
    in0[927]=32'h1e8dcda7; in1[927]=32'hbc0865f9; out[927]=32'hbb47ea6f;
    in0[928]=32'h62a04d42; in1[928]=32'he3e3e90c; out[928]=32'h8d5ab118;
    in0[929]=32'h0a5b33a2; in1[929]=32'h09137d43; out[929]=32'hc51a9d66;
    in0[930]=32'hf761404b; in1[930]=32'h1f37f967; out[930]=32'h04c6d12d;
    in0[931]=32'h33125917; in1[931]=32'hae27a759; out[931]=32'hedfff9ff;
    in0[932]=32'h94591673; in1[932]=32'hbef9009f; out[932]=32'h532ff16d;
    in0[933]=32'ha8bcc9ca; in1[933]=32'h95f13469; out[933]=32'h1795cbda;
    in0[934]=32'h6d5f8168; in1[934]=32'hf7c01f9e; out[934]=32'h779d7630;
    in0[935]=32'h84e791f1; in1[935]=32'hbc85e823; out[935]=32'hd6205bf3;
    in0[936]=32'h81136a65; in1[936]=32'hb39ec118; out[936]=32'h065e1e78;
    in0[937]=32'h6b98237a; in1[937]=32'he9bbf4c2; out[937]=32'h7f392a74;
    in0[938]=32'hfbc88922; in1[938]=32'h585bcdbc; out[938]=32'hec2aeef8;
    in0[939]=32'h51aaea89; in1[939]=32'h29ab689f; out[939]=32'hc2f25317;
    in0[940]=32'h1e52d098; in1[940]=32'h2897a1a5; out[940]=32'h6a3809f8;
    in0[941]=32'h4951ce7a; in1[941]=32'h8892eead; out[941]=32'h2bd1f472;
    in0[942]=32'h3a773ceb; in1[942]=32'h686a0506; out[942]=32'h644a0482;
    in0[943]=32'h28b26b37; in1[943]=32'ha915122b; out[943]=32'h7c04e03d;
    in0[944]=32'hbb62d718; in1[944]=32'hbd9c98ad; out[944]=32'h1c219b38;
    in0[945]=32'h0e1b6b25; in1[945]=32'hd6634915; out[945]=32'h571c5709;
    in0[946]=32'h8a12f39b; in1[946]=32'h8fe8a50d; out[946]=32'h937145df;
    in0[947]=32'hace3497f; in1[947]=32'hc792cbae; out[947]=32'h6131a952;
    in0[948]=32'hf1e33f32; in1[948]=32'h5041bdea; out[948]=32'h8b11adb4;
    in0[949]=32'hfb13090f; in1[949]=32'hec3582d7; out[949]=32'h3bb13999;
    in0[950]=32'h0f0e6582; in1[950]=32'hc8c343c6; out[950]=32'h4bb9888c;
    in0[951]=32'hb934822e; in1[951]=32'ha01052e9; out[951]=32'h455d37de;
    in0[952]=32'hc9ea3217; in1[952]=32'h9bc9c080; out[952]=32'hdbb94b80;
    in0[953]=32'h46dcad91; in1[953]=32'h1ed38538; out[953]=32'h32f54cb8;
    in0[954]=32'h822ceb31; in1[954]=32'hfb95f346; out[954]=32'h2a0cd266;
    in0[955]=32'ha5c9f9a2; in1[955]=32'hce261c59; out[955]=32'h24918152;
    in0[956]=32'he049c89c; in1[956]=32'hfabaec4b; out[956]=32'hd3e595b4;
    in0[957]=32'hc18fc20c; in1[957]=32'h0f637478; out[957]=32'h9df465a0;
    in0[958]=32'h8d9b3ff9; in1[958]=32'h111a5551; out[958]=32'h62a6eac9;
    in0[959]=32'h09c9adb0; in1[959]=32'hf87aba4c; out[959]=32'hb5f17040;
    in0[960]=32'h26c959fa; in1[960]=32'hee68e73b; out[960]=32'h9a28529e;
    in0[961]=32'h468e3a8f; in1[961]=32'h6ae13517; out[961]=32'h7695ddd9;
    in0[962]=32'hfdaa8e92; in1[962]=32'h8b61e5f6; out[962]=32'h9ebf9a4c;
    in0[963]=32'hb5a8d252; in1[963]=32'h291d87e1; out[963]=32'ha5941812;
    in0[964]=32'h5a75b528; in1[964]=32'h1e436362; out[964]=32'h3f95d150;
    in0[965]=32'haf4aca69; in1[965]=32'h9570d177; out[965]=32'h35f3cfcf;
    in0[966]=32'h5477dba9; in1[966]=32'h068a4325; out[966]=32'hf2e9fa6d;
    in0[967]=32'h49380ddb; in1[967]=32'h291a7e5f; out[967]=32'h3ddcee45;
    in0[968]=32'h6311b748; in1[968]=32'hf394b902; out[968]=32'he1367690;
    in0[969]=32'h9dca68b1; in1[969]=32'hc286eee4; out[969]=32'ha43fcba4;
    in0[970]=32'h4cc0cbc9; in1[970]=32'h4178dbb4; out[970]=32'h751c3c54;
    in0[971]=32'h2c44a9e5; in1[971]=32'h81a61118; out[971]=32'h45362278;
    in0[972]=32'hf6eb60ca; in1[972]=32'hb323a9dc; out[972]=32'h0eca8798;
    in0[973]=32'h64fe0070; in1[973]=32'hec0eb6e7; out[973]=32'hfba20510;
    in0[974]=32'h570918e2; in1[974]=32'he740a2f6; out[974]=32'h8afced2c;
    in0[975]=32'hf5c0beaa; in1[975]=32'ha3bd4293; out[975]=32'hd0574f9e;
    in0[976]=32'hca884cb9; in1[976]=32'hb712fab6; out[976]=32'hbbd53586;
    in0[977]=32'h7183f4f5; in1[977]=32'hcb6bd8a3; out[977]=32'h471aafff;
    in0[978]=32'h32c090c8; in1[978]=32'he3805d9b; out[978]=32'h6b305118;
    in0[979]=32'h27a01739; in1[979]=32'ha85b5cc6; out[979]=32'hd76d7216;
    in0[980]=32'hca1ecd06; in1[980]=32'h1f6324cf; out[980]=32'hc70e9fda;
    in0[981]=32'h93e0efb0; in1[981]=32'h43c8dc61; out[981]=32'ha7b611b0;
    in0[982]=32'h54508e7c; in1[982]=32'h0ce4ea44; out[982]=32'hbe1330f0;
    in0[983]=32'h98b644c4; in1[983]=32'h48e914cd; out[983]=32'h3db860f4;
    in0[984]=32'h48afee7f; in1[984]=32'h0431950c; out[984]=32'h705e18f4;
    in0[985]=32'hcd7fb32e; in1[985]=32'hb53707cc; out[985]=32'h448b0aa8;
    in0[986]=32'hed11e356; in1[986]=32'h7399c6de; out[986]=32'hebbda894;
    in0[987]=32'hdbf49b9c; in1[987]=32'h38c12e37; out[987]=32'ha61f7684;
    in0[988]=32'h7962888e; in1[988]=32'hb46b88fe; out[988]=32'hb3a8ece4;
    in0[989]=32'h260a77ed; in1[989]=32'ha4ddc857; out[989]=32'h76d8e98b;
    in0[990]=32'hf4b1b206; in1[990]=32'he64ab8d3; out[990]=32'h40260af2;
    in0[991]=32'h45b35df2; in1[991]=32'h801d317f; out[991]=32'h8d60ed0e;
    in0[992]=32'h67ab1a9e; in1[992]=32'hb324b580; out[992]=32'h07970500;
    in0[993]=32'h49845ba5; in1[993]=32'h73ee210b; out[993]=32'h8ae63517;
    in0[994]=32'he547b72d; in1[994]=32'hd8ed9d9e; out[994]=32'h0a42a6c6;
    in0[995]=32'h2c79afab; in1[995]=32'h30e71b97; out[995]=32'ha49aa6dd;
    in0[996]=32'h598abf4b; in1[996]=32'h87a7ad1c; out[996]=32'he55f9b34;
    in0[997]=32'hda26caf5; in1[997]=32'hb2840d76; out[997]=32'h8683fdee;
    in0[998]=32'h8f6579b8; in1[998]=32'h0c42201d; out[998]=32'hef25c9d8;
    in0[999]=32'hfe455497; in1[999]=32'h344d1e55; out[999]=32'haa59c823;
  end
  // Initial Block
  initial begin
    // Reset signal
    #10 reset = 1'b0;
    // Parse Arguments
    if ( !$value$plusargs( "nmults=%d", nmults ) ) begin
      $display( "No nmults specified!  Example: ./simv +nmults=10" ); $finish;
    end
    if ( !$value$plusargs( "verbose=%d", verbose ) ) begin
      verbose = 0;
    end
    // Set request valid high
    src_val = 1'b1;
    // Always end simulation after a set time to prevent renegade simulations
    // from filling up our drives with a huge VCD file...
    #100000000000
    $display( "###  ERROR: Simulation timed out!!!  ###" );
    $finish;
  end
  // Begin Sim Loop
  reg        busy = 1'b0;
  reg [31:0] cycle_count = 32'd0;
  always @ ( * ) begin
    src_msg_a <= in0[ idx % 1000 ];
    src_msg_b <= in1[ idx % 1000 ];
  end
  always @ ( posedge clk ) begin
    // Line Trace
    //$display( "%d ( %h %h | %h )",
    //              cycle_count,
    //              imul.dpath.a_reg, imul.dpath.b_reg,
    //              imul.dpath.result_reg[31:0] );
    // Computation has started
    if ( muldivreq_go ) begin
      busy <= 1'b1;
    end
    // Result is ready, display output, increment index.
    else if ( muldivresp_go ) begin
      // Weird first one fails, second passes... hmm.
      //$display( "%h, %d", sink_msg, sink_msg );
      //$display( "%h, %d", out[idx], out[idx] );
      //$display( "%h, %d", src_msg_a * src_msg_b, src_msg_a * src_msg_b );
      //`VC_TEST_EQ( "MulVar", sink_msg, out[ idx ])
      //`VC_TEST_EQ( "MulVar", sink_msg, src_msg_a*src_msg_b)
      //$display( "%h * %h = %h", src_msg_a, src_msg_b, sink_msg );
      `VC_TEST_EQ( "MulVar", sink_msg, out[ idx % 1000 ])
      idx = idx + 1;
    end
    // We've done all the multiplies! Print cycle count and terminate.
    if ( idx == nmults ) begin
      $display( "Cycle Count = %d", cycle_count );
      $finish;
    end
    // Reset val signal after operands have been accepted
    //if ( src_val ) begin
    //  src_val <= 1'b0;
    //end
    // If computation has started, start counting cycles. We need to
    // count starting the clock edge when new operands are flopped in to
    // accurately measure the total clock cycles since the simulation
    // terminates before the final clock cycle can be flopped into the register.
    if ( muldivreq_go || busy ) begin
      cycle_count <= cycle_count + 1;
    end
  end
endmodule