module CapSense_CSD_P4_v2_0_3 (
    sclk2);
    output      sclk2;
          wire  Net_534;
          wire  Net_474;
          wire  Net_540;
          wire  Net_329;
          wire  Net_312;
          wire  Net_104;
          wire  Net_328;
    electrical  Net_398;
    electrical  Net_241;
    electrical  Net_246;
          wire  Net_420;
          wire  Net_429;
    electrical [3:0] Net_245;
          wire  Net_248;
    electrical  Net_270;
    cy_psoc4_csd_v1_0 CSD_FFB (
        .source(Net_245[3:0]),
        .csh(Net_246),
        .shield(Net_241),
        .cmod(Net_398),
        .sample_out(Net_328),
        .sense_in(Net_104),
        .clk1(Net_429),
        .clk2(Net_420),
        .irq(Net_248),
        .sample_in(Net_312),
        .sense_out(Net_329),
        .amuxa(Net_270));
    defparam CSD_FFB.sensors_count = 4;
    defparam CSD_FFB.shield_count = 1;
	cy_clock_v1_0
		#(.id("3c8c7eac-aaf5-41b9-9d0a-e31e77bfd8ce/74063576-f256-4f8f-8a82-9abdee876261"),
		  .source_clock_id("413DE2EF-D9F2-4233-A808-DFAF137FD877"),
		  .divisor(255),
		  .period("0"),
		  .is_direct(0),
		  .is_digital(0))
		SampleClk
		 (.clock_out(Net_420));
	wire [0:0] tmpOE__Cmod_net;
	wire [0:0] tmpFB_0__Cmod_net;
	wire [0:0] tmpIO_0__Cmod_net;
	wire [0:0] tmpINTERRUPT_0__Cmod_net;
	electrical [0:0] tmpSIOVREF__Cmod_net;
	cy_psoc3_pins_v1_10
		#(.id("3c8c7eac-aaf5-41b9-9d0a-e31e77bfd8ce/899719c0-e797-4403-a44f-07a66de2cbeb"),
		  .drive_mode(3'b000),
		  .ibuf_enabled(1'b0),
		  .init_dr_st(1'b1),
		  .input_clk_en(0),
		  .input_sync(1'b1),
		  .input_sync_mode(1'b0),
		  .intr_mode(2'b00),
		  .invert_in_clock(0),
		  .invert_in_clock_en(0),
		  .invert_in_reset(0),
		  .invert_out_clock(0),
		  .invert_out_clock_en(0),
		  .invert_out_reset(0),
		  .io_voltage(""),
		  .layout_mode("CONTIGUOUS"),
		  .oe_conn(1'b0),
		  .oe_reset(0),
		  .oe_sync(1'b0),
		  .output_clk_en(0),
		  .output_clock_mode(1'b0),
		  .output_conn(1'b0),
		  .output_mode(1'b0),
		  .output_reset(0),
		  .output_sync(1'b0),
		  .pa_in_clock(-1),
		  .pa_in_clock_en(-1),
		  .pa_in_reset(-1),
		  .pa_out_clock(-1),
		  .pa_out_clock_en(-1),
		  .pa_out_reset(-1),
		  .pin_aliases("Cmod"),
		  .pin_mode("A"),
		  .por_state(4),
		  .sio_group_cnt(0),
		  .sio_hyst(1'b0),
		  .sio_ibuf(""),
		  .sio_info(2'b00),
		  .sio_obuf(""),
		  .sio_refsel(""),
		  .sio_vtrip(""),
		  .slew_rate(1'b0),
		  .spanning(0),
		  .use_annotation(1'b0),
		  .vtrip(2'b10),
		  .width(1))
		Cmod
		 (.oe(tmpOE__Cmod_net),
		  .y({1'b0}),
		  .fb({tmpFB_0__Cmod_net[0:0]}),
		  .analog({Net_398}),
		  .io({tmpIO_0__Cmod_net[0:0]}),
		  .siovref(tmpSIOVREF__Cmod_net),
		  .interrupt({tmpINTERRUPT_0__Cmod_net[0:0]}),
		  .in_clock({1'b0}),
		  .in_clock_en({1'b1}),
		  .in_reset({1'b0}),
		  .out_clock({1'b0}),
		  .out_clock_en({1'b1}),
		  .out_reset({1'b0}));
	assign tmpOE__Cmod_net = (`CYDEV_CHIP_MEMBER_USED == `CYDEV_CHIP_MEMBER_3A && `CYDEV_CHIP_REVISION_USED < `CYDEV_CHIP_REVISION_3A_ES3) ? ~{1'b1} : {1'b1};
	cy_isr_v1_0
		#(.int_type(2'b10))
		ISR
		 (.int_signal(Net_248));
    IDAC_P4_v1_0_1 IDAC2 (
        .Iout(Net_270));
	wire [3:0] tmpOE__Sns_net;
	wire [3:0] tmpFB_3__Sns_net;
	wire [3:0] tmpIO_3__Sns_net;
	wire [0:0] tmpINTERRUPT_0__Sns_net;
	electrical [0:0] tmpSIOVREF__Sns_net;
	cy_psoc3_pins_v1_10
		#(.id("3c8c7eac-aaf5-41b9-9d0a-e31e77bfd8ce/73b612cd-240c-4d8e-8340-ea28aabf4b11"),
		  .drive_mode(12'b000_000_000_000),
		  .ibuf_enabled(4'b0_0_0_0),
		  .init_dr_st(4'b1_1_1_1),
		  .input_clk_en(0),
		  .input_sync(4'b1_1_1_1),
		  .input_sync_mode(4'b0_0_0_0),
		  .intr_mode(8'b00_00_00_00),
		  .invert_in_clock(0),
		  .invert_in_clock_en(0),
		  .invert_in_reset(0),
		  .invert_out_clock(0),
		  .invert_out_clock_en(0),
		  .invert_out_reset(0),
		  .io_voltage(",,,"),
		  .layout_mode("NONCONTIGUOUS"),
		  .oe_conn(4'b0_0_0_0),
		  .oe_reset(0),
		  .oe_sync(4'b0_0_0_0),
		  .output_clk_en(0),
		  .output_clock_mode(4'b0_0_0_0),
		  .output_conn(4'b0_0_0_0),
		  .output_mode(4'b0_0_0_0),
		  .output_reset(0),
		  .output_sync(4'b0_0_0_0),
		  .pa_in_clock(-1),
		  .pa_in_clock_en(-1),
		  .pa_in_reset(-1),
		  .pa_out_clock(-1),
		  .pa_out_clock_en(-1),
		  .pa_out_reset(-1),
		  .pin_aliases("Button0__BTN,Button1__BTN,Button2__BTN,Button3__BTN"),
		  .pin_mode("AAAA"),
		  .por_state(4),
		  .sio_group_cnt(0),
		  .sio_hyst(4'b0_0_0_0),
		  .sio_ibuf(""),
		  .sio_info(8'b00_00_00_00),
		  .sio_obuf(""),
		  .sio_refsel(""),
		  .sio_vtrip(""),
		  .slew_rate(4'b0_0_0_0),
		  .spanning(1),
		  .use_annotation(4'b0_0_0_0),
		  .vtrip(8'b10_10_10_10),
		  .width(4))
		Sns
		 (.oe(tmpOE__Sns_net),
		  .y({4'b0}),
		  .fb({tmpFB_3__Sns_net[3:0]}),
		  .analog({Net_245[3:0]}),
		  .io({tmpIO_3__Sns_net[3:0]}),
		  .siovref(tmpSIOVREF__Sns_net),
		  .interrupt({tmpINTERRUPT_0__Sns_net[0:0]}),
		  .in_clock({1'b0}),
		  .in_clock_en({1'b1}),
		  .in_reset({1'b0}),
		  .out_clock({1'b0}),
		  .out_clock_en({1'b1}),
		  .out_reset({1'b0}));
	assign tmpOE__Sns_net = (`CYDEV_CHIP_MEMBER_USED == `CYDEV_CHIP_MEMBER_3A && `CYDEV_CHIP_REVISION_USED < `CYDEV_CHIP_REVISION_3A_ES3) ? ~{4'b1111} : {4'b1111};
    IDAC_P4_v1_0_2 IDAC1 (
        .Iout(Net_270));
    ZeroTerminal ZeroTerminal_1 (
        .z(Net_312));
    ZeroTerminal ZeroTerminal_2 (
        .z(Net_104));
    assign sclk2 = Net_420 | Net_474;
    ZeroTerminal ZeroTerminal_7 (
        .z(Net_474));
	cy_clock_v1_0
		#(.id("3c8c7eac-aaf5-41b9-9d0a-e31e77bfd8ce/9a635726-510c-483c-9c5c-3e233ee2906a"),
		  .source_clock_id("413DE2EF-D9F2-4233-A808-DFAF137FD877"),
		  .divisor(255),
		  .period("0"),
		  .is_direct(0),
		  .is_digital(0))
		SenseClk
		 (.clock_out(Net_429));
endmodule