module without the
   // following additional dead code
   wire    a;
   assign		a = | in;
`endif
endmodule