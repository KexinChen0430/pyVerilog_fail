module ADC_SAR_SEQ_P4_v1_10_1 (
    soc,
    aclk,
    Vref,
    sdone,
    eoc,
    vinPlus0);
    input       soc;
    input       aclk;
    inout       Vref;
    electrical  Vref;
    output      sdone;
    output      eoc;
    inout       vinPlus0;
    electrical  vinPlus0;
          wire  Net_3093;
          wire  Net_3090;
          wire  Net_2786;
    electrical  Net_2785;
    electrical  Net_2784;
    electrical  Net_2783;
          wire  Net_2782;
    electrical  Net_2781;
    electrical  Net_2780;
    electrical  Net_2779;
    electrical  Net_2575;
    electrical  Net_2574;
    electrical  Net_2573;
    electrical  Net_2572;
    electrical  Net_2571;
    electrical  Net_2570;
    electrical  Net_2569;
    electrical  Net_2568;
    electrical  Net_2567;
    electrical  Net_2566;
    electrical  Net_2565;
    electrical  Net_2564;
    electrical  muxout_plus;
    electrical  Net_2563;
    electrical  Net_2562;
    electrical  Net_2561;
    electrical  Net_2560;
    electrical  Net_2559;
    electrical  Net_2557;
    electrical  Net_2556;
    electrical  Net_2555;
    electrical  Net_2554;
    electrical  muxout_minus;
    electrical  Net_2553;
    electrical  Net_2552;
    electrical  Net_2551;
    electrical  Net_2550;
    electrical  Net_2549;
    electrical  Net_2548;
    electrical  Net_2547;
    electrical [16:0] mux_bus_minus;
    electrical [16:0] mux_bus_plus;
    electrical  Net_2546;
    electrical  Net_2545;
    electrical  Net_2544;
    electrical  Net_2542;
    electrical  Net_2541;
          wire  Net_2221;
    electrical  Net_1849;
    electrical  Net_1848;
    electrical  Net_1846;
          wire  Net_2273;
          wire [11:0] Net_2272;
          wire  Net_2271;
          wire [3:0] Net_2270;
          wire  Net_2269;
          wire  Net_15;
          wire  Net_13;
          wire  Net_14;
          wire  Net_11;
          wire  Net_26;
    electrical  Net_2793;
    electrical  Net_2794;
          wire  Net_1845;
    electrical [0:0] Net_1450;
    electrical [0:0] Net_2375;
    electrical  Net_1851;
    electrical  Net_2580;
    electrical  Net_3046;
    electrical  Net_3016;
    electrical  Net_2020;
    electrical  Net_124;
    electrical  Net_2102;
    electrical  Net_2099;
          wire [1:0] Net_1963;
          wire  Net_17;
    electrical  Net_8;
    electrical  Net_43;
    cy_psoc4_sar_v1_0 cy_psoc4_sar (
        .vplus(Net_2020),
        .vminus(Net_124),
        .vref(Net_8),
        .ext_vref(Net_43),
        .clock(Net_17),
        .sw_negvref(Net_26),
        .cfg_st_sel(Net_1963[1:0]),
        .cfg_average(Net_11),
        .cfg_resolution(Net_14),
        .cfg_differential(Net_13),
        .trigger(soc),
        .data_hilo_sel(Net_15),
        .sample_done(sdone),
        .chan_id_valid(Net_2269),
        .chan_id(Net_2270[3:0]),
        .data_valid(Net_2271),
        .eos_intr(eoc),
        .data(Net_2272[11:0]),
        .irq(Net_2273));
	// clk_src_sel (cy_virtualmux_v1_0)
	assign Net_17 = Net_1845;
	// int_vref_sel (cy_analog_virtualmux_v1_0)
	cy_connect_v1_0 int_vref_sel_connect(Net_8, Net_1846);
	defparam int_vref_sel_connect.sig_width = 1;
	// ext_vref_sel (cy_analog_virtualmux_v1_0)
	cy_connect_v1_0 ext_vref_sel_connect(Net_43, Net_1849);
	defparam ext_vref_sel_connect.sig_width = 1;
    cy_analog_noconnect_v1_0 cy_analog_noconnect_1 (
        .noconnect(Net_1846));
    ZeroTerminal ZeroTerminal_3 (
        .z(Net_14));
    ZeroTerminal ZeroTerminal_4 (
        .z(Net_13));
    ZeroTerminal ZeroTerminal_5 (
        .z(Net_15));
    ZeroTerminal ZeroTerminal_6 (
        .z(Net_1963[0]));
    ZeroTerminal ZeroTerminal_7 (
        .z(Net_1963[1]));
	cy_clock_v1_0
		#(.id("b0574397-86aa-4552-91b4-736ae77c7a57/a12a1691-924f-48e5-a017-176d592c3b32"),
		  .source_clock_id(""),
		  .divisor(0),
		  .period("333334666.672"),
		  .is_direct(0),
		  .is_digital(0))
		intClock
		 (.clock_out(Net_1845));
    ZeroTerminal ZeroTerminal_2 (
        .z(Net_11));
    ZeroTerminal ZeroTerminal_1 (
        .z(Net_26));
	wire [0:0] tmpOE__ExtVref_net;
	wire [0:0] tmpFB_0__ExtVref_net;
	wire [0:0] tmpIO_0__ExtVref_net;
	wire [0:0] tmpINTERRUPT_0__ExtVref_net;
	electrical [0:0] tmpSIOVREF__ExtVref_net;
	cy_psoc3_pins_v1_10
		#(.id("b0574397-86aa-4552-91b4-736ae77c7a57/05a9c8de-3ba2-4909-8250-95fdc61c0bf4"),
		  .drive_mode(3'b000),
		  .ibuf_enabled(1'b0),
		  .init_dr_st(1'b1),
		  .input_clk_en(0),
		  .input_sync(1'b1),
		  .input_sync_mode(1'b0),
		  .intr_mode(2'b00),
		  .invert_in_clock(0),
		  .invert_in_clock_en(0),
		  .invert_in_reset(0),
		  .invert_out_clock(0),
		  .invert_out_clock_en(0),
		  .invert_out_reset(0),
		  .io_voltage(""),
		  .layout_mode("CONTIGUOUS"),
		  .oe_conn(1'b0),
		  .oe_reset(0),
		  .oe_sync(1'b0),
		  .output_clk_en(0),
		  .output_clock_mode(1'b0),
		  .output_conn(1'b0),
		  .output_mode(1'b0),
		  .output_reset(0),
		  .output_sync(1'b0),
		  .pa_in_clock(-1),
		  .pa_in_clock_en(-1),
		  .pa_in_reset(-1),
		  .pa_out_clock(-1),
		  .pa_out_clock_en(-1),
		  .pa_out_reset(-1),
		  .pin_aliases(""),
		  .pin_mode("A"),
		  .por_state(4),
		  .sio_group_cnt(0),
		  .sio_hyst(1'b0),
		  .sio_ibuf(""),
		  .sio_info(2'b00),
		  .sio_obuf(""),
		  .sio_refsel(""),
		  .sio_vtrip(""),
		  .slew_rate(1'b0),
		  .spanning(0),
		  .use_annotation(1'b0),
		  .vtrip(2'b10),
		  .width(1))
		ExtVref
		 (.oe(tmpOE__ExtVref_net),
		  .y({1'b0}),
		  .fb({tmpFB_0__ExtVref_net[0:0]}),
		  .analog({Net_1849}),
		  .io({tmpIO_0__ExtVref_net[0:0]}),
		  .siovref(tmpSIOVREF__ExtVref_net),
		  .interrupt({tmpINTERRUPT_0__ExtVref_net[0:0]}),
		  .in_clock({1'b0}),
		  .in_clock_en({1'b1}),
		  .in_reset({1'b0}),
		  .out_clock({1'b0}),
		  .out_clock_en({1'b1}),
		  .out_reset({1'b0}));
	assign tmpOE__ExtVref_net = (`CYDEV_CHIP_MEMBER_USED == `CYDEV_CHIP_MEMBER_3A && `CYDEV_CHIP_REVISION_USED < `CYDEV_CHIP_REVISION_3A_ES3) ? ~{1'b1} : {1'b1};
	// ext_vneg_sel (cy_analog_virtualmux_v1_0)
	cy_connect_v1_0 ext_vneg_sel_connect(Net_2580, Net_1851);
	defparam ext_vneg_sel_connect.sig_width = 1;
    cy_analog_noconnect_v1_0 cy_analog_noconnect_3 (
        .noconnect(Net_1851));
	// cy_analog_virtualmux_vplus9 (cy_analog_virtualmux_v1_0)
	cy_connect_v1_0 cy_analog_virtualmux_vplus9_connect(mux_bus_plus[9], Net_2541);
	defparam cy_analog_virtualmux_vplus9_connect.sig_width = 1;
	// cy_analog_virtualmux_vplus8 (cy_analog_virtualmux_v1_0)
	cy_connect_v1_0 cy_analog_virtualmux_vplus8_connect(mux_bus_plus[8], Net_2542);
	defparam cy_analog_virtualmux_vplus8_connect.sig_width = 1;
	// cy_analog_virtualmux_vplus1 (cy_analog_virtualmux_v1_0)
	cy_connect_v1_0 cy_analog_virtualmux_vplus1_connect(mux_bus_plus[1], Net_2544);
	defparam cy_analog_virtualmux_vplus1_connect.sig_width = 1;
	// cy_analog_virtualmux_vplus2 (cy_analog_virtualmux_v1_0)
	cy_connect_v1_0 cy_analog_virtualmux_vplus2_connect(mux_bus_plus[2], Net_2545);
	defparam cy_analog_virtualmux_vplus2_connect.sig_width = 1;
	// cy_analog_virtualmux_vplus3 (cy_analog_virtualmux_v1_0)
	cy_connect_v1_0 cy_analog_virtualmux_vplus3_connect(mux_bus_plus[3], Net_2546);
	defparam cy_analog_virtualmux_vplus3_connect.sig_width = 1;
	// cy_analog_virtualmux_vplus4 (cy_analog_virtualmux_v1_0)
	cy_connect_v1_0 cy_analog_virtualmux_vplus4_connect(mux_bus_plus[4], Net_2547);
	defparam cy_analog_virtualmux_vplus4_connect.sig_width = 1;
	// cy_analog_virtualmux_vplus6 (cy_analog_virtualmux_v1_0)
	cy_connect_v1_0 cy_analog_virtualmux_vplus6_connect(mux_bus_plus[6], Net_2548);
	defparam cy_analog_virtualmux_vplus6_connect.sig_width = 1;
	// cy_analog_virtualmux_vplus7 (cy_analog_virtualmux_v1_0)
	cy_connect_v1_0 cy_analog_virtualmux_vplus7_connect(mux_bus_plus[7], Net_2549);
	defparam cy_analog_virtualmux_vplus7_connect.sig_width = 1;
    Bus_Connect_v1_10 Connect_1 (
        .in_bus(mux_bus_plus[16:0]),
        .out_bus(Net_1450[0:0]));
    defparam Connect_1.in_width = 17;
    defparam Connect_1.out_width = 1;
	// cy_analog_virtualmux_vplus5 (cy_analog_virtualmux_v1_0)
	cy_connect_v1_0 cy_analog_virtualmux_vplus5_connect(mux_bus_plus[5], Net_2550);
	defparam cy_analog_virtualmux_vplus5_connect.sig_width = 1;
	// cy_analog_virtualmux_vplus10 (cy_analog_virtualmux_v1_0)
	cy_connect_v1_0 cy_analog_virtualmux_vplus10_connect(mux_bus_plus[10], Net_2551);
	defparam cy_analog_virtualmux_vplus10_connect.sig_width = 1;
	// cy_analog_virtualmux_vplus11 (cy_analog_virtualmux_v1_0)
	cy_connect_v1_0 cy_analog_virtualmux_vplus11_connect(mux_bus_plus[11], Net_2552);
	defparam cy_analog_virtualmux_vplus11_connect.sig_width = 1;
	// cy_analog_virtualmux_vplus12 (cy_analog_virtualmux_v1_0)
	cy_connect_v1_0 cy_analog_virtualmux_vplus12_connect(mux_bus_plus[12], Net_2553);
	defparam cy_analog_virtualmux_vplus12_connect.sig_width = 1;
	// cy_analog_virtualmux_vplus13 (cy_analog_virtualmux_v1_0)
	cy_connect_v1_0 cy_analog_virtualmux_vplus13_connect(mux_bus_plus[13], Net_2554);
	defparam cy_analog_virtualmux_vplus13_connect.sig_width = 1;
	// cy_analog_virtualmux_vplus14 (cy_analog_virtualmux_v1_0)
	cy_connect_v1_0 cy_analog_virtualmux_vplus14_connect(mux_bus_plus[14], Net_2555);
	defparam cy_analog_virtualmux_vplus14_connect.sig_width = 1;
	// cy_analog_virtualmux_vplus15 (cy_analog_virtualmux_v1_0)
	cy_connect_v1_0 cy_analog_virtualmux_vplus15_connect(mux_bus_plus[15], Net_2556);
	defparam cy_analog_virtualmux_vplus15_connect.sig_width = 1;
	// cy_analog_virtualmux_vplus_inj (cy_analog_virtualmux_v1_0)
	cy_connect_v1_0 cy_analog_virtualmux_vplus_inj_connect(Net_3016, Net_2557);
	defparam cy_analog_virtualmux_vplus_inj_connect.sig_width = 1;
    cy_analog_noconnect_v1_0 cy_analog_noconnect_6 (
        .noconnect(Net_2544));
    cy_analog_noconnect_v1_0 cy_analog_noconnect_7 (
        .noconnect(Net_2545));
    cy_analog_noconnect_v1_0 cy_analog_noconnect_8 (
        .noconnect(Net_2546));
    cy_analog_noconnect_v1_0 cy_analog_noconnect_9 (
        .noconnect(Net_2547));
    cy_analog_noconnect_v1_0 cy_analog_noconnect_10 (
        .noconnect(Net_2550));
    cy_analog_noconnect_v1_0 cy_analog_noconnect_11 (
        .noconnect(Net_2548));
    cy_analog_noconnect_v1_0 cy_analog_noconnect_12 (
        .noconnect(Net_2549));
    cy_analog_noconnect_v1_0 cy_analog_noconnect_13 (
        .noconnect(Net_2542));
    cy_analog_noconnect_v1_0 cy_analog_noconnect_14 (
        .noconnect(Net_2541));
    cy_analog_noconnect_v1_0 cy_analog_noconnect_15 (
        .noconnect(Net_2551));
    cy_analog_noconnect_v1_0 cy_analog_noconnect_16 (
        .noconnect(Net_2552));
    cy_analog_noconnect_v1_0 cy_analog_noconnect_17 (
        .noconnect(Net_2553));
    cy_analog_noconnect_v1_0 cy_analog_noconnect_18 (
        .noconnect(Net_2554));
    cy_analog_noconnect_v1_0 cy_analog_noconnect_19 (
        .noconnect(Net_2555));
    cy_analog_noconnect_v1_0 cy_analog_noconnect_20 (
        .noconnect(Net_2556));
    cy_analog_noconnect_v1_0 cy_analog_noconnect_21 (
        .noconnect(Net_2557));
	// cy_analog_virtualmux_37 (cy_analog_virtualmux_v1_0)
	cy_connect_v1_0 cy_analog_virtualmux_37_connect(Net_3016, mux_bus_plus[1]);
	defparam cy_analog_virtualmux_37_connect.sig_width = 1;
	// cy_analog_virtualmux_vminus0 (cy_analog_virtualmux_v1_0)
	cy_connect_v1_0 cy_analog_virtualmux_vminus0_connect(mux_bus_minus[0], Net_2559);
	defparam cy_analog_virtualmux_vminus0_connect.sig_width = 1;
	// cy_analog_virtualmux_vminus1 (cy_analog_virtualmux_v1_0)
	cy_connect_v1_0 cy_analog_virtualmux_vminus1_connect(mux_bus_minus[1], Net_2560);
	defparam cy_analog_virtualmux_vminus1_connect.sig_width = 1;
	// cy_analog_virtualmux_vminus2 (cy_analog_virtualmux_v1_0)
	cy_connect_v1_0 cy_analog_virtualmux_vminus2_connect(mux_bus_minus[2], Net_2561);
	defparam cy_analog_virtualmux_vminus2_connect.sig_width = 1;
	// cy_analog_virtualmux_vminus3 (cy_analog_virtualmux_v1_0)
	cy_connect_v1_0 cy_analog_virtualmux_vminus3_connect(mux_bus_minus[3], Net_2562);
	defparam cy_analog_virtualmux_vminus3_connect.sig_width = 1;
	// cy_analog_virtualmux_vminus4 (cy_analog_virtualmux_v1_0)
	cy_connect_v1_0 cy_analog_virtualmux_vminus4_connect(mux_bus_minus[4], Net_2563);
	defparam cy_analog_virtualmux_vminus4_connect.sig_width = 1;
	// cy_analog_virtualmux_vminus5 (cy_analog_virtualmux_v1_0)
	cy_connect_v1_0 cy_analog_virtualmux_vminus5_connect(mux_bus_minus[5], Net_2564);
	defparam cy_analog_virtualmux_vminus5_connect.sig_width = 1;
	// cy_analog_virtualmux_vminus6 (cy_analog_virtualmux_v1_0)
	cy_connect_v1_0 cy_analog_virtualmux_vminus6_connect(mux_bus_minus[6], Net_2565);
	defparam cy_analog_virtualmux_vminus6_connect.sig_width = 1;
	// cy_analog_virtualmux_vminus7 (cy_analog_virtualmux_v1_0)
	cy_connect_v1_0 cy_analog_virtualmux_vminus7_connect(mux_bus_minus[7], Net_2566);
	defparam cy_analog_virtualmux_vminus7_connect.sig_width = 1;
	// cy_analog_virtualmux_vminus8 (cy_analog_virtualmux_v1_0)
	cy_connect_v1_0 cy_analog_virtualmux_vminus8_connect(mux_bus_minus[8], Net_2567);
	defparam cy_analog_virtualmux_vminus8_connect.sig_width = 1;
	// cy_analog_virtualmux_vminus9 (cy_analog_virtualmux_v1_0)
	cy_connect_v1_0 cy_analog_virtualmux_vminus9_connect(mux_bus_minus[9], Net_2568);
	defparam cy_analog_virtualmux_vminus9_connect.sig_width = 1;
	// cy_analog_virtualmux_vminus10 (cy_analog_virtualmux_v1_0)
	cy_connect_v1_0 cy_analog_virtualmux_vminus10_connect(mux_bus_minus[10], Net_2569);
	defparam cy_analog_virtualmux_vminus10_connect.sig_width = 1;
	// cy_analog_virtualmux_vminus11 (cy_analog_virtualmux_v1_0)
	cy_connect_v1_0 cy_analog_virtualmux_vminus11_connect(mux_bus_minus[11], Net_2570);
	defparam cy_analog_virtualmux_vminus11_connect.sig_width = 1;
	// cy_analog_virtualmux_vminus12 (cy_analog_virtualmux_v1_0)
	cy_connect_v1_0 cy_analog_virtualmux_vminus12_connect(mux_bus_minus[12], Net_2571);
	defparam cy_analog_virtualmux_vminus12_connect.sig_width = 1;
	// cy_analog_virtualmux_vminus13 (cy_analog_virtualmux_v1_0)
	cy_connect_v1_0 cy_analog_virtualmux_vminus13_connect(mux_bus_minus[13], Net_2572);
	defparam cy_analog_virtualmux_vminus13_connect.sig_width = 1;
	// cy_analog_virtualmux_vminus14 (cy_analog_virtualmux_v1_0)
	cy_connect_v1_0 cy_analog_virtualmux_vminus14_connect(mux_bus_minus[14], Net_2573);
	defparam cy_analog_virtualmux_vminus14_connect.sig_width = 1;
	// cy_analog_virtualmux_vminus15 (cy_analog_virtualmux_v1_0)
	cy_connect_v1_0 cy_analog_virtualmux_vminus15_connect(mux_bus_minus[15], Net_2574);
	defparam cy_analog_virtualmux_vminus15_connect.sig_width = 1;
	// cy_analog_virtualmux_vminus_inj (cy_analog_virtualmux_v1_0)
	cy_connect_v1_0 cy_analog_virtualmux_vminus_inj_connect(Net_3046, Net_2575);
	defparam cy_analog_virtualmux_vminus_inj_connect.sig_width = 1;
    cy_analog_noconnect_v1_0 cy_analog_noconnect_37 (
        .noconnect(Net_2575));
	// cy_analog_virtualmux_36 (cy_analog_virtualmux_v1_0)
	cy_connect_v1_0 cy_analog_virtualmux_36_connect(Net_3046, mux_bus_minus[1]);
	defparam cy_analog_virtualmux_36_connect.sig_width = 1;
	// cy_analog_virtualmux_42 (cy_analog_virtualmux_v1_0)
	cy_connect_v1_0 cy_analog_virtualmux_42_connect(Net_2020, muxout_plus);
	defparam cy_analog_virtualmux_42_connect.sig_width = 1;
	// cy_analog_virtualmux_43 (cy_analog_virtualmux_v1_0)
	cy_connect_v1_0 cy_analog_virtualmux_43_connect(Net_124, muxout_minus);
	defparam cy_analog_virtualmux_43_connect.sig_width = 1;
    cy_analog_noconnect_v1_0 cy_analog_noconnect_39 (
        .noconnect(Net_2779));
    cy_analog_noconnect_v1_0 cy_analog_noconnect_40 (
        .noconnect(Net_2783));
    cy_analog_noconnect_v1_0 cy_analog_noconnect_38 (
        .noconnect(Net_2780));
    cy_analog_noconnect_v1_0 cy_analog_noconnect_41 (
        .noconnect(Net_2781));
    cy_analog_noconnect_v1_0 cy_analog_noconnect_43 (
        .noconnect(Net_2784));
    cy_analog_noconnect_v1_0 cy_analog_noconnect_44 (
        .noconnect(Net_2785));
    Bus_Connect_v1_10 Connect_2 (
        .in_bus(mux_bus_minus[16:0]),
        .out_bus(Net_2375[0:0]));
    defparam Connect_2.in_width = 17;
    defparam Connect_2.out_width = 1;
    cy_analog_noconnect_v1_0 cy_analog_noconnect_2 (
        .noconnect(Net_2559));
    cy_analog_noconnect_v1_0 cy_analog_noconnect_4 (
        .noconnect(Net_2560));
    cy_analog_noconnect_v1_0 cy_analog_noconnect_22 (
        .noconnect(Net_2561));
    cy_analog_noconnect_v1_0 cy_analog_noconnect_23 (
        .noconnect(Net_2562));
    cy_analog_noconnect_v1_0 cy_analog_noconnect_24 (
        .noconnect(Net_2563));
    cy_analog_noconnect_v1_0 cy_analog_noconnect_25 (
        .noconnect(Net_2564));
    cy_analog_noconnect_v1_0 cy_analog_noconnect_26 (
        .noconnect(Net_2565));
    cy_analog_noconnect_v1_0 cy_analog_noconnect_27 (
        .noconnect(Net_2566));
    cy_analog_noconnect_v1_0 cy_analog_noconnect_28 (
        .noconnect(Net_2567));
    cy_analog_noconnect_v1_0 cy_analog_noconnect_29 (
        .noconnect(Net_2568));
    cy_analog_noconnect_v1_0 cy_analog_noconnect_30 (
        .noconnect(Net_2569));
    cy_analog_noconnect_v1_0 cy_analog_noconnect_31 (
        .noconnect(Net_2570));
    cy_analog_noconnect_v1_0 cy_analog_noconnect_32 (
        .noconnect(Net_2571));
    cy_analog_noconnect_v1_0 cy_analog_noconnect_33 (
        .noconnect(Net_2572));
    cy_analog_noconnect_v1_0 cy_analog_noconnect_34 (
        .noconnect(Net_2573));
    cy_analog_noconnect_v1_0 cy_analog_noconnect_35 (
        .noconnect(Net_2574));
	cy_isr_v1_0
		#(.int_type(2'b10))
		IRQ
		 (.int_signal(Net_2273));
    assign Net_3093 = Net_1845 | Net_3090;
    ZeroTerminal ZeroTerminal_8 (
        .z(Net_3090));
	// adc_plus_in_sel (cy_analog_virtualmux_v1_0)
	cy_connect_v1_0 adc_plus_in_sel_connect(muxout_plus, mux_bus_plus[0]);
	defparam adc_plus_in_sel_connect.sig_width = 1;
	// adc_minus_in_sel (cy_analog_virtualmux_v1_0)
	cy_connect_v1_0 adc_minus_in_sel_connect(muxout_minus, mux_bus_minus[0]);
	defparam adc_minus_in_sel_connect.sig_width = 1;
    cy_connect_v1_0 vinPlus0__cy_connect_v1_0(vinPlus0, mux_bus_plus[0]);
    defparam vinPlus0__cy_connect_v1_0.sig_width = 1;
endmodule