module floating_point_v5_0 (
  clk, a, b, operation, result
)/* synthesis syn_black_box syn_noprune=1 */;
  input clk;
  input [63 : 0] a;
  input [63 : 0] b;
  input [5 : 0] operation;
  output [63 : 0] result;
  // synthesis translate_off
  wire \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/sign_op ;
  wire sig00000001;
  wire sig00000002;
  wire sig00000003;
  wire sig00000004;
  wire sig00000005;
  wire sig00000006;
  wire sig00000007;
  wire sig00000008;
  wire sig00000009;
  wire sig0000000a;
  wire sig0000000b;
  wire sig0000000c;
  wire sig0000000d;
  wire sig0000000e;
  wire sig0000000f;
  wire sig00000010;
  wire sig00000011;
  wire sig00000012;
  wire sig00000013;
  wire sig00000014;
  wire sig00000015;
  wire sig00000016;
  wire sig00000017;
  wire sig00000018;
  wire sig00000019;
  wire sig0000001a;
  wire sig0000001b;
  wire sig0000001c;
  wire sig0000001d;
  wire sig0000001e;
  wire sig0000001f;
  wire sig00000020;
  wire sig00000021;
  wire sig00000022;
  wire sig00000023;
  wire sig00000024;
  wire sig00000025;
  wire sig00000026;
  wire sig00000027;
  wire sig00000028;
  wire sig00000029;
  wire sig0000002a;
  wire sig0000002b;
  wire sig0000002c;
  wire sig0000002d;
  wire sig0000002e;
  wire sig0000002f;
  wire sig00000030;
  wire sig00000031;
  wire sig00000032;
  wire sig00000033;
  wire sig00000034;
  wire sig00000035;
  wire sig00000036;
  wire sig00000037;
  wire sig00000038;
  wire sig00000039;
  wire sig0000003a;
  wire sig0000003b;
  wire sig0000003c;
  wire sig0000003d;
  wire sig0000003e;
  wire sig0000003f;
  wire sig00000040;
  wire sig00000041;
  wire sig00000042;
  wire sig00000043;
  wire sig00000044;
  wire sig00000045;
  wire sig00000046;
  wire sig00000047;
  wire sig00000048;
  wire sig00000049;
  wire sig0000004a;
  wire sig0000004b;
  wire sig0000004c;
  wire sig0000004d;
  wire sig0000004e;
  wire sig0000004f;
  wire sig00000050;
  wire sig00000051;
  wire sig00000052;
  wire sig00000053;
  wire sig00000054;
  wire sig00000055;
  wire sig00000056;
  wire sig00000057;
  wire sig00000058;
  wire sig00000059;
  wire sig0000005a;
  wire sig0000005b;
  wire sig0000005c;
  wire sig0000005d;
  wire sig0000005e;
  wire sig0000005f;
  wire sig00000060;
  wire sig00000061;
  wire sig00000062;
  wire sig00000063;
  wire sig00000064;
  wire sig00000065;
  wire sig00000066;
  wire sig00000067;
  wire sig00000068;
  wire sig00000069;
  wire sig0000006a;
  wire sig0000006b;
  wire sig0000006c;
  wire sig0000006d;
  wire sig0000006e;
  wire sig0000006f;
  wire sig00000070;
  wire sig00000071;
  wire sig00000072;
  wire sig00000073;
  wire sig00000074;
  wire sig00000075;
  wire sig00000076;
  wire sig00000077;
  wire sig00000078;
  wire sig00000079;
  wire sig0000007a;
  wire sig0000007b;
  wire sig0000007c;
  wire sig0000007d;
  wire sig0000007e;
  wire sig0000007f;
  wire sig00000080;
  wire sig00000081;
  wire sig00000082;
  wire sig00000083;
  wire sig00000084;
  wire sig00000085;
  wire sig00000086;
  wire sig00000087;
  wire sig00000088;
  wire sig00000089;
  wire sig0000008a;
  wire sig0000008b;
  wire sig0000008c;
  wire sig0000008d;
  wire sig0000008e;
  wire sig0000008f;
  wire sig00000090;
  wire sig00000091;
  wire sig00000092;
  wire sig00000093;
  wire sig00000094;
  wire sig00000095;
  wire sig00000096;
  wire sig00000097;
  wire sig00000098;
  wire sig00000099;
  wire sig0000009a;
  wire sig0000009b;
  wire sig0000009c;
  wire sig0000009d;
  wire sig0000009e;
  wire sig0000009f;
  wire sig000000a0;
  wire sig000000a1;
  wire sig000000a2;
  wire sig000000a3;
  wire sig000000a4;
  wire sig000000a5;
  wire sig000000a6;
  wire sig000000a7;
  wire sig000000a8;
  wire sig000000a9;
  wire sig000000aa;
  wire sig000000ab;
  wire sig000000ac;
  wire sig000000ad;
  wire sig000000ae;
  wire sig000000af;
  wire sig000000b0;
  wire sig000000b1;
  wire sig000000b2;
  wire sig000000b3;
  wire sig000000b4;
  wire sig000000b5;
  wire sig000000b6;
  wire sig000000b7;
  wire sig000000b8;
  wire sig000000b9;
  wire sig000000ba;
  wire sig000000bb;
  wire sig000000bc;
  wire sig000000bd;
  wire sig000000be;
  wire sig000000bf;
  wire sig000000c0;
  wire sig000000c1;
  wire sig000000c2;
  wire sig000000c3;
  wire sig000000c4;
  wire sig000000c5;
  wire sig000000c6;
  wire sig000000c7;
  wire sig000000c8;
  wire sig000000c9;
  wire sig000000ca;
  wire sig000000cb;
  wire sig000000cc;
  wire sig000000cd;
  wire sig000000ce;
  wire sig000000cf;
  wire sig000000d0;
  wire sig000000d1;
  wire sig000000d2;
  wire sig000000d3;
  wire sig000000d4;
  wire sig000000d5;
  wire sig000000d6;
  wire sig000000d7;
  wire sig000000d8;
  wire sig000000d9;
  wire sig000000da;
  wire sig000000db;
  wire sig000000dc;
  wire sig000000dd;
  wire sig000000de;
  wire sig000000df;
  wire sig000000e0;
  wire sig000000e1;
  wire sig000000e2;
  wire sig000000e3;
  wire sig000000e4;
  wire sig000000e5;
  wire sig000000e6;
  wire sig000000e7;
  wire sig000000e8;
  wire sig000000e9;
  wire sig000000ea;
  wire sig000000eb;
  wire sig000000ec;
  wire sig000000ed;
  wire sig000000ee;
  wire sig000000ef;
  wire sig000000f0;
  wire sig000000f1;
  wire sig000000f2;
  wire sig000000f3;
  wire sig000000f4;
  wire sig000000f5;
  wire sig000000f6;
  wire sig000000f7;
  wire sig000000f8;
  wire sig000000f9;
  wire sig000000fa;
  wire sig000000fb;
  wire sig000000fc;
  wire sig000000fd;
  wire sig000000fe;
  wire sig000000ff;
  wire sig00000100;
  wire sig00000101;
  wire sig00000102;
  wire sig00000103;
  wire sig00000104;
  wire sig00000105;
  wire sig00000106;
  wire sig00000107;
  wire sig00000108;
  wire sig00000109;
  wire sig0000010a;
  wire sig0000010b;
  wire sig0000010c;
  wire sig0000010d;
  wire sig0000010e;
  wire sig0000010f;
  wire sig00000110;
  wire sig00000111;
  wire sig00000112;
  wire sig00000113;
  wire sig00000114;
  wire sig00000115;
  wire sig00000116;
  wire sig00000117;
  wire sig00000118;
  wire sig00000119;
  wire sig0000011a;
  wire sig0000011b;
  wire sig0000011c;
  wire sig0000011d;
  wire sig0000011e;
  wire sig0000011f;
  wire sig00000120;
  wire sig00000121;
  wire sig00000122;
  wire sig00000123;
  wire sig00000124;
  wire sig00000125;
  wire sig00000126;
  wire sig00000127;
  wire sig00000128;
  wire sig00000129;
  wire sig0000012a;
  wire sig0000012b;
  wire sig0000012c;
  wire sig0000012d;
  wire sig0000012e;
  wire sig0000012f;
  wire sig00000130;
  wire sig00000131;
  wire sig00000132;
  wire sig00000133;
  wire sig00000134;
  wire sig00000135;
  wire sig00000136;
  wire sig00000137;
  wire sig00000138;
  wire sig00000139;
  wire sig0000013a;
  wire sig0000013b;
  wire sig0000013c;
  wire sig0000013d;
  wire sig0000013e;
  wire sig0000013f;
  wire sig00000140;
  wire sig00000141;
  wire sig00000142;
  wire sig00000143;
  wire sig00000144;
  wire sig00000145;
  wire sig00000146;
  wire sig00000147;
  wire sig00000148;
  wire sig00000149;
  wire sig0000014a;
  wire sig0000014b;
  wire sig0000014c;
  wire sig0000014d;
  wire sig0000014e;
  wire sig0000014f;
  wire sig00000150;
  wire sig00000151;
  wire sig00000152;
  wire sig00000153;
  wire sig00000154;
  wire sig00000155;
  wire sig00000156;
  wire sig00000157;
  wire sig00000158;
  wire sig00000159;
  wire sig0000015a;
  wire sig0000015b;
  wire sig0000015c;
  wire sig0000015d;
  wire sig0000015e;
  wire sig0000015f;
  wire sig00000160;
  wire sig00000161;
  wire sig00000162;
  wire sig00000163;
  wire sig00000164;
  wire sig00000165;
  wire sig00000166;
  wire sig00000167;
  wire sig00000168;
  wire sig00000169;
  wire sig0000016a;
  wire sig0000016b;
  wire sig0000016c;
  wire sig0000016d;
  wire sig0000016e;
  wire sig0000016f;
  wire sig00000170;
  wire sig00000171;
  wire sig00000172;
  wire sig00000173;
  wire sig00000174;
  wire sig00000175;
  wire sig00000176;
  wire sig00000177;
  wire sig00000178;
  wire sig00000179;
  wire sig0000017a;
  wire sig0000017b;
  wire sig0000017c;
  wire sig0000017d;
  wire sig0000017e;
  wire sig0000017f;
  wire sig00000180;
  wire sig00000181;
  wire sig00000182;
  wire sig00000183;
  wire sig00000184;
  wire sig00000185;
  wire sig00000186;
  wire sig00000187;
  wire sig00000188;
  wire sig00000189;
  wire sig0000018a;
  wire sig0000018b;
  wire sig0000018c;
  wire sig0000018d;
  wire sig0000018e;
  wire sig0000018f;
  wire sig00000190;
  wire sig00000191;
  wire sig00000192;
  wire sig00000193;
  wire sig00000194;
  wire sig00000195;
  wire sig00000196;
  wire sig00000197;
  wire sig00000198;
  wire sig00000199;
  wire sig0000019a;
  wire sig0000019b;
  wire sig0000019c;
  wire sig0000019d;
  wire sig0000019e;
  wire sig0000019f;
  wire sig000001a0;
  wire sig000001a1;
  wire sig000001a2;
  wire sig000001a3;
  wire sig000001a4;
  wire sig000001a5;
  wire sig000001a6;
  wire sig000001a7;
  wire sig000001a8;
  wire sig000001a9;
  wire sig000001aa;
  wire sig000001ab;
  wire sig000001ac;
  wire sig000001ad;
  wire sig000001ae;
  wire sig000001af;
  wire sig000001b0;
  wire sig000001b1;
  wire sig000001b2;
  wire sig000001b3;
  wire sig000001b4;
  wire sig000001b5;
  wire sig000001b6;
  wire sig000001b7;
  wire sig000001b8;
  wire sig000001b9;
  wire sig000001ba;
  wire sig000001bb;
  wire sig000001bc;
  wire sig000001bd;
  wire sig000001be;
  wire sig000001bf;
  wire sig000001c0;
  wire sig000001c1;
  wire sig000001c2;
  wire sig000001c3;
  wire sig000001c4;
  wire sig000001c5;
  wire sig000001c6;
  wire sig000001c7;
  wire sig000001c8;
  wire sig000001c9;
  wire sig000001ca;
  wire sig000001cb;
  wire sig000001cc;
  wire sig000001cd;
  wire sig000001ce;
  wire sig000001cf;
  wire sig000001d0;
  wire sig000001d1;
  wire sig000001d2;
  wire sig000001d3;
  wire sig000001d4;
  wire sig000001d5;
  wire sig000001d6;
  wire sig000001d7;
  wire sig000001d8;
  wire sig000001d9;
  wire sig000001da;
  wire sig000001db;
  wire sig000001dc;
  wire sig000001dd;
  wire sig000001de;
  wire sig000001df;
  wire sig000001e0;
  wire sig000001e1;
  wire sig000001e2;
  wire sig000001e3;
  wire sig000001e4;
  wire sig000001e5;
  wire sig000001e6;
  wire sig000001e7;
  wire sig000001e8;
  wire sig000001e9;
  wire sig000001ea;
  wire sig000001eb;
  wire sig000001ec;
  wire sig000001ed;
  wire sig000001ee;
  wire sig000001ef;
  wire sig000001f0;
  wire sig000001f1;
  wire sig000001f2;
  wire sig000001f3;
  wire sig000001f4;
  wire sig000001f5;
  wire sig000001f6;
  wire sig000001f7;
  wire sig000001f8;
  wire sig000001f9;
  wire sig000001fa;
  wire sig000001fb;
  wire sig000001fc;
  wire sig000001fd;
  wire sig000001fe;
  wire sig000001ff;
  wire sig00000200;
  wire sig00000201;
  wire sig00000202;
  wire sig00000203;
  wire sig00000204;
  wire sig00000205;
  wire sig00000206;
  wire sig00000207;
  wire sig00000208;
  wire sig00000209;
  wire sig0000020a;
  wire sig0000020b;
  wire sig0000020c;
  wire sig0000020d;
  wire sig0000020e;
  wire sig0000020f;
  wire sig00000210;
  wire sig00000211;
  wire sig00000212;
  wire sig00000213;
  wire sig00000214;
  wire sig00000215;
  wire sig00000216;
  wire sig00000217;
  wire sig00000218;
  wire sig00000219;
  wire sig0000021a;
  wire sig0000021b;
  wire sig0000021c;
  wire sig0000021d;
  wire sig0000021e;
  wire sig0000021f;
  wire sig00000220;
  wire sig00000221;
  wire sig00000222;
  wire sig00000223;
  wire sig00000224;
  wire sig00000225;
  wire sig00000226;
  wire sig00000227;
  wire sig00000228;
  wire sig00000229;
  wire sig0000022a;
  wire sig0000022b;
  wire sig0000022c;
  wire sig0000022d;
  wire sig0000022e;
  wire sig0000022f;
  wire sig00000230;
  wire sig00000231;
  wire sig00000232;
  wire sig00000233;
  wire sig00000234;
  wire sig00000235;
  wire sig00000236;
  wire sig00000237;
  wire sig00000238;
  wire sig00000239;
  wire sig0000023a;
  wire sig0000023b;
  wire sig0000023c;
  wire sig0000023d;
  wire sig0000023e;
  wire sig0000023f;
  wire sig00000240;
  wire sig00000241;
  wire sig00000242;
  wire sig00000243;
  wire sig00000244;
  wire sig00000245;
  wire sig00000246;
  wire sig00000247;
  wire sig00000248;
  wire sig00000249;
  wire sig0000024a;
  wire sig0000024b;
  wire sig0000024c;
  wire sig0000024d;
  wire sig0000024e;
  wire sig0000024f;
  wire sig00000250;
  wire sig00000251;
  wire sig00000252;
  wire sig00000253;
  wire sig00000254;
  wire sig00000255;
  wire sig00000256;
  wire sig00000257;
  wire sig00000258;
  wire sig00000259;
  wire sig0000025a;
  wire sig0000025b;
  wire sig0000025c;
  wire sig0000025d;
  wire sig0000025e;
  wire sig0000025f;
  wire sig00000260;
  wire sig00000261;
  wire sig00000262;
  wire sig00000263;
  wire sig00000264;
  wire sig00000265;
  wire sig00000266;
  wire sig00000267;
  wire sig00000268;
  wire sig00000269;
  wire sig0000026a;
  wire sig0000026b;
  wire sig0000026c;
  wire sig0000026d;
  wire sig0000026e;
  wire sig0000026f;
  wire sig00000270;
  wire sig00000271;
  wire sig00000272;
  wire sig00000273;
  wire sig00000274;
  wire sig00000275;
  wire sig00000276;
  wire sig00000277;
  wire sig00000278;
  wire sig00000279;
  wire sig0000027a;
  wire sig0000027b;
  wire sig0000027c;
  wire sig0000027d;
  wire sig0000027e;
  wire sig0000027f;
  wire sig00000280;
  wire sig00000281;
  wire sig00000282;
  wire sig00000283;
  wire sig00000284;
  wire sig00000285;
  wire sig00000286;
  wire sig00000287;
  wire sig00000288;
  wire sig00000289;
  wire sig0000028a;
  wire sig0000028b;
  wire sig0000028c;
  wire sig0000028d;
  wire sig0000028e;
  wire sig0000028f;
  wire sig00000290;
  wire sig00000291;
  wire sig00000292;
  wire sig00000293;
  wire sig00000294;
  wire sig00000295;
  wire sig00000296;
  wire sig00000297;
  wire sig00000298;
  wire sig00000299;
  wire sig0000029a;
  wire sig0000029b;
  wire sig0000029c;
  wire sig0000029d;
  wire sig0000029e;
  wire sig0000029f;
  wire sig000002a0;
  wire sig000002a1;
  wire sig000002a2;
  wire sig000002a3;
  wire sig000002a4;
  wire sig000002a5;
  wire sig000002a6;
  wire sig000002a7;
  wire sig000002a8;
  wire sig000002a9;
  wire sig000002aa;
  wire sig000002ab;
  wire sig000002ac;
  wire sig000002ad;
  wire sig000002ae;
  wire sig000002af;
  wire sig000002b0;
  wire sig000002b1;
  wire sig000002b2;
  wire sig000002b3;
  wire sig000002b4;
  wire sig000002b5;
  wire sig000002b6;
  wire sig000002b7;
  wire sig000002b8;
  wire sig000002b9;
  wire sig000002ba;
  wire sig000002bb;
  wire sig000002bc;
  wire sig000002bd;
  wire sig000002be;
  wire sig000002bf;
  wire sig000002c0;
  wire sig000002c1;
  wire sig000002c2;
  wire sig000002c3;
  wire sig000002c4;
  wire sig000002c5;
  wire sig000002c6;
  wire sig000002c7;
  wire sig000002c8;
  wire sig000002c9;
  wire sig000002ca;
  wire sig000002cb;
  wire sig000002cc;
  wire sig000002cd;
  wire sig000002ce;
  wire sig000002cf;
  wire sig000002d0;
  wire sig000002d1;
  wire sig000002d2;
  wire sig000002d3;
  wire sig000002d4;
  wire sig000002d5;
  wire sig000002d6;
  wire sig000002d7;
  wire sig000002d8;
  wire sig000002d9;
  wire sig000002da;
  wire sig000002db;
  wire sig000002dc;
  wire sig000002dd;
  wire sig000002de;
  wire sig000002df;
  wire sig000002e0;
  wire sig000002e1;
  wire sig000002e2;
  wire sig000002e3;
  wire sig000002e4;
  wire sig000002e5;
  wire sig000002e6;
  wire sig000002e7;
  wire sig000002e8;
  wire sig000002e9;
  wire sig000002ea;
  wire sig000002eb;
  wire sig000002ec;
  wire sig000002ed;
  wire sig000002ee;
  wire sig000002ef;
  wire sig000002f0;
  wire sig000002f1;
  wire sig000002f2;
  wire sig000002f3;
  wire sig000002f4;
  wire sig000002f5;
  wire sig000002f6;
  wire sig000002f7;
  wire sig000002f8;
  wire sig000002f9;
  wire sig000002fa;
  wire sig000002fb;
  wire sig000002fc;
  wire sig000002fd;
  wire sig000002fe;
  wire sig000002ff;
  wire sig00000300;
  wire sig00000301;
  wire sig00000302;
  wire sig00000303;
  wire sig00000304;
  wire sig00000305;
  wire sig00000306;
  wire sig00000307;
  wire sig00000308;
  wire sig00000309;
  wire sig0000030a;
  wire sig0000030b;
  wire sig0000030c;
  wire sig0000030d;
  wire sig0000030e;
  wire sig0000030f;
  wire sig00000310;
  wire sig00000311;
  wire sig00000312;
  wire sig00000313;
  wire sig00000314;
  wire sig00000315;
  wire sig00000316;
  wire sig00000317;
  wire sig00000318;
  wire sig00000319;
  wire sig0000031a;
  wire sig0000031b;
  wire sig0000031c;
  wire sig0000031d;
  wire sig0000031e;
  wire sig0000031f;
  wire sig00000320;
  wire sig00000321;
  wire sig00000322;
  wire sig00000323;
  wire sig00000324;
  wire sig00000325;
  wire sig00000326;
  wire sig00000327;
  wire sig00000328;
  wire sig00000329;
  wire sig0000032a;
  wire sig0000032b;
  wire sig0000032c;
  wire sig0000032d;
  wire sig0000032e;
  wire sig0000032f;
  wire sig00000330;
  wire sig00000331;
  wire sig00000332;
  wire sig00000333;
  wire sig00000334;
  wire sig00000335;
  wire sig00000336;
  wire sig00000337;
  wire sig00000338;
  wire sig00000339;
  wire sig0000033a;
  wire sig0000033b;
  wire sig0000033c;
  wire sig0000033d;
  wire sig0000033e;
  wire sig0000033f;
  wire sig00000340;
  wire sig00000341;
  wire sig00000342;
  wire sig00000343;
  wire sig00000344;
  wire sig00000345;
  wire sig00000346;
  wire sig00000347;
  wire sig00000348;
  wire sig00000349;
  wire sig0000034a;
  wire sig0000034b;
  wire sig0000034c;
  wire sig0000034d;
  wire sig0000034e;
  wire sig0000034f;
  wire sig00000350;
  wire sig00000351;
  wire sig00000352;
  wire sig00000353;
  wire sig00000354;
  wire sig00000355;
  wire sig00000356;
  wire sig00000357;
  wire sig00000358;
  wire sig00000359;
  wire sig0000035a;
  wire sig0000035b;
  wire sig0000035c;
  wire sig0000035d;
  wire sig0000035e;
  wire sig0000035f;
  wire sig00000360;
  wire sig00000361;
  wire sig00000362;
  wire sig00000363;
  wire sig00000364;
  wire sig00000365;
  wire sig00000366;
  wire sig00000367;
  wire sig00000368;
  wire sig00000369;
  wire sig0000036a;
  wire sig0000036b;
  wire sig0000036c;
  wire sig0000036d;
  wire sig0000036e;
  wire sig0000036f;
  wire sig00000370;
  wire sig00000371;
  wire sig00000372;
  wire sig00000373;
  wire sig00000374;
  wire sig00000375;
  wire sig00000376;
  wire sig00000377;
  wire sig00000378;
  wire sig00000379;
  wire sig0000037a;
  wire sig0000037b;
  wire sig0000037c;
  wire sig0000037d;
  wire sig0000037e;
  wire sig0000037f;
  wire sig00000380;
  wire sig00000381;
  wire sig00000382;
  wire sig00000383;
  wire sig00000384;
  wire sig00000385;
  wire sig00000386;
  wire sig00000387;
  wire sig00000388;
  wire sig00000389;
  wire sig0000038a;
  wire sig0000038b;
  wire sig0000038c;
  wire sig0000038d;
  wire sig0000038e;
  wire sig0000038f;
  wire sig00000390;
  wire sig00000391;
  wire sig00000392;
  wire sig00000393;
  wire sig00000394;
  wire sig00000395;
  wire sig00000396;
  wire sig00000397;
  wire sig00000398;
  wire sig00000399;
  wire sig0000039a;
  wire sig0000039b;
  wire sig0000039c;
  wire sig0000039d;
  wire sig0000039e;
  wire sig0000039f;
  wire sig000003a0;
  wire sig000003a1;
  wire sig000003a2;
  wire sig000003a3;
  wire sig000003a4;
  wire sig000003a5;
  wire sig000003a6;
  wire sig000003a7;
  wire sig000003a8;
  wire sig000003a9;
  wire sig000003aa;
  wire sig000003ab;
  wire sig000003ac;
  wire sig000003ad;
  wire sig000003ae;
  wire sig000003af;
  wire sig000003b0;
  wire sig000003b1;
  wire sig000003b2;
  wire sig000003b3;
  wire sig000003b4;
  wire sig000003b5;
  wire sig000003b6;
  wire sig000003b7;
  wire sig000003b8;
  wire sig000003b9;
  wire sig000003ba;
  wire sig000003bb;
  wire sig000003bc;
  wire sig000003bd;
  wire sig000003be;
  wire sig000003bf;
  wire sig000003c0;
  wire sig000003c1;
  wire sig000003c2;
  wire sig000003c3;
  wire sig000003c4;
  wire sig000003c5;
  wire sig000003c6;
  wire sig000003c7;
  wire sig000003c8;
  wire sig000003c9;
  wire sig000003ca;
  wire sig000003cb;
  wire sig000003cc;
  wire sig000003cd;
  wire sig000003ce;
  wire sig000003cf;
  wire sig000003d0;
  wire sig000003d1;
  wire sig000003d2;
  wire sig000003d3;
  wire sig000003d4;
  wire sig000003d5;
  wire sig000003d6;
  wire sig000003d7;
  wire sig000003d8;
  wire sig000003d9;
  wire sig000003da;
  wire sig000003db;
  wire sig000003dc;
  wire sig000003dd;
  wire sig000003de;
  wire sig000003df;
  wire sig000003e0;
  wire sig000003e1;
  wire sig000003e2;
  wire sig000003e3;
  wire sig000003e4;
  wire sig000003e5;
  wire sig000003e6;
  wire sig000003e7;
  wire sig000003e8;
  wire sig000003e9;
  wire sig000003ea;
  wire sig000003eb;
  wire sig000003ec;
  wire sig000003ed;
  wire sig000003ee;
  wire sig000003ef;
  wire sig000003f0;
  wire sig000003f1;
  wire sig000003f2;
  wire sig000003f3;
  wire sig000003f4;
  wire sig000003f5;
  wire sig000003f6;
  wire sig000003f7;
  wire sig000003f8;
  wire sig000003f9;
  wire sig000003fa;
  wire sig000003fb;
  wire sig000003fc;
  wire sig000003fd;
  wire sig000003fe;
  wire sig000003ff;
  wire sig00000400;
  wire sig00000401;
  wire sig00000402;
  wire sig00000403;
  wire sig00000404;
  wire sig00000405;
  wire sig00000406;
  wire sig00000407;
  wire sig00000408;
  wire sig00000409;
  wire sig0000040a;
  wire sig0000040b;
  wire sig0000040c;
  wire sig0000040d;
  wire sig0000040e;
  wire sig0000040f;
  wire sig00000410;
  wire sig00000411;
  wire sig00000412;
  wire sig00000413;
  wire sig00000414;
  wire sig00000415;
  wire sig00000416;
  wire sig00000417;
  wire sig00000418;
  wire sig00000419;
  wire sig0000041a;
  wire sig0000041b;
  wire sig0000041c;
  wire sig0000041d;
  wire sig0000041e;
  wire sig0000041f;
  wire sig00000420;
  wire sig00000421;
  wire sig00000422;
  wire sig00000423;
  wire sig00000424;
  wire sig00000425;
  wire sig00000426;
  wire sig00000427;
  wire sig00000428;
  wire sig00000429;
  wire sig0000042a;
  wire sig0000042b;
  wire sig0000042c;
  wire sig0000042d;
  wire sig0000042e;
  wire sig0000042f;
  wire sig00000430;
  wire sig00000431;
  wire sig00000432;
  wire sig00000433;
  wire sig00000434;
  wire sig00000435;
  wire sig00000436;
  wire sig00000437;
  wire sig00000438;
  wire sig00000439;
  wire sig0000043a;
  wire sig0000043b;
  wire sig0000043c;
  wire sig0000043d;
  wire sig0000043e;
  wire sig0000043f;
  wire sig00000440;
  wire sig00000441;
  wire sig00000442;
  wire sig00000443;
  wire sig00000444;
  wire sig00000445;
  wire sig00000446;
  wire sig00000447;
  wire sig00000448;
  wire sig00000449;
  wire sig0000044a;
  wire sig0000044b;
  wire sig0000044c;
  wire sig0000044d;
  wire sig0000044e;
  wire sig0000044f;
  wire sig00000450;
  wire sig00000451;
  wire sig00000452;
  wire sig00000453;
  wire sig00000454;
  wire sig00000455;
  wire sig00000456;
  wire sig00000457;
  wire sig00000458;
  wire sig00000459;
  wire sig0000045a;
  wire sig0000045b;
  wire sig0000045c;
  wire sig0000045d;
  wire sig0000045e;
  wire sig0000045f;
  wire sig00000460;
  wire sig00000461;
  wire sig00000462;
  wire sig00000463;
  wire sig00000464;
  wire sig00000465;
  wire sig00000466;
  wire sig00000467;
  wire sig00000468;
  wire sig00000469;
  wire sig0000046a;
  wire sig0000046b;
  wire sig0000046c;
  wire sig0000046d;
  wire sig0000046e;
  wire sig0000046f;
  wire sig00000470;
  wire sig00000471;
  wire sig00000472;
  wire sig00000473;
  wire sig00000474;
  wire sig00000475;
  wire sig00000476;
  wire sig00000477;
  wire sig00000478;
  wire sig00000479;
  wire sig0000047a;
  wire sig0000047b;
  wire sig0000047c;
  wire sig0000047d;
  wire sig0000047e;
  wire sig0000047f;
  wire sig00000480;
  wire sig00000481;
  wire sig00000482;
  wire sig00000483;
  wire sig00000484;
  wire sig00000485;
  wire sig00000486;
  wire sig00000487;
  wire sig00000488;
  wire sig00000489;
  wire sig0000048a;
  wire sig0000048b;
  wire sig0000048c;
  wire sig0000048d;
  wire sig0000048e;
  wire sig0000048f;
  wire sig00000490;
  wire sig00000491;
  wire sig00000492;
  wire sig00000493;
  wire sig00000494;
  wire sig00000495;
  wire sig00000496;
  wire sig00000497;
  wire sig00000498;
  wire sig00000499;
  wire sig0000049a;
  wire sig0000049b;
  wire sig0000049c;
  wire sig0000049d;
  wire sig0000049e;
  wire sig0000049f;
  wire sig000004a0;
  wire sig000004a1;
  wire sig000004a2;
  wire sig000004a3;
  wire sig000004a4;
  wire sig000004a5;
  wire sig000004a6;
  wire sig000004a7;
  wire sig000004a8;
  wire sig000004a9;
  wire sig000004aa;
  wire sig000004ab;
  wire sig000004ac;
  wire sig000004ad;
  wire sig000004ae;
  wire sig000004af;
  wire sig000004b0;
  wire sig000004b1;
  wire sig000004b2;
  wire sig000004b3;
  wire sig000004b4;
  wire sig000004b5;
  wire sig000004b6;
  wire sig000004b7;
  wire sig000004b8;
  wire sig000004b9;
  wire sig000004ba;
  wire sig000004bb;
  wire sig000004bc;
  wire sig000004bd;
  wire sig000004be;
  wire sig000004bf;
  wire sig000004c0;
  wire sig000004c1;
  wire sig000004c2;
  wire sig000004c3;
  wire sig000004c4;
  wire sig000004c5;
  wire sig000004c6;
  wire sig000004c7;
  wire sig000004c8;
  wire sig000004c9;
  wire sig000004ca;
  wire sig000004cb;
  wire sig000004cc;
  wire sig000004cd;
  wire sig000004ce;
  wire sig000004cf;
  wire sig000004d0;
  wire sig000004d1;
  wire sig000004d2;
  wire sig000004d3;
  wire sig000004d4;
  wire sig000004d5;
  wire sig000004d6;
  wire sig000004d7;
  wire sig000004d8;
  wire sig000004d9;
  wire sig000004da;
  wire sig000004db;
  wire sig000004dc;
  wire sig000004dd;
  wire sig000004de;
  wire sig000004df;
  wire sig000004e0;
  wire sig000004e1;
  wire sig000004e2;
  wire sig000004e3;
  wire sig000004e4;
  wire sig000004e5;
  wire sig000004e6;
  wire sig000004e7;
  wire sig000004e8;
  wire sig000004e9;
  wire sig000004ea;
  wire sig000004eb;
  wire sig000004ec;
  wire sig000004ed;
  wire sig000004ee;
  wire sig000004ef;
  wire sig000004f0;
  wire sig000004f1;
  wire sig000004f2;
  wire sig000004f3;
  wire sig000004f4;
  wire sig000004f5;
  wire sig000004f6;
  wire sig000004f7;
  wire sig000004f8;
  wire sig000004f9;
  wire sig000004fa;
  wire sig000004fb;
  wire sig000004fc;
  wire sig000004fd;
  wire sig000004fe;
  wire sig000004ff;
  wire sig00000500;
  wire sig00000501;
  wire sig00000502;
  wire sig00000503;
  wire sig00000504;
  wire sig00000505;
  wire sig00000506;
  wire sig00000507;
  wire sig00000508;
  wire sig00000509;
  wire sig0000050a;
  wire sig0000050b;
  wire sig0000050c;
  wire sig0000050d;
  wire sig0000050e;
  wire sig0000050f;
  wire sig00000510;
  wire sig00000511;
  wire sig00000512;
  wire sig00000513;
  wire sig00000514;
  wire sig00000515;
  wire sig00000516;
  wire sig00000517;
  wire sig00000518;
  wire sig00000519;
  wire sig0000051a;
  wire sig0000051b;
  wire sig0000051c;
  wire sig0000051d;
  wire sig0000051e;
  wire sig0000051f;
  wire sig00000520;
  wire sig00000521;
  wire sig00000522;
  wire sig00000523;
  wire sig00000524;
  wire sig00000525;
  wire sig00000526;
  wire sig00000527;
  wire sig00000528;
  wire sig00000529;
  wire sig0000052a;
  wire sig0000052b;
  wire sig0000052c;
  wire sig0000052d;
  wire sig0000052e;
  wire sig0000052f;
  wire sig00000530;
  wire sig00000531;
  wire sig00000532;
  wire sig00000533;
  wire sig00000534;
  wire sig00000535;
  wire sig00000536;
  wire sig00000537;
  wire sig00000538;
  wire sig00000539;
  wire sig0000053a;
  wire sig0000053b;
  wire sig0000053c;
  wire sig0000053d;
  wire sig0000053e;
  wire sig0000053f;
  wire sig00000540;
  wire sig00000541;
  wire sig00000542;
  wire sig00000543;
  wire sig00000544;
  wire sig00000545;
  wire sig00000546;
  wire sig00000547;
  wire sig00000548;
  wire sig00000549;
  wire sig0000054a;
  wire sig0000054b;
  wire sig0000054c;
  wire sig0000054d;
  wire sig0000054e;
  wire sig0000054f;
  wire sig00000550;
  wire sig00000551;
  wire sig00000552;
  wire sig00000553;
  wire sig00000554;
  wire sig00000555;
  wire sig00000556;
  wire sig00000557;
  wire sig00000558;
  wire sig00000559;
  wire sig0000055a;
  wire sig0000055b;
  wire sig0000055c;
  wire sig0000055d;
  wire sig0000055e;
  wire sig0000055f;
  wire sig00000560;
  wire sig00000561;
  wire sig00000562;
  wire sig00000563;
  wire sig00000564;
  wire sig00000565;
  wire sig00000566;
  wire sig00000567;
  wire sig00000568;
  wire sig00000569;
  wire sig0000056a;
  wire sig0000056b;
  wire sig0000056c;
  wire sig0000056d;
  wire sig0000056e;
  wire sig0000056f;
  wire sig00000570;
  wire sig00000571;
  wire sig00000572;
  wire sig00000573;
  wire sig00000574;
  wire sig00000575;
  wire sig00000576;
  wire sig00000577;
  wire sig00000578;
  wire sig00000579;
  wire sig0000057a;
  wire sig0000057b;
  wire sig0000057c;
  wire sig0000057d;
  wire sig0000057e;
  wire sig0000057f;
  wire sig00000580;
  wire sig00000581;
  wire sig00000582;
  wire sig00000583;
  wire sig00000584;
  wire sig00000585;
  wire sig00000586;
  wire sig00000587;
  wire sig00000588;
  wire sig00000589;
  wire sig0000058a;
  wire sig0000058b;
  wire sig0000058c;
  wire sig0000058d;
  wire sig0000058e;
  wire sig0000058f;
  wire sig00000590;
  wire sig00000591;
  wire sig00000592;
  wire sig00000593;
  wire sig00000594;
  wire sig00000595;
  wire sig00000596;
  wire sig00000597;
  wire sig00000598;
  wire sig00000599;
  wire sig0000059a;
  wire sig0000059b;
  wire sig0000059c;
  wire sig0000059d;
  wire sig0000059e;
  wire sig0000059f;
  wire sig000005a0;
  wire sig000005a1;
  wire sig000005a2;
  wire sig000005a3;
  wire sig000005a4;
  wire sig000005a5;
  wire sig000005a6;
  wire sig000005a7;
  wire sig000005a8;
  wire sig000005a9;
  wire sig000005aa;
  wire sig000005ab;
  wire sig000005ac;
  wire sig000005ad;
  wire sig000005ae;
  wire sig000005af;
  wire sig000005b0;
  wire sig000005b1;
  wire sig000005b2;
  wire sig000005b3;
  wire sig000005b4;
  wire sig000005b5;
  wire sig000005b6;
  wire sig000005b7;
  wire sig000005b8;
  wire sig000005b9;
  wire sig000005ba;
  wire sig000005bb;
  wire sig000005bc;
  wire sig000005bd;
  wire sig000005be;
  wire sig000005bf;
  wire sig000005c0;
  wire sig000005c1;
  wire sig000005c2;
  wire sig000005c3;
  wire sig000005c4;
  wire sig000005c5;
  wire sig000005c6;
  wire sig000005c7;
  wire sig000005c8;
  wire sig000005c9;
  wire sig000005ca;
  wire sig000005cb;
  wire sig000005cc;
  wire sig000005cd;
  wire sig000005ce;
  wire sig000005cf;
  wire sig000005d0;
  wire sig000005d1;
  wire sig000005d2;
  wire sig000005d3;
  wire sig000005d4;
  wire sig000005d5;
  wire sig000005d6;
  wire sig000005d7;
  wire sig000005d8;
  wire sig000005d9;
  wire sig000005da;
  wire sig000005db;
  wire sig000005dc;
  wire sig000005dd;
  wire sig000005de;
  wire sig000005df;
  wire sig000005e0;
  wire sig000005e1;
  wire sig000005e2;
  wire sig000005e3;
  wire sig000005e4;
  wire sig000005e5;
  wire sig000005e6;
  wire sig000005e7;
  wire sig000005e8;
  wire sig000005e9;
  wire sig000005ea;
  wire sig000005eb;
  wire sig000005ec;
  wire sig000005ed;
  wire sig000005ee;
  wire sig000005ef;
  wire sig000005f0;
  wire sig000005f1;
  wire sig000005f2;
  wire sig000005f3;
  wire sig000005f4;
  wire sig000005f5;
  wire sig000005f6;
  wire sig000005f7;
  wire sig000005f8;
  wire sig000005f9;
  wire sig000005fa;
  wire sig000005fb;
  wire sig000005fc;
  wire sig000005fd;
  wire sig000005fe;
  wire sig000005ff;
  wire sig00000600;
  wire sig00000601;
  wire sig00000602;
  wire sig00000603;
  wire sig00000604;
  wire sig00000605;
  wire sig00000606;
  wire sig00000607;
  wire sig00000608;
  wire sig00000609;
  wire sig0000060a;
  wire sig0000060b;
  wire sig0000060c;
  wire sig0000060d;
  wire sig0000060e;
  wire sig0000060f;
  wire sig00000610;
  wire sig00000611;
  wire sig00000612;
  wire sig00000613;
  wire sig00000614;
  wire sig00000615;
  wire sig00000616;
  wire sig00000617;
  wire sig00000618;
  wire sig00000619;
  wire sig0000061a;
  wire sig0000061b;
  wire sig0000061c;
  wire sig0000061d;
  wire sig0000061e;
  wire sig0000061f;
  wire sig00000620;
  wire sig00000621;
  wire sig00000622;
  wire sig00000623;
  wire sig00000624;
  wire sig00000625;
  wire sig00000626;
  wire sig00000627;
  wire sig00000628;
  wire sig00000629;
  wire sig0000062a;
  wire sig0000062b;
  wire sig0000062c;
  wire sig0000062d;
  wire sig0000062e;
  wire sig0000062f;
  wire sig00000630;
  wire sig00000631;
  wire sig00000632;
  wire sig00000633;
  wire sig00000634;
  wire sig00000635;
  wire sig00000636;
  wire sig00000637;
  wire sig00000638;
  wire sig00000639;
  wire sig0000063a;
  wire sig0000063b;
  wire sig0000063c;
  wire sig0000063d;
  wire sig0000063e;
  wire sig0000063f;
  wire sig00000640;
  wire sig00000641;
  wire sig00000642;
  wire sig00000643;
  wire sig00000644;
  wire sig00000645;
  wire sig00000646;
  wire sig00000647;
  wire sig00000648;
  wire sig00000649;
  wire sig0000064a;
  wire sig0000064b;
  wire sig0000064c;
  wire sig0000064d;
  wire sig0000064e;
  wire sig0000064f;
  wire sig00000650;
  wire sig00000651;
  wire sig00000652;
  wire sig00000653;
  wire sig00000654;
  wire sig00000655;
  wire sig00000656;
  wire sig00000657;
  wire sig00000658;
  wire sig00000659;
  wire sig0000065a;
  wire sig0000065b;
  wire sig0000065c;
  wire sig0000065d;
  wire sig0000065e;
  wire sig0000065f;
  wire sig00000660;
  wire sig00000661;
  wire sig00000662;
  wire sig00000663;
  wire sig00000664;
  wire sig00000665;
  wire sig00000666;
  wire sig00000667;
  wire sig00000668;
  wire sig00000669;
  wire sig0000066a;
  wire sig0000066b;
  wire sig0000066c;
  wire sig0000066d;
  wire sig0000066e;
  wire sig0000066f;
  wire sig00000670;
  wire sig00000671;
  wire sig00000672;
  wire sig00000673;
  wire sig00000674;
  wire sig00000675;
  wire sig00000676;
  wire sig00000677;
  wire sig00000678;
  wire sig00000679;
  wire sig0000067a;
  wire sig0000067b;
  wire sig0000067c;
  wire sig0000067d;
  wire sig0000067e;
  wire sig0000067f;
  wire sig00000680;
  wire sig00000681;
  wire sig00000682;
  wire sig00000683;
  wire sig00000684;
  wire sig00000685;
  wire sig00000686;
  wire sig00000687;
  wire sig00000688;
  wire sig00000689;
  wire sig0000068a;
  wire sig0000068b;
  wire sig0000068c;
  wire sig0000068d;
  wire sig0000068e;
  wire sig0000068f;
  wire sig00000690;
  wire sig00000691;
  wire sig00000692;
  wire sig00000693;
  wire sig00000694;
  wire sig00000695;
  wire sig00000696;
  wire sig00000697;
  wire sig00000698;
  wire sig00000699;
  wire sig0000069a;
  wire sig0000069b;
  wire sig0000069c;
  wire sig0000069d;
  wire sig0000069e;
  wire sig0000069f;
  wire sig000006a0;
  wire sig000006a1;
  wire sig000006a2;
  wire sig000006a3;
  wire sig000006a4;
  wire sig000006a5;
  wire sig000006a6;
  wire sig000006a7;
  wire sig000006a8;
  wire sig000006a9;
  wire sig000006aa;
  wire sig000006ab;
  wire sig000006ac;
  wire sig000006ad;
  wire sig000006ae;
  wire sig000006af;
  wire sig000006b0;
  wire sig000006b1;
  wire sig000006b2;
  wire sig000006b3;
  wire sig000006b4;
  wire sig000006b5;
  wire sig000006b6;
  wire sig000006b7;
  wire sig000006b8;
  wire sig000006b9;
  wire sig000006ba;
  wire sig000006bb;
  wire sig000006bc;
  wire sig000006bd;
  wire sig000006be;
  wire sig000006bf;
  wire sig000006c0;
  wire sig000006c1;
  wire sig000006c2;
  wire sig000006c3;
  wire sig000006c4;
  wire sig000006c5;
  wire sig000006c6;
  wire sig000006c7;
  wire sig000006c8;
  wire sig000006c9;
  wire sig000006ca;
  wire sig000006cb;
  wire sig000006cc;
  wire sig000006cd;
  wire sig000006ce;
  wire sig000006cf;
  wire sig000006d0;
  wire sig000006d1;
  wire sig000006d2;
  wire sig000006d3;
  wire sig000006d4;
  wire sig000006d5;
  wire sig000006d6;
  wire sig000006d7;
  wire sig000006d8;
  wire sig000006d9;
  wire sig000006da;
  wire sig000006db;
  wire sig000006dc;
  wire sig000006dd;
  wire sig000006de;
  wire sig000006df;
  wire sig000006e0;
  wire sig000006e1;
  wire sig000006e2;
  wire sig000006e3;
  wire sig000006e4;
  wire sig000006e5;
  wire sig000006e6;
  wire sig000006e7;
  wire sig000006e8;
  wire sig000006e9;
  wire sig000006ea;
  wire sig000006eb;
  wire sig000006ec;
  wire sig000006ed;
  wire sig000006ee;
  wire sig000006ef;
  wire sig000006f0;
  wire sig000006f1;
  wire sig000006f2;
  wire sig000006f3;
  wire sig000006f4;
  wire sig000006f5;
  wire sig000006f6;
  wire sig000006f7;
  wire sig000006f8;
  wire sig000006f9;
  wire sig000006fa;
  wire sig000006fb;
  wire sig000006fc;
  wire sig000006fd;
  wire sig000006fe;
  wire sig000006ff;
  wire sig00000700;
  wire sig00000701;
  wire sig00000702;
  wire sig00000703;
  wire sig00000704;
  wire sig00000705;
  wire sig00000706;
  wire sig00000707;
  wire sig00000708;
  wire sig00000709;
  wire sig0000070a;
  wire sig0000070b;
  wire sig0000070c;
  wire sig0000070d;
  wire sig0000070e;
  wire sig0000070f;
  wire sig00000710;
  wire sig00000711;
  wire sig00000712;
  wire sig00000713;
  wire sig00000714;
  wire sig00000715;
  wire sig00000716;
  wire sig00000717;
  wire sig00000718;
  wire sig00000719;
  wire sig0000071a;
  wire sig0000071b;
  wire sig0000071c;
  wire sig0000071d;
  wire sig0000071e;
  wire sig0000071f;
  wire sig00000720;
  wire sig00000721;
  wire sig00000722;
  wire sig00000723;
  wire sig00000724;
  wire sig00000725;
  wire sig00000726;
  wire sig00000727;
  wire sig00000728;
  wire sig00000729;
  wire sig0000072a;
  wire sig0000072b;
  wire sig0000072c;
  wire sig0000072d;
  wire sig0000072e;
  wire sig0000072f;
  wire sig00000730;
  wire sig00000731;
  wire sig00000732;
  wire sig00000733;
  wire sig00000734;
  wire sig00000735;
  wire sig00000736;
  wire sig00000737;
  wire sig00000738;
  wire sig00000739;
  wire sig0000073a;
  wire sig0000073b;
  wire sig0000073c;
  wire sig0000073d;
  wire sig0000073e;
  wire sig0000073f;
  wire sig00000740;
  wire sig00000741;
  wire sig00000742;
  wire sig00000743;
  wire sig00000744;
  wire sig00000745;
  wire sig00000746;
  wire sig00000747;
  wire sig00000748;
  wire sig00000749;
  wire sig0000074a;
  wire sig0000074b;
  wire sig0000074c;
  wire sig0000074d;
  wire sig0000074e;
  wire sig0000074f;
  wire sig00000750;
  wire sig00000751;
  wire sig00000752;
  wire sig00000753;
  wire sig00000754;
  wire sig00000755;
  wire sig00000756;
  wire sig00000757;
  wire sig00000758;
  wire sig00000759;
  wire sig0000075a;
  wire sig0000075b;
  wire sig0000075c;
  wire sig0000075d;
  wire sig0000075e;
  wire sig0000075f;
  wire sig00000760;
  wire sig00000761;
  wire sig00000762;
  wire sig00000763;
  wire sig00000764;
  wire sig00000765;
  wire sig00000766;
  wire sig00000767;
  wire sig00000768;
  wire sig00000769;
  wire sig0000076a;
  wire sig0000076b;
  wire sig0000076c;
  wire sig0000076d;
  wire sig0000076e;
  wire sig0000076f;
  wire sig00000770;
  wire sig00000771;
  wire sig00000772;
  wire sig00000773;
  wire sig00000774;
  wire sig00000775;
  wire sig00000776;
  wire sig00000777;
  wire sig00000778;
  wire sig00000779;
  wire sig0000077a;
  wire sig0000077b;
  wire sig0000077c;
  wire sig0000077d;
  wire sig0000077e;
  wire sig0000077f;
  wire sig00000780;
  wire sig00000781;
  wire sig00000782;
  wire sig00000783;
  wire sig00000784;
  wire sig00000785;
  wire sig00000786;
  wire sig00000787;
  wire sig00000788;
  wire sig00000789;
  wire sig0000078a;
  wire sig0000078b;
  wire sig0000078c;
  wire sig0000078d;
  wire sig0000078e;
  wire sig0000078f;
  wire sig00000790;
  wire sig00000791;
  wire sig00000792;
  wire sig00000793;
  wire sig00000794;
  wire sig00000795;
  wire sig00000796;
  wire sig00000797;
  wire sig00000798;
  wire sig00000799;
  wire sig0000079a;
  wire sig0000079b;
  wire sig0000079c;
  wire sig0000079d;
  wire sig0000079e;
  wire sig0000079f;
  wire sig000007a0;
  wire sig000007a1;
  wire sig000007a2;
  wire sig000007a3;
  wire sig000007a4;
  wire sig000007a5;
  wire sig000007a6;
  wire sig000007a7;
  wire sig000007a8;
  wire sig000007a9;
  wire sig000007aa;
  wire sig000007ab;
  wire sig000007ac;
  wire sig000007ad;
  wire sig000007ae;
  wire sig000007af;
  wire sig000007b0;
  wire sig000007b1;
  wire sig000007b2;
  wire sig000007b3;
  wire sig000007b4;
  wire sig000007b5;
  wire sig000007b6;
  wire sig000007b7;
  wire sig000007b8;
  wire sig000007b9;
  wire sig000007ba;
  wire sig000007bb;
  wire sig000007bc;
  wire sig000007bd;
  wire sig000007be;
  wire sig000007bf;
  wire sig000007c0;
  wire sig000007c1;
  wire sig000007c2;
  wire sig000007c3;
  wire sig000007c4;
  wire sig000007c5;
  wire sig000007c6;
  wire sig000007c7;
  wire sig000007c8;
  wire sig000007c9;
  wire sig000007ca;
  wire sig000007cb;
  wire sig000007cc;
  wire sig000007cd;
  wire sig000007ce;
  wire sig000007cf;
  wire sig000007d0;
  wire sig000007d1;
  wire sig000007d2;
  wire sig000007d3;
  wire sig000007d4;
  wire sig000007d5;
  wire sig000007d6;
  wire sig000007d7;
  wire sig000007d8;
  wire sig000007d9;
  wire sig000007da;
  wire sig000007db;
  wire sig000007dc;
  wire sig000007dd;
  wire sig000007de;
  wire sig000007df;
  wire sig000007e0;
  wire sig000007e1;
  wire sig000007e2;
  wire sig000007e3;
  wire sig000007e4;
  wire sig000007e5;
  wire sig000007e6;
  wire sig000007e7;
  wire sig000007e8;
  wire sig000007e9;
  wire sig000007ea;
  wire sig000007eb;
  wire sig000007ec;
  wire sig000007ed;
  wire sig000007ee;
  wire sig000007ef;
  wire sig000007f0;
  wire sig000007f1;
  wire sig000007f2;
  wire sig000007f3;
  wire sig000007f4;
  wire sig000007f5;
  wire sig000007f6;
  wire sig000007f7;
  wire sig000007f8;
  wire sig000007f9;
  wire sig000007fa;
  wire sig000007fb;
  wire sig000007fc;
  wire sig000007fd;
  wire sig000007fe;
  wire sig000007ff;
  wire sig00000800;
  wire sig00000801;
  wire sig00000802;
  wire sig00000803;
  wire sig00000804;
  wire sig00000805;
  wire sig00000806;
  wire sig00000807;
  wire sig00000808;
  wire sig00000809;
  wire sig0000080a;
  wire sig0000080b;
  wire sig0000080c;
  wire sig0000080d;
  wire sig0000080e;
  wire sig0000080f;
  wire sig00000810;
  wire sig00000811;
  wire sig00000812;
  wire sig00000813;
  wire sig00000814;
  wire sig00000815;
  wire sig00000816;
  wire sig00000817;
  wire sig00000818;
  wire sig00000819;
  wire sig0000081a;
  wire sig0000081b;
  wire sig0000081c;
  wire sig0000081d;
  wire sig0000081e;
  wire sig0000081f;
  wire sig00000820;
  wire sig00000821;
  wire sig00000822;
  wire sig00000823;
  wire sig00000824;
  wire sig00000825;
  wire sig00000826;
  wire sig00000827;
  wire sig00000828;
  wire sig00000829;
  wire sig0000082a;
  wire sig0000082b;
  wire sig0000082c;
  wire sig0000082d;
  wire sig0000082e;
  wire sig0000082f;
  wire sig00000830;
  wire sig00000831;
  wire sig00000832;
  wire sig00000833;
  wire sig00000834;
  wire sig00000835;
  wire sig00000836;
  wire sig00000837;
  wire sig00000838;
  wire sig00000839;
  wire sig0000083a;
  wire sig0000083b;
  wire sig0000083c;
  wire sig0000083d;
  wire sig0000083e;
  wire sig0000083f;
  wire sig00000840;
  wire sig00000841;
  wire sig00000842;
  wire sig00000843;
  wire sig00000844;
  wire sig00000845;
  wire NLW_blk000003c6_O_UNCONNECTED;
  wire NLW_blk000003cc_O_UNCONNECTED;
  wire NLW_blk00000416_O_UNCONNECTED;
  wire NLW_blk00000418_O_UNCONNECTED;
  wire NLW_blk0000041a_O_UNCONNECTED;
  wire NLW_blk0000041c_O_UNCONNECTED;
  wire NLW_blk0000041e_O_UNCONNECTED;
  wire NLW_blk00000420_O_UNCONNECTED;
  wire NLW_blk00000422_O_UNCONNECTED;
  wire NLW_blk00000424_O_UNCONNECTED;
  wire NLW_blk00000426_O_UNCONNECTED;
  wire NLW_blk00000428_O_UNCONNECTED;
  wire NLW_blk0000042a_O_UNCONNECTED;
  wire NLW_blk0000042c_O_UNCONNECTED;
  wire NLW_blk0000042d_O_UNCONNECTED;
  wire NLW_blk0000043b_O_UNCONNECTED;
  wire NLW_blk0000043f_O_UNCONNECTED;
  wire NLW_blk00000441_O_UNCONNECTED;
  wire NLW_blk00000443_O_UNCONNECTED;
  wire NLW_blk00000445_O_UNCONNECTED;
  wire NLW_blk00000447_O_UNCONNECTED;
  wire NLW_blk00000449_O_UNCONNECTED;
  wire NLW_blk0000044b_O_UNCONNECTED;
  wire NLW_blk0000044d_O_UNCONNECTED;
  wire NLW_blk0000044f_O_UNCONNECTED;
  wire NLW_blk00000451_O_UNCONNECTED;
  wire NLW_blk00000452_O_UNCONNECTED;
  wire NLW_blk000007d8_Q15_UNCONNECTED;
  wire NLW_blk000007da_Q15_UNCONNECTED;
  wire NLW_blk000007dc_Q15_UNCONNECTED;
  wire NLW_blk000007de_Q15_UNCONNECTED;
  wire NLW_blk000007e0_Q15_UNCONNECTED;
  wire NLW_blk000007e2_Q15_UNCONNECTED;
  wire NLW_blk000007e4_Q15_UNCONNECTED;
  wire NLW_blk000007e6_Q15_UNCONNECTED;
  wire NLW_blk000007e8_Q15_UNCONNECTED;
  wire NLW_blk000007ea_Q15_UNCONNECTED;
  wire NLW_blk000007ec_Q15_UNCONNECTED;
  wire NLW_blk000007ee_Q15_UNCONNECTED;
  wire NLW_blk000007f0_Q15_UNCONNECTED;
  wire NLW_blk000007f2_Q15_UNCONNECTED;
  wire NLW_blk000007f4_Q15_UNCONNECTED;
  wire NLW_blk000007f6_Q15_UNCONNECTED;
  wire NLW_blk000007f8_Q15_UNCONNECTED;
  wire NLW_blk000007fa_Q15_UNCONNECTED;
  wire NLW_blk000007fc_Q15_UNCONNECTED;
  wire NLW_blk000007fe_Q15_UNCONNECTED;
  wire NLW_blk00000800_Q15_UNCONNECTED;
  wire NLW_blk00000802_Q15_UNCONNECTED;
  wire NLW_blk00000804_Q15_UNCONNECTED;
  wire NLW_blk00000806_Q15_UNCONNECTED;
  wire NLW_blk00000808_Q15_UNCONNECTED;
  wire NLW_blk0000080a_Q15_UNCONNECTED;
  wire NLW_blk0000080c_Q15_UNCONNECTED;
  wire NLW_blk0000080e_Q15_UNCONNECTED;
  wire NLW_blk00000810_Q15_UNCONNECTED;
  wire NLW_blk00000812_PATTERNBDETECT_UNCONNECTED;
  wire NLW_blk00000812_MULTSIGNOUT_UNCONNECTED;
  wire NLW_blk00000812_CARRYCASCOUT_UNCONNECTED;
  wire NLW_blk00000812_UNDERFLOW_UNCONNECTED;
  wire NLW_blk00000812_PATTERNDETECT_UNCONNECTED;
  wire NLW_blk00000812_OVERFLOW_UNCONNECTED;
  wire \NLW_blk00000812_ACOUT<29>_UNCONNECTED ;
  wire \NLW_blk00000812_ACOUT<28>_UNCONNECTED ;
  wire \NLW_blk00000812_ACOUT<27>_UNCONNECTED ;
  wire \NLW_blk00000812_ACOUT<26>_UNCONNECTED ;
  wire \NLW_blk00000812_ACOUT<25>_UNCONNECTED ;
  wire \NLW_blk00000812_ACOUT<24>_UNCONNECTED ;
  wire \NLW_blk00000812_ACOUT<23>_UNCONNECTED ;
  wire \NLW_blk00000812_ACOUT<22>_UNCONNECTED ;
  wire \NLW_blk00000812_ACOUT<21>_UNCONNECTED ;
  wire \NLW_blk00000812_ACOUT<20>_UNCONNECTED ;
  wire \NLW_blk00000812_ACOUT<19>_UNCONNECTED ;
  wire \NLW_blk00000812_ACOUT<18>_UNCONNECTED ;
  wire \NLW_blk00000812_ACOUT<17>_UNCONNECTED ;
  wire \NLW_blk00000812_ACOUT<16>_UNCONNECTED ;
  wire \NLW_blk00000812_ACOUT<15>_UNCONNECTED ;
  wire \NLW_blk00000812_ACOUT<14>_UNCONNECTED ;
  wire \NLW_blk00000812_ACOUT<13>_UNCONNECTED ;
  wire \NLW_blk00000812_ACOUT<12>_UNCONNECTED ;
  wire \NLW_blk00000812_ACOUT<11>_UNCONNECTED ;
  wire \NLW_blk00000812_ACOUT<10>_UNCONNECTED ;
  wire \NLW_blk00000812_ACOUT<9>_UNCONNECTED ;
  wire \NLW_blk00000812_ACOUT<8>_UNCONNECTED ;
  wire \NLW_blk00000812_ACOUT<7>_UNCONNECTED ;
  wire \NLW_blk00000812_ACOUT<6>_UNCONNECTED ;
  wire \NLW_blk00000812_ACOUT<5>_UNCONNECTED ;
  wire \NLW_blk00000812_ACOUT<4>_UNCONNECTED ;
  wire \NLW_blk00000812_ACOUT<3>_UNCONNECTED ;
  wire \NLW_blk00000812_ACOUT<2>_UNCONNECTED ;
  wire \NLW_blk00000812_ACOUT<1>_UNCONNECTED ;
  wire \NLW_blk00000812_ACOUT<0>_UNCONNECTED ;
  wire \NLW_blk00000812_CARRYOUT<3>_UNCONNECTED ;
  wire \NLW_blk00000812_CARRYOUT<2>_UNCONNECTED ;
  wire \NLW_blk00000812_CARRYOUT<1>_UNCONNECTED ;
  wire \NLW_blk00000812_CARRYOUT<0>_UNCONNECTED ;
  wire \NLW_blk00000812_BCOUT<17>_UNCONNECTED ;
  wire \NLW_blk00000812_BCOUT<16>_UNCONNECTED ;
  wire \NLW_blk00000812_BCOUT<15>_UNCONNECTED ;
  wire \NLW_blk00000812_BCOUT<14>_UNCONNECTED ;
  wire \NLW_blk00000812_BCOUT<13>_UNCONNECTED ;
  wire \NLW_blk00000812_BCOUT<12>_UNCONNECTED ;
  wire \NLW_blk00000812_BCOUT<11>_UNCONNECTED ;
  wire \NLW_blk00000812_BCOUT<10>_UNCONNECTED ;
  wire \NLW_blk00000812_BCOUT<9>_UNCONNECTED ;
  wire \NLW_blk00000812_BCOUT<8>_UNCONNECTED ;
  wire \NLW_blk00000812_BCOUT<7>_UNCONNECTED ;
  wire \NLW_blk00000812_BCOUT<6>_UNCONNECTED ;
  wire \NLW_blk00000812_BCOUT<5>_UNCONNECTED ;
  wire \NLW_blk00000812_BCOUT<4>_UNCONNECTED ;
  wire \NLW_blk00000812_BCOUT<3>_UNCONNECTED ;
  wire \NLW_blk00000812_BCOUT<2>_UNCONNECTED ;
  wire \NLW_blk00000812_BCOUT<1>_UNCONNECTED ;
  wire \NLW_blk00000812_BCOUT<0>_UNCONNECTED ;
  wire \NLW_blk00000812_P<47>_UNCONNECTED ;
  wire \NLW_blk00000812_P<46>_UNCONNECTED ;
  wire \NLW_blk00000812_P<45>_UNCONNECTED ;
  wire \NLW_blk00000812_P<44>_UNCONNECTED ;
  wire \NLW_blk00000812_P<43>_UNCONNECTED ;
  wire \NLW_blk00000812_P<42>_UNCONNECTED ;
  wire \NLW_blk00000812_P<41>_UNCONNECTED ;
  wire \NLW_blk00000812_P<40>_UNCONNECTED ;
  wire \NLW_blk00000812_P<39>_UNCONNECTED ;
  wire \NLW_blk00000812_P<38>_UNCONNECTED ;
  wire \NLW_blk00000812_P<37>_UNCONNECTED ;
  wire \NLW_blk00000812_P<36>_UNCONNECTED ;
  wire \NLW_blk00000812_P<35>_UNCONNECTED ;
  wire \NLW_blk00000812_P<34>_UNCONNECTED ;
  wire \NLW_blk00000812_P<33>_UNCONNECTED ;
  wire \NLW_blk00000812_P<32>_UNCONNECTED ;
  wire \NLW_blk00000812_P<31>_UNCONNECTED ;
  wire \NLW_blk00000812_P<30>_UNCONNECTED ;
  wire \NLW_blk00000812_P<29>_UNCONNECTED ;
  wire \NLW_blk00000812_P<28>_UNCONNECTED ;
  wire \NLW_blk00000812_P<27>_UNCONNECTED ;
  wire \NLW_blk00000812_P<26>_UNCONNECTED ;
  wire \NLW_blk00000812_P<25>_UNCONNECTED ;
  wire \NLW_blk00000812_P<24>_UNCONNECTED ;
  wire \NLW_blk00000812_P<23>_UNCONNECTED ;
  wire \NLW_blk00000812_P<22>_UNCONNECTED ;
  wire \NLW_blk00000812_P<21>_UNCONNECTED ;
  wire \NLW_blk00000812_P<20>_UNCONNECTED ;
  wire \NLW_blk00000812_P<19>_UNCONNECTED ;
  wire \NLW_blk00000812_P<18>_UNCONNECTED ;
  wire \NLW_blk00000812_P<17>_UNCONNECTED ;
  wire \NLW_blk00000812_P<16>_UNCONNECTED ;
  wire \NLW_blk00000812_P<15>_UNCONNECTED ;
  wire \NLW_blk00000812_P<14>_UNCONNECTED ;
  wire \NLW_blk00000812_P<13>_UNCONNECTED ;
  wire \NLW_blk00000812_P<12>_UNCONNECTED ;
  wire \NLW_blk00000812_P<11>_UNCONNECTED ;
  wire \NLW_blk00000812_P<10>_UNCONNECTED ;
  wire \NLW_blk00000812_P<9>_UNCONNECTED ;
  wire \NLW_blk00000812_P<8>_UNCONNECTED ;
  wire \NLW_blk00000812_P<7>_UNCONNECTED ;
  wire \NLW_blk00000812_P<6>_UNCONNECTED ;
  wire \NLW_blk00000812_P<5>_UNCONNECTED ;
  wire \NLW_blk00000812_P<4>_UNCONNECTED ;
  wire \NLW_blk00000812_P<3>_UNCONNECTED ;
  wire \NLW_blk00000812_P<2>_UNCONNECTED ;
  wire \NLW_blk00000812_P<1>_UNCONNECTED ;
  wire \NLW_blk00000812_P<0>_UNCONNECTED ;
  wire NLW_blk00000813_PATTERNBDETECT_UNCONNECTED;
  wire NLW_blk00000813_MULTSIGNOUT_UNCONNECTED;
  wire NLW_blk00000813_CARRYCASCOUT_UNCONNECTED;
  wire NLW_blk00000813_UNDERFLOW_UNCONNECTED;
  wire NLW_blk00000813_PATTERNDETECT_UNCONNECTED;
  wire NLW_blk00000813_OVERFLOW_UNCONNECTED;
  wire \NLW_blk00000813_ACOUT<29>_UNCONNECTED ;
  wire \NLW_blk00000813_ACOUT<28>_UNCONNECTED ;
  wire \NLW_blk00000813_ACOUT<27>_UNCONNECTED ;
  wire \NLW_blk00000813_ACOUT<26>_UNCONNECTED ;
  wire \NLW_blk00000813_ACOUT<25>_UNCONNECTED ;
  wire \NLW_blk00000813_ACOUT<24>_UNCONNECTED ;
  wire \NLW_blk00000813_ACOUT<23>_UNCONNECTED ;
  wire \NLW_blk00000813_ACOUT<22>_UNCONNECTED ;
  wire \NLW_blk00000813_ACOUT<21>_UNCONNECTED ;
  wire \NLW_blk00000813_ACOUT<20>_UNCONNECTED ;
  wire \NLW_blk00000813_ACOUT<19>_UNCONNECTED ;
  wire \NLW_blk00000813_ACOUT<18>_UNCONNECTED ;
  wire \NLW_blk00000813_ACOUT<17>_UNCONNECTED ;
  wire \NLW_blk00000813_ACOUT<16>_UNCONNECTED ;
  wire \NLW_blk00000813_ACOUT<15>_UNCONNECTED ;
  wire \NLW_blk00000813_ACOUT<14>_UNCONNECTED ;
  wire \NLW_blk00000813_ACOUT<13>_UNCONNECTED ;
  wire \NLW_blk00000813_ACOUT<12>_UNCONNECTED ;
  wire \NLW_blk00000813_ACOUT<11>_UNCONNECTED ;
  wire \NLW_blk00000813_ACOUT<10>_UNCONNECTED ;
  wire \NLW_blk00000813_ACOUT<9>_UNCONNECTED ;
  wire \NLW_blk00000813_ACOUT<8>_UNCONNECTED ;
  wire \NLW_blk00000813_ACOUT<7>_UNCONNECTED ;
  wire \NLW_blk00000813_ACOUT<6>_UNCONNECTED ;
  wire \NLW_blk00000813_ACOUT<5>_UNCONNECTED ;
  wire \NLW_blk00000813_ACOUT<4>_UNCONNECTED ;
  wire \NLW_blk00000813_ACOUT<3>_UNCONNECTED ;
  wire \NLW_blk00000813_ACOUT<2>_UNCONNECTED ;
  wire \NLW_blk00000813_ACOUT<1>_UNCONNECTED ;
  wire \NLW_blk00000813_ACOUT<0>_UNCONNECTED ;
  wire \NLW_blk00000813_CARRYOUT<3>_UNCONNECTED ;
  wire \NLW_blk00000813_CARRYOUT<2>_UNCONNECTED ;
  wire \NLW_blk00000813_CARRYOUT<1>_UNCONNECTED ;
  wire \NLW_blk00000813_CARRYOUT<0>_UNCONNECTED ;
  wire \NLW_blk00000813_BCOUT<17>_UNCONNECTED ;
  wire \NLW_blk00000813_BCOUT<16>_UNCONNECTED ;
  wire \NLW_blk00000813_BCOUT<15>_UNCONNECTED ;
  wire \NLW_blk00000813_BCOUT<14>_UNCONNECTED ;
  wire \NLW_blk00000813_BCOUT<13>_UNCONNECTED ;
  wire \NLW_blk00000813_BCOUT<12>_UNCONNECTED ;
  wire \NLW_blk00000813_BCOUT<11>_UNCONNECTED ;
  wire \NLW_blk00000813_BCOUT<10>_UNCONNECTED ;
  wire \NLW_blk00000813_BCOUT<9>_UNCONNECTED ;
  wire \NLW_blk00000813_BCOUT<8>_UNCONNECTED ;
  wire \NLW_blk00000813_BCOUT<7>_UNCONNECTED ;
  wire \NLW_blk00000813_BCOUT<6>_UNCONNECTED ;
  wire \NLW_blk00000813_BCOUT<5>_UNCONNECTED ;
  wire \NLW_blk00000813_BCOUT<4>_UNCONNECTED ;
  wire \NLW_blk00000813_BCOUT<3>_UNCONNECTED ;
  wire \NLW_blk00000813_BCOUT<2>_UNCONNECTED ;
  wire \NLW_blk00000813_BCOUT<1>_UNCONNECTED ;
  wire \NLW_blk00000813_BCOUT<0>_UNCONNECTED ;
  wire \NLW_blk00000813_PCOUT<47>_UNCONNECTED ;
  wire \NLW_blk00000813_PCOUT<46>_UNCONNECTED ;
  wire \NLW_blk00000813_PCOUT<45>_UNCONNECTED ;
  wire \NLW_blk00000813_PCOUT<44>_UNCONNECTED ;
  wire \NLW_blk00000813_PCOUT<43>_UNCONNECTED ;
  wire \NLW_blk00000813_PCOUT<42>_UNCONNECTED ;
  wire \NLW_blk00000813_PCOUT<41>_UNCONNECTED ;
  wire \NLW_blk00000813_PCOUT<40>_UNCONNECTED ;
  wire \NLW_blk00000813_PCOUT<39>_UNCONNECTED ;
  wire \NLW_blk00000813_PCOUT<38>_UNCONNECTED ;
  wire \NLW_blk00000813_PCOUT<37>_UNCONNECTED ;
  wire \NLW_blk00000813_PCOUT<36>_UNCONNECTED ;
  wire \NLW_blk00000813_PCOUT<35>_UNCONNECTED ;
  wire \NLW_blk00000813_PCOUT<34>_UNCONNECTED ;
  wire \NLW_blk00000813_PCOUT<33>_UNCONNECTED ;
  wire \NLW_blk00000813_PCOUT<32>_UNCONNECTED ;
  wire \NLW_blk00000813_PCOUT<31>_UNCONNECTED ;
  wire \NLW_blk00000813_PCOUT<30>_UNCONNECTED ;
  wire \NLW_blk00000813_PCOUT<29>_UNCONNECTED ;
  wire \NLW_blk00000813_PCOUT<28>_UNCONNECTED ;
  wire \NLW_blk00000813_PCOUT<27>_UNCONNECTED ;
  wire \NLW_blk00000813_PCOUT<26>_UNCONNECTED ;
  wire \NLW_blk00000813_PCOUT<25>_UNCONNECTED ;
  wire \NLW_blk00000813_PCOUT<24>_UNCONNECTED ;
  wire \NLW_blk00000813_PCOUT<23>_UNCONNECTED ;
  wire \NLW_blk00000813_PCOUT<22>_UNCONNECTED ;
  wire \NLW_blk00000813_PCOUT<21>_UNCONNECTED ;
  wire \NLW_blk00000813_PCOUT<20>_UNCONNECTED ;
  wire \NLW_blk00000813_PCOUT<19>_UNCONNECTED ;
  wire \NLW_blk00000813_PCOUT<18>_UNCONNECTED ;
  wire \NLW_blk00000813_PCOUT<17>_UNCONNECTED ;
  wire \NLW_blk00000813_PCOUT<16>_UNCONNECTED ;
  wire \NLW_blk00000813_PCOUT<15>_UNCONNECTED ;
  wire \NLW_blk00000813_PCOUT<14>_UNCONNECTED ;
  wire \NLW_blk00000813_PCOUT<13>_UNCONNECTED ;
  wire \NLW_blk00000813_PCOUT<12>_UNCONNECTED ;
  wire \NLW_blk00000813_PCOUT<11>_UNCONNECTED ;
  wire \NLW_blk00000813_PCOUT<10>_UNCONNECTED ;
  wire \NLW_blk00000813_PCOUT<9>_UNCONNECTED ;
  wire \NLW_blk00000813_PCOUT<8>_UNCONNECTED ;
  wire \NLW_blk00000813_PCOUT<7>_UNCONNECTED ;
  wire \NLW_blk00000813_PCOUT<6>_UNCONNECTED ;
  wire \NLW_blk00000813_PCOUT<5>_UNCONNECTED ;
  wire \NLW_blk00000813_PCOUT<4>_UNCONNECTED ;
  wire \NLW_blk00000813_PCOUT<3>_UNCONNECTED ;
  wire \NLW_blk00000813_PCOUT<2>_UNCONNECTED ;
  wire \NLW_blk00000813_PCOUT<1>_UNCONNECTED ;
  wire \NLW_blk00000813_PCOUT<0>_UNCONNECTED ;
  wire NLW_blk00000814_PATTERNBDETECT_UNCONNECTED;
  wire NLW_blk00000814_MULTSIGNOUT_UNCONNECTED;
  wire NLW_blk00000814_CARRYCASCOUT_UNCONNECTED;
  wire NLW_blk00000814_UNDERFLOW_UNCONNECTED;
  wire NLW_blk00000814_PATTERNDETECT_UNCONNECTED;
  wire NLW_blk00000814_OVERFLOW_UNCONNECTED;
  wire \NLW_blk00000814_ACOUT<29>_UNCONNECTED ;
  wire \NLW_blk00000814_ACOUT<28>_UNCONNECTED ;
  wire \NLW_blk00000814_ACOUT<27>_UNCONNECTED ;
  wire \NLW_blk00000814_ACOUT<26>_UNCONNECTED ;
  wire \NLW_blk00000814_ACOUT<25>_UNCONNECTED ;
  wire \NLW_blk00000814_ACOUT<24>_UNCONNECTED ;
  wire \NLW_blk00000814_ACOUT<23>_UNCONNECTED ;
  wire \NLW_blk00000814_ACOUT<22>_UNCONNECTED ;
  wire \NLW_blk00000814_ACOUT<21>_UNCONNECTED ;
  wire \NLW_blk00000814_ACOUT<20>_UNCONNECTED ;
  wire \NLW_blk00000814_ACOUT<19>_UNCONNECTED ;
  wire \NLW_blk00000814_ACOUT<18>_UNCONNECTED ;
  wire \NLW_blk00000814_ACOUT<17>_UNCONNECTED ;
  wire \NLW_blk00000814_ACOUT<16>_UNCONNECTED ;
  wire \NLW_blk00000814_ACOUT<15>_UNCONNECTED ;
  wire \NLW_blk00000814_ACOUT<14>_UNCONNECTED ;
  wire \NLW_blk00000814_ACOUT<13>_UNCONNECTED ;
  wire \NLW_blk00000814_ACOUT<12>_UNCONNECTED ;
  wire \NLW_blk00000814_ACOUT<11>_UNCONNECTED ;
  wire \NLW_blk00000814_ACOUT<10>_UNCONNECTED ;
  wire \NLW_blk00000814_ACOUT<9>_UNCONNECTED ;
  wire \NLW_blk00000814_ACOUT<8>_UNCONNECTED ;
  wire \NLW_blk00000814_ACOUT<7>_UNCONNECTED ;
  wire \NLW_blk00000814_ACOUT<6>_UNCONNECTED ;
  wire \NLW_blk00000814_ACOUT<5>_UNCONNECTED ;
  wire \NLW_blk00000814_ACOUT<4>_UNCONNECTED ;
  wire \NLW_blk00000814_ACOUT<3>_UNCONNECTED ;
  wire \NLW_blk00000814_ACOUT<2>_UNCONNECTED ;
  wire \NLW_blk00000814_ACOUT<1>_UNCONNECTED ;
  wire \NLW_blk00000814_ACOUT<0>_UNCONNECTED ;
  wire \NLW_blk00000814_CARRYOUT<3>_UNCONNECTED ;
  wire \NLW_blk00000814_CARRYOUT<2>_UNCONNECTED ;
  wire \NLW_blk00000814_CARRYOUT<1>_UNCONNECTED ;
  wire \NLW_blk00000814_CARRYOUT<0>_UNCONNECTED ;
  wire \NLW_blk00000814_BCOUT<17>_UNCONNECTED ;
  wire \NLW_blk00000814_BCOUT<16>_UNCONNECTED ;
  wire \NLW_blk00000814_BCOUT<15>_UNCONNECTED ;
  wire \NLW_blk00000814_BCOUT<14>_UNCONNECTED ;
  wire \NLW_blk00000814_BCOUT<13>_UNCONNECTED ;
  wire \NLW_blk00000814_BCOUT<12>_UNCONNECTED ;
  wire \NLW_blk00000814_BCOUT<11>_UNCONNECTED ;
  wire \NLW_blk00000814_BCOUT<10>_UNCONNECTED ;
  wire \NLW_blk00000814_BCOUT<9>_UNCONNECTED ;
  wire \NLW_blk00000814_BCOUT<8>_UNCONNECTED ;
  wire \NLW_blk00000814_BCOUT<7>_UNCONNECTED ;
  wire \NLW_blk00000814_BCOUT<6>_UNCONNECTED ;
  wire \NLW_blk00000814_BCOUT<5>_UNCONNECTED ;
  wire \NLW_blk00000814_BCOUT<4>_UNCONNECTED ;
  wire \NLW_blk00000814_BCOUT<3>_UNCONNECTED ;
  wire \NLW_blk00000814_BCOUT<2>_UNCONNECTED ;
  wire \NLW_blk00000814_BCOUT<1>_UNCONNECTED ;
  wire \NLW_blk00000814_BCOUT<0>_UNCONNECTED ;
  wire \NLW_blk00000814_P<0>_UNCONNECTED ;
  wire \NLW_blk00000814_PCOUT<47>_UNCONNECTED ;
  wire \NLW_blk00000814_PCOUT<46>_UNCONNECTED ;
  wire \NLW_blk00000814_PCOUT<45>_UNCONNECTED ;
  wire \NLW_blk00000814_PCOUT<44>_UNCONNECTED ;
  wire \NLW_blk00000814_PCOUT<43>_UNCONNECTED ;
  wire \NLW_blk00000814_PCOUT<42>_UNCONNECTED ;
  wire \NLW_blk00000814_PCOUT<41>_UNCONNECTED ;
  wire \NLW_blk00000814_PCOUT<40>_UNCONNECTED ;
  wire \NLW_blk00000814_PCOUT<39>_UNCONNECTED ;
  wire \NLW_blk00000814_PCOUT<38>_UNCONNECTED ;
  wire \NLW_blk00000814_PCOUT<37>_UNCONNECTED ;
  wire \NLW_blk00000814_PCOUT<36>_UNCONNECTED ;
  wire \NLW_blk00000814_PCOUT<35>_UNCONNECTED ;
  wire \NLW_blk00000814_PCOUT<34>_UNCONNECTED ;
  wire \NLW_blk00000814_PCOUT<33>_UNCONNECTED ;
  wire \NLW_blk00000814_PCOUT<32>_UNCONNECTED ;
  wire \NLW_blk00000814_PCOUT<31>_UNCONNECTED ;
  wire \NLW_blk00000814_PCOUT<30>_UNCONNECTED ;
  wire \NLW_blk00000814_PCOUT<29>_UNCONNECTED ;
  wire \NLW_blk00000814_PCOUT<28>_UNCONNECTED ;
  wire \NLW_blk00000814_PCOUT<27>_UNCONNECTED ;
  wire \NLW_blk00000814_PCOUT<26>_UNCONNECTED ;
  wire \NLW_blk00000814_PCOUT<25>_UNCONNECTED ;
  wire \NLW_blk00000814_PCOUT<24>_UNCONNECTED ;
  wire \NLW_blk00000814_PCOUT<23>_UNCONNECTED ;
  wire \NLW_blk00000814_PCOUT<22>_UNCONNECTED ;
  wire \NLW_blk00000814_PCOUT<21>_UNCONNECTED ;
  wire \NLW_blk00000814_PCOUT<20>_UNCONNECTED ;
  wire \NLW_blk00000814_PCOUT<19>_UNCONNECTED ;
  wire \NLW_blk00000814_PCOUT<18>_UNCONNECTED ;
  wire \NLW_blk00000814_PCOUT<17>_UNCONNECTED ;
  wire \NLW_blk00000814_PCOUT<16>_UNCONNECTED ;
  wire \NLW_blk00000814_PCOUT<15>_UNCONNECTED ;
  wire \NLW_blk00000814_PCOUT<14>_UNCONNECTED ;
  wire \NLW_blk00000814_PCOUT<13>_UNCONNECTED ;
  wire \NLW_blk00000814_PCOUT<12>_UNCONNECTED ;
  wire \NLW_blk00000814_PCOUT<11>_UNCONNECTED ;
  wire \NLW_blk00000814_PCOUT<10>_UNCONNECTED ;
  wire \NLW_blk00000814_PCOUT<9>_UNCONNECTED ;
  wire \NLW_blk00000814_PCOUT<8>_UNCONNECTED ;
  wire \NLW_blk00000814_PCOUT<7>_UNCONNECTED ;
  wire \NLW_blk00000814_PCOUT<6>_UNCONNECTED ;
  wire \NLW_blk00000814_PCOUT<5>_UNCONNECTED ;
  wire \NLW_blk00000814_PCOUT<4>_UNCONNECTED ;
  wire \NLW_blk00000814_PCOUT<3>_UNCONNECTED ;
  wire \NLW_blk00000814_PCOUT<2>_UNCONNECTED ;
  wire \NLW_blk00000814_PCOUT<1>_UNCONNECTED ;
  wire \NLW_blk00000814_PCOUT<0>_UNCONNECTED ;
  wire [10 : 0] \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/exp_op ;
  wire [51 : 0] \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op ;
  assign
    result[63] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/sign_op ,
    result[62] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/exp_op [10],
    result[61] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/exp_op [9],
    result[60] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/exp_op [8],
    result[59] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/exp_op [7],
    result[58] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/exp_op [6],
    result[57] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/exp_op [5],
    result[56] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/exp_op [4],
    result[55] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/exp_op [3],
    result[54] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/exp_op [2],
    result[53] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/exp_op [1],
    result[52] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/exp_op [0],
    result[51] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [51],
    result[50] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [50],
    result[49] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [49],
    result[48] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [48],
    result[47] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [47],
    result[46] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [46],
    result[45] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [45],
    result[44] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [44],
    result[43] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [43],
    result[42] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [42],
    result[41] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [41],
    result[40] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [40],
    result[39] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [39],
    result[38] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [38],
    result[37] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [37],
    result[36] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [36],
    result[35] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [35],
    result[34] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [34],
    result[33] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [33],
    result[32] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [32],
    result[31] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [31],
    result[30] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [30],
    result[29] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [29],
    result[28] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [28],
    result[27] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [27],
    result[26] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [26],
    result[25] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [25],
    result[24] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [24],
    result[23] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [23],
    result[22] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [22],
    result[21] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [21],
    result[20] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [20],
    result[19] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [19],
    result[18] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [18],
    result[17] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [17],
    result[16] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [16],
    result[15] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [15],
    result[14] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [14],
    result[13] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [13],
    result[12] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [12],
    result[11] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [11],
    result[10] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [10],
    result[9] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [9],
    result[8] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [8],
    result[7] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [7],
    result[6] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [6],
    result[5] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [5],
    result[4] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [4],
    result[3] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [3],
    result[2] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [2],
    result[1] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [1],
    result[0] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [0];
  VCC   blk00000001 (
    .P(sig00000001)
  );
  GND   blk00000002 (
    .G(sig000006c3)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000003 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000156),
    .Q(sig0000023f)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000004 (
    .C(clk),
    .D(sig00000279),
    .Q(sig0000023b)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000005 (
    .C(clk),
    .D(sig00000278),
    .Q(sig0000023c)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000006 (
    .C(clk),
    .D(sig00000277),
    .Q(sig0000023e)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000007 (
    .C(clk),
    .D(sig000002b6),
    .Q(sig0000023a)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000008 (
    .C(clk),
    .D(sig000002b7),
    .Q(sig0000023d)
  );
  XORCY   blk00000009 (
    .CI(sig0000024b),
    .LI(sig00000001),
    .O(sig000002aa)
  );
  XORCY   blk0000000a (
    .CI(sig0000024d),
    .LI(sig0000024c),
    .O(sig000002b5)
  );
  MUXCY   blk0000000b (
    .CI(sig0000024d),
    .DI(sig000002d1),
    .S(sig0000024c),
    .O(sig0000024b)
  );
  XORCY   blk0000000c (
    .CI(sig0000024f),
    .LI(sig0000024e),
    .O(sig000002b4)
  );
  MUXCY   blk0000000d (
    .CI(sig0000024f),
    .DI(sig000002d0),
    .S(sig0000024e),
    .O(sig0000024d)
  );
  XORCY   blk0000000e (
    .CI(sig00000251),
    .LI(sig00000250),
    .O(sig000002b3)
  );
  MUXCY   blk0000000f (
    .CI(sig00000251),
    .DI(sig000002cf),
    .S(sig00000250),
    .O(sig0000024f)
  );
  XORCY   blk00000010 (
    .CI(sig00000253),
    .LI(sig00000252),
    .O(sig000002b2)
  );
  MUXCY   blk00000011 (
    .CI(sig00000253),
    .DI(sig000002ce),
    .S(sig00000252),
    .O(sig00000251)
  );
  XORCY   blk00000012 (
    .CI(sig00000255),
    .LI(sig00000254),
    .O(sig000002b1)
  );
  MUXCY   blk00000013 (
    .CI(sig00000255),
    .DI(sig000002cd),
    .S(sig00000254),
    .O(sig00000253)
  );
  XORCY   blk00000014 (
    .CI(sig00000257),
    .LI(sig00000256),
    .O(sig000002b0)
  );
  MUXCY   blk00000015 (
    .CI(sig00000257),
    .DI(sig000002cc),
    .S(sig00000256),
    .O(sig00000255)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000016 (
    .I0(sig000002cc),
    .I1(sig00000189),
    .O(sig00000256)
  );
  XORCY   blk00000017 (
    .CI(sig00000259),
    .LI(sig00000258),
    .O(sig000002af)
  );
  MUXCY   blk00000018 (
    .CI(sig00000259),
    .DI(sig000002cb),
    .S(sig00000258),
    .O(sig00000257)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000019 (
    .I0(sig000002cb),
    .I1(sig00000188),
    .O(sig00000258)
  );
  XORCY   blk0000001a (
    .CI(sig0000025b),
    .LI(sig0000025a),
    .O(sig000002ae)
  );
  MUXCY   blk0000001b (
    .CI(sig0000025b),
    .DI(sig000002ca),
    .S(sig0000025a),
    .O(sig00000259)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk0000001c (
    .I0(sig000002ca),
    .I1(sig00000187),
    .O(sig0000025a)
  );
  XORCY   blk0000001d (
    .CI(sig0000025d),
    .LI(sig0000025c),
    .O(sig000002ad)
  );
  MUXCY   blk0000001e (
    .CI(sig0000025d),
    .DI(sig000002c9),
    .S(sig0000025c),
    .O(sig0000025b)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk0000001f (
    .I0(sig000002c9),
    .I1(sig00000186),
    .O(sig0000025c)
  );
  XORCY   blk00000020 (
    .CI(sig0000025f),
    .LI(sig0000025e),
    .O(sig000002ac)
  );
  MUXCY   blk00000021 (
    .CI(sig0000025f),
    .DI(sig000002c8),
    .S(sig0000025e),
    .O(sig0000025d)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000022 (
    .I0(sig000002c8),
    .I1(sig0000011c),
    .O(sig0000025e)
  );
  XORCY   blk00000023 (
    .CI(sig00000001),
    .LI(sig00000260),
    .O(sig000002ab)
  );
  MUXCY   blk00000024 (
    .CI(sig00000001),
    .DI(sig000002c7),
    .S(sig00000260),
    .O(sig0000025f)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000025 (
    .I0(sig000002c7),
    .I1(sig0000011d),
    .O(sig00000260)
  );
  XORCY   blk00000026 (
    .CI(sig00000261),
    .LI(sig00000001),
    .O(sig0000029e)
  );
  XORCY   blk00000027 (
    .CI(sig00000263),
    .LI(sig00000262),
    .O(sig0000029d)
  );
  MUXCY   blk00000028 (
    .CI(sig00000263),
    .DI(b[62]),
    .S(sig00000262),
    .O(sig00000261)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000029 (
    .I0(b[62]),
    .I1(a[62]),
    .O(sig00000262)
  );
  XORCY   blk0000002a (
    .CI(sig00000265),
    .LI(sig00000264),
    .O(sig0000029c)
  );
  MUXCY   blk0000002b (
    .CI(sig00000265),
    .DI(b[61]),
    .S(sig00000264),
    .O(sig00000263)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk0000002c (
    .I0(b[61]),
    .I1(a[61]),
    .O(sig00000264)
  );
  XORCY   blk0000002d (
    .CI(sig00000267),
    .LI(sig00000266),
    .O(sig0000029b)
  );
  MUXCY   blk0000002e (
    .CI(sig00000267),
    .DI(b[60]),
    .S(sig00000266),
    .O(sig00000265)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk0000002f (
    .I0(b[60]),
    .I1(a[60]),
    .O(sig00000266)
  );
  XORCY   blk00000030 (
    .CI(sig00000269),
    .LI(sig00000268),
    .O(sig0000029a)
  );
  MUXCY   blk00000031 (
    .CI(sig00000269),
    .DI(b[59]),
    .S(sig00000268),
    .O(sig00000267)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000032 (
    .I0(b[59]),
    .I1(a[59]),
    .O(sig00000268)
  );
  XORCY   blk00000033 (
    .CI(sig0000026b),
    .LI(sig0000026a),
    .O(sig00000299)
  );
  MUXCY   blk00000034 (
    .CI(sig0000026b),
    .DI(b[58]),
    .S(sig0000026a),
    .O(sig00000269)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000035 (
    .I0(b[58]),
    .I1(a[58]),
    .O(sig0000026a)
  );
  XORCY   blk00000036 (
    .CI(sig0000026d),
    .LI(sig0000026c),
    .O(sig00000298)
  );
  MUXCY   blk00000037 (
    .CI(sig0000026d),
    .DI(b[57]),
    .S(sig0000026c),
    .O(sig0000026b)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000038 (
    .I0(b[57]),
    .I1(a[57]),
    .O(sig0000026c)
  );
  XORCY   blk00000039 (
    .CI(sig0000026f),
    .LI(sig0000026e),
    .O(sig00000297)
  );
  MUXCY   blk0000003a (
    .CI(sig0000026f),
    .DI(b[56]),
    .S(sig0000026e),
    .O(sig0000026d)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk0000003b (
    .I0(b[56]),
    .I1(a[56]),
    .O(sig0000026e)
  );
  XORCY   blk0000003c (
    .CI(sig00000271),
    .LI(sig00000270),
    .O(sig00000296)
  );
  MUXCY   blk0000003d (
    .CI(sig00000271),
    .DI(b[55]),
    .S(sig00000270),
    .O(sig0000026f)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk0000003e (
    .I0(b[55]),
    .I1(a[55]),
    .O(sig00000270)
  );
  XORCY   blk0000003f (
    .CI(sig00000273),
    .LI(sig00000272),
    .O(sig00000295)
  );
  MUXCY   blk00000040 (
    .CI(sig00000273),
    .DI(b[54]),
    .S(sig00000272),
    .O(sig00000271)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000041 (
    .I0(b[54]),
    .I1(a[54]),
    .O(sig00000272)
  );
  XORCY   blk00000042 (
    .CI(sig00000275),
    .LI(sig00000274),
    .O(sig00000294)
  );
  MUXCY   blk00000043 (
    .CI(sig00000275),
    .DI(b[53]),
    .S(sig00000274),
    .O(sig00000273)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000044 (
    .I0(b[53]),
    .I1(a[53]),
    .O(sig00000274)
  );
  MUXCY   blk00000045 (
    .CI(sig00000001),
    .DI(b[52]),
    .S(sig00000276),
    .O(sig00000275)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000046 (
    .I0(b[52]),
    .I1(a[52]),
    .O(sig00000276)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000047 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000002a1),
    .Q(sig000002b6)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000048 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000002a2),
    .Q(sig000002b7)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000049 (
    .C(clk),
    .CE(sig00000001),
    .D(a[63]),
    .Q(sig000002f5)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000004a (
    .C(clk),
    .CE(sig00000001),
    .D(sig000002a9),
    .Q(sig000002f4)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000004b (
    .C(clk),
    .CE(sig00000001),
    .D(sig000002aa),
    .Q(sig000002b8)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000004c (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000157),
    .Q(sig0000027d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000004d (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000027d),
    .Q(sig0000030c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000004e (
    .C(clk),
    .CE(sig00000001),
    .D(sig000002a0),
    .Q(sig0000027e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000004f (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000027e),
    .Q(sig0000022b)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000050 (
    .C(clk),
    .D(sig000001c2),
    .Q(sig0000027f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000051 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000022d),
    .Q(sig000002f3)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000052 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000291),
    .Q(sig000002f2)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000053 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000293),
    .Q(sig000002f1)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000054 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000292),
    .Q(sig000002ef)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000055 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000290),
    .Q(sig000004b6)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000056 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000002a6),
    .Q(sig000002ee)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000057 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000002a7),
    .Q(sig000002f0)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000058 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000002a8),
    .Q(sig000002ed)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000059 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000029f),
    .Q(sig000002c5)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000005a (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000030e),
    .Q(sig000002c4)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000005b (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000283),
    .Q(sig0000030f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000005c (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000282),
    .Q(sig00000310)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000005d (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000281),
    .Q(sig00000312)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000005e (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000280),
    .Q(sig00000313)
  );
  MUXCY   blk0000005f (
    .CI(sig00000328),
    .DI(sig000006c3),
    .S(sig00000326),
    .O(sig00000327)
  );
  MUXCY   blk00000060 (
    .CI(sig00000329),
    .DI(sig000006c3),
    .S(sig0000031e),
    .O(sig00000328)
  );
  MUXCY   blk00000061 (
    .CI(sig0000032a),
    .DI(sig000006c3),
    .S(sig0000031f),
    .O(sig00000329)
  );
  MUXCY   blk00000062 (
    .CI(sig0000032b),
    .DI(sig000006c3),
    .S(sig00000320),
    .O(sig0000032a)
  );
  MUXCY   blk00000063 (
    .CI(sig0000032c),
    .DI(sig000006c3),
    .S(sig00000321),
    .O(sig0000032b)
  );
  MUXCY   blk00000064 (
    .CI(sig0000032d),
    .DI(sig000006c3),
    .S(sig00000322),
    .O(sig0000032c)
  );
  MUXCY   blk00000065 (
    .CI(sig0000032e),
    .DI(sig000006c3),
    .S(sig00000323),
    .O(sig0000032d)
  );
  MUXCY   blk00000066 (
    .CI(sig0000032f),
    .DI(sig000006c3),
    .S(sig00000324),
    .O(sig0000032e)
  );
  MUXCY   blk00000067 (
    .CI(sig00000001),
    .DI(sig000006c3),
    .S(sig00000325),
    .O(sig0000032f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000068 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000327),
    .Q(sig00000311)
  );
  MUXCY   blk00000069 (
    .CI(sig00000331),
    .DI(sig000006c3),
    .S(sig0000031d),
    .O(sig00000330)
  );
  MUXCY   blk0000006a (
    .CI(sig00000332),
    .DI(sig000006c3),
    .S(sig00000315),
    .O(sig00000331)
  );
  MUXCY   blk0000006b (
    .CI(sig00000333),
    .DI(sig000006c3),
    .S(sig00000316),
    .O(sig00000332)
  );
  MUXCY   blk0000006c (
    .CI(sig00000334),
    .DI(sig000006c3),
    .S(sig00000317),
    .O(sig00000333)
  );
  MUXCY   blk0000006d (
    .CI(sig00000335),
    .DI(sig000006c3),
    .S(sig00000318),
    .O(sig00000334)
  );
  MUXCY   blk0000006e (
    .CI(sig00000336),
    .DI(sig000006c3),
    .S(sig00000319),
    .O(sig00000335)
  );
  MUXCY   blk0000006f (
    .CI(sig00000337),
    .DI(sig000006c3),
    .S(sig0000031a),
    .O(sig00000336)
  );
  MUXCY   blk00000070 (
    .CI(sig00000338),
    .DI(sig000006c3),
    .S(sig0000031b),
    .O(sig00000337)
  );
  MUXCY   blk00000071 (
    .CI(sig00000001),
    .DI(sig000006c3),
    .S(sig0000031c),
    .O(sig00000338)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000072 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000330),
    .Q(sig00000314)
  );
  MUXCY   blk00000073 (
    .CI(sig0000037a),
    .DI(sig00000359),
    .S(sig0000035a),
    .O(sig00000379)
  );
  MUXCY   blk00000074 (
    .CI(sig0000037b),
    .DI(sig0000035b),
    .S(sig0000035c),
    .O(sig0000037a)
  );
  MUXCY   blk00000075 (
    .CI(sig0000037c),
    .DI(sig0000035d),
    .S(sig0000035e),
    .O(sig0000037b)
  );
  MUXCY   blk00000076 (
    .CI(sig0000037d),
    .DI(sig0000035f),
    .S(sig00000360),
    .O(sig0000037c)
  );
  MUXCY   blk00000077 (
    .CI(sig0000037e),
    .DI(sig00000361),
    .S(sig00000362),
    .O(sig0000037d)
  );
  MUXCY   blk00000078 (
    .CI(sig0000037f),
    .DI(sig00000363),
    .S(sig00000364),
    .O(sig0000037e)
  );
  MUXCY   blk00000079 (
    .CI(sig00000380),
    .DI(sig00000365),
    .S(sig00000366),
    .O(sig0000037f)
  );
  MUXCY   blk0000007a (
    .CI(sig00000381),
    .DI(sig00000367),
    .S(sig00000368),
    .O(sig00000380)
  );
  MUXCY   blk0000007b (
    .CI(sig00000382),
    .DI(sig00000369),
    .S(sig0000036a),
    .O(sig00000381)
  );
  MUXCY   blk0000007c (
    .CI(sig00000383),
    .DI(sig0000036b),
    .S(sig0000036c),
    .O(sig00000382)
  );
  MUXCY   blk0000007d (
    .CI(sig00000384),
    .DI(sig0000036d),
    .S(sig0000036e),
    .O(sig00000383)
  );
  MUXCY   blk0000007e (
    .CI(sig00000385),
    .DI(sig0000036f),
    .S(sig00000370),
    .O(sig00000384)
  );
  MUXCY   blk0000007f (
    .CI(sig00000386),
    .DI(sig00000371),
    .S(sig00000372),
    .O(sig00000385)
  );
  MUXCY   blk00000080 (
    .CI(sig00000387),
    .DI(sig00000373),
    .S(sig00000374),
    .O(sig00000386)
  );
  MUXCY   blk00000081 (
    .CI(sig00000388),
    .DI(sig00000375),
    .S(sig00000376),
    .O(sig00000387)
  );
  MUXCY   blk00000082 (
    .CI(sig000006c3),
    .DI(sig00000377),
    .S(sig00000378),
    .O(sig00000388)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000083 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000379),
    .Q(sig0000027b)
  );
  MUXCY   blk00000084 (
    .CI(sig0000038a),
    .DI(sig00000339),
    .S(sig0000033a),
    .O(sig00000389)
  );
  MUXCY   blk00000085 (
    .CI(sig0000038b),
    .DI(sig0000033b),
    .S(sig0000033c),
    .O(sig0000038a)
  );
  MUXCY   blk00000086 (
    .CI(sig0000038c),
    .DI(sig0000033d),
    .S(sig0000033e),
    .O(sig0000038b)
  );
  MUXCY   blk00000087 (
    .CI(sig0000038d),
    .DI(sig0000033f),
    .S(sig00000340),
    .O(sig0000038c)
  );
  MUXCY   blk00000088 (
    .CI(sig0000038e),
    .DI(sig00000341),
    .S(sig00000342),
    .O(sig0000038d)
  );
  MUXCY   blk00000089 (
    .CI(sig0000038f),
    .DI(sig00000343),
    .S(sig00000344),
    .O(sig0000038e)
  );
  MUXCY   blk0000008a (
    .CI(sig00000390),
    .DI(sig00000345),
    .S(sig00000346),
    .O(sig0000038f)
  );
  MUXCY   blk0000008b (
    .CI(sig00000391),
    .DI(sig00000347),
    .S(sig00000348),
    .O(sig00000390)
  );
  MUXCY   blk0000008c (
    .CI(sig00000392),
    .DI(sig00000349),
    .S(sig0000034a),
    .O(sig00000391)
  );
  MUXCY   blk0000008d (
    .CI(sig00000393),
    .DI(sig0000034b),
    .S(sig0000034c),
    .O(sig00000392)
  );
  MUXCY   blk0000008e (
    .CI(sig00000394),
    .DI(sig0000034d),
    .S(sig0000034e),
    .O(sig00000393)
  );
  MUXCY   blk0000008f (
    .CI(sig00000395),
    .DI(sig0000034f),
    .S(sig00000350),
    .O(sig00000394)
  );
  MUXCY   blk00000090 (
    .CI(sig00000396),
    .DI(sig00000351),
    .S(sig00000352),
    .O(sig00000395)
  );
  MUXCY   blk00000091 (
    .CI(sig00000397),
    .DI(sig00000353),
    .S(sig00000354),
    .O(sig00000396)
  );
  MUXCY   blk00000092 (
    .CI(sig00000398),
    .DI(sig00000355),
    .S(sig00000356),
    .O(sig00000397)
  );
  MUXCY   blk00000093 (
    .CI(sig000006c3),
    .DI(sig00000357),
    .S(sig00000358),
    .O(sig00000398)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000094 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000389),
    .Q(sig0000027a)
  );
  MUXCY   blk00000095 (
    .CI(sig000003a5),
    .DI(sig000006c3),
    .S(sig00000399),
    .O(sig000003a4)
  );
  MUXCY   blk00000096 (
    .CI(sig000003a6),
    .DI(sig000006c3),
    .S(sig0000039a),
    .O(sig000003a5)
  );
  MUXCY   blk00000097 (
    .CI(sig000003a7),
    .DI(sig000006c3),
    .S(sig0000039b),
    .O(sig000003a6)
  );
  MUXCY   blk00000098 (
    .CI(sig000003a8),
    .DI(sig000006c3),
    .S(sig0000039c),
    .O(sig000003a7)
  );
  MUXCY   blk00000099 (
    .CI(sig000003a9),
    .DI(sig000006c3),
    .S(sig0000039d),
    .O(sig000003a8)
  );
  MUXCY   blk0000009a (
    .CI(sig000003aa),
    .DI(sig000006c3),
    .S(sig0000039e),
    .O(sig000003a9)
  );
  MUXCY   blk0000009b (
    .CI(sig000003ab),
    .DI(sig000006c3),
    .S(sig0000039f),
    .O(sig000003aa)
  );
  MUXCY   blk0000009c (
    .CI(sig000003ac),
    .DI(sig000006c3),
    .S(sig000003a0),
    .O(sig000003ab)
  );
  MUXCY   blk0000009d (
    .CI(sig000003ad),
    .DI(sig000006c3),
    .S(sig000003a1),
    .O(sig000003ac)
  );
  MUXCY   blk0000009e (
    .CI(sig000003ae),
    .DI(sig000006c3),
    .S(sig000003a2),
    .O(sig000003ad)
  );
  MUXCY   blk0000009f (
    .CI(sig00000001),
    .DI(sig000006c3),
    .S(sig000003a3),
    .O(sig000003ae)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000a0 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000003a4),
    .Q(sig0000027c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000a1 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000002b5),
    .Q(sig000002c3)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000a2 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000002b4),
    .Q(sig000002c2)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000a3 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000002b3),
    .Q(sig000002c1)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000a4 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000002b2),
    .Q(sig000002c0)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000a5 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000002b1),
    .Q(sig000002bf)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000a6 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000002b0),
    .Q(sig000002be)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000a7 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000002af),
    .Q(sig000002bd)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000a8 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000002ae),
    .Q(sig000002bc)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000a9 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000002ad),
    .Q(sig000002bb)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000aa (
    .C(clk),
    .CE(sig00000001),
    .D(sig000002ac),
    .Q(sig000002ba)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000ab (
    .C(clk),
    .CE(sig00000001),
    .D(sig000002ab),
    .Q(sig000002b9)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000ac (
    .C(clk),
    .CE(sig00000001),
    .D(b[62]),
    .Q(sig00000300)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000ad (
    .C(clk),
    .CE(sig00000001),
    .D(b[61]),
    .Q(sig000002ff)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000ae (
    .C(clk),
    .CE(sig00000001),
    .D(b[60]),
    .Q(sig000002fe)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000af (
    .C(clk),
    .CE(sig00000001),
    .D(b[59]),
    .Q(sig000002fd)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000b0 (
    .C(clk),
    .CE(sig00000001),
    .D(b[58]),
    .Q(sig000002fc)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000b1 (
    .C(clk),
    .CE(sig00000001),
    .D(b[57]),
    .Q(sig000002fb)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000b2 (
    .C(clk),
    .CE(sig00000001),
    .D(b[56]),
    .Q(sig000002fa)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000b3 (
    .C(clk),
    .CE(sig00000001),
    .D(b[55]),
    .Q(sig000002f9)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000b4 (
    .C(clk),
    .CE(sig00000001),
    .D(b[54]),
    .Q(sig000002f8)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000b5 (
    .C(clk),
    .CE(sig00000001),
    .D(b[53]),
    .Q(sig000002f7)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000b6 (
    .C(clk),
    .CE(sig00000001),
    .D(b[52]),
    .Q(sig000002f6)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000b7 (
    .C(clk),
    .CE(sig00000001),
    .D(a[62]),
    .Q(sig0000030b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000b8 (
    .C(clk),
    .CE(sig00000001),
    .D(a[61]),
    .Q(sig0000030a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000b9 (
    .C(clk),
    .CE(sig00000001),
    .D(a[60]),
    .Q(sig00000309)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000ba (
    .C(clk),
    .CE(sig00000001),
    .D(a[59]),
    .Q(sig00000308)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000bb (
    .C(clk),
    .CE(sig00000001),
    .D(a[58]),
    .Q(sig00000307)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000bc (
    .C(clk),
    .CE(sig00000001),
    .D(a[57]),
    .Q(sig00000306)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000bd (
    .C(clk),
    .CE(sig00000001),
    .D(a[56]),
    .Q(sig00000305)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000be (
    .C(clk),
    .CE(sig00000001),
    .D(a[55]),
    .Q(sig00000304)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000bf (
    .C(clk),
    .CE(sig00000001),
    .D(a[54]),
    .Q(sig00000303)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000c0 (
    .C(clk),
    .CE(sig00000001),
    .D(a[53]),
    .Q(sig00000302)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000c1 (
    .C(clk),
    .CE(sig00000001),
    .D(a[52]),
    .Q(sig00000301)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000000c2 (
    .C(clk),
    .D(sig0000029e),
    .Q(sig0000024a)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000000c3 (
    .C(clk),
    .D(sig0000029d),
    .Q(sig00000249)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000000c4 (
    .C(clk),
    .D(sig0000029c),
    .Q(sig00000248)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000000c5 (
    .C(clk),
    .D(sig0000029b),
    .Q(sig00000247)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000000c6 (
    .C(clk),
    .D(sig0000029a),
    .Q(sig00000246)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000000c7 (
    .C(clk),
    .D(sig00000299),
    .Q(sig00000245)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000000c8 (
    .C(clk),
    .D(sig00000298),
    .Q(sig00000244)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000000c9 (
    .C(clk),
    .D(sig00000297),
    .Q(sig00000243)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000000ca (
    .C(clk),
    .D(sig00000296),
    .Q(sig00000242)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000000cb (
    .C(clk),
    .D(sig00000295),
    .Q(sig00000241)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000000cc (
    .C(clk),
    .D(sig00000294),
    .Q(sig00000240)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000000cd (
    .C(clk),
    .D(sig000002a5),
    .Q(sig000003b0)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000000ce (
    .C(clk),
    .D(sig000002a4),
    .Q(sig000003af)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000000cf (
    .C(clk),
    .D(sig000002a3),
    .Q(sig000003b1)
  );
  XORCY   blk000000d0 (
    .CI(sig000003b2),
    .LI(sig000006c3),
    .O(sig000002e9)
  );
  XORCY   blk000000d1 (
    .CI(sig000003b3),
    .LI(sig0000028e),
    .O(sig000002e8)
  );
  MUXCY   blk000000d2 (
    .CI(sig000003b3),
    .DI(sig000006c3),
    .S(sig0000028e),
    .O(sig000003b2)
  );
  XORCY   blk000000d3 (
    .CI(sig000003b4),
    .LI(sig0000028d),
    .O(sig000002e7)
  );
  MUXCY   blk000000d4 (
    .CI(sig000003b4),
    .DI(sig000006c3),
    .S(sig0000028d),
    .O(sig000003b3)
  );
  XORCY   blk000000d5 (
    .CI(sig000003b5),
    .LI(sig0000028c),
    .O(sig000002e6)
  );
  MUXCY   blk000000d6 (
    .CI(sig000003b5),
    .DI(sig000006c3),
    .S(sig0000028c),
    .O(sig000003b4)
  );
  XORCY   blk000000d7 (
    .CI(sig000003b6),
    .LI(sig0000028b),
    .O(sig000002e5)
  );
  MUXCY   blk000000d8 (
    .CI(sig000003b6),
    .DI(sig000006c3),
    .S(sig0000028b),
    .O(sig000003b5)
  );
  XORCY   blk000000d9 (
    .CI(sig000003b7),
    .LI(sig0000028a),
    .O(sig000002e4)
  );
  MUXCY   blk000000da (
    .CI(sig000003b7),
    .DI(sig000006c3),
    .S(sig0000028a),
    .O(sig000003b6)
  );
  XORCY   blk000000db (
    .CI(sig000003b8),
    .LI(sig00000289),
    .O(sig000002e3)
  );
  MUXCY   blk000000dc (
    .CI(sig000003b8),
    .DI(sig000006c3),
    .S(sig00000289),
    .O(sig000003b7)
  );
  XORCY   blk000000dd (
    .CI(sig000003b9),
    .LI(sig00000288),
    .O(sig000002e2)
  );
  MUXCY   blk000000de (
    .CI(sig000003b9),
    .DI(sig000006c3),
    .S(sig00000288),
    .O(sig000003b8)
  );
  XORCY   blk000000df (
    .CI(sig000003ba),
    .LI(sig00000287),
    .O(sig000002e1)
  );
  MUXCY   blk000000e0 (
    .CI(sig000003ba),
    .DI(sig000006c3),
    .S(sig00000287),
    .O(sig000003b9)
  );
  XORCY   blk000000e1 (
    .CI(sig000003bb),
    .LI(sig00000286),
    .O(sig000002e0)
  );
  MUXCY   blk000000e2 (
    .CI(sig000003bb),
    .DI(sig000006c3),
    .S(sig00000286),
    .O(sig000003ba)
  );
  XORCY   blk000000e3 (
    .CI(sig000003bc),
    .LI(sig00000285),
    .O(sig000002df)
  );
  MUXCY   blk000000e4 (
    .CI(sig000003bc),
    .DI(sig000006c3),
    .S(sig00000285),
    .O(sig000003bb)
  );
  XORCY   blk000000e5 (
    .CI(sig000006c3),
    .LI(sig00000284),
    .O(sig000002de)
  );
  MUXCY   blk000000e6 (
    .CI(sig000006c3),
    .DI(sig00000001),
    .S(sig00000284),
    .O(sig000003bc)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000000e7 (
    .C(clk),
    .D(sig000002e9),
    .Q(sig000002dd)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000000e8 (
    .C(clk),
    .D(sig000002e8),
    .Q(sig000002dc)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000000e9 (
    .C(clk),
    .D(sig000002e7),
    .Q(sig000002db)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000000ea (
    .C(clk),
    .D(sig000002e6),
    .Q(sig000002da)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000000eb (
    .C(clk),
    .D(sig000002e5),
    .Q(sig000002d9)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000000ec (
    .C(clk),
    .D(sig000002e4),
    .Q(sig000002d8)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000000ed (
    .C(clk),
    .D(sig000002e3),
    .Q(sig000002d7)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000000ee (
    .C(clk),
    .D(sig000002e2),
    .Q(sig000002d6)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000000ef (
    .C(clk),
    .D(sig000002e1),
    .Q(sig000002d5)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000000f0 (
    .C(clk),
    .D(sig000002e0),
    .Q(sig000002d4)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000000f1 (
    .C(clk),
    .D(sig000002df),
    .Q(sig000002d3)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000000f2 (
    .C(clk),
    .D(sig000002de),
    .Q(sig000002d2)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000000f3 (
    .C(clk),
    .D(sig0000028f),
    .Q(sig000003bd)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000000f4 (
    .C(clk),
    .D(sig000003c8),
    .Q(sig00000239)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000000f5 (
    .C(clk),
    .D(sig000003c7),
    .Q(sig00000238)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000000f6 (
    .C(clk),
    .D(sig000003c6),
    .Q(sig00000237)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000000f7 (
    .C(clk),
    .D(sig000003c5),
    .Q(sig00000236)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000000f8 (
    .C(clk),
    .D(sig000003c4),
    .Q(sig00000235)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000000f9 (
    .C(clk),
    .D(sig000003c3),
    .Q(sig00000234)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000000fa (
    .C(clk),
    .D(sig000003c2),
    .Q(sig00000233)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000000fb (
    .C(clk),
    .D(sig000003c1),
    .Q(sig00000232)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000000fc (
    .C(clk),
    .D(sig000003c0),
    .Q(sig00000231)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000000fd (
    .C(clk),
    .D(sig000003bf),
    .Q(sig00000230)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000000fe (
    .C(clk),
    .D(sig000003be),
    .Q(sig0000022f)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000000ff (
    .C(clk),
    .D(sig000002c3),
    .Q(sig000003c8)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000100 (
    .C(clk),
    .D(sig000002c2),
    .Q(sig000003c7)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000101 (
    .C(clk),
    .D(sig000002c1),
    .Q(sig000003c6)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000102 (
    .C(clk),
    .D(sig000002c0),
    .Q(sig000003c5)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000103 (
    .C(clk),
    .D(sig000002bf),
    .Q(sig000003c4)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000104 (
    .C(clk),
    .D(sig000002be),
    .Q(sig000003c3)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000105 (
    .C(clk),
    .D(sig000002bd),
    .Q(sig000003c2)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000106 (
    .C(clk),
    .D(sig000002bc),
    .Q(sig000003c1)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000107 (
    .C(clk),
    .D(sig000002bb),
    .Q(sig000003c0)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000108 (
    .C(clk),
    .D(sig000002ba),
    .Q(sig000003bf)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000109 (
    .C(clk),
    .D(sig000002b9),
    .Q(sig000003be)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000010a (
    .C(clk),
    .CE(sig00000001),
    .D(b[51]),
    .Q(sig000001f6)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000010b (
    .C(clk),
    .CE(sig00000001),
    .D(b[50]),
    .Q(sig000001f5)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000010c (
    .C(clk),
    .CE(sig00000001),
    .D(b[49]),
    .Q(sig000001f4)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000010d (
    .C(clk),
    .CE(sig00000001),
    .D(b[48]),
    .Q(sig000001f3)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000010e (
    .C(clk),
    .CE(sig00000001),
    .D(b[47]),
    .Q(sig000001f2)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000010f (
    .C(clk),
    .CE(sig00000001),
    .D(b[46]),
    .Q(sig000001f1)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000110 (
    .C(clk),
    .CE(sig00000001),
    .D(b[45]),
    .Q(sig000001f0)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000111 (
    .C(clk),
    .CE(sig00000001),
    .D(b[44]),
    .Q(sig000001ef)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000112 (
    .C(clk),
    .CE(sig00000001),
    .D(b[43]),
    .Q(sig000001ee)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000113 (
    .C(clk),
    .CE(sig00000001),
    .D(b[42]),
    .Q(sig000001ed)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000114 (
    .C(clk),
    .CE(sig00000001),
    .D(b[41]),
    .Q(sig000001ec)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000115 (
    .C(clk),
    .CE(sig00000001),
    .D(b[40]),
    .Q(sig000001eb)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000116 (
    .C(clk),
    .CE(sig00000001),
    .D(b[39]),
    .Q(sig000001ea)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000117 (
    .C(clk),
    .CE(sig00000001),
    .D(b[38]),
    .Q(sig000001e9)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000118 (
    .C(clk),
    .CE(sig00000001),
    .D(b[37]),
    .Q(sig000001e8)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000119 (
    .C(clk),
    .CE(sig00000001),
    .D(b[36]),
    .Q(sig000001e7)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000011a (
    .C(clk),
    .CE(sig00000001),
    .D(b[35]),
    .Q(sig000001e6)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000011b (
    .C(clk),
    .CE(sig00000001),
    .D(b[34]),
    .Q(sig000001e5)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000011c (
    .C(clk),
    .CE(sig00000001),
    .D(b[33]),
    .Q(sig000001e4)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000011d (
    .C(clk),
    .CE(sig00000001),
    .D(b[32]),
    .Q(sig000001e3)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000011e (
    .C(clk),
    .CE(sig00000001),
    .D(b[31]),
    .Q(sig000001e2)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000011f (
    .C(clk),
    .CE(sig00000001),
    .D(b[30]),
    .Q(sig000001e1)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000120 (
    .C(clk),
    .CE(sig00000001),
    .D(b[29]),
    .Q(sig000001e0)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000121 (
    .C(clk),
    .CE(sig00000001),
    .D(b[28]),
    .Q(sig000001df)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000122 (
    .C(clk),
    .CE(sig00000001),
    .D(b[27]),
    .Q(sig000001de)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000123 (
    .C(clk),
    .CE(sig00000001),
    .D(b[26]),
    .Q(sig000001dd)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000124 (
    .C(clk),
    .CE(sig00000001),
    .D(b[25]),
    .Q(sig000001dc)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000125 (
    .C(clk),
    .CE(sig00000001),
    .D(b[24]),
    .Q(sig000001db)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000126 (
    .C(clk),
    .CE(sig00000001),
    .D(b[23]),
    .Q(sig000001da)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000127 (
    .C(clk),
    .CE(sig00000001),
    .D(b[22]),
    .Q(sig000001d9)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000128 (
    .C(clk),
    .CE(sig00000001),
    .D(b[21]),
    .Q(sig000001d8)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000129 (
    .C(clk),
    .CE(sig00000001),
    .D(b[20]),
    .Q(sig000001d7)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000012a (
    .C(clk),
    .CE(sig00000001),
    .D(b[19]),
    .Q(sig000001d6)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000012b (
    .C(clk),
    .CE(sig00000001),
    .D(b[18]),
    .Q(sig000001d5)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000012c (
    .C(clk),
    .CE(sig00000001),
    .D(b[17]),
    .Q(sig000001d4)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000012d (
    .C(clk),
    .CE(sig00000001),
    .D(b[16]),
    .Q(sig000001d3)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000012e (
    .C(clk),
    .CE(sig00000001),
    .D(b[15]),
    .Q(sig000001d2)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000012f (
    .C(clk),
    .CE(sig00000001),
    .D(b[14]),
    .Q(sig000001d1)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000130 (
    .C(clk),
    .CE(sig00000001),
    .D(b[13]),
    .Q(sig000001d0)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000131 (
    .C(clk),
    .CE(sig00000001),
    .D(b[12]),
    .Q(sig000001cf)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000132 (
    .C(clk),
    .CE(sig00000001),
    .D(b[11]),
    .Q(sig000001ce)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000133 (
    .C(clk),
    .CE(sig00000001),
    .D(b[10]),
    .Q(sig000001cd)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000134 (
    .C(clk),
    .CE(sig00000001),
    .D(b[9]),
    .Q(sig000001cc)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000135 (
    .C(clk),
    .CE(sig00000001),
    .D(b[8]),
    .Q(sig000001cb)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000136 (
    .C(clk),
    .CE(sig00000001),
    .D(b[7]),
    .Q(sig000001ca)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000137 (
    .C(clk),
    .CE(sig00000001),
    .D(b[6]),
    .Q(sig000001c9)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000138 (
    .C(clk),
    .CE(sig00000001),
    .D(b[5]),
    .Q(sig000001c8)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000139 (
    .C(clk),
    .CE(sig00000001),
    .D(b[4]),
    .Q(sig000001c7)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000013a (
    .C(clk),
    .CE(sig00000001),
    .D(b[3]),
    .Q(sig000001c6)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000013b (
    .C(clk),
    .CE(sig00000001),
    .D(b[2]),
    .Q(sig000001c5)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000013c (
    .C(clk),
    .CE(sig00000001),
    .D(b[1]),
    .Q(sig000001c4)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000013d (
    .C(clk),
    .CE(sig00000001),
    .D(b[0]),
    .Q(sig000001c3)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000013e (
    .C(clk),
    .CE(sig00000001),
    .D(a[51]),
    .Q(sig0000022a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000013f (
    .C(clk),
    .CE(sig00000001),
    .D(a[50]),
    .Q(sig00000229)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000140 (
    .C(clk),
    .CE(sig00000001),
    .D(a[49]),
    .Q(sig00000228)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000141 (
    .C(clk),
    .CE(sig00000001),
    .D(a[48]),
    .Q(sig00000227)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000142 (
    .C(clk),
    .CE(sig00000001),
    .D(a[47]),
    .Q(sig00000226)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000143 (
    .C(clk),
    .CE(sig00000001),
    .D(a[46]),
    .Q(sig00000225)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000144 (
    .C(clk),
    .CE(sig00000001),
    .D(a[45]),
    .Q(sig00000224)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000145 (
    .C(clk),
    .CE(sig00000001),
    .D(a[44]),
    .Q(sig00000223)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000146 (
    .C(clk),
    .CE(sig00000001),
    .D(a[43]),
    .Q(sig00000222)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000147 (
    .C(clk),
    .CE(sig00000001),
    .D(a[42]),
    .Q(sig00000221)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000148 (
    .C(clk),
    .CE(sig00000001),
    .D(a[41]),
    .Q(sig00000220)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000149 (
    .C(clk),
    .CE(sig00000001),
    .D(a[40]),
    .Q(sig0000021f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000014a (
    .C(clk),
    .CE(sig00000001),
    .D(a[39]),
    .Q(sig0000021e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000014b (
    .C(clk),
    .CE(sig00000001),
    .D(a[38]),
    .Q(sig0000021d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000014c (
    .C(clk),
    .CE(sig00000001),
    .D(a[37]),
    .Q(sig0000021c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000014d (
    .C(clk),
    .CE(sig00000001),
    .D(a[36]),
    .Q(sig0000021b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000014e (
    .C(clk),
    .CE(sig00000001),
    .D(a[35]),
    .Q(sig0000021a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000014f (
    .C(clk),
    .CE(sig00000001),
    .D(a[34]),
    .Q(sig00000219)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000150 (
    .C(clk),
    .CE(sig00000001),
    .D(a[33]),
    .Q(sig00000218)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000151 (
    .C(clk),
    .CE(sig00000001),
    .D(a[32]),
    .Q(sig00000217)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000152 (
    .C(clk),
    .CE(sig00000001),
    .D(a[31]),
    .Q(sig00000216)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000153 (
    .C(clk),
    .CE(sig00000001),
    .D(a[30]),
    .Q(sig00000215)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000154 (
    .C(clk),
    .CE(sig00000001),
    .D(a[29]),
    .Q(sig00000214)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000155 (
    .C(clk),
    .CE(sig00000001),
    .D(a[28]),
    .Q(sig00000213)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000156 (
    .C(clk),
    .CE(sig00000001),
    .D(a[27]),
    .Q(sig00000212)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000157 (
    .C(clk),
    .CE(sig00000001),
    .D(a[26]),
    .Q(sig00000211)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000158 (
    .C(clk),
    .CE(sig00000001),
    .D(a[25]),
    .Q(sig00000210)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000159 (
    .C(clk),
    .CE(sig00000001),
    .D(a[24]),
    .Q(sig0000020f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000015a (
    .C(clk),
    .CE(sig00000001),
    .D(a[23]),
    .Q(sig0000020e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000015b (
    .C(clk),
    .CE(sig00000001),
    .D(a[22]),
    .Q(sig0000020d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000015c (
    .C(clk),
    .CE(sig00000001),
    .D(a[21]),
    .Q(sig0000020c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000015d (
    .C(clk),
    .CE(sig00000001),
    .D(a[20]),
    .Q(sig0000020b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000015e (
    .C(clk),
    .CE(sig00000001),
    .D(a[19]),
    .Q(sig0000020a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000015f (
    .C(clk),
    .CE(sig00000001),
    .D(a[18]),
    .Q(sig00000209)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000160 (
    .C(clk),
    .CE(sig00000001),
    .D(a[17]),
    .Q(sig00000208)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000161 (
    .C(clk),
    .CE(sig00000001),
    .D(a[16]),
    .Q(sig00000207)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000162 (
    .C(clk),
    .CE(sig00000001),
    .D(a[15]),
    .Q(sig00000206)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000163 (
    .C(clk),
    .CE(sig00000001),
    .D(a[14]),
    .Q(sig00000205)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000164 (
    .C(clk),
    .CE(sig00000001),
    .D(a[13]),
    .Q(sig00000204)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000165 (
    .C(clk),
    .CE(sig00000001),
    .D(a[12]),
    .Q(sig00000203)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000166 (
    .C(clk),
    .CE(sig00000001),
    .D(a[11]),
    .Q(sig00000202)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000167 (
    .C(clk),
    .CE(sig00000001),
    .D(a[10]),
    .Q(sig00000201)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000168 (
    .C(clk),
    .CE(sig00000001),
    .D(a[9]),
    .Q(sig00000200)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000169 (
    .C(clk),
    .CE(sig00000001),
    .D(a[8]),
    .Q(sig000001ff)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000016a (
    .C(clk),
    .CE(sig00000001),
    .D(a[7]),
    .Q(sig000001fe)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000016b (
    .C(clk),
    .CE(sig00000001),
    .D(a[6]),
    .Q(sig000001fd)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000016c (
    .C(clk),
    .CE(sig00000001),
    .D(a[5]),
    .Q(sig000001fc)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000016d (
    .C(clk),
    .CE(sig00000001),
    .D(a[4]),
    .Q(sig000001fb)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000016e (
    .C(clk),
    .CE(sig00000001),
    .D(a[3]),
    .Q(sig000001fa)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000016f (
    .C(clk),
    .CE(sig00000001),
    .D(a[2]),
    .Q(sig000001f9)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000170 (
    .C(clk),
    .CE(sig00000001),
    .D(a[1]),
    .Q(sig000001f8)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000171 (
    .C(clk),
    .CE(sig00000001),
    .D(a[0]),
    .Q(sig000001f7)
  );
  XORCY   blk00000172 (
    .CI(sig000003c9),
    .LI(sig00000583),
    .O(sig000004c6)
  );
  XORCY   blk00000173 (
    .CI(sig000003ca),
    .LI(sig00000582),
    .O(sig000004c5)
  );
  MUXCY   blk00000174 (
    .CI(sig000003ca),
    .DI(sig000006c3),
    .S(sig00000582),
    .O(sig000003c9)
  );
  XORCY   blk00000175 (
    .CI(sig000003cb),
    .LI(sig00000581),
    .O(sig000004c4)
  );
  MUXCY   blk00000176 (
    .CI(sig000003cb),
    .DI(sig000006c3),
    .S(sig00000581),
    .O(sig000003ca)
  );
  XORCY   blk00000177 (
    .CI(sig000003cc),
    .LI(sig00000580),
    .O(sig000004c3)
  );
  MUXCY   blk00000178 (
    .CI(sig000003cc),
    .DI(sig000006c3),
    .S(sig00000580),
    .O(sig000003cb)
  );
  XORCY   blk00000179 (
    .CI(sig000003cd),
    .LI(sig0000057f),
    .O(sig000004c2)
  );
  MUXCY   blk0000017a (
    .CI(sig000003cd),
    .DI(sig000006c3),
    .S(sig0000057f),
    .O(sig000003cc)
  );
  XORCY   blk0000017b (
    .CI(sig000003ce),
    .LI(sig0000057e),
    .O(sig000004c1)
  );
  MUXCY   blk0000017c (
    .CI(sig000003ce),
    .DI(sig000006c3),
    .S(sig0000057e),
    .O(sig000003cd)
  );
  XORCY   blk0000017d (
    .CI(sig000003cf),
    .LI(sig0000057d),
    .O(sig000004c0)
  );
  MUXCY   blk0000017e (
    .CI(sig000003cf),
    .DI(sig000006c3),
    .S(sig0000057d),
    .O(sig000003ce)
  );
  XORCY   blk0000017f (
    .CI(sig000003d0),
    .LI(sig0000057c),
    .O(sig000004bf)
  );
  MUXCY   blk00000180 (
    .CI(sig000003d0),
    .DI(sig000006c3),
    .S(sig0000057c),
    .O(sig000003cf)
  );
  XORCY   blk00000181 (
    .CI(sig000003d1),
    .LI(sig0000057b),
    .O(sig000004be)
  );
  MUXCY   blk00000182 (
    .CI(sig000003d1),
    .DI(sig000006c3),
    .S(sig0000057b),
    .O(sig000003d0)
  );
  XORCY   blk00000183 (
    .CI(sig000003d2),
    .LI(sig0000057a),
    .O(sig000004bd)
  );
  MUXCY   blk00000184 (
    .CI(sig000003d2),
    .DI(sig000006c3),
    .S(sig0000057a),
    .O(sig000003d1)
  );
  XORCY   blk00000185 (
    .CI(sig000006c3),
    .LI(sig00000828),
    .O(sig000004bc)
  );
  MUXCY   blk00000186 (
    .CI(sig000006c3),
    .DI(sig0000024a),
    .S(sig00000828),
    .O(sig000003d2)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000187 (
    .C(clk),
    .D(sig000004b8),
    .Q(sig000004c7)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000188 (
    .C(clk),
    .D(sig000004b7),
    .Q(sig000004c8)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000189 (
    .C(clk),
    .D(sig000004ba),
    .Q(sig000004c9)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000018a (
    .C(clk),
    .D(sig000004cc),
    .Q(sig000003d3)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000018b (
    .C(clk),
    .CE(sig00000001),
    .D(sig000004d0),
    .Q(sig0000040e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000018c (
    .C(clk),
    .CE(sig00000001),
    .D(sig000004d1),
    .Q(sig0000040d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000018d (
    .C(clk),
    .CE(sig00000001),
    .D(sig000004b4),
    .Q(sig0000050d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000018e (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000022c),
    .Q(sig000004b5)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000018f (
    .C(clk),
    .CE(sig00000001),
    .D(sig000004b5),
    .Q(sig00000544)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000190 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000004b6),
    .Q(sig000004b4)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000191 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000004cf),
    .Q(sig000004cb)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000192 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000004b9),
    .Q(sig000004cd)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000193 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000004bb),
    .Q(sig000004ca)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000194 (
    .C(clk),
    .D(sig00000543),
    .Q(sig0000050c)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000195 (
    .C(clk),
    .D(sig00000542),
    .Q(sig0000050b)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000196 (
    .C(clk),
    .D(sig00000541),
    .Q(sig0000050a)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000197 (
    .C(clk),
    .D(sig00000540),
    .Q(sig00000509)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000198 (
    .C(clk),
    .D(sig0000053f),
    .Q(sig00000508)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000199 (
    .C(clk),
    .D(sig0000053e),
    .Q(sig00000507)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000019a (
    .C(clk),
    .D(sig0000053d),
    .Q(sig00000506)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000019b (
    .C(clk),
    .D(sig0000053c),
    .Q(sig00000505)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000019c (
    .C(clk),
    .D(sig0000053b),
    .Q(sig00000504)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000019d (
    .C(clk),
    .D(sig0000053a),
    .Q(sig00000503)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000019e (
    .C(clk),
    .D(sig00000539),
    .Q(sig00000502)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000019f (
    .C(clk),
    .D(sig00000538),
    .Q(sig00000501)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001a0 (
    .C(clk),
    .D(sig00000537),
    .Q(sig00000500)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001a1 (
    .C(clk),
    .D(sig00000536),
    .Q(sig000004ff)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001a2 (
    .C(clk),
    .D(sig00000535),
    .Q(sig000004fe)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001a3 (
    .C(clk),
    .D(sig00000534),
    .Q(sig000004fd)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001a4 (
    .C(clk),
    .D(sig00000533),
    .Q(sig000004fc)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001a5 (
    .C(clk),
    .D(sig00000532),
    .Q(sig000004fb)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001a6 (
    .C(clk),
    .D(sig00000531),
    .Q(sig000004fa)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001a7 (
    .C(clk),
    .D(sig00000530),
    .Q(sig000004f9)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001a8 (
    .C(clk),
    .D(sig0000052f),
    .Q(sig000004f8)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001a9 (
    .C(clk),
    .D(sig0000052e),
    .Q(sig000004f7)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001aa (
    .C(clk),
    .D(sig0000052d),
    .Q(sig000004f6)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001ab (
    .C(clk),
    .D(sig0000052c),
    .Q(sig000004f5)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001ac (
    .C(clk),
    .D(sig0000052b),
    .Q(sig000004f4)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001ad (
    .C(clk),
    .D(sig0000052a),
    .Q(sig000004f3)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001ae (
    .C(clk),
    .D(sig00000529),
    .Q(sig000004f2)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001af (
    .C(clk),
    .D(sig00000528),
    .Q(sig000004f1)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001b0 (
    .C(clk),
    .D(sig00000527),
    .Q(sig000004f0)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001b1 (
    .C(clk),
    .D(sig00000526),
    .Q(sig000004ef)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001b2 (
    .C(clk),
    .D(sig00000525),
    .Q(sig000004ee)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001b3 (
    .C(clk),
    .D(sig00000524),
    .Q(sig000004ed)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001b4 (
    .C(clk),
    .D(sig00000523),
    .Q(sig000004ec)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001b5 (
    .C(clk),
    .D(sig00000522),
    .Q(sig000004eb)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001b6 (
    .C(clk),
    .D(sig00000521),
    .Q(sig000004ea)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001b7 (
    .C(clk),
    .D(sig00000520),
    .Q(sig000004e9)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001b8 (
    .C(clk),
    .D(sig0000051f),
    .Q(sig000004e8)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001b9 (
    .C(clk),
    .D(sig0000051e),
    .Q(sig000004e7)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001ba (
    .C(clk),
    .D(sig0000051d),
    .Q(sig000004e6)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001bb (
    .C(clk),
    .D(sig0000051c),
    .Q(sig000004e5)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001bc (
    .C(clk),
    .D(sig0000051b),
    .Q(sig000004e4)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001bd (
    .C(clk),
    .D(sig0000051a),
    .Q(sig000004e3)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001be (
    .C(clk),
    .D(sig00000519),
    .Q(sig000004e2)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001bf (
    .C(clk),
    .D(sig00000518),
    .Q(sig000004e1)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001c0 (
    .C(clk),
    .D(sig00000517),
    .Q(sig000004e0)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001c1 (
    .C(clk),
    .D(sig00000516),
    .Q(sig000004df)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001c2 (
    .C(clk),
    .D(sig00000515),
    .Q(sig000004de)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001c3 (
    .C(clk),
    .D(sig00000514),
    .Q(sig000004dd)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001c4 (
    .C(clk),
    .D(sig00000513),
    .Q(sig000004dc)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001c5 (
    .C(clk),
    .D(sig00000512),
    .Q(sig000004db)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001c6 (
    .C(clk),
    .D(sig00000511),
    .Q(sig000004da)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001c7 (
    .C(clk),
    .D(sig00000510),
    .Q(sig000004d9)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001c8 (
    .C(clk),
    .D(sig0000050f),
    .Q(sig000004d8)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001c9 (
    .C(clk),
    .D(sig0000050e),
    .Q(sig000004d7)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001ca (
    .C(clk),
    .D(sig000004c6),
    .Q(sig000004d6)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001cb (
    .C(clk),
    .D(sig000004c5),
    .Q(sig000004d5)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001cc (
    .C(clk),
    .D(sig000004c4),
    .Q(sig000004d4)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001cd (
    .C(clk),
    .D(sig000004c3),
    .Q(sig000004d3)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001ce (
    .C(clk),
    .D(sig000004c2),
    .Q(sig000004d2)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001cf (
    .C(clk),
    .D(sig000004c1),
    .Q(sig000003d4)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001d0 (
    .C(clk),
    .D(sig000004c0),
    .Q(sig000003d5)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001d1 (
    .C(clk),
    .D(sig000004bf),
    .Q(sig000004d1)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001d2 (
    .C(clk),
    .D(sig000004be),
    .Q(sig000004d0)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001d3 (
    .C(clk),
    .D(sig000004bd),
    .Q(sig000004cf)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000001d4 (
    .C(clk),
    .D(sig000004bc),
    .Q(sig000004ce)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001d5 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000040f),
    .Q(sig000003d6)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001d6 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000410),
    .Q(sig000003d7)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001d7 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000411),
    .Q(sig000003d8)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001d8 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000412),
    .Q(sig000003d9)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001d9 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000413),
    .Q(sig000003da)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001da (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000414),
    .Q(sig000003db)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001db (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000415),
    .Q(sig000003dc)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001dc (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000416),
    .Q(sig000003dd)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001dd (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000417),
    .Q(sig000003de)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001de (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000418),
    .Q(sig000003df)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001df (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000419),
    .Q(sig000003e0)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001e0 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000041a),
    .Q(sig000003e1)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001e1 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000041b),
    .Q(sig000003e2)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001e2 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000041c),
    .Q(sig000003e3)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001e3 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000041d),
    .Q(sig000003e4)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001e4 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000041e),
    .Q(sig000003e5)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001e5 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000041f),
    .Q(sig000003e6)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001e6 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000420),
    .Q(sig000003e7)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001e7 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000421),
    .Q(sig000003e8)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001e8 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000422),
    .Q(sig000003e9)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001e9 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000423),
    .Q(sig000003ea)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001ea (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000424),
    .Q(sig000003eb)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001eb (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000425),
    .Q(sig000003ec)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001ec (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000426),
    .Q(sig000003ed)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001ed (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000427),
    .Q(sig000003ee)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001ee (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000428),
    .Q(sig000003ef)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001ef (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000429),
    .Q(sig000003f0)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001f0 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000042a),
    .Q(sig000003f1)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001f1 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000042b),
    .Q(sig000003f2)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001f2 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000042c),
    .Q(sig000003f3)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001f3 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000042d),
    .Q(sig000003f4)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001f4 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000042e),
    .Q(sig000003f5)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001f5 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000042f),
    .Q(sig000003f6)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001f6 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000430),
    .Q(sig000003f7)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001f7 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000431),
    .Q(sig000003f8)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001f8 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000432),
    .Q(sig000003f9)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001f9 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000433),
    .Q(sig000003fa)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001fa (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000434),
    .Q(sig000003fb)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001fb (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000435),
    .Q(sig000003fc)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001fc (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000436),
    .Q(sig000003fd)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001fd (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000437),
    .Q(sig000003fe)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001fe (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000438),
    .Q(sig000003ff)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000001ff (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000439),
    .Q(sig00000400)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000200 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000043a),
    .Q(sig00000401)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000201 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000043b),
    .Q(sig00000402)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000202 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000043c),
    .Q(sig00000403)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000203 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000043d),
    .Q(sig00000404)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000204 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000043e),
    .Q(sig00000405)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000205 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000043f),
    .Q(sig00000406)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000206 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000440),
    .Q(sig00000407)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000207 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000441),
    .Q(sig00000408)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000208 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000442),
    .Q(sig00000409)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000209 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000443),
    .Q(sig0000040a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000020a (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000444),
    .Q(sig0000040b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000020b (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000445),
    .Q(sig0000040c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000020c (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000446),
    .Q(sig0000047d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000020d (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000447),
    .Q(sig0000047e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000020e (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000448),
    .Q(sig0000047f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000020f (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000449),
    .Q(sig00000480)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000210 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000044a),
    .Q(sig00000481)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000211 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000044b),
    .Q(sig00000482)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000212 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000044c),
    .Q(sig00000483)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000213 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000044d),
    .Q(sig00000484)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000214 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000044e),
    .Q(sig00000485)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000215 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000044f),
    .Q(sig00000486)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000216 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000450),
    .Q(sig00000487)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000217 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000451),
    .Q(sig00000488)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000218 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000452),
    .Q(sig00000489)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000219 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000453),
    .Q(sig0000048a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000021a (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000454),
    .Q(sig0000048b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000021b (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000455),
    .Q(sig0000048c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000021c (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000456),
    .Q(sig0000048d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000021d (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000457),
    .Q(sig0000048e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000021e (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000458),
    .Q(sig0000048f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000021f (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000459),
    .Q(sig00000490)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000220 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000045a),
    .Q(sig00000491)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000221 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000045b),
    .Q(sig00000492)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000222 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000045c),
    .Q(sig00000493)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000223 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000045d),
    .Q(sig00000494)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000224 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000045e),
    .Q(sig00000495)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000225 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000045f),
    .Q(sig00000496)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000226 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000460),
    .Q(sig00000497)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000227 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000461),
    .Q(sig00000498)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000228 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000462),
    .Q(sig00000499)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000229 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000463),
    .Q(sig0000049a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000022a (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000464),
    .Q(sig0000049b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000022b (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000465),
    .Q(sig0000049c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000022c (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000466),
    .Q(sig0000049d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000022d (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000467),
    .Q(sig0000049e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000022e (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000468),
    .Q(sig0000049f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000022f (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000469),
    .Q(sig000004a0)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000230 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000046a),
    .Q(sig000004a1)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000231 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000046b),
    .Q(sig000004a2)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000232 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000046c),
    .Q(sig000004a3)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000233 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000046d),
    .Q(sig000004a4)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000234 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000046e),
    .Q(sig000004a5)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000235 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000046f),
    .Q(sig000004a6)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000236 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000470),
    .Q(sig000004a7)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000237 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000471),
    .Q(sig000004a8)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000238 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000472),
    .Q(sig000004a9)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000239 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000473),
    .Q(sig000004aa)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000023a (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000474),
    .Q(sig000004ab)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000023b (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000475),
    .Q(sig000004ac)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000023c (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000476),
    .Q(sig000004ad)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000023d (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000477),
    .Q(sig000004ae)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000023e (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000478),
    .Q(sig000004af)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000023f (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000479),
    .Q(sig000004b0)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000240 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000047a),
    .Q(sig000004b1)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000241 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000047b),
    .Q(sig000004b2)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000242 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000047c),
    .Q(sig000004b3)
  );
  MUXF8   blk00000243 (
    .I0(sig00000586),
    .I1(sig00000585),
    .S(sig00000595),
    .O(sig00000584)
  );
  MUXF7   blk00000244 (
    .I0(sig00000598),
    .I1(sig00000597),
    .S(sig00000596),
    .O(sig00000585)
  );
  MUXF7   blk00000245 (
    .I0(sig0000059a),
    .I1(sig00000599),
    .S(sig00000596),
    .O(sig00000586)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000246 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000003d5),
    .Q(sig00000596)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000247 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000003d4),
    .Q(sig00000595)
  );
  MUXCY   blk00000248 (
    .CI(sig000005c7),
    .DI(sig000006c3),
    .S(sig000005b7),
    .O(sig000005c6)
  );
  MUXCY   blk00000249 (
    .CI(sig000005c8),
    .DI(sig000006c3),
    .S(sig000005b8),
    .O(sig000005c7)
  );
  MUXCY   blk0000024a (
    .CI(sig000005c9),
    .DI(sig000006c3),
    .S(sig000005b9),
    .O(sig000005c8)
  );
  MUXCY   blk0000024b (
    .CI(sig000005ca),
    .DI(sig000006c3),
    .S(sig000005ba),
    .O(sig000005c9)
  );
  MUXCY   blk0000024c (
    .CI(sig000005cb),
    .DI(sig000006c3),
    .S(sig000005bb),
    .O(sig000005ca)
  );
  MUXCY   blk0000024d (
    .CI(sig000005cc),
    .DI(sig000006c3),
    .S(sig000005bc),
    .O(sig000005cb)
  );
  MUXCY   blk0000024e (
    .CI(sig000005cd),
    .DI(sig000006c3),
    .S(sig000005bd),
    .O(sig000005cc)
  );
  MUXCY   blk0000024f (
    .CI(sig000005ce),
    .DI(sig000006c3),
    .S(sig000005be),
    .O(sig000005cd)
  );
  MUXCY   blk00000250 (
    .CI(sig000005cf),
    .DI(sig000006c3),
    .S(sig000005bf),
    .O(sig000005ce)
  );
  MUXCY   blk00000251 (
    .CI(sig000005d0),
    .DI(sig000006c3),
    .S(sig000005c0),
    .O(sig000005cf)
  );
  MUXCY   blk00000252 (
    .CI(sig000005d1),
    .DI(sig000006c3),
    .S(sig000005c1),
    .O(sig000005d0)
  );
  MUXCY   blk00000253 (
    .CI(sig000005d2),
    .DI(sig000006c3),
    .S(sig000005c2),
    .O(sig000005d1)
  );
  MUXCY   blk00000254 (
    .CI(sig000005d3),
    .DI(sig000006c3),
    .S(sig000005c3),
    .O(sig000005d2)
  );
  MUXCY   blk00000255 (
    .CI(sig00000001),
    .DI(sig000006c3),
    .S(sig000005c4),
    .O(sig000005d3)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000256 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000005c6),
    .Q(sig000005c5)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000257 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000005c7),
    .Q(sig000005ab)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000258 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000005c8),
    .Q(sig000005aa)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000259 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000005c9),
    .Q(sig000005ad)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000025a (
    .C(clk),
    .CE(sig00000001),
    .D(sig000005ca),
    .Q(sig000005ae)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000025b (
    .C(clk),
    .CE(sig00000001),
    .D(sig000005cb),
    .Q(sig000005af)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000025c (
    .C(clk),
    .CE(sig00000001),
    .D(sig000005cc),
    .Q(sig000005ac)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000025d (
    .C(clk),
    .CE(sig00000001),
    .D(sig000005cd),
    .Q(sig000005b1)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000025e (
    .C(clk),
    .CE(sig00000001),
    .D(sig000005ce),
    .Q(sig000005b2)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000025f (
    .C(clk),
    .CE(sig00000001),
    .D(sig000005cf),
    .Q(sig000005b3)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000260 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000005d0),
    .Q(sig000005b0)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000261 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000005d1),
    .Q(sig000005b4)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000262 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000005d2),
    .Q(sig000005b5)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000263 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000005d3),
    .Q(sig000005b6)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000264 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000584),
    .Q(sig000004cc)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000265 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000001),
    .Q(sig0000059c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000266 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000587),
    .Q(sig0000059d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000267 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000588),
    .Q(sig0000059b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000268 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000589),
    .Q(sig0000059f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000269 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000058a),
    .Q(sig000005a0)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000026a (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000058b),
    .Q(sig000005a1)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000026b (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000058c),
    .Q(sig0000059e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000026c (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000058d),
    .Q(sig000005a3)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000026d (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000058e),
    .Q(sig000005a4)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000026e (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000058f),
    .Q(sig000005a5)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000026f (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000590),
    .Q(sig000005a2)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000270 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000591),
    .Q(sig000005a7)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000271 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000592),
    .Q(sig000005a8)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000272 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000593),
    .Q(sig000005a9)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000273 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000594),
    .Q(sig000005a6)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000274 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000004ca),
    .Q(sig00000697)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000275 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000050d),
    .Q(sig00000696)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000276 (
    .C(clk),
    .D(sig00000571),
    .Q(sig00000665)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000277 (
    .C(clk),
    .D(sig00000570),
    .Q(sig00000664)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000278 (
    .C(clk),
    .D(sig0000056f),
    .Q(sig00000663)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000279 (
    .C(clk),
    .D(sig0000056e),
    .Q(sig00000662)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000027a (
    .C(clk),
    .D(sig0000056d),
    .Q(sig00000661)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000027b (
    .C(clk),
    .D(sig0000056c),
    .Q(sig00000660)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000027c (
    .C(clk),
    .D(sig0000056b),
    .Q(sig0000065f)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000027d (
    .C(clk),
    .D(sig0000056a),
    .Q(sig0000065e)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000027e (
    .C(clk),
    .D(sig00000569),
    .Q(sig0000065d)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000027f (
    .C(clk),
    .D(sig00000568),
    .Q(sig0000065c)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000280 (
    .C(clk),
    .D(sig00000567),
    .Q(sig0000065b)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000281 (
    .C(clk),
    .D(sig00000566),
    .Q(sig0000065a)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000282 (
    .C(clk),
    .D(sig00000565),
    .Q(sig00000659)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000283 (
    .C(clk),
    .D(sig00000564),
    .Q(sig00000658)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000284 (
    .C(clk),
    .D(sig00000563),
    .Q(sig00000657)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000285 (
    .C(clk),
    .D(sig00000562),
    .Q(sig00000656)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000286 (
    .C(clk),
    .D(sig00000561),
    .Q(sig00000655)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000287 (
    .C(clk),
    .D(sig00000560),
    .Q(sig00000654)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000288 (
    .C(clk),
    .D(sig0000055f),
    .Q(sig00000653)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000289 (
    .C(clk),
    .D(sig0000055e),
    .Q(sig00000652)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000028a (
    .C(clk),
    .D(sig0000055d),
    .Q(sig00000651)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000028b (
    .C(clk),
    .D(sig0000055c),
    .Q(sig00000650)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000028c (
    .C(clk),
    .D(sig0000055b),
    .Q(sig0000064f)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000028d (
    .C(clk),
    .D(sig0000055a),
    .Q(sig0000064e)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000028e (
    .C(clk),
    .D(sig00000559),
    .Q(sig0000064d)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000028f (
    .C(clk),
    .D(sig00000558),
    .Q(sig0000064c)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000290 (
    .C(clk),
    .D(sig00000557),
    .Q(sig0000064b)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000291 (
    .C(clk),
    .D(sig00000556),
    .Q(sig0000064a)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000292 (
    .C(clk),
    .D(sig00000555),
    .Q(sig00000649)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000293 (
    .C(clk),
    .D(sig00000554),
    .Q(sig00000648)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000294 (
    .C(clk),
    .D(sig00000553),
    .Q(sig00000647)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000295 (
    .C(clk),
    .D(sig00000552),
    .Q(sig00000646)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000296 (
    .C(clk),
    .D(sig00000551),
    .Q(sig00000645)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000297 (
    .C(clk),
    .D(sig00000550),
    .Q(sig00000644)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000298 (
    .C(clk),
    .D(sig0000054f),
    .Q(sig00000643)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000299 (
    .C(clk),
    .D(sig0000054e),
    .Q(sig00000642)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000029a (
    .C(clk),
    .D(sig0000054d),
    .Q(sig00000641)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000029b (
    .C(clk),
    .D(sig0000054c),
    .Q(sig00000640)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000029c (
    .C(clk),
    .D(sig0000054b),
    .Q(sig0000063f)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000029d (
    .C(clk),
    .D(sig0000054a),
    .Q(sig0000063e)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000029e (
    .C(clk),
    .D(sig00000549),
    .Q(sig0000063d)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000029f (
    .C(clk),
    .D(sig00000548),
    .Q(sig0000063c)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000002a0 (
    .C(clk),
    .D(sig00000547),
    .Q(sig0000063b)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000002a1 (
    .C(clk),
    .D(sig00000546),
    .Q(sig0000063a)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000002a2 (
    .C(clk),
    .D(sig00000545),
    .Q(sig00000639)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000002a3 (
    .C(clk),
    .D(sig00000579),
    .Q(sig0000069f)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000002a4 (
    .C(clk),
    .D(sig00000578),
    .Q(sig0000069e)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000002a5 (
    .C(clk),
    .D(sig00000577),
    .Q(sig0000069d)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000002a6 (
    .C(clk),
    .D(sig00000576),
    .Q(sig0000069c)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000002a7 (
    .C(clk),
    .D(sig00000575),
    .Q(sig0000069b)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000002a8 (
    .C(clk),
    .D(sig00000574),
    .Q(sig0000069a)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000002a9 (
    .C(clk),
    .D(sig00000573),
    .Q(sig00000699)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000002aa (
    .C(clk),
    .D(sig00000572),
    .Q(sig00000698)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000002ab (
    .C(clk),
    .D(sig0000047d),
    .Q(sig00000600)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000002ac (
    .C(clk),
    .D(sig0000047e),
    .Q(sig000005ff)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000002ad (
    .C(clk),
    .D(sig0000047f),
    .Q(sig000005fe)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000002ae (
    .C(clk),
    .D(sig00000480),
    .Q(sig000005fd)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000002af (
    .C(clk),
    .D(sig00000481),
    .Q(sig000005fc)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000002b0 (
    .C(clk),
    .D(sig00000482),
    .Q(sig000005fb)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000002b1 (
    .C(clk),
    .D(sig00000483),
    .Q(sig000005fa)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000002b2 (
    .C(clk),
    .D(sig00000484),
    .Q(sig000005f9)
  );
  XORCY   blk000002b3 (
    .CI(sig000006a2),
    .LI(sig00000827),
    .O(sig000006a0)
  );
  XORCY   blk000002b4 (
    .CI(sig000006a4),
    .LI(sig00000811),
    .O(sig000006a1)
  );
  MUXCY   blk000002b5 (
    .CI(sig000006a4),
    .DI(sig00000608),
    .S(sig00000811),
    .O(sig000006a2)
  );
  XORCY   blk000002b6 (
    .CI(sig000006a6),
    .LI(sig00000812),
    .O(sig000006a3)
  );
  MUXCY   blk000002b7 (
    .CI(sig000006a6),
    .DI(sig00000607),
    .S(sig00000812),
    .O(sig000006a4)
  );
  XORCY   blk000002b8 (
    .CI(sig000006a8),
    .LI(sig00000813),
    .O(sig000006a5)
  );
  MUXCY   blk000002b9 (
    .CI(sig000006a8),
    .DI(sig00000606),
    .S(sig00000813),
    .O(sig000006a6)
  );
  XORCY   blk000002ba (
    .CI(sig000006aa),
    .LI(sig00000814),
    .O(sig000006a7)
  );
  MUXCY   blk000002bb (
    .CI(sig000006aa),
    .DI(sig00000605),
    .S(sig00000814),
    .O(sig000006a8)
  );
  XORCY   blk000002bc (
    .CI(sig000006ac),
    .LI(sig00000815),
    .O(sig000006a9)
  );
  MUXCY   blk000002bd (
    .CI(sig000006ac),
    .DI(sig00000604),
    .S(sig00000815),
    .O(sig000006aa)
  );
  XORCY   blk000002be (
    .CI(sig000006ae),
    .LI(sig00000816),
    .O(sig000006ab)
  );
  MUXCY   blk000002bf (
    .CI(sig000006ae),
    .DI(sig00000603),
    .S(sig00000816),
    .O(sig000006ac)
  );
  XORCY   blk000002c0 (
    .CI(sig000006b0),
    .LI(sig00000817),
    .O(sig000006ad)
  );
  MUXCY   blk000002c1 (
    .CI(sig000006b0),
    .DI(sig00000602),
    .S(sig00000817),
    .O(sig000006ae)
  );
  XORCY   blk000002c2 (
    .CI(sig00000001),
    .LI(sig00000818),
    .O(sig000006af)
  );
  MUXCY   blk000002c3 (
    .CI(sig00000001),
    .DI(sig00000601),
    .S(sig00000818),
    .O(sig000006b0)
  );
  XORCY   blk000002c4 (
    .CI(sig000006b3),
    .LI(sig000005dc),
    .O(sig000006b1)
  );
  XORCY   blk000002c5 (
    .CI(sig000006b5),
    .LI(sig000005db),
    .O(sig000006b2)
  );
  MUXCY   blk000002c6 (
    .CI(sig000006b5),
    .DI(sig00000608),
    .S(sig000005db),
    .O(sig000006b3)
  );
  XORCY   blk000002c7 (
    .CI(sig000006b7),
    .LI(sig000005da),
    .O(sig000006b4)
  );
  MUXCY   blk000002c8 (
    .CI(sig000006b7),
    .DI(sig00000607),
    .S(sig000005da),
    .O(sig000006b5)
  );
  XORCY   blk000002c9 (
    .CI(sig000006b9),
    .LI(sig000005d9),
    .O(sig000006b6)
  );
  MUXCY   blk000002ca (
    .CI(sig000006b9),
    .DI(sig00000606),
    .S(sig000005d9),
    .O(sig000006b7)
  );
  XORCY   blk000002cb (
    .CI(sig000006bb),
    .LI(sig000005d8),
    .O(sig000006b8)
  );
  MUXCY   blk000002cc (
    .CI(sig000006bb),
    .DI(sig00000605),
    .S(sig000005d8),
    .O(sig000006b9)
  );
  XORCY   blk000002cd (
    .CI(sig000006bd),
    .LI(sig000005d7),
    .O(sig000006ba)
  );
  MUXCY   blk000002ce (
    .CI(sig000006bd),
    .DI(sig00000604),
    .S(sig000005d7),
    .O(sig000006bb)
  );
  XORCY   blk000002cf (
    .CI(sig000006bf),
    .LI(sig000005d6),
    .O(sig000006bc)
  );
  MUXCY   blk000002d0 (
    .CI(sig000006bf),
    .DI(sig00000603),
    .S(sig000005d6),
    .O(sig000006bd)
  );
  XORCY   blk000002d1 (
    .CI(sig000006c1),
    .LI(sig000005d5),
    .O(sig000006be)
  );
  MUXCY   blk000002d2 (
    .CI(sig000006c1),
    .DI(sig00000602),
    .S(sig000005d5),
    .O(sig000006bf)
  );
  XORCY   blk000002d3 (
    .CI(sig000006c3),
    .LI(sig000005d4),
    .O(sig000006c0)
  );
  MUXCY   blk000002d4 (
    .CI(sig000006c3),
    .DI(sig00000601),
    .S(sig000005d4),
    .O(sig000006c1)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002d5 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000006b1),
    .Q(sig000005f7)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002d6 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000006b2),
    .Q(sig000005f6)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002d7 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000006b4),
    .Q(sig000005f5)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002d8 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000006b6),
    .Q(sig000005f4)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002d9 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000006b8),
    .Q(sig000005f3)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002da (
    .C(clk),
    .CE(sig00000001),
    .D(sig000006ba),
    .Q(sig000005f2)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002db (
    .C(clk),
    .CE(sig00000001),
    .D(sig000006bc),
    .Q(sig000005f1)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002dc (
    .C(clk),
    .CE(sig00000001),
    .D(sig000006be),
    .Q(sig000005f0)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002dd (
    .C(clk),
    .CE(sig00000001),
    .D(sig000006c0),
    .Q(sig000005ef)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002de (
    .C(clk),
    .CE(sig00000001),
    .D(sig000006a0),
    .Q(sig000005ee)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002df (
    .C(clk),
    .CE(sig00000001),
    .D(sig000006a1),
    .Q(sig000005ed)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002e0 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000006a3),
    .Q(sig000005ec)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002e1 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000006a5),
    .Q(sig000005eb)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002e2 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000006a7),
    .Q(sig000005ea)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002e3 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000006a9),
    .Q(sig000005e9)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002e4 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000006ab),
    .Q(sig000005e8)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002e5 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000006ad),
    .Q(sig000005e7)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002e6 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000006af),
    .Q(sig000005e6)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002e7 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000005e5),
    .Q(sig000001c2)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002e8 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000005e4),
    .Q(sig000001c1)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002e9 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000005e3),
    .Q(sig000001c0)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002ea (
    .C(clk),
    .CE(sig00000001),
    .D(sig000005e2),
    .Q(sig000001bf)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002eb (
    .C(clk),
    .CE(sig00000001),
    .D(sig000005e1),
    .Q(sig000001be)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002ec (
    .C(clk),
    .CE(sig00000001),
    .D(sig000005e0),
    .Q(sig000001bd)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002ed (
    .C(clk),
    .CE(sig00000001),
    .D(sig000005df),
    .Q(sig000001bc)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002ee (
    .C(clk),
    .CE(sig00000001),
    .D(sig000005de),
    .Q(sig000001bb)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002ef (
    .C(clk),
    .CE(sig00000001),
    .D(sig000005dd),
    .Q(sig000001ba)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002f0 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000695),
    .Q(sig000001b9)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002f1 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000694),
    .Q(sig000001b8)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002f2 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000693),
    .Q(sig000001b7)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002f3 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000692),
    .Q(sig000001b6)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002f4 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000691),
    .Q(sig000001b5)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002f5 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000690),
    .Q(sig000001b4)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002f6 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000068f),
    .Q(sig000001b3)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002f7 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000068e),
    .Q(sig000001b2)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002f8 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000068d),
    .Q(sig000001b1)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002f9 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000068c),
    .Q(sig000001b0)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002fa (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000068b),
    .Q(sig000001af)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002fb (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000068a),
    .Q(sig000001ae)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002fc (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000689),
    .Q(sig000001ad)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002fd (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000688),
    .Q(sig000001ac)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002fe (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000687),
    .Q(sig000001ab)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002ff (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000686),
    .Q(sig000001aa)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000300 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000685),
    .Q(sig000001a9)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000301 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000684),
    .Q(sig000001a8)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000302 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000683),
    .Q(sig000001a7)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000303 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000682),
    .Q(sig000001a6)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000304 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000681),
    .Q(sig000001a5)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000305 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000680),
    .Q(sig000001a4)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000306 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000067f),
    .Q(sig000001a3)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000307 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000067e),
    .Q(sig000001a2)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000308 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000067d),
    .Q(sig000001a1)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000309 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000067c),
    .Q(sig000001a0)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000030a (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000067b),
    .Q(sig0000019f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000030b (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000067a),
    .Q(sig0000019e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000030c (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000679),
    .Q(sig0000019d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000030d (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000678),
    .Q(sig0000019c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000030e (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000677),
    .Q(sig0000019b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000030f (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000676),
    .Q(sig0000019a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000310 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000675),
    .Q(sig00000199)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000311 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000674),
    .Q(sig00000198)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000312 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000673),
    .Q(sig00000197)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000313 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000672),
    .Q(sig00000196)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000314 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000671),
    .Q(sig00000195)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000315 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000670),
    .Q(sig00000194)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000316 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000066f),
    .Q(sig00000193)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000317 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000066e),
    .Q(sig00000192)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000318 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000066d),
    .Q(sig00000191)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000319 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000066c),
    .Q(sig00000190)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000031a (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000066b),
    .Q(sig0000018f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000031b (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000066a),
    .Q(sig0000018e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000031c (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000669),
    .Q(sig0000018d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000031d (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000668),
    .Q(sig0000018c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000031e (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000667),
    .Q(sig0000018b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000031f (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000072),
    .Q(sig00000002)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000320 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000073),
    .Q(sig00000003)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000321 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000074),
    .Q(sig00000004)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000322 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000075),
    .Q(sig00000005)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000323 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000076),
    .Q(sig00000006)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000324 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000077),
    .Q(sig00000007)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000325 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000078),
    .Q(sig00000008)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000326 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000079),
    .Q(sig00000009)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000327 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000007a),
    .Q(sig0000000a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000328 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000007b),
    .Q(sig0000000b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000329 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000007c),
    .Q(sig0000000c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000032a (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000007d),
    .Q(sig0000000d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000032b (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000007e),
    .Q(sig0000000e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000032c (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000007f),
    .Q(sig0000000f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000032d (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000080),
    .Q(sig00000010)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000032e (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000081),
    .Q(sig00000011)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000032f (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000082),
    .Q(sig00000012)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000330 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000083),
    .Q(sig00000013)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000331 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000084),
    .Q(sig00000014)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000332 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000085),
    .Q(sig00000015)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000333 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000086),
    .Q(sig00000016)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000334 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000087),
    .Q(sig00000017)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000335 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000088),
    .Q(sig00000018)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000336 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000089),
    .Q(sig00000019)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000337 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000008a),
    .Q(sig0000001a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000338 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000008b),
    .Q(sig0000001b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000339 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000008c),
    .Q(sig0000001c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000033a (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000008d),
    .Q(sig0000001d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000033b (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000008e),
    .Q(sig0000001e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000033c (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000008f),
    .Q(sig0000001f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000033d (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000090),
    .Q(sig00000020)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000033e (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000091),
    .Q(sig00000021)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000033f (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000092),
    .Q(sig00000022)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000340 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000093),
    .Q(sig00000023)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000341 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000094),
    .Q(sig00000024)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000342 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000095),
    .Q(sig00000025)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000343 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000096),
    .Q(sig00000026)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000344 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000097),
    .Q(sig00000027)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000345 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000098),
    .Q(sig00000028)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000346 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000099),
    .Q(sig00000029)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000347 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000009a),
    .Q(sig0000002a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000348 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000009b),
    .Q(sig0000002b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000349 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000009c),
    .Q(sig0000002c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000034a (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000009d),
    .Q(sig0000002d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000034b (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000009e),
    .Q(sig0000002e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000034c (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000009f),
    .Q(sig0000002f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000034d (
    .C(clk),
    .CE(sig00000001),
    .D(sig000000a0),
    .Q(sig00000030)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000034e (
    .C(clk),
    .CE(sig00000001),
    .D(sig000000a1),
    .Q(sig00000031)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000034f (
    .C(clk),
    .CE(sig00000001),
    .D(sig000000a2),
    .Q(sig00000032)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000350 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000000a3),
    .Q(sig00000033)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000351 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000000a4),
    .Q(sig00000034)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000352 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000000a5),
    .Q(sig00000035)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000353 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000000a6),
    .Q(sig00000036)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000354 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000000a7),
    .Q(sig00000037)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000355 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000000a8),
    .Q(sig00000038)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000356 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000000a9),
    .Q(sig00000039)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000357 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000000aa),
    .Q(sig0000003a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000358 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000000ab),
    .Q(sig0000003b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000359 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000000ac),
    .Q(sig0000003c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000035a (
    .C(clk),
    .CE(sig00000001),
    .D(sig000000ad),
    .Q(sig0000003d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000035b (
    .C(clk),
    .CE(sig00000001),
    .D(sig000000ae),
    .Q(sig0000003e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000035c (
    .C(clk),
    .CE(sig00000001),
    .D(sig000000af),
    .Q(sig0000003f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000035d (
    .C(clk),
    .CE(sig00000001),
    .D(sig000000b0),
    .Q(sig00000040)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000035e (
    .C(clk),
    .CE(sig00000001),
    .D(sig000000b1),
    .Q(sig00000041)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000035f (
    .C(clk),
    .CE(sig00000001),
    .D(sig000000b2),
    .Q(sig00000042)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000360 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000000b3),
    .Q(sig00000043)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000361 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000000b4),
    .Q(sig00000044)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000362 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000000b5),
    .Q(sig00000045)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000363 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000000b6),
    .Q(sig00000046)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000364 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000000b7),
    .Q(sig00000047)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000365 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000000b8),
    .Q(sig00000048)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000366 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000000b9),
    .Q(sig00000049)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000367 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000000ba),
    .Q(sig0000004a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000368 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000000bb),
    .Q(sig0000004b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000369 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000000bc),
    .Q(sig0000004c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000036a (
    .C(clk),
    .CE(sig00000001),
    .D(sig000000bd),
    .Q(sig0000004d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000036b (
    .C(clk),
    .CE(sig00000001),
    .D(sig000000be),
    .Q(sig0000004e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000036c (
    .C(clk),
    .CE(sig00000001),
    .D(sig000000bf),
    .Q(sig0000004f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000036d (
    .C(clk),
    .CE(sig00000001),
    .D(sig000000c0),
    .Q(sig00000050)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000036e (
    .C(clk),
    .CE(sig00000001),
    .D(sig000000c1),
    .Q(sig00000051)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000036f (
    .C(clk),
    .CE(sig00000001),
    .D(sig000000c2),
    .Q(sig00000052)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000370 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000000c3),
    .Q(sig00000053)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000371 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000000c4),
    .Q(sig00000054)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000372 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000000c5),
    .Q(sig00000055)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000373 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000000c6),
    .Q(sig00000056)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000374 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000000c7),
    .Q(sig00000057)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000375 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000000c8),
    .Q(sig00000058)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000376 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000000c9),
    .Q(sig00000059)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000377 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000000ca),
    .Q(sig0000005a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000378 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000000cb),
    .Q(sig0000005b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000379 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000000cc),
    .Q(sig0000005c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000037a (
    .C(clk),
    .CE(sig00000001),
    .D(sig000000cd),
    .Q(sig0000005d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000037b (
    .C(clk),
    .CE(sig00000001),
    .D(sig000000ce),
    .Q(sig0000005e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000037c (
    .C(clk),
    .CE(sig00000001),
    .D(sig000000cf),
    .Q(sig0000005f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000037d (
    .C(clk),
    .CE(sig00000001),
    .D(sig000000d0),
    .Q(sig00000060)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000037e (
    .C(clk),
    .CE(sig00000001),
    .D(sig000000d1),
    .Q(sig00000061)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000037f (
    .C(clk),
    .CE(sig00000001),
    .D(sig000000d2),
    .Q(sig00000062)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000380 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000000d3),
    .Q(sig00000063)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000381 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000000d4),
    .Q(sig00000064)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000382 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000000d5),
    .Q(sig00000065)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000383 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000000d6),
    .Q(sig00000066)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000384 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000000d7),
    .Q(sig00000067)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000385 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000000d8),
    .Q(sig00000068)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000386 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000000d9),
    .Q(sig00000069)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000387 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000000da),
    .Q(sig0000006a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000388 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000000db),
    .Q(sig0000006b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000389 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000000dc),
    .Q(sig0000006c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000038a (
    .C(clk),
    .CE(sig00000001),
    .D(sig000000dd),
    .Q(sig0000006d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000038b (
    .C(clk),
    .CE(sig00000001),
    .D(sig000000de),
    .Q(sig0000006e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000038c (
    .C(clk),
    .CE(sig00000001),
    .D(sig000000df),
    .Q(sig0000006f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000038d (
    .C(clk),
    .CE(sig00000001),
    .D(sig000000e0),
    .Q(sig00000070)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000038e (
    .C(clk),
    .CE(sig00000001),
    .D(sig000000e1),
    .Q(sig00000071)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000038f (
    .C(clk),
    .CE(sig00000001),
    .D(sig000001c1),
    .Q(sig0000011e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000390 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000001c0),
    .Q(sig0000011f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000391 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000001bf),
    .Q(sig00000120)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000392 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000001be),
    .Q(sig00000121)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000393 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000001bd),
    .Q(sig00000122)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000394 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000001bc),
    .Q(sig00000123)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000395 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000001bb),
    .Q(sig00000124)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000396 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000001ba),
    .Q(sig00000125)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000397 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000001b9),
    .Q(sig00000126)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000398 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000001b8),
    .Q(sig00000127)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000399 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000001b7),
    .Q(sig00000128)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000039a (
    .C(clk),
    .CE(sig00000001),
    .D(sig000001b6),
    .Q(sig00000129)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000039b (
    .C(clk),
    .CE(sig00000001),
    .D(sig000001b5),
    .Q(sig0000012a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000039c (
    .C(clk),
    .CE(sig00000001),
    .D(sig000001b4),
    .Q(sig0000012b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000039d (
    .C(clk),
    .CE(sig00000001),
    .D(sig000001b3),
    .Q(sig0000012c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000039e (
    .C(clk),
    .CE(sig00000001),
    .D(sig000001b2),
    .Q(sig0000012d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000039f (
    .C(clk),
    .CE(sig00000001),
    .D(sig000001b1),
    .Q(sig0000012e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003a0 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000001b0),
    .Q(sig0000012f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003a1 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000001af),
    .Q(sig00000130)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003a2 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000001ae),
    .Q(sig00000131)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003a3 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000001ad),
    .Q(sig00000132)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003a4 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000001ac),
    .Q(sig00000133)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003a5 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000001ab),
    .Q(sig00000134)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003a6 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000001aa),
    .Q(sig00000135)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003a7 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000001a9),
    .Q(sig00000136)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003a8 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000001a8),
    .Q(sig00000137)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003a9 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000001a7),
    .Q(sig00000138)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003aa (
    .C(clk),
    .CE(sig00000001),
    .D(sig000001a6),
    .Q(sig00000139)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003ab (
    .C(clk),
    .CE(sig00000001),
    .D(sig000001a5),
    .Q(sig0000013a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003ac (
    .C(clk),
    .CE(sig00000001),
    .D(sig000001a4),
    .Q(sig0000013b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003ad (
    .C(clk),
    .CE(sig00000001),
    .D(sig000001a3),
    .Q(sig0000013c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003ae (
    .C(clk),
    .CE(sig00000001),
    .D(sig000001a2),
    .Q(sig0000013d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003af (
    .C(clk),
    .CE(sig00000001),
    .D(sig000001a1),
    .Q(sig0000013e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003b0 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000001a0),
    .Q(sig0000013f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003b1 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000019f),
    .Q(sig00000140)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003b2 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000019e),
    .Q(sig00000141)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003b3 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000019d),
    .Q(sig00000142)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003b4 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000019c),
    .Q(sig00000143)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003b5 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000019b),
    .Q(sig00000144)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003b6 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000019a),
    .Q(sig00000145)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003b7 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000199),
    .Q(sig00000146)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003b8 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000198),
    .Q(sig00000147)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003b9 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000197),
    .Q(sig00000148)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003ba (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000196),
    .Q(sig00000149)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003bb (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000195),
    .Q(sig0000014a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003bc (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000194),
    .Q(sig0000014b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003bd (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000193),
    .Q(sig0000014c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003be (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000192),
    .Q(sig0000014d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003bf (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000191),
    .Q(sig0000014e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003c0 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000190),
    .Q(sig0000014f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003c1 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000018f),
    .Q(sig00000150)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003c2 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000018e),
    .Q(sig00000151)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003c3 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000018d),
    .Q(sig00000152)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003c4 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000018c),
    .Q(sig00000153)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003c5 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000018b),
    .Q(sig00000154)
  );
  MUXF7   blk000003c6 (
    .I0(sig000006c2),
    .I1(sig000006c3),
    .S(sig0000011a),
    .O(NLW_blk000003c6_O_UNCONNECTED)
  );
  MUXF7   blk000003c7 (
    .I0(sig000006c4),
    .I1(sig000006c6),
    .S(sig0000011a),
    .O(sig000006c8)
  );
  MUXF7   blk000003c8 (
    .I0(sig000006c5),
    .I1(sig000006c7),
    .S(sig0000011a),
    .O(sig000006c9)
  );
  MUXF7   blk000003c9 (
    .I0(sig000006ca),
    .I1(sig000006ce),
    .S(sig00000118),
    .O(sig000006d1)
  );
  MUXF7   blk000003ca (
    .I0(sig000006cb),
    .I1(sig000006cf),
    .S(sig00000118),
    .O(sig000006d2)
  );
  MUXF7   blk000003cb (
    .I0(sig000006cc),
    .I1(sig000006d0),
    .S(sig00000118),
    .O(sig000006d3)
  );
  MUXF7   blk000003cc (
    .I0(sig000006cd),
    .I1(sig000006c3),
    .S(sig00000118),
    .O(NLW_blk000003cc_O_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003cd (
    .C(clk),
    .CE(sig00000001),
    .D(sig000006c9),
    .Q(sig0000011c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003ce (
    .C(clk),
    .CE(sig00000001),
    .D(sig000006c8),
    .Q(sig0000011d)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000003cf (
    .C(clk),
    .D(sig000006d1),
    .Q(sig000006e4)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000003d0 (
    .C(clk),
    .D(sig000006d2),
    .Q(sig0000011a)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000003d1 (
    .C(clk),
    .D(sig000006d3),
    .Q(sig000006e3)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003d2 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000011a),
    .Q(sig00000187)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003d3 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000011b),
    .Q(sig00000186)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003d4 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000006d4),
    .Q(sig00000157)
  );
  MUXCY   blk000003d5 (
    .CI(sig000006fb),
    .DI(sig000006c3),
    .S(sig000006dc),
    .O(sig000006fa)
  );
  MUXCY   blk000003d6 (
    .CI(sig000006fc),
    .DI(sig000006c3),
    .S(sig000006db),
    .O(sig000006fb)
  );
  MUXCY   blk000003d7 (
    .CI(sig000006fd),
    .DI(sig000006c3),
    .S(sig000006da),
    .O(sig000006fc)
  );
  MUXCY   blk000003d8 (
    .CI(sig000006fe),
    .DI(sig000006c3),
    .S(sig000006d9),
    .O(sig000006fd)
  );
  MUXCY   blk000003d9 (
    .CI(sig000006ff),
    .DI(sig000006c3),
    .S(sig000006d8),
    .O(sig000006fe)
  );
  MUXCY   blk000003da (
    .CI(sig00000700),
    .DI(sig000006c3),
    .S(sig000006d7),
    .O(sig000006ff)
  );
  MUXCY   blk000003db (
    .CI(sig00000701),
    .DI(sig000006c3),
    .S(sig000006d6),
    .O(sig00000700)
  );
  MUXCY   blk000003dc (
    .CI(sig00000001),
    .DI(sig000006c3),
    .S(sig000006d5),
    .O(sig00000701)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003dd (
    .C(clk),
    .CE(sig00000001),
    .D(sig000006fa),
    .Q(sig00000118)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003de (
    .C(clk),
    .CE(sig00000001),
    .D(sig000006fb),
    .Q(sig000006f5)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003df (
    .C(clk),
    .CE(sig00000001),
    .D(sig000006fc),
    .Q(sig000006f4)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003e0 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000006fd),
    .Q(sig000006f3)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003e1 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000006fe),
    .Q(sig000006f9)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003e2 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000006ff),
    .Q(sig000006f8)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003e3 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000700),
    .Q(sig000006f7)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003e4 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000701),
    .Q(sig000006f6)
  );
  MUXCY   blk000003e5 (
    .CI(sig00000703),
    .DI(sig000006c3),
    .S(sig000006e2),
    .O(sig00000702)
  );
  MUXCY   blk000003e6 (
    .CI(sig00000704),
    .DI(sig000006c3),
    .S(sig000006e1),
    .O(sig00000703)
  );
  MUXCY   blk000003e7 (
    .CI(sig00000705),
    .DI(sig000006c3),
    .S(sig000006e0),
    .O(sig00000704)
  );
  MUXCY   blk000003e8 (
    .CI(sig00000706),
    .DI(sig000006c3),
    .S(sig000006df),
    .O(sig00000705)
  );
  MUXCY   blk000003e9 (
    .CI(sig00000707),
    .DI(sig000006c3),
    .S(sig000006de),
    .O(sig00000706)
  );
  MUXCY   blk000003ea (
    .CI(sig00000001),
    .DI(sig000006c3),
    .S(sig000006dd),
    .O(sig00000707)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003eb (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000702),
    .Q(sig000006f2)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003ec (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000703),
    .Q(sig000006ed)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003ed (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000704),
    .Q(sig000006f1)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003ee (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000705),
    .Q(sig000006f0)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003ef (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000706),
    .Q(sig000006ef)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003f0 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000707),
    .Q(sig000006ee)
  );
  MUXF7   blk000003f1 (
    .I0(sig00000718),
    .I1(sig00000710),
    .S(sig00000118),
    .O(sig00000708)
  );
  MUXF7   blk000003f2 (
    .I0(sig00000719),
    .I1(sig00000711),
    .S(sig00000118),
    .O(sig00000709)
  );
  MUXF7   blk000003f3 (
    .I0(sig0000071a),
    .I1(sig00000712),
    .S(sig00000118),
    .O(sig0000070a)
  );
  MUXF7   blk000003f4 (
    .I0(sig0000071b),
    .I1(sig00000713),
    .S(sig00000118),
    .O(sig0000070b)
  );
  MUXF7   blk000003f5 (
    .I0(sig0000071c),
    .I1(sig00000714),
    .S(sig00000118),
    .O(sig0000070c)
  );
  MUXF7   blk000003f6 (
    .I0(sig0000071d),
    .I1(sig00000715),
    .S(sig00000118),
    .O(sig0000070d)
  );
  MUXF7   blk000003f7 (
    .I0(sig0000071e),
    .I1(sig00000716),
    .S(sig00000118),
    .O(sig0000070e)
  );
  MUXF7   blk000003f8 (
    .I0(sig0000071f),
    .I1(sig00000717),
    .S(sig00000118),
    .O(sig0000070f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003f9 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000708),
    .Q(sig000006e6)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003fa (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000709),
    .Q(sig000006e5)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003fb (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000070a),
    .Q(sig000006e8)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003fc (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000070b),
    .Q(sig000006e7)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003fd (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000070c),
    .Q(sig000006ea)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003fe (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000070d),
    .Q(sig000006e9)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003ff (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000070e),
    .Q(sig000006ec)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000400 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000070f),
    .Q(sig000006eb)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000401 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000769),
    .Q(sig00000761)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000402 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000076a),
    .Q(sig00000762)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000403 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000076b),
    .Q(sig00000763)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000404 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000076c),
    .Q(sig00000764)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000405 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000076d),
    .Q(sig00000765)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000406 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000076e),
    .Q(sig00000766)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000407 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000076f),
    .Q(sig00000760)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000408 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000720),
    .Q(sig00000768)
  );
  MUXCY   blk00000409 (
    .CI(sig000006c3),
    .DI(sig000006c3),
    .S(sig00000819),
    .O(sig00000721)
  );
  XORCY   blk0000040a (
    .CI(sig000006c3),
    .LI(sig00000819),
    .O(sig00000722)
  );
  MUXCY   blk0000040b (
    .CI(sig00000721),
    .DI(sig000006c3),
    .S(sig0000081a),
    .O(sig00000723)
  );
  XORCY   blk0000040c (
    .CI(sig00000721),
    .LI(sig0000081a),
    .O(sig00000724)
  );
  MUXCY   blk0000040d (
    .CI(sig00000723),
    .DI(sig000006c3),
    .S(sig0000081b),
    .O(sig00000725)
  );
  XORCY   blk0000040e (
    .CI(sig00000723),
    .LI(sig0000081b),
    .O(sig00000726)
  );
  MUXCY   blk0000040f (
    .CI(sig00000725),
    .DI(sig000006c3),
    .S(sig0000081c),
    .O(sig00000727)
  );
  XORCY   blk00000410 (
    .CI(sig00000725),
    .LI(sig0000081c),
    .O(sig00000728)
  );
  MUXCY   blk00000411 (
    .CI(sig00000727),
    .DI(sig000006c3),
    .S(sig0000081d),
    .O(sig00000729)
  );
  XORCY   blk00000412 (
    .CI(sig00000727),
    .LI(sig0000081d),
    .O(sig0000072a)
  );
  MUXCY   blk00000413 (
    .CI(sig00000729),
    .DI(sig000006c3),
    .S(sig0000081e),
    .O(sig0000072b)
  );
  XORCY   blk00000414 (
    .CI(sig00000729),
    .LI(sig0000081e),
    .O(sig0000072c)
  );
  MUXCY   blk00000415 (
    .CI(sig0000072b),
    .DI(sig000006c3),
    .S(sig0000081f),
    .O(sig0000072d)
  );
  XORCY   blk00000416 (
    .CI(sig0000072b),
    .LI(sig0000081f),
    .O(NLW_blk00000416_O_UNCONNECTED)
  );
  MUXCY   blk00000417 (
    .CI(sig0000072d),
    .DI(sig00000001),
    .S(sig00000001),
    .O(sig0000072e)
  );
  XORCY   blk00000418 (
    .CI(sig0000072d),
    .LI(sig00000001),
    .O(NLW_blk00000418_O_UNCONNECTED)
  );
  MUXCY   blk00000419 (
    .CI(sig0000072e),
    .DI(sig000006c3),
    .S(sig000006c3),
    .O(sig0000072f)
  );
  XORCY   blk0000041a (
    .CI(sig0000072e),
    .LI(sig000006c3),
    .O(NLW_blk0000041a_O_UNCONNECTED)
  );
  MUXCY   blk0000041b (
    .CI(sig0000072f),
    .DI(sig000006c3),
    .S(sig000006c3),
    .O(sig00000730)
  );
  XORCY   blk0000041c (
    .CI(sig0000072f),
    .LI(sig000006c3),
    .O(NLW_blk0000041c_O_UNCONNECTED)
  );
  MUXCY   blk0000041d (
    .CI(sig00000730),
    .DI(sig000006c3),
    .S(sig000006c3),
    .O(sig00000731)
  );
  XORCY   blk0000041e (
    .CI(sig00000730),
    .LI(sig000006c3),
    .O(NLW_blk0000041e_O_UNCONNECTED)
  );
  MUXCY   blk0000041f (
    .CI(sig00000731),
    .DI(sig000006c3),
    .S(sig000006c3),
    .O(sig00000732)
  );
  XORCY   blk00000420 (
    .CI(sig00000731),
    .LI(sig000006c3),
    .O(NLW_blk00000420_O_UNCONNECTED)
  );
  MUXCY   blk00000421 (
    .CI(sig00000732),
    .DI(sig000006c3),
    .S(sig000006c3),
    .O(sig00000733)
  );
  XORCY   blk00000422 (
    .CI(sig00000732),
    .LI(sig000006c3),
    .O(NLW_blk00000422_O_UNCONNECTED)
  );
  MUXCY   blk00000423 (
    .CI(sig00000733),
    .DI(sig000006c3),
    .S(sig000006c3),
    .O(sig00000734)
  );
  XORCY   blk00000424 (
    .CI(sig00000733),
    .LI(sig000006c3),
    .O(NLW_blk00000424_O_UNCONNECTED)
  );
  MUXCY   blk00000425 (
    .CI(sig00000734),
    .DI(sig000006c3),
    .S(sig000006c3),
    .O(sig00000735)
  );
  XORCY   blk00000426 (
    .CI(sig00000734),
    .LI(sig000006c3),
    .O(NLW_blk00000426_O_UNCONNECTED)
  );
  MUXCY   blk00000427 (
    .CI(sig00000735),
    .DI(sig000006c3),
    .S(sig000006c3),
    .O(sig00000736)
  );
  XORCY   blk00000428 (
    .CI(sig00000735),
    .LI(sig000006c3),
    .O(NLW_blk00000428_O_UNCONNECTED)
  );
  MUXCY   blk00000429 (
    .CI(sig00000736),
    .DI(sig000006c3),
    .S(sig000006c3),
    .O(sig00000737)
  );
  XORCY   blk0000042a (
    .CI(sig00000736),
    .LI(sig000006c3),
    .O(NLW_blk0000042a_O_UNCONNECTED)
  );
  MUXCY   blk0000042b (
    .CI(sig00000737),
    .DI(sig000006c3),
    .S(sig000006c3),
    .O(sig00000738)
  );
  XORCY   blk0000042c (
    .CI(sig00000737),
    .LI(sig000006c3),
    .O(NLW_blk0000042c_O_UNCONNECTED)
  );
  XORCY   blk0000042d (
    .CI(sig00000738),
    .LI(sig000006c3),
    .O(NLW_blk0000042d_O_UNCONNECTED)
  );
  MUXCY   blk0000042e (
    .CI(sig00000001),
    .DI(sig000006c3),
    .S(sig00000820),
    .O(sig00000739)
  );
  XORCY   blk0000042f (
    .CI(sig00000001),
    .LI(sig00000820),
    .O(sig0000073a)
  );
  MUXCY   blk00000430 (
    .CI(sig00000739),
    .DI(sig000006c3),
    .S(sig00000821),
    .O(sig0000073b)
  );
  XORCY   blk00000431 (
    .CI(sig00000739),
    .LI(sig00000821),
    .O(sig0000073c)
  );
  MUXCY   blk00000432 (
    .CI(sig0000073b),
    .DI(sig000006c3),
    .S(sig00000822),
    .O(sig0000073d)
  );
  XORCY   blk00000433 (
    .CI(sig0000073b),
    .LI(sig00000822),
    .O(sig0000073e)
  );
  MUXCY   blk00000434 (
    .CI(sig0000073d),
    .DI(sig000006c3),
    .S(sig00000823),
    .O(sig0000073f)
  );
  XORCY   blk00000435 (
    .CI(sig0000073d),
    .LI(sig00000823),
    .O(sig00000740)
  );
  MUXCY   blk00000436 (
    .CI(sig0000073f),
    .DI(sig000006c3),
    .S(sig00000824),
    .O(sig00000741)
  );
  XORCY   blk00000437 (
    .CI(sig0000073f),
    .LI(sig00000824),
    .O(sig00000742)
  );
  MUXCY   blk00000438 (
    .CI(sig00000741),
    .DI(sig000006c3),
    .S(sig00000825),
    .O(sig00000743)
  );
  XORCY   blk00000439 (
    .CI(sig00000741),
    .LI(sig00000825),
    .O(sig00000744)
  );
  MUXCY   blk0000043a (
    .CI(sig00000743),
    .DI(sig000006c3),
    .S(sig00000826),
    .O(sig00000745)
  );
  XORCY   blk0000043b (
    .CI(sig00000743),
    .LI(sig00000826),
    .O(NLW_blk0000043b_O_UNCONNECTED)
  );
  MUXCY   blk0000043c (
    .CI(sig00000745),
    .DI(sig00000001),
    .S(sig00000001),
    .O(sig00000746)
  );
  XORCY   blk0000043d (
    .CI(sig00000745),
    .LI(sig00000001),
    .O(sig00000747)
  );
  MUXCY   blk0000043e (
    .CI(sig00000746),
    .DI(sig000006c3),
    .S(sig000006c3),
    .O(sig00000748)
  );
  XORCY   blk0000043f (
    .CI(sig00000746),
    .LI(sig000006c3),
    .O(NLW_blk0000043f_O_UNCONNECTED)
  );
  MUXCY   blk00000440 (
    .CI(sig00000748),
    .DI(sig000006c3),
    .S(sig000006c3),
    .O(sig00000749)
  );
  XORCY   blk00000441 (
    .CI(sig00000748),
    .LI(sig000006c3),
    .O(NLW_blk00000441_O_UNCONNECTED)
  );
  MUXCY   blk00000442 (
    .CI(sig00000749),
    .DI(sig000006c3),
    .S(sig000006c3),
    .O(sig0000074a)
  );
  XORCY   blk00000443 (
    .CI(sig00000749),
    .LI(sig000006c3),
    .O(NLW_blk00000443_O_UNCONNECTED)
  );
  MUXCY   blk00000444 (
    .CI(sig0000074a),
    .DI(sig000006c3),
    .S(sig000006c3),
    .O(sig0000074b)
  );
  XORCY   blk00000445 (
    .CI(sig0000074a),
    .LI(sig000006c3),
    .O(NLW_blk00000445_O_UNCONNECTED)
  );
  MUXCY   blk00000446 (
    .CI(sig0000074b),
    .DI(sig000006c3),
    .S(sig000006c3),
    .O(sig0000074c)
  );
  XORCY   blk00000447 (
    .CI(sig0000074b),
    .LI(sig000006c3),
    .O(NLW_blk00000447_O_UNCONNECTED)
  );
  MUXCY   blk00000448 (
    .CI(sig0000074c),
    .DI(sig000006c3),
    .S(sig000006c3),
    .O(sig0000074d)
  );
  XORCY   blk00000449 (
    .CI(sig0000074c),
    .LI(sig000006c3),
    .O(NLW_blk00000449_O_UNCONNECTED)
  );
  MUXCY   blk0000044a (
    .CI(sig0000074d),
    .DI(sig000006c3),
    .S(sig000006c3),
    .O(sig0000074e)
  );
  XORCY   blk0000044b (
    .CI(sig0000074d),
    .LI(sig000006c3),
    .O(NLW_blk0000044b_O_UNCONNECTED)
  );
  MUXCY   blk0000044c (
    .CI(sig0000074e),
    .DI(sig000006c3),
    .S(sig000006c3),
    .O(sig0000074f)
  );
  XORCY   blk0000044d (
    .CI(sig0000074e),
    .LI(sig000006c3),
    .O(NLW_blk0000044d_O_UNCONNECTED)
  );
  MUXCY   blk0000044e (
    .CI(sig0000074f),
    .DI(sig000006c3),
    .S(sig000006c3),
    .O(sig00000750)
  );
  XORCY   blk0000044f (
    .CI(sig0000074f),
    .LI(sig000006c3),
    .O(NLW_blk0000044f_O_UNCONNECTED)
  );
  MUXCY   blk00000450 (
    .CI(sig00000750),
    .DI(sig000006c3),
    .S(sig000006c3),
    .O(sig00000751)
  );
  XORCY   blk00000451 (
    .CI(sig00000750),
    .LI(sig000006c3),
    .O(NLW_blk00000451_O_UNCONNECTED)
  );
  XORCY   blk00000452 (
    .CI(sig00000751),
    .LI(sig000006c3),
    .O(NLW_blk00000452_O_UNCONNECTED)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000453 (
    .C(clk),
    .D(sig00000117),
    .Q(sig0000076f)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000454 (
    .C(clk),
    .D(sig00000116),
    .Q(sig0000076e)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000455 (
    .C(clk),
    .D(sig00000115),
    .Q(sig0000076d)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000456 (
    .C(clk),
    .D(sig00000114),
    .Q(sig0000076c)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000457 (
    .C(clk),
    .D(sig00000113),
    .Q(sig0000076b)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000458 (
    .C(clk),
    .D(sig00000112),
    .Q(sig0000076a)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000459 (
    .C(clk),
    .D(sig00000111),
    .Q(sig00000769)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000045a (
    .C(clk),
    .D(sig00000110),
    .Q(sig00000752)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000045b (
    .C(clk),
    .D(sig0000010f),
    .Q(sig0000079d)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000045c (
    .C(clk),
    .D(sig0000010e),
    .Q(sig0000079c)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000045d (
    .C(clk),
    .D(sig0000010d),
    .Q(sig0000079b)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000045e (
    .C(clk),
    .D(sig0000010c),
    .Q(sig0000079a)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000045f (
    .C(clk),
    .D(sig0000010b),
    .Q(sig00000799)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000460 (
    .C(clk),
    .D(sig0000010a),
    .Q(sig00000798)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000461 (
    .C(clk),
    .D(sig00000109),
    .Q(sig00000797)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000462 (
    .C(clk),
    .D(sig00000108),
    .Q(sig00000796)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000463 (
    .C(clk),
    .D(sig00000107),
    .Q(sig00000795)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000464 (
    .C(clk),
    .D(sig00000106),
    .Q(sig00000794)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000465 (
    .C(clk),
    .D(sig00000105),
    .Q(sig00000793)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000466 (
    .C(clk),
    .D(sig00000104),
    .Q(sig00000792)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000467 (
    .C(clk),
    .D(sig00000103),
    .Q(sig00000791)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000468 (
    .C(clk),
    .D(sig00000102),
    .Q(sig00000790)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000469 (
    .C(clk),
    .D(sig00000101),
    .Q(sig0000078f)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000046a (
    .C(clk),
    .D(sig00000100),
    .Q(sig0000078e)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000046b (
    .C(clk),
    .D(sig000000ff),
    .Q(sig0000078d)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000046c (
    .C(clk),
    .D(sig000000fe),
    .Q(sig0000078c)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000046d (
    .C(clk),
    .D(sig000000fd),
    .Q(sig0000078b)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000046e (
    .C(clk),
    .D(sig000000fc),
    .Q(sig0000078a)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000046f (
    .C(clk),
    .D(sig000000fb),
    .Q(sig00000789)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000470 (
    .C(clk),
    .D(sig000000fa),
    .Q(sig00000788)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000471 (
    .C(clk),
    .D(sig000000f9),
    .Q(sig00000787)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000472 (
    .C(clk),
    .D(sig000000f8),
    .Q(sig00000786)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000473 (
    .C(clk),
    .D(sig000000f7),
    .Q(sig00000785)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000474 (
    .C(clk),
    .D(sig000000f6),
    .Q(sig00000784)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000475 (
    .C(clk),
    .D(sig000000f5),
    .Q(sig00000783)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000476 (
    .C(clk),
    .D(sig000000f4),
    .Q(sig00000782)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000477 (
    .C(clk),
    .D(sig000000f3),
    .Q(sig00000781)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000478 (
    .C(clk),
    .D(sig000000f2),
    .Q(sig00000780)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000479 (
    .C(clk),
    .D(sig000000f1),
    .Q(sig0000077f)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000047a (
    .C(clk),
    .D(sig000000f0),
    .Q(sig0000077e)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000047b (
    .C(clk),
    .D(sig000000ef),
    .Q(sig0000077d)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000047c (
    .C(clk),
    .D(sig000000ee),
    .Q(sig0000077c)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000047d (
    .C(clk),
    .D(sig000000ed),
    .Q(sig0000077b)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000047e (
    .C(clk),
    .D(sig000000ec),
    .Q(sig0000077a)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000047f (
    .C(clk),
    .D(sig000000eb),
    .Q(sig00000779)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000480 (
    .C(clk),
    .D(sig000000ea),
    .Q(sig00000778)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000481 (
    .C(clk),
    .D(sig000000e9),
    .Q(sig00000777)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000482 (
    .C(clk),
    .D(sig000000e8),
    .Q(sig00000776)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000483 (
    .C(clk),
    .D(sig000000e7),
    .Q(sig00000775)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000484 (
    .C(clk),
    .D(sig000000e6),
    .Q(sig00000774)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000485 (
    .C(clk),
    .D(sig000000e5),
    .Q(sig00000773)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000486 (
    .C(clk),
    .D(sig000000e4),
    .Q(sig00000772)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000487 (
    .C(clk),
    .D(sig000000e3),
    .Q(sig00000771)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000488 (
    .C(clk),
    .D(sig000000e2),
    .Q(sig00000770)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000489 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000072c),
    .Q(sig0000075f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000048a (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000072a),
    .Q(sig0000075e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000048b (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000728),
    .Q(sig0000075d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000048c (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000726),
    .Q(sig0000075c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000048d (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000724),
    .Q(sig0000075b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000048e (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000722),
    .Q(sig0000075a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000048f (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000747),
    .Q(sig00000759)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000490 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000744),
    .Q(sig00000758)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000491 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000742),
    .Q(sig00000757)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000492 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000740),
    .Q(sig00000756)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000493 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000073e),
    .Q(sig00000755)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000494 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000073c),
    .Q(sig00000754)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000495 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000073a),
    .Q(sig00000753)
  );
  XORCY   blk00000496 (
    .CI(sig0000079e),
    .LI(sig000007f2),
    .O(sig000007b3)
  );
  XORCY   blk00000497 (
    .CI(sig0000079f),
    .LI(sig000007f1),
    .O(sig000007b2)
  );
  MUXCY   blk00000498 (
    .CI(sig0000079f),
    .DI(sig000006c3),
    .S(sig000007f1),
    .O(sig0000079e)
  );
  XORCY   blk00000499 (
    .CI(sig000007a0),
    .LI(sig000007f0),
    .O(sig000007b1)
  );
  MUXCY   blk0000049a (
    .CI(sig000007a0),
    .DI(sig000006c3),
    .S(sig000007f0),
    .O(sig0000079f)
  );
  XORCY   blk0000049b (
    .CI(sig000007a1),
    .LI(sig000007ef),
    .O(sig000007b0)
  );
  MUXCY   blk0000049c (
    .CI(sig000007a1),
    .DI(sig000006c3),
    .S(sig000007ef),
    .O(sig000007a0)
  );
  XORCY   blk0000049d (
    .CI(sig000007a2),
    .LI(sig000007ee),
    .O(sig000007af)
  );
  MUXCY   blk0000049e (
    .CI(sig000007a2),
    .DI(sig000006c3),
    .S(sig000007ee),
    .O(sig000007a1)
  );
  XORCY   blk0000049f (
    .CI(sig000007a3),
    .LI(sig000007ed),
    .O(sig000007ae)
  );
  MUXCY   blk000004a0 (
    .CI(sig000007a3),
    .DI(sig000006c3),
    .S(sig000007ed),
    .O(sig000007a2)
  );
  XORCY   blk000004a1 (
    .CI(sig000007a4),
    .LI(sig000007ec),
    .O(sig000007ad)
  );
  MUXCY   blk000004a2 (
    .CI(sig000007a4),
    .DI(sig000006c3),
    .S(sig000007ec),
    .O(sig000007a3)
  );
  XORCY   blk000004a3 (
    .CI(sig000007a5),
    .LI(sig000007eb),
    .O(sig000007ac)
  );
  MUXCY   blk000004a4 (
    .CI(sig000007a5),
    .DI(sig000006c3),
    .S(sig000007eb),
    .O(sig000007a4)
  );
  XORCY   blk000004a5 (
    .CI(sig000007a6),
    .LI(sig000007ea),
    .O(sig000007ab)
  );
  MUXCY   blk000004a6 (
    .CI(sig000007a6),
    .DI(sig000006c3),
    .S(sig000007ea),
    .O(sig000007a5)
  );
  XORCY   blk000004a7 (
    .CI(sig000007a7),
    .LI(sig000007e9),
    .O(sig000007aa)
  );
  MUXCY   blk000004a8 (
    .CI(sig000007a7),
    .DI(sig000006c3),
    .S(sig000007e9),
    .O(sig000007a6)
  );
  XORCY   blk000004a9 (
    .CI(sig000006c3),
    .LI(sig000007a8),
    .O(sig000007a9)
  );
  MUXCY   blk000004aa (
    .CI(sig000006c3),
    .DI(sig000007e8),
    .S(sig000007a8),
    .O(sig000007a7)
  );
  FD   blk000004ab (
    .C(clk),
    .D(sig000007b3),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/exp_op [10])
  );
  FD   blk000004ac (
    .C(clk),
    .D(sig000007b2),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/exp_op [9])
  );
  FD   blk000004ad (
    .C(clk),
    .D(sig000007b1),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/exp_op [8])
  );
  FD   blk000004ae (
    .C(clk),
    .D(sig000007b0),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/exp_op [7])
  );
  FD   blk000004af (
    .C(clk),
    .D(sig000007af),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/exp_op [6])
  );
  FD   blk000004b0 (
    .C(clk),
    .D(sig000007ae),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/exp_op [5])
  );
  FD   blk000004b1 (
    .C(clk),
    .D(sig000007ad),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/exp_op [4])
  );
  FD   blk000004b2 (
    .C(clk),
    .D(sig000007ac),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/exp_op [3])
  );
  FD   blk000004b3 (
    .C(clk),
    .D(sig000007ab),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/exp_op [2])
  );
  FD   blk000004b4 (
    .C(clk),
    .D(sig000007aa),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/exp_op [1])
  );
  FD   blk000004b5 (
    .C(clk),
    .D(sig000007a9),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/exp_op [0])
  );
  FD   blk000004b6 (
    .C(clk),
    .D(sig000007e7),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [51])
  );
  FD   blk000004b7 (
    .C(clk),
    .D(sig000007e6),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [50])
  );
  FD   blk000004b8 (
    .C(clk),
    .D(sig000007e5),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [49])
  );
  FD   blk000004b9 (
    .C(clk),
    .D(sig000007e4),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [48])
  );
  FD   blk000004ba (
    .C(clk),
    .D(sig000007e3),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [47])
  );
  FD   blk000004bb (
    .C(clk),
    .D(sig000007e2),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [46])
  );
  FD   blk000004bc (
    .C(clk),
    .D(sig000007e1),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [45])
  );
  FD   blk000004bd (
    .C(clk),
    .D(sig000007e0),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [44])
  );
  FD   blk000004be (
    .C(clk),
    .D(sig000007df),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [43])
  );
  FD   blk000004bf (
    .C(clk),
    .D(sig000007de),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [42])
  );
  FD   blk000004c0 (
    .C(clk),
    .D(sig000007dd),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [41])
  );
  FD   blk000004c1 (
    .C(clk),
    .D(sig000007dc),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [40])
  );
  FD   blk000004c2 (
    .C(clk),
    .D(sig000007db),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [39])
  );
  FD   blk000004c3 (
    .C(clk),
    .D(sig000007da),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [38])
  );
  FD   blk000004c4 (
    .C(clk),
    .D(sig000007d9),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [37])
  );
  FD   blk000004c5 (
    .C(clk),
    .D(sig000007d8),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [36])
  );
  FD   blk000004c6 (
    .C(clk),
    .D(sig000007d7),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [35])
  );
  FD   blk000004c7 (
    .C(clk),
    .D(sig000007d6),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [34])
  );
  FD   blk000004c8 (
    .C(clk),
    .D(sig000007d5),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [33])
  );
  FD   blk000004c9 (
    .C(clk),
    .D(sig000007d4),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [32])
  );
  FD   blk000004ca (
    .C(clk),
    .D(sig000007d3),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [31])
  );
  FD   blk000004cb (
    .C(clk),
    .D(sig000007d2),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [30])
  );
  FD   blk000004cc (
    .C(clk),
    .D(sig000007d1),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [29])
  );
  FD   blk000004cd (
    .C(clk),
    .D(sig000007d0),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [28])
  );
  FD   blk000004ce (
    .C(clk),
    .D(sig000007cf),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [27])
  );
  FD   blk000004cf (
    .C(clk),
    .D(sig000007ce),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [26])
  );
  FD   blk000004d0 (
    .C(clk),
    .D(sig000007cd),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [25])
  );
  FD   blk000004d1 (
    .C(clk),
    .D(sig000007cc),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [24])
  );
  FD   blk000004d2 (
    .C(clk),
    .D(sig000007cb),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [23])
  );
  FD   blk000004d3 (
    .C(clk),
    .D(sig000007ca),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [22])
  );
  FD   blk000004d4 (
    .C(clk),
    .D(sig000007c9),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [21])
  );
  FD   blk000004d5 (
    .C(clk),
    .D(sig000007c8),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [20])
  );
  FD   blk000004d6 (
    .C(clk),
    .D(sig000007c7),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [19])
  );
  FD   blk000004d7 (
    .C(clk),
    .D(sig000007c6),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [18])
  );
  FD   blk000004d8 (
    .C(clk),
    .D(sig000007c5),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [17])
  );
  FD   blk000004d9 (
    .C(clk),
    .D(sig000007c4),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [16])
  );
  FD   blk000004da (
    .C(clk),
    .D(sig000007c3),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [15])
  );
  FD   blk000004db (
    .C(clk),
    .D(sig000007c2),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [14])
  );
  FD   blk000004dc (
    .C(clk),
    .D(sig000007c1),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [13])
  );
  FD   blk000004dd (
    .C(clk),
    .D(sig000007c0),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [12])
  );
  FD   blk000004de (
    .C(clk),
    .D(sig000007bf),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [11])
  );
  FD   blk000004df (
    .C(clk),
    .D(sig000007be),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [10])
  );
  FD   blk000004e0 (
    .C(clk),
    .D(sig000007bd),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [9])
  );
  FD   blk000004e1 (
    .C(clk),
    .D(sig000007bc),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [8])
  );
  FD   blk000004e2 (
    .C(clk),
    .D(sig000007bb),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [7])
  );
  FD   blk000004e3 (
    .C(clk),
    .D(sig000007ba),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [6])
  );
  FD   blk000004e4 (
    .C(clk),
    .D(sig000007b9),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [5])
  );
  FD   blk000004e5 (
    .C(clk),
    .D(sig000007b8),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [4])
  );
  FD   blk000004e6 (
    .C(clk),
    .D(sig000007b7),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [3])
  );
  FD   blk000004e7 (
    .C(clk),
    .D(sig000007b6),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [2])
  );
  FD   blk000004e8 (
    .C(clk),
    .D(sig000007b5),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [1])
  );
  FD   blk000004e9 (
    .C(clk),
    .D(sig000007b4),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/mant_op [0])
  );
  LUT6 #(
    .INIT ( 64'hFF00CCCCF0F0AAAA ))
  blk000004ea (
    .I0(sig00000124),
    .I1(sig00000134),
    .I2(sig00000144),
    .I3(sig00000154),
    .I4(sig00000118),
    .I5(sig00000119),
    .O(sig000000a2)
  );
  LUT6 #(
    .INIT ( 64'hFF00CCCCF0F0AAAA ))
  blk000004eb (
    .I0(sig00000123),
    .I1(sig00000133),
    .I2(sig00000143),
    .I3(sig00000153),
    .I4(sig00000118),
    .I5(sig00000119),
    .O(sig000000a3)
  );
  LUT6 #(
    .INIT ( 64'hFF00CCCCF0F0AAAA ))
  blk000004ec (
    .I0(sig0000027f),
    .I1(sig0000012d),
    .I2(sig0000013d),
    .I3(sig0000014d),
    .I4(sig00000118),
    .I5(sig00000119),
    .O(sig000000a9)
  );
  LUT6 #(
    .INIT ( 64'hFF00CCCCF0F0AAAA ))
  blk000004ed (
    .I0(sig00000122),
    .I1(sig00000132),
    .I2(sig00000142),
    .I3(sig00000152),
    .I4(sig00000118),
    .I5(sig00000119),
    .O(sig000000a4)
  );
  LUT6 #(
    .INIT ( 64'hFF00CCCCF0F0AAAA ))
  blk000004ee (
    .I0(sig00000121),
    .I1(sig00000131),
    .I2(sig00000141),
    .I3(sig00000151),
    .I4(sig00000118),
    .I5(sig00000119),
    .O(sig000000a5)
  );
  LUT6 #(
    .INIT ( 64'hFF00CCCCF0F0AAAA ))
  blk000004ef (
    .I0(sig00000120),
    .I1(sig00000130),
    .I2(sig00000140),
    .I3(sig00000150),
    .I4(sig00000118),
    .I5(sig00000119),
    .O(sig000000a6)
  );
  LUT6 #(
    .INIT ( 64'hFF00CCCCF0F0AAAA ))
  blk000004f0 (
    .I0(sig0000011f),
    .I1(sig0000012f),
    .I2(sig0000013f),
    .I3(sig0000014f),
    .I4(sig00000118),
    .I5(sig00000119),
    .O(sig000000a7)
  );
  LUT6 #(
    .INIT ( 64'hFF00CCCCF0F0AAAA ))
  blk000004f1 (
    .I0(sig0000011e),
    .I1(sig0000012e),
    .I2(sig0000013e),
    .I3(sig0000014e),
    .I4(sig00000118),
    .I5(sig00000119),
    .O(sig000000a8)
  );
  LUT6 #(
    .INIT ( 64'hF0F0FF00CCCCAAAA ))
  blk000004f2 (
    .I0(sig0000000e),
    .I1(sig00000006),
    .I2(sig00000002),
    .I3(sig0000000a),
    .I4(sig0000011a),
    .I5(sig0000011b),
    .O(sig000000b6)
  );
  LUT6 #(
    .INIT ( 64'hF0F0FF00CCCCAAAA ))
  blk000004f3 (
    .I0(sig0000000f),
    .I1(sig00000007),
    .I2(sig00000003),
    .I3(sig0000000b),
    .I4(sig0000011a),
    .I5(sig0000011b),
    .O(sig000000b7)
  );
  LUT6 #(
    .INIT ( 64'hF0F0FF00CCCCAAAA ))
  blk000004f4 (
    .I0(sig00000010),
    .I1(sig00000008),
    .I2(sig00000004),
    .I3(sig0000000c),
    .I4(sig0000011a),
    .I5(sig0000011b),
    .O(sig000000b8)
  );
  LUT6 #(
    .INIT ( 64'hF0F0FF00CCCCAAAA ))
  blk000004f5 (
    .I0(sig00000011),
    .I1(sig00000009),
    .I2(sig00000005),
    .I3(sig0000000d),
    .I4(sig0000011a),
    .I5(sig0000011b),
    .O(sig000000b9)
  );
  LUT6 #(
    .INIT ( 64'hF0F0FF00CCCCAAAA ))
  blk000004f6 (
    .I0(sig00000012),
    .I1(sig0000000a),
    .I2(sig00000006),
    .I3(sig0000000e),
    .I4(sig0000011a),
    .I5(sig0000011b),
    .O(sig000000ba)
  );
  LUT6 #(
    .INIT ( 64'hF0F0FF00CCCCAAAA ))
  blk000004f7 (
    .I0(sig00000016),
    .I1(sig0000000e),
    .I2(sig0000000a),
    .I3(sig00000012),
    .I4(sig0000011a),
    .I5(sig0000011b),
    .O(sig000000be)
  );
  LUT6 #(
    .INIT ( 64'hF0F0FF00CCCCAAAA ))
  blk000004f8 (
    .I0(sig00000017),
    .I1(sig0000000f),
    .I2(sig0000000b),
    .I3(sig00000013),
    .I4(sig0000011a),
    .I5(sig0000011b),
    .O(sig000000bf)
  );
  LUT6 #(
    .INIT ( 64'hF0F0FF00CCCCAAAA ))
  blk000004f9 (
    .I0(sig00000018),
    .I1(sig00000010),
    .I2(sig0000000c),
    .I3(sig00000014),
    .I4(sig0000011a),
    .I5(sig0000011b),
    .O(sig000000c0)
  );
  LUT6 #(
    .INIT ( 64'hF0F0FF00CCCCAAAA ))
  blk000004fa (
    .I0(sig00000019),
    .I1(sig00000011),
    .I2(sig0000000d),
    .I3(sig00000015),
    .I4(sig0000011a),
    .I5(sig0000011b),
    .O(sig000000c1)
  );
  LUT6 #(
    .INIT ( 64'hF0F0FF00CCCCAAAA ))
  blk000004fb (
    .I0(sig0000001a),
    .I1(sig00000012),
    .I2(sig0000000e),
    .I3(sig00000016),
    .I4(sig0000011a),
    .I5(sig0000011b),
    .O(sig000000c2)
  );
  LUT6 #(
    .INIT ( 64'hF0F0FF00CCCCAAAA ))
  blk000004fc (
    .I0(sig0000001f),
    .I1(sig00000017),
    .I2(sig00000013),
    .I3(sig0000001b),
    .I4(sig0000011a),
    .I5(sig0000011b),
    .O(sig000000c7)
  );
  LUT6 #(
    .INIT ( 64'hF0F0FF00CCCCAAAA ))
  blk000004fd (
    .I0(sig00000020),
    .I1(sig00000018),
    .I2(sig00000014),
    .I3(sig0000001c),
    .I4(sig0000011a),
    .I5(sig0000011b),
    .O(sig000000c8)
  );
  LUT6 #(
    .INIT ( 64'hF0F0FF00CCCCAAAA ))
  blk000004fe (
    .I0(sig00000021),
    .I1(sig00000019),
    .I2(sig00000015),
    .I3(sig0000001d),
    .I4(sig0000011a),
    .I5(sig0000011b),
    .O(sig000000c9)
  );
  LUT6 #(
    .INIT ( 64'hF0F0FF00CCCCAAAA ))
  blk000004ff (
    .I0(sig00000013),
    .I1(sig0000000b),
    .I2(sig00000007),
    .I3(sig0000000f),
    .I4(sig0000011a),
    .I5(sig0000011b),
    .O(sig000000bb)
  );
  LUT6 #(
    .INIT ( 64'hF0F0FF00CCCCAAAA ))
  blk00000500 (
    .I0(sig00000022),
    .I1(sig0000001a),
    .I2(sig00000016),
    .I3(sig0000001e),
    .I4(sig0000011a),
    .I5(sig0000011b),
    .O(sig000000ca)
  );
  LUT6 #(
    .INIT ( 64'hF0F0FF00CCCCAAAA ))
  blk00000501 (
    .I0(sig0000001b),
    .I1(sig00000013),
    .I2(sig0000000f),
    .I3(sig00000017),
    .I4(sig0000011a),
    .I5(sig0000011b),
    .O(sig000000c3)
  );
  LUT6 #(
    .INIT ( 64'hF0F0FF00CCCCAAAA ))
  blk00000502 (
    .I0(sig00000023),
    .I1(sig0000001b),
    .I2(sig00000017),
    .I3(sig0000001f),
    .I4(sig0000011a),
    .I5(sig0000011b),
    .O(sig000000cb)
  );
  LUT6 #(
    .INIT ( 64'hF0F0FF00CCCCAAAA ))
  blk00000503 (
    .I0(sig00000024),
    .I1(sig0000001c),
    .I2(sig00000018),
    .I3(sig00000020),
    .I4(sig0000011a),
    .I5(sig0000011b),
    .O(sig000000cc)
  );
  LUT6 #(
    .INIT ( 64'hF0F0FF00CCCCAAAA ))
  blk00000504 (
    .I0(sig0000001c),
    .I1(sig00000014),
    .I2(sig00000010),
    .I3(sig00000018),
    .I4(sig0000011a),
    .I5(sig0000011b),
    .O(sig000000c4)
  );
  LUT6 #(
    .INIT ( 64'hF0F0FF00CCCCAAAA ))
  blk00000505 (
    .I0(sig00000025),
    .I1(sig0000001d),
    .I2(sig00000019),
    .I3(sig00000021),
    .I4(sig0000011a),
    .I5(sig0000011b),
    .O(sig000000cd)
  );
  LUT6 #(
    .INIT ( 64'hF0F0FF00CCCCAAAA ))
  blk00000506 (
    .I0(sig0000001d),
    .I1(sig00000015),
    .I2(sig00000011),
    .I3(sig00000019),
    .I4(sig0000011a),
    .I5(sig0000011b),
    .O(sig000000c5)
  );
  LUT6 #(
    .INIT ( 64'hF0F0FF00CCCCAAAA ))
  blk00000507 (
    .I0(sig00000026),
    .I1(sig0000001e),
    .I2(sig0000001a),
    .I3(sig00000022),
    .I4(sig0000011a),
    .I5(sig0000011b),
    .O(sig000000ce)
  );
  LUT6 #(
    .INIT ( 64'hF0F0FF00CCCCAAAA ))
  blk00000508 (
    .I0(sig0000001e),
    .I1(sig00000016),
    .I2(sig00000012),
    .I3(sig0000001a),
    .I4(sig0000011a),
    .I5(sig0000011b),
    .O(sig000000c6)
  );
  LUT6 #(
    .INIT ( 64'hF0F0FF00CCCCAAAA ))
  blk00000509 (
    .I0(sig00000027),
    .I1(sig0000001f),
    .I2(sig0000001b),
    .I3(sig00000023),
    .I4(sig0000011a),
    .I5(sig0000011b),
    .O(sig000000cf)
  );
  LUT6 #(
    .INIT ( 64'hF0F0FF00CCCCAAAA ))
  blk0000050a (
    .I0(sig00000028),
    .I1(sig00000020),
    .I2(sig0000001c),
    .I3(sig00000024),
    .I4(sig0000011a),
    .I5(sig0000011b),
    .O(sig000000d0)
  );
  LUT6 #(
    .INIT ( 64'hF0F0FF00CCCCAAAA ))
  blk0000050b (
    .I0(sig00000029),
    .I1(sig00000021),
    .I2(sig0000001d),
    .I3(sig00000025),
    .I4(sig0000011a),
    .I5(sig0000011b),
    .O(sig000000d1)
  );
  LUT6 #(
    .INIT ( 64'hF0F0FF00CCCCAAAA ))
  blk0000050c (
    .I0(sig0000002a),
    .I1(sig00000022),
    .I2(sig0000001e),
    .I3(sig00000026),
    .I4(sig0000011a),
    .I5(sig0000011b),
    .O(sig000000d2)
  );
  LUT6 #(
    .INIT ( 64'hF0F0FF00CCCCAAAA ))
  blk0000050d (
    .I0(sig00000014),
    .I1(sig0000000c),
    .I2(sig00000008),
    .I3(sig00000010),
    .I4(sig0000011a),
    .I5(sig0000011b),
    .O(sig000000bc)
  );
  LUT6 #(
    .INIT ( 64'hF0F0FF00CCCCAAAA ))
  blk0000050e (
    .I0(sig0000002b),
    .I1(sig00000023),
    .I2(sig0000001f),
    .I3(sig00000027),
    .I4(sig0000011a),
    .I5(sig0000011b),
    .O(sig000000d3)
  );
  LUT6 #(
    .INIT ( 64'hF0F0FF00CCCCAAAA ))
  blk0000050f (
    .I0(sig0000002c),
    .I1(sig00000024),
    .I2(sig00000020),
    .I3(sig00000028),
    .I4(sig0000011a),
    .I5(sig0000011b),
    .O(sig000000d4)
  );
  LUT6 #(
    .INIT ( 64'hF0F0FF00CCCCAAAA ))
  blk00000510 (
    .I0(sig0000002d),
    .I1(sig00000025),
    .I2(sig00000021),
    .I3(sig00000029),
    .I4(sig0000011a),
    .I5(sig0000011b),
    .O(sig000000d5)
  );
  LUT6 #(
    .INIT ( 64'hF0F0FF00CCCCAAAA ))
  blk00000511 (
    .I0(sig0000002e),
    .I1(sig00000026),
    .I2(sig00000022),
    .I3(sig0000002a),
    .I4(sig0000011a),
    .I5(sig0000011b),
    .O(sig000000d6)
  );
  LUT6 #(
    .INIT ( 64'hF0F0FF00CCCCAAAA ))
  blk00000512 (
    .I0(sig0000002f),
    .I1(sig00000027),
    .I2(sig00000023),
    .I3(sig0000002b),
    .I4(sig0000011a),
    .I5(sig0000011b),
    .O(sig000000d7)
  );
  LUT6 #(
    .INIT ( 64'hF0F0FF00CCCCAAAA ))
  blk00000513 (
    .I0(sig00000030),
    .I1(sig00000028),
    .I2(sig00000024),
    .I3(sig0000002c),
    .I4(sig0000011a),
    .I5(sig0000011b),
    .O(sig000000d8)
  );
  LUT6 #(
    .INIT ( 64'hFF00CCCCF0F0AAAA ))
  blk00000514 (
    .I0(sig00000038),
    .I1(sig00000034),
    .I2(sig00000030),
    .I3(sig0000002c),
    .I4(sig0000011a),
    .I5(sig0000011b),
    .O(sig000000e0)
  );
  LUT6 #(
    .INIT ( 64'hF0F0FF00CCCCAAAA ))
  blk00000515 (
    .I0(sig00000031),
    .I1(sig00000029),
    .I2(sig00000025),
    .I3(sig0000002d),
    .I4(sig0000011a),
    .I5(sig0000011b),
    .O(sig000000d9)
  );
  LUT6 #(
    .INIT ( 64'hFF00CCCCF0F0AAAA ))
  blk00000516 (
    .I0(sig00000032),
    .I1(sig0000002e),
    .I2(sig0000002a),
    .I3(sig00000026),
    .I4(sig0000011a),
    .I5(sig0000011b),
    .O(sig000000da)
  );
  LUT6 #(
    .INIT ( 64'hFF00CCCCF0F0AAAA ))
  blk00000517 (
    .I0(sig00000039),
    .I1(sig00000035),
    .I2(sig00000031),
    .I3(sig0000002d),
    .I4(sig0000011a),
    .I5(sig0000011b),
    .O(sig000000e1)
  );
  LUT6 #(
    .INIT ( 64'hF0F0FF00CCCCAAAA ))
  blk00000518 (
    .I0(sig00000015),
    .I1(sig0000000d),
    .I2(sig00000009),
    .I3(sig00000011),
    .I4(sig0000011a),
    .I5(sig0000011b),
    .O(sig000000bd)
  );
  LUT6 #(
    .INIT ( 64'hFF00CCCCF0F0AAAA ))
  blk00000519 (
    .I0(sig00000033),
    .I1(sig0000002f),
    .I2(sig0000002b),
    .I3(sig00000027),
    .I4(sig0000011a),
    .I5(sig0000011b),
    .O(sig000000db)
  );
  LUT6 #(
    .INIT ( 64'hFF00CCCCF0F0AAAA ))
  blk0000051a (
    .I0(sig00000034),
    .I1(sig00000030),
    .I2(sig0000002c),
    .I3(sig00000028),
    .I4(sig0000011a),
    .I5(sig0000011b),
    .O(sig000000dc)
  );
  LUT6 #(
    .INIT ( 64'hFF00CCCCF0F0AAAA ))
  blk0000051b (
    .I0(sig00000035),
    .I1(sig00000031),
    .I2(sig0000002d),
    .I3(sig00000029),
    .I4(sig0000011a),
    .I5(sig0000011b),
    .O(sig000000dd)
  );
  LUT6 #(
    .INIT ( 64'hFF00CCCCF0F0AAAA ))
  blk0000051c (
    .I0(sig00000036),
    .I1(sig00000032),
    .I2(sig0000002e),
    .I3(sig0000002a),
    .I4(sig0000011a),
    .I5(sig0000011b),
    .O(sig000000de)
  );
  LUT6 #(
    .INIT ( 64'hFF00CCCCF0F0AAAA ))
  blk0000051d (
    .I0(sig00000037),
    .I1(sig00000033),
    .I2(sig0000002f),
    .I3(sig0000002b),
    .I4(sig0000011a),
    .I5(sig0000011b),
    .O(sig000000df)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk0000051e (
    .I0(sig0000011d),
    .I1(sig0000011c),
    .I2(sig0000006d),
    .I3(sig0000006b),
    .I4(sig0000006c),
    .I5(sig0000006e),
    .O(sig00000114)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk0000051f (
    .I0(sig0000011d),
    .I1(sig0000011c),
    .I2(sig0000006b),
    .I3(sig00000069),
    .I4(sig0000006a),
    .I5(sig0000006c),
    .O(sig00000112)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk00000520 (
    .I0(sig0000011d),
    .I1(sig0000011c),
    .I2(sig00000041),
    .I3(sig0000003f),
    .I4(sig00000040),
    .I5(sig00000042),
    .O(sig000000e8)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk00000521 (
    .I0(sig0000011d),
    .I1(sig0000011c),
    .I2(sig0000003f),
    .I3(sig0000003d),
    .I4(sig0000003e),
    .I5(sig00000040),
    .O(sig000000e6)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk00000522 (
    .I0(sig0000011d),
    .I1(sig0000011c),
    .I2(sig00000042),
    .I3(sig00000040),
    .I4(sig00000041),
    .I5(sig00000043),
    .O(sig000000e9)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk00000523 (
    .I0(sig0000011d),
    .I1(sig0000011c),
    .I2(sig00000040),
    .I3(sig0000003e),
    .I4(sig0000003f),
    .I5(sig00000041),
    .O(sig000000e7)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk00000524 (
    .I0(sig0000011d),
    .I1(sig0000011c),
    .I2(sig00000043),
    .I3(sig00000041),
    .I4(sig00000042),
    .I5(sig00000044),
    .O(sig000000ea)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk00000525 (
    .I0(sig0000011d),
    .I1(sig0000011c),
    .I2(sig00000048),
    .I3(sig00000046),
    .I4(sig00000047),
    .I5(sig00000049),
    .O(sig000000ef)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk00000526 (
    .I0(sig0000011d),
    .I1(sig0000011c),
    .I2(sig00000046),
    .I3(sig00000044),
    .I4(sig00000045),
    .I5(sig00000047),
    .O(sig000000ed)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk00000527 (
    .I0(sig0000011d),
    .I1(sig0000011c),
    .I2(sig00000049),
    .I3(sig00000047),
    .I4(sig00000048),
    .I5(sig0000004a),
    .O(sig000000f0)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk00000528 (
    .I0(sig0000011d),
    .I1(sig0000011c),
    .I2(sig00000047),
    .I3(sig00000045),
    .I4(sig00000046),
    .I5(sig00000048),
    .O(sig000000ee)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk00000529 (
    .I0(sig0000011d),
    .I1(sig0000011c),
    .I2(sig0000004a),
    .I3(sig00000048),
    .I4(sig00000049),
    .I5(sig0000004b),
    .O(sig000000f1)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk0000052a (
    .I0(sig0000011d),
    .I1(sig0000011c),
    .I2(sig0000006e),
    .I3(sig0000006c),
    .I4(sig0000006d),
    .I5(sig0000006f),
    .O(sig00000115)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk0000052b (
    .I0(sig0000011d),
    .I1(sig0000011c),
    .I2(sig0000006c),
    .I3(sig0000006a),
    .I4(sig0000006b),
    .I5(sig0000006d),
    .O(sig00000113)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk0000052c (
    .I0(sig0000011d),
    .I1(sig0000011c),
    .I2(sig00000044),
    .I3(sig00000042),
    .I4(sig00000043),
    .I5(sig00000045),
    .O(sig000000eb)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk0000052d (
    .I0(sig0000011d),
    .I1(sig0000011c),
    .I2(sig00000051),
    .I3(sig0000004f),
    .I4(sig00000050),
    .I5(sig00000052),
    .O(sig000000f8)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk0000052e (
    .I0(sig0000011d),
    .I1(sig0000011c),
    .I2(sig0000004f),
    .I3(sig0000004d),
    .I4(sig0000004e),
    .I5(sig00000050),
    .O(sig000000f6)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk0000052f (
    .I0(sig0000011d),
    .I1(sig0000011c),
    .I2(sig00000052),
    .I3(sig00000050),
    .I4(sig00000051),
    .I5(sig00000053),
    .O(sig000000f9)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk00000530 (
    .I0(sig0000011d),
    .I1(sig0000011c),
    .I2(sig00000050),
    .I3(sig0000004e),
    .I4(sig0000004f),
    .I5(sig00000051),
    .O(sig000000f7)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk00000531 (
    .I0(sig0000011d),
    .I1(sig0000011c),
    .I2(sig00000053),
    .I3(sig00000051),
    .I4(sig00000052),
    .I5(sig00000054),
    .O(sig000000fa)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk00000532 (
    .I0(sig0000011d),
    .I1(sig0000011c),
    .I2(sig00000054),
    .I3(sig00000052),
    .I4(sig00000053),
    .I5(sig00000055),
    .O(sig000000fb)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk00000533 (
    .I0(sig0000011d),
    .I1(sig0000011c),
    .I2(sig0000004b),
    .I3(sig00000049),
    .I4(sig0000004a),
    .I5(sig0000004c),
    .O(sig000000f2)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk00000534 (
    .I0(sig0000011d),
    .I1(sig0000011c),
    .I2(sig0000006f),
    .I3(sig0000006d),
    .I4(sig0000006e),
    .I5(sig00000070),
    .O(sig00000116)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk00000535 (
    .I0(sig0000011d),
    .I1(sig0000011c),
    .I2(sig00000055),
    .I3(sig00000053),
    .I4(sig00000054),
    .I5(sig00000056),
    .O(sig000000fc)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk00000536 (
    .I0(sig0000011d),
    .I1(sig0000011c),
    .I2(sig00000056),
    .I3(sig00000054),
    .I4(sig00000055),
    .I5(sig00000057),
    .O(sig000000fd)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk00000537 (
    .I0(sig0000011d),
    .I1(sig0000011c),
    .I2(sig00000057),
    .I3(sig00000055),
    .I4(sig00000056),
    .I5(sig00000058),
    .O(sig000000fe)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk00000538 (
    .I0(sig0000011d),
    .I1(sig0000011c),
    .I2(sig00000058),
    .I3(sig00000056),
    .I4(sig00000057),
    .I5(sig00000059),
    .O(sig000000ff)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk00000539 (
    .I0(sig0000011d),
    .I1(sig0000011c),
    .I2(sig00000045),
    .I3(sig00000043),
    .I4(sig00000044),
    .I5(sig00000046),
    .O(sig000000ec)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk0000053a (
    .I0(sig0000011d),
    .I1(sig0000011c),
    .I2(sig00000059),
    .I3(sig00000057),
    .I4(sig00000058),
    .I5(sig0000005a),
    .O(sig00000100)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk0000053b (
    .I0(sig0000011d),
    .I1(sig0000011c),
    .I2(sig0000005a),
    .I3(sig00000058),
    .I4(sig00000059),
    .I5(sig0000005b),
    .O(sig00000101)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk0000053c (
    .I0(sig0000011d),
    .I1(sig0000011c),
    .I2(sig0000005b),
    .I3(sig00000059),
    .I4(sig0000005a),
    .I5(sig0000005c),
    .O(sig00000102)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk0000053d (
    .I0(sig0000011d),
    .I1(sig0000011c),
    .I2(sig0000005c),
    .I3(sig0000005a),
    .I4(sig0000005b),
    .I5(sig0000005d),
    .O(sig00000103)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk0000053e (
    .I0(sig0000011d),
    .I1(sig0000011c),
    .I2(sig0000005d),
    .I3(sig0000005b),
    .I4(sig0000005c),
    .I5(sig0000005e),
    .O(sig00000104)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk0000053f (
    .I0(sig0000011d),
    .I1(sig0000011c),
    .I2(sig0000004c),
    .I3(sig0000004a),
    .I4(sig0000004b),
    .I5(sig0000004d),
    .O(sig000000f3)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk00000540 (
    .I0(sig0000011d),
    .I1(sig0000011c),
    .I2(sig0000005e),
    .I3(sig0000005c),
    .I4(sig0000005d),
    .I5(sig0000005f),
    .O(sig00000105)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk00000541 (
    .I0(sig0000011d),
    .I1(sig0000011c),
    .I2(sig0000005f),
    .I3(sig0000005d),
    .I4(sig0000005e),
    .I5(sig00000060),
    .O(sig00000106)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk00000542 (
    .I0(sig0000011d),
    .I1(sig0000011c),
    .I2(sig00000060),
    .I3(sig0000005e),
    .I4(sig0000005f),
    .I5(sig00000061),
    .O(sig00000107)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk00000543 (
    .I0(sig0000011d),
    .I1(sig0000011c),
    .I2(sig00000061),
    .I3(sig0000005f),
    .I4(sig00000060),
    .I5(sig00000062),
    .O(sig00000108)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk00000544 (
    .I0(sig0000011d),
    .I1(sig0000011c),
    .I2(sig00000062),
    .I3(sig00000060),
    .I4(sig00000061),
    .I5(sig00000063),
    .O(sig00000109)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk00000545 (
    .I0(sig0000011d),
    .I1(sig0000011c),
    .I2(sig00000063),
    .I3(sig00000061),
    .I4(sig00000062),
    .I5(sig00000064),
    .O(sig0000010a)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk00000546 (
    .I0(sig0000011d),
    .I1(sig0000011c),
    .I2(sig00000064),
    .I3(sig00000062),
    .I4(sig00000063),
    .I5(sig00000065),
    .O(sig0000010b)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk00000547 (
    .I0(sig0000011d),
    .I1(sig0000011c),
    .I2(sig00000070),
    .I3(sig0000006e),
    .I4(sig0000006f),
    .I5(sig00000071),
    .O(sig00000117)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk00000548 (
    .I0(sig0000011d),
    .I1(sig0000011c),
    .I2(sig00000065),
    .I3(sig00000063),
    .I4(sig00000064),
    .I5(sig00000066),
    .O(sig0000010c)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk00000549 (
    .I0(sig0000011d),
    .I1(sig0000011c),
    .I2(sig00000066),
    .I3(sig00000064),
    .I4(sig00000065),
    .I5(sig00000067),
    .O(sig0000010d)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk0000054a (
    .I0(sig0000011d),
    .I1(sig0000011c),
    .I2(sig0000004d),
    .I3(sig0000004b),
    .I4(sig0000004c),
    .I5(sig0000004e),
    .O(sig000000f4)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk0000054b (
    .I0(sig0000011d),
    .I1(sig0000011c),
    .I2(sig00000067),
    .I3(sig00000065),
    .I4(sig00000066),
    .I5(sig00000068),
    .O(sig0000010e)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk0000054c (
    .I0(sig0000011d),
    .I1(sig0000011c),
    .I2(sig00000068),
    .I3(sig00000066),
    .I4(sig00000067),
    .I5(sig00000069),
    .O(sig0000010f)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk0000054d (
    .I0(sig0000011d),
    .I1(sig0000011c),
    .I2(sig00000069),
    .I3(sig00000067),
    .I4(sig00000068),
    .I5(sig0000006a),
    .O(sig00000110)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk0000054e (
    .I0(sig0000011d),
    .I1(sig0000011c),
    .I2(sig0000006a),
    .I3(sig00000068),
    .I4(sig00000069),
    .I5(sig0000006b),
    .O(sig00000111)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk0000054f (
    .I0(sig0000011d),
    .I1(sig0000011c),
    .I2(sig0000003c),
    .I3(sig0000003a),
    .I4(sig0000003b),
    .I5(sig0000003d),
    .O(sig000000e3)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk00000550 (
    .I0(sig0000011d),
    .I1(sig0000011c),
    .I2(sig0000003d),
    .I3(sig0000003b),
    .I4(sig0000003c),
    .I5(sig0000003e),
    .O(sig000000e4)
  );
  LUT5 #(
    .INIT ( 32'h00AAF0CC ))
  blk00000551 (
    .I0(sig0000003a),
    .I1(sig0000003c),
    .I2(sig0000003b),
    .I3(sig0000011d),
    .I4(sig0000011c),
    .O(sig000000e2)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk00000552 (
    .I0(sig0000011d),
    .I1(sig0000011c),
    .I2(sig0000003e),
    .I3(sig0000003c),
    .I4(sig0000003d),
    .I5(sig0000003f),
    .O(sig000000e5)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk00000553 (
    .I0(sig0000011d),
    .I1(sig0000011c),
    .I2(sig0000004e),
    .I3(sig0000004c),
    .I4(sig0000004d),
    .I5(sig0000004f),
    .O(sig000000f5)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000554 (
    .I0(a[52]),
    .I1(b[52]),
    .O(sig00000156)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000555 (
    .I0(b[63]),
    .I1(operation[0]),
    .O(sig000002a9)
  );
  LUT3 #(
    .INIT ( 8'hF8 ))
  blk00000556 (
    .I0(sig0000027c),
    .I1(sig0000027a),
    .I2(sig0000027b),
    .O(sig0000022e)
  );
  LUT5 #(
    .INIT ( 32'hFEEE0222 ))
  blk00000557 (
    .I0(sig000002f5),
    .I1(sig0000027b),
    .I2(sig0000027c),
    .I3(sig0000027a),
    .I4(sig000002f4),
    .O(sig000002a8)
  );
  LUT4 #(
    .INIT ( 16'hAA8A ))
  blk00000558 (
    .I0(sig000002ea),
    .I1(sig000002eb),
    .I2(sig0000030c),
    .I3(sig000002ec),
    .O(sig000002a0)
  );
  LUT4 #(
    .INIT ( 16'hEA2A ))
  blk00000559 (
    .I0(sig000002f4),
    .I1(sig00000313),
    .I2(sig00000314),
    .I3(sig000002f5),
    .O(sig000002a6)
  );
  LUT4 #(
    .INIT ( 16'h8000 ))
  blk0000055a (
    .I0(sig00000313),
    .I1(sig00000314),
    .I2(sig00000310),
    .I3(sig00000311),
    .O(sig00000293)
  );
  LUT4 #(
    .INIT ( 16'hF888 ))
  blk0000055b (
    .I0(sig00000313),
    .I1(sig00000314),
    .I2(sig00000310),
    .I3(sig00000311),
    .O(sig00000292)
  );
  LUT5 #(
    .INIT ( 32'hFFFF1504 ))
  blk0000055c (
    .I0(sig000002f2),
    .I1(sig000002f1),
    .I2(sig000004b6),
    .I3(sig000002ef),
    .I4(sig000002f3),
    .O(sig000002a5)
  );
  LUT4 #(
    .INIT ( 16'h5554 ))
  blk0000055d (
    .I0(sig000002f3),
    .I1(sig000002f1),
    .I2(sig000002ef),
    .I3(sig000002f2),
    .O(sig000002a4)
  );
  LUT6 #(
    .INIT ( 64'hFFFFFFFF55555554 ))
  blk0000055e (
    .I0(sig000002eb),
    .I1(sig0000030c),
    .I2(sig000002b8),
    .I3(sig000002c5),
    .I4(sig000002c4),
    .I5(sig000002ec),
    .O(sig000002a2)
  );
  LUT6 #(
    .INIT ( 64'hAAAAAAAAAAAAABAA ))
  blk0000055f (
    .I0(sig000002eb),
    .I1(sig0000030c),
    .I2(sig000002ec),
    .I3(sig000002c5),
    .I4(sig000002b8),
    .I5(sig000002c4),
    .O(sig000002a1)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk00000560 (
    .I0(sig0000024a),
    .I1(sig0000030b),
    .I2(sig00000300),
    .O(sig0000028e)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000561 (
    .I0(sig000002f7),
    .I1(sig00000302),
    .I2(sig0000024a),
    .O(sig00000285)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000562 (
    .I0(sig000002f8),
    .I1(sig00000303),
    .I2(sig0000024a),
    .O(sig00000286)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000563 (
    .I0(sig000002f9),
    .I1(sig00000304),
    .I2(sig0000024a),
    .O(sig00000287)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000564 (
    .I0(sig000002fa),
    .I1(sig00000305),
    .I2(sig0000024a),
    .O(sig00000288)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000565 (
    .I0(sig000002fb),
    .I1(sig00000306),
    .I2(sig0000024a),
    .O(sig00000289)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000566 (
    .I0(sig000002fc),
    .I1(sig00000307),
    .I2(sig0000024a),
    .O(sig0000028a)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk00000567 (
    .I0(sig0000024a),
    .I1(sig00000308),
    .I2(sig000002fd),
    .O(sig0000028b)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk00000568 (
    .I0(sig0000024a),
    .I1(sig00000309),
    .I2(sig000002fe),
    .O(sig0000028c)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk00000569 (
    .I0(sig0000024a),
    .I1(sig0000030a),
    .I2(sig000002ff),
    .O(sig0000028d)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk0000056a (
    .I0(sig000002f5),
    .I1(sig000002f4),
    .O(sig00000290)
  );
  LUT3 #(
    .INIT ( 8'h53 ))
  blk0000056b (
    .I0(sig00000301),
    .I1(sig000002f6),
    .I2(sig0000024a),
    .O(sig00000284)
  );
  LUT2 #(
    .INIT ( 4'hE ))
  blk0000056c (
    .I0(sig000002b7),
    .I1(sig000002b6),
    .O(sig00000277)
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  blk0000056d (
    .I0(sig000002b6),
    .I1(sig000002b7),
    .O(sig00000278)
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  blk0000056e (
    .I0(sig000002b7),
    .I1(sig000002b6),
    .O(sig00000279)
  );
  LUT4 #(
    .INIT ( 16'h22F2 ))
  blk0000056f (
    .I0(sig00000313),
    .I1(sig00000314),
    .I2(sig00000310),
    .I3(sig00000311),
    .O(sig00000291)
  );
  LUT2 #(
    .INIT ( 4'h8 ))
  blk00000570 (
    .I0(sig000002c6),
    .I1(sig0000030d),
    .O(sig0000029f)
  );
  LUT2 #(
    .INIT ( 4'h8 ))
  blk00000571 (
    .I0(sig000002f5),
    .I1(sig000002f4),
    .O(sig000002a7)
  );
  LUT2 #(
    .INIT ( 4'hE ))
  blk00000572 (
    .I0(sig0000030f),
    .I1(sig00000312),
    .O(sig0000022c)
  );
  LUT2 #(
    .INIT ( 4'h8 ))
  blk00000573 (
    .I0(sig0000030f),
    .I1(sig00000312),
    .O(sig0000022d)
  );
  LUT6 #(
    .INIT ( 64'h0000000000000001 ))
  blk00000574 (
    .I0(a[42]),
    .I1(a[43]),
    .I2(a[44]),
    .I3(a[45]),
    .I4(a[46]),
    .I5(a[47]),
    .O(sig00000315)
  );
  LUT6 #(
    .INIT ( 64'h0000000000000001 ))
  blk00000575 (
    .I0(a[36]),
    .I1(a[37]),
    .I2(a[38]),
    .I3(a[39]),
    .I4(a[40]),
    .I5(a[41]),
    .O(sig00000316)
  );
  LUT6 #(
    .INIT ( 64'h0000000000000001 ))
  blk00000576 (
    .I0(a[30]),
    .I1(a[31]),
    .I2(a[32]),
    .I3(a[33]),
    .I4(a[34]),
    .I5(a[35]),
    .O(sig00000317)
  );
  LUT6 #(
    .INIT ( 64'h0000000000000001 ))
  blk00000577 (
    .I0(a[24]),
    .I1(a[25]),
    .I2(a[26]),
    .I3(a[27]),
    .I4(a[28]),
    .I5(a[29]),
    .O(sig00000318)
  );
  LUT6 #(
    .INIT ( 64'h0000000000000001 ))
  blk00000578 (
    .I0(a[18]),
    .I1(a[19]),
    .I2(a[20]),
    .I3(a[21]),
    .I4(a[22]),
    .I5(a[23]),
    .O(sig00000319)
  );
  LUT6 #(
    .INIT ( 64'h0000000000000001 ))
  blk00000579 (
    .I0(a[12]),
    .I1(a[13]),
    .I2(a[14]),
    .I3(a[15]),
    .I4(a[16]),
    .I5(a[17]),
    .O(sig0000031a)
  );
  LUT6 #(
    .INIT ( 64'h0000000000000001 ))
  blk0000057a (
    .I0(a[6]),
    .I1(a[7]),
    .I2(a[8]),
    .I3(a[9]),
    .I4(a[10]),
    .I5(a[11]),
    .O(sig0000031b)
  );
  LUT6 #(
    .INIT ( 64'h0000000000000001 ))
  blk0000057b (
    .I0(a[0]),
    .I1(a[1]),
    .I2(a[2]),
    .I3(a[3]),
    .I4(a[4]),
    .I5(a[5]),
    .O(sig0000031c)
  );
  LUT4 #(
    .INIT ( 16'h0001 ))
  blk0000057c (
    .I0(a[48]),
    .I1(a[49]),
    .I2(a[50]),
    .I3(a[51]),
    .O(sig0000031d)
  );
  LUT6 #(
    .INIT ( 64'h0000000000000001 ))
  blk0000057d (
    .I0(b[42]),
    .I1(b[43]),
    .I2(b[44]),
    .I3(b[45]),
    .I4(b[46]),
    .I5(b[47]),
    .O(sig0000031e)
  );
  LUT6 #(
    .INIT ( 64'h0000000000000001 ))
  blk0000057e (
    .I0(b[36]),
    .I1(b[37]),
    .I2(b[38]),
    .I3(b[39]),
    .I4(b[40]),
    .I5(b[41]),
    .O(sig0000031f)
  );
  LUT6 #(
    .INIT ( 64'h0000000000000001 ))
  blk0000057f (
    .I0(b[30]),
    .I1(b[31]),
    .I2(b[32]),
    .I3(b[33]),
    .I4(b[34]),
    .I5(b[35]),
    .O(sig00000320)
  );
  LUT6 #(
    .INIT ( 64'h0000000000000001 ))
  blk00000580 (
    .I0(b[24]),
    .I1(b[25]),
    .I2(b[26]),
    .I3(b[27]),
    .I4(b[28]),
    .I5(b[29]),
    .O(sig00000321)
  );
  LUT6 #(
    .INIT ( 64'h0000000000000001 ))
  blk00000581 (
    .I0(b[18]),
    .I1(b[19]),
    .I2(b[20]),
    .I3(b[21]),
    .I4(b[22]),
    .I5(b[23]),
    .O(sig00000322)
  );
  LUT6 #(
    .INIT ( 64'h0000000000000001 ))
  blk00000582 (
    .I0(b[12]),
    .I1(b[13]),
    .I2(b[14]),
    .I3(b[15]),
    .I4(b[16]),
    .I5(b[17]),
    .O(sig00000323)
  );
  LUT6 #(
    .INIT ( 64'h0000000000000001 ))
  blk00000583 (
    .I0(b[6]),
    .I1(b[7]),
    .I2(b[8]),
    .I3(b[9]),
    .I4(b[10]),
    .I5(b[11]),
    .O(sig00000324)
  );
  LUT6 #(
    .INIT ( 64'h0000000000000001 ))
  blk00000584 (
    .I0(b[0]),
    .I1(b[1]),
    .I2(b[2]),
    .I3(b[3]),
    .I4(b[4]),
    .I5(b[5]),
    .O(sig00000325)
  );
  LUT4 #(
    .INIT ( 16'h0001 ))
  blk00000585 (
    .I0(b[48]),
    .I1(b[49]),
    .I2(b[50]),
    .I3(b[51]),
    .O(sig00000326)
  );
  LUT4 #(
    .INIT ( 16'h9009 ))
  blk00000586 (
    .I0(b[19]),
    .I1(a[19]),
    .I2(b[18]),
    .I3(a[18]),
    .O(sig00000346)
  );
  LUT4 #(
    .INIT ( 16'h9009 ))
  blk00000587 (
    .I0(b[17]),
    .I1(a[17]),
    .I2(b[16]),
    .I3(a[16]),
    .O(sig00000348)
  );
  LUT4 #(
    .INIT ( 16'h9009 ))
  blk00000588 (
    .I0(b[15]),
    .I1(a[15]),
    .I2(b[14]),
    .I3(a[14]),
    .O(sig0000034a)
  );
  LUT4 #(
    .INIT ( 16'h9009 ))
  blk00000589 (
    .I0(b[13]),
    .I1(a[13]),
    .I2(b[12]),
    .I3(a[12]),
    .O(sig0000034c)
  );
  LUT4 #(
    .INIT ( 16'h9009 ))
  blk0000058a (
    .I0(b[11]),
    .I1(a[11]),
    .I2(b[10]),
    .I3(a[10]),
    .O(sig0000034e)
  );
  LUT4 #(
    .INIT ( 16'h9009 ))
  blk0000058b (
    .I0(b[9]),
    .I1(a[9]),
    .I2(b[8]),
    .I3(a[8]),
    .O(sig00000350)
  );
  LUT4 #(
    .INIT ( 16'h9009 ))
  blk0000058c (
    .I0(b[7]),
    .I1(a[7]),
    .I2(b[6]),
    .I3(a[6]),
    .O(sig00000352)
  );
  LUT4 #(
    .INIT ( 16'h9009 ))
  blk0000058d (
    .I0(b[5]),
    .I1(a[5]),
    .I2(b[4]),
    .I3(a[4]),
    .O(sig00000354)
  );
  LUT4 #(
    .INIT ( 16'h9009 ))
  blk0000058e (
    .I0(b[3]),
    .I1(a[3]),
    .I2(b[2]),
    .I3(a[2]),
    .O(sig00000356)
  );
  LUT4 #(
    .INIT ( 16'h9009 ))
  blk0000058f (
    .I0(b[31]),
    .I1(a[31]),
    .I2(b[30]),
    .I3(a[30]),
    .O(sig0000033a)
  );
  LUT4 #(
    .INIT ( 16'h9009 ))
  blk00000590 (
    .I0(b[29]),
    .I1(a[29]),
    .I2(b[28]),
    .I3(a[28]),
    .O(sig0000033c)
  );
  LUT4 #(
    .INIT ( 16'h9009 ))
  blk00000591 (
    .I0(b[27]),
    .I1(a[27]),
    .I2(b[26]),
    .I3(a[26]),
    .O(sig0000033e)
  );
  LUT4 #(
    .INIT ( 16'h9009 ))
  blk00000592 (
    .I0(b[25]),
    .I1(a[25]),
    .I2(b[24]),
    .I3(a[24]),
    .O(sig00000340)
  );
  LUT4 #(
    .INIT ( 16'h9009 ))
  blk00000593 (
    .I0(b[23]),
    .I1(a[23]),
    .I2(b[22]),
    .I3(a[22]),
    .O(sig00000342)
  );
  LUT4 #(
    .INIT ( 16'h9009 ))
  blk00000594 (
    .I0(b[21]),
    .I1(a[21]),
    .I2(b[20]),
    .I3(a[20]),
    .O(sig00000344)
  );
  LUT4 #(
    .INIT ( 16'h9009 ))
  blk00000595 (
    .I0(b[1]),
    .I1(a[1]),
    .I2(b[0]),
    .I3(a[0]),
    .O(sig00000358)
  );
  LUT4 #(
    .INIT ( 16'h22B2 ))
  blk00000596 (
    .I0(b[31]),
    .I1(a[31]),
    .I2(b[30]),
    .I3(a[30]),
    .O(sig00000339)
  );
  LUT4 #(
    .INIT ( 16'h22B2 ))
  blk00000597 (
    .I0(b[29]),
    .I1(a[29]),
    .I2(b[28]),
    .I3(a[28]),
    .O(sig0000033b)
  );
  LUT4 #(
    .INIT ( 16'h22B2 ))
  blk00000598 (
    .I0(b[27]),
    .I1(a[27]),
    .I2(b[26]),
    .I3(a[26]),
    .O(sig0000033d)
  );
  LUT4 #(
    .INIT ( 16'h22B2 ))
  blk00000599 (
    .I0(b[25]),
    .I1(a[25]),
    .I2(b[24]),
    .I3(a[24]),
    .O(sig0000033f)
  );
  LUT4 #(
    .INIT ( 16'h22B2 ))
  blk0000059a (
    .I0(b[23]),
    .I1(a[23]),
    .I2(b[22]),
    .I3(a[22]),
    .O(sig00000341)
  );
  LUT4 #(
    .INIT ( 16'h22B2 ))
  blk0000059b (
    .I0(b[21]),
    .I1(a[21]),
    .I2(b[20]),
    .I3(a[20]),
    .O(sig00000343)
  );
  LUT4 #(
    .INIT ( 16'h22B2 ))
  blk0000059c (
    .I0(b[19]),
    .I1(a[19]),
    .I2(b[18]),
    .I3(a[18]),
    .O(sig00000345)
  );
  LUT4 #(
    .INIT ( 16'h22B2 ))
  blk0000059d (
    .I0(b[17]),
    .I1(a[17]),
    .I2(b[16]),
    .I3(a[16]),
    .O(sig00000347)
  );
  LUT4 #(
    .INIT ( 16'h22B2 ))
  blk0000059e (
    .I0(b[15]),
    .I1(a[15]),
    .I2(b[14]),
    .I3(a[14]),
    .O(sig00000349)
  );
  LUT4 #(
    .INIT ( 16'h22B2 ))
  blk0000059f (
    .I0(b[13]),
    .I1(a[13]),
    .I2(b[12]),
    .I3(a[12]),
    .O(sig0000034b)
  );
  LUT4 #(
    .INIT ( 16'h22B2 ))
  blk000005a0 (
    .I0(b[11]),
    .I1(a[11]),
    .I2(b[10]),
    .I3(a[10]),
    .O(sig0000034d)
  );
  LUT4 #(
    .INIT ( 16'h22B2 ))
  blk000005a1 (
    .I0(b[9]),
    .I1(a[9]),
    .I2(b[8]),
    .I3(a[8]),
    .O(sig0000034f)
  );
  LUT4 #(
    .INIT ( 16'h22B2 ))
  blk000005a2 (
    .I0(b[7]),
    .I1(a[7]),
    .I2(b[6]),
    .I3(a[6]),
    .O(sig00000351)
  );
  LUT4 #(
    .INIT ( 16'h22B2 ))
  blk000005a3 (
    .I0(b[5]),
    .I1(a[5]),
    .I2(b[4]),
    .I3(a[4]),
    .O(sig00000353)
  );
  LUT4 #(
    .INIT ( 16'h22B2 ))
  blk000005a4 (
    .I0(b[3]),
    .I1(a[3]),
    .I2(b[2]),
    .I3(a[2]),
    .O(sig00000355)
  );
  LUT4 #(
    .INIT ( 16'h22B2 ))
  blk000005a5 (
    .I0(b[1]),
    .I1(a[1]),
    .I2(b[0]),
    .I3(a[0]),
    .O(sig00000357)
  );
  LUT4 #(
    .INIT ( 16'h9009 ))
  blk000005a6 (
    .I0(b[51]),
    .I1(a[51]),
    .I2(b[50]),
    .I3(a[50]),
    .O(sig00000366)
  );
  LUT4 #(
    .INIT ( 16'h9009 ))
  blk000005a7 (
    .I0(b[49]),
    .I1(a[49]),
    .I2(b[48]),
    .I3(a[48]),
    .O(sig00000368)
  );
  LUT4 #(
    .INIT ( 16'h9009 ))
  blk000005a8 (
    .I0(b[47]),
    .I1(a[47]),
    .I2(b[46]),
    .I3(a[46]),
    .O(sig0000036a)
  );
  LUT4 #(
    .INIT ( 16'h9009 ))
  blk000005a9 (
    .I0(b[45]),
    .I1(a[45]),
    .I2(b[44]),
    .I3(a[44]),
    .O(sig0000036c)
  );
  LUT4 #(
    .INIT ( 16'h9009 ))
  blk000005aa (
    .I0(b[43]),
    .I1(a[43]),
    .I2(b[42]),
    .I3(a[42]),
    .O(sig0000036e)
  );
  LUT4 #(
    .INIT ( 16'h9009 ))
  blk000005ab (
    .I0(b[41]),
    .I1(a[41]),
    .I2(b[40]),
    .I3(a[40]),
    .O(sig00000370)
  );
  LUT4 #(
    .INIT ( 16'h9009 ))
  blk000005ac (
    .I0(b[39]),
    .I1(a[39]),
    .I2(b[38]),
    .I3(a[38]),
    .O(sig00000372)
  );
  LUT4 #(
    .INIT ( 16'h9009 ))
  blk000005ad (
    .I0(b[37]),
    .I1(a[37]),
    .I2(b[36]),
    .I3(a[36]),
    .O(sig00000374)
  );
  LUT4 #(
    .INIT ( 16'h9009 ))
  blk000005ae (
    .I0(b[35]),
    .I1(a[35]),
    .I2(b[34]),
    .I3(a[34]),
    .O(sig00000376)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk000005af (
    .I0(b[62]),
    .I1(a[62]),
    .O(sig0000035a)
  );
  LUT4 #(
    .INIT ( 16'h9009 ))
  blk000005b0 (
    .I0(b[61]),
    .I1(a[61]),
    .I2(b[60]),
    .I3(a[60]),
    .O(sig0000035c)
  );
  LUT4 #(
    .INIT ( 16'h9009 ))
  blk000005b1 (
    .I0(b[59]),
    .I1(a[59]),
    .I2(b[58]),
    .I3(a[58]),
    .O(sig0000035e)
  );
  LUT4 #(
    .INIT ( 16'h9009 ))
  blk000005b2 (
    .I0(b[57]),
    .I1(a[57]),
    .I2(b[56]),
    .I3(a[56]),
    .O(sig00000360)
  );
  LUT4 #(
    .INIT ( 16'h9009 ))
  blk000005b3 (
    .I0(b[55]),
    .I1(a[55]),
    .I2(b[54]),
    .I3(a[54]),
    .O(sig00000362)
  );
  LUT4 #(
    .INIT ( 16'h9009 ))
  blk000005b4 (
    .I0(b[53]),
    .I1(a[53]),
    .I2(b[52]),
    .I3(a[52]),
    .O(sig00000364)
  );
  LUT4 #(
    .INIT ( 16'h9009 ))
  blk000005b5 (
    .I0(b[33]),
    .I1(a[33]),
    .I2(b[32]),
    .I3(a[32]),
    .O(sig00000378)
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  blk000005b6 (
    .I0(b[62]),
    .I1(a[62]),
    .O(sig00000359)
  );
  LUT4 #(
    .INIT ( 16'h22B2 ))
  blk000005b7 (
    .I0(b[61]),
    .I1(a[61]),
    .I2(b[60]),
    .I3(a[60]),
    .O(sig0000035b)
  );
  LUT4 #(
    .INIT ( 16'h22B2 ))
  blk000005b8 (
    .I0(b[59]),
    .I1(a[59]),
    .I2(b[58]),
    .I3(a[58]),
    .O(sig0000035d)
  );
  LUT4 #(
    .INIT ( 16'h22B2 ))
  blk000005b9 (
    .I0(b[57]),
    .I1(a[57]),
    .I2(b[56]),
    .I3(a[56]),
    .O(sig0000035f)
  );
  LUT4 #(
    .INIT ( 16'h22B2 ))
  blk000005ba (
    .I0(b[55]),
    .I1(a[55]),
    .I2(b[54]),
    .I3(a[54]),
    .O(sig00000361)
  );
  LUT4 #(
    .INIT ( 16'h22B2 ))
  blk000005bb (
    .I0(b[53]),
    .I1(a[53]),
    .I2(b[52]),
    .I3(a[52]),
    .O(sig00000363)
  );
  LUT4 #(
    .INIT ( 16'h22B2 ))
  blk000005bc (
    .I0(b[51]),
    .I1(a[51]),
    .I2(b[50]),
    .I3(a[50]),
    .O(sig00000365)
  );
  LUT4 #(
    .INIT ( 16'h22B2 ))
  blk000005bd (
    .I0(b[49]),
    .I1(a[49]),
    .I2(b[48]),
    .I3(a[48]),
    .O(sig00000367)
  );
  LUT4 #(
    .INIT ( 16'h22B2 ))
  blk000005be (
    .I0(b[47]),
    .I1(a[47]),
    .I2(b[46]),
    .I3(a[46]),
    .O(sig00000369)
  );
  LUT4 #(
    .INIT ( 16'h22B2 ))
  blk000005bf (
    .I0(b[45]),
    .I1(a[45]),
    .I2(b[44]),
    .I3(a[44]),
    .O(sig0000036b)
  );
  LUT4 #(
    .INIT ( 16'h22B2 ))
  blk000005c0 (
    .I0(b[43]),
    .I1(a[43]),
    .I2(b[42]),
    .I3(a[42]),
    .O(sig0000036d)
  );
  LUT4 #(
    .INIT ( 16'h22B2 ))
  blk000005c1 (
    .I0(b[41]),
    .I1(a[41]),
    .I2(b[40]),
    .I3(a[40]),
    .O(sig0000036f)
  );
  LUT4 #(
    .INIT ( 16'h22B2 ))
  blk000005c2 (
    .I0(b[39]),
    .I1(a[39]),
    .I2(b[38]),
    .I3(a[38]),
    .O(sig00000371)
  );
  LUT4 #(
    .INIT ( 16'h22B2 ))
  blk000005c3 (
    .I0(b[37]),
    .I1(a[37]),
    .I2(b[36]),
    .I3(a[36]),
    .O(sig00000373)
  );
  LUT4 #(
    .INIT ( 16'h22B2 ))
  blk000005c4 (
    .I0(b[35]),
    .I1(a[35]),
    .I2(b[34]),
    .I3(a[34]),
    .O(sig00000375)
  );
  LUT4 #(
    .INIT ( 16'h22B2 ))
  blk000005c5 (
    .I0(b[33]),
    .I1(a[33]),
    .I2(b[32]),
    .I3(a[32]),
    .O(sig00000377)
  );
  LUT6 #(
    .INIT ( 64'h9009000000009009 ))
  blk000005c6 (
    .I0(b[59]),
    .I1(a[59]),
    .I2(b[61]),
    .I3(a[61]),
    .I4(b[60]),
    .I5(a[60]),
    .O(sig0000039a)
  );
  LUT6 #(
    .INIT ( 64'h9009000000009009 ))
  blk000005c7 (
    .I0(b[56]),
    .I1(a[56]),
    .I2(b[58]),
    .I3(a[58]),
    .I4(b[57]),
    .I5(a[57]),
    .O(sig0000039b)
  );
  LUT6 #(
    .INIT ( 64'h9009000000009009 ))
  blk000005c8 (
    .I0(b[53]),
    .I1(a[53]),
    .I2(b[55]),
    .I3(a[55]),
    .I4(b[54]),
    .I5(a[54]),
    .O(sig0000039c)
  );
  LUT6 #(
    .INIT ( 64'h9009000000009009 ))
  blk000005c9 (
    .I0(b[50]),
    .I1(a[50]),
    .I2(b[52]),
    .I3(a[52]),
    .I4(b[51]),
    .I5(a[51]),
    .O(sig0000039d)
  );
  LUT6 #(
    .INIT ( 64'h9009000000009009 ))
  blk000005ca (
    .I0(b[47]),
    .I1(a[47]),
    .I2(b[49]),
    .I3(a[49]),
    .I4(b[48]),
    .I5(a[48]),
    .O(sig0000039e)
  );
  LUT6 #(
    .INIT ( 64'h9009000000009009 ))
  blk000005cb (
    .I0(b[44]),
    .I1(a[44]),
    .I2(b[46]),
    .I3(a[46]),
    .I4(b[45]),
    .I5(a[45]),
    .O(sig0000039f)
  );
  LUT6 #(
    .INIT ( 64'h9009000000009009 ))
  blk000005cc (
    .I0(b[42]),
    .I1(a[42]),
    .I2(b[41]),
    .I3(a[41]),
    .I4(b[43]),
    .I5(a[43]),
    .O(sig000003a0)
  );
  LUT6 #(
    .INIT ( 64'h9009000000009009 ))
  blk000005cd (
    .I0(b[38]),
    .I1(a[38]),
    .I2(b[40]),
    .I3(a[40]),
    .I4(b[39]),
    .I5(a[39]),
    .O(sig000003a1)
  );
  LUT6 #(
    .INIT ( 64'h9009000000009009 ))
  blk000005ce (
    .I0(b[35]),
    .I1(a[35]),
    .I2(b[37]),
    .I3(a[37]),
    .I4(b[36]),
    .I5(a[36]),
    .O(sig000003a2)
  );
  LUT6 #(
    .INIT ( 64'h9009000000009009 ))
  blk000005cf (
    .I0(b[32]),
    .I1(a[32]),
    .I2(b[34]),
    .I3(a[34]),
    .I4(b[33]),
    .I5(a[33]),
    .O(sig000003a3)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk000005d0 (
    .I0(a[62]),
    .I1(b[62]),
    .O(sig00000399)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk000005d1 (
    .I0(sig000003d5),
    .I1(sig000003d4),
    .I2(sig000004ec),
    .I3(sig0000050c),
    .I4(sig000004fc),
    .I5(sig000004dc),
    .O(sig0000043f)
  );
  LUT4 #(
    .INIT ( 16'h5410 ))
  blk000005d2 (
    .I0(sig000003d4),
    .I1(sig000003d5),
    .I2(sig000004fc),
    .I3(sig0000050c),
    .O(sig0000041f)
  );
  LUT5 #(
    .INIT ( 32'hE6C4A280 ))
  blk000005d3 (
    .I0(sig000003d4),
    .I1(sig000003d5),
    .I2(sig00000506),
    .I3(sig000004f6),
    .I4(sig000004e6),
    .O(sig00000445)
  );
  LUT4 #(
    .INIT ( 16'h5410 ))
  blk000005d4 (
    .I0(sig000003d4),
    .I1(sig000003d5),
    .I2(sig000004f6),
    .I3(sig00000506),
    .O(sig00000425)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk000005d5 (
    .I0(sig000003d5),
    .I1(sig000003d4),
    .I2(sig000004eb),
    .I3(sig0000050b),
    .I4(sig000004fb),
    .I5(sig000004db),
    .O(sig00000440)
  );
  LUT4 #(
    .INIT ( 16'h5410 ))
  blk000005d6 (
    .I0(sig000003d4),
    .I1(sig000003d5),
    .I2(sig000004fb),
    .I3(sig0000050b),
    .O(sig00000420)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk000005d7 (
    .I0(sig000003d5),
    .I1(sig000003d4),
    .I2(sig000004ea),
    .I3(sig0000050a),
    .I4(sig000004fa),
    .I5(sig000004da),
    .O(sig00000441)
  );
  LUT4 #(
    .INIT ( 16'h5410 ))
  blk000005d8 (
    .I0(sig000003d4),
    .I1(sig000003d5),
    .I2(sig000004fa),
    .I3(sig0000050a),
    .O(sig00000421)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk000005d9 (
    .I0(sig000003d5),
    .I1(sig000003d4),
    .I2(sig000004e8),
    .I3(sig00000508),
    .I4(sig000004f8),
    .I5(sig000004d8),
    .O(sig00000443)
  );
  LUT4 #(
    .INIT ( 16'h5410 ))
  blk000005da (
    .I0(sig000003d4),
    .I1(sig000003d5),
    .I2(sig000004f8),
    .I3(sig00000508),
    .O(sig00000423)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk000005db (
    .I0(sig000003d5),
    .I1(sig000003d4),
    .I2(sig000004e9),
    .I3(sig00000509),
    .I4(sig000004f9),
    .I5(sig000004d9),
    .O(sig00000442)
  );
  LUT4 #(
    .INIT ( 16'h5410 ))
  blk000005dc (
    .I0(sig000003d4),
    .I1(sig000003d5),
    .I2(sig000004f9),
    .I3(sig00000509),
    .O(sig00000422)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk000005dd (
    .I0(sig000003d5),
    .I1(sig000003d4),
    .I2(sig000004e7),
    .I3(sig00000507),
    .I4(sig000004f7),
    .I5(sig000004d7),
    .O(sig00000444)
  );
  LUT4 #(
    .INIT ( 16'h5410 ))
  blk000005de (
    .I0(sig000003d4),
    .I1(sig000003d5),
    .I2(sig000004f7),
    .I3(sig00000507),
    .O(sig00000424)
  );
  LUT6 #(
    .INIT ( 64'hF0F0FF00CCCCAAAA ))
  blk000005df (
    .I0(sig000001ea),
    .I1(sig000001eb),
    .I2(sig0000021f),
    .I3(sig0000021e),
    .I4(sig0000023f),
    .I5(sig0000022e),
    .O(sig00000536)
  );
  LUT6 #(
    .INIT ( 64'hF0F0FF00CCCCAAAA ))
  blk000005e0 (
    .I0(sig000001eb),
    .I1(sig000001ec),
    .I2(sig00000220),
    .I3(sig0000021f),
    .I4(sig0000023f),
    .I5(sig0000022e),
    .O(sig00000537)
  );
  LUT6 #(
    .INIT ( 64'hF0F0FF00CCCCAAAA ))
  blk000005e1 (
    .I0(sig000001e9),
    .I1(sig000001ea),
    .I2(sig0000021e),
    .I3(sig0000021d),
    .I4(sig0000023f),
    .I5(sig0000022e),
    .O(sig00000535)
  );
  LUT6 #(
    .INIT ( 64'hF0F0FF00CCCCAAAA ))
  blk000005e2 (
    .I0(sig000001e8),
    .I1(sig000001e9),
    .I2(sig0000021d),
    .I3(sig0000021c),
    .I4(sig0000023f),
    .I5(sig0000022e),
    .O(sig00000534)
  );
  LUT6 #(
    .INIT ( 64'hF0F0FF00CCCCAAAA ))
  blk000005e3 (
    .I0(sig000001e7),
    .I1(sig000001e8),
    .I2(sig0000021c),
    .I3(sig0000021b),
    .I4(sig0000023f),
    .I5(sig0000022e),
    .O(sig00000533)
  );
  LUT6 #(
    .INIT ( 64'hF0F0FF00CCCCAAAA ))
  blk000005e4 (
    .I0(sig000001e3),
    .I1(sig000001e4),
    .I2(sig00000218),
    .I3(sig00000217),
    .I4(sig0000023f),
    .I5(sig0000022e),
    .O(sig0000052f)
  );
  LUT6 #(
    .INIT ( 64'hF0F0FF00CCCCAAAA ))
  blk000005e5 (
    .I0(sig000001e4),
    .I1(sig000001e5),
    .I2(sig00000219),
    .I3(sig00000218),
    .I4(sig0000023f),
    .I5(sig0000022e),
    .O(sig00000530)
  );
  LUT6 #(
    .INIT ( 64'hF0F0FF00CCCCAAAA ))
  blk000005e6 (
    .I0(sig000001e2),
    .I1(sig000001e3),
    .I2(sig00000217),
    .I3(sig00000216),
    .I4(sig0000023f),
    .I5(sig0000022e),
    .O(sig0000052e)
  );
  LUT6 #(
    .INIT ( 64'hF0F0FF00CCCCAAAA ))
  blk000005e7 (
    .I0(sig000001e6),
    .I1(sig000001e7),
    .I2(sig0000021b),
    .I3(sig0000021a),
    .I4(sig0000023f),
    .I5(sig0000022e),
    .O(sig00000532)
  );
  LUT6 #(
    .INIT ( 64'hF0F0FF00CCCCAAAA ))
  blk000005e8 (
    .I0(sig000001e1),
    .I1(sig000001e2),
    .I2(sig00000216),
    .I3(sig00000215),
    .I4(sig0000023f),
    .I5(sig0000022e),
    .O(sig0000052d)
  );
  LUT6 #(
    .INIT ( 64'hF0F0FF00CCCCAAAA ))
  blk000005e9 (
    .I0(sig000001e0),
    .I1(sig000001e1),
    .I2(sig00000215),
    .I3(sig00000214),
    .I4(sig0000023f),
    .I5(sig0000022e),
    .O(sig0000052c)
  );
  LUT6 #(
    .INIT ( 64'hF0F0FF00CCCCAAAA ))
  blk000005ea (
    .I0(sig000001da),
    .I1(sig000001db),
    .I2(sig0000020f),
    .I3(sig0000020e),
    .I4(sig0000023f),
    .I5(sig0000022e),
    .O(sig00000526)
  );
  LUT6 #(
    .INIT ( 64'hF0F0FF00CCCCAAAA ))
  blk000005eb (
    .I0(sig000001db),
    .I1(sig000001dc),
    .I2(sig00000210),
    .I3(sig0000020f),
    .I4(sig0000023f),
    .I5(sig0000022e),
    .O(sig00000527)
  );
  LUT6 #(
    .INIT ( 64'hF0F0FF00CCCCAAAA ))
  blk000005ec (
    .I0(sig000001d9),
    .I1(sig000001da),
    .I2(sig0000020e),
    .I3(sig0000020d),
    .I4(sig0000023f),
    .I5(sig0000022e),
    .O(sig00000525)
  );
  LUT6 #(
    .INIT ( 64'hF0F0FF00CCCCAAAA ))
  blk000005ed (
    .I0(sig000001df),
    .I1(sig000001e0),
    .I2(sig00000214),
    .I3(sig00000213),
    .I4(sig0000023f),
    .I5(sig0000022e),
    .O(sig0000052b)
  );
  LUT6 #(
    .INIT ( 64'hF0F0FF00CCCCAAAA ))
  blk000005ee (
    .I0(sig000001d8),
    .I1(sig000001d9),
    .I2(sig0000020d),
    .I3(sig0000020c),
    .I4(sig0000023f),
    .I5(sig0000022e),
    .O(sig00000524)
  );
  LUT6 #(
    .INIT ( 64'hF0F0FF00CCCCAAAA ))
  blk000005ef (
    .I0(sig000001d7),
    .I1(sig000001d8),
    .I2(sig0000020c),
    .I3(sig0000020b),
    .I4(sig0000023f),
    .I5(sig0000022e),
    .O(sig00000523)
  );
  LUT6 #(
    .INIT ( 64'hF0F0FF00CCCCAAAA ))
  blk000005f0 (
    .I0(sig000001d6),
    .I1(sig000001d7),
    .I2(sig0000020b),
    .I3(sig0000020a),
    .I4(sig0000023f),
    .I5(sig0000022e),
    .O(sig00000522)
  );
  LUT6 #(
    .INIT ( 64'hF0F0FF00CCCCAAAA ))
  blk000005f1 (
    .I0(sig000001d5),
    .I1(sig000001d6),
    .I2(sig0000020a),
    .I3(sig00000209),
    .I4(sig0000023f),
    .I5(sig0000022e),
    .O(sig00000521)
  );
  LUT6 #(
    .INIT ( 64'hF0F0FF00CCCCAAAA ))
  blk000005f2 (
    .I0(sig000001d4),
    .I1(sig000001d5),
    .I2(sig00000209),
    .I3(sig00000208),
    .I4(sig0000023f),
    .I5(sig0000022e),
    .O(sig00000520)
  );
  LUT6 #(
    .INIT ( 64'hF0F0FF00CCCCAAAA ))
  blk000005f3 (
    .I0(sig000001e5),
    .I1(sig000001e6),
    .I2(sig0000021a),
    .I3(sig00000219),
    .I4(sig0000023f),
    .I5(sig0000022e),
    .O(sig00000531)
  );
  LUT6 #(
    .INIT ( 64'hF0F0FF00CCCCAAAA ))
  blk000005f4 (
    .I0(sig000001d3),
    .I1(sig000001d4),
    .I2(sig00000208),
    .I3(sig00000207),
    .I4(sig0000023f),
    .I5(sig0000022e),
    .O(sig0000051f)
  );
  LUT6 #(
    .INIT ( 64'hF0F0FF00CCCCAAAA ))
  blk000005f5 (
    .I0(sig000001d2),
    .I1(sig000001d3),
    .I2(sig00000207),
    .I3(sig00000206),
    .I4(sig0000023f),
    .I5(sig0000022e),
    .O(sig0000051e)
  );
  LUT6 #(
    .INIT ( 64'hF0F0FF00CCCCAAAA ))
  blk000005f6 (
    .I0(sig000001d1),
    .I1(sig000001d2),
    .I2(sig00000206),
    .I3(sig00000205),
    .I4(sig0000023f),
    .I5(sig0000022e),
    .O(sig0000051d)
  );
  LUT6 #(
    .INIT ( 64'hF0F0FF00CCCCAAAA ))
  blk000005f7 (
    .I0(sig000001c3),
    .I1(sig000001c4),
    .I2(sig000001f8),
    .I3(sig000001f7),
    .I4(sig0000023f),
    .I5(sig0000022e),
    .O(sig0000050f)
  );
  LUT6 #(
    .INIT ( 64'hF0F0FF00CCCCAAAA ))
  blk000005f8 (
    .I0(sig000001c4),
    .I1(sig000001c5),
    .I2(sig000001f9),
    .I3(sig000001f8),
    .I4(sig0000023f),
    .I5(sig0000022e),
    .O(sig00000510)
  );
  LUT6 #(
    .INIT ( 64'hF0F0FF00CCCCAAAA ))
  blk000005f9 (
    .I0(sig000001d0),
    .I1(sig000001d1),
    .I2(sig00000205),
    .I3(sig00000204),
    .I4(sig0000023f),
    .I5(sig0000022e),
    .O(sig0000051c)
  );
  LUT6 #(
    .INIT ( 64'hF0F0FF00CCCCAAAA ))
  blk000005fa (
    .I0(sig000001de),
    .I1(sig000001df),
    .I2(sig00000213),
    .I3(sig00000212),
    .I4(sig0000023f),
    .I5(sig0000022e),
    .O(sig0000052a)
  );
  LUT6 #(
    .INIT ( 64'hF0F0FF00CCCCAAAA ))
  blk000005fb (
    .I0(sig000001cf),
    .I1(sig000001d0),
    .I2(sig00000204),
    .I3(sig00000203),
    .I4(sig0000023f),
    .I5(sig0000022e),
    .O(sig0000051b)
  );
  LUT6 #(
    .INIT ( 64'hF0F0FF00CCCCAAAA ))
  blk000005fc (
    .I0(sig000001ce),
    .I1(sig000001cf),
    .I2(sig00000203),
    .I3(sig00000202),
    .I4(sig0000023f),
    .I5(sig0000022e),
    .O(sig0000051a)
  );
  LUT6 #(
    .INIT ( 64'hF0F0FF00CCCCAAAA ))
  blk000005fd (
    .I0(sig000001cd),
    .I1(sig000001ce),
    .I2(sig00000202),
    .I3(sig00000201),
    .I4(sig0000023f),
    .I5(sig0000022e),
    .O(sig00000519)
  );
  LUT6 #(
    .INIT ( 64'hF0F0FF00CCCCAAAA ))
  blk000005fe (
    .I0(sig000001cc),
    .I1(sig000001cd),
    .I2(sig00000201),
    .I3(sig00000200),
    .I4(sig0000023f),
    .I5(sig0000022e),
    .O(sig00000518)
  );
  LUT6 #(
    .INIT ( 64'hF0F0FF00CCCCAAAA ))
  blk000005ff (
    .I0(sig000001c6),
    .I1(sig000001c7),
    .I2(sig000001fb),
    .I3(sig000001fa),
    .I4(sig0000023f),
    .I5(sig0000022e),
    .O(sig00000512)
  );
  LUT6 #(
    .INIT ( 64'hF0F0FF00CCCCAAAA ))
  blk00000600 (
    .I0(sig000001c5),
    .I1(sig000001c6),
    .I2(sig000001fa),
    .I3(sig000001f9),
    .I4(sig0000023f),
    .I5(sig0000022e),
    .O(sig00000511)
  );
  LUT6 #(
    .INIT ( 64'hF0F0FF00CCCCAAAA ))
  blk00000601 (
    .I0(sig000001cb),
    .I1(sig000001cc),
    .I2(sig00000200),
    .I3(sig000001ff),
    .I4(sig0000023f),
    .I5(sig0000022e),
    .O(sig00000517)
  );
  LUT6 #(
    .INIT ( 64'hF0F0FF00CCCCAAAA ))
  blk00000602 (
    .I0(sig000001ca),
    .I1(sig000001cb),
    .I2(sig000001ff),
    .I3(sig000001fe),
    .I4(sig0000023f),
    .I5(sig0000022e),
    .O(sig00000516)
  );
  LUT6 #(
    .INIT ( 64'hF0F0FF00CCCCAAAA ))
  blk00000603 (
    .I0(sig000001c9),
    .I1(sig000001ca),
    .I2(sig000001fe),
    .I3(sig000001fd),
    .I4(sig0000023f),
    .I5(sig0000022e),
    .O(sig00000515)
  );
  LUT6 #(
    .INIT ( 64'hF0F0FF00CCCCAAAA ))
  blk00000604 (
    .I0(sig000001c8),
    .I1(sig000001c9),
    .I2(sig000001fd),
    .I3(sig000001fc),
    .I4(sig0000023f),
    .I5(sig0000022e),
    .O(sig00000514)
  );
  LUT6 #(
    .INIT ( 64'hF0F0FF00CCCCAAAA ))
  blk00000605 (
    .I0(sig000001c7),
    .I1(sig000001c8),
    .I2(sig000001fc),
    .I3(sig000001fb),
    .I4(sig0000023f),
    .I5(sig0000022e),
    .O(sig00000513)
  );
  LUT6 #(
    .INIT ( 64'hF0F0FF00CCCCAAAA ))
  blk00000606 (
    .I0(sig000001f5),
    .I1(sig000001f6),
    .I2(sig0000022a),
    .I3(sig00000229),
    .I4(sig0000023f),
    .I5(sig0000022e),
    .O(sig00000541)
  );
  LUT6 #(
    .INIT ( 64'hF0F0FF00CCCCAAAA ))
  blk00000607 (
    .I0(sig000001dd),
    .I1(sig000001de),
    .I2(sig00000212),
    .I3(sig00000211),
    .I4(sig0000023f),
    .I5(sig0000022e),
    .O(sig00000529)
  );
  LUT6 #(
    .INIT ( 64'hF0F0FF00CCCCAAAA ))
  blk00000608 (
    .I0(sig000001f4),
    .I1(sig000001f5),
    .I2(sig00000229),
    .I3(sig00000228),
    .I4(sig0000023f),
    .I5(sig0000022e),
    .O(sig00000540)
  );
  LUT6 #(
    .INIT ( 64'hF0F0FF00CCCCAAAA ))
  blk00000609 (
    .I0(sig000001f3),
    .I1(sig000001f4),
    .I2(sig00000228),
    .I3(sig00000227),
    .I4(sig0000023f),
    .I5(sig0000022e),
    .O(sig0000053f)
  );
  LUT6 #(
    .INIT ( 64'hF0F0FF00CCCCAAAA ))
  blk0000060a (
    .I0(sig000001f2),
    .I1(sig000001f3),
    .I2(sig00000227),
    .I3(sig00000226),
    .I4(sig0000023f),
    .I5(sig0000022e),
    .O(sig0000053e)
  );
  LUT6 #(
    .INIT ( 64'hF0F0FF00CCCCAAAA ))
  blk0000060b (
    .I0(sig000001f1),
    .I1(sig000001f2),
    .I2(sig00000226),
    .I3(sig00000225),
    .I4(sig0000023f),
    .I5(sig0000022e),
    .O(sig0000053d)
  );
  LUT6 #(
    .INIT ( 64'hF0F0FF00CCCCAAAA ))
  blk0000060c (
    .I0(sig000001f0),
    .I1(sig000001f1),
    .I2(sig00000225),
    .I3(sig00000224),
    .I4(sig0000023f),
    .I5(sig0000022e),
    .O(sig0000053c)
  );
  LUT6 #(
    .INIT ( 64'hF0F0FF00CCCCAAAA ))
  blk0000060d (
    .I0(sig000001ef),
    .I1(sig000001f0),
    .I2(sig00000224),
    .I3(sig00000223),
    .I4(sig0000023f),
    .I5(sig0000022e),
    .O(sig0000053b)
  );
  LUT6 #(
    .INIT ( 64'hF0F0FF00CCCCAAAA ))
  blk0000060e (
    .I0(sig000001ee),
    .I1(sig000001ef),
    .I2(sig00000223),
    .I3(sig00000222),
    .I4(sig0000023f),
    .I5(sig0000022e),
    .O(sig0000053a)
  );
  LUT6 #(
    .INIT ( 64'hF0F0FF00CCCCAAAA ))
  blk0000060f (
    .I0(sig000001ed),
    .I1(sig000001ee),
    .I2(sig00000222),
    .I3(sig00000221),
    .I4(sig0000023f),
    .I5(sig0000022e),
    .O(sig00000539)
  );
  LUT6 #(
    .INIT ( 64'hF0F0FF00CCCCAAAA ))
  blk00000610 (
    .I0(sig000001dc),
    .I1(sig000001dd),
    .I2(sig00000211),
    .I3(sig00000210),
    .I4(sig0000023f),
    .I5(sig0000022e),
    .O(sig00000528)
  );
  LUT6 #(
    .INIT ( 64'hF0F0FF00CCCCAAAA ))
  blk00000611 (
    .I0(sig000001ec),
    .I1(sig000001ed),
    .I2(sig00000221),
    .I3(sig00000220),
    .I4(sig0000023f),
    .I5(sig0000022e),
    .O(sig00000538)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk00000612 (
    .I0(sig0000040e),
    .I1(sig0000040d),
    .I2(sig000003de),
    .I3(sig000003d6),
    .I4(sig000003da),
    .I5(sig000003e2),
    .O(sig00000452)
  );
  LUT4 #(
    .INIT ( 16'h5410 ))
  blk00000613 (
    .I0(sig0000040d),
    .I1(sig0000040e),
    .I2(sig000003da),
    .I3(sig000003d6),
    .O(sig0000044a)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk00000614 (
    .I0(sig0000040e),
    .I1(sig0000040d),
    .I2(sig000003df),
    .I3(sig000003d7),
    .I4(sig000003db),
    .I5(sig000003e3),
    .O(sig00000453)
  );
  LUT4 #(
    .INIT ( 16'h5410 ))
  blk00000615 (
    .I0(sig0000040d),
    .I1(sig0000040e),
    .I2(sig000003db),
    .I3(sig000003d7),
    .O(sig0000044b)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk00000616 (
    .I0(sig0000040e),
    .I1(sig0000040d),
    .I2(sig000003e0),
    .I3(sig000003d8),
    .I4(sig000003dc),
    .I5(sig000003e4),
    .O(sig00000454)
  );
  LUT4 #(
    .INIT ( 16'h5410 ))
  blk00000617 (
    .I0(sig0000040d),
    .I1(sig0000040e),
    .I2(sig000003dc),
    .I3(sig000003d8),
    .O(sig0000044c)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk00000618 (
    .I0(sig0000040e),
    .I1(sig0000040d),
    .I2(sig000003e1),
    .I3(sig000003d9),
    .I4(sig000003dd),
    .I5(sig000003e5),
    .O(sig00000455)
  );
  LUT4 #(
    .INIT ( 16'h5410 ))
  blk00000619 (
    .I0(sig0000040d),
    .I1(sig0000040e),
    .I2(sig000003dd),
    .I3(sig000003d9),
    .O(sig0000044d)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk0000061a (
    .I0(sig0000040e),
    .I1(sig0000040d),
    .I2(sig000003e5),
    .I3(sig000003dd),
    .I4(sig000003e1),
    .I5(sig000003e9),
    .O(sig00000459)
  );
  LUT5 #(
    .INIT ( 32'h73625140 ))
  blk0000061b (
    .I0(sig0000040d),
    .I1(sig0000040e),
    .I2(sig000003dd),
    .I3(sig000003e1),
    .I4(sig000003d9),
    .O(sig00000451)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk0000061c (
    .I0(sig0000040e),
    .I1(sig0000040d),
    .I2(sig000003e6),
    .I3(sig000003de),
    .I4(sig000003e2),
    .I5(sig000003ea),
    .O(sig0000045a)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk0000061d (
    .I0(sig0000040e),
    .I1(sig0000040d),
    .I2(sig000003e7),
    .I3(sig000003df),
    .I4(sig000003e3),
    .I5(sig000003eb),
    .O(sig0000045b)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk0000061e (
    .I0(sig0000040e),
    .I1(sig0000040d),
    .I2(sig000003e8),
    .I3(sig000003e0),
    .I4(sig000003e4),
    .I5(sig000003ec),
    .O(sig0000045c)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk0000061f (
    .I0(sig0000040e),
    .I1(sig0000040d),
    .I2(sig000003e9),
    .I3(sig000003e1),
    .I4(sig000003e5),
    .I5(sig000003ed),
    .O(sig0000045d)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk00000620 (
    .I0(sig0000040e),
    .I1(sig0000040d),
    .I2(sig000003ee),
    .I3(sig000003e6),
    .I4(sig000003ea),
    .I5(sig000003f2),
    .O(sig00000462)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk00000621 (
    .I0(sig0000040e),
    .I1(sig0000040d),
    .I2(sig000003ef),
    .I3(sig000003e7),
    .I4(sig000003eb),
    .I5(sig000003f3),
    .O(sig00000463)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk00000622 (
    .I0(sig0000040e),
    .I1(sig0000040d),
    .I2(sig000003e2),
    .I3(sig000003da),
    .I4(sig000003de),
    .I5(sig000003e6),
    .O(sig00000456)
  );
  LUT5 #(
    .INIT ( 32'h73625140 ))
  blk00000623 (
    .I0(sig0000040d),
    .I1(sig0000040e),
    .I2(sig000003da),
    .I3(sig000003de),
    .I4(sig000003d6),
    .O(sig0000044e)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk00000624 (
    .I0(sig0000040e),
    .I1(sig0000040d),
    .I2(sig000003f0),
    .I3(sig000003e8),
    .I4(sig000003ec),
    .I5(sig000003f4),
    .O(sig00000464)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk00000625 (
    .I0(sig0000040e),
    .I1(sig0000040d),
    .I2(sig000003f1),
    .I3(sig000003e9),
    .I4(sig000003ed),
    .I5(sig000003f5),
    .O(sig00000465)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk00000626 (
    .I0(sig0000040e),
    .I1(sig0000040d),
    .I2(sig000003ea),
    .I3(sig000003e2),
    .I4(sig000003e6),
    .I5(sig000003ee),
    .O(sig0000045e)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk00000627 (
    .I0(sig0000040e),
    .I1(sig0000040d),
    .I2(sig000003f2),
    .I3(sig000003ea),
    .I4(sig000003ee),
    .I5(sig000003f6),
    .O(sig00000466)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk00000628 (
    .I0(sig0000040e),
    .I1(sig0000040d),
    .I2(sig000003f3),
    .I3(sig000003eb),
    .I4(sig000003ef),
    .I5(sig000003f7),
    .O(sig00000467)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk00000629 (
    .I0(sig0000040e),
    .I1(sig0000040d),
    .I2(sig000003eb),
    .I3(sig000003e3),
    .I4(sig000003e7),
    .I5(sig000003ef),
    .O(sig0000045f)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk0000062a (
    .I0(sig0000040e),
    .I1(sig0000040d),
    .I2(sig000003f4),
    .I3(sig000003ec),
    .I4(sig000003f0),
    .I5(sig000003f8),
    .O(sig00000468)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk0000062b (
    .I0(sig0000040e),
    .I1(sig0000040d),
    .I2(sig000003ec),
    .I3(sig000003e4),
    .I4(sig000003e8),
    .I5(sig000003f0),
    .O(sig00000460)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk0000062c (
    .I0(sig0000040e),
    .I1(sig0000040d),
    .I2(sig000003f5),
    .I3(sig000003ed),
    .I4(sig000003f1),
    .I5(sig000003f9),
    .O(sig00000469)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk0000062d (
    .I0(sig0000040e),
    .I1(sig0000040d),
    .I2(sig000003ed),
    .I3(sig000003e5),
    .I4(sig000003e9),
    .I5(sig000003f1),
    .O(sig00000461)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk0000062e (
    .I0(sig0000040e),
    .I1(sig0000040d),
    .I2(sig000003f6),
    .I3(sig000003ee),
    .I4(sig000003f2),
    .I5(sig000003fa),
    .O(sig0000046a)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk0000062f (
    .I0(sig0000040e),
    .I1(sig0000040d),
    .I2(sig000003f7),
    .I3(sig000003ef),
    .I4(sig000003f3),
    .I5(sig000003fb),
    .O(sig0000046b)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk00000630 (
    .I0(sig0000040e),
    .I1(sig0000040d),
    .I2(sig000003f8),
    .I3(sig000003f0),
    .I4(sig000003f4),
    .I5(sig000003fc),
    .O(sig0000046c)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk00000631 (
    .I0(sig0000040e),
    .I1(sig0000040d),
    .I2(sig000003e3),
    .I3(sig000003db),
    .I4(sig000003df),
    .I5(sig000003e7),
    .O(sig00000457)
  );
  LUT5 #(
    .INIT ( 32'h73625140 ))
  blk00000632 (
    .I0(sig0000040d),
    .I1(sig0000040e),
    .I2(sig000003db),
    .I3(sig000003df),
    .I4(sig000003d7),
    .O(sig0000044f)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk00000633 (
    .I0(sig0000040e),
    .I1(sig0000040d),
    .I2(sig000003f9),
    .I3(sig000003f1),
    .I4(sig000003f5),
    .I5(sig000003fd),
    .O(sig0000046d)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk00000634 (
    .I0(sig0000040e),
    .I1(sig0000040d),
    .I2(sig000003fa),
    .I3(sig000003f2),
    .I4(sig000003f6),
    .I5(sig000003fe),
    .O(sig0000046e)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk00000635 (
    .I0(sig0000040e),
    .I1(sig0000040d),
    .I2(sig000003fb),
    .I3(sig000003f3),
    .I4(sig000003f7),
    .I5(sig000003ff),
    .O(sig0000046f)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk00000636 (
    .I0(sig0000040e),
    .I1(sig0000040d),
    .I2(sig000003fc),
    .I3(sig000003f4),
    .I4(sig000003f8),
    .I5(sig00000400),
    .O(sig00000470)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk00000637 (
    .I0(sig0000040e),
    .I1(sig0000040d),
    .I2(sig000003fd),
    .I3(sig000003f5),
    .I4(sig000003f9),
    .I5(sig00000401),
    .O(sig00000471)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk00000638 (
    .I0(sig0000040e),
    .I1(sig0000040d),
    .I2(sig000003fe),
    .I3(sig000003f6),
    .I4(sig000003fa),
    .I5(sig00000402),
    .O(sig00000472)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk00000639 (
    .I0(sig0000040e),
    .I1(sig0000040d),
    .I2(sig000003ff),
    .I3(sig000003f7),
    .I4(sig000003fb),
    .I5(sig00000403),
    .O(sig00000473)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk0000063a (
    .I0(sig0000040e),
    .I1(sig0000040d),
    .I2(sig00000407),
    .I3(sig000003ff),
    .I4(sig00000403),
    .I5(sig0000040b),
    .O(sig0000047b)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk0000063b (
    .I0(sig0000040e),
    .I1(sig0000040d),
    .I2(sig00000400),
    .I3(sig000003f8),
    .I4(sig000003fc),
    .I5(sig00000404),
    .O(sig00000474)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk0000063c (
    .I0(sig0000040e),
    .I1(sig0000040d),
    .I2(sig00000401),
    .I3(sig000003f9),
    .I4(sig000003fd),
    .I5(sig00000405),
    .O(sig00000475)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk0000063d (
    .I0(sig0000040e),
    .I1(sig0000040d),
    .I2(sig000003e4),
    .I3(sig000003dc),
    .I4(sig000003e0),
    .I5(sig000003e8),
    .O(sig00000458)
  );
  LUT5 #(
    .INIT ( 32'h73625140 ))
  blk0000063e (
    .I0(sig0000040d),
    .I1(sig0000040e),
    .I2(sig000003dc),
    .I3(sig000003e0),
    .I4(sig000003d8),
    .O(sig00000450)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk0000063f (
    .I0(sig0000040e),
    .I1(sig0000040d),
    .I2(sig00000408),
    .I3(sig00000400),
    .I4(sig00000404),
    .I5(sig0000040c),
    .O(sig0000047c)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk00000640 (
    .I0(sig0000040e),
    .I1(sig0000040d),
    .I2(sig00000402),
    .I3(sig000003fa),
    .I4(sig000003fe),
    .I5(sig00000406),
    .O(sig00000476)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk00000641 (
    .I0(sig0000040e),
    .I1(sig0000040d),
    .I2(sig00000403),
    .I3(sig000003fb),
    .I4(sig000003ff),
    .I5(sig00000407),
    .O(sig00000477)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk00000642 (
    .I0(sig0000040e),
    .I1(sig0000040d),
    .I2(sig00000404),
    .I3(sig000003fc),
    .I4(sig00000400),
    .I5(sig00000408),
    .O(sig00000478)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk00000643 (
    .I0(sig0000040e),
    .I1(sig0000040d),
    .I2(sig00000405),
    .I3(sig000003fd),
    .I4(sig00000401),
    .I5(sig00000409),
    .O(sig00000479)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk00000644 (
    .I0(sig0000040e),
    .I1(sig0000040d),
    .I2(sig00000406),
    .I3(sig000003fe),
    .I4(sig00000402),
    .I5(sig0000040a),
    .O(sig0000047a)
  );
  LUT5 #(
    .INIT ( 32'h73625140 ))
  blk00000645 (
    .I0(sig000003d4),
    .I1(sig000003d5),
    .I2(sig000004f0),
    .I3(sig000004e0),
    .I4(sig00000500),
    .O(sig0000043b)
  );
  LUT5 #(
    .INIT ( 32'h73625140 ))
  blk00000646 (
    .I0(sig000003d4),
    .I1(sig000003d5),
    .I2(sig000004f1),
    .I3(sig000004e1),
    .I4(sig00000501),
    .O(sig0000043a)
  );
  LUT5 #(
    .INIT ( 32'h73625140 ))
  blk00000647 (
    .I0(sig000003d4),
    .I1(sig000003d5),
    .I2(sig000004f2),
    .I3(sig000004e2),
    .I4(sig00000502),
    .O(sig00000439)
  );
  LUT5 #(
    .INIT ( 32'h73625140 ))
  blk00000648 (
    .I0(sig000003d4),
    .I1(sig000003d5),
    .I2(sig000004f3),
    .I3(sig000004e3),
    .I4(sig00000503),
    .O(sig00000438)
  );
  LUT5 #(
    .INIT ( 32'h73625140 ))
  blk00000649 (
    .I0(sig000003d4),
    .I1(sig000003d5),
    .I2(sig000004f4),
    .I3(sig000004e4),
    .I4(sig00000504),
    .O(sig00000437)
  );
  LUT5 #(
    .INIT ( 32'h73625140 ))
  blk0000064a (
    .I0(sig000003d4),
    .I1(sig000003d5),
    .I2(sig000004f5),
    .I3(sig000004e5),
    .I4(sig00000505),
    .O(sig00000436)
  );
  LUT5 #(
    .INIT ( 32'h73625140 ))
  blk0000064b (
    .I0(sig000003d4),
    .I1(sig000003d5),
    .I2(sig000004f6),
    .I3(sig000004e6),
    .I4(sig00000506),
    .O(sig00000435)
  );
  LUT5 #(
    .INIT ( 32'h73625140 ))
  blk0000064c (
    .I0(sig000003d4),
    .I1(sig000003d5),
    .I2(sig000004f7),
    .I3(sig000004e7),
    .I4(sig00000507),
    .O(sig00000434)
  );
  LUT5 #(
    .INIT ( 32'h73625140 ))
  blk0000064d (
    .I0(sig000003d4),
    .I1(sig000003d5),
    .I2(sig000004f8),
    .I3(sig000004e8),
    .I4(sig00000508),
    .O(sig00000433)
  );
  LUT5 #(
    .INIT ( 32'h73625140 ))
  blk0000064e (
    .I0(sig000003d4),
    .I1(sig000003d5),
    .I2(sig000004f9),
    .I3(sig000004e9),
    .I4(sig00000509),
    .O(sig00000432)
  );
  LUT5 #(
    .INIT ( 32'h73625140 ))
  blk0000064f (
    .I0(sig000003d4),
    .I1(sig000003d5),
    .I2(sig000004fa),
    .I3(sig000004ea),
    .I4(sig0000050a),
    .O(sig00000431)
  );
  LUT5 #(
    .INIT ( 32'h73625140 ))
  blk00000650 (
    .I0(sig000003d4),
    .I1(sig000003d5),
    .I2(sig000004fb),
    .I3(sig000004eb),
    .I4(sig0000050b),
    .O(sig00000430)
  );
  LUT5 #(
    .INIT ( 32'h73625140 ))
  blk00000651 (
    .I0(sig000003d4),
    .I1(sig000003d5),
    .I2(sig000004fc),
    .I3(sig000004ec),
    .I4(sig0000050c),
    .O(sig0000042f)
  );
  LUT4 #(
    .INIT ( 16'h5410 ))
  blk00000652 (
    .I0(sig000003d4),
    .I1(sig000003d5),
    .I2(sig000004ed),
    .I3(sig000004fd),
    .O(sig0000042e)
  );
  LUT4 #(
    .INIT ( 16'h5410 ))
  blk00000653 (
    .I0(sig000003d4),
    .I1(sig000003d5),
    .I2(sig000004ee),
    .I3(sig000004fe),
    .O(sig0000042d)
  );
  LUT4 #(
    .INIT ( 16'h5410 ))
  blk00000654 (
    .I0(sig000003d4),
    .I1(sig000003d5),
    .I2(sig000004ef),
    .I3(sig000004ff),
    .O(sig0000042c)
  );
  LUT4 #(
    .INIT ( 16'h5410 ))
  blk00000655 (
    .I0(sig000003d4),
    .I1(sig000003d5),
    .I2(sig000004f0),
    .I3(sig00000500),
    .O(sig0000042b)
  );
  LUT4 #(
    .INIT ( 16'h5410 ))
  blk00000656 (
    .I0(sig000003d4),
    .I1(sig000003d5),
    .I2(sig000004f1),
    .I3(sig00000501),
    .O(sig0000042a)
  );
  LUT4 #(
    .INIT ( 16'h5410 ))
  blk00000657 (
    .I0(sig000003d4),
    .I1(sig000003d5),
    .I2(sig000004f2),
    .I3(sig00000502),
    .O(sig00000429)
  );
  LUT4 #(
    .INIT ( 16'h5410 ))
  blk00000658 (
    .I0(sig000003d4),
    .I1(sig000003d5),
    .I2(sig000004f3),
    .I3(sig00000503),
    .O(sig00000428)
  );
  LUT4 #(
    .INIT ( 16'h5410 ))
  blk00000659 (
    .I0(sig000003d4),
    .I1(sig000003d5),
    .I2(sig000004f4),
    .I3(sig00000504),
    .O(sig00000427)
  );
  LUT4 #(
    .INIT ( 16'h5410 ))
  blk0000065a (
    .I0(sig000003d4),
    .I1(sig000003d5),
    .I2(sig000004f5),
    .I3(sig00000505),
    .O(sig00000426)
  );
  LUT5 #(
    .INIT ( 32'h73625140 ))
  blk0000065b (
    .I0(sig000003d4),
    .I1(sig000003d5),
    .I2(sig000004ed),
    .I3(sig000004dd),
    .I4(sig000004fd),
    .O(sig0000043e)
  );
  LUT5 #(
    .INIT ( 32'h73625140 ))
  blk0000065c (
    .I0(sig000003d4),
    .I1(sig000003d5),
    .I2(sig000004ee),
    .I3(sig000004de),
    .I4(sig000004fe),
    .O(sig0000043d)
  );
  LUT5 #(
    .INIT ( 32'h73625140 ))
  blk0000065d (
    .I0(sig000003d4),
    .I1(sig000003d5),
    .I2(sig000004ef),
    .I3(sig000004df),
    .I4(sig000004ff),
    .O(sig0000043c)
  );
  LUT3 #(
    .INIT ( 8'h10 ))
  blk0000065e (
    .I0(sig0000040d),
    .I1(sig0000040e),
    .I2(sig000003d9),
    .O(sig00000449)
  );
  LUT3 #(
    .INIT ( 8'h10 ))
  blk0000065f (
    .I0(sig0000040d),
    .I1(sig0000040e),
    .I2(sig000003d8),
    .O(sig00000448)
  );
  LUT3 #(
    .INIT ( 8'h10 ))
  blk00000660 (
    .I0(sig0000040d),
    .I1(sig0000040e),
    .I2(sig000003d7),
    .O(sig00000447)
  );
  LUT3 #(
    .INIT ( 8'h10 ))
  blk00000661 (
    .I0(sig0000040d),
    .I1(sig0000040e),
    .I2(sig000003d6),
    .O(sig00000446)
  );
  LUT3 #(
    .INIT ( 8'h10 ))
  blk00000662 (
    .I0(sig000003d4),
    .I1(sig000003d5),
    .I2(sig000004fd),
    .O(sig0000041e)
  );
  LUT3 #(
    .INIT ( 8'h10 ))
  blk00000663 (
    .I0(sig000003d4),
    .I1(sig000003d5),
    .I2(sig000004fe),
    .O(sig0000041d)
  );
  LUT3 #(
    .INIT ( 8'h10 ))
  blk00000664 (
    .I0(sig000003d4),
    .I1(sig000003d5),
    .I2(sig000004ff),
    .O(sig0000041c)
  );
  LUT3 #(
    .INIT ( 8'h10 ))
  blk00000665 (
    .I0(sig000003d4),
    .I1(sig000003d5),
    .I2(sig00000500),
    .O(sig0000041b)
  );
  LUT3 #(
    .INIT ( 8'h10 ))
  blk00000666 (
    .I0(sig000003d4),
    .I1(sig000003d5),
    .I2(sig00000501),
    .O(sig0000041a)
  );
  LUT3 #(
    .INIT ( 8'h10 ))
  blk00000667 (
    .I0(sig000003d4),
    .I1(sig000003d5),
    .I2(sig00000502),
    .O(sig00000419)
  );
  LUT3 #(
    .INIT ( 8'h10 ))
  blk00000668 (
    .I0(sig000003d4),
    .I1(sig000003d5),
    .I2(sig00000503),
    .O(sig00000418)
  );
  LUT3 #(
    .INIT ( 8'h10 ))
  blk00000669 (
    .I0(sig000003d4),
    .I1(sig000003d5),
    .I2(sig00000504),
    .O(sig00000417)
  );
  LUT3 #(
    .INIT ( 8'h10 ))
  blk0000066a (
    .I0(sig000003d4),
    .I1(sig000003d5),
    .I2(sig00000505),
    .O(sig00000416)
  );
  LUT3 #(
    .INIT ( 8'h10 ))
  blk0000066b (
    .I0(sig000003d4),
    .I1(sig000003d5),
    .I2(sig00000506),
    .O(sig00000415)
  );
  LUT3 #(
    .INIT ( 8'h10 ))
  blk0000066c (
    .I0(sig000003d4),
    .I1(sig000003d5),
    .I2(sig00000507),
    .O(sig00000414)
  );
  LUT3 #(
    .INIT ( 8'h10 ))
  blk0000066d (
    .I0(sig000003d4),
    .I1(sig000003d5),
    .I2(sig00000508),
    .O(sig00000413)
  );
  LUT3 #(
    .INIT ( 8'h10 ))
  blk0000066e (
    .I0(sig000003d4),
    .I1(sig000003d5),
    .I2(sig00000509),
    .O(sig00000412)
  );
  LUT3 #(
    .INIT ( 8'h10 ))
  blk0000066f (
    .I0(sig000003d4),
    .I1(sig000003d5),
    .I2(sig0000050a),
    .O(sig00000411)
  );
  LUT3 #(
    .INIT ( 8'h10 ))
  blk00000670 (
    .I0(sig000003d4),
    .I1(sig000003d5),
    .I2(sig0000050b),
    .O(sig00000410)
  );
  LUT3 #(
    .INIT ( 8'h10 ))
  blk00000671 (
    .I0(sig000003d4),
    .I1(sig000003d5),
    .I2(sig0000050c),
    .O(sig0000040f)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000672 (
    .I0(sig00000249),
    .I1(sig0000024a),
    .O(sig00000583)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000673 (
    .I0(sig00000240),
    .I1(sig0000024a),
    .O(sig0000057a)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000674 (
    .I0(sig00000241),
    .I1(sig0000024a),
    .O(sig0000057b)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000675 (
    .I0(sig00000242),
    .I1(sig0000024a),
    .O(sig0000057c)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000676 (
    .I0(sig00000243),
    .I1(sig0000024a),
    .O(sig0000057d)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000677 (
    .I0(sig00000244),
    .I1(sig0000024a),
    .O(sig0000057e)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000678 (
    .I0(sig00000245),
    .I1(sig0000024a),
    .O(sig0000057f)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000679 (
    .I0(sig00000246),
    .I1(sig0000024a),
    .O(sig00000580)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk0000067a (
    .I0(sig00000247),
    .I1(sig0000024a),
    .O(sig00000581)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk0000067b (
    .I0(sig00000248),
    .I1(sig0000024a),
    .O(sig00000582)
  );
  LUT2 #(
    .INIT ( 4'hE ))
  blk0000067c (
    .I0(sig000004cd),
    .I1(sig00000544),
    .O(sig000004bb)
  );
  LUT3 #(
    .INIT ( 8'h1F ))
  blk0000067d (
    .I0(sig0000050b),
    .I1(sig0000050a),
    .I2(sig000004cf),
    .O(sig00000587)
  );
  LUT3 #(
    .INIT ( 8'h1F ))
  blk0000067e (
    .I0(sig00000507),
    .I1(sig00000506),
    .I2(sig000004cf),
    .O(sig00000588)
  );
  LUT3 #(
    .INIT ( 8'h1F ))
  blk0000067f (
    .I0(sig000004ff),
    .I1(sig000004fe),
    .I2(sig000004cf),
    .O(sig0000058a)
  );
  LUT3 #(
    .INIT ( 8'h1F ))
  blk00000680 (
    .I0(sig000004fb),
    .I1(sig000004fa),
    .I2(sig000004cf),
    .O(sig0000058b)
  );
  LUT3 #(
    .INIT ( 8'h1F ))
  blk00000681 (
    .I0(sig00000503),
    .I1(sig00000502),
    .I2(sig000004cf),
    .O(sig00000589)
  );
  LUT3 #(
    .INIT ( 8'h1F ))
  blk00000682 (
    .I0(sig000004f3),
    .I1(sig000004f2),
    .I2(sig000004cf),
    .O(sig0000058d)
  );
  LUT3 #(
    .INIT ( 8'h1F ))
  blk00000683 (
    .I0(sig000004ef),
    .I1(sig000004ee),
    .I2(sig000004cf),
    .O(sig0000058e)
  );
  LUT3 #(
    .INIT ( 8'h1F ))
  blk00000684 (
    .I0(sig000004f7),
    .I1(sig000004f6),
    .I2(sig000004cf),
    .O(sig0000058c)
  );
  LUT3 #(
    .INIT ( 8'h1F ))
  blk00000685 (
    .I0(sig000004e7),
    .I1(sig000004e6),
    .I2(sig000004cf),
    .O(sig00000590)
  );
  LUT3 #(
    .INIT ( 8'h1F ))
  blk00000686 (
    .I0(sig000004e3),
    .I1(sig000004e2),
    .I2(sig000004cf),
    .O(sig00000591)
  );
  LUT3 #(
    .INIT ( 8'h1F ))
  blk00000687 (
    .I0(sig000004eb),
    .I1(sig000004ea),
    .I2(sig000004cf),
    .O(sig0000058f)
  );
  LUT3 #(
    .INIT ( 8'h1F ))
  blk00000688 (
    .I0(sig000004db),
    .I1(sig000004da),
    .I2(sig000004cf),
    .O(sig00000593)
  );
  LUT2 #(
    .INIT ( 4'h7 ))
  blk00000689 (
    .I0(sig000004cf),
    .I1(sig000004d7),
    .O(sig00000594)
  );
  LUT3 #(
    .INIT ( 8'h1F ))
  blk0000068a (
    .I0(sig000004df),
    .I1(sig000004de),
    .I2(sig000004cf),
    .O(sig00000592)
  );
  LUT3 #(
    .INIT ( 8'h01 ))
  blk0000068b (
    .I0(sig0000050a),
    .I1(sig0000050b),
    .I2(sig0000050c),
    .O(sig000005b7)
  );
  LUT4 #(
    .INIT ( 16'h0001 ))
  blk0000068c (
    .I0(sig00000506),
    .I1(sig00000507),
    .I2(sig00000508),
    .I3(sig00000509),
    .O(sig000005b8)
  );
  LUT4 #(
    .INIT ( 16'h0001 ))
  blk0000068d (
    .I0(sig00000502),
    .I1(sig00000503),
    .I2(sig00000504),
    .I3(sig00000505),
    .O(sig000005b9)
  );
  LUT4 #(
    .INIT ( 16'h0001 ))
  blk0000068e (
    .I0(sig000004fe),
    .I1(sig000004ff),
    .I2(sig00000500),
    .I3(sig00000501),
    .O(sig000005ba)
  );
  LUT4 #(
    .INIT ( 16'h0001 ))
  blk0000068f (
    .I0(sig000004fa),
    .I1(sig000004fb),
    .I2(sig000004fc),
    .I3(sig000004fd),
    .O(sig000005bb)
  );
  LUT4 #(
    .INIT ( 16'h0001 ))
  blk00000690 (
    .I0(sig000004f6),
    .I1(sig000004f7),
    .I2(sig000004f8),
    .I3(sig000004f9),
    .O(sig000005bc)
  );
  LUT4 #(
    .INIT ( 16'h0001 ))
  blk00000691 (
    .I0(sig000004f2),
    .I1(sig000004f3),
    .I2(sig000004f4),
    .I3(sig000004f5),
    .O(sig000005bd)
  );
  LUT4 #(
    .INIT ( 16'h0001 ))
  blk00000692 (
    .I0(sig000004ee),
    .I1(sig000004ef),
    .I2(sig000004f0),
    .I3(sig000004f1),
    .O(sig000005be)
  );
  LUT4 #(
    .INIT ( 16'h0001 ))
  blk00000693 (
    .I0(sig000004ea),
    .I1(sig000004eb),
    .I2(sig000004ec),
    .I3(sig000004ed),
    .O(sig000005bf)
  );
  LUT4 #(
    .INIT ( 16'h0001 ))
  blk00000694 (
    .I0(sig000004e6),
    .I1(sig000004e7),
    .I2(sig000004e8),
    .I3(sig000004e9),
    .O(sig000005c0)
  );
  LUT4 #(
    .INIT ( 16'h0001 ))
  blk00000695 (
    .I0(sig000004e2),
    .I1(sig000004e3),
    .I2(sig000004e4),
    .I3(sig000004e5),
    .O(sig000005c1)
  );
  LUT4 #(
    .INIT ( 16'h0001 ))
  blk00000696 (
    .I0(sig000004de),
    .I1(sig000004df),
    .I2(sig000004e0),
    .I3(sig000004e1),
    .O(sig000005c2)
  );
  LUT4 #(
    .INIT ( 16'h0001 ))
  blk00000697 (
    .I0(sig000004da),
    .I1(sig000004db),
    .I2(sig000004dc),
    .I3(sig000004dd),
    .O(sig000005c3)
  );
  LUT3 #(
    .INIT ( 8'h01 ))
  blk00000698 (
    .I0(sig000004d7),
    .I1(sig000004d8),
    .I2(sig000004d9),
    .O(sig000005c4)
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  blk00000699 (
    .I0(sig00000696),
    .I1(sig00000697),
    .O(sig000005dc)
  );
  LUT6 #(
    .INIT ( 64'hCCCCCCCCC3993C66 ))
  blk0000069a (
    .I0(sig000005f9),
    .I1(sig00000601),
    .I2(sig000005fb),
    .I3(sig000005f8),
    .I4(sig00000696),
    .I5(sig00000697),
    .O(sig000005d4)
  );
  LUT6 #(
    .INIT ( 64'hCCCCCCCCC3993C66 ))
  blk0000069b (
    .I0(sig000005fa),
    .I1(sig00000602),
    .I2(sig000005fc),
    .I3(sig000005f8),
    .I4(sig00000696),
    .I5(sig00000697),
    .O(sig000005d5)
  );
  LUT6 #(
    .INIT ( 64'hAAAAAAAAA5995A66 ))
  blk0000069c (
    .I0(sig00000603),
    .I1(sig000005fb),
    .I2(sig000005fd),
    .I3(sig000005f8),
    .I4(sig00000696),
    .I5(sig00000697),
    .O(sig000005d6)
  );
  LUT6 #(
    .INIT ( 64'hAAAAAAAAA5995A66 ))
  blk0000069d (
    .I0(sig00000604),
    .I1(sig000005fc),
    .I2(sig000005fe),
    .I3(sig000005f8),
    .I4(sig00000696),
    .I5(sig00000697),
    .O(sig000005d7)
  );
  LUT6 #(
    .INIT ( 64'hAAAAAAAAA5995A66 ))
  blk0000069e (
    .I0(sig00000605),
    .I1(sig000005fd),
    .I2(sig000005ff),
    .I3(sig000005f8),
    .I4(sig00000696),
    .I5(sig00000697),
    .O(sig000005d8)
  );
  LUT6 #(
    .INIT ( 64'hAAAAAAAAA5995A66 ))
  blk0000069f (
    .I0(sig00000606),
    .I1(sig000005fe),
    .I2(sig00000600),
    .I3(sig000005f8),
    .I4(sig00000696),
    .I5(sig00000697),
    .O(sig000005d9)
  );
  LUT5 #(
    .INIT ( 32'hAAAA59A6 ))
  blk000006a0 (
    .I0(sig00000607),
    .I1(sig000005ff),
    .I2(sig000005f8),
    .I3(sig00000696),
    .I4(sig00000697),
    .O(sig000005da)
  );
  LUT5 #(
    .INIT ( 32'hAAAA59A6 ))
  blk000006a1 (
    .I0(sig00000608),
    .I1(sig00000600),
    .I2(sig000005f8),
    .I3(sig00000696),
    .I4(sig00000697),
    .O(sig000005db)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk000006a2 (
    .I0(sig00000666),
    .I1(sig000005e6),
    .I2(sig000005ef),
    .O(sig000005dd)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk000006a3 (
    .I0(sig00000666),
    .I1(sig000005e7),
    .I2(sig000005f0),
    .O(sig000005de)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk000006a4 (
    .I0(sig00000666),
    .I1(sig000005e8),
    .I2(sig000005f1),
    .O(sig000005df)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk000006a5 (
    .I0(sig00000666),
    .I1(sig000005e9),
    .I2(sig000005f2),
    .O(sig000005e0)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk000006a6 (
    .I0(sig00000666),
    .I1(sig000005ea),
    .I2(sig000005f3),
    .O(sig000005e1)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk000006a7 (
    .I0(sig00000666),
    .I1(sig000005eb),
    .I2(sig000005f4),
    .O(sig000005e2)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk000006a8 (
    .I0(sig00000666),
    .I1(sig000005ec),
    .I2(sig000005f5),
    .O(sig000005e3)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk000006a9 (
    .I0(sig00000666),
    .I1(sig000005ed),
    .I2(sig000005f6),
    .O(sig000005e4)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk000006aa (
    .I0(sig00000666),
    .I1(sig000005ee),
    .I2(sig000005f7),
    .O(sig000005e5)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk000006ab (
    .I0(sig000006e4),
    .I1(sig000006e9),
    .I2(sig000006eb),
    .O(sig000006c4)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk000006ac (
    .I0(sig000006e4),
    .I1(sig000006ea),
    .I2(sig000006ec),
    .O(sig000006c5)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk000006ad (
    .I0(sig000006e3),
    .I1(sig000006e5),
    .I2(sig000006e7),
    .O(sig000006c6)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk000006ae (
    .I0(sig000006e3),
    .I1(sig000006e6),
    .I2(sig000006e8),
    .O(sig000006c7)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk000006af (
    .I0(sig000006f9),
    .I1(sig000006f3),
    .I2(sig000006f6),
    .O(sig000006ca)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk000006b0 (
    .I0(sig000006f9),
    .I1(sig000006f4),
    .I2(sig000006f7),
    .O(sig000006cb)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk000006b1 (
    .I0(sig000006f9),
    .I1(sig000006f5),
    .I2(sig000006f8),
    .O(sig000006cc)
  );
  LUT2 #(
    .INIT ( 4'h8 ))
  blk000006b2 (
    .I0(sig000006f9),
    .I1(sig00000118),
    .O(sig000006cd)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk000006b3 (
    .I0(sig000006f1),
    .I1(sig000006ed),
    .I2(sig000006ee),
    .O(sig000006ce)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk000006b4 (
    .I0(sig000006f1),
    .I1(sig000006f2),
    .I2(sig000006ef),
    .O(sig000006cf)
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  blk000006b5 (
    .I0(sig000006f0),
    .I1(sig000006f1),
    .O(sig000006d0)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk000006b6 (
    .I0(sig00000118),
    .I1(sig000006f1),
    .I2(sig000006f9),
    .O(sig00000119)
  );
  LUT3 #(
    .INIT ( 8'hAC ))
  blk000006b7 (
    .I0(sig000006e3),
    .I1(sig000006e4),
    .I2(sig0000011a),
    .O(sig0000011b)
  );
  LUT2 #(
    .INIT ( 4'h8 ))
  blk000006b8 (
    .I0(sig0000011a),
    .I1(sig000006e4),
    .O(sig000006c2)
  );
  LUT2 #(
    .INIT ( 4'h8 ))
  blk000006b9 (
    .I0(sig00000118),
    .I1(sig000006f2),
    .O(sig000006d4)
  );
  LUT4 #(
    .INIT ( 16'h0001 ))
  blk000006ba (
    .I0(sig000001c2),
    .I1(sig000001c1),
    .I2(sig000001c0),
    .I3(sig000001bf),
    .O(sig000006d5)
  );
  LUT4 #(
    .INIT ( 16'h0001 ))
  blk000006bb (
    .I0(sig000001be),
    .I1(sig000001bd),
    .I2(sig000001bc),
    .I3(sig000001bb),
    .O(sig000006d6)
  );
  LUT4 #(
    .INIT ( 16'h0001 ))
  blk000006bc (
    .I0(sig000001b8),
    .I1(sig000001b7),
    .I2(sig000001ba),
    .I3(sig000001b9),
    .O(sig000006d7)
  );
  LUT4 #(
    .INIT ( 16'h0001 ))
  blk000006bd (
    .I0(sig000001b6),
    .I1(sig000001b5),
    .I2(sig000001b4),
    .I3(sig000001b3),
    .O(sig000006d8)
  );
  LUT4 #(
    .INIT ( 16'h0001 ))
  blk000006be (
    .I0(sig000001b2),
    .I1(sig000001b1),
    .I2(sig000001b0),
    .I3(sig000001af),
    .O(sig000006d9)
  );
  LUT4 #(
    .INIT ( 16'h0001 ))
  blk000006bf (
    .I0(sig000001ae),
    .I1(sig000001ad),
    .I2(sig000001ac),
    .I3(sig000001ab),
    .O(sig000006da)
  );
  LUT4 #(
    .INIT ( 16'h0001 ))
  blk000006c0 (
    .I0(sig000001aa),
    .I1(sig000001a9),
    .I2(sig000001a8),
    .I3(sig000001a7),
    .O(sig000006db)
  );
  LUT4 #(
    .INIT ( 16'h0001 ))
  blk000006c1 (
    .I0(sig000001a6),
    .I1(sig000001a5),
    .I2(sig000001a4),
    .I3(sig000001a3),
    .O(sig000006dc)
  );
  LUT4 #(
    .INIT ( 16'h0001 ))
  blk000006c2 (
    .I0(sig000001a2),
    .I1(sig000001a1),
    .I2(sig000001a0),
    .I3(sig0000019f),
    .O(sig000006dd)
  );
  LUT4 #(
    .INIT ( 16'h0001 ))
  blk000006c3 (
    .I0(sig0000019e),
    .I1(sig0000019d),
    .I2(sig0000019c),
    .I3(sig0000019b),
    .O(sig000006de)
  );
  LUT4 #(
    .INIT ( 16'h0001 ))
  blk000006c4 (
    .I0(sig0000019a),
    .I1(sig00000199),
    .I2(sig00000198),
    .I3(sig00000197),
    .O(sig000006df)
  );
  LUT4 #(
    .INIT ( 16'h0001 ))
  blk000006c5 (
    .I0(sig00000196),
    .I1(sig00000195),
    .I2(sig00000194),
    .I3(sig00000193),
    .O(sig000006e0)
  );
  LUT4 #(
    .INIT ( 16'h0001 ))
  blk000006c6 (
    .I0(sig00000192),
    .I1(sig00000191),
    .I2(sig00000190),
    .I3(sig0000018f),
    .O(sig000006e1)
  );
  LUT4 #(
    .INIT ( 16'h0001 ))
  blk000006c7 (
    .I0(sig0000018e),
    .I1(sig0000018d),
    .I2(sig0000018c),
    .I3(sig0000018b),
    .O(sig000006e2)
  );
  LUT5 #(
    .INIT ( 32'h11110010 ))
  blk000006c8 (
    .I0(sig000006f1),
    .I1(sig00000145),
    .I2(sig00000148),
    .I3(sig00000147),
    .I4(sig00000146),
    .O(sig00000713)
  );
  LUT5 #(
    .INIT ( 32'h01010100 ))
  blk000006c9 (
    .I0(sig000006f1),
    .I1(sig00000146),
    .I2(sig00000145),
    .I3(sig00000148),
    .I4(sig00000147),
    .O(sig00000712)
  );
  LUT5 #(
    .INIT ( 32'h11110010 ))
  blk000006ca (
    .I0(sig000006f1),
    .I1(sig00000149),
    .I2(sig0000014c),
    .I3(sig0000014b),
    .I4(sig0000014a),
    .O(sig00000711)
  );
  LUT5 #(
    .INIT ( 32'h01010100 ))
  blk000006cb (
    .I0(sig000006f1),
    .I1(sig0000014a),
    .I2(sig00000149),
    .I3(sig0000014c),
    .I4(sig0000014b),
    .O(sig00000710)
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  blk000006cc (
    .I0(sig00000158),
    .I1(sig0000023e),
    .O(sig000007b4)
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  blk000006cd (
    .I0(sig00000159),
    .I1(sig0000023e),
    .O(sig000007b5)
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  blk000006ce (
    .I0(sig0000015b),
    .I1(sig0000023e),
    .O(sig000007b7)
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  blk000006cf (
    .I0(sig0000015c),
    .I1(sig0000023e),
    .O(sig000007b8)
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  blk000006d0 (
    .I0(sig0000015a),
    .I1(sig0000023e),
    .O(sig000007b6)
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  blk000006d1 (
    .I0(sig0000015e),
    .I1(sig0000023e),
    .O(sig000007ba)
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  blk000006d2 (
    .I0(sig0000015f),
    .I1(sig0000023e),
    .O(sig000007bb)
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  blk000006d3 (
    .I0(sig0000015d),
    .I1(sig0000023e),
    .O(sig000007b9)
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  blk000006d4 (
    .I0(sig00000160),
    .I1(sig0000023e),
    .O(sig000007bc)
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  blk000006d5 (
    .I0(sig00000161),
    .I1(sig0000023e),
    .O(sig000007bd)
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  blk000006d6 (
    .I0(sig00000162),
    .I1(sig0000023e),
    .O(sig000007be)
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  blk000006d7 (
    .I0(sig00000163),
    .I1(sig0000023e),
    .O(sig000007bf)
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  blk000006d8 (
    .I0(sig00000165),
    .I1(sig0000023e),
    .O(sig000007c1)
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  blk000006d9 (
    .I0(sig00000166),
    .I1(sig0000023e),
    .O(sig000007c2)
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  blk000006da (
    .I0(sig00000164),
    .I1(sig0000023e),
    .O(sig000007c0)
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  blk000006db (
    .I0(sig00000167),
    .I1(sig0000023e),
    .O(sig000007c3)
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  blk000006dc (
    .I0(sig00000168),
    .I1(sig0000023e),
    .O(sig000007c4)
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  blk000006dd (
    .I0(sig00000169),
    .I1(sig0000023e),
    .O(sig000007c5)
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  blk000006de (
    .I0(sig0000016a),
    .I1(sig0000023e),
    .O(sig000007c6)
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  blk000006df (
    .I0(sig0000016c),
    .I1(sig0000023e),
    .O(sig000007c8)
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  blk000006e0 (
    .I0(sig0000016d),
    .I1(sig0000023e),
    .O(sig000007c9)
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  blk000006e1 (
    .I0(sig0000016b),
    .I1(sig0000023e),
    .O(sig000007c7)
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  blk000006e2 (
    .I0(sig0000016e),
    .I1(sig0000023e),
    .O(sig000007ca)
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  blk000006e3 (
    .I0(sig0000016f),
    .I1(sig0000023e),
    .O(sig000007cb)
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  blk000006e4 (
    .I0(sig00000170),
    .I1(sig0000023e),
    .O(sig000007cc)
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  blk000006e5 (
    .I0(sig00000171),
    .I1(sig0000023e),
    .O(sig000007cd)
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  blk000006e6 (
    .I0(sig00000173),
    .I1(sig0000023e),
    .O(sig000007cf)
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  blk000006e7 (
    .I0(sig00000174),
    .I1(sig0000023e),
    .O(sig000007d0)
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  blk000006e8 (
    .I0(sig00000172),
    .I1(sig0000023e),
    .O(sig000007ce)
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  blk000006e9 (
    .I0(sig00000176),
    .I1(sig0000023e),
    .O(sig000007d2)
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  blk000006ea (
    .I0(sig00000177),
    .I1(sig0000023e),
    .O(sig000007d3)
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  blk000006eb (
    .I0(sig00000175),
    .I1(sig0000023e),
    .O(sig000007d1)
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  blk000006ec (
    .I0(sig00000179),
    .I1(sig0000023e),
    .O(sig000007d5)
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  blk000006ed (
    .I0(sig0000017a),
    .I1(sig0000023e),
    .O(sig000007d6)
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  blk000006ee (
    .I0(sig00000178),
    .I1(sig0000023e),
    .O(sig000007d4)
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  blk000006ef (
    .I0(sig0000017b),
    .I1(sig0000023e),
    .O(sig000007d7)
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  blk000006f0 (
    .I0(sig0000017c),
    .I1(sig0000023e),
    .O(sig000007d8)
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  blk000006f1 (
    .I0(sig0000017d),
    .I1(sig0000023e),
    .O(sig000007d9)
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  blk000006f2 (
    .I0(sig0000017e),
    .I1(sig0000023e),
    .O(sig000007da)
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  blk000006f3 (
    .I0(sig00000180),
    .I1(sig0000023e),
    .O(sig000007dc)
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  blk000006f4 (
    .I0(sig00000181),
    .I1(sig0000023e),
    .O(sig000007dd)
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  blk000006f5 (
    .I0(sig0000017f),
    .I1(sig0000023e),
    .O(sig000007db)
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  blk000006f6 (
    .I0(sig00000182),
    .I1(sig0000023e),
    .O(sig000007de)
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  blk000006f7 (
    .I0(sig00000183),
    .I1(sig0000023e),
    .O(sig000007df)
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  blk000006f8 (
    .I0(sig00000184),
    .I1(sig0000023e),
    .O(sig000007e0)
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  blk000006f9 (
    .I0(sig00000185),
    .I1(sig0000023e),
    .O(sig000007e1)
  );
  LUT4 #(
    .INIT ( 16'h5410 ))
  blk000006fa (
    .I0(sig0000023e),
    .I1(sig00000767),
    .I2(sig0000075b),
    .I3(sig00000754),
    .O(sig000007e3)
  );
  LUT4 #(
    .INIT ( 16'h5410 ))
  blk000006fb (
    .I0(sig0000023e),
    .I1(sig00000767),
    .I2(sig0000075c),
    .I3(sig00000755),
    .O(sig000007e4)
  );
  LUT4 #(
    .INIT ( 16'h5410 ))
  blk000006fc (
    .I0(sig0000023e),
    .I1(sig00000767),
    .I2(sig0000075a),
    .I3(sig00000753),
    .O(sig000007e2)
  );
  LUT4 #(
    .INIT ( 16'h5410 ))
  blk000006fd (
    .I0(sig0000023e),
    .I1(sig00000767),
    .I2(sig0000075d),
    .I3(sig00000756),
    .O(sig000007e5)
  );
  LUT4 #(
    .INIT ( 16'h5410 ))
  blk000006fe (
    .I0(sig0000023e),
    .I1(sig00000767),
    .I2(sig0000075e),
    .I3(sig00000757),
    .O(sig000007e6)
  );
  LUT5 #(
    .INIT ( 32'h55555410 ))
  blk000006ff (
    .I0(sig0000023d),
    .I1(sig00000767),
    .I2(sig0000075f),
    .I3(sig00000758),
    .I4(sig0000023c),
    .O(sig000007e7)
  );
  LUT3 #(
    .INIT ( 8'h0E ))
  blk00000700 (
    .I0(sig0000022f),
    .I1(sig0000023a),
    .I2(sig0000023b),
    .O(sig000007e8)
  );
  LUT3 #(
    .INIT ( 8'h54 ))
  blk00000701 (
    .I0(sig0000023b),
    .I1(sig0000023a),
    .I2(sig00000239),
    .O(sig000007f2)
  );
  LUT3 #(
    .INIT ( 8'h0E ))
  blk00000702 (
    .I0(sig00000230),
    .I1(sig0000023a),
    .I2(sig0000023b),
    .O(sig000007e9)
  );
  LUT3 #(
    .INIT ( 8'h0E ))
  blk00000703 (
    .I0(sig00000231),
    .I1(sig0000023a),
    .I2(sig0000023b),
    .O(sig000007ea)
  );
  LUT3 #(
    .INIT ( 8'h54 ))
  blk00000704 (
    .I0(sig0000023b),
    .I1(sig0000023a),
    .I2(sig00000232),
    .O(sig000007eb)
  );
  LUT3 #(
    .INIT ( 8'h54 ))
  blk00000705 (
    .I0(sig0000023b),
    .I1(sig0000023a),
    .I2(sig00000233),
    .O(sig000007ec)
  );
  LUT3 #(
    .INIT ( 8'h54 ))
  blk00000706 (
    .I0(sig0000023b),
    .I1(sig0000023a),
    .I2(sig00000234),
    .O(sig000007ed)
  );
  LUT3 #(
    .INIT ( 8'h54 ))
  blk00000707 (
    .I0(sig0000023b),
    .I1(sig0000023a),
    .I2(sig00000235),
    .O(sig000007ee)
  );
  LUT3 #(
    .INIT ( 8'h54 ))
  blk00000708 (
    .I0(sig0000023b),
    .I1(sig0000023a),
    .I2(sig00000236),
    .O(sig000007ef)
  );
  LUT3 #(
    .INIT ( 8'h54 ))
  blk00000709 (
    .I0(sig0000023b),
    .I1(sig0000023a),
    .I2(sig00000237),
    .O(sig000007f0)
  );
  LUT3 #(
    .INIT ( 8'h54 ))
  blk0000070a (
    .I0(sig0000023b),
    .I1(sig0000023a),
    .I2(sig00000238),
    .O(sig000007f1)
  );
  LUT6 #(
    .INIT ( 64'h0001000000000001 ))
  blk0000070b (
    .I0(sig000002d0),
    .I1(sig000002cf),
    .I2(sig000002ce),
    .I3(sig000002d1),
    .I4(sig000002cc),
    .I5(sig00000189),
    .O(sig000007f3)
  );
  LUT4 #(
    .INIT ( 16'h9009 ))
  blk0000070c (
    .I0(sig00000188),
    .I1(sig000002cb),
    .I2(sig000002c7),
    .I3(sig0000011d),
    .O(sig000007f4)
  );
  LUT5 #(
    .INIT ( 32'h00009009 ))
  blk0000070d (
    .I0(sig000002c9),
    .I1(sig00000186),
    .I2(sig000002c8),
    .I3(sig0000011c),
    .I4(sig000002cd),
    .O(sig000007f5)
  );
  LUT5 #(
    .INIT ( 32'h90000000 ))
  blk0000070e (
    .I0(sig00000187),
    .I1(sig000002ca),
    .I2(sig000007f5),
    .I3(sig000007f3),
    .I4(sig000007f4),
    .O(sig0000030e)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk0000070f (
    .I0(sig000002ef),
    .I1(sig000002ee),
    .I2(sig000002ed),
    .O(sig000007f6)
  );
  LUT5 #(
    .INIT ( 32'hAA0BAA08 ))
  blk00000710 (
    .I0(sig000002f0),
    .I1(sig000002f1),
    .I2(sig000002f2),
    .I3(sig000002f3),
    .I4(sig000007f6),
    .O(sig000002a3)
  );
  LUT6 #(
    .INIT ( 64'h8000000000000000 ))
  blk00000711 (
    .I0(a[57]),
    .I1(a[56]),
    .I2(a[55]),
    .I3(a[54]),
    .I4(a[53]),
    .I5(a[52]),
    .O(sig000007f7)
  );
  LUT6 #(
    .INIT ( 64'h8000000000000000 ))
  blk00000712 (
    .I0(a[62]),
    .I1(a[61]),
    .I2(a[60]),
    .I3(a[59]),
    .I4(a[58]),
    .I5(sig000007f7),
    .O(sig00000280)
  );
  LUT6 #(
    .INIT ( 64'hFFFFFFFFFFFFFFFE ))
  blk00000713 (
    .I0(a[57]),
    .I1(a[56]),
    .I2(a[55]),
    .I3(a[54]),
    .I4(a[53]),
    .I5(a[52]),
    .O(sig000007f8)
  );
  LUT6 #(
    .INIT ( 64'h0000000000000001 ))
  blk00000714 (
    .I0(a[62]),
    .I1(a[61]),
    .I2(a[60]),
    .I3(a[59]),
    .I4(a[58]),
    .I5(sig000007f8),
    .O(sig00000281)
  );
  LUT6 #(
    .INIT ( 64'h8000000000000000 ))
  blk00000715 (
    .I0(b[57]),
    .I1(b[56]),
    .I2(b[55]),
    .I3(b[54]),
    .I4(b[53]),
    .I5(b[52]),
    .O(sig000007f9)
  );
  LUT6 #(
    .INIT ( 64'h8000000000000000 ))
  blk00000716 (
    .I0(b[62]),
    .I1(b[61]),
    .I2(b[60]),
    .I3(b[59]),
    .I4(b[58]),
    .I5(sig000007f9),
    .O(sig00000282)
  );
  LUT6 #(
    .INIT ( 64'hFFFFFFFFFFFFFFFE ))
  blk00000717 (
    .I0(b[57]),
    .I1(b[56]),
    .I2(b[55]),
    .I3(b[54]),
    .I4(b[53]),
    .I5(b[52]),
    .O(sig000007fa)
  );
  LUT6 #(
    .INIT ( 64'h0000000000000001 ))
  blk00000718 (
    .I0(b[62]),
    .I1(b[61]),
    .I2(b[60]),
    .I3(b[59]),
    .I4(b[58]),
    .I5(sig000007fa),
    .O(sig00000283)
  );
  LUT5 #(
    .INIT ( 32'h40000000 ))
  blk00000719 (
    .I0(sig000002dd),
    .I1(sig000002d2),
    .I2(sig000002d5),
    .I3(sig000002d4),
    .I4(sig000002d3),
    .O(sig000007fb)
  );
  LUT5 #(
    .INIT ( 32'h80000000 ))
  blk0000071a (
    .I0(sig000002d9),
    .I1(sig000002d8),
    .I2(sig000002dc),
    .I3(sig000002db),
    .I4(sig000002da),
    .O(sig000007fc)
  );
  LUT4 #(
    .INIT ( 16'h8000 ))
  blk0000071b (
    .I0(sig000002d7),
    .I1(sig000002d6),
    .I2(sig000007fc),
    .I3(sig000007fb),
    .O(sig0000028f)
  );
  LUT6 #(
    .INIT ( 64'h8888888880000000 ))
  blk0000071c (
    .I0(sig000003d5),
    .I1(sig000003d4),
    .I2(sig000004ce),
    .I3(sig000004cf),
    .I4(sig000004d0),
    .I5(sig000004d1),
    .O(sig000007fd)
  );
  LUT6 #(
    .INIT ( 64'hFFFFFFFFFFFFFFFE ))
  blk0000071d (
    .I0(sig000004d4),
    .I1(sig000004d5),
    .I2(sig000004d6),
    .I3(sig000004d2),
    .I4(sig000004d3),
    .I5(sig000007fd),
    .O(sig000004b9)
  );
  LUT5 #(
    .INIT ( 32'h0FFF7777 ))
  blk0000071e (
    .I0(sig0000059b),
    .I1(sig000005aa),
    .I2(sig000005ab),
    .I3(sig0000059d),
    .I4(sig0000040e),
    .O(sig000007fe)
  );
  LUT5 #(
    .INIT ( 32'h8880BBB3 ))
  blk0000071f (
    .I0(sig0000059c),
    .I1(sig0000040d),
    .I2(sig0000040e),
    .I3(sig000005c5),
    .I4(sig000007fe),
    .O(sig00000597)
  );
  LUT5 #(
    .INIT ( 32'h8888F000 ))
  blk00000720 (
    .I0(sig000005b4),
    .I1(sig000005a7),
    .I2(sig000005b6),
    .I3(sig000005a9),
    .I4(sig0000040d),
    .O(sig000007ff)
  );
  LUT6 #(
    .INIT ( 64'hFBBBEAAA51114000 ))
  blk00000721 (
    .I0(sig0000040e),
    .I1(sig0000040d),
    .I2(sig000005a8),
    .I3(sig000005b5),
    .I4(sig000005a6),
    .I5(sig000007ff),
    .O(sig0000059a)
  );
  LUT5 #(
    .INIT ( 32'h8888F000 ))
  blk00000722 (
    .I0(sig000005ad),
    .I1(sig0000059f),
    .I2(sig000005af),
    .I3(sig000005a1),
    .I4(sig0000040d),
    .O(sig00000800)
  );
  LUT5 #(
    .INIT ( 32'h8888F000 ))
  blk00000723 (
    .I0(sig000005ae),
    .I1(sig000005a0),
    .I2(sig000005ac),
    .I3(sig0000059e),
    .I4(sig0000040d),
    .O(sig00000801)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk00000724 (
    .I0(sig0000040e),
    .I1(sig00000800),
    .I2(sig00000801),
    .O(sig00000598)
  );
  LUT5 #(
    .INIT ( 32'h8888F000 ))
  blk00000725 (
    .I0(sig000005b1),
    .I1(sig000005a3),
    .I2(sig000005b3),
    .I3(sig000005a5),
    .I4(sig0000040d),
    .O(sig00000802)
  );
  LUT5 #(
    .INIT ( 32'h8888F000 ))
  blk00000726 (
    .I0(sig000005b2),
    .I1(sig000005a4),
    .I2(sig000005b0),
    .I3(sig000005a2),
    .I4(sig0000040d),
    .O(sig00000803)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk00000727 (
    .I0(sig0000040e),
    .I1(sig00000802),
    .I2(sig00000803),
    .O(sig00000599)
  );
  LUT4 #(
    .INIT ( 16'hFF45 ))
  blk00000728 (
    .I0(sig0000013e),
    .I1(sig0000013f),
    .I2(sig00000140),
    .I3(sig0000013d),
    .O(sig00000804)
  );
  LUT6 #(
    .INIT ( 64'h2222020077775755 ))
  blk00000729 (
    .I0(sig000006f1),
    .I1(sig0000014d),
    .I2(sig0000014f),
    .I3(sig00000150),
    .I4(sig0000014e),
    .I5(sig00000804),
    .O(sig00000717)
  );
  LUT4 #(
    .INIT ( 16'hFFAB ))
  blk0000072a (
    .I0(sig0000013e),
    .I1(sig0000013f),
    .I2(sig00000140),
    .I3(sig0000013d),
    .O(sig00000805)
  );
  LUT6 #(
    .INIT ( 64'h0404040037373733 ))
  blk0000072b (
    .I0(sig0000014d),
    .I1(sig000006f1),
    .I2(sig0000014e),
    .I3(sig00000150),
    .I4(sig0000014f),
    .I5(sig00000805),
    .O(sig00000716)
  );
  LUT4 #(
    .INIT ( 16'hFF45 ))
  blk0000072c (
    .I0(sig00000142),
    .I1(sig00000143),
    .I2(sig00000144),
    .I3(sig00000141),
    .O(sig00000806)
  );
  LUT6 #(
    .INIT ( 64'h2222020077775755 ))
  blk0000072d (
    .I0(sig000006f1),
    .I1(sig00000151),
    .I2(sig00000153),
    .I3(sig00000154),
    .I4(sig00000152),
    .I5(sig00000806),
    .O(sig00000715)
  );
  LUT4 #(
    .INIT ( 16'hFFAB ))
  blk0000072e (
    .I0(sig00000142),
    .I1(sig00000143),
    .I2(sig00000144),
    .I3(sig00000141),
    .O(sig00000807)
  );
  LUT6 #(
    .INIT ( 64'h0404040037373733 ))
  blk0000072f (
    .I0(sig00000151),
    .I1(sig000006f1),
    .I2(sig00000152),
    .I3(sig00000154),
    .I4(sig00000153),
    .I5(sig00000807),
    .O(sig00000714)
  );
  LUT4 #(
    .INIT ( 16'hFF45 ))
  blk00000730 (
    .I0(sig0000012e),
    .I1(sig0000012f),
    .I2(sig00000130),
    .I3(sig0000012d),
    .O(sig00000808)
  );
  LUT6 #(
    .INIT ( 64'h10111010BABBBABA ))
  blk00000731 (
    .I0(sig000006f9),
    .I1(sig0000027f),
    .I2(sig0000011e),
    .I3(sig0000011f),
    .I4(sig00000120),
    .I5(sig00000808),
    .O(sig0000071f)
  );
  LUT4 #(
    .INIT ( 16'hFFAB ))
  blk00000732 (
    .I0(sig0000012d),
    .I1(sig0000012f),
    .I2(sig00000130),
    .I3(sig0000012e),
    .O(sig00000809)
  );
  LUT6 #(
    .INIT ( 64'h01010100CDCDCDCC ))
  blk00000733 (
    .I0(sig0000027f),
    .I1(sig000006f9),
    .I2(sig0000011e),
    .I3(sig00000120),
    .I4(sig0000011f),
    .I5(sig00000809),
    .O(sig0000071e)
  );
  LUT4 #(
    .INIT ( 16'hFF45 ))
  blk00000734 (
    .I0(sig00000132),
    .I1(sig00000133),
    .I2(sig00000134),
    .I3(sig00000131),
    .O(sig0000080a)
  );
  LUT6 #(
    .INIT ( 64'h10111010BABBBABA ))
  blk00000735 (
    .I0(sig000006f9),
    .I1(sig00000121),
    .I2(sig00000122),
    .I3(sig00000123),
    .I4(sig00000124),
    .I5(sig0000080a),
    .O(sig0000071d)
  );
  LUT4 #(
    .INIT ( 16'hFFAB ))
  blk00000736 (
    .I0(sig00000131),
    .I1(sig00000133),
    .I2(sig00000134),
    .I3(sig00000132),
    .O(sig0000080b)
  );
  LUT6 #(
    .INIT ( 64'h01010100CDCDCDCC ))
  blk00000737 (
    .I0(sig00000122),
    .I1(sig000006f9),
    .I2(sig00000121),
    .I3(sig00000124),
    .I4(sig00000123),
    .I5(sig0000080b),
    .O(sig0000071c)
  );
  LUT4 #(
    .INIT ( 16'hFF45 ))
  blk00000738 (
    .I0(sig00000136),
    .I1(sig00000137),
    .I2(sig00000138),
    .I3(sig00000135),
    .O(sig0000080c)
  );
  LUT6 #(
    .INIT ( 64'h10111010BABBBABA ))
  blk00000739 (
    .I0(sig000006f9),
    .I1(sig00000125),
    .I2(sig00000126),
    .I3(sig00000127),
    .I4(sig00000128),
    .I5(sig0000080c),
    .O(sig0000071b)
  );
  LUT4 #(
    .INIT ( 16'hFFAB ))
  blk0000073a (
    .I0(sig00000135),
    .I1(sig00000137),
    .I2(sig00000138),
    .I3(sig00000136),
    .O(sig0000080d)
  );
  LUT6 #(
    .INIT ( 64'h01010100CDCDCDCC ))
  blk0000073b (
    .I0(sig00000126),
    .I1(sig000006f9),
    .I2(sig00000125),
    .I3(sig00000128),
    .I4(sig00000127),
    .I5(sig0000080d),
    .O(sig0000071a)
  );
  LUT4 #(
    .INIT ( 16'hFF45 ))
  blk0000073c (
    .I0(sig0000013a),
    .I1(sig0000013b),
    .I2(sig0000013c),
    .I3(sig00000139),
    .O(sig0000080e)
  );
  LUT6 #(
    .INIT ( 64'h10111010BABBBABA ))
  blk0000073d (
    .I0(sig000006f9),
    .I1(sig00000129),
    .I2(sig0000012a),
    .I3(sig0000012b),
    .I4(sig0000012c),
    .I5(sig0000080e),
    .O(sig00000719)
  );
  LUT4 #(
    .INIT ( 16'hFFAB ))
  blk0000073e (
    .I0(sig00000139),
    .I1(sig0000013b),
    .I2(sig0000013c),
    .I3(sig0000013a),
    .O(sig0000080f)
  );
  LUT6 #(
    .INIT ( 64'h01010100CDCDCDCC ))
  blk0000073f (
    .I0(sig0000012a),
    .I1(sig000006f9),
    .I2(sig00000129),
    .I3(sig0000012c),
    .I4(sig0000012b),
    .I5(sig0000080f),
    .O(sig00000718)
  );
  LUT2 #(
    .INIT ( 4'hD ))
  blk00000740 (
    .I0(sig0000003b),
    .I1(sig0000011d),
    .O(sig00000810)
  );
  LUT6 #(
    .INIT ( 64'hFFFF00005D5F0000 ))
  blk00000741 (
    .I0(sig00000155),
    .I1(sig0000003a),
    .I2(sig0000011c),
    .I3(sig00000810),
    .I4(sig000000e2),
    .I5(sig000000e3),
    .O(sig00000720)
  );
  FD   blk00000742 (
    .C(clk),
    .D(sig0000022b),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.LOGIC.OP/OP/sign_op )
  );
  LUT5 #(
    .INIT ( 32'hAAAA59A6 ))
  blk00000743 (
    .I0(sig00000608),
    .I1(sig00000600),
    .I2(sig000005f8),
    .I3(sig00000696),
    .I4(sig00000697),
    .O(sig00000811)
  );
  LUT5 #(
    .INIT ( 32'hAAAA59A6 ))
  blk00000744 (
    .I0(sig00000607),
    .I1(sig000005ff),
    .I2(sig000005f8),
    .I3(sig00000696),
    .I4(sig00000697),
    .O(sig00000812)
  );
  LUT6 #(
    .INIT ( 64'hAAAAAAAAA5995A66 ))
  blk00000745 (
    .I0(sig00000606),
    .I1(sig000005fe),
    .I2(sig00000600),
    .I3(sig000005f8),
    .I4(sig00000696),
    .I5(sig00000697),
    .O(sig00000813)
  );
  LUT6 #(
    .INIT ( 64'hAAAAAAAAA5995A66 ))
  blk00000746 (
    .I0(sig00000605),
    .I1(sig000005fd),
    .I2(sig000005ff),
    .I3(sig000005f8),
    .I4(sig00000696),
    .I5(sig00000697),
    .O(sig00000814)
  );
  LUT6 #(
    .INIT ( 64'hAAAAAAAAA5995A66 ))
  blk00000747 (
    .I0(sig00000604),
    .I1(sig000005fc),
    .I2(sig000005fe),
    .I3(sig000005f8),
    .I4(sig00000696),
    .I5(sig00000697),
    .O(sig00000815)
  );
  LUT6 #(
    .INIT ( 64'hAAAAAAAAA5995A66 ))
  blk00000748 (
    .I0(sig00000603),
    .I1(sig000005fb),
    .I2(sig000005fd),
    .I3(sig000005f8),
    .I4(sig00000696),
    .I5(sig00000697),
    .O(sig00000816)
  );
  LUT6 #(
    .INIT ( 64'hCCCCCCCCC3993C66 ))
  blk00000749 (
    .I0(sig000005fa),
    .I1(sig00000602),
    .I2(sig000005fc),
    .I3(sig000005f8),
    .I4(sig00000696),
    .I5(sig00000697),
    .O(sig00000817)
  );
  LUT6 #(
    .INIT ( 64'hCCCCCCCCC3993C66 ))
  blk0000074a (
    .I0(sig000005f9),
    .I1(sig00000601),
    .I2(sig000005fb),
    .I3(sig000005f8),
    .I4(sig00000696),
    .I5(sig00000697),
    .O(sig00000818)
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  blk0000074b (
    .I0(sig00000761),
    .O(sig00000819)
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  blk0000074c (
    .I0(sig00000762),
    .O(sig0000081a)
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  blk0000074d (
    .I0(sig00000763),
    .O(sig0000081b)
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  blk0000074e (
    .I0(sig00000764),
    .O(sig0000081c)
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  blk0000074f (
    .I0(sig00000765),
    .O(sig0000081d)
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  blk00000750 (
    .I0(sig00000766),
    .O(sig0000081e)
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  blk00000751 (
    .I0(sig00000760),
    .O(sig0000081f)
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  blk00000752 (
    .I0(sig00000761),
    .O(sig00000820)
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  blk00000753 (
    .I0(sig00000762),
    .O(sig00000821)
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  blk00000754 (
    .I0(sig00000763),
    .O(sig00000822)
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  blk00000755 (
    .I0(sig00000764),
    .O(sig00000823)
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  blk00000756 (
    .I0(sig00000765),
    .O(sig00000824)
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  blk00000757 (
    .I0(sig00000766),
    .O(sig00000825)
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  blk00000758 (
    .I0(sig00000760),
    .O(sig00000826)
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  blk00000759 (
    .I0(sig00000696),
    .I1(sig00000697),
    .O(sig00000827)
  );
  LUT6 #(
    .INIT ( 64'h0000FFA50000FFC3 ))
  blk0000075a (
    .I0(sig00000759),
    .I1(sig0000059c),
    .I2(sig0000022f),
    .I3(sig0000023a),
    .I4(sig0000023b),
    .I5(sig00000767),
    .O(sig000007a8)
  );
  LUT4 #(
    .INIT ( 16'h5410 ))
  blk0000075b (
    .I0(sig00000118),
    .I1(sig000006f9),
    .I2(sig00000144),
    .I3(sig00000154),
    .O(sig00000082)
  );
  LUT4 #(
    .INIT ( 16'h5410 ))
  blk0000075c (
    .I0(sig00000118),
    .I1(sig000006f9),
    .I2(sig00000143),
    .I3(sig00000153),
    .O(sig00000083)
  );
  LUT4 #(
    .INIT ( 16'h5410 ))
  blk0000075d (
    .I0(sig00000118),
    .I1(sig000006f9),
    .I2(sig0000013d),
    .I3(sig0000014d),
    .O(sig00000089)
  );
  LUT4 #(
    .INIT ( 16'h5410 ))
  blk0000075e (
    .I0(sig00000118),
    .I1(sig000006f9),
    .I2(sig00000142),
    .I3(sig00000152),
    .O(sig00000084)
  );
  LUT4 #(
    .INIT ( 16'h5410 ))
  blk0000075f (
    .I0(sig00000118),
    .I1(sig000006f9),
    .I2(sig00000141),
    .I3(sig00000151),
    .O(sig00000085)
  );
  LUT4 #(
    .INIT ( 16'h5410 ))
  blk00000760 (
    .I0(sig00000118),
    .I1(sig000006f9),
    .I2(sig00000140),
    .I3(sig00000150),
    .O(sig00000086)
  );
  LUT4 #(
    .INIT ( 16'h5410 ))
  blk00000761 (
    .I0(sig00000118),
    .I1(sig000006f9),
    .I2(sig0000013f),
    .I3(sig0000014f),
    .O(sig00000087)
  );
  LUT4 #(
    .INIT ( 16'h5410 ))
  blk00000762 (
    .I0(sig00000118),
    .I1(sig000006f9),
    .I2(sig0000013e),
    .I3(sig0000014e),
    .O(sig00000088)
  );
  LUT4 #(
    .INIT ( 16'h5410 ))
  blk00000763 (
    .I0(sig0000011a),
    .I1(sig000006e4),
    .I2(sig00000006),
    .I3(sig00000002),
    .O(sig000000ae)
  );
  LUT4 #(
    .INIT ( 16'h5410 ))
  blk00000764 (
    .I0(sig0000011a),
    .I1(sig000006e4),
    .I2(sig00000007),
    .I3(sig00000003),
    .O(sig000000af)
  );
  LUT4 #(
    .INIT ( 16'h5410 ))
  blk00000765 (
    .I0(sig0000011a),
    .I1(sig000006e4),
    .I2(sig00000008),
    .I3(sig00000004),
    .O(sig000000b0)
  );
  LUT4 #(
    .INIT ( 16'h5410 ))
  blk00000766 (
    .I0(sig0000011a),
    .I1(sig000006e4),
    .I2(sig00000009),
    .I3(sig00000005),
    .O(sig000000b1)
  );
  LUT4 #(
    .INIT ( 16'h5410 ))
  blk00000767 (
    .I0(sig00000118),
    .I1(sig000006f9),
    .I2(sig00000135),
    .I3(sig00000145),
    .O(sig00000091)
  );
  LUT4 #(
    .INIT ( 16'h5410 ))
  blk00000768 (
    .I0(sig00000118),
    .I1(sig000006f9),
    .I2(sig00000136),
    .I3(sig00000146),
    .O(sig00000090)
  );
  LUT4 #(
    .INIT ( 16'h5410 ))
  blk00000769 (
    .I0(sig00000118),
    .I1(sig000006f9),
    .I2(sig00000137),
    .I3(sig00000147),
    .O(sig0000008f)
  );
  LUT4 #(
    .INIT ( 16'h5410 ))
  blk0000076a (
    .I0(sig00000118),
    .I1(sig000006f9),
    .I2(sig00000138),
    .I3(sig00000148),
    .O(sig0000008e)
  );
  LUT4 #(
    .INIT ( 16'h5410 ))
  blk0000076b (
    .I0(sig00000118),
    .I1(sig000006f9),
    .I2(sig00000139),
    .I3(sig00000149),
    .O(sig0000008d)
  );
  LUT4 #(
    .INIT ( 16'h5410 ))
  blk0000076c (
    .I0(sig00000118),
    .I1(sig000006f9),
    .I2(sig0000013a),
    .I3(sig0000014a),
    .O(sig0000008c)
  );
  LUT4 #(
    .INIT ( 16'h5410 ))
  blk0000076d (
    .I0(sig00000118),
    .I1(sig000006f9),
    .I2(sig0000013b),
    .I3(sig0000014b),
    .O(sig0000008b)
  );
  LUT4 #(
    .INIT ( 16'h5410 ))
  blk0000076e (
    .I0(sig00000118),
    .I1(sig000006f9),
    .I2(sig0000013c),
    .I3(sig0000014c),
    .O(sig0000008a)
  );
  LUT3 #(
    .INIT ( 8'h10 ))
  blk0000076f (
    .I0(sig0000011a),
    .I1(sig000006e4),
    .I2(sig00000005),
    .O(sig000000ad)
  );
  LUT3 #(
    .INIT ( 8'h10 ))
  blk00000770 (
    .I0(sig0000011a),
    .I1(sig000006e4),
    .I2(sig00000004),
    .O(sig000000ac)
  );
  LUT3 #(
    .INIT ( 8'h10 ))
  blk00000771 (
    .I0(sig0000011a),
    .I1(sig000006e4),
    .I2(sig00000003),
    .O(sig000000ab)
  );
  LUT3 #(
    .INIT ( 8'h10 ))
  blk00000772 (
    .I0(sig0000011a),
    .I1(sig000006e4),
    .I2(sig00000002),
    .O(sig000000aa)
  );
  LUT3 #(
    .INIT ( 8'h10 ))
  blk00000773 (
    .I0(sig00000118),
    .I1(sig000006f9),
    .I2(sig00000145),
    .O(sig00000081)
  );
  LUT3 #(
    .INIT ( 8'h10 ))
  blk00000774 (
    .I0(sig00000118),
    .I1(sig000006f9),
    .I2(sig00000146),
    .O(sig00000080)
  );
  LUT3 #(
    .INIT ( 8'h10 ))
  blk00000775 (
    .I0(sig00000118),
    .I1(sig000006f9),
    .I2(sig00000147),
    .O(sig0000007f)
  );
  LUT3 #(
    .INIT ( 8'h10 ))
  blk00000776 (
    .I0(sig00000118),
    .I1(sig000006f9),
    .I2(sig00000148),
    .O(sig0000007e)
  );
  LUT3 #(
    .INIT ( 8'h10 ))
  blk00000777 (
    .I0(sig00000118),
    .I1(sig000006f9),
    .I2(sig00000149),
    .O(sig0000007d)
  );
  LUT3 #(
    .INIT ( 8'h10 ))
  blk00000778 (
    .I0(sig00000118),
    .I1(sig000006f9),
    .I2(sig0000014a),
    .O(sig0000007c)
  );
  LUT3 #(
    .INIT ( 8'h10 ))
  blk00000779 (
    .I0(sig00000118),
    .I1(sig000006f9),
    .I2(sig0000014b),
    .O(sig0000007b)
  );
  LUT3 #(
    .INIT ( 8'h10 ))
  blk0000077a (
    .I0(sig00000118),
    .I1(sig000006f9),
    .I2(sig0000014c),
    .O(sig0000007a)
  );
  LUT3 #(
    .INIT ( 8'h10 ))
  blk0000077b (
    .I0(sig00000118),
    .I1(sig000006f9),
    .I2(sig0000014d),
    .O(sig00000079)
  );
  LUT3 #(
    .INIT ( 8'h10 ))
  blk0000077c (
    .I0(sig00000118),
    .I1(sig000006f9),
    .I2(sig0000014e),
    .O(sig00000078)
  );
  LUT3 #(
    .INIT ( 8'h10 ))
  blk0000077d (
    .I0(sig00000118),
    .I1(sig000006f9),
    .I2(sig0000014f),
    .O(sig00000077)
  );
  LUT3 #(
    .INIT ( 8'h10 ))
  blk0000077e (
    .I0(sig00000118),
    .I1(sig000006f9),
    .I2(sig00000150),
    .O(sig00000076)
  );
  LUT3 #(
    .INIT ( 8'h10 ))
  blk0000077f (
    .I0(sig00000118),
    .I1(sig000006f9),
    .I2(sig00000151),
    .O(sig00000075)
  );
  LUT3 #(
    .INIT ( 8'h10 ))
  blk00000780 (
    .I0(sig00000118),
    .I1(sig000006f9),
    .I2(sig00000152),
    .O(sig00000074)
  );
  LUT3 #(
    .INIT ( 8'h10 ))
  blk00000781 (
    .I0(sig00000118),
    .I1(sig000006f9),
    .I2(sig00000153),
    .O(sig00000073)
  );
  LUT3 #(
    .INIT ( 8'h10 ))
  blk00000782 (
    .I0(sig00000118),
    .I1(sig000006f9),
    .I2(sig00000154),
    .O(sig00000072)
  );
  LUT6 #(
    .INIT ( 64'h5410FEBA54105410 ))
  blk00000783 (
    .I0(sig0000011a),
    .I1(sig000006e4),
    .I2(sig0000000a),
    .I3(sig00000006),
    .I4(sig000006e3),
    .I5(sig00000002),
    .O(sig000000b2)
  );
  LUT6 #(
    .INIT ( 64'h5410FEBA54105410 ))
  blk00000784 (
    .I0(sig0000011a),
    .I1(sig000006e4),
    .I2(sig0000000b),
    .I3(sig00000007),
    .I4(sig000006e3),
    .I5(sig00000003),
    .O(sig000000b3)
  );
  LUT6 #(
    .INIT ( 64'h5410FEBA54105410 ))
  blk00000785 (
    .I0(sig0000011a),
    .I1(sig000006e4),
    .I2(sig0000000c),
    .I3(sig00000008),
    .I4(sig000006e3),
    .I5(sig00000004),
    .O(sig000000b4)
  );
  LUT6 #(
    .INIT ( 64'h5410FEBA54105410 ))
  blk00000786 (
    .I0(sig0000011a),
    .I1(sig000006e4),
    .I2(sig0000000d),
    .I3(sig00000009),
    .I4(sig000006e3),
    .I5(sig00000005),
    .O(sig000000b5)
  );
  LUT6 #(
    .INIT ( 64'h5410FEBA54105410 ))
  blk00000787 (
    .I0(sig00000118),
    .I1(sig000006f9),
    .I2(sig00000127),
    .I3(sig00000137),
    .I4(sig000006f1),
    .I5(sig00000147),
    .O(sig0000009f)
  );
  LUT6 #(
    .INIT ( 64'h5410FEBA54105410 ))
  blk00000788 (
    .I0(sig00000118),
    .I1(sig000006f9),
    .I2(sig00000128),
    .I3(sig00000138),
    .I4(sig000006f1),
    .I5(sig00000148),
    .O(sig0000009e)
  );
  LUT6 #(
    .INIT ( 64'h5410FEBA54105410 ))
  blk00000789 (
    .I0(sig00000118),
    .I1(sig000006f9),
    .I2(sig00000129),
    .I3(sig00000139),
    .I4(sig000006f1),
    .I5(sig00000149),
    .O(sig0000009d)
  );
  LUT6 #(
    .INIT ( 64'h5410FEBA54105410 ))
  blk0000078a (
    .I0(sig00000118),
    .I1(sig000006f9),
    .I2(sig0000012a),
    .I3(sig0000013a),
    .I4(sig000006f1),
    .I5(sig0000014a),
    .O(sig0000009c)
  );
  LUT6 #(
    .INIT ( 64'h5410FEBA54105410 ))
  blk0000078b (
    .I0(sig00000118),
    .I1(sig000006f9),
    .I2(sig0000012b),
    .I3(sig0000013b),
    .I4(sig000006f1),
    .I5(sig0000014b),
    .O(sig0000009b)
  );
  LUT6 #(
    .INIT ( 64'h5410FEBA54105410 ))
  blk0000078c (
    .I0(sig00000118),
    .I1(sig000006f9),
    .I2(sig0000012c),
    .I3(sig0000013c),
    .I4(sig000006f1),
    .I5(sig0000014c),
    .O(sig0000009a)
  );
  LUT6 #(
    .INIT ( 64'h5410FEBA54105410 ))
  blk0000078d (
    .I0(sig00000118),
    .I1(sig000006f9),
    .I2(sig0000012d),
    .I3(sig0000013d),
    .I4(sig000006f1),
    .I5(sig0000014d),
    .O(sig00000099)
  );
  LUT6 #(
    .INIT ( 64'h5410FEBA54105410 ))
  blk0000078e (
    .I0(sig00000118),
    .I1(sig000006f9),
    .I2(sig0000012e),
    .I3(sig0000013e),
    .I4(sig000006f1),
    .I5(sig0000014e),
    .O(sig00000098)
  );
  LUT6 #(
    .INIT ( 64'h5410FEBA54105410 ))
  blk0000078f (
    .I0(sig00000118),
    .I1(sig000006f9),
    .I2(sig0000012f),
    .I3(sig0000013f),
    .I4(sig000006f1),
    .I5(sig0000014f),
    .O(sig00000097)
  );
  LUT6 #(
    .INIT ( 64'h5410FEBA54105410 ))
  blk00000790 (
    .I0(sig00000118),
    .I1(sig000006f9),
    .I2(sig00000130),
    .I3(sig00000140),
    .I4(sig000006f1),
    .I5(sig00000150),
    .O(sig00000096)
  );
  LUT6 #(
    .INIT ( 64'h5410FEBA54105410 ))
  blk00000791 (
    .I0(sig00000118),
    .I1(sig000006f9),
    .I2(sig00000131),
    .I3(sig00000141),
    .I4(sig000006f1),
    .I5(sig00000151),
    .O(sig00000095)
  );
  LUT6 #(
    .INIT ( 64'h5410FEBA54105410 ))
  blk00000792 (
    .I0(sig00000118),
    .I1(sig000006f9),
    .I2(sig00000132),
    .I3(sig00000142),
    .I4(sig000006f1),
    .I5(sig00000152),
    .O(sig00000094)
  );
  LUT6 #(
    .INIT ( 64'h5410FEBA54105410 ))
  blk00000793 (
    .I0(sig00000118),
    .I1(sig000006f9),
    .I2(sig00000133),
    .I3(sig00000143),
    .I4(sig000006f1),
    .I5(sig00000153),
    .O(sig00000093)
  );
  LUT6 #(
    .INIT ( 64'h5410FEBA54105410 ))
  blk00000794 (
    .I0(sig00000118),
    .I1(sig000006f9),
    .I2(sig00000134),
    .I3(sig00000144),
    .I4(sig000006f1),
    .I5(sig00000154),
    .O(sig00000092)
  );
  LUT6 #(
    .INIT ( 64'h5410FEBA54105410 ))
  blk00000795 (
    .I0(sig00000118),
    .I1(sig000006f9),
    .I2(sig00000125),
    .I3(sig00000135),
    .I4(sig000006f1),
    .I5(sig00000145),
    .O(sig000000a1)
  );
  LUT6 #(
    .INIT ( 64'h5410FEBA54105410 ))
  blk00000796 (
    .I0(sig00000118),
    .I1(sig000006f9),
    .I2(sig00000126),
    .I3(sig00000136),
    .I4(sig000006f1),
    .I5(sig00000146),
    .O(sig000000a0)
  );
  LUT6 #(
    .INIT ( 64'hFFFFFFFFFEEE0444 ))
  blk00000797 (
    .I0(sig0000027b),
    .I1(sig000001f6),
    .I2(sig0000027a),
    .I3(sig0000027c),
    .I4(sig0000022a),
    .I5(sig0000023f),
    .O(sig00000542)
  );
  LUT6 #(
    .INIT ( 64'hAAA8A8A800202020 ))
  blk00000798 (
    .I0(sig0000023f),
    .I1(sig0000027b),
    .I2(sig000001c3),
    .I3(sig0000027a),
    .I4(sig0000027c),
    .I5(sig000001f7),
    .O(sig0000050e)
  );
  LUT2 #(
    .INIT ( 4'h7 ))
  blk00000799 (
    .I0(sig0000030f),
    .I1(sig00000312),
    .O(sig00000579)
  );
  LUT3 #(
    .INIT ( 8'h01 ))
  blk0000079a (
    .I0(sig000004cb),
    .I1(sig000004cd),
    .I2(sig00000544),
    .O(sig000004b7)
  );
  LUT3 #(
    .INIT ( 8'h10 ))
  blk0000079b (
    .I0(sig000004cd),
    .I1(sig00000544),
    .I2(sig000004cb),
    .O(sig000004b8)
  );
  LUT3 #(
    .INIT ( 8'h10 ))
  blk0000079c (
    .I0(sig000004cd),
    .I1(sig00000544),
    .I2(sig000004b4),
    .O(sig000004ba)
  );
  LUT5 #(
    .INIT ( 32'h0AAA0CCC ))
  blk0000079d (
    .I0(sig000001c3),
    .I1(sig000001f7),
    .I2(sig00000312),
    .I3(sig0000030f),
    .I4(sig0000022e),
    .O(sig00000545)
  );
  LUT5 #(
    .INIT ( 32'h0AAA0CCC ))
  blk0000079e (
    .I0(sig000001cd),
    .I1(sig00000201),
    .I2(sig00000312),
    .I3(sig0000030f),
    .I4(sig0000022e),
    .O(sig0000054f)
  );
  LUT5 #(
    .INIT ( 32'h0AAA0CCC ))
  blk0000079f (
    .I0(sig000001ce),
    .I1(sig00000202),
    .I2(sig00000312),
    .I3(sig0000030f),
    .I4(sig0000022e),
    .O(sig00000550)
  );
  LUT5 #(
    .INIT ( 32'h0AAA0CCC ))
  blk000007a0 (
    .I0(sig000001cf),
    .I1(sig00000203),
    .I2(sig00000312),
    .I3(sig0000030f),
    .I4(sig0000022e),
    .O(sig00000551)
  );
  LUT5 #(
    .INIT ( 32'h0AAA0CCC ))
  blk000007a1 (
    .I0(sig000001d0),
    .I1(sig00000204),
    .I2(sig00000312),
    .I3(sig0000030f),
    .I4(sig0000022e),
    .O(sig00000552)
  );
  LUT5 #(
    .INIT ( 32'h0AAA0CCC ))
  blk000007a2 (
    .I0(sig000001d1),
    .I1(sig00000205),
    .I2(sig00000312),
    .I3(sig0000030f),
    .I4(sig0000022e),
    .O(sig00000553)
  );
  LUT5 #(
    .INIT ( 32'h0AAA0CCC ))
  blk000007a3 (
    .I0(sig000001d2),
    .I1(sig00000206),
    .I2(sig00000312),
    .I3(sig0000030f),
    .I4(sig0000022e),
    .O(sig00000554)
  );
  LUT5 #(
    .INIT ( 32'h0AAA0CCC ))
  blk000007a4 (
    .I0(sig000001d3),
    .I1(sig00000207),
    .I2(sig00000312),
    .I3(sig0000030f),
    .I4(sig0000022e),
    .O(sig00000555)
  );
  LUT5 #(
    .INIT ( 32'h0AAA0CCC ))
  blk000007a5 (
    .I0(sig000001d4),
    .I1(sig00000208),
    .I2(sig00000312),
    .I3(sig0000030f),
    .I4(sig0000022e),
    .O(sig00000556)
  );
  LUT5 #(
    .INIT ( 32'h0AAA0CCC ))
  blk000007a6 (
    .I0(sig000001d5),
    .I1(sig00000209),
    .I2(sig00000312),
    .I3(sig0000030f),
    .I4(sig0000022e),
    .O(sig00000557)
  );
  LUT5 #(
    .INIT ( 32'h0AAA0CCC ))
  blk000007a7 (
    .I0(sig000001d6),
    .I1(sig0000020a),
    .I2(sig00000312),
    .I3(sig0000030f),
    .I4(sig0000022e),
    .O(sig00000558)
  );
  LUT5 #(
    .INIT ( 32'h0AAA0CCC ))
  blk000007a8 (
    .I0(sig000001c4),
    .I1(sig000001f8),
    .I2(sig00000312),
    .I3(sig0000030f),
    .I4(sig0000022e),
    .O(sig00000546)
  );
  LUT5 #(
    .INIT ( 32'h0AAA0CCC ))
  blk000007a9 (
    .I0(sig000001d7),
    .I1(sig0000020b),
    .I2(sig00000312),
    .I3(sig0000030f),
    .I4(sig0000022e),
    .O(sig00000559)
  );
  LUT5 #(
    .INIT ( 32'h0AAA0CCC ))
  blk000007aa (
    .I0(sig000001d8),
    .I1(sig0000020c),
    .I2(sig00000312),
    .I3(sig0000030f),
    .I4(sig0000022e),
    .O(sig0000055a)
  );
  LUT5 #(
    .INIT ( 32'h0AAA0CCC ))
  blk000007ab (
    .I0(sig000001d9),
    .I1(sig0000020d),
    .I2(sig00000312),
    .I3(sig0000030f),
    .I4(sig0000022e),
    .O(sig0000055b)
  );
  LUT5 #(
    .INIT ( 32'h0AAA0CCC ))
  blk000007ac (
    .I0(sig000001da),
    .I1(sig0000020e),
    .I2(sig00000312),
    .I3(sig0000030f),
    .I4(sig0000022e),
    .O(sig0000055c)
  );
  LUT5 #(
    .INIT ( 32'h0AAA0CCC ))
  blk000007ad (
    .I0(sig000001db),
    .I1(sig0000020f),
    .I2(sig00000312),
    .I3(sig0000030f),
    .I4(sig0000022e),
    .O(sig0000055d)
  );
  LUT5 #(
    .INIT ( 32'h0AAA0CCC ))
  blk000007ae (
    .I0(sig000001dc),
    .I1(sig00000210),
    .I2(sig00000312),
    .I3(sig0000030f),
    .I4(sig0000022e),
    .O(sig0000055e)
  );
  LUT5 #(
    .INIT ( 32'h0AAA0CCC ))
  blk000007af (
    .I0(sig000001dd),
    .I1(sig00000211),
    .I2(sig00000312),
    .I3(sig0000030f),
    .I4(sig0000022e),
    .O(sig0000055f)
  );
  LUT5 #(
    .INIT ( 32'h0AAA0CCC ))
  blk000007b0 (
    .I0(sig000001de),
    .I1(sig00000212),
    .I2(sig00000312),
    .I3(sig0000030f),
    .I4(sig0000022e),
    .O(sig00000560)
  );
  LUT5 #(
    .INIT ( 32'h0AAA0CCC ))
  blk000007b1 (
    .I0(sig000001df),
    .I1(sig00000213),
    .I2(sig00000312),
    .I3(sig0000030f),
    .I4(sig0000022e),
    .O(sig00000561)
  );
  LUT5 #(
    .INIT ( 32'h0AAA0CCC ))
  blk000007b2 (
    .I0(sig000001e0),
    .I1(sig00000214),
    .I2(sig00000312),
    .I3(sig0000030f),
    .I4(sig0000022e),
    .O(sig00000562)
  );
  LUT5 #(
    .INIT ( 32'h0AAA0CCC ))
  blk000007b3 (
    .I0(sig000001c5),
    .I1(sig000001f9),
    .I2(sig00000312),
    .I3(sig0000030f),
    .I4(sig0000022e),
    .O(sig00000547)
  );
  LUT5 #(
    .INIT ( 32'h0AAA0CCC ))
  blk000007b4 (
    .I0(sig000001e1),
    .I1(sig00000215),
    .I2(sig00000312),
    .I3(sig0000030f),
    .I4(sig0000022e),
    .O(sig00000563)
  );
  LUT5 #(
    .INIT ( 32'h0AAA0CCC ))
  blk000007b5 (
    .I0(sig000001e2),
    .I1(sig00000216),
    .I2(sig00000312),
    .I3(sig0000030f),
    .I4(sig0000022e),
    .O(sig00000564)
  );
  LUT5 #(
    .INIT ( 32'h0AAA0CCC ))
  blk000007b6 (
    .I0(sig000001e3),
    .I1(sig00000217),
    .I2(sig00000312),
    .I3(sig0000030f),
    .I4(sig0000022e),
    .O(sig00000565)
  );
  LUT5 #(
    .INIT ( 32'h0AAA0CCC ))
  blk000007b7 (
    .I0(sig000001e4),
    .I1(sig00000218),
    .I2(sig00000312),
    .I3(sig0000030f),
    .I4(sig0000022e),
    .O(sig00000566)
  );
  LUT5 #(
    .INIT ( 32'h0AAA0CCC ))
  blk000007b8 (
    .I0(sig000001e5),
    .I1(sig00000219),
    .I2(sig00000312),
    .I3(sig0000030f),
    .I4(sig0000022e),
    .O(sig00000567)
  );
  LUT5 #(
    .INIT ( 32'h0AAA0CCC ))
  blk000007b9 (
    .I0(sig000001e6),
    .I1(sig0000021a),
    .I2(sig00000312),
    .I3(sig0000030f),
    .I4(sig0000022e),
    .O(sig00000568)
  );
  LUT5 #(
    .INIT ( 32'h0AAA0CCC ))
  blk000007ba (
    .I0(sig000001e7),
    .I1(sig0000021b),
    .I2(sig00000312),
    .I3(sig0000030f),
    .I4(sig0000022e),
    .O(sig00000569)
  );
  LUT5 #(
    .INIT ( 32'h0AAA0CCC ))
  blk000007bb (
    .I0(sig000001e8),
    .I1(sig0000021c),
    .I2(sig00000312),
    .I3(sig0000030f),
    .I4(sig0000022e),
    .O(sig0000056a)
  );
  LUT5 #(
    .INIT ( 32'h0AAA0CCC ))
  blk000007bc (
    .I0(sig000001e9),
    .I1(sig0000021d),
    .I2(sig00000312),
    .I3(sig0000030f),
    .I4(sig0000022e),
    .O(sig0000056b)
  );
  LUT5 #(
    .INIT ( 32'h0AAA0CCC ))
  blk000007bd (
    .I0(sig000001ea),
    .I1(sig0000021e),
    .I2(sig00000312),
    .I3(sig0000030f),
    .I4(sig0000022e),
    .O(sig0000056c)
  );
  LUT5 #(
    .INIT ( 32'h0AAA0CCC ))
  blk000007be (
    .I0(sig000001c6),
    .I1(sig000001fa),
    .I2(sig00000312),
    .I3(sig0000030f),
    .I4(sig0000022e),
    .O(sig00000548)
  );
  LUT5 #(
    .INIT ( 32'h0AAA0CCC ))
  blk000007bf (
    .I0(sig000001eb),
    .I1(sig0000021f),
    .I2(sig00000312),
    .I3(sig0000030f),
    .I4(sig0000022e),
    .O(sig0000056d)
  );
  LUT5 #(
    .INIT ( 32'h0AAA0CCC ))
  blk000007c0 (
    .I0(sig000001ec),
    .I1(sig00000220),
    .I2(sig00000312),
    .I3(sig0000030f),
    .I4(sig0000022e),
    .O(sig0000056e)
  );
  LUT5 #(
    .INIT ( 32'h0AAA0CCC ))
  blk000007c1 (
    .I0(sig000001ed),
    .I1(sig00000221),
    .I2(sig00000312),
    .I3(sig0000030f),
    .I4(sig0000022e),
    .O(sig0000056f)
  );
  LUT5 #(
    .INIT ( 32'h0AAA0CCC ))
  blk000007c2 (
    .I0(sig000001ee),
    .I1(sig00000222),
    .I2(sig00000312),
    .I3(sig0000030f),
    .I4(sig0000022e),
    .O(sig00000570)
  );
  LUT5 #(
    .INIT ( 32'h0AAA0CCC ))
  blk000007c3 (
    .I0(sig000001ef),
    .I1(sig00000223),
    .I2(sig00000312),
    .I3(sig0000030f),
    .I4(sig0000022e),
    .O(sig00000571)
  );
  LUT5 #(
    .INIT ( 32'h0AAA0CCC ))
  blk000007c4 (
    .I0(sig000001f0),
    .I1(sig00000224),
    .I2(sig00000312),
    .I3(sig0000030f),
    .I4(sig0000022e),
    .O(sig00000572)
  );
  LUT5 #(
    .INIT ( 32'h0AAA0CCC ))
  blk000007c5 (
    .I0(sig000001f1),
    .I1(sig00000225),
    .I2(sig00000312),
    .I3(sig0000030f),
    .I4(sig0000022e),
    .O(sig00000573)
  );
  LUT5 #(
    .INIT ( 32'h0AAA0CCC ))
  blk000007c6 (
    .I0(sig000001f2),
    .I1(sig00000226),
    .I2(sig00000312),
    .I3(sig0000030f),
    .I4(sig0000022e),
    .O(sig00000574)
  );
  LUT5 #(
    .INIT ( 32'h0AAA0CCC ))
  blk000007c7 (
    .I0(sig000001f3),
    .I1(sig00000227),
    .I2(sig00000312),
    .I3(sig0000030f),
    .I4(sig0000022e),
    .O(sig00000575)
  );
  LUT5 #(
    .INIT ( 32'h0AAA0CCC ))
  blk000007c8 (
    .I0(sig000001f4),
    .I1(sig00000228),
    .I2(sig00000312),
    .I3(sig0000030f),
    .I4(sig0000022e),
    .O(sig00000576)
  );
  LUT5 #(
    .INIT ( 32'h0AAA0CCC ))
  blk000007c9 (
    .I0(sig000001c7),
    .I1(sig000001fb),
    .I2(sig00000312),
    .I3(sig0000030f),
    .I4(sig0000022e),
    .O(sig00000549)
  );
  LUT5 #(
    .INIT ( 32'h0AAA0CCC ))
  blk000007ca (
    .I0(sig000001f5),
    .I1(sig00000229),
    .I2(sig00000312),
    .I3(sig0000030f),
    .I4(sig0000022e),
    .O(sig00000577)
  );
  LUT5 #(
    .INIT ( 32'h0AAA0CCC ))
  blk000007cb (
    .I0(sig000001f6),
    .I1(sig0000022a),
    .I2(sig00000312),
    .I3(sig0000030f),
    .I4(sig0000022e),
    .O(sig00000578)
  );
  LUT5 #(
    .INIT ( 32'h0AAA0CCC ))
  blk000007cc (
    .I0(sig000001c8),
    .I1(sig000001fc),
    .I2(sig00000312),
    .I3(sig0000030f),
    .I4(sig0000022e),
    .O(sig0000054a)
  );
  LUT5 #(
    .INIT ( 32'h0AAA0CCC ))
  blk000007cd (
    .I0(sig000001c9),
    .I1(sig000001fd),
    .I2(sig00000312),
    .I3(sig0000030f),
    .I4(sig0000022e),
    .O(sig0000054b)
  );
  LUT5 #(
    .INIT ( 32'h0AAA0CCC ))
  blk000007ce (
    .I0(sig000001ca),
    .I1(sig000001fe),
    .I2(sig00000312),
    .I3(sig0000030f),
    .I4(sig0000022e),
    .O(sig0000054c)
  );
  LUT5 #(
    .INIT ( 32'h0AAA0CCC ))
  blk000007cf (
    .I0(sig000001cb),
    .I1(sig000001ff),
    .I2(sig00000312),
    .I3(sig0000030f),
    .I4(sig0000022e),
    .O(sig0000054d)
  );
  LUT5 #(
    .INIT ( 32'h0AAA0CCC ))
  blk000007d0 (
    .I0(sig000001cc),
    .I1(sig00000200),
    .I2(sig00000312),
    .I3(sig0000030f),
    .I4(sig0000022e),
    .O(sig0000054e)
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  blk000007d1 (
    .I0(sig0000023f),
    .O(sig00000828)
  );
  INV   blk000007d2 (
    .I(sig0000023f),
    .O(sig00000543)
  );
  INV   blk000007d3 (
    .I(sig000002d1),
    .O(sig0000024c)
  );
  INV   blk000007d4 (
    .I(sig000002cd),
    .O(sig00000254)
  );
  INV   blk000007d5 (
    .I(sig000002ce),
    .O(sig00000252)
  );
  INV   blk000007d6 (
    .I(sig000002cf),
    .O(sig00000250)
  );
  INV   blk000007d7 (
    .I(sig000002d0),
    .O(sig0000024e)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000007d8 (
    .A0(sig000006c3),
    .A1(sig000006c3),
    .A2(sig000006c3),
    .A3(sig000006c3),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig0000027f),
    .Q(sig00000829),
    .Q15(NLW_blk000007d8_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000007d9 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000829),
    .Q(sig0000030d)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000007da (
    .A0(sig000006c3),
    .A1(sig00000001),
    .A2(sig00000001),
    .A3(sig000006c3),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000003b0),
    .Q(sig0000082a),
    .Q15(NLW_blk000007da_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000007db (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000082a),
    .Q(sig000002ec)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000007dc (
    .A0(sig000006c3),
    .A1(sig00000001),
    .A2(sig00000001),
    .A3(sig000006c3),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000003af),
    .Q(sig0000082b),
    .Q15(NLW_blk000007dc_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000007dd (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000082b),
    .Q(sig000002eb)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000007de (
    .A0(sig000006c3),
    .A1(sig00000001),
    .A2(sig00000001),
    .A3(sig000006c3),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000003b1),
    .Q(sig0000082c),
    .Q15(NLW_blk000007de_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000007df (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000082c),
    .Q(sig000002ea)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000007e0 (
    .A0(sig000006c3),
    .A1(sig00000001),
    .A2(sig00000001),
    .A3(sig000006c3),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000002dc),
    .Q(sig0000082d),
    .Q15(NLW_blk000007e0_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000007e1 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000082d),
    .Q(sig000002d1)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000007e2 (
    .A0(sig000006c3),
    .A1(sig00000001),
    .A2(sig00000001),
    .A3(sig000006c3),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000002db),
    .Q(sig0000082e),
    .Q15(NLW_blk000007e2_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000007e3 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000082e),
    .Q(sig000002d0)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000007e4 (
    .A0(sig000006c3),
    .A1(sig00000001),
    .A2(sig00000001),
    .A3(sig000006c3),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000002da),
    .Q(sig0000082f),
    .Q15(NLW_blk000007e4_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000007e5 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000082f),
    .Q(sig000002cf)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000007e6 (
    .A0(sig000006c3),
    .A1(sig00000001),
    .A2(sig00000001),
    .A3(sig000006c3),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000002d9),
    .Q(sig00000830),
    .Q15(NLW_blk000007e6_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000007e7 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000830),
    .Q(sig000002ce)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000007e8 (
    .A0(sig000006c3),
    .A1(sig00000001),
    .A2(sig00000001),
    .A3(sig000006c3),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000002d8),
    .Q(sig00000831),
    .Q15(NLW_blk000007e8_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000007e9 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000831),
    .Q(sig000002cd)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000007ea (
    .A0(sig000006c3),
    .A1(sig00000001),
    .A2(sig00000001),
    .A3(sig000006c3),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000002d7),
    .Q(sig00000832),
    .Q15(NLW_blk000007ea_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000007eb (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000832),
    .Q(sig000002cc)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000007ec (
    .A0(sig000006c3),
    .A1(sig00000001),
    .A2(sig00000001),
    .A3(sig000006c3),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000002d6),
    .Q(sig00000833),
    .Q15(NLW_blk000007ec_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000007ed (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000833),
    .Q(sig000002cb)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000007ee (
    .A0(sig000006c3),
    .A1(sig00000001),
    .A2(sig00000001),
    .A3(sig000006c3),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000002d3),
    .Q(sig00000834),
    .Q15(NLW_blk000007ee_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000007ef (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000834),
    .Q(sig000002c8)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000007f0 (
    .A0(sig000006c3),
    .A1(sig00000001),
    .A2(sig00000001),
    .A3(sig000006c3),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000002d5),
    .Q(sig00000835),
    .Q15(NLW_blk000007f0_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000007f1 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000835),
    .Q(sig000002ca)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000007f2 (
    .A0(sig000006c3),
    .A1(sig00000001),
    .A2(sig00000001),
    .A3(sig000006c3),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000002d4),
    .Q(sig00000836),
    .Q15(NLW_blk000007f2_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000007f3 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000836),
    .Q(sig000002c9)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000007f4 (
    .A0(sig000006c3),
    .A1(sig00000001),
    .A2(sig00000001),
    .A3(sig000006c3),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000002d2),
    .Q(sig00000837),
    .Q15(NLW_blk000007f4_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000007f5 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000837),
    .Q(sig000002c7)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000007f6 (
    .A0(sig00000001),
    .A1(sig000006c3),
    .A2(sig00000001),
    .A3(sig000006c3),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000003bd),
    .Q(sig00000838),
    .Q15(NLW_blk000007f6_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000007f7 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000838),
    .Q(sig000002c6)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000007f8 (
    .A0(sig000006c3),
    .A1(sig000006c3),
    .A2(sig000006c3),
    .A3(sig000006c3),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000003d3),
    .Q(sig00000839),
    .Q15(NLW_blk000007f8_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000007f9 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000839),
    .Q(sig0000018a)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000007fa (
    .A0(sig000006c3),
    .A1(sig000006c3),
    .A2(sig000006c3),
    .A3(sig000006c3),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000004cb),
    .Q(sig0000083a),
    .Q15(NLW_blk000007fa_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000007fb (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000083a),
    .Q(sig000005f8)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000007fc (
    .A0(sig00000001),
    .A1(sig000006c3),
    .A2(sig000006c3),
    .A3(sig000006c3),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig0000069d),
    .Q(sig0000083b),
    .Q15(NLW_blk000007fc_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000007fd (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000083b),
    .Q(sig00000606)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000007fe (
    .A0(sig00000001),
    .A1(sig000006c3),
    .A2(sig000006c3),
    .A3(sig000006c3),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig0000069f),
    .Q(sig0000083c),
    .Q15(NLW_blk000007fe_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000007ff (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000083c),
    .Q(sig00000608)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000800 (
    .A0(sig00000001),
    .A1(sig000006c3),
    .A2(sig000006c3),
    .A3(sig000006c3),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig0000069e),
    .Q(sig0000083d),
    .Q15(NLW_blk00000800_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000801 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000083d),
    .Q(sig00000607)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000802 (
    .A0(sig00000001),
    .A1(sig000006c3),
    .A2(sig000006c3),
    .A3(sig000006c3),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig0000069c),
    .Q(sig0000083e),
    .Q15(NLW_blk00000802_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000803 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000083e),
    .Q(sig00000605)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000804 (
    .A0(sig00000001),
    .A1(sig000006c3),
    .A2(sig000006c3),
    .A3(sig000006c3),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig0000069b),
    .Q(sig0000083f),
    .Q15(NLW_blk00000804_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000805 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000083f),
    .Q(sig00000604)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000806 (
    .A0(sig00000001),
    .A1(sig000006c3),
    .A2(sig000006c3),
    .A3(sig000006c3),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig0000069a),
    .Q(sig00000840),
    .Q15(NLW_blk00000806_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000807 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000840),
    .Q(sig00000603)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000808 (
    .A0(sig00000001),
    .A1(sig000006c3),
    .A2(sig000006c3),
    .A3(sig000006c3),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig00000699),
    .Q(sig00000841),
    .Q15(NLW_blk00000808_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000809 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000841),
    .Q(sig00000602)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk0000080a (
    .A0(sig000006c3),
    .A1(sig000006c3),
    .A2(sig000006c3),
    .A3(sig000006c3),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig00000119),
    .Q(sig00000842),
    .Q15(NLW_blk0000080a_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000080b (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000842),
    .Q(sig00000188)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk0000080c (
    .A0(sig00000001),
    .A1(sig000006c3),
    .A2(sig000006c3),
    .A3(sig000006c3),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig00000698),
    .Q(sig00000843),
    .Q15(NLW_blk0000080c_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000080d (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000843),
    .Q(sig00000601)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk0000080e (
    .A0(sig000006c3),
    .A1(sig000006c3),
    .A2(sig000006c3),
    .A3(sig000006c3),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig00000118),
    .Q(sig00000844),
    .Q15(NLW_blk0000080e_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000080f (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000844),
    .Q(sig00000189)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000810 (
    .A0(sig00000001),
    .A1(sig000006c3),
    .A2(sig000006c3),
    .A3(sig000006c3),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig0000018a),
    .Q(sig00000845),
    .Q15(NLW_blk00000810_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000811 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000845),
    .Q(sig00000155)
  );
  DSP48E #(
    .ACASCREG ( 2 ),
    .ALUMODEREG ( 0 ),
    .AREG ( 2 ),
    .AUTORESET_PATTERN_DETECT ( "FALSE" ),
    .AUTORESET_PATTERN_DETECT_OPTINV ( "MATCH" ),
    .A_INPUT ( "DIRECT" ),
    .BCASCREG ( 2 ),
    .BREG ( 2 ),
    .B_INPUT ( "DIRECT" ),
    .CARRYINREG ( 0 ),
    .CARRYINSELREG ( 0 ),
    .CREG ( 0 ),
    .MASK ( 48'h3FFFFFFFFFFF ),
    .MREG ( 0 ),
    .MULTCARRYINREG ( 0 ),
    .OPMODEREG ( 0 ),
    .PATTERN ( 48'h000000000000 ),
    .PREG ( 1 ),
    .SEL_MASK ( "MASK" ),
    .SEL_PATTERN ( "PATTERN" ),
    .SEL_ROUNDING_MASK ( "SEL_MASK" ),
    .SIM_MODE ( "SAFE" ),
    .USE_MULT ( "NONE" ),
    .USE_PATTERN_DETECT ( "NO_PATDET" ),
    .USE_SIMD ( "ONE48" ))
  blk00000812 (
    .CLK(clk),
    .PATTERNBDETECT(NLW_blk00000812_PATTERNBDETECT_UNCONNECTED),
    .RSTC(sig000006c3),
    .CEB1(sig00000001),
    .MULTSIGNOUT(NLW_blk00000812_MULTSIGNOUT_UNCONNECTED),
    .CEC(sig000006c3),
    .RSTM(sig000006c3),
    .MULTSIGNIN(sig000006c3),
    .CEB2(sig00000001),
    .RSTCTRL(sig000006c3),
    .CEP(sig00000001),
    .CARRYCASCOUT(NLW_blk00000812_CARRYCASCOUT_UNCONNECTED),
    .RSTA(sig000006c3),
    .CECARRYIN(sig000006c3),
    .UNDERFLOW(NLW_blk00000812_UNDERFLOW_UNCONNECTED),
    .PATTERNDETECT(NLW_blk00000812_PATTERNDETECT_UNCONNECTED),
    .RSTALUMODE(sig000006c3),
    .RSTALLCARRYIN(sig000006c3),
    .CEALUMODE(sig000006c3),
    .CEA2(sig00000001),
    .CEA1(sig00000001),
    .RSTB(sig000006c3),
    .CEMULTCARRYIN(sig000006c3),
    .OVERFLOW(NLW_blk00000812_OVERFLOW_UNCONNECTED),
    .CECTRL(sig000006c3),
    .CEM(sig000006c3),
    .CARRYIN(sig000006c3),
    .CARRYCASCIN(sig000006c3),
    .RSTP(sig000006c3),
    .CARRYINSEL({sig000006c3, sig000006c3, sig000006c3}),
    .OPMODE({sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig00000001, sig00000001}),
    .B({sig00000648, sig00000647, sig00000646, sig00000645, sig00000644, sig00000643, sig00000642, sig00000641, sig00000640, sig0000063f, sig0000063e
, sig0000063d, sig0000063c, sig0000063b, sig0000063a, sig00000639, sig000006c3, sig000006c3}),
    .A({sig000006c3, sig00000665, sig00000664, sig00000663, sig00000662, sig00000661, sig00000660, sig0000065f, sig0000065e, sig0000065d, sig0000065c
, sig0000065b, sig0000065a, sig00000659, sig00000658, sig00000657, sig00000656, sig00000655, sig00000654, sig00000653, sig00000652, sig00000651,
sig00000650, sig0000064f, sig0000064e, sig0000064d, sig0000064c, sig0000064b, sig0000064a, sig00000649}),
    .PCOUT({sig00000638, sig00000637, sig00000636, sig00000635, sig00000634, sig00000633, sig00000632, sig00000631, sig00000630, sig0000062f,
sig0000062e, sig0000062d, sig0000062c, sig0000062b, sig0000062a, sig00000629, sig00000628, sig00000627, sig00000626, sig00000625, sig00000624,
sig00000623, sig00000622, sig00000621, sig00000620, sig0000061f, sig0000061e, sig0000061d, sig0000061c, sig0000061b, sig0000061a, sig00000619,
sig00000618, sig00000617, sig00000616, sig00000615, sig00000614, sig00000613, sig00000612, sig00000611, sig00000610, sig0000060f, sig0000060e,
sig0000060d, sig0000060c, sig0000060b, sig0000060a, sig00000609}),
    .ACOUT({\NLW_blk00000812_ACOUT<29>_UNCONNECTED , \NLW_blk00000812_ACOUT<28>_UNCONNECTED , \NLW_blk00000812_ACOUT<27>_UNCONNECTED ,
\NLW_blk00000812_ACOUT<26>_UNCONNECTED , \NLW_blk00000812_ACOUT<25>_UNCONNECTED , \NLW_blk00000812_ACOUT<24>_UNCONNECTED ,
\NLW_blk00000812_ACOUT<23>_UNCONNECTED , \NLW_blk00000812_ACOUT<22>_UNCONNECTED , \NLW_blk00000812_ACOUT<21>_UNCONNECTED ,
\NLW_blk00000812_ACOUT<20>_UNCONNECTED , \NLW_blk00000812_ACOUT<19>_UNCONNECTED , \NLW_blk00000812_ACOUT<18>_UNCONNECTED ,
\NLW_blk00000812_ACOUT<17>_UNCONNECTED , \NLW_blk00000812_ACOUT<16>_UNCONNECTED , \NLW_blk00000812_ACOUT<15>_UNCONNECTED ,
\NLW_blk00000812_ACOUT<14>_UNCONNECTED , \NLW_blk00000812_ACOUT<13>_UNCONNECTED , \NLW_blk00000812_ACOUT<12>_UNCONNECTED ,
\NLW_blk00000812_ACOUT<11>_UNCONNECTED , \NLW_blk00000812_ACOUT<10>_UNCONNECTED , \NLW_blk00000812_ACOUT<9>_UNCONNECTED ,
\NLW_blk00000812_ACOUT<8>_UNCONNECTED , \NLW_blk00000812_ACOUT<7>_UNCONNECTED , \NLW_blk00000812_ACOUT<6>_UNCONNECTED ,
\NLW_blk00000812_ACOUT<5>_UNCONNECTED , \NLW_blk00000812_ACOUT<4>_UNCONNECTED , \NLW_blk00000812_ACOUT<3>_UNCONNECTED ,
\NLW_blk00000812_ACOUT<2>_UNCONNECTED , \NLW_blk00000812_ACOUT<1>_UNCONNECTED , \NLW_blk00000812_ACOUT<0>_UNCONNECTED }),
    .PCIN({sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3,
sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3,
sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3,
sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3,
sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3}),
    .ALUMODE({sig000006c3, sig000006c3, sig000006c3, sig000006c3}),
    .C({sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3
, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3,
sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3,
sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3,
sig000006c3, sig000006c3, sig000006c3, sig000006c3}),
    .CARRYOUT({\NLW_blk00000812_CARRYOUT<3>_UNCONNECTED , \NLW_blk00000812_CARRYOUT<2>_UNCONNECTED , \NLW_blk00000812_CARRYOUT<1>_UNCONNECTED ,
\NLW_blk00000812_CARRYOUT<0>_UNCONNECTED }),
    .BCIN({sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3,
sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3}),
    .BCOUT({\NLW_blk00000812_BCOUT<17>_UNCONNECTED , \NLW_blk00000812_BCOUT<16>_UNCONNECTED , \NLW_blk00000812_BCOUT<15>_UNCONNECTED ,
\NLW_blk00000812_BCOUT<14>_UNCONNECTED , \NLW_blk00000812_BCOUT<13>_UNCONNECTED , \NLW_blk00000812_BCOUT<12>_UNCONNECTED ,
\NLW_blk00000812_BCOUT<11>_UNCONNECTED , \NLW_blk00000812_BCOUT<10>_UNCONNECTED , \NLW_blk00000812_BCOUT<9>_UNCONNECTED ,
\NLW_blk00000812_BCOUT<8>_UNCONNECTED , \NLW_blk00000812_BCOUT<7>_UNCONNECTED , \NLW_blk00000812_BCOUT<6>_UNCONNECTED ,
\NLW_blk00000812_BCOUT<5>_UNCONNECTED , \NLW_blk00000812_BCOUT<4>_UNCONNECTED , \NLW_blk00000812_BCOUT<3>_UNCONNECTED ,
\NLW_blk00000812_BCOUT<2>_UNCONNECTED , \NLW_blk00000812_BCOUT<1>_UNCONNECTED , \NLW_blk00000812_BCOUT<0>_UNCONNECTED }),
    .P({\NLW_blk00000812_P<47>_UNCONNECTED , \NLW_blk00000812_P<46>_UNCONNECTED , \NLW_blk00000812_P<45>_UNCONNECTED ,
\NLW_blk00000812_P<44>_UNCONNECTED , \NLW_blk00000812_P<43>_UNCONNECTED , \NLW_blk00000812_P<42>_UNCONNECTED , \NLW_blk00000812_P<41>_UNCONNECTED ,
\NLW_blk00000812_P<40>_UNCONNECTED , \NLW_blk00000812_P<39>_UNCONNECTED , \NLW_blk00000812_P<38>_UNCONNECTED , \NLW_blk00000812_P<37>_UNCONNECTED ,
\NLW_blk00000812_P<36>_UNCONNECTED , \NLW_blk00000812_P<35>_UNCONNECTED , \NLW_blk00000812_P<34>_UNCONNECTED , \NLW_blk00000812_P<33>_UNCONNECTED ,
\NLW_blk00000812_P<32>_UNCONNECTED , \NLW_blk00000812_P<31>_UNCONNECTED , \NLW_blk00000812_P<30>_UNCONNECTED , \NLW_blk00000812_P<29>_UNCONNECTED ,
\NLW_blk00000812_P<28>_UNCONNECTED , \NLW_blk00000812_P<27>_UNCONNECTED , \NLW_blk00000812_P<26>_UNCONNECTED , \NLW_blk00000812_P<25>_UNCONNECTED ,
\NLW_blk00000812_P<24>_UNCONNECTED , \NLW_blk00000812_P<23>_UNCONNECTED , \NLW_blk00000812_P<22>_UNCONNECTED , \NLW_blk00000812_P<21>_UNCONNECTED ,
\NLW_blk00000812_P<20>_UNCONNECTED , \NLW_blk00000812_P<19>_UNCONNECTED , \NLW_blk00000812_P<18>_UNCONNECTED , \NLW_blk00000812_P<17>_UNCONNECTED ,
\NLW_blk00000812_P<16>_UNCONNECTED , \NLW_blk00000812_P<15>_UNCONNECTED , \NLW_blk00000812_P<14>_UNCONNECTED , \NLW_blk00000812_P<13>_UNCONNECTED ,
\NLW_blk00000812_P<12>_UNCONNECTED , \NLW_blk00000812_P<11>_UNCONNECTED , \NLW_blk00000812_P<10>_UNCONNECTED , \NLW_blk00000812_P<9>_UNCONNECTED ,
\NLW_blk00000812_P<8>_UNCONNECTED , \NLW_blk00000812_P<7>_UNCONNECTED , \NLW_blk00000812_P<6>_UNCONNECTED , \NLW_blk00000812_P<5>_UNCONNECTED ,
\NLW_blk00000812_P<4>_UNCONNECTED , \NLW_blk00000812_P<3>_UNCONNECTED , \NLW_blk00000812_P<2>_UNCONNECTED , \NLW_blk00000812_P<1>_UNCONNECTED ,
\NLW_blk00000812_P<0>_UNCONNECTED }),
    .ACIN({sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3,
sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3,
sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3})
  );
  DSP48E #(
    .ACASCREG ( 1 ),
    .ALUMODEREG ( 1 ),
    .AREG ( 1 ),
    .AUTORESET_PATTERN_DETECT ( "FALSE" ),
    .AUTORESET_PATTERN_DETECT_OPTINV ( "MATCH" ),
    .A_INPUT ( "DIRECT" ),
    .BCASCREG ( 1 ),
    .BREG ( 1 ),
    .B_INPUT ( "DIRECT" ),
    .CARRYINREG ( 1 ),
    .CARRYINSELREG ( 1 ),
    .CREG ( 1 ),
    .MASK ( 48'h3FFFFFFFFFFF ),
    .MREG ( 0 ),
    .MULTCARRYINREG ( 0 ),
    .OPMODEREG ( 1 ),
    .PATTERN ( 48'h000000000000 ),
    .PREG ( 1 ),
    .SEL_MASK ( "MASK" ),
    .SEL_PATTERN ( "PATTERN" ),
    .SEL_ROUNDING_MASK ( "SEL_MASK" ),
    .SIM_MODE ( "SAFE" ),
    .USE_MULT ( "NONE" ),
    .USE_PATTERN_DETECT ( "NO_PATDET" ),
    .USE_SIMD ( "ONE48" ))
  blk00000813 (
    .RSTALLCARRYIN(sig000004cc),
    .CLK(clk),
    .CARRYIN(sig0000050d),
    .PATTERNBDETECT(NLW_blk00000813_PATTERNBDETECT_UNCONNECTED),
    .RSTC(sig000006c3),
    .CEB1(sig000006c3),
    .MULTSIGNOUT(NLW_blk00000813_MULTSIGNOUT_UNCONNECTED),
    .CEC(sig00000001),
    .RSTM(sig000006c3),
    .MULTSIGNIN(sig000006c3),
    .CEB2(sig00000001),
    .RSTCTRL(sig000006c3),
    .CEP(sig00000001),
    .CARRYCASCOUT(NLW_blk00000813_CARRYCASCOUT_UNCONNECTED),
    .RSTA(sig000006c3),
    .CECARRYIN(sig00000001),
    .UNDERFLOW(NLW_blk00000813_UNDERFLOW_UNCONNECTED),
    .PATTERNDETECT(NLW_blk00000813_PATTERNDETECT_UNCONNECTED),
    .RSTALUMODE(sig000006c3),
    .CEALUMODE(sig00000001),
    .CEA2(sig00000001),
    .CEA1(sig000006c3),
    .RSTB(sig000006c3),
    .CEMULTCARRYIN(sig000006c3),
    .OVERFLOW(NLW_blk00000813_OVERFLOW_UNCONNECTED),
    .CECTRL(sig00000001),
    .CEM(sig000006c3),
    .CARRYCASCIN(sig000006c3),
    .RSTP(sig000006c3),
    .CARRYINSEL({sig000006c3, sig000006c3, sig000006c3}),
    .OPMODE({sig000006c3, sig000006c3, sig00000001, sig000004c7, sig000004c7, sig000004c8, sig000004c8}),
    .PCIN({sig00000638, sig00000637, sig00000636, sig00000635, sig00000634, sig00000633, sig00000632, sig00000631, sig00000630, sig0000062f,
sig0000062e, sig0000062d, sig0000062c, sig0000062b, sig0000062a, sig00000629, sig00000628, sig00000627, sig00000626, sig00000625, sig00000624,
sig00000623, sig00000622, sig00000621, sig00000620, sig0000061f, sig0000061e, sig0000061d, sig0000061c, sig0000061b, sig0000061a, sig00000619,
sig00000618, sig00000617, sig00000616, sig00000615, sig00000614, sig00000613, sig00000612, sig00000611, sig00000610, sig0000060f, sig0000060e,
sig0000060d, sig0000060c, sig0000060b, sig0000060a, sig00000609}),
    .A({sig000004c9, sig00000485, sig00000486, sig00000487, sig00000488, sig00000489, sig0000048a, sig0000048b, sig0000048c, sig0000048d, sig0000048e
, sig0000048f, sig00000490, sig00000491, sig00000492, sig00000493, sig00000494, sig00000495, sig00000496, sig00000497, sig00000498, sig00000499,
sig0000049a, sig0000049b, sig0000049c, sig0000049d, sig0000049e, sig0000049f, sig000004a0, sig000004a1}),
    .C({sig000004c9, sig00000483, sig00000484, sig00000485, sig00000486, sig00000487, sig00000488, sig00000489, sig0000048a, sig0000048b, sig0000048c
, sig0000048d, sig0000048e, sig0000048f, sig00000490, sig00000491, sig00000492, sig00000493, sig00000494, sig00000495, sig00000496, sig00000497,
sig00000498, sig00000499, sig0000049a, sig0000049b, sig0000049c, sig0000049d, sig0000049e, sig0000049f, sig000004a0, sig000004a1, sig000004a2,
sig000004a3, sig000004a4, sig000004a5, sig000004a6, sig000004a7, sig000004a8, sig000004a9, sig000004aa, sig000004ab, sig000004ac, sig000004ad,
sig000004ae, sig000004af, sig000004b0, sig000004b1}),
    .B({sig000004a2, sig000004a3, sig000004a4, sig000004a5, sig000004a6, sig000004a7, sig000004a8, sig000004a9, sig000004aa, sig000004ab, sig000004ac
, sig000004ad, sig000004ae, sig000004af, sig000004b0, sig000004b1, sig000004b2, sig000004b3}),
    .P({sig00000666, sig00000695, sig00000694, sig00000693, sig00000692, sig00000691, sig00000690, sig0000068f, sig0000068e, sig0000068d, sig0000068c
, sig0000068b, sig0000068a, sig00000689, sig00000688, sig00000687, sig00000686, sig00000685, sig00000684, sig00000683, sig00000682, sig00000681,
sig00000680, sig0000067f, sig0000067e, sig0000067d, sig0000067c, sig0000067b, sig0000067a, sig00000679, sig00000678, sig00000677, sig00000676,
sig00000675, sig00000674, sig00000673, sig00000672, sig00000671, sig00000670, sig0000066f, sig0000066e, sig0000066d, sig0000066c, sig0000066b,
sig0000066a, sig00000669, sig00000668, sig00000667}),
    .ACOUT({\NLW_blk00000813_ACOUT<29>_UNCONNECTED , \NLW_blk00000813_ACOUT<28>_UNCONNECTED , \NLW_blk00000813_ACOUT<27>_UNCONNECTED ,
\NLW_blk00000813_ACOUT<26>_UNCONNECTED , \NLW_blk00000813_ACOUT<25>_UNCONNECTED , \NLW_blk00000813_ACOUT<24>_UNCONNECTED ,
\NLW_blk00000813_ACOUT<23>_UNCONNECTED , \NLW_blk00000813_ACOUT<22>_UNCONNECTED , \NLW_blk00000813_ACOUT<21>_UNCONNECTED ,
\NLW_blk00000813_ACOUT<20>_UNCONNECTED , \NLW_blk00000813_ACOUT<19>_UNCONNECTED , \NLW_blk00000813_ACOUT<18>_UNCONNECTED ,
\NLW_blk00000813_ACOUT<17>_UNCONNECTED , \NLW_blk00000813_ACOUT<16>_UNCONNECTED , \NLW_blk00000813_ACOUT<15>_UNCONNECTED ,
\NLW_blk00000813_ACOUT<14>_UNCONNECTED , \NLW_blk00000813_ACOUT<13>_UNCONNECTED , \NLW_blk00000813_ACOUT<12>_UNCONNECTED ,
\NLW_blk00000813_ACOUT<11>_UNCONNECTED , \NLW_blk00000813_ACOUT<10>_UNCONNECTED , \NLW_blk00000813_ACOUT<9>_UNCONNECTED ,
\NLW_blk00000813_ACOUT<8>_UNCONNECTED , \NLW_blk00000813_ACOUT<7>_UNCONNECTED , \NLW_blk00000813_ACOUT<6>_UNCONNECTED ,
\NLW_blk00000813_ACOUT<5>_UNCONNECTED , \NLW_blk00000813_ACOUT<4>_UNCONNECTED , \NLW_blk00000813_ACOUT<3>_UNCONNECTED ,
\NLW_blk00000813_ACOUT<2>_UNCONNECTED , \NLW_blk00000813_ACOUT<1>_UNCONNECTED , \NLW_blk00000813_ACOUT<0>_UNCONNECTED }),
    .ALUMODE({sig000006c3, sig000006c3, sig000004c9, sig000004c9}),
    .CARRYOUT({\NLW_blk00000813_CARRYOUT<3>_UNCONNECTED , \NLW_blk00000813_CARRYOUT<2>_UNCONNECTED , \NLW_blk00000813_CARRYOUT<1>_UNCONNECTED ,
\NLW_blk00000813_CARRYOUT<0>_UNCONNECTED }),
    .BCIN({sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3,
sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3}),
    .BCOUT({\NLW_blk00000813_BCOUT<17>_UNCONNECTED , \NLW_blk00000813_BCOUT<16>_UNCONNECTED , \NLW_blk00000813_BCOUT<15>_UNCONNECTED ,
\NLW_blk00000813_BCOUT<14>_UNCONNECTED , \NLW_blk00000813_BCOUT<13>_UNCONNECTED , \NLW_blk00000813_BCOUT<12>_UNCONNECTED ,
\NLW_blk00000813_BCOUT<11>_UNCONNECTED , \NLW_blk00000813_BCOUT<10>_UNCONNECTED , \NLW_blk00000813_BCOUT<9>_UNCONNECTED ,
\NLW_blk00000813_BCOUT<8>_UNCONNECTED , \NLW_blk00000813_BCOUT<7>_UNCONNECTED , \NLW_blk00000813_BCOUT<6>_UNCONNECTED ,
\NLW_blk00000813_BCOUT<5>_UNCONNECTED , \NLW_blk00000813_BCOUT<4>_UNCONNECTED , \NLW_blk00000813_BCOUT<3>_UNCONNECTED ,
\NLW_blk00000813_BCOUT<2>_UNCONNECTED , \NLW_blk00000813_BCOUT<1>_UNCONNECTED , \NLW_blk00000813_BCOUT<0>_UNCONNECTED }),
    .PCOUT({\NLW_blk00000813_PCOUT<47>_UNCONNECTED , \NLW_blk00000813_PCOUT<46>_UNCONNECTED , \NLW_blk00000813_PCOUT<45>_UNCONNECTED ,
\NLW_blk00000813_PCOUT<44>_UNCONNECTED , \NLW_blk00000813_PCOUT<43>_UNCONNECTED , \NLW_blk00000813_PCOUT<42>_UNCONNECTED ,
\NLW_blk00000813_PCOUT<41>_UNCONNECTED , \NLW_blk00000813_PCOUT<40>_UNCONNECTED , \NLW_blk00000813_PCOUT<39>_UNCONNECTED ,
\NLW_blk00000813_PCOUT<38>_UNCONNECTED , \NLW_blk00000813_PCOUT<37>_UNCONNECTED , \NLW_blk00000813_PCOUT<36>_UNCONNECTED ,
\NLW_blk00000813_PCOUT<35>_UNCONNECTED , \NLW_blk00000813_PCOUT<34>_UNCONNECTED , \NLW_blk00000813_PCOUT<33>_UNCONNECTED ,
\NLW_blk00000813_PCOUT<32>_UNCONNECTED , \NLW_blk00000813_PCOUT<31>_UNCONNECTED , \NLW_blk00000813_PCOUT<30>_UNCONNECTED ,
\NLW_blk00000813_PCOUT<29>_UNCONNECTED , \NLW_blk00000813_PCOUT<28>_UNCONNECTED , \NLW_blk00000813_PCOUT<27>_UNCONNECTED ,
\NLW_blk00000813_PCOUT<26>_UNCONNECTED , \NLW_blk00000813_PCOUT<25>_UNCONNECTED , \NLW_blk00000813_PCOUT<24>_UNCONNECTED ,
\NLW_blk00000813_PCOUT<23>_UNCONNECTED , \NLW_blk00000813_PCOUT<22>_UNCONNECTED , \NLW_blk00000813_PCOUT<21>_UNCONNECTED ,
\NLW_blk00000813_PCOUT<20>_UNCONNECTED , \NLW_blk00000813_PCOUT<19>_UNCONNECTED , \NLW_blk00000813_PCOUT<18>_UNCONNECTED ,
\NLW_blk00000813_PCOUT<17>_UNCONNECTED , \NLW_blk00000813_PCOUT<16>_UNCONNECTED , \NLW_blk00000813_PCOUT<15>_UNCONNECTED ,
\NLW_blk00000813_PCOUT<14>_UNCONNECTED , \NLW_blk00000813_PCOUT<13>_UNCONNECTED , \NLW_blk00000813_PCOUT<12>_UNCONNECTED ,
\NLW_blk00000813_PCOUT<11>_UNCONNECTED , \NLW_blk00000813_PCOUT<10>_UNCONNECTED , \NLW_blk00000813_PCOUT<9>_UNCONNECTED ,
\NLW_blk00000813_PCOUT<8>_UNCONNECTED , \NLW_blk00000813_PCOUT<7>_UNCONNECTED , \NLW_blk00000813_PCOUT<6>_UNCONNECTED ,
\NLW_blk00000813_PCOUT<5>_UNCONNECTED , \NLW_blk00000813_PCOUT<4>_UNCONNECTED , \NLW_blk00000813_PCOUT<3>_UNCONNECTED ,
\NLW_blk00000813_PCOUT<2>_UNCONNECTED , \NLW_blk00000813_PCOUT<1>_UNCONNECTED , \NLW_blk00000813_PCOUT<0>_UNCONNECTED }),
    .ACIN({sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3,
sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3,
sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3})
  );
  DSP48E #(
    .ACASCREG ( 0 ),
    .ALUMODEREG ( 1 ),
    .AREG ( 0 ),
    .AUTORESET_PATTERN_DETECT ( "FALSE" ),
    .AUTORESET_PATTERN_DETECT_OPTINV ( "MATCH" ),
    .A_INPUT ( "DIRECT" ),
    .BCASCREG ( 1 ),
    .BREG ( 1 ),
    .B_INPUT ( "DIRECT" ),
    .CARRYINREG ( 1 ),
    .CARRYINSELREG ( 1 ),
    .CREG ( 1 ),
    .MASK ( 48'h3FFFFFFFFFFF ),
    .MREG ( 0 ),
    .MULTCARRYINREG ( 0 ),
    .OPMODEREG ( 1 ),
    .PATTERN ( 48'h000000000000 ),
    .PREG ( 1 ),
    .SEL_MASK ( "MASK" ),
    .SEL_PATTERN ( "PATTERN" ),
    .SEL_ROUNDING_MASK ( "SEL_MASK" ),
    .SIM_MODE ( "SAFE" ),
    .USE_MULT ( "NONE" ),
    .USE_PATTERN_DETECT ( "NO_PATDET" ),
    .USE_SIMD ( "ONE48" ))
  blk00000814 (
    .CLK(clk),
    .PATTERNBDETECT(NLW_blk00000814_PATTERNBDETECT_UNCONNECTED),
    .RSTC(sig000006c3),
    .CEB1(sig000006c3),
    .MULTSIGNOUT(NLW_blk00000814_MULTSIGNOUT_UNCONNECTED),
    .CEC(sig00000001),
    .RSTM(sig000006c3),
    .MULTSIGNIN(sig000006c3),
    .CEB2(sig00000001),
    .RSTCTRL(sig000006c3),
    .CEP(sig00000001),
    .CARRYCASCOUT(NLW_blk00000814_CARRYCASCOUT_UNCONNECTED),
    .RSTA(sig000006c3),
    .CECARRYIN(sig00000001),
    .UNDERFLOW(NLW_blk00000814_UNDERFLOW_UNCONNECTED),
    .PATTERNDETECT(NLW_blk00000814_PATTERNDETECT_UNCONNECTED),
    .RSTALUMODE(sig000006c3),
    .RSTALLCARRYIN(sig000006c3),
    .CEALUMODE(sig00000001),
    .CEA2(sig000006c3),
    .CEA1(sig000006c3),
    .RSTB(sig000006c3),
    .CEMULTCARRYIN(sig000006c3),
    .OVERFLOW(NLW_blk00000814_OVERFLOW_UNCONNECTED),
    .CECTRL(sig00000001),
    .CEM(sig000006c3),
    .CARRYIN(sig000006c3),
    .CARRYCASCIN(sig000006c3),
    .RSTP(sig000006c3),
    .CARRYINSEL({sig000006c3, sig000006c3, sig000006c3}),
    .OPMODE({sig000006c3, sig00000001, sig00000001, sig000006c3, sig000006c3, sig00000001, sig00000001}),
    .C({sig000006c3, sig00000752, sig0000079d, sig0000079c, sig0000079b, sig0000079a, sig00000799, sig00000798, sig00000797, sig00000796, sig00000795
, sig00000794, sig00000793, sig00000792, sig00000791, sig00000790, sig0000078f, sig0000078e, sig0000078d, sig0000078c, sig0000078b, sig0000078a,
sig00000789, sig00000788, sig00000787, sig00000786, sig00000785, sig00000784, sig00000783, sig00000782, sig00000781, sig00000780, sig0000077f,
sig0000077e, sig0000077d, sig0000077c, sig0000077b, sig0000077a, sig00000779, sig00000778, sig00000777, sig00000776, sig00000775, sig00000774,
sig00000773, sig00000772, sig00000771, sig00000770}),
    .B({sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3
, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig00000768, sig000006c3}),
    .P({sig00000767, sig00000185, sig00000184, sig00000183, sig00000182, sig00000181, sig00000180, sig0000017f, sig0000017e, sig0000017d, sig0000017c
, sig0000017b, sig0000017a, sig00000179, sig00000178, sig00000177, sig00000176, sig00000175, sig00000174, sig00000173, sig00000172, sig00000171,
sig00000170, sig0000016f, sig0000016e, sig0000016d, sig0000016c, sig0000016b, sig0000016a, sig00000169, sig00000168, sig00000167, sig00000166,
sig00000165, sig00000164, sig00000163, sig00000162, sig00000161, sig00000160, sig0000015f, sig0000015e, sig0000015d, sig0000015c, sig0000015b,
sig0000015a, sig00000159, sig00000158, \NLW_blk00000814_P<0>_UNCONNECTED }),
    .ACOUT({\NLW_blk00000814_ACOUT<29>_UNCONNECTED , \NLW_blk00000814_ACOUT<28>_UNCONNECTED , \NLW_blk00000814_ACOUT<27>_UNCONNECTED ,
\NLW_blk00000814_ACOUT<26>_UNCONNECTED , \NLW_blk00000814_ACOUT<25>_UNCONNECTED , \NLW_blk00000814_ACOUT<24>_UNCONNECTED ,
\NLW_blk00000814_ACOUT<23>_UNCONNECTED , \NLW_blk00000814_ACOUT<22>_UNCONNECTED , \NLW_blk00000814_ACOUT<21>_UNCONNECTED ,
\NLW_blk00000814_ACOUT<20>_UNCONNECTED , \NLW_blk00000814_ACOUT<19>_UNCONNECTED , \NLW_blk00000814_ACOUT<18>_UNCONNECTED ,
\NLW_blk00000814_ACOUT<17>_UNCONNECTED , \NLW_blk00000814_ACOUT<16>_UNCONNECTED , \NLW_blk00000814_ACOUT<15>_UNCONNECTED ,
\NLW_blk00000814_ACOUT<14>_UNCONNECTED , \NLW_blk00000814_ACOUT<13>_UNCONNECTED , \NLW_blk00000814_ACOUT<12>_UNCONNECTED ,
\NLW_blk00000814_ACOUT<11>_UNCONNECTED , \NLW_blk00000814_ACOUT<10>_UNCONNECTED , \NLW_blk00000814_ACOUT<9>_UNCONNECTED ,
\NLW_blk00000814_ACOUT<8>_UNCONNECTED , \NLW_blk00000814_ACOUT<7>_UNCONNECTED , \NLW_blk00000814_ACOUT<6>_UNCONNECTED ,
\NLW_blk00000814_ACOUT<5>_UNCONNECTED , \NLW_blk00000814_ACOUT<4>_UNCONNECTED , \NLW_blk00000814_ACOUT<3>_UNCONNECTED ,
\NLW_blk00000814_ACOUT<2>_UNCONNECTED , \NLW_blk00000814_ACOUT<1>_UNCONNECTED , \NLW_blk00000814_ACOUT<0>_UNCONNECTED }),
    .PCIN({sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3,
sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3,
sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3,
sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3,
sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3}),
    .ALUMODE({sig000006c3, sig000006c3, sig000006c3, sig000006c3}),
    .CARRYOUT({\NLW_blk00000814_CARRYOUT<3>_UNCONNECTED , \NLW_blk00000814_CARRYOUT<2>_UNCONNECTED , \NLW_blk00000814_CARRYOUT<1>_UNCONNECTED ,
\NLW_blk00000814_CARRYOUT<0>_UNCONNECTED }),
    .BCIN({sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3,
sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3}),
    .BCOUT({\NLW_blk00000814_BCOUT<17>_UNCONNECTED , \NLW_blk00000814_BCOUT<16>_UNCONNECTED , \NLW_blk00000814_BCOUT<15>_UNCONNECTED ,
\NLW_blk00000814_BCOUT<14>_UNCONNECTED , \NLW_blk00000814_BCOUT<13>_UNCONNECTED , \NLW_blk00000814_BCOUT<12>_UNCONNECTED ,
\NLW_blk00000814_BCOUT<11>_UNCONNECTED , \NLW_blk00000814_BCOUT<10>_UNCONNECTED , \NLW_blk00000814_BCOUT<9>_UNCONNECTED ,
\NLW_blk00000814_BCOUT<8>_UNCONNECTED , \NLW_blk00000814_BCOUT<7>_UNCONNECTED , \NLW_blk00000814_BCOUT<6>_UNCONNECTED ,
\NLW_blk00000814_BCOUT<5>_UNCONNECTED , \NLW_blk00000814_BCOUT<4>_UNCONNECTED , \NLW_blk00000814_BCOUT<3>_UNCONNECTED ,
\NLW_blk00000814_BCOUT<2>_UNCONNECTED , \NLW_blk00000814_BCOUT<1>_UNCONNECTED , \NLW_blk00000814_BCOUT<0>_UNCONNECTED }),
    .A({sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3
, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3,
sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3}),
    .PCOUT({\NLW_blk00000814_PCOUT<47>_UNCONNECTED , \NLW_blk00000814_PCOUT<46>_UNCONNECTED , \NLW_blk00000814_PCOUT<45>_UNCONNECTED ,
\NLW_blk00000814_PCOUT<44>_UNCONNECTED , \NLW_blk00000814_PCOUT<43>_UNCONNECTED , \NLW_blk00000814_PCOUT<42>_UNCONNECTED ,
\NLW_blk00000814_PCOUT<41>_UNCONNECTED , \NLW_blk00000814_PCOUT<40>_UNCONNECTED , \NLW_blk00000814_PCOUT<39>_UNCONNECTED ,
\NLW_blk00000814_PCOUT<38>_UNCONNECTED , \NLW_blk00000814_PCOUT<37>_UNCONNECTED , \NLW_blk00000814_PCOUT<36>_UNCONNECTED ,
\NLW_blk00000814_PCOUT<35>_UNCONNECTED , \NLW_blk00000814_PCOUT<34>_UNCONNECTED , \NLW_blk00000814_PCOUT<33>_UNCONNECTED ,
\NLW_blk00000814_PCOUT<32>_UNCONNECTED , \NLW_blk00000814_PCOUT<31>_UNCONNECTED , \NLW_blk00000814_PCOUT<30>_UNCONNECTED ,
\NLW_blk00000814_PCOUT<29>_UNCONNECTED , \NLW_blk00000814_PCOUT<28>_UNCONNECTED , \NLW_blk00000814_PCOUT<27>_UNCONNECTED ,
\NLW_blk00000814_PCOUT<26>_UNCONNECTED , \NLW_blk00000814_PCOUT<25>_UNCONNECTED , \NLW_blk00000814_PCOUT<24>_UNCONNECTED ,
\NLW_blk00000814_PCOUT<23>_UNCONNECTED , \NLW_blk00000814_PCOUT<22>_UNCONNECTED , \NLW_blk00000814_PCOUT<21>_UNCONNECTED ,
\NLW_blk00000814_PCOUT<20>_UNCONNECTED , \NLW_blk00000814_PCOUT<19>_UNCONNECTED , \NLW_blk00000814_PCOUT<18>_UNCONNECTED ,
\NLW_blk00000814_PCOUT<17>_UNCONNECTED , \NLW_blk00000814_PCOUT<16>_UNCONNECTED , \NLW_blk00000814_PCOUT<15>_UNCONNECTED ,
\NLW_blk00000814_PCOUT<14>_UNCONNECTED , \NLW_blk00000814_PCOUT<13>_UNCONNECTED , \NLW_blk00000814_PCOUT<12>_UNCONNECTED ,
\NLW_blk00000814_PCOUT<11>_UNCONNECTED , \NLW_blk00000814_PCOUT<10>_UNCONNECTED , \NLW_blk00000814_PCOUT<9>_UNCONNECTED ,
\NLW_blk00000814_PCOUT<8>_UNCONNECTED , \NLW_blk00000814_PCOUT<7>_UNCONNECTED , \NLW_blk00000814_PCOUT<6>_UNCONNECTED ,
\NLW_blk00000814_PCOUT<5>_UNCONNECTED , \NLW_blk00000814_PCOUT<4>_UNCONNECTED , \NLW_blk00000814_PCOUT<3>_UNCONNECTED ,
\NLW_blk00000814_PCOUT<2>_UNCONNECTED , \NLW_blk00000814_PCOUT<1>_UNCONNECTED , \NLW_blk00000814_PCOUT<0>_UNCONNECTED }),
    .ACIN({sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3,
sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3,
sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3, sig000006c3})
  );
// synthesis translate_on
endmodule