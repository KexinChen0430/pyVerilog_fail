module srio_gen2_0_GT #
(
    // Simulation attributes
    parameter   GT_SIM_GTRESET_SPEEDUP   =   "FALSE",       // Set to "TRUE" to speed up sim reset;
    parameter   RX_DFE_KL_CFG2_IN        =   32'h301148AC,
    parameter   PMA_RSV_IN               =   32'h00018480,
    parameter   PCS_RSVD_ATTR_IN         =   48'h000000000000
)
(
    output          cpllfbclklost_out,
    output          cplllock_out,
    input           cplllockdetclk_in,
    output          cpllrefclklost_out,
    input           cpllreset_in,
    input           gtrefclk0_in,
    input   [8:0]   drpaddr_in,
    input           drpclk_in,
    input   [15:0]  drpdi_in,
    output  [15:0]  drpdo_out,
    input           drpen_in,
    output          drprdy_out,
    input           drpwe_in,
    input           qpllclk_in,
    input           qpllrefclk_in,
    output  [7:0]   dmonitorout_out,
    input   [2:0]   loopback_in,
    input           eyescanreset_in,
    input           rxuserrdy_in,
    output          eyescandataerror_out,
    input           eyescantrigger_in,
    input           rxcdrhold_in,
    output  [1:0]   rxclkcorcnt_out,
    input           rxusrclk_in,
    input           rxusrclk2_in,
    output  [31:0]  rxdata_out,
    output          rxprbserr_out,
    input   [2:0]   rxprbssel_in,
    input           rxprbscntreset_in,
    output  [3:0]   rxdisperr_out,
    output  [3:0]   rxnotintable_out,
    input           gtxrxp_in,
    input           gtxrxn_in,
    input           rxbufreset_in,
    output  [2:0]   rxbufstatus_out,
    output          rxbyteisaligned_out,
    output          rxbyterealign_out,
    output          rxcommadet_out,
    input           rxmcommaalignen_in,
    input           rxpcommaalignen_in,
    output          rxchanbondseq_out,
    input           rxchbonden_in,
    input   [2:0]   rxchbondlevel_in,
    input           rxchbondmaster_in,
    output  [4:0]   rxchbondo_out,
    input           rxchbondslave_in,
    output          rxchanisaligned_out,
    output          rxchanrealign_out,
    input           rxdfeagchold_in,
    input           rxdfelfhold_in,
    input           rxdfelpmreset_in,
    output  [6:0]   rxmonitorout_out,
    input   [1:0]   rxmonitorsel_in,
    output          rxoutclk_out,
    input           gtrxreset_in,
    input           rxpcsreset_in,
    input           rxpmareset_in,
    input           rxlpmen_in,
    input           rxpolarity_in,
    output  [3:0]   rxchariscomma_out,
    output  [3:0]   rxcharisk_out,
    input   [4:0]   rxchbondi_in,
    output          rxresetdone_out,
    input   [4:0]   txpostcursor_in,
    input   [4:0]   txprecursor_in,
    input           gttxreset_in,
    input           txuserrdy_in,
    input           txusrclk_in,
    input           txusrclk2_in,
    input           txprbsforceerr_in,
    output  [1:0]   txbufstatus_out,
    input   [3:0]   txdiffctrl_in,
    input           txinhibit_in,
    input   [31:0]  txdata_in,
    output          gtxtxn_out,
    output          gtxtxp_out,
    output          txoutclk_out,
    output          txoutclkfabric_out,
    output          txoutclkpcs_out,
    input   [3:0]   txcharisk_in,
    input           txpcsreset_in,
    input           txpmareset_in,
    output          txresetdone_out,
    input           txpolarity_in,
    input   [2:0]   txprbssel_in
);
    // ground and vcc signals
wire            tied_to_ground_i;
wire    [63:0]  tied_to_ground_vec_i;
wire            tied_to_vcc_i;
wire    [63:0]  tied_to_vcc_vec_i;
    //RX Datapath signals
wire    [63:0]  rxdata_i;
wire    [3:0]   rxchariscomma_float_i;
wire    [3:0]   rxcharisk_float_i;
wire    [3:0]   rxdisperr_float_i;
wire    [3:0]   rxnotintable_float_i;
wire    [3:0]   rxrundisp_float_i;
    //TX Datapath signals
wire    [63:0]  txdata_i;
wire    [3:0]   txkerr_float_i;
wire    [3:0]   txrundisp_float_i;
wire            rxstartofseq_float_i;
(* equivalent_register_removal="no" *) reg [95:0]   cpllpd_wait    =  96'hFFFFFFFFFFFFFFFFFFFFFFFF;
(* equivalent_register_removal="no" *) reg [127:0]  cpllreset_wait = 128'h000000000000000000000000000000FF;
wire    cpllpd_ovrd_i ;
wire    cpllreset_ovrd_i ;
wire    cpll_reset_i;
wire    cpllreset_sync;
wire    cpllpd_sync;
wire    cpll_pd_i;
wire    ack_i;
reg     flag = 1'b0;
reg     flag2 = 1'b0;
reg     ack_flag = 1'b0;
  // Internal Signals
  wire data_sync1;
  wire data_sync2;
  wire data_sync3;
  wire data_sync4;
  wire data_sync5;
  wire data_sync6;
  wire ack_sync1;
  wire ack_sync2;
  wire ack_sync3;
  wire ack_sync4;
  wire ack_sync5;
  wire ack_sync6;
    assign tied_to_ground_i             = 1'b0;
    assign tied_to_ground_vec_i         = 64'h0000000000000000;
    assign tied_to_vcc_i                = 1'b1;
    assign tied_to_vcc_vec_i            = 64'hffffffffffffffff;
    assign  rxdata_out    =   rxdata_i[31:0];
    // The GT transmits little endian data (TXDATA[7:0] transmitted first)
    assign  txdata_i    =   {tied_to_ground_vec_i[31:0],txdata_in};
        GTXE2_CHANNEL #
        (
            //_______________________ Simulation-Only Attributes __________________
            .SIM_RECEIVER_DETECT_PASS   ("TRUE"),
            .SIM_TX_EIDLE_DRIVE_LEVEL   ("X"),
            .SIM_RESET_SPEEDUP          (GT_SIM_GTRESET_SPEEDUP),
            .SIM_CPLLREFCLK_SEL         (3'b001),
            .SIM_VERSION                ("4.0"),
            .ALIGN_COMMA_DOUBLE                     ("FALSE"),
            .ALIGN_COMMA_ENABLE                     (10'b1111111111),
            .ALIGN_COMMA_WORD                       (1),
            .ALIGN_MCOMMA_DET                       ("TRUE"),
            .ALIGN_MCOMMA_VALUE                     (10'b1010000011),
            .ALIGN_PCOMMA_DET                       ("TRUE"),
            .ALIGN_PCOMMA_VALUE                     (10'b0101111100),
            .SHOW_REALIGN_COMMA                     ("TRUE"),
            .RXSLIDE_AUTO_WAIT                      (7),
            .RXSLIDE_MODE                           ("OFF"),
            .RX_SIG_VALID_DLY                       (10),
            .RX_DISPERR_SEQ_MATCH                   ("TRUE"),
            .DEC_MCOMMA_DETECT                      ("TRUE"),
            .DEC_PCOMMA_DETECT                      ("TRUE"),
            .DEC_VALID_COMMA_ONLY                   ("TRUE"),
            .CBCC_DATA_SOURCE_SEL                   ("DECODED"),
            .CLK_COR_SEQ_2_USE                      ("FALSE"),
            .CLK_COR_KEEP_IDLE                      ("FALSE"),
            .CLK_COR_MAX_LAT                        (36),
            .CLK_COR_MIN_LAT                        (31),
            .CLK_COR_PRECEDENCE                     ("TRUE"),
            .CLK_COR_REPEAT_WAIT                    (0),
            .CLK_COR_SEQ_LEN                        (2),
            .CLK_COR_SEQ_1_ENABLE                   (4'b0011),
            .CLK_COR_SEQ_1_1                        (10'b0111111101),
            .CLK_COR_SEQ_1_2                        (10'b0111111101),
            .CLK_COR_SEQ_1_3                        (10'b0000000000),
            .CLK_COR_SEQ_1_4                        (10'b0000000000),
            .CLK_CORRECT_USE                        ("TRUE"),
            .CLK_COR_SEQ_2_ENABLE                   (4'b1111),
            .CLK_COR_SEQ_2_1                        (10'b0000000000),
            .CLK_COR_SEQ_2_2                        (10'b0000000000),
            .CLK_COR_SEQ_2_3                        (10'b0000000000),
            .CLK_COR_SEQ_2_4                        (10'b0000000000),
            .CHAN_BOND_KEEP_ALIGN                   ("FALSE"),
            .CHAN_BOND_MAX_SKEW                     (8),
            .CHAN_BOND_SEQ_LEN                      (1),
            .CHAN_BOND_SEQ_1_1                      (10'b0111111011),
            .CHAN_BOND_SEQ_1_2                      (10'b0000000000),
            .CHAN_BOND_SEQ_1_3                      (10'b0000000000),
            .CHAN_BOND_SEQ_1_4                      (10'b0000000000),
            .CHAN_BOND_SEQ_1_ENABLE                 (4'b0001),
            .CHAN_BOND_SEQ_2_1                      (10'b0000000000),
            .CHAN_BOND_SEQ_2_2                      (10'b0000000000),
            .CHAN_BOND_SEQ_2_3                      (10'b0000000000),
            .CHAN_BOND_SEQ_2_4                      (10'b0000000000),
            .CHAN_BOND_SEQ_2_ENABLE                 (4'b1111),
            .CHAN_BOND_SEQ_2_USE                    ("FALSE"),
            .FTS_DESKEW_SEQ_ENABLE                  (4'b1111),
            .FTS_LANE_DESKEW_CFG                    (4'b1111),
            .FTS_LANE_DESKEW_EN                     ("FALSE"),
            .ES_CONTROL                             (6'b000000),
            .ES_ERRDET_EN                           ("FALSE"),
            .ES_EYE_SCAN_EN                         ("TRUE"),
            .ES_HORZ_OFFSET                         (12'h000),
            .ES_PMA_CFG                             (10'b0000000000),
            .ES_PRESCALE                            (5'b00000),
            .ES_QUALIFIER                           (80'h00000000000000000000),
            .ES_QUAL_MASK                           (80'h00000000000000000000),
            .ES_SDATA_MASK                          (80'h00000000000000000000),
            .ES_VERT_OFFSET                         (9'b000000000),
            .RX_DATA_WIDTH                          (40),
            .OUTREFCLK_SEL_INV                      (2'b11),
            .PMA_RSV                                (PMA_RSV_IN),
            .PMA_RSV2                               (16'h2050),
            .PMA_RSV3                               (2'b00),
            .PMA_RSV4                               (32'h00000000),
            .RX_BIAS_CFG                            (12'b000000000100),
            .DMONITOR_CFG                           (24'h000A00),
            .RX_CM_SEL                              (2'b11),
            .RX_CM_TRIM                             (3'b010),
            .RX_DEBUG_CFG                           (12'b000000000000),
            .RX_OS_CFG                              (13'b0000010000000),
            .TERM_RCAL_CFG                          (5'b10000),
            .TERM_RCAL_OVRD                         (1'b0),
            .TST_RSV                                (32'h00000000),
            .RX_CLK25_DIV                           (7),
            .TX_CLK25_DIV                           (7),
            .UCODEER_CLR                            (1'b0),
            .PCS_PCIE_EN                            ("FALSE"),
            .PCS_RSVD_ATTR                          (PCS_RSVD_ATTR_IN),
            .RXBUF_ADDR_MODE                        ("FULL"),
            .RXBUF_EIDLE_HI_CNT                     (4'b1000),
            .RXBUF_EIDLE_LO_CNT                     (4'b0000),
            .RXBUF_EN                               ("TRUE"),
            .RX_BUFFER_CFG                          (6'b000000),
            .RXBUF_RESET_ON_CB_CHANGE               ("TRUE"),
            .RXBUF_RESET_ON_COMMAALIGN              ("FALSE"),
            .RXBUF_RESET_ON_EIDLE                   ("FALSE"),
            .RXBUF_RESET_ON_RATE_CHANGE             ("TRUE"),
            .RXBUFRESET_TIME                        (5'b00001),
            .RXBUF_THRESH_OVFLW                     (61),
            .RXBUF_THRESH_OVRD                      ("FALSE"),
            .RXBUF_THRESH_UNDFLW                    (4),
            .RXDLY_CFG                              (16'h001F),
            .RXDLY_LCFG                             (9'h030),
            .RXDLY_TAP_CFG                          (16'h0000),
            .RXPH_CFG                               (24'h000000),
            .RXPHDLY_CFG                            (24'h084020),
            .RXPH_MONITOR_SEL                       (5'b00000),
            .RX_XCLK_SEL                            ("RXREC"),
            .RX_DDI_SEL                             (6'b000000),
            .RX_DEFER_RESET_BUF_EN                  ("TRUE"),
           //For Display Port, HBR/RBR- set RXCDR_CFG=72'h0380008bff40200008
           //For Display Port, HBR2 -   set RXCDR_CFG=72'h038c008bff20200010
           //For SATA Gen1- set RXCDR_CFG=72'h03_8000_8BFF_4010_0008
           //For SATA Gen2- set RXCDR_CFG=72'h03_8800_8BFF_4020_0008
           //For SATA Gen3- set RXCDR_CFG=72'h03_8000_8BFF_1020_0010
            .RXCDR_CFG                              (72'h03000023ff40200020),
            .RXCDR_FR_RESET_ON_EIDLE                (1'b0),
            .RXCDR_HOLD_DURING_EIDLE                (1'b0),
            .RXCDR_PH_RESET_ON_EIDLE                (1'b0),
            .RXCDR_LOCK_CFG                         (6'b010101),
            .RXCDRFREQRESET_TIME                    (5'b00001),
            .RXCDRPHRESET_TIME                      (5'b00001),
            .RXISCANRESET_TIME                      (5'b00001),
            .RXPCSRESET_TIME                        (5'b00001),
            .RXPMARESET_TIME                        (5'b00011),
            .RXOOB_CFG                              (7'b0000110),
            .RXGEARBOX_EN                           ("FALSE"),
            .GEARBOX_MODE                           (3'b000),
            .RXPRBS_ERR_LOOPBACK                    (1'b0),
            .PD_TRANS_TIME_FROM_P2                  (12'h03c),
            .PD_TRANS_TIME_NONE_P2                  (8'h19),
            .PD_TRANS_TIME_TO_P2                    (8'h64),
            .SAS_MAX_COM                            (64),
            .SAS_MIN_COM                            (36),
            .SATA_BURST_SEQ_LEN                     (4'b0101),
            .SATA_BURST_VAL                         (3'b100),
            .SATA_EIDLE_VAL                         (3'b100),
            .SATA_MAX_BURST                         (8),
            .SATA_MAX_INIT                          (21),
            .SATA_MAX_WAKE                          (7),
            .SATA_MIN_BURST                         (4),
            .SATA_MIN_INIT                          (12),
            .SATA_MIN_WAKE                          (4),
            .TRANS_TIME_RATE                        (8'h0E),
            .TXBUF_EN                               ("TRUE"),
            .TXBUF_RESET_ON_RATE_CHANGE             ("TRUE"),
            .TXDLY_CFG                              (16'h001F),
            .TXDLY_LCFG                             (9'h030),
            .TXDLY_TAP_CFG                          (16'h0000),
            .TXPH_CFG                               (16'h0780),
            .TXPHDLY_CFG                            (24'h084020),
            .TXPH_MONITOR_SEL                       (5'b00000),
            .TX_XCLK_SEL                            ("TXOUT"),
            .TX_DATA_WIDTH                          (40),
            .TX_DEEMPH0                             (5'b00000),
            .TX_DEEMPH1                             (5'b00000),
            .TX_EIDLE_ASSERT_DELAY                  (3'b110),
            .TX_EIDLE_DEASSERT_DELAY                (3'b100),
            .TX_LOOPBACK_DRIVE_HIZ                  ("FALSE"),
            .TX_MAINCURSOR_SEL                      (1'b0),
            .TX_DRIVE_MODE                          ("DIRECT"),
            .TX_MARGIN_FULL_0                       (7'b1001110),
            .TX_MARGIN_FULL_1                       (7'b1001001),
            .TX_MARGIN_FULL_2                       (7'b1000101),
            .TX_MARGIN_FULL_3                       (7'b1000010),
            .TX_MARGIN_FULL_4                       (7'b1000000),
            .TX_MARGIN_LOW_0                        (7'b1000110),
            .TX_MARGIN_LOW_1                        (7'b1000100),
            .TX_MARGIN_LOW_2                        (7'b1000010),
            .TX_MARGIN_LOW_3                        (7'b1000000),
            .TX_MARGIN_LOW_4                        (7'b1000000),
            .TXGEARBOX_EN                           ("FALSE"),
            .TXPCSRESET_TIME                        (5'b00001),
            .TXPMARESET_TIME                        (5'b00001),
            .TX_RXDETECT_CFG                        (14'h1832),
            .TX_RXDETECT_REF                        (3'b100),
            .CPLL_CFG                               (24'hBC07DC),
            .CPLL_FBDIV                             (4),
            .CPLL_FBDIV_45                          (5),
            .CPLL_INIT_CFG                          (24'h00001E),
            .CPLL_LOCK_CFG                          (16'h01E8),
            .CPLL_REFCLK_DIV                        (1),
            .RXOUT_DIV                              (2),
            .TXOUT_DIV                              (2),
            .SATA_CPLL_CFG                          ("VCO_3000MHZ"),
            .RXDFELPMRESET_TIME                     (7'b0001111),
            .RXLPM_HF_CFG                           (14'b00000011110000),
            .RXLPM_LF_CFG                           (14'b00000011110000),
            .RX_DFE_GAIN_CFG                        (23'h020FEA),
            .RX_DFE_H2_CFG                          (12'b000000000000),
            .RX_DFE_H3_CFG                          (12'b000001000000),
            .RX_DFE_H4_CFG                          (11'b00011110000),
            .RX_DFE_H5_CFG                          (11'b00011100000),
            .RX_DFE_KL_CFG                          (13'b0000011111110),
            .RX_DFE_LPM_CFG                         (16'h0954),
            .RX_DFE_LPM_HOLD_DURING_EIDLE           (1'b0),
            .RX_DFE_UT_CFG                          (17'b10001111000000000),
            .RX_DFE_VP_CFG                          (17'b00011111100000011),
            .RX_CLKMUX_PD                           (1'b1),
            .TX_CLKMUX_PD                           (1'b1),
            .RX_INT_DATAWIDTH                       (0),
            .TX_INT_DATAWIDTH                       (0),
            .TX_QPI_STATUS_EN                       (1'b0),
            .RX_DFE_KL_CFG2                         (RX_DFE_KL_CFG2_IN),
            .RX_DFE_XYD_CFG                         (13'b0000000000000),
            .TX_PREDRIVER_MODE                      (1'b0)
        )
        gtxe2_i
        (
        .CPLLFBCLKLOST                  (cpllfbclklost_out),
        .CPLLLOCK                       (cplllock_out),
        .CPLLLOCKDETCLK                 (cplllockdetclk_in),
        .CPLLLOCKEN                     (tied_to_vcc_i),
        .CPLLPD                         (cpll_pd_i),
        .CPLLREFCLKLOST                 (cpllrefclklost_out),
        .CPLLREFCLKSEL                  (3'b001),
        .CPLLRESET                      (cpll_reset_i),
        .GTRSVD                         (16'b0000000000000000),
        .PCSRSVDIN                      (16'b0000000000000000),
        .PCSRSVDIN2                     (5'b00000),
        .PMARSVDIN                      (5'b00000),
        .PMARSVDIN2                     (5'b00000),
        .TSTIN                          (20'b11111111111111111111),
        .TSTOUT                         (),
        .CLKRSVD                        (4'b0000),
        .GTGREFCLK                      (tied_to_ground_i),
        .GTNORTHREFCLK0                 (tied_to_ground_i),
        .GTNORTHREFCLK1                 (tied_to_ground_i),
        .GTREFCLK0                      (gtrefclk0_in),
        .GTREFCLK1                      (tied_to_ground_i),
        .GTSOUTHREFCLK0                 (tied_to_ground_i),
        .GTSOUTHREFCLK1                 (tied_to_ground_i),
        .DRPADDR                        (drpaddr_in),
        .DRPCLK                         (drpclk_in),
        .DRPDI                          (drpdi_in),
        .DRPDO                          (drpdo_out),
        .DRPEN                          (drpen_in),
        .DRPRDY                         (drprdy_out),
        .DRPWE                          (drpwe_in),
        .GTREFCLKMONITOR                (),
        .QPLLCLK                        (qpllclk_in),
        .QPLLREFCLK                     (qpllrefclk_in),
        .RXSYSCLKSEL                    (2'b00),
        .TXSYSCLKSEL                    (2'b00),
        .DMONITOROUT                    (dmonitorout_out),
        .TX8B10BEN                      (tied_to_vcc_i),
        .LOOPBACK                       (loopback_in),
        .PHYSTATUS                      (),
        .RXRATE                         (tied_to_ground_vec_i[2:0]),
        .RXVALID                        (),
        .RXPD                           (2'b00),
        .TXPD                           (2'b00),
        .SETERRSTATUS                   (tied_to_ground_i),
        .EYESCANRESET                   (eyescanreset_in),
        .RXUSERRDY                      (rxuserrdy_in),
        .EYESCANDATAERROR               (eyescandataerror_out),
        .EYESCANMODE                    (tied_to_ground_i),
        .EYESCANTRIGGER                 (eyescantrigger_in),
        .RXCDRFREQRESET                 (tied_to_ground_i),
        .RXCDRHOLD                      (rxcdrhold_in),
        .RXCDRLOCK                      (),
        .RXCDROVRDEN                    (tied_to_ground_i),
        .RXCDRRESET                     (tied_to_ground_i),
        .RXCDRRESETRSV                  (tied_to_ground_i),
        .RXCLKCORCNT                    (rxclkcorcnt_out),
        .RX8B10BEN                      (tied_to_vcc_i),
        .RXUSRCLK                       (rxusrclk_in),
        .RXUSRCLK2                      (rxusrclk2_in),
        .RXDATA                         (rxdata_i),
        .RXPRBSERR                      (rxprbserr_out),
        .RXPRBSSEL                      (rxprbssel_in),
        .RXPRBSCNTRESET                 (rxprbscntreset_in),
        .RXDFEXYDEN                     (tied_to_vcc_i),
        .RXDFEXYDHOLD                   (tied_to_ground_i),
        .RXDFEXYDOVRDEN                 (tied_to_ground_i),
        .RXDISPERR                      ({rxdisperr_float_i,rxdisperr_out}),
        .RXNOTINTABLE                   ({rxnotintable_float_i,rxnotintable_out}),
        .GTXRXP                         (gtxrxp_in),
        .GTXRXN                         (gtxrxn_in),
        .RXBUFRESET                     (rxbufreset_in),
        .RXBUFSTATUS                    (rxbufstatus_out),
        .RXDDIEN                        (tied_to_ground_i),
        .RXDLYBYPASS                    (tied_to_vcc_i),
        .RXDLYEN                        (tied_to_ground_i),
        .RXDLYOVRDEN                    (tied_to_ground_i),
        .RXDLYSRESET                    (tied_to_ground_i),
        .RXDLYSRESETDONE                (),
        .RXPHALIGN                      (tied_to_ground_i),
        .RXPHALIGNDONE                  (),
        .RXPHALIGNEN                    (tied_to_ground_i),
        .RXPHDLYPD                      (tied_to_ground_i),
        .RXPHDLYRESET                   (tied_to_ground_i),
        .RXPHMONITOR                    (),
        .RXPHOVRDEN                     (tied_to_ground_i),
        .RXPHSLIPMONITOR                (),
        .RXSTATUS                       (),
        .RXBYTEISALIGNED                (rxbyteisaligned_out),
        .RXBYTEREALIGN                  (rxbyterealign_out),
        .RXCOMMADET                     (rxcommadet_out),
        .RXCOMMADETEN                   (tied_to_vcc_i),
        .RXMCOMMAALIGNEN                (rxmcommaalignen_in),
        .RXPCOMMAALIGNEN                (rxpcommaalignen_in),
        .RXCHANBONDSEQ                  (rxchanbondseq_out),
        .RXCHBONDEN                     (rxchbonden_in),
        .RXCHBONDLEVEL                  (rxchbondlevel_in),
        .RXCHBONDMASTER                 (rxchbondmaster_in),
        .RXCHBONDO                      (rxchbondo_out),
        .RXCHBONDSLAVE                  (rxchbondslave_in),
        .RXCHANISALIGNED                (rxchanisaligned_out),
        .RXCHANREALIGN                  (rxchanrealign_out),
        .RXLPMHFHOLD                    (tied_to_ground_i),
        .RXLPMHFOVRDEN                  (tied_to_ground_i),
        .RXLPMLFHOLD                    (tied_to_ground_i),
        .RXDFEAGCHOLD                   (rxdfeagchold_in),
        .RXDFEAGCOVRDEN                 (tied_to_ground_i),
        .RXDFECM1EN                     (tied_to_ground_i),
        .RXDFELFHOLD                    (rxdfelfhold_in),
        .RXDFELFOVRDEN                  (tied_to_vcc_i),
        .RXDFELPMRESET                  (rxdfelpmreset_in),
        .RXDFETAP2HOLD                  (tied_to_ground_i),
        .RXDFETAP2OVRDEN                (tied_to_ground_i),
        .RXDFETAP3HOLD                  (tied_to_ground_i),
        .RXDFETAP3OVRDEN                (tied_to_ground_i),
        .RXDFETAP4HOLD                  (tied_to_ground_i),
        .RXDFETAP4OVRDEN                (tied_to_ground_i),
        .RXDFETAP5HOLD                  (tied_to_ground_i),
        .RXDFETAP5OVRDEN                (tied_to_ground_i),
        .RXDFEUTHOLD                    (tied_to_ground_i),
        .RXDFEUTOVRDEN                  (tied_to_ground_i),
        .RXDFEVPHOLD                    (tied_to_ground_i),
        .RXDFEVPOVRDEN                  (tied_to_ground_i),
        .RXDFEVSEN                      (tied_to_ground_i),
        .RXLPMLFKLOVRDEN                (tied_to_ground_i),
        .RXMONITOROUT                   (rxmonitorout_out),
        .RXMONITORSEL                   (rxmonitorsel_in),
        .RXOSHOLD                       (tied_to_ground_i),
        .RXOSOVRDEN                     (tied_to_ground_i),
        .RXRATEDONE                     (),
        .RXOUTCLK                       (rxoutclk_out),
        .RXOUTCLKFABRIC                 (),
        .RXOUTCLKPCS                    (),
        .RXOUTCLKSEL                    (3'b010),
        .RXDATAVALID                    (),
        .RXHEADER                       (),
        .RXHEADERVALID                  (),
        .RXSTARTOFSEQ                   (),
        .RXGEARBOXSLIP                  (tied_to_ground_i),
        .GTRXRESET                      (gtrxreset_in),
        .RXOOBRESET                     (tied_to_ground_i),
        .RXPCSRESET                     (rxpcsreset_in),
        .RXPMARESET                     (rxpmareset_in),
        .RXLPMEN                        (rxlpmen_in),
        .RXCOMSASDET                    (),
        .RXCOMWAKEDET                   (),
        .RXCOMINITDET                   (),
        .RXELECIDLE                     (),
        .RXELECIDLEMODE                 (2'b11),
        .RXPOLARITY                     (rxpolarity_in),
        .RXSLIDE                        (tied_to_ground_i),
        .RXCHARISCOMMA                  ({rxchariscomma_float_i,rxchariscomma_out}),
        .RXCHARISK                      ({rxcharisk_float_i,rxcharisk_out}),
        .RXCHBONDI                      (rxchbondi_in),
        .RXRESETDONE                    (rxresetdone_out),
        .RXQPIEN                        (tied_to_ground_i),
        .RXQPISENN                      (),
        .RXQPISENP                      (),
        .TXPHDLYTSTCLK                  (tied_to_ground_i),
        .TXPOSTCURSOR                   (txpostcursor_in),
        .TXPOSTCURSORINV                (tied_to_ground_i),
        .TXPRECURSOR                    (txprecursor_in),
        .TXPRECURSORINV                 (tied_to_ground_i),
        .TXQPIBIASEN                    (tied_to_ground_i),
        .TXQPISTRONGPDOWN               (tied_to_ground_i),
        .TXQPIWEAKPUP                   (tied_to_ground_i),
        .CFGRESET                       (tied_to_ground_i),
        .GTTXRESET                      (gttxreset_in),
        .PCSRSVDOUT                     (),
        .TXUSERRDY                      (txuserrdy_in),
        .GTRESETSEL                     (tied_to_ground_i),
        .RESETOVRD                      (tied_to_ground_i),
        .TXCHARDISPMODE                 (tied_to_ground_vec_i[7:0]),
        .TXCHARDISPVAL                  (tied_to_ground_vec_i[7:0]),
        .TXUSRCLK                       (txusrclk_in),
        .TXUSRCLK2                      (txusrclk2_in),
        .TXELECIDLE                     (tied_to_ground_i),
        .TXMARGIN                       (tied_to_ground_vec_i[2:0]),
        .TXRATE                         (tied_to_ground_vec_i[2:0]),
        .TXSWING                        (tied_to_ground_i),
        .TXPRBSFORCEERR                 (txprbsforceerr_in),
        .TXDLYBYPASS                    (tied_to_vcc_i),
        .TXDLYEN                        (tied_to_ground_i),
        .TXDLYHOLD                      (tied_to_ground_i),
        .TXDLYOVRDEN                    (tied_to_ground_i),
        .TXDLYSRESET                    (tied_to_ground_i),
        .TXDLYSRESETDONE                (),
        .TXDLYUPDOWN                    (tied_to_ground_i),
        .TXPHALIGN                      (tied_to_ground_i),
        .TXPHALIGNDONE                  (),
        .TXPHALIGNEN                    (tied_to_ground_i),
        .TXPHDLYPD                      (tied_to_ground_i),
        .TXPHDLYRESET                   (tied_to_ground_i),
        .TXPHINIT                       (tied_to_ground_i),
        .TXPHINITDONE                   (),
        .TXPHOVRDEN                     (tied_to_ground_i),
        .TXBUFSTATUS                    (txbufstatus_out),
        .TXBUFDIFFCTRL                  (3'b100),
        .TXDEEMPH                       (tied_to_ground_i),
        .TXDIFFCTRL                     (txdiffctrl_in),
        .TXDIFFPD                       (tied_to_ground_i),
        .TXINHIBIT                      (txinhibit_in),
        .TXMAINCURSOR                   (7'b0000000),
        .TXPISOPD                       (tied_to_ground_i),
        .TXDATA                         (txdata_i),
        .GTXTXN                         (gtxtxn_out),
        .GTXTXP                         (gtxtxp_out),
        .TXOUTCLK                       (txoutclk_out),
        .TXOUTCLKFABRIC                 (txoutclkfabric_out),
        .TXOUTCLKPCS                    (txoutclkpcs_out),
        .TXOUTCLKSEL                    (3'b010),
        .TXRATEDONE                     (),
        .TXCHARISK                      ({tied_to_ground_vec_i[3:0],txcharisk_in}),
        .TXGEARBOXREADY                 (),
        .TXHEADER                       (tied_to_ground_vec_i[2:0]),
        .TXSEQUENCE                     (tied_to_ground_vec_i[6:0]),
        .TXSTARTSEQ                     (tied_to_ground_i),
        .TXPCSRESET                     (txpcsreset_in),
        .TXPMARESET                     (txpmareset_in),
        .TXRESETDONE                    (txresetdone_out),
        .TXCOMFINISH                    (),
        .TXCOMINIT                      (tied_to_ground_i),
        .TXCOMSAS                       (tied_to_ground_i),
        .TXCOMWAKE                      (tied_to_ground_i),
        .TXPDELECIDLEMODE               (tied_to_ground_i),
        .TXPOLARITY                     (txpolarity_in),
        .TXDETECTRX                     (tied_to_ground_i),
        .TX8B10BBYPASS                  (tied_to_ground_vec_i[7:0]),
        .TXPRBSSEL                      (txprbssel_in),
        .TXQPISENN                      (),
        .TXQPISENP                      ()
     );
always @(posedge gtrefclk0_in)
begin
  cpllpd_wait <= {cpllpd_wait[94:0], 1'b0};
  cpllreset_wait <= {cpllreset_wait[126:0], 1'b0};
end
assign cpllpd_ovrd_i = cpllpd_wait[95];
assign cpllreset_ovrd_i = cpllreset_wait[127];
assign cpll_pd_i = cpllpd_ovrd_i;
always @(posedge drpclk_in)
begin
if(cpllreset_in == 1'b1 && ack_flag == 1'b0)
begin
    flag <= !flag;
    flag2 <= 1'b1;
end
else
begin
    flag <= flag;
    flag2 <= 1'b0;
end
end
always @(posedge drpclk_in)
begin
if(flag2 == 1'b1)
 ack_flag <= 1'b1;
else if(ack_i == 1'b1)
 ack_flag <= 1'b0;
end
  (* shreg_extract = "no", ASYNC_REG = "TRUE" *)
  FD #(
    .INIT (1'b0)
  ) data_sync_reg1 (
    .C  (gtrefclk0_in),
    .D  (flag),
    .Q  (data_sync1)
  );
  (* shreg_extract = "no", ASYNC_REG = "TRUE" *)
  FD #(
   .INIT (1'b0)
  ) data_sync_reg2 (
  .C  (gtrefclk0_in),
  .D  (data_sync1),
  .Q  (data_sync2)
  );
  (* shreg_extract = "no", ASYNC_REG = "TRUE" *)
  FD #(
   .INIT (1'b0)
  ) data_sync_reg3 (
  .C  (gtrefclk0_in),
  .D  (data_sync2),
  .Q  (data_sync3)
  );
  (* shreg_extract = "no", ASYNC_REG = "TRUE" *)
  FD #(
   .INIT (1'b0)
  ) data_sync_reg4 (
  .C  (gtrefclk0_in),
  .D  (data_sync3),
  .Q  (data_sync4)
  );
  (* shreg_extract = "no", ASYNC_REG = "TRUE" *)
  FD #(
   .INIT (1'b0)
  ) data_sync_reg5 (
  .C  (gtrefclk0_in),
  .D  (data_sync4),
  .Q  (data_sync5)
  );
  (* shreg_extract = "no", ASYNC_REG = "TRUE" *)
  FD #(
   .INIT (1'b0)
  ) data_sync_reg6 (
  .C  (gtrefclk0_in),
  .D  (data_sync5),
  .Q  (data_sync6)
  );
assign cpllreset_sync = data_sync5 ^ data_sync6;
  (* shreg_extract = "no", ASYNC_REG = "TRUE" *)
  FD #(
   .INIT (1'b0)
  ) ack_sync_reg1 (
  .C  (drpclk_in),
  .D  (data_sync6),
  .Q  (ack_sync1)
  );
  (* shreg_extract = "no", ASYNC_REG = "TRUE" *)
  FD #(
   .INIT (1'b0)
  ) ack_sync_reg2 (
  .C  (drpclk_in),
  .D  (ack_sync1),
  .Q  (ack_sync2)
  );
  (* shreg_extract = "no", ASYNC_REG = "TRUE" *)
  FD #(
   .INIT (1'b0)
  ) ack_sync_reg3 (
  .C  (drpclk_in),
  .D  (ack_sync2),
  .Q  (ack_sync3)
  );
  (* shreg_extract = "no", ASYNC_REG = "TRUE" *)
  FD #(
   .INIT (1'b0)
  ) ack_sync_reg4 (
  .C  (drpclk_in),
  .D  (ack_sync3),
  .Q  (ack_sync4)
  );
  (* shreg_extract = "no", ASYNC_REG = "TRUE" *)
  FD #(
   .INIT (1'b0)
  ) ack_sync_reg5 (
  .C  (drpclk_in),
  .D  (ack_sync4),
  .Q  (ack_sync5)
  );
  (* shreg_extract = "no", ASYNC_REG = "TRUE" *)
  FD #(
   .INIT (1'b0)
  ) ack_sync_reg6 (
  .C  (drpclk_in),
  .D  (ack_sync5),
  .Q  (ack_sync6)
  );
assign ack_i = ack_sync5 ^ ack_sync6;
assign cpll_reset_i = cpllreset_sync || cpllreset_ovrd_i;
endmodule