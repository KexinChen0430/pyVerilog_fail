module topkeyboard(PS2_CLK, PS2_DAT, LEDR);
  synthkeyboard(clock
endmodule