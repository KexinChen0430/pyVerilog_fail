module top ;
          wire  Net_163;
          wire  Net_162;
          wire  Net_161;
          wire  Net_154;
          wire  Net_139;
          wire  Net_153;
          wire  Net_137;
          wire  Net_152;
          wire  Net_151;
          wire  Net_150;
          wire  Net_149;
          wire  Net_148;
          wire  Net_147;
          wire  Net_146;
          wire  Net_145;
          wire  Net_144;
          wire  Net_69;
          wire  Net_102;
          wire  Net_101;
          wire  Net_100;
          wire  Net_99;
          wire  Net_98;
          wire  Net_87;
          wire  Net_97;
          wire  Net_96;
          wire  Net_95;
          wire  Net_94;
          wire  Net_93;
          wire  Net_104;
          wire  Net_68;
          wire  Net_46;
	wire [0:0] tmpOE__Btn0_net;
	wire [0:0] tmpFB_0__Btn0_net;
	wire [0:0] tmpIO_0__Btn0_net;
	electrical [0:0] tmpSIOVREF__Btn0_net;
	cy_psoc3_pins_v1_10
		#(.id("552faf00-97dc-47bf-ad14-15574b2c6e9b"),
		  .drive_mode(3'b010),
		  .ibuf_enabled(1'b1),
		  .init_dr_st(1'b1),
		  .input_clk_en(0),
		  .input_sync(1'b1),
		  .input_sync_mode(1'b0),
		  .intr_mode(2'b10),
		  .invert_in_clock(0),
		  .invert_in_clock_en(0),
		  .invert_in_reset(0),
		  .invert_out_clock(0),
		  .invert_out_clock_en(0),
		  .invert_out_reset(0),
		  .io_voltage(""),
		  .layout_mode("CONTIGUOUS"),
		  .oe_conn(1'b0),
		  .oe_reset(0),
		  .oe_sync(1'b0),
		  .output_clk_en(0),
		  .output_clock_mode(1'b0),
		  .output_conn(1'b0),
		  .output_mode(1'b0),
		  .output_reset(0),
		  .output_sync(1'b0),
		  .pa_in_clock(-1),
		  .pa_in_clock_en(-1),
		  .pa_in_reset(-1),
		  .pa_out_clock(-1),
		  .pa_out_clock_en(-1),
		  .pa_out_reset(-1),
		  .pin_aliases(""),
		  .pin_mode("I"),
		  .por_state(4),
		  .sio_group_cnt(0),
		  .sio_hyst(1'b0),
		  .sio_ibuf(""),
		  .sio_info(2'b00),
		  .sio_obuf(""),
		  .sio_refsel(""),
		  .sio_vtrip(""),
		  .slew_rate(1'b0),
		  .spanning(0),
		  .use_annotation(1'b0),
		  .vtrip(2'b00),
		  .width(1))
		Btn0
		 (.oe(tmpOE__Btn0_net),
		  .y({1'b0}),
		  .fb({tmpFB_0__Btn0_net[0:0]}),
		  .io({tmpIO_0__Btn0_net[0:0]}),
		  .siovref(tmpSIOVREF__Btn0_net),
		  .interrupt({Net_46}),
		  .in_clock({1'b0}),
		  .in_clock_en({1'b1}),
		  .in_reset({1'b0}),
		  .out_clock({1'b0}),
		  .out_clock_en({1'b1}),
		  .out_reset({1'b0}));
	assign tmpOE__Btn0_net = (`CYDEV_CHIP_MEMBER_USED == `CYDEV_CHIP_MEMBER_3A && `CYDEV_CHIP_REVISION_USED < `CYDEV_CHIP_REVISION_3A_ES3) ? ~{1'b1} : {1'b1};
	wire [0:0] tmpOE__LED_net;
	wire [0:0] tmpFB_0__LED_net;
	wire [0:0] tmpIO_0__LED_net;
	wire [0:0] tmpINTERRUPT_0__LED_net;
	electrical [0:0] tmpSIOVREF__LED_net;
	cy_psoc3_pins_v1_10
		#(.id("b0f37199-6c06-4e0a-98e7-b2170ef91497"),
		  .drive_mode(3'b110),
		  .ibuf_enabled(1'b1),
		  .init_dr_st(1'b0),
		  .input_clk_en(0),
		  .input_sync(1'b1),
		  .input_sync_mode(1'b0),
		  .intr_mode(2'b00),
		  .invert_in_clock(0),
		  .invert_in_clock_en(0),
		  .invert_in_reset(0),
		  .invert_out_clock(0),
		  .invert_out_clock_en(0),
		  .invert_out_reset(0),
		  .io_voltage(""),
		  .layout_mode("CONTIGUOUS"),
		  .oe_conn(1'b0),
		  .oe_reset(0),
		  .oe_sync(1'b0),
		  .output_clk_en(0),
		  .output_clock_mode(1'b0),
		  .output_conn(1'b0),
		  .output_mode(1'b0),
		  .output_reset(0),
		  .output_sync(1'b0),
		  .pa_in_clock(-1),
		  .pa_in_clock_en(-1),
		  .pa_in_reset(-1),
		  .pa_out_clock(-1),
		  .pa_out_clock_en(-1),
		  .pa_out_reset(-1),
		  .pin_aliases(""),
		  .pin_mode("O"),
		  .por_state(4),
		  .sio_group_cnt(0),
		  .sio_hyst(1'b0),
		  .sio_ibuf(""),
		  .sio_info(2'b00),
		  .sio_obuf(""),
		  .sio_refsel(""),
		  .sio_vtrip(""),
		  .slew_rate(1'b0),
		  .spanning(0),
		  .use_annotation(1'b0),
		  .vtrip(2'b10),
		  .width(1))
		LED
		 (.oe(tmpOE__LED_net),
		  .y({1'b0}),
		  .fb({tmpFB_0__LED_net[0:0]}),
		  .io({tmpIO_0__LED_net[0:0]}),
		  .siovref(tmpSIOVREF__LED_net),
		  .interrupt({tmpINTERRUPT_0__LED_net[0:0]}),
		  .in_clock({1'b0}),
		  .in_clock_en({1'b1}),
		  .in_reset({1'b0}),
		  .out_clock({1'b0}),
		  .out_clock_en({1'b1}),
		  .out_reset({1'b0}));
	assign tmpOE__LED_net = (`CYDEV_CHIP_MEMBER_USED == `CYDEV_CHIP_MEMBER_3A && `CYDEV_CHIP_REVISION_USED < `CYDEV_CHIP_REVISION_3A_ES3) ? ~{1'b1} : {1'b1};
	wire [0:0] tmpOE__Btn1_net;
	wire [0:0] tmpFB_0__Btn1_net;
	wire [0:0] tmpIO_0__Btn1_net;
	electrical [0:0] tmpSIOVREF__Btn1_net;
	cy_psoc3_pins_v1_10
		#(.id("bab6a988-52aa-4376-a76e-7dbb3ddd8f50"),
		  .drive_mode(3'b010),
		  .ibuf_enabled(1'b1),
		  .init_dr_st(1'b1),
		  .input_clk_en(0),
		  .input_sync(1'b1),
		  .input_sync_mode(1'b0),
		  .intr_mode(2'b10),
		  .invert_in_clock(0),
		  .invert_in_clock_en(0),
		  .invert_in_reset(0),
		  .invert_out_clock(0),
		  .invert_out_clock_en(0),
		  .invert_out_reset(0),
		  .io_voltage(""),
		  .layout_mode("CONTIGUOUS"),
		  .oe_conn(1'b0),
		  .oe_reset(0),
		  .oe_sync(1'b0),
		  .output_clk_en(0),
		  .output_clock_mode(1'b0),
		  .output_conn(1'b0),
		  .output_mode(1'b0),
		  .output_reset(0),
		  .output_sync(1'b0),
		  .pa_in_clock(-1),
		  .pa_in_clock_en(-1),
		  .pa_in_reset(-1),
		  .pa_out_clock(-1),
		  .pa_out_clock_en(-1),
		  .pa_out_reset(-1),
		  .pin_aliases(""),
		  .pin_mode("I"),
		  .por_state(4),
		  .sio_group_cnt(0),
		  .sio_hyst(1'b0),
		  .sio_ibuf(""),
		  .sio_info(2'b00),
		  .sio_obuf(""),
		  .sio_refsel(""),
		  .sio_vtrip(""),
		  .slew_rate(1'b0),
		  .spanning(0),
		  .use_annotation(1'b0),
		  .vtrip(2'b00),
		  .width(1))
		Btn1
		 (.oe(tmpOE__Btn1_net),
		  .y({1'b0}),
		  .fb({tmpFB_0__Btn1_net[0:0]}),
		  .io({tmpIO_0__Btn1_net[0:0]}),
		  .siovref(tmpSIOVREF__Btn1_net),
		  .interrupt({Net_104}),
		  .in_clock({1'b0}),
		  .in_clock_en({1'b1}),
		  .in_reset({1'b0}),
		  .out_clock({1'b0}),
		  .out_clock_en({1'b1}),
		  .out_reset({1'b0}));
	assign tmpOE__Btn1_net = (`CYDEV_CHIP_MEMBER_USED == `CYDEV_CHIP_MEMBER_3A && `CYDEV_CHIP_REVISION_USED < `CYDEV_CHIP_REVISION_3A_ES3) ? ~{1'b1} : {1'b1};
    TCPWM_P4_v1_10_0 Timer1 (
        .stop(1'b0),
        .reload(1'b0),
        .start(1'b0),
        .count(1'b1),
        .capture(1'b0),
        .interrupt(Net_87),
        .ov(Net_98),
        .un(Net_99),
        .cc(Net_100),
        .line(Net_101),
        .line_n(Net_102),
        .clock(Net_68));
    defparam Timer1.PWMCountMode = 3;
    defparam Timer1.PWMReloadMode = 0;
    defparam Timer1.PWMReloadPresent = 0;
    defparam Timer1.PWMStartMode = 0;
    defparam Timer1.PWMStopMode = 0;
    defparam Timer1.PWMSwitchMode = 0;
    defparam Timer1.QuadIndexMode = 0;
    defparam Timer1.QuadPhiAMode = 3;
    defparam Timer1.QuadPhiBMode = 3;
    defparam Timer1.QuadStopMode = 0;
    defparam Timer1.TCCaptureMode = 0;
    defparam Timer1.TCCountMode = 3;
    defparam Timer1.TCReloadMode = 0;
    defparam Timer1.TCStartMode = 0;
    defparam Timer1.TCStopMode = 0;
	cy_clock_v1_0
		#(.id("c4d993e1-c103-4e85-b1df-bc9c6402cfed"),
		  .source_clock_id(""),
		  .divisor(0),
		  .period("1000000000"),
		  .is_direct(0),
		  .is_digital(0))
		Clock_1
		 (.clock_out(Net_68));
	cy_isr_v1_0
		#(.int_type(2'b10))
		ISR_Btn0
		 (.int_signal(Net_46));
	cy_isr_v1_0
		#(.int_type(2'b10))
		ISR_Timer1
		 (.int_signal(Net_87));
	wire [0:0] tmpOE__LED1_net;
	wire [0:0] tmpFB_0__LED1_net;
	wire [0:0] tmpIO_0__LED1_net;
	wire [0:0] tmpINTERRUPT_0__LED1_net;
	electrical [0:0] tmpSIOVREF__LED1_net;
	cy_psoc3_pins_v1_10
		#(.id("0e0c9380-6965-4440-8709-ce08a91e474c"),
		  .drive_mode(3'b110),
		  .ibuf_enabled(1'b1),
		  .init_dr_st(1'b0),
		  .input_clk_en(0),
		  .input_sync(1'b1),
		  .input_sync_mode(1'b0),
		  .intr_mode(2'b00),
		  .invert_in_clock(0),
		  .invert_in_clock_en(0),
		  .invert_in_reset(0),
		  .invert_out_clock(0),
		  .invert_out_clock_en(0),
		  .invert_out_reset(0),
		  .io_voltage(""),
		  .layout_mode("CONTIGUOUS"),
		  .oe_conn(1'b0),
		  .oe_reset(0),
		  .oe_sync(1'b0),
		  .output_clk_en(0),
		  .output_clock_mode(1'b0),
		  .output_conn(1'b0),
		  .output_mode(1'b0),
		  .output_reset(0),
		  .output_sync(1'b0),
		  .pa_in_clock(-1),
		  .pa_in_clock_en(-1),
		  .pa_in_reset(-1),
		  .pa_out_clock(-1),
		  .pa_out_clock_en(-1),
		  .pa_out_reset(-1),
		  .pin_aliases(""),
		  .pin_mode("O"),
		  .por_state(4),
		  .sio_group_cnt(0),
		  .sio_hyst(1'b0),
		  .sio_ibuf(""),
		  .sio_info(2'b00),
		  .sio_obuf(""),
		  .sio_refsel(""),
		  .sio_vtrip(""),
		  .slew_rate(1'b0),
		  .spanning(0),
		  .use_annotation(1'b0),
		  .vtrip(2'b10),
		  .width(1))
		LED1
		 (.oe(tmpOE__LED1_net),
		  .y({1'b0}),
		  .fb({tmpFB_0__LED1_net[0:0]}),
		  .io({tmpIO_0__LED1_net[0:0]}),
		  .siovref(tmpSIOVREF__LED1_net),
		  .interrupt({tmpINTERRUPT_0__LED1_net[0:0]}),
		  .in_clock({1'b0}),
		  .in_clock_en({1'b1}),
		  .in_reset({1'b0}),
		  .out_clock({1'b0}),
		  .out_clock_en({1'b1}),
		  .out_reset({1'b0}));
	assign tmpOE__LED1_net = (`CYDEV_CHIP_MEMBER_USED == `CYDEV_CHIP_MEMBER_3A && `CYDEV_CHIP_REVISION_USED < `CYDEV_CHIP_REVISION_3A_ES3) ? ~{1'b1} : {1'b1};
	cy_isr_v1_0
		#(.int_type(2'b10))
		ISR_Bnt1
		 (.int_signal(Net_104));
    TCPWM_P4_v1_10_1 PWM_Servo (
        .stop(1'b0),
        .reload(1'b0),
        .start(1'b0),
        .count(1'b1),
        .capture(1'b0),
        .interrupt(Net_149),
        .ov(Net_150),
        .un(Net_151),
        .cc(Net_152),
        .line(Net_137),
        .line_n(Net_153),
        .clock(Net_139));
    defparam PWM_Servo.PWMCountMode = 3;
    defparam PWM_Servo.PWMReloadMode = 0;
    defparam PWM_Servo.PWMReloadPresent = 0;
    defparam PWM_Servo.PWMStartMode = 0;
    defparam PWM_Servo.PWMStopMode = 0;
    defparam PWM_Servo.PWMSwitchMode = 0;
    defparam PWM_Servo.QuadIndexMode = 0;
    defparam PWM_Servo.QuadPhiAMode = 3;
    defparam PWM_Servo.QuadPhiBMode = 3;
    defparam PWM_Servo.QuadStopMode = 0;
    defparam PWM_Servo.TCCaptureMode = 0;
    defparam PWM_Servo.TCCountMode = 3;
    defparam PWM_Servo.TCReloadMode = 0;
    defparam PWM_Servo.TCStartMode = 0;
    defparam PWM_Servo.TCStopMode = 0;
	cy_clock_v1_0
		#(.id("2f98ca16-0407-4eeb-a907-2282a5b81a79"),
		  .source_clock_id(""),
		  .divisor(0),
		  .period("1000000000"),
		  .is_direct(0),
		  .is_digital(0))
		Clock_2
		 (.clock_out(Net_139));
	wire [0:0] tmpOE__Servo_1_net;
	wire [0:0] tmpFB_0__Servo_1_net;
	wire [0:0] tmpIO_0__Servo_1_net;
	wire [0:0] tmpINTERRUPT_0__Servo_1_net;
	electrical [0:0] tmpSIOVREF__Servo_1_net;
	cy_psoc3_pins_v1_10
		#(.id("e4e9a0b1-0370-4889-90ef-76026e833f55"),
		  .drive_mode(3'b110),
		  .ibuf_enabled(1'b1),
		  .init_dr_st(1'b1),
		  .input_clk_en(0),
		  .input_sync(1'b1),
		  .input_sync_mode(1'b0),
		  .intr_mode(2'b00),
		  .invert_in_clock(0),
		  .invert_in_clock_en(0),
		  .invert_in_reset(0),
		  .invert_out_clock(0),
		  .invert_out_clock_en(0),
		  .invert_out_reset(0),
		  .io_voltage(""),
		  .layout_mode("CONTIGUOUS"),
		  .oe_conn(1'b0),
		  .oe_reset(0),
		  .oe_sync(1'b0),
		  .output_clk_en(0),
		  .output_clock_mode(1'b0),
		  .output_conn(1'b1),
		  .output_mode(1'b0),
		  .output_reset(0),
		  .output_sync(1'b0),
		  .pa_in_clock(-1),
		  .pa_in_clock_en(-1),
		  .pa_in_reset(-1),
		  .pa_out_clock(-1),
		  .pa_out_clock_en(-1),
		  .pa_out_reset(-1),
		  .pin_aliases(""),
		  .pin_mode("O"),
		  .por_state(4),
		  .sio_group_cnt(0),
		  .sio_hyst(1'b0),
		  .sio_ibuf(""),
		  .sio_info(2'b00),
		  .sio_obuf(""),
		  .sio_refsel(""),
		  .sio_vtrip(""),
		  .slew_rate(1'b0),
		  .spanning(0),
		  .use_annotation(1'b0),
		  .vtrip(2'b10),
		  .width(1))
		Servo_1
		 (.oe(tmpOE__Servo_1_net),
		  .y({Net_137}),
		  .fb({tmpFB_0__Servo_1_net[0:0]}),
		  .io({tmpIO_0__Servo_1_net[0:0]}),
		  .siovref(tmpSIOVREF__Servo_1_net),
		  .interrupt({tmpINTERRUPT_0__Servo_1_net[0:0]}),
		  .in_clock({1'b0}),
		  .in_clock_en({1'b1}),
		  .in_reset({1'b0}),
		  .out_clock({1'b0}),
		  .out_clock_en({1'b1}),
		  .out_reset({1'b0}));
	assign tmpOE__Servo_1_net = (`CYDEV_CHIP_MEMBER_USED == `CYDEV_CHIP_MEMBER_3A && `CYDEV_CHIP_REVISION_USED < `CYDEV_CHIP_REVISION_3A_ES3) ? ~{1'b1} : {1'b1};
    SCB_P4_v1_20_2 UART_1 (
        .sclk(Net_161),
        .interrupt(Net_162),
        .clock(1'b0));
	cy_isr_v1_0
		#(.int_type(2'b10))
		ISR_UART_Rx
		 (.int_signal(Net_162));
endmodule