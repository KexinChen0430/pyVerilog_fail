module header
	// Internal signals
		// Generated Signal List
		// End of Generated Signal List
	// %COMPILER_OPTS%
	// Generated Signal Assignments
	// Generated Instances
	// wiring ...
	// Generated Instances and Port Mappings
		// Generated Instance Port Map for dut
		avfb_chip dut (
		);
		// End of Generated Instance Port Map for dut
endmodule