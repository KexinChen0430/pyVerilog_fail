module
CAPB3l
(
input
[
16
:
0
]
CAPB3OI,
input
[
31
:
0
]
PRDATAS0,
input
[
31
:
0
]
PRDATAS1,
input
[
31
:
0
]
PRDATAS2,
input
[
31
:
0
]
PRDATAS3,
input
[
31
:
0
]
PRDATAS4,
input
[
31
:
0
]
PRDATAS5,
input
[
31
:
0
]
PRDATAS6,
input
[
31
:
0
]
PRDATAS7,
input
[
31
:
0
]
PRDATAS8,
input
[
31
:
0
]
PRDATAS9,
input
[
31
:
0
]
PRDATAS10,
input
[
31
:
0
]
PRDATAS11,
input
[
31
:
0
]
PRDATAS12,
input
[
31
:
0
]
PRDATAS13,
input
[
31
:
0
]
PRDATAS14,
input
[
31
:
0
]
PRDATAS15,
input
[
31
:
0
]
PRDATAS16,
input
[
16
:
0
]
CAPB3II,
input
[
16
:
0
]
CAPB3lI,
output
wire
PREADY,
output
wire
PSLVERR,
output
wire
[
31
:
0
]
PRDATA
)
;
localparam
[
4
:
0
]
CAPB3Ol
=
5
'b
00000
;
localparam
[
4
:
0
]
CAPB3Il
=
5
'b
00001
;
localparam
[
4
:
0
]
CAPB3ll
=
5
'b
00010
;
localparam
[
4
:
0
]
CAPB3O0
=
5
'b
00011
;
localparam
[
4
:
0
]
CAPB3I0
=
5
'b
00100
;
localparam
[
4
:
0
]
CAPB3l0
=
5
'b
00101
;
localparam
[
4
:
0
]
CAPB3O1
=
5
'b
00110
;
localparam
[
4
:
0
]
CAPB3I1
=
5
'b
00111
;
localparam
[
4
:
0
]
CAPB3l1
=
5
'b
01000
;
localparam
[
4
:
0
]
CAPB3OOI
=
5
'b
01001
;
localparam
[
4
:
0
]
CAPB3IOI
=
5
'b
01010
;
localparam
[
4
:
0
]
CAPB3lOI
=
5
'b
01011
;
localparam
[
4
:
0
]
CAPB3OII
=
5
'b
01100
;
localparam
[
4
:
0
]
CAPB3III
=
5
'b
01101
;
localparam
[
4
:
0
]
CAPB3lII
=
5
'b
01110
;
localparam
[
4
:
0
]
CAPB3OlI
=
5
'b
01111
;
localparam
[
4
:
0
]
CAPB3IlI
=
5
'b
10000
;
reg
CAPB3llI
;
reg
CAPB3O0I
;
reg
[
31
:
0
]
CAPB3I0I
;
wire
[
4
:
0
]
CAPB3l0I
;
wire
[
31
:
0
]
CAPB3O1I
;
assign
CAPB3O1I
=
32
'b
0
;
assign
CAPB3l0I
[
4
]
=
CAPB3OI
[
16
]
;
assign
CAPB3l0I
[
3
]
=
CAPB3OI
[
15
]
|
CAPB3OI
[
14
]
|
CAPB3OI
[
13
]
|
CAPB3OI
[
12
]
|
CAPB3OI
[
11
]
|
CAPB3OI
[
10
]
|
CAPB3OI
[
9
]
|
CAPB3OI
[
8
]
;
assign
CAPB3l0I
[
2
]
=
CAPB3OI
[
15
]
|
CAPB3OI
[
14
]
|
CAPB3OI
[
13
]
|
CAPB3OI
[
12
]
|
CAPB3OI
[
7
]
|
CAPB3OI
[
6
]
|
CAPB3OI
[
5
]
|
CAPB3OI
[
4
]
;
assign
CAPB3l0I
[
1
]
=
CAPB3OI
[
15
]
|
CAPB3OI
[
14
]
|
CAPB3OI
[
11
]
|
CAPB3OI
[
10
]
|
CAPB3OI
[
7
]
|
CAPB3OI
[
6
]
|
CAPB3OI
[
3
]
|
CAPB3OI
[
2
]
;
assign
CAPB3l0I
[
0
]
=
CAPB3OI
[
15
]
|
CAPB3OI
[
13
]
|
CAPB3OI
[
11
]
|
CAPB3OI
[
9
]
|
CAPB3OI
[
7
]
|
CAPB3OI
[
5
]
|
CAPB3OI
[
3
]
|
CAPB3OI
[
1
]
;
always
@(*)
begin
case
(
CAPB3l0I
)
CAPB3Ol
:
if
(
CAPB3OI
[
0
]
)
CAPB3I0I
[
31
:
0
]
=
PRDATAS0
[
31
:
0
]
;
else
CAPB3I0I
[
31
:
0
]
=
CAPB3O1I
[
31
:
0
]
;
CAPB3Il
:
CAPB3I0I
[
31
:
0
]
=
PRDATAS1
[
31
:
0
]
;
CAPB3ll
:
CAPB3I0I
[
31
:
0
]
=
PRDATAS2
[
31
:
0
]
;
CAPB3O0
:
CAPB3I0I
[
31
:
0
]
=
PRDATAS3
[
31
:
0
]
;
CAPB3I0
:
CAPB3I0I
[
31
:
0
]
=
PRDATAS4
[
31
:
0
]
;
CAPB3l0
:
CAPB3I0I
[
31
:
0
]
=
PRDATAS5
[
31
:
0
]
;
CAPB3O1
:
CAPB3I0I
[
31
:
0
]
=
PRDATAS6
[
31
:
0
]
;
CAPB3I1
:
CAPB3I0I
[
31
:
0
]
=
PRDATAS7
[
31
:
0
]
;
CAPB3l1
:
CAPB3I0I
[
31
:
0
]
=
PRDATAS8
[
31
:
0
]
;
CAPB3OOI
:
CAPB3I0I
[
31
:
0
]
=
PRDATAS9
[
31
:
0
]
;
CAPB3IOI
:
CAPB3I0I
[
31
:
0
]
=
PRDATAS10
[
31
:
0
]
;
CAPB3lOI
:
CAPB3I0I
[
31
:
0
]
=
PRDATAS11
[
31
:
0
]
;
CAPB3OII
:
CAPB3I0I
[
31
:
0
]
=
PRDATAS12
[
31
:
0
]
;
CAPB3III
:
CAPB3I0I
[
31
:
0
]
=
PRDATAS13
[
31
:
0
]
;
CAPB3lII
:
CAPB3I0I
[
31
:
0
]
=
PRDATAS14
[
31
:
0
]
;
CAPB3OlI
:
CAPB3I0I
[
31
:
0
]
=
PRDATAS15
[
31
:
0
]
;
CAPB3IlI
:
CAPB3I0I
[
31
:
0
]
=
PRDATAS16
[
31
:
0
]
;
default
:
CAPB3I0I
[
31
:
0
]
=
CAPB3O1I
[
31
:
0
]
;
endcase
end
always
@(*)
begin
case
(
CAPB3l0I
)
CAPB3Ol
:
if
(
CAPB3OI
[
0
]
)
CAPB3llI
=
CAPB3II
[
0
]
;
else
CAPB3llI
=
1
'b
1
;
CAPB3Il
:
CAPB3llI
=
CAPB3II
[
1
]
;
CAPB3ll
:
CAPB3llI
=
CAPB3II
[
2
]
;
CAPB3O0
:
CAPB3llI
=
CAPB3II
[
3
]
;
CAPB3I0
:
CAPB3llI
=
CAPB3II
[
4
]
;
CAPB3l0
:
CAPB3llI
=
CAPB3II
[
5
]
;
CAPB3O1
:
CAPB3llI
=
CAPB3II
[
6
]
;
CAPB3I1
:
CAPB3llI
=
CAPB3II
[
7
]
;
CAPB3l1
:
CAPB3llI
=
CAPB3II
[
8
]
;
CAPB3OOI
:
CAPB3llI
=
CAPB3II
[
9
]
;
CAPB3IOI
:
CAPB3llI
=
CAPB3II
[
10
]
;
CAPB3lOI
:
CAPB3llI
=
CAPB3II
[
11
]
;
CAPB3OII
:
CAPB3llI
=
CAPB3II
[
12
]
;
CAPB3III
:
CAPB3llI
=
CAPB3II
[
13
]
;
CAPB3lII
:
CAPB3llI
=
CAPB3II
[
14
]
;
CAPB3OlI
:
CAPB3llI
=
CAPB3II
[
15
]
;
CAPB3IlI
:
CAPB3llI
=
CAPB3II
[
16
]
;
default
:
CAPB3llI
=
1
'b
1
;
endcase
end
always
@(*)
begin
case
(
CAPB3l0I
)
CAPB3Ol
:
if
(
CAPB3OI
[
0
]
)
CAPB3O0I
=
CAPB3lI
[
0
]
;
else
CAPB3O0I
=
1
'b
0
;
CAPB3Il
:
CAPB3O0I
=
CAPB3lI
[
1
]
;
CAPB3ll
:
CAPB3O0I
=
CAPB3lI
[
2
]
;
CAPB3O0
:
CAPB3O0I
=
CAPB3lI
[
3
]
;
CAPB3I0
:
CAPB3O0I
=
CAPB3lI
[
4
]
;
CAPB3l0
:
CAPB3O0I
=
CAPB3lI
[
5
]
;
CAPB3O1
:
CAPB3O0I
=
CAPB3lI
[
6
]
;
CAPB3I1
:
CAPB3O0I
=
CAPB3lI
[
7
]
;
CAPB3l1
:
CAPB3O0I
=
CAPB3lI
[
8
]
;
CAPB3OOI
:
CAPB3O0I
=
CAPB3lI
[
9
]
;
CAPB3IOI
:
CAPB3O0I
=
CAPB3lI
[
10
]
;
CAPB3lOI
:
CAPB3O0I
=
CAPB3lI
[
11
]
;
CAPB3OII
:
CAPB3O0I
=
CAPB3lI
[
12
]
;
CAPB3III
:
CAPB3O0I
=
CAPB3lI
[
13
]
;
CAPB3lII
:
CAPB3O0I
=
CAPB3lI
[
14
]
;
CAPB3OlI
:
CAPB3O0I
=
CAPB3lI
[
15
]
;
CAPB3IlI
:
CAPB3O0I
=
CAPB3lI
[
16
]
;
default
:
CAPB3O0I
=
1
'b
0
;
endcase
end
assign
PREADY
=
CAPB3llI
;
assign
PSLVERR
=
CAPB3O0I
;
assign
PRDATA
=
CAPB3I0I
[
31
:
0
]
;
endmodule