module outputs
  wire [63 : 0] word_fst;
  wire [4 : 0] word_snd;
  wire RDY_set_verbosity, valid;
  // inlined wires
  reg [68 : 0] dw_result$wget;
  wire dw_valid$wget, dw_valid$whas;
  // register cfg_verbosity
  reg [3 : 0] cfg_verbosity;
  wire [3 : 0] cfg_verbosity$D_IN;
  wire cfg_verbosity$EN;
  // register requestR
  reg [214 : 0] requestR;
  wire [214 : 0] requestR$D_IN;
  wire requestR$EN;
  // register resultR
  reg [69 : 0] resultR;
  reg [69 : 0] resultR$D_IN;
  wire resultR$EN;
  // register stateR
  reg [1 : 0] stateR;
  reg [1 : 0] stateR$D_IN;
  wire stateR$EN;
  // ports of submodule fpu
  reg [201 : 0] fpu$request_put;
  wire [69 : 0] fpu$response_get;
  wire fpu$EN_request_put,
       fpu$EN_response_get,
       fpu$RDY_request_put,
       fpu$RDY_response_get;
  // ports of submodule frmFpuF
  wire frmFpuF$CLR, frmFpuF$DEQ, frmFpuF$D_IN, frmFpuF$ENQ;
  // rule scheduling signals
  wire CAN_FIRE_RL_doFADD_D,
       CAN_FIRE_RL_doFADD_S,
       CAN_FIRE_RL_doFCLASS_D,
       CAN_FIRE_RL_doFCLASS_S,
       CAN_FIRE_RL_doFCVT_D_L,
       CAN_FIRE_RL_doFCVT_D_LU,
       CAN_FIRE_RL_doFCVT_D_S,
       CAN_FIRE_RL_doFCVT_D_W,
       CAN_FIRE_RL_doFCVT_D_WU,
       CAN_FIRE_RL_doFCVT_LU_D,
       CAN_FIRE_RL_doFCVT_LU_S,
       CAN_FIRE_RL_doFCVT_L_D,
       CAN_FIRE_RL_doFCVT_L_S,
       CAN_FIRE_RL_doFCVT_S_D,
       CAN_FIRE_RL_doFCVT_S_L,
       CAN_FIRE_RL_doFCVT_S_LU,
       CAN_FIRE_RL_doFCVT_S_W,
       CAN_FIRE_RL_doFCVT_S_WU,
       CAN_FIRE_RL_doFCVT_WU_D,
       CAN_FIRE_RL_doFCVT_WU_S,
       CAN_FIRE_RL_doFCVT_W_D,
       CAN_FIRE_RL_doFCVT_W_S,
       CAN_FIRE_RL_doFEQ_D,
       CAN_FIRE_RL_doFEQ_S,
       CAN_FIRE_RL_doFLE_D,
       CAN_FIRE_RL_doFLE_S,
       CAN_FIRE_RL_doFLT_D,
       CAN_FIRE_RL_doFLT_S,
       CAN_FIRE_RL_doFMADD_D,
       CAN_FIRE_RL_doFMADD_S,
       CAN_FIRE_RL_doFMAX_D,
       CAN_FIRE_RL_doFMAX_S,
       CAN_FIRE_RL_doFMIN_D,
       CAN_FIRE_RL_doFMIN_S,
       CAN_FIRE_RL_doFMSUB_D,
       CAN_FIRE_RL_doFMSUB_S,
       CAN_FIRE_RL_doFMUL_D,
       CAN_FIRE_RL_doFMUL_S,
       CAN_FIRE_RL_doFMV_D_X,
       CAN_FIRE_RL_doFMV_W_X,
       CAN_FIRE_RL_doFMV_X_D,
       CAN_FIRE_RL_doFMV_X_W,
       CAN_FIRE_RL_doFNMADD_D,
       CAN_FIRE_RL_doFNMADD_S,
       CAN_FIRE_RL_doFNMSUB_D,
       CAN_FIRE_RL_doFNMSUB_S,
       CAN_FIRE_RL_doFSGNJN_D,
       CAN_FIRE_RL_doFSGNJN_S,
       CAN_FIRE_RL_doFSGNJX_D,
       CAN_FIRE_RL_doFSGNJX_S,
       CAN_FIRE_RL_doFSGNJ_D,
       CAN_FIRE_RL_doFSGNJ_S,
       CAN_FIRE_RL_doFSUB_D,
       CAN_FIRE_RL_doFSUB_S,
       CAN_FIRE_RL_rl_drive_fpu_result,
       CAN_FIRE_RL_rl_get_fpu_result,
       CAN_FIRE_req,
       CAN_FIRE_set_verbosity,
       WILL_FIRE_RL_doFADD_D,
       WILL_FIRE_RL_doFADD_S,
       WILL_FIRE_RL_doFCLASS_D,
       WILL_FIRE_RL_doFCLASS_S,
       WILL_FIRE_RL_doFCVT_D_L,
       WILL_FIRE_RL_doFCVT_D_LU,
       WILL_FIRE_RL_doFCVT_D_S,
       WILL_FIRE_RL_doFCVT_D_W,
       WILL_FIRE_RL_doFCVT_D_WU,
       WILL_FIRE_RL_doFCVT_LU_D,
       WILL_FIRE_RL_doFCVT_LU_S,
       WILL_FIRE_RL_doFCVT_L_D,
       WILL_FIRE_RL_doFCVT_L_S,
       WILL_FIRE_RL_doFCVT_S_D,
       WILL_FIRE_RL_doFCVT_S_L,
       WILL_FIRE_RL_doFCVT_S_LU,
       WILL_FIRE_RL_doFCVT_S_W,
       WILL_FIRE_RL_doFCVT_S_WU,
       WILL_FIRE_RL_doFCVT_WU_D,
       WILL_FIRE_RL_doFCVT_WU_S,
       WILL_FIRE_RL_doFCVT_W_D,
       WILL_FIRE_RL_doFCVT_W_S,
       WILL_FIRE_RL_doFEQ_D,
       WILL_FIRE_RL_doFEQ_S,
       WILL_FIRE_RL_doFLE_D,
       WILL_FIRE_RL_doFLE_S,
       WILL_FIRE_RL_doFLT_D,
       WILL_FIRE_RL_doFLT_S,
       WILL_FIRE_RL_doFMADD_D,
       WILL_FIRE_RL_doFMADD_S,
       WILL_FIRE_RL_doFMAX_D,
       WILL_FIRE_RL_doFMAX_S,
       WILL_FIRE_RL_doFMIN_D,
       WILL_FIRE_RL_doFMIN_S,
       WILL_FIRE_RL_doFMSUB_D,
       WILL_FIRE_RL_doFMSUB_S,
       WILL_FIRE_RL_doFMUL_D,
       WILL_FIRE_RL_doFMUL_S,
       WILL_FIRE_RL_doFMV_D_X,
       WILL_FIRE_RL_doFMV_W_X,
       WILL_FIRE_RL_doFMV_X_D,
       WILL_FIRE_RL_doFMV_X_W,
       WILL_FIRE_RL_doFNMADD_D,
       WILL_FIRE_RL_doFNMADD_S,
       WILL_FIRE_RL_doFNMSUB_D,
       WILL_FIRE_RL_doFNMSUB_S,
       WILL_FIRE_RL_doFSGNJN_D,
       WILL_FIRE_RL_doFSGNJN_S,
       WILL_FIRE_RL_doFSGNJX_D,
       WILL_FIRE_RL_doFSGNJX_S,
       WILL_FIRE_RL_doFSGNJ_D,
       WILL_FIRE_RL_doFSGNJ_S,
       WILL_FIRE_RL_doFSUB_D,
       WILL_FIRE_RL_doFSUB_S,
       WILL_FIRE_RL_rl_drive_fpu_result,
       WILL_FIRE_RL_rl_get_fpu_result,
       WILL_FIRE_req,
       WILL_FIRE_set_verbosity;
  // inputs to muxes for submodule ports
  wire [201 : 0] MUX_fpu$request_put_1__VAL_1,
		 MUX_fpu$request_put_1__VAL_10,
		 MUX_fpu$request_put_1__VAL_11,
		 MUX_fpu$request_put_1__VAL_12,
		 MUX_fpu$request_put_1__VAL_13,
		 MUX_fpu$request_put_1__VAL_14,
		 MUX_fpu$request_put_1__VAL_2,
		 MUX_fpu$request_put_1__VAL_3,
		 MUX_fpu$request_put_1__VAL_4,
		 MUX_fpu$request_put_1__VAL_5,
		 MUX_fpu$request_put_1__VAL_6,
		 MUX_fpu$request_put_1__VAL_7,
		 MUX_fpu$request_put_1__VAL_8,
		 MUX_fpu$request_put_1__VAL_9;
  wire [69 : 0] MUX_resultR$write_1__VAL_10,
		MUX_resultR$write_1__VAL_11,
		MUX_resultR$write_1__VAL_12,
		MUX_resultR$write_1__VAL_13,
		MUX_resultR$write_1__VAL_14,
		MUX_resultR$write_1__VAL_15,
		MUX_resultR$write_1__VAL_16,
		MUX_resultR$write_1__VAL_17,
		MUX_resultR$write_1__VAL_18,
		MUX_resultR$write_1__VAL_19,
		MUX_resultR$write_1__VAL_2,
		MUX_resultR$write_1__VAL_20,
		MUX_resultR$write_1__VAL_21,
		MUX_resultR$write_1__VAL_22,
		MUX_resultR$write_1__VAL_23,
		MUX_resultR$write_1__VAL_24,
		MUX_resultR$write_1__VAL_25,
		MUX_resultR$write_1__VAL_26,
		MUX_resultR$write_1__VAL_27,
		MUX_resultR$write_1__VAL_28,
		MUX_resultR$write_1__VAL_29,
		MUX_resultR$write_1__VAL_3,
		MUX_resultR$write_1__VAL_30,
		MUX_resultR$write_1__VAL_31,
		MUX_resultR$write_1__VAL_32,
		MUX_resultR$write_1__VAL_33,
		MUX_resultR$write_1__VAL_34,
		MUX_resultR$write_1__VAL_35,
		MUX_resultR$write_1__VAL_36,
		MUX_resultR$write_1__VAL_37,
		MUX_resultR$write_1__VAL_38,
		MUX_resultR$write_1__VAL_39,
		MUX_resultR$write_1__VAL_4,
		MUX_resultR$write_1__VAL_40,
		MUX_resultR$write_1__VAL_41,
		MUX_resultR$write_1__VAL_42,
		MUX_resultR$write_1__VAL_6,
		MUX_resultR$write_1__VAL_7,
		MUX_resultR$write_1__VAL_8,
		MUX_resultR$write_1__VAL_9;
  wire [68 : 0] MUX_dw_result$wset_1__VAL_1,
		MUX_dw_result$wset_1__VAL_10,
		MUX_dw_result$wset_1__VAL_11,
		MUX_dw_result$wset_1__VAL_12,
		MUX_dw_result$wset_1__VAL_13,
		MUX_dw_result$wset_1__VAL_14,
		MUX_dw_result$wset_1__VAL_15,
		MUX_dw_result$wset_1__VAL_16,
		MUX_dw_result$wset_1__VAL_17,
		MUX_dw_result$wset_1__VAL_18,
		MUX_dw_result$wset_1__VAL_19,
		MUX_dw_result$wset_1__VAL_2,
		MUX_dw_result$wset_1__VAL_20,
		MUX_dw_result$wset_1__VAL_21,
		MUX_dw_result$wset_1__VAL_22,
		MUX_dw_result$wset_1__VAL_23,
		MUX_dw_result$wset_1__VAL_24,
		MUX_dw_result$wset_1__VAL_25,
		MUX_dw_result$wset_1__VAL_26,
		MUX_dw_result$wset_1__VAL_27,
		MUX_dw_result$wset_1__VAL_28,
		MUX_dw_result$wset_1__VAL_29,
		MUX_dw_result$wset_1__VAL_3,
		MUX_dw_result$wset_1__VAL_30,
		MUX_dw_result$wset_1__VAL_31,
		MUX_dw_result$wset_1__VAL_32,
		MUX_dw_result$wset_1__VAL_33,
		MUX_dw_result$wset_1__VAL_34,
		MUX_dw_result$wset_1__VAL_35,
		MUX_dw_result$wset_1__VAL_36,
		MUX_dw_result$wset_1__VAL_37,
		MUX_dw_result$wset_1__VAL_38,
		MUX_dw_result$wset_1__VAL_39,
		MUX_dw_result$wset_1__VAL_4,
		MUX_dw_result$wset_1__VAL_40,
		MUX_dw_result$wset_1__VAL_5,
		MUX_dw_result$wset_1__VAL_6,
		MUX_dw_result$wset_1__VAL_7,
		MUX_dw_result$wset_1__VAL_8,
		MUX_dw_result$wset_1__VAL_9;
  wire MUX_dw_result$wset_1__SEL_1,
       MUX_dw_result$wset_1__SEL_2,
       MUX_dw_result$wset_1__SEL_38;
  // remaining internal signals
  reg [51 : 0] CASE_guard0287_0b0_sfd___30277_BITS_54_TO_3_0b_ETC__q79,
	       CASE_guard0287_0b0_sfd___30277_BITS_54_TO_3_0b_ETC__q80,
	       CASE_guard0712_0b0_sfd___39973_BITS_53_TO_2_0b_ETC__q88,
	       CASE_guard0712_0b0_sfd___39973_BITS_53_TO_2_0b_ETC__q89,
	       CASE_guard1017_0b0_sfd___30277_BITS_53_TO_2_0b_ETC__q75,
	       CASE_guard1017_0b0_sfd___30277_BITS_53_TO_2_0b_ETC__q76,
	       CASE_guard3828_0b0_sfd___31835_BITS_63_TO_12_0_ETC__q104,
	       CASE_guard3828_0b0_sfd___31835_BITS_63_TO_12_0_ETC__q105,
	       CASE_guard4558_0b0_sfd___31835_BITS_62_TO_11_0_ETC__q100,
	       CASE_guard4558_0b0_sfd___31835_BITS_62_TO_11_0_ETC__q101,
	       CASE_guard4840_0b0_sfd___32457_BITS_63_TO_12_0_ETC__q110,
	       CASE_guard4840_0b0_sfd___32457_BITS_63_TO_12_0_ETC__q111,
	       CASE_guard5569_0b0_sfd___32457_BITS_62_TO_11_0_ETC__q108,
	       CASE_guard5569_0b0_sfd___32457_BITS_62_TO_11_0_ETC__q109,
	       CASE_guard61118_0b0_theResult___snd69030_BITS__ETC__q168,
	       CASE_guard61118_0b0_theResult___snd69030_BITS__ETC__q169,
	       CASE_guard70426_0b0_sfdin78646_BITS_56_TO_5_0b_ETC__q170,
	       CASE_guard70426_0b0_sfdin78646_BITS_56_TO_5_0b_ETC__q171,
	       CASE_guard79493_0b0_theResult___snd87429_BITS__ETC__q172,
	       CASE_guard79493_0b0_theResult___snd87429_BITS__ETC__q173,
	       CASE_guard9983_0b0_sfd___39973_BITS_54_TO_3_0b_ETC__q90,
	       CASE_guard9983_0b0_sfd___39973_BITS_54_TO_3_0b_ETC__q91,
	       CASE_requestR_BITS_194_TO_192_0x1_450359962737_ETC__q5,
	       IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d2365,
	       IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d2383,
	       IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d2551,
	       IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d2566,
	       IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d2900,
	       IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d2918,
	       IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d3056,
	       IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d3071,
	       IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d4982,
	       IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d5009,
	       IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d5028;
  reg [22 : 0] CASE_guard11367_0b0_sfdin19458_BITS_56_TO_34_0_ETC__q134,
	       CASE_guard11367_0b0_sfdin19458_BITS_56_TO_34_0_ETC__q135,
	       CASE_guard1845_0b0_sfd___31835_BITS_63_TO_41_0_ETC__q18,
	       CASE_guard1845_0b0_sfd___31835_BITS_63_TO_41_0_ETC__q19,
	       CASE_guard20102_0b0_theResult___snd28101_BITS__ETC__q132,
	       CASE_guard20102_0b0_theResult___snd28101_BITS__ETC__q133,
	       CASE_guard2375_0b0_sfd___31835_BITS_62_TO_40_0_ETC__q20,
	       CASE_guard2375_0b0_sfd___31835_BITS_62_TO_40_0_ETC__q21,
	       CASE_guard2467_0b0_sfd___32457_BITS_63_TO_41_0_ETC__q36,
	       CASE_guard2467_0b0_sfd___32457_BITS_63_TO_41_0_ETC__q37,
	       CASE_guard29091_0b0_sfdin37311_BITS_56_TO_34_0_ETC__q136,
	       CASE_guard29091_0b0_sfdin37311_BITS_56_TO_34_0_ETC__q137,
	       CASE_guard2993_0b0_sfd___32457_BITS_62_TO_40_0_ETC__q34,
	       CASE_guard2993_0b0_sfd___32457_BITS_62_TO_40_0_ETC__q35,
	       CASE_guard37955_0b0_theResult___snd45978_BITS__ETC__q138,
	       CASE_guard37955_0b0_theResult___snd45978_BITS__ETC__q139,
	       CASE_guard5065_0b0_sfd___35055_BITS_31_TO_9_0b_ETC__q61,
	       CASE_guard5065_0b0_sfd___35055_BITS_31_TO_9_0b_ETC__q62,
	       CASE_guard5591_0b0_sfd___35055_BITS_30_TO_8_0b_ETC__q59,
	       CASE_guard5591_0b0_sfd___35055_BITS_30_TO_8_0b_ETC__q60,
	       CASE_guard8894_0b0_sfd___38884_BITS_31_TO_9_0b_ETC__q48,
	       CASE_guard8894_0b0_sfd___38884_BITS_31_TO_9_0b_ETC__q49,
	       CASE_guard9421_0b0_sfd___38884_BITS_30_TO_8_0b_ETC__q50,
	       CASE_guard9421_0b0_sfd___38884_BITS_30_TO_8_0b_ETC__q51,
	       CASE_requestR_BITS_194_TO_192_0x1_8388607_0x2__ETC__q3,
	       IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d1008,
	       IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d1023,
	       IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d1390,
	       IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d1408,
	       IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d1613,
	       IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d1628,
	       IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d4149,
	       IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d4168,
	       IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d4195,
	       IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d4214,
	       IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d531,
	       IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d549;
  reg [10 : 0] CASE_guard0287_0b0_0_0b1_0_0b10_out_exp0906_0b_ETC__q78,
	       CASE_guard0287_0b0_0_0b1_theResult___exp0903_0_ETC__q77,
	       CASE_guard0712_0b0_x0727_BITS_10_TO_0_0b1_theR_ETC__q86,
	       CASE_guard0712_0b0_x0727_BITS_10_TO_0_0b1_x072_ETC__q87,
	       CASE_guard1017_0b0_x1032_BITS_10_TO_0_0b1_theR_ETC__q73,
	       CASE_guard1017_0b0_x1032_BITS_10_TO_0_0b1_x103_ETC__q74,
	       CASE_guard3828_0b0_0_0b1_0_0b10_out_exp4447_0b_ETC__q103,
	       CASE_guard3828_0b0_0_0b1_theResult___exp4444_0_ETC__q102,
	       CASE_guard4558_0b0_x4573_BITS_10_TO_0_0b1_theR_ETC__q98,
	       CASE_guard4558_0b0_x4573_BITS_10_TO_0_0b1_x457_ETC__q99,
	       CASE_guard4840_0b0_0_0b1_0_0b10_out_exp5459_0b_ETC__q29,
	       CASE_guard4840_0b0_0_0b1_theResult___exp5456_0_ETC__q30,
	       CASE_guard5569_0b0_x5584_BITS_10_TO_0_0b1_theR_ETC__q106,
	       CASE_guard5569_0b0_x5584_BITS_10_TO_0_0b1_x558_ETC__q107,
	       CASE_guard61118_0b0_theResult___fst_exp69079_0_ETC__q156,
	       CASE_guard61118_0b0_theResult___fst_exp69079_0_ETC__q157,
	       CASE_guard70426_0b0_theResult___fst_exp78652_0_ETC__q158,
	       CASE_guard70426_0b0_theResult___fst_exp78652_0_ETC__q159,
	       CASE_guard79493_0b0_theResult___fst_exp87483_0_ETC__q160,
	       CASE_guard79493_0b0_theResult___fst_exp87483_0_ETC__q161,
	       CASE_guard9983_0b0_0_0b1_0_0b10_out_exp0602_0b_ETC__q83,
	       CASE_guard9983_0b0_0_0b1_theResult___exp0599_0_ETC__q84,
	       CASE_requestR_BITS_194_TO_192_0x1_2046_0x2_IF__ETC__q4,
	       CASE_requestR_BITS_194_TO_192_0x3_IF_guard4840_ETC__q31,
	       CASE_requestR_BITS_194_TO_192_0x3_IF_guard9983_ETC__q85,
	       IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d2313,
	       IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d2342,
	       IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d2529,
	       IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d2848,
	       IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d2877,
	       IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d3033,
	       IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d4555,
	       IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d4880,
	       IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d4949;
  reg [7 : 0] CASE_guard11367_0b0_theResult___fst_exp19464_0_ETC__q124,
	      CASE_guard11367_0b0_theResult___fst_exp19464_0_ETC__q125,
	      CASE_guard1845_0b0_0_0b1_0_0b10_out_exp2264_0b_ETC__q15,
	      CASE_guard1845_0b0_0_0b1_theResult___exp2261_0_ETC__q14,
	      CASE_guard20102_0b0_theResult___fst_exp28150_0_ETC__q126,
	      CASE_guard20102_0b0_theResult___fst_exp28150_0_ETC__q127,
	      CASE_guard2375_0b0_x2390_BITS_7_TO_0_0b1_theRe_ETC__q16,
	      CASE_guard2375_0b0_x2390_BITS_7_TO_0_0b1_x2390_ETC__q17,
	      CASE_guard2467_0b0_0_0b1_0_0b10_out_exp2883_0b_ETC__q26,
	      CASE_guard2467_0b0_0_0b1_theResult___exp2880_0_ETC__q27,
	      CASE_guard29091_0b0_theResult___fst_exp37317_0_ETC__q128,
	      CASE_guard29091_0b0_theResult___fst_exp37317_0_ETC__q129,
	      CASE_guard2993_0b0_x3008_BITS_7_TO_0_0b1_theRe_ETC__q32,
	      CASE_guard2993_0b0_x3008_BITS_7_TO_0_0b1_x3008_ETC__q33,
	      CASE_guard37955_0b0_theResult___fst_exp46032_0_ETC__q130,
	      CASE_guard37955_0b0_theResult___fst_exp46032_0_ETC__q131,
	      CASE_guard5065_0b0_0_0b1_0_0b10_out_exp5481_0b_ETC__q54,
	      CASE_guard5065_0b0_0_0b1_theResult___exp5478_0_ETC__q55,
	      CASE_guard5591_0b0_x5606_BITS_7_TO_0_0b1_theRe_ETC__q57,
	      CASE_guard5591_0b0_x5606_BITS_7_TO_0_0b1_x5606_ETC__q58,
	      CASE_guard8894_0b0_0_0b1_0_0b10_out_exp9310_0b_ETC__q45,
	      CASE_guard8894_0b0_0_0b1_theResult___exp9307_0_ETC__q44,
	      CASE_guard9421_0b0_x9436_BITS_7_TO_0_0b1_theRe_ETC__q46,
	      CASE_guard9421_0b0_x9436_BITS_7_TO_0_0b1_x9436_ETC__q47,
	      CASE_requestR_BITS_194_TO_192_0x1_254_0x2_IF_r_ETC__q2,
	      CASE_requestR_BITS_194_TO_192_0x3_IF_guard2467_ETC__q28,
	      CASE_requestR_BITS_194_TO_192_0x3_IF_guard5065_ETC__q56,
	      IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d1338,
	      IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d1367,
	      IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d1590,
	      IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d3602,
	      IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d3719,
	      IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d4046,
	      IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d4115,
	      IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d479,
	      IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d508,
	      IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d985;
  reg [2 : 0] IF_requestR_BITS_194_TO_192_0_EQ_0x0_1_THEN_re_ETC___d40;
  reg CASE_guard0287_0b0_requestR_BIT_159_0b1_reques_ETC__q69,
      CASE_guard1017_0b0_requestR_BIT_159_0b1_reques_ETC__q71,
      CASE_guard11367_0b0_requestR_BIT_191_0b1_reque_ETC__q140,
      CASE_guard1845_0b0_requestR_BIT_191_0b1_reques_ETC__q10,
      CASE_guard20102_0b0_requestR_BIT_191_0b1_reque_ETC__q142,
      CASE_guard2375_0b0_requestR_BIT_191_0b1_reques_ETC__q12,
      CASE_guard29091_0b0_requestR_BIT_191_0b1_reque_ETC__q144,
      CASE_guard37955_0b0_requestR_BIT_191_0b1_reque_ETC__q146,
      CASE_guard3828_0b0_requestR_BIT_191_0b1_reques_ETC__q94,
      CASE_guard4558_0b0_requestR_BIT_191_0b1_reques_ETC__q96,
      CASE_guard61118_0b0_requestR_BITS_191_TO_160_E_ETC__q162,
      CASE_guard70426_0b0_requestR_BITS_191_TO_160_E_ETC__q164,
      CASE_guard79493_0b0_requestR_BITS_191_TO_160_E_ETC__q166,
      CASE_guard8894_0b0_requestR_BIT_159_0b1_reques_ETC__q40,
      CASE_guard9421_0b0_requestR_BIT_159_0b1_reques_ETC__q42,
      CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q11,
      CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q13,
      CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q141,
      CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q143,
      CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q145,
      CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q147,
      CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q163,
      CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q165,
      CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q167,
      CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q41,
      CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q43,
      CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q70,
      CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q72,
      CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q95,
      CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q97;
  wire [117 : 0] IF_requestR_BIT_191_27_THEN_NEG_0b0_CONCAT_NOT_ETC___d3109,
		 b__h96976,
		 x__h97876,
		 x__h99175;
  wire [88 : 0] IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d1689,
		b__h36799,
		x__h37699,
		x__h39015;
  wire [85 : 0] IF_requestR_BIT_191_27_THEN_NEG_0b0_CONCAT_NOT_ETC___d2620,
		b__h72122,
		x__h72798,
		x__h73876;
  wire [68 : 0] ab__h206728;
  wire [64 : 0] _1_CONCAT_DONTCARE_CONCAT_requestR_BITS_63_TO_3_ETC___d68,
		_theResult_____2__h36734,
		_theResult_____2__h96911,
		out1___1__h37450,
		out1___1__h97627;
  wire [63 : 0] IF_IF_requestR_BITS_127_TO_96_2_EQ_0xFFFFFFFF__ETC___d2040,
		IF_IF_requestR_BITS_127_TO_96_2_EQ_0xFFFFFFFF__ETC___d2056,
		IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_ETC___d1748,
		IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_ETC___d1807,
		IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_ETC___d2039,
		IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_ETC___d2041,
		IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_ETC___d2055,
		IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_ETC___d2057,
		IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_ETC___d2127,
		IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_ETC___d2128,
		IF_NEG_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0_ETC___d1744,
		IF_NEG_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0_ETC___d1746,
		IF_NEG_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0_ETC___d1805,
		IF_NEG_SEXT_requestR_BITS_190_TO_180_599_MINUS_ETC___d3164,
		IF_NEG_SEXT_requestR_BITS_190_TO_180_599_MINUS_ETC___d3166,
		IF_NEG_SEXT_requestR_BITS_190_TO_180_599_MINUS_ETC___d3219,
		IF_requestR_BITS_126_TO_116_166_EQ_2047_167_AN_ETC___d5214,
		IF_requestR_BITS_190_TO_180_599_EQ_0_609_AND_r_ETC___d3221,
		IF_requestR_BITS_190_TO_180_599_EQ_0_609_AND_r_ETC___d5228,
		IF_requestR_BITS_190_TO_180_599_EQ_0_609_AND_r_ETC___d5299,
		IF_requestR_BITS_190_TO_180_599_EQ_2047_600_AN_ETC___d3168,
		IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d1677,
		IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d1809,
		IF_requestR_BIT_191_27_THEN_922337203685477580_ETC___d3105,
		res___1__h205637,
		res___1__h206075,
		res___1__h206085,
		res___1__h206104,
		res___1__h50736,
		res___1__h50972,
		res___1__h50982,
		res___1__h51001,
		res__h147098,
		res__h188903,
		res__h193345,
		res__h197893,
		res__h200597,
		res__h203292,
		res__h205169,
		res__h206120,
		res__h206301,
		res__h42340,
		res__h42577,
		res__h47949,
		res__h49432,
		res__h50501,
		res__h51017,
		sfd___3__h11835,
		sfd___3__h22457,
		sfd__h2230,
		x__h13371,
		x__h148202,
		x__h1781,
		x__h189928,
		x__h1927,
		x__h194476,
		x__h198920,
		x__h201615,
		x__h203492,
		x__h205619,
		x__h2061,
		x__h206269,
		x__h2209,
		x__h23959,
		x__h30414,
		x__h36556,
		x__h38594,
		x__h39336,
		x__h40912,
		x__h41662,
		x__h44296,
		x__h46821,
		x__h46942,
		x__h47080,
		x__h48563,
		x__h49632,
		x__h50718,
		x__h51885,
		x__h52007,
		x__h52131,
		x__h52261,
		x__h62209,
		x__h71876,
		x__h73452,
		x__h74198,
		x__h85750,
		x__h96733,
		x__h98754,
		x__h99497;
  wire [56 : 0] IF_0_CONCAT_IF_IF_0b0_CONCAT_NOT_requestR_BITS_ETC__q114,
		IF_0_CONCAT_IF_IF_3074_MINUS_SEXT_IF_requestR__ETC__q151,
		IF_0_CONCAT_IF_IF_3970_MINUS_SEXT_requestR_BIT_ETC__q119,
		IF_0_CONCAT_IF_IF_requestR_BITS_191_TO_160_4_E_ETC__q148,
		IF_0_CONCAT_IF_IF_requestR_BITS_191_TO_160_4_E_ETC__q154,
		IF_0_CONCAT_IF_requestR_BITS_190_TO_180_599_EQ_ETC__q116,
		IF_0_CONCAT_IF_requestR_BITS_190_TO_180_599_EQ_ETC__q122,
		IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d1838,
		_0b0_CONCAT_NOT_IF_requestR_BITS_191_TO_160_4_E_ETC___d4573,
		_0b0_CONCAT_NOT_requestR_BITS_190_TO_180_599_EQ_ETC___d3741,
		_theResult____h111357,
		_theResult____h129081,
		_theResult____h170416,
		_theResult___snd__h119475,
		_theResult___snd__h119486,
		_theResult___snd__h119488,
		_theResult___snd__h119498,
		_theResult___snd__h119504,
		_theResult___snd__h119527,
		_theResult___snd__h128101,
		_theResult___snd__h128103,
		_theResult___snd__h128110,
		_theResult___snd__h128116,
		_theResult___snd__h128139,
		_theResult___snd__h137328,
		_theResult___snd__h137339,
		_theResult___snd__h137341,
		_theResult___snd__h137351,
		_theResult___snd__h137357,
		_theResult___snd__h137380,
		_theResult___snd__h145978,
		_theResult___snd__h145992,
		_theResult___snd__h145998,
		_theResult___snd__h146016,
		_theResult___snd__h169030,
		_theResult___snd__h169032,
		_theResult___snd__h169039,
		_theResult___snd__h169045,
		_theResult___snd__h169068,
		_theResult___snd__h178663,
		_theResult___snd__h178674,
		_theResult___snd__h178676,
		_theResult___snd__h178686,
		_theResult___snd__h178692,
		_theResult___snd__h178715,
		_theResult___snd__h187429,
		_theResult___snd__h187443,
		_theResult___snd__h187449,
		_theResult___snd__h187467,
		b__h39582,
		result__h129694,
		result__h171029,
		sfd__h103727,
		sfdin__h119458,
		sfdin__h137311,
		sfdin__h178646,
		x__h129789,
		x__h171124,
		x__h40258,
		x__h41336;
  wire [54 : 0] sfd___3__h60277, sfd___3__h69973, sfd__h52276, sfd__h62221;
  wire [53 : 0] sfd__h169097,
		sfd__h178744,
		sfd__h187502,
		sfd__h60304,
		sfd__h61047,
		sfd__h70000,
		sfd__h70742,
		sfd__h83845,
		sfd__h84588,
		sfd__h94857,
		sfd__h95599,
		value__h72124;
  wire [51 : 0] IF_IF_IF_IF_3074_MINUS_SEXT_IF_requestR_BITS_1_ETC___d5003,
		IF_IF_IF_IF_3074_MINUS_SEXT_IF_requestR_BITS_1_ETC___d5005,
		IF_IF_IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFF_ETC___d4976,
		IF_IF_IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFF_ETC___d4978,
		IF_IF_IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFF_ETC___d5022,
		IF_IF_IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFF_ETC___d5024,
		IF_IF_IF_requestR_BIT_159_6_THEN_NEG_requestR__ETC___d2359,
		IF_IF_IF_requestR_BIT_159_6_THEN_NEG_requestR__ETC___d2361,
		IF_IF_IF_requestR_BIT_159_6_THEN_NEG_requestR__ETC___d2377,
		IF_IF_IF_requestR_BIT_159_6_THEN_NEG_requestR__ETC___d2379,
		IF_IF_IF_requestR_BIT_191_27_THEN_NEG_requestR_ETC___d2894,
		IF_IF_IF_requestR_BIT_191_27_THEN_NEG_requestR_ETC___d2896,
		IF_IF_IF_requestR_BIT_191_27_THEN_NEG_requestR_ETC___d2912,
		IF_IF_IF_requestR_BIT_191_27_THEN_NEG_requestR_ETC___d2914,
		IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_ETC___d5035,
		IF_requestR_BITS_159_TO_128_121_EQ_0_122_OR_NO_ETC___d2387,
		IF_requestR_BITS_159_TO_128_121_EQ_0_122_OR_NO_ETC___d2570,
		_theResult___fst_sfd__h100023,
		_theResult___fst_sfd__h154007,
		_theResult___fst_sfd__h169833,
		_theResult___fst_sfd__h169836,
		_theResult___fst_sfd__h179480,
		_theResult___fst_sfd__h179483,
		_theResult___fst_sfd__h188262,
		_theResult___fst_sfd__h188265,
		_theResult___fst_sfd__h188274,
		_theResult___fst_sfd__h188280,
		_theResult___fst_sfd__h61001,
		_theResult___fst_sfd__h61757,
		_theResult___fst_sfd__h61760,
		_theResult___fst_sfd__h70696,
		_theResult___fst_sfd__h71451,
		_theResult___fst_sfd__h71454,
		_theResult___fst_sfd__h84542,
		_theResult___fst_sfd__h85298,
		_theResult___fst_sfd__h85301,
		_theResult___fst_sfd__h95553,
		_theResult___fst_sfd__h96308,
		_theResult___fst_sfd__h96311,
		_theResult___sfd__h169735,
		_theResult___sfd__h179382,
		_theResult___sfd__h188164,
		_theResult___sfd__h60904,
		_theResult___sfd__h61660,
		_theResult___sfd__h70600,
		_theResult___sfd__h71355,
		_theResult___sfd__h84445,
		_theResult___sfd__h85201,
		_theResult___sfd__h95457,
		_theResult___sfd__h96212,
		_theResult___snd_fst_sfd__h150153,
		_theResult___snd_fst_sfd__h169839,
		_theResult___snd_fst_sfd__h188268,
		_theResult___snd_fst_sfd__h61763,
		_theResult___snd_fst_sfd__h71457,
		_theResult___snd_fst_sfd__h85304,
		_theResult___snd_fst_sfd__h96314,
		out___1_sfd__h148267,
		out_sfd__h169738,
		out_sfd__h179385,
		out_sfd__h188167,
		out_sfd__h60907,
		out_sfd__h61663,
		out_sfd__h70603,
		out_sfd__h71358,
		out_sfd__h84448,
		out_sfd__h85204,
		out_sfd__h95460,
		out_sfd__h96215,
		value__h99566;
  wire [32 : 0] _theResult_____2__h39517,
		_theResult_____2__h72057,
		out1___1__h40009,
		out1___1__h72549;
  wire [31 : 0] IF_IF_requestR_BITS_127_TO_96_2_EQ_0xFFFFFFFF__ETC___d2036,
		IF_IF_requestR_BITS_127_TO_96_2_EQ_0xFFFFFFFF__ETC___d2050,
		IF_IF_requestR_BITS_127_TO_96_2_EQ_0xFFFFFFFF__ETC___d2052,
		IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_ETC___d1897,
		IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_ETC___d1951,
		IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_ETC___d2037,
		IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_ETC___d2053,
		IF_NEG_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0_ETC___d1893,
		IF_NEG_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0_ETC___d1895,
		IF_NEG_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0_ETC___d1949,
		IF_NEG_SEXT_requestR_BITS_190_TO_180_599_MINUS_ETC___d2675,
		IF_NEG_SEXT_requestR_BITS_190_TO_180_599_MINUS_ETC___d2677,
		IF_NEG_SEXT_requestR_BITS_190_TO_180_599_MINUS_ETC___d2737,
		IF_NOT_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFF_ETC___d2034,
		IF_NOT_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFF_ETC___d2049,
		IF_requestR_BITS_190_TO_180_599_EQ_0_609_AND_r_ETC___d2739,
		IF_requestR_BITS_190_TO_180_599_EQ_2047_600_AN_ETC___d2679,
		IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d1834,
		IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d1953,
		IF_requestR_BIT_191_27_THEN_2147483648_ELSE_21_ETC___d2608,
		requestR_BITS_127_TO_96_2_EQ_0xFFFFFFFF_3_AND__ETC___d28,
		requestR_BITS_159_TO_128__q1,
		sfd___3__h28884,
		sfd___3__h35055,
		sfd__h23980,
		x__h147104,
		x__h1787,
		x__h1933,
		x__h2067,
		x__h2215,
		x__h23965,
		x__h39339,
		x__h40915,
		x__h71879,
		x__h73455;
  wire [30 : 0] IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d19;
  wire [24 : 0] sfd__h11862,
		sfd__h119556,
		sfd__h12405,
		sfd__h128168,
		sfd__h137409,
		sfd__h146051,
		sfd__h22484,
		sfd__h23023,
		sfd__h28911,
		sfd__h29451,
		sfd__h35082,
		sfd__h35621,
		value__h36801;
  wire [23 : 0] NEG_SEXT_requestR_BITS_190_TO_180_599_MINUS_10_ETC___d2613,
		NEG_SEXT_requestR_BITS_190_TO_180_599_MINUS_10_ETC___d2645,
		NEG_SEXT_requestR_BITS_190_TO_180_599_MINUS_10_ETC___d2646,
		NEG_SEXT_requestR_BITS_190_TO_180_599_MINUS_10_ETC___d2710,
		NEG_SEXT_requestR_BITS_190_TO_180_599_MINUS_10_ETC___d3134,
		NEG_SEXT_requestR_BITS_190_TO_180_599_MINUS_10_ETC___d3135,
		NEG_SEXT_requestR_BITS_190_TO_180_599_MINUS_10_ETC___d3192;
  wire [22 : 0] IF_IF_IF_IF_0b0_CONCAT_NOT_requestR_BITS_190_T_ETC___d4143,
		IF_IF_IF_IF_0b0_CONCAT_NOT_requestR_BITS_190_T_ETC___d4145,
		IF_IF_IF_IF_3970_MINUS_SEXT_requestR_BITS_190__ETC___d4189,
		IF_IF_IF_IF_3970_MINUS_SEXT_requestR_BITS_190__ETC___d4191,
		IF_IF_IF_requestR_BITS_190_TO_180_599_EQ_0_609_ETC___d4162,
		IF_IF_IF_requestR_BITS_190_TO_180_599_EQ_0_609_ETC___d4164,
		IF_IF_IF_requestR_BITS_190_TO_180_599_EQ_0_609_ETC___d4208,
		IF_IF_IF_requestR_BITS_190_TO_180_599_EQ_0_609_ETC___d4210,
		IF_IF_IF_requestR_BIT_159_6_THEN_NEG_requestR__ETC___d1384,
		IF_IF_IF_requestR_BIT_159_6_THEN_NEG_requestR__ETC___d1386,
		IF_IF_IF_requestR_BIT_159_6_THEN_NEG_requestR__ETC___d1402,
		IF_IF_IF_requestR_BIT_159_6_THEN_NEG_requestR__ETC___d1404,
		IF_IF_IF_requestR_BIT_191_27_THEN_NEG_requestR_ETC___d525,
		IF_IF_IF_requestR_BIT_191_27_THEN_NEG_requestR_ETC___d527,
		IF_IF_IF_requestR_BIT_191_27_THEN_NEG_requestR_ETC___d543,
		IF_IF_IF_requestR_BIT_191_27_THEN_NEG_requestR_ETC___d545,
		IF_requestR_BITS_190_TO_180_599_EQ_2047_600_AN_ETC___d4221,
		_theResult___fst_sfd__h111340,
		_theResult___fst_sfd__h120089,
		_theResult___fst_sfd__h120092,
		_theResult___fst_sfd__h12359,
		_theResult___fst_sfd__h128701,
		_theResult___fst_sfd__h128704,
		_theResult___fst_sfd__h12912,
		_theResult___fst_sfd__h12915,
		_theResult___fst_sfd__h137942,
		_theResult___fst_sfd__h137945,
		_theResult___fst_sfd__h146608,
		_theResult___fst_sfd__h146611,
		_theResult___fst_sfd__h146620,
		_theResult___fst_sfd__h146626,
		_theResult___fst_sfd__h148525,
		_theResult___fst_sfd__h22977,
		_theResult___fst_sfd__h23529,
		_theResult___fst_sfd__h23532,
		_theResult___fst_sfd__h29405,
		_theResult___fst_sfd__h29958,
		_theResult___fst_sfd__h29961,
		_theResult___fst_sfd__h35575,
		_theResult___fst_sfd__h36127,
		_theResult___fst_sfd__h36130,
		_theResult___sfd__h119991,
		_theResult___sfd__h12262,
		_theResult___sfd__h12815,
		_theResult___sfd__h128603,
		_theResult___sfd__h137844,
		_theResult___sfd__h146510,
		_theResult___sfd__h22881,
		_theResult___sfd__h23433,
		_theResult___sfd__h29308,
		_theResult___sfd__h29861,
		_theResult___sfd__h35479,
		_theResult___sfd__h36031,
		_theResult___snd_fst_sfd__h103681,
		_theResult___snd_fst_sfd__h128707,
		_theResult___snd_fst_sfd__h12918,
		_theResult___snd_fst_sfd__h146614,
		_theResult___snd_fst_sfd__h23535,
		_theResult___snd_fst_sfd__h29964,
		_theResult___snd_fst_sfd__h36133,
		out_sfd__h119994,
		out_sfd__h12265,
		out_sfd__h12818,
		out_sfd__h128606,
		out_sfd__h137847,
		out_sfd__h146513,
		out_sfd__h22884,
		out_sfd__h23436,
		out_sfd__h29311,
		out_sfd__h29864,
		out_sfd__h35482,
		out_sfd__h36034,
		sV1_sfd__h824,
		sV2_sfd__h927,
		value__h148270;
  wire [19 : 0] NEG_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFF_ETC___d1682,
		NEG_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFF_ETC___d1714,
		NEG_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFF_ETC___d1715,
		NEG_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFF_ETC___d1778,
		NEG_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFF_ETC___d1863,
		NEG_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFF_ETC___d1864,
		NEG_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFF_ETC___d1922;
  wire [11 : 0] IF_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFFF_ETC___d4889,
		SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFF_ETC___d4566,
		SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFF_ETC__q150,
		SEXT_requestR_BITS_190_TO_180_599_MINUS_1023_611___d3734,
		SEXT_requestR_BITS_190_TO_180_599_MINUS_1023_6_ETC__q118,
		_3074_MINUS_0_CONCAT_IF_requestR_BIT_179_71_THE_ETC___d3303,
		_3074_MINUS_SEXT_IF_requestR_BITS_191_TO_160_4__ETC___d4569,
		_32_MINUS_0_CONCAT_IF_IF_requestR_BIT_159_6_THE_ETC___d2233,
		_32_MINUS_0_CONCAT_IF_requestR_BIT_159_6_THEN_0_ETC___d2448,
		_3970_MINUS_0_CONCAT_IF_IF_requestR_BITS_191_TO_ETC___d4423,
		_3970_MINUS_SEXT_requestR_BITS_190_TO_180_599_M_ETC___d3737,
		_64_MINUS_0_CONCAT_IF_IF_requestR_BIT_191_27_TH_ETC___d2769,
		_64_MINUS_0_CONCAT_IF_requestR_BIT_191_27_THEN__ETC___d2954,
		x__h129822,
		x__h171157,
		x__h61032,
		x__h70727,
		x__h84573,
		x__h95584;
  wire [10 : 0] IF_IF_IF_IF_3074_MINUS_SEXT_IF_requestR_BITS_1_ETC___d4874,
		IF_IF_IF_IF_3074_MINUS_SEXT_IF_requestR_BITS_1_ETC___d4876,
		IF_IF_IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFF_ETC___d4549,
		IF_IF_IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFF_ETC___d4551,
		IF_IF_IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFF_ETC___d4943,
		IF_IF_IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFF_ETC___d4945,
		IF_IF_IF_requestR_BIT_159_6_THEN_NEG_requestR__ETC___d2310,
		IF_IF_IF_requestR_BIT_159_6_THEN_NEG_requestR__ETC___d2336,
		IF_IF_IF_requestR_BIT_159_6_THEN_NEG_requestR__ETC___d2338,
		IF_IF_IF_requestR_BIT_191_27_THEN_NEG_requestR_ETC___d2845,
		IF_IF_IF_requestR_BIT_191_27_THEN_NEG_requestR_ETC___d2871,
		IF_IF_IF_requestR_BIT_191_27_THEN_NEG_requestR_ETC___d2873,
		IF_requestR_BITS_191_TO_128_24_EQ_0_25_OR_NOT__ETC___d2883,
		SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFF_ETC__q153,
		_theResult___exp__h169734,
		_theResult___exp__h179381,
		_theResult___exp__h188163,
		_theResult___exp__h60903,
		_theResult___exp__h61659,
		_theResult___exp__h70599,
		_theResult___exp__h71354,
		_theResult___exp__h84444,
		_theResult___exp__h85200,
		_theResult___exp__h95456,
		_theResult___exp__h96211,
		_theResult___fst_exp__h154006,
		_theResult___fst_exp__h169070,
		_theResult___fst_exp__h169076,
		_theResult___fst_exp__h169079,
		_theResult___fst_exp__h169832,
		_theResult___fst_exp__h169835,
		_theResult___fst_exp__h178652,
		_theResult___fst_exp__h178717,
		_theResult___fst_exp__h178723,
		_theResult___fst_exp__h178726,
		_theResult___fst_exp__h179479,
		_theResult___fst_exp__h179482,
		_theResult___fst_exp__h187435,
		_theResult___fst_exp__h187474,
		_theResult___fst_exp__h187480,
		_theResult___fst_exp__h187483,
		_theResult___fst_exp__h188261,
		_theResult___fst_exp__h188264,
		_theResult___fst_exp__h188273,
		_theResult___fst_exp__h188276,
		_theResult___fst_exp__h61000,
		_theResult___fst_exp__h61756,
		_theResult___fst_exp__h61759,
		_theResult___fst_exp__h70695,
		_theResult___fst_exp__h71450,
		_theResult___fst_exp__h71453,
		_theResult___fst_exp__h84541,
		_theResult___fst_exp__h85297,
		_theResult___fst_exp__h85300,
		_theResult___fst_exp__h95552,
		_theResult___fst_exp__h96307,
		_theResult___fst_exp__h96310,
		_theResult___snd_fst_exp__h169838,
		_theResult___snd_fst_exp__h188267,
		_theResult___snd_fst_exp__h61762,
		_theResult___snd_fst_exp__h61765,
		_theResult___snd_fst_exp__h61768,
		_theResult___snd_fst_exp__h71456,
		_theResult___snd_fst_exp__h71459,
		_theResult___snd_fst_exp__h71462,
		_theResult___snd_fst_exp__h85303,
		_theResult___snd_fst_exp__h85306,
		_theResult___snd_fst_exp__h85309,
		_theResult___snd_fst_exp__h96313,
		_theResult___snd_fst_exp__h96316,
		_theResult___snd_fst_exp__h96319,
		din_inc___2_exp__h188299,
		din_inc___2_exp__h188329,
		din_inc___2_exp__h188353,
		din_inc___2_exp__h61802,
		din_inc___2_exp__h71492,
		din_inc___2_exp__h85343,
		din_inc___2_exp__h96349,
		out_exp__h169737,
		out_exp__h179384,
		out_exp__h188166,
		out_exp__h60906,
		out_exp__h61662,
		out_exp__h70602,
		out_exp__h71357,
		out_exp__h84447,
		out_exp__h85203,
		out_exp__h95459,
		out_exp__h96214,
		requestR_BITS_190_TO_180_599_MINUS_1023___d2611,
		x__h148211;
  wire [8 : 0] IF_SEXT_requestR_BITS_190_TO_180_599_MINUS_102_ETC___d4055,
	       _32_MINUS_0_CONCAT_IF_IF_requestR_BIT_159_6_THE_ETC___d1255,
	       _32_MINUS_0_CONCAT_IF_requestR_BIT_159_6_THEN_0_ETC___d1510,
	       _64_MINUS_0_CONCAT_IF_IF_requestR_BIT_191_27_TH_ETC___d387,
	       _64_MINUS_0_CONCAT_IF_requestR_BIT_191_27_THEN__ETC___d904,
	       x__h12390,
	       x__h23008,
	       x__h29436,
	       x__h35606;
  wire [7 : 0] IF_IF_IF_IF_0b0_CONCAT_NOT_requestR_BITS_190_T_ETC___d3596,
	       IF_IF_IF_IF_0b0_CONCAT_NOT_requestR_BITS_190_T_ETC___d3598,
	       IF_IF_IF_IF_3970_MINUS_SEXT_requestR_BITS_190__ETC___d4040,
	       IF_IF_IF_IF_3970_MINUS_SEXT_requestR_BITS_190__ETC___d4042,
	       IF_IF_IF_requestR_BITS_190_TO_180_599_EQ_0_609_ETC___d3713,
	       IF_IF_IF_requestR_BITS_190_TO_180_599_EQ_0_609_ETC___d3715,
	       IF_IF_IF_requestR_BITS_190_TO_180_599_EQ_0_609_ETC___d4109,
	       IF_IF_IF_requestR_BITS_190_TO_180_599_EQ_0_609_ETC___d4111,
	       IF_IF_IF_requestR_BIT_159_6_THEN_NEG_requestR__ETC___d1335,
	       IF_IF_IF_requestR_BIT_159_6_THEN_NEG_requestR__ETC___d1361,
	       IF_IF_IF_requestR_BIT_159_6_THEN_NEG_requestR__ETC___d1363,
	       IF_IF_IF_requestR_BIT_191_27_THEN_NEG_requestR_ETC___d476,
	       IF_IF_IF_requestR_BIT_191_27_THEN_NEG_requestR_ETC___d502,
	       IF_IF_IF_requestR_BIT_191_27_THEN_NEG_requestR_ETC___d504,
	       IF_requestR_BITS_159_TO_128_121_EQ_0_122_OR_NO_ETC___d1373,
	       IF_requestR_BITS_159_TO_128_121_EQ_0_122_OR_NO_ETC___d1596,
	       IF_requestR_BITS_191_TO_128_24_EQ_0_25_OR_NOT__ETC___d514,
	       IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d1680,
	       SEXT_requestR_BITS_190_TO_180_599_MINUS_1023_6_ETC__q121,
	       _theResult___exp__h119990,
	       _theResult___exp__h12261,
	       _theResult___exp__h12814,
	       _theResult___exp__h128602,
	       _theResult___exp__h137843,
	       _theResult___exp__h146509,
	       _theResult___exp__h22880,
	       _theResult___exp__h23432,
	       _theResult___exp__h29307,
	       _theResult___exp__h29860,
	       _theResult___exp__h35478,
	       _theResult___exp__h36030,
	       _theResult___fst_exp__h111339,
	       _theResult___fst_exp__h119464,
	       _theResult___fst_exp__h119529,
	       _theResult___fst_exp__h119535,
	       _theResult___fst_exp__h119538,
	       _theResult___fst_exp__h120088,
	       _theResult___fst_exp__h120091,
	       _theResult___fst_exp__h12358,
	       _theResult___fst_exp__h128141,
	       _theResult___fst_exp__h128147,
	       _theResult___fst_exp__h128150,
	       _theResult___fst_exp__h128700,
	       _theResult___fst_exp__h128703,
	       _theResult___fst_exp__h12911,
	       _theResult___fst_exp__h12914,
	       _theResult___fst_exp__h137317,
	       _theResult___fst_exp__h137382,
	       _theResult___fst_exp__h137388,
	       _theResult___fst_exp__h137391,
	       _theResult___fst_exp__h137941,
	       _theResult___fst_exp__h137944,
	       _theResult___fst_exp__h145984,
	       _theResult___fst_exp__h146023,
	       _theResult___fst_exp__h146029,
	       _theResult___fst_exp__h146032,
	       _theResult___fst_exp__h146607,
	       _theResult___fst_exp__h146610,
	       _theResult___fst_exp__h146619,
	       _theResult___fst_exp__h146622,
	       _theResult___fst_exp__h22976,
	       _theResult___fst_exp__h23528,
	       _theResult___fst_exp__h23531,
	       _theResult___fst_exp__h29404,
	       _theResult___fst_exp__h29957,
	       _theResult___fst_exp__h29960,
	       _theResult___fst_exp__h35574,
	       _theResult___fst_exp__h36126,
	       _theResult___fst_exp__h36129,
	       _theResult___snd_fst_exp__h128706,
	       _theResult___snd_fst_exp__h12917,
	       _theResult___snd_fst_exp__h12920,
	       _theResult___snd_fst_exp__h12923,
	       _theResult___snd_fst_exp__h146613,
	       _theResult___snd_fst_exp__h23534,
	       _theResult___snd_fst_exp__h23537,
	       _theResult___snd_fst_exp__h23540,
	       _theResult___snd_fst_exp__h29963,
	       _theResult___snd_fst_exp__h29966,
	       _theResult___snd_fst_exp__h29969,
	       _theResult___snd_fst_exp__h36132,
	       _theResult___snd_fst_exp__h36135,
	       _theResult___snd_fst_exp__h36138,
	       din_inc___2_exp__h12957,
	       din_inc___2_exp__h146641,
	       din_inc___2_exp__h146665,
	       din_inc___2_exp__h146695,
	       din_inc___2_exp__h146719,
	       din_inc___2_exp__h23570,
	       din_inc___2_exp__h30003,
	       din_inc___2_exp__h36168,
	       out_exp__h119993,
	       out_exp__h12264,
	       out_exp__h12817,
	       out_exp__h128605,
	       out_exp__h137846,
	       out_exp__h146512,
	       out_exp__h22883,
	       out_exp__h23435,
	       out_exp__h29310,
	       out_exp__h29863,
	       out_exp__h35481,
	       out_exp__h36033,
	       sV1_exp__h823,
	       sV2_exp__h926,
	       x__h99506;
  wire [6 : 0] IF_IF_requestR_BIT_191_27_THEN_NEG_requestR_BI_ETC___d384,
	       IF_requestR_BIT_191_27_THEN_0_ELSE_IF_requestR_ETC___d901;
  wire [5 : 0] IF_IF_0b0_CONCAT_NOT_requestR_BITS_190_TO_180__ETC___d3537,
	       IF_IF_3074_MINUS_SEXT_IF_requestR_BITS_191_TO__ETC___d4815,
	       IF_IF_3970_MINUS_SEXT_requestR_BITS_190_TO_180_ETC___d3981,
	       IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_ETC___d4495,
	       IF_IF_requestR_BIT_159_6_THEN_NEG_requestR_BIT_ETC___d1252,
	       IF_IF_requestR_BIT_159_6_THEN_NEG_requestR_BIT_ETC___d2230,
	       IF_requestR_BITS_190_TO_180_599_EQ_0_609_THEN__ETC___d3659,
	       IF_requestR_BIT_159_6_THEN_0_ELSE_IF_requestR__ETC___d1507,
	       IF_requestR_BIT_159_6_THEN_0_ELSE_IF_requestR__ETC___d2445;
  wire [4 : 0] _0_CONCAT_IF_IF_0b0_CONCAT_NOT_requestR_BITS_19_ETC___d4279,
	       _0_CONCAT_IF_IF_3074_MINUS_SEXT_IF_requestR_BIT_ETC___d5102,
	       _0_CONCAT_IF_IF_3970_MINUS_SEXT_requestR_BITS_1_ETC___d4308,
	       _0_CONCAT_IF_IF_requestR_BITS_191_TO_160_4_EQ_0_ETC___d5085,
	       _0_CONCAT_IF_requestR_BITS_190_TO_180_599_EQ_0__ETC___d4291,
	       x__h13083,
	       x__h147219,
	       x__h189005,
	       x__h193477,
	       x__h203311,
	       x__h23674,
	       x__h30129,
	       x__h36272,
	       x__h38337,
	       x__h39093,
	       x__h40655,
	       x__h41414,
	       x__h43701,
	       x__h49451,
	       x__h61924,
	       x__h71592,
	       x__h73195,
	       x__h73954,
	       x__h85465,
	       x__h96449,
	       x__h98497,
	       x__h99253;
  wire [1 : 0] IF_sfd___30277_BIT_1_THEN_2_ELSE_0__q68,
	       IF_sfd___30277_BIT_2_THEN_2_ELSE_0__q67,
	       IF_sfd___31835_BIT_10_THEN_2_ELSE_0__q9,
	       IF_sfd___31835_BIT_11_THEN_2_ELSE_0__q8,
	       IF_sfd___31835_BIT_39_THEN_2_ELSE_0__q7,
	       IF_sfd___31835_BIT_40_THEN_2_ELSE_0__q6,
	       IF_sfd___32457_BIT_10_THEN_2_ELSE_0__q25,
	       IF_sfd___32457_BIT_11_THEN_2_ELSE_0__q24,
	       IF_sfd___32457_BIT_39_THEN_2_ELSE_0__q23,
	       IF_sfd___32457_BIT_40_THEN_2_ELSE_0__q22,
	       IF_sfd___35055_BIT_7_THEN_2_ELSE_0__q53,
	       IF_sfd___35055_BIT_8_THEN_2_ELSE_0__q52,
	       IF_sfd___38884_BIT_7_THEN_2_ELSE_0__q39,
	       IF_sfd___38884_BIT_8_THEN_2_ELSE_0__q38,
	       IF_sfd___39973_BIT_1_THEN_2_ELSE_0__q82,
	       IF_sfd___39973_BIT_2_THEN_2_ELSE_0__q81,
	       IF_sfdin19458_BIT_33_THEN_2_ELSE_0__q115,
	       IF_sfdin37311_BIT_33_THEN_2_ELSE_0__q120,
	       IF_sfdin78646_BIT_4_THEN_2_ELSE_0__q152,
	       IF_theResult___snd28101_BIT_33_THEN_2_ELSE_0__q117,
	       IF_theResult___snd45978_BIT_33_THEN_2_ELSE_0__q123,
	       IF_theResult___snd69030_BIT_4_THEN_2_ELSE_0__q149,
	       IF_theResult___snd87429_BIT_4_THEN_2_ELSE_0__q155,
	       IF_x0258_BIT_24_THEN_2_ELSE_0__q65,
	       IF_x1336_BIT_24_THEN_2_ELSE_0__q66,
	       IF_x2798_BIT_53_THEN_2_ELSE_0__q92,
	       IF_x3876_BIT_53_THEN_2_ELSE_0__q93,
	       IF_x7699_BIT_24_THEN_2_ELSE_0__q63,
	       IF_x7876_BIT_53_THEN_2_ELSE_0__q112,
	       IF_x9015_BIT_24_THEN_2_ELSE_0__q64,
	       IF_x9175_BIT_53_THEN_2_ELSE_0__q113,
	       guard__h111367,
	       guard__h11845,
	       guard__h120102,
	       guard__h12375,
	       guard__h129091,
	       guard__h137955,
	       guard__h161118,
	       guard__h170426,
	       guard__h179493,
	       guard__h22467,
	       guard__h22993,
	       guard__h28894,
	       guard__h29421,
	       guard__h35065,
	       guard__h35591,
	       guard__h36732,
	       guard__h37510,
	       guard__h38794,
	       guard__h39515,
	       guard__h40069,
	       guard__h41115,
	       guard__h60287,
	       guard__h61017,
	       guard__h69983,
	       guard__h70712,
	       guard__h72055,
	       guard__h72609,
	       guard__h73655,
	       guard__h83828,
	       guard__h84558,
	       guard__h94840,
	       guard__h95569,
	       guard__h96909,
	       guard__h97687,
	       guard__h98954;
  wire IF_3074_MINUS_0_CONCAT_IF_requestR_BIT_179_71__ETC___d4241,
       IF_32_MINUS_0_CONCAT_IF_IF_requestR_BIT_159_6__ETC___d1313,
       IF_32_MINUS_0_CONCAT_IF_IF_requestR_BIT_159_6__ETC___d1463,
       IF_32_MINUS_0_CONCAT_IF_IF_requestR_BIT_159_6__ETC___d2289,
       IF_32_MINUS_0_CONCAT_IF_IF_requestR_BIT_159_6__ETC___d2404,
       IF_32_MINUS_0_CONCAT_IF_requestR_BIT_159_6_THE_ETC___d1651,
       IF_32_MINUS_0_CONCAT_IF_requestR_BIT_159_6_THE_ETC___d2587,
       IF_64_MINUS_0_CONCAT_IF_IF_requestR_BIT_191_27_ETC___d2824,
       IF_64_MINUS_0_CONCAT_IF_IF_requestR_BIT_191_27_ETC___d2941,
       IF_64_MINUS_0_CONCAT_IF_IF_requestR_BIT_191_27_ETC___d454,
       IF_64_MINUS_0_CONCAT_IF_IF_requestR_BIT_191_27_ETC___d636,
       IF_64_MINUS_0_CONCAT_IF_requestR_BIT_191_27_TH_ETC___d1109,
       IF_64_MINUS_0_CONCAT_IF_requestR_BIT_191_27_TH_ETC___d3094,
       IF_IF_IF_3074_MINUS_SEXT_IF_requestR_BITS_191__ETC___d5059,
       IF_IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFF_ETC___d5067,
       IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_ETC___d5071,
       IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_ETC___d5106,
       IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_ETC___d5109,
       IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_ETC___d5116,
       IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_ETC___d5130,
       IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_ETC___d5142,
       IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_ETC___d5154,
       IF_NEG_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0_ETC___d1769,
       IF_NEG_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0_ETC___d1913,
       IF_NEG_SEXT_requestR_BITS_190_TO_180_599_MINUS_ETC___d2701,
       IF_NEG_SEXT_requestR_BITS_190_TO_180_599_MINUS_ETC___d3183,
       IF_NOT_32_MINUS_0_CONCAT_IF_IF_requestR_BIT_15_ETC___d2290,
       IF_NOT_3970_MINUS_0_CONCAT_IF_IF_requestR_BITS_ETC___d5051,
       IF_NOT_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFF_ETC___d2029,
       IF_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFFF_ETC___d5069,
       IF_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFFF_ETC___d5128,
       IF_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFFF_ETC___d5140,
       IF_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFFF_ETC___d5152,
       IF_SEXT_requestR_BITS_190_TO_180_599_MINUS_102_ETC___d4259,
       IF_SEXT_requestR_BITS_190_TO_180_599_MINUS_102_ETC___d4337,
       IF_SEXT_requestR_BITS_190_TO_180_599_MINUS_102_ETC___d4350,
       IF_SEXT_requestR_BITS_190_TO_180_599_MINUS_102_ETC___d4363,
       IF_requestR_BITS_127_TO_96_2_EQ_0xFFFFFFFF_3_T_ETC___d2009,
       IF_requestR_BITS_190_TO_180_599_EQ_0_609_THEN__ETC___d4261,
       IF_requestR_BITS_190_TO_180_599_EQ_0_609_THEN__ETC___d4312,
       IF_requestR_BITS_190_TO_180_599_EQ_0_609_THEN__ETC___d4323,
       IF_requestR_BITS_190_TO_180_599_EQ_0_609_THEN__ETC___d4339,
       IF_requestR_BITS_190_TO_180_599_EQ_0_609_THEN__ETC___d4352,
       IF_requestR_BITS_190_TO_180_599_EQ_0_609_THEN__ETC___d4365,
       IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d1676,
       IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d1815,
       IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d1827,
       IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d1828,
       IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d1960,
       IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d1972,
       IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d1973,
       IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d1995,
       IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d2005,
       IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d2018,
       IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d2019,
       IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d2020,
       IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d2023,
       IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d2025,
       IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d2043,
       IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d2080,
       IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d2091,
       IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d2095,
       IF_requestR_BITS_194_TO_192_0_EQ_0x0_1_OR_NOT__ETC___d1706,
       IF_requestR_BITS_194_TO_192_0_EQ_0x0_1_OR_NOT__ETC___d1738,
       IF_requestR_BITS_194_TO_192_0_EQ_0x0_1_OR_NOT__ETC___d1799,
       IF_requestR_BITS_194_TO_192_0_EQ_0x0_1_OR_NOT__ETC___d1855,
       IF_requestR_BITS_194_TO_192_0_EQ_0x0_1_OR_NOT__ETC___d1887,
       IF_requestR_BITS_194_TO_192_0_EQ_0x0_1_OR_NOT__ETC___d1943,
       IF_requestR_BITS_194_TO_192_0_EQ_0x0_1_OR_NOT__ETC___d2637,
       IF_requestR_BITS_194_TO_192_0_EQ_0x0_1_OR_NOT__ETC___d2669,
       IF_requestR_BITS_194_TO_192_0_EQ_0x0_1_OR_NOT__ETC___d2731,
       IF_requestR_BITS_194_TO_192_0_EQ_0x0_1_OR_NOT__ETC___d3126,
       IF_requestR_BITS_194_TO_192_0_EQ_0x0_1_OR_NOT__ETC___d3158,
       IF_requestR_BITS_194_TO_192_0_EQ_0x0_1_OR_NOT__ETC___d3213,
       IF_requestR_BIT_159_6_THEN_NEG_requestR_BITS_1_ETC___d1454,
       IF_requestR_BIT_159_6_THEN_NEG_requestR_BITS_1_ETC___d1457,
       IF_requestR_BIT_159_6_THEN_NEG_requestR_BITS_1_ETC___d1466,
       IF_requestR_BIT_191_27_THEN_NEG_requestR_BITS__ETC___d2932,
       IF_requestR_BIT_191_27_THEN_NEG_requestR_BITS__ETC___d2935,
       IF_requestR_BIT_191_27_THEN_NEG_requestR_BITS__ETC___d2944,
       IF_requestR_BIT_191_27_THEN_NEG_requestR_BITS__ETC___d627,
       IF_requestR_BIT_191_27_THEN_NEG_requestR_BITS__ETC___d630,
       IF_requestR_BIT_191_27_THEN_NEG_requestR_BITS__ETC___d639,
       IF_requestR_BIT_191_27_THEN_NOT_requestR_BITS__ETC___d5207,
       NEG_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFF_ETC___d1717,
       NEG_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFF_ETC___d1780,
       NEG_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFF_ETC___d1866,
       NEG_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFF_ETC___d1924,
       NEG_SEXT_requestR_BITS_190_TO_180_599_MINUS_10_ETC___d2648,
       NEG_SEXT_requestR_BITS_190_TO_180_599_MINUS_10_ETC___d2712,
       NEG_SEXT_requestR_BITS_190_TO_180_599_MINUS_10_ETC___d3137,
       NEG_SEXT_requestR_BITS_190_TO_180_599_MINUS_10_ETC___d3194,
       NOT_3074_MINUS_0_CONCAT_IF_requestR_BIT_179_71_ETC___d4331,
       NOT_3074_MINUS_0_CONCAT_IF_requestR_BIT_179_71_ETC___d4359,
       NOT_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFF_ETC___d1758,
       NOT_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFF_ETC___d1821,
       NOT_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFF_ETC___d1905,
       NOT_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFF_ETC___d1966,
       NOT_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFF_ETC___d2032,
       NOT_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFF_ETC___d2033,
       NOT_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFF_ETC___d2090,
       NOT_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFF_ETC___d2096,
       NOT_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFF_ETC___d2114,
       NOT_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFF_ETC___d4468,
       NOT_IF_requestR_BIT_159_6_THEN_NEG_requestR_BI_ETC___d1260,
       NOT_IF_requestR_BIT_191_27_THEN_NEG_requestR_B_ETC___d2774,
       NOT_IF_requestR_BIT_191_27_THEN_NEG_requestR_B_ETC___d392,
       NOT_requestR_BITS_159_TO_128_121_EQ_0_122_123__ETC___d1643,
       NOT_requestR_BITS_190_TO_180_599_EQ_0_609_615__ETC___d2690,
       NOT_requestR_BITS_190_TO_180_599_EQ_0_609_615__ETC___d2754,
       NOT_requestR_BITS_190_TO_180_599_EQ_0_609_615__ETC___d3175,
       NOT_requestR_BITS_190_TO_180_599_EQ_0_609_615__ETC___d3235,
       NOT_requestR_BITS_190_TO_180_599_EQ_2047_600_6_ETC___d5211,
       NOT_requestR_BITS_190_TO_180_599_EQ_2047_600_6_ETC___d5276,
       NOT_requestR_BITS_190_TO_180_599_ULT_requestR__ETC___d5253,
       NOT_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5_ETC___d2094,
       NOT_requestR_BIT_158_12_13_AND_NOT_requestR_BI_ETC___d803,
       NOT_requestR_BIT_179_71_72_AND_NOT_requestR_BI_ETC___d824,
       NOT_requestR_BIT_191_27_48_AND_NOT_requestR_BI_ETC___d3042,
       NOT_requestR_BIT_191_27_48_AND_NOT_requestR_BI_ETC___d994,
       SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFF_ETC___d4567,
       SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFF_ETC___d4568,
       SEXT_requestR_BITS_190_TO_180_599_MINUS_1023_6_ETC___d3735,
       SEXT_requestR_BITS_190_TO_180_599_MINUS_1023_6_ETC___d3736,
       _0_CONCAT_IF_IF_0b0_CONCAT_NOT_requestR_BITS_19_ETC___d3539,
       _0_CONCAT_IF_IF_3074_MINUS_SEXT_IF_requestR_BIT_ETC___d4817,
       _0_CONCAT_IF_IF_3970_MINUS_SEXT_requestR_BITS_1_ETC___d3983,
       _0_CONCAT_IF_IF_requestR_BITS_191_TO_160_4_EQ_0_ETC___d4497,
       _0_CONCAT_IF_IF_requestR_BITS_191_TO_160_4_EQ_0_ETC___d4890,
       _0_CONCAT_IF_requestR_BITS_190_TO_180_599_EQ_0__ETC___d3661,
       _0_CONCAT_IF_requestR_BITS_190_TO_180_599_EQ_0__ETC___d4056,
       _3074_MINUS_0_CONCAT_IF_requestR_BIT_179_71_THE_ETC___d3304,
       _3074_MINUS_0_CONCAT_IF_requestR_BIT_179_71_THE_ETC___d3305,
       _3074_MINUS_0_CONCAT_IF_requestR_BIT_179_71_THE_ETC___d4294,
       _3074_MINUS_0_CONCAT_IF_requestR_BIT_179_71_THE_ETC___d4319,
       _3074_MINUS_0_CONCAT_IF_requestR_BIT_179_71_THE_ETC___d4346,
       _32_MINUS_0_CONCAT_IF_IF_requestR_BIT_159_6_THE_ETC___d1256,
       _32_MINUS_0_CONCAT_IF_IF_requestR_BIT_159_6_THE_ETC___d1258,
       _32_MINUS_0_CONCAT_IF_IF_requestR_BIT_159_6_THE_ETC___d1261,
       _32_MINUS_0_CONCAT_IF_IF_requestR_BIT_159_6_THE_ETC___d2234,
       _32_MINUS_0_CONCAT_IF_IF_requestR_BIT_159_6_THE_ETC___d2236,
       _32_MINUS_0_CONCAT_IF_IF_requestR_BIT_159_6_THE_ETC___d2238,
       _32_MINUS_0_CONCAT_IF_requestR_BIT_159_6_THEN_0_ETC___d1511,
       _32_MINUS_0_CONCAT_IF_requestR_BIT_159_6_THEN_0_ETC___d1512,
       _32_MINUS_0_CONCAT_IF_requestR_BIT_159_6_THEN_0_ETC___d1513,
       _32_MINUS_0_CONCAT_IF_requestR_BIT_159_6_THEN_0_ETC___d2449,
       _32_MINUS_0_CONCAT_IF_requestR_BIT_159_6_THEN_0_ETC___d2450,
       _32_MINUS_0_CONCAT_IF_requestR_BIT_159_6_THEN_0_ETC___d2451,
       _3970_MINUS_0_CONCAT_IF_IF_requestR_BITS_191_TO_ETC___d4424,
       _3970_MINUS_0_CONCAT_IF_IF_requestR_BITS_191_TO_ETC___d4425,
       _64_MINUS_0_CONCAT_IF_IF_requestR_BIT_191_27_TH_ETC___d2770,
       _64_MINUS_0_CONCAT_IF_IF_requestR_BIT_191_27_TH_ETC___d2772,
       _64_MINUS_0_CONCAT_IF_IF_requestR_BIT_191_27_TH_ETC___d2775,
       _64_MINUS_0_CONCAT_IF_IF_requestR_BIT_191_27_TH_ETC___d388,
       _64_MINUS_0_CONCAT_IF_IF_requestR_BIT_191_27_TH_ETC___d390,
       _64_MINUS_0_CONCAT_IF_IF_requestR_BIT_191_27_TH_ETC___d393,
       _64_MINUS_0_CONCAT_IF_requestR_BIT_191_27_THEN__ETC___d2955,
       _64_MINUS_0_CONCAT_IF_requestR_BIT_191_27_THEN__ETC___d2956,
       _64_MINUS_0_CONCAT_IF_requestR_BIT_191_27_THEN__ETC___d2957,
       _64_MINUS_0_CONCAT_IF_requestR_BIT_191_27_THEN__ETC___d905,
       _64_MINUS_0_CONCAT_IF_requestR_BIT_191_27_THEN__ETC___d906,
       _64_MINUS_0_CONCAT_IF_requestR_BIT_191_27_THEN__ETC___d907,
       guard__h129689,
       guard__h171024,
       requestR_BITS_126_TO_116_166_EQ_0_180_AND_requ_ETC___d5187,
       requestR_BITS_179_TO_128_601_ULE_requestR_BITS_ETC___d5199,
       requestR_BITS_179_TO_128_601_ULT_requestR_BITS_ETC___d5204,
       requestR_BITS_190_TO_180_599_EQ_0_609_AND_requ_ETC___d5183,
       requestR_BITS_190_TO_180_599_EQ_0_609_AND_requ_ETC___d5257,
       requestR_BITS_190_TO_180_599_EQ_2047_600_AND_0_ETC___d2749,
       requestR_BITS_190_TO_180_599_EQ_2047_600_AND_0_ETC___d2760,
       requestR_BITS_190_TO_180_599_EQ_2047_600_AND_0_ETC___d3230,
       requestR_BITS_190_TO_180_599_EQ_2047_600_AND_0_ETC___d3241,
       requestR_BITS_190_TO_180_599_EQ_2047_600_AND_N_ETC___d5175,
       requestR_BITS_190_TO_180_599_EQ_2047_600_AND_N_ETC___d5220,
       requestR_BITS_190_TO_180_599_EQ_2047_600_AND_N_ETC___d5242,
       requestR_BITS_190_TO_180_599_EQ_requestR_BITS__ETC___d5198,
       requestR_BITS_190_TO_180_599_ULE_requestR_BITS_ETC___d5196,
       requestR_BITS_190_TO_180_599_ULE_requestR_BITS_ETC___d5252,
       requestR_BITS_190_TO_180_599_ULT_requestR_BITS_ETC___d5203,
       requestR_BITS_191_TO_128_24_EQ_0_25_OR_NOT_req_ETC___d837,
       requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5_AND_ETC___d2031,
       requestR_BIT_158_12_OR_requestR_BIT_157_14_OR__ETC___d1058,
       requestR_BIT_159_6_OR_requestR_BIT_158_12_OR_r_ETC___d1654,
       requestR_BIT_179_71_OR_requestR_BIT_178_73_OR__ETC___d1079,
       requestR_BIT_191_27_OR_requestR_BIT_190_49_OR__ETC___d1100,
       requestR_BIT_191_27_OR_requestR_BIT_190_49_OR__ETC___d1103,
       requestR_BIT_191_27_OR_requestR_BIT_190_49_OR__ETC___d1112,
       requestR_BIT_191_27_OR_requestR_BIT_190_49_OR__ETC___d3085,
       requestR_BIT_191_27_OR_requestR_BIT_190_49_OR__ETC___d3088,
       requestR_BIT_191_27_OR_requestR_BIT_190_49_OR__ETC___d3097,
       value_BIT_23___h161776;
  // action method set_verbosity
  assign RDY_set_verbosity = 1'd1 ;
  assign CAN_FIRE_set_verbosity = 1'd1 ;
  assign WILL_FIRE_set_verbosity = EN_set_verbosity ;
  // action method req
  assign CAN_FIRE_req = 1'd1 ;
  assign WILL_FIRE_req = EN_req ;
  // value method valid
  assign valid = dw_valid$whas && dw_valid$wget ;
  // value method word_fst
  assign word_fst = ab__h206728[68:5] ;
  // value method word_snd
  assign word_snd = ab__h206728[4:0] ;
  // submodule fpu
  mkFPU fpu(.CLK(CLK),
	    .RST_N(RST_N),
	    .request_put(fpu$request_put),
	    .EN_request_put(fpu$EN_request_put),
	    .EN_response_get(fpu$EN_response_get),
	    .RDY_request_put(fpu$RDY_request_put),
	    .response_get(fpu$response_get),
	    .RDY_response_get(fpu$RDY_response_get));
  // submodule frmFpuF
  FIFO2 #(.width(32'd1), .guarded(32'd1)) frmFpuF(.RST(RST_N),
						  .CLK(CLK),
						  .D_IN(frmFpuF$D_IN),
						  .ENQ(frmFpuF$ENQ),
						  .DEQ(frmFpuF$DEQ),
						  .CLR(frmFpuF$CLR),
						  .D_OUT(),
						  .FULL_N(),
						  .EMPTY_N());
  // rule RL_doFADD_S
  assign CAN_FIRE_RL_doFADD_S =
	     fpu$RDY_request_put && requestR[214] && stateR == 2'd0 &&
	     requestR[213:207] == 7'b1010011 &&
	     requestR[206:200] == 7'h0 ;
  assign WILL_FIRE_RL_doFADD_S = CAN_FIRE_RL_doFADD_S ;
  // rule RL_doFSUB_S
  assign CAN_FIRE_RL_doFSUB_S =
	     fpu$RDY_request_put && requestR[214] && stateR == 2'd0 &&
	     requestR[213:207] == 7'b1010011 &&
	     requestR[206:200] == 7'h04 ;
  assign WILL_FIRE_RL_doFSUB_S = CAN_FIRE_RL_doFSUB_S ;
  // rule RL_doFMUL_S
  assign CAN_FIRE_RL_doFMUL_S =
	     fpu$RDY_request_put && requestR[214] && stateR == 2'd0 &&
	     requestR[213:207] == 7'b1010011 &&
	     requestR[206:200] == 7'h08 ;
  assign WILL_FIRE_RL_doFMUL_S = CAN_FIRE_RL_doFMUL_S ;
  // rule RL_doFMADD_S
  assign CAN_FIRE_RL_doFMADD_S =
	     fpu$RDY_request_put && requestR[214] && stateR == 2'd0 &&
	     requestR[213:207] == 7'b1000011 &&
	     requestR[201:200] == 2'd0 ;
  assign WILL_FIRE_RL_doFMADD_S = CAN_FIRE_RL_doFMADD_S ;
  // rule RL_doFMSUB_S
  assign CAN_FIRE_RL_doFMSUB_S =
	     fpu$RDY_request_put && requestR[214] && stateR == 2'd0 &&
	     requestR[213:207] == 7'b1000111 &&
	     requestR[201:200] == 2'd0 ;
  assign WILL_FIRE_RL_doFMSUB_S = CAN_FIRE_RL_doFMSUB_S ;
  // rule RL_doFNMADD_S
  assign CAN_FIRE_RL_doFNMADD_S =
	     fpu$RDY_request_put && requestR[214] && stateR == 2'd0 &&
	     requestR[213:207] == 7'b1001111 &&
	     requestR[201:200] == 2'd0 ;
  assign WILL_FIRE_RL_doFNMADD_S = CAN_FIRE_RL_doFNMADD_S ;
  // rule RL_doFNMSUB_S
  assign CAN_FIRE_RL_doFNMSUB_S =
	     fpu$RDY_request_put && requestR[214] && stateR == 2'd0 &&
	     requestR[213:207] == 7'b1001011 &&
	     requestR[201:200] == 2'd0 ;
  assign WILL_FIRE_RL_doFNMSUB_S = CAN_FIRE_RL_doFNMSUB_S ;
  // rule RL_doFSGNJ_S
  assign CAN_FIRE_RL_doFSGNJ_S = MUX_dw_result$wset_1__SEL_2 ;
  assign WILL_FIRE_RL_doFSGNJ_S = MUX_dw_result$wset_1__SEL_2 ;
  // rule RL_doFSGNJN_S
  assign CAN_FIRE_RL_doFSGNJN_S = MUX_dw_result$wset_1__SEL_1 ;
  assign WILL_FIRE_RL_doFSGNJN_S = MUX_dw_result$wset_1__SEL_1 ;
  // rule RL_doFSGNJX_S
  assign CAN_FIRE_RL_doFSGNJX_S =
	     requestR[214] && stateR == 2'd0 &&
	     requestR[213:207] == 7'b1010011 &&
	     requestR[206:200] == 7'h10 &&
	     requestR[194:192] == 3'h2 ;
  assign WILL_FIRE_RL_doFSGNJX_S = CAN_FIRE_RL_doFSGNJX_S ;
  // rule RL_doFCVT_S_L
  assign CAN_FIRE_RL_doFCVT_S_L =
	     requestR[214] && stateR == 2'd0 &&
	     requestR[213:207] == 7'b1010011 &&
	     requestR[206:200] == 7'h68 &&
	     requestR[199:195] == 5'd2 ;
  assign WILL_FIRE_RL_doFCVT_S_L = CAN_FIRE_RL_doFCVT_S_L ;
  // rule RL_doFCVT_S_LU
  assign CAN_FIRE_RL_doFCVT_S_LU =
	     requestR[214] && stateR == 2'd0 &&
	     requestR[213:207] == 7'b1010011 &&
	     requestR[206:200] == 7'h68 &&
	     requestR[199:195] == 5'd3 ;
  assign WILL_FIRE_RL_doFCVT_S_LU = CAN_FIRE_RL_doFCVT_S_LU ;
  // rule RL_doFCVT_S_W
  assign CAN_FIRE_RL_doFCVT_S_W =
	     requestR[214] && stateR == 2'd0 &&
	     requestR[213:207] == 7'b1010011 &&
	     requestR[206:200] == 7'h68 &&
	     requestR[199:195] == 5'd0 ;
  assign WILL_FIRE_RL_doFCVT_S_W = CAN_FIRE_RL_doFCVT_S_W ;
  // rule RL_doFCVT_S_WU
  assign CAN_FIRE_RL_doFCVT_S_WU =
	     requestR[214] && stateR == 2'd0 &&
	     requestR[213:207] == 7'b1010011 &&
	     requestR[206:200] == 7'h68 &&
	     requestR[199:195] == 5'd1 ;
  assign WILL_FIRE_RL_doFCVT_S_WU = CAN_FIRE_RL_doFCVT_S_WU ;
  // rule RL_doFCVT_L_S
  assign CAN_FIRE_RL_doFCVT_L_S =
	     requestR[214] && stateR == 2'd0 &&
	     requestR[213:207] == 7'b1010011 &&
	     requestR[206:200] == 7'h60 &&
	     requestR[199:195] == 5'd2 ;
  assign WILL_FIRE_RL_doFCVT_L_S = CAN_FIRE_RL_doFCVT_L_S ;
  // rule RL_doFCVT_LU_S
  assign CAN_FIRE_RL_doFCVT_LU_S =
	     requestR[214] && stateR == 2'd0 &&
	     requestR[213:207] == 7'b1010011 &&
	     requestR[206:200] == 7'h60 &&
	     requestR[199:195] == 5'd3 ;
  assign WILL_FIRE_RL_doFCVT_LU_S = CAN_FIRE_RL_doFCVT_LU_S ;
  // rule RL_doFCVT_W_S
  assign CAN_FIRE_RL_doFCVT_W_S =
	     requestR[214] && stateR == 2'd0 &&
	     requestR[213:207] == 7'b1010011 &&
	     requestR[206:200] == 7'h60 &&
	     requestR[199:195] == 5'd0 ;
  assign WILL_FIRE_RL_doFCVT_W_S = CAN_FIRE_RL_doFCVT_W_S ;
  // rule RL_doFCVT_WU_S
  assign CAN_FIRE_RL_doFCVT_WU_S =
	     requestR[214] && stateR == 2'd0 &&
	     requestR[213:207] == 7'b1010011 &&
	     requestR[206:200] == 7'h60 &&
	     requestR[199:195] == 5'd1 ;
  assign WILL_FIRE_RL_doFCVT_WU_S = CAN_FIRE_RL_doFCVT_WU_S ;
  // rule RL_doFMIN_S
  assign CAN_FIRE_RL_doFMIN_S =
	     requestR[214] && stateR == 2'd0 &&
	     requestR[213:207] == 7'b1010011 &&
	     requestR[206:200] == 7'h14 &&
	     requestR[194:192] == 3'h0 ;
  assign WILL_FIRE_RL_doFMIN_S = CAN_FIRE_RL_doFMIN_S ;
  // rule RL_doFMAX_S
  assign CAN_FIRE_RL_doFMAX_S =
	     requestR[214] && stateR == 2'd0 &&
	     requestR[213:207] == 7'b1010011 &&
	     requestR[206:200] == 7'h14 &&
	     requestR[194:192] == 3'h1 ;
  assign WILL_FIRE_RL_doFMAX_S = CAN_FIRE_RL_doFMAX_S ;
  // rule RL_doFMV_W_X
  assign CAN_FIRE_RL_doFMV_W_X =
	     requestR[214] && stateR == 2'd0 &&
	     requestR[213:207] == 7'b1010011 &&
	     requestR[206:200] == 7'h78 &&
	     requestR[194:192] == 3'h0 ;
  assign WILL_FIRE_RL_doFMV_W_X = CAN_FIRE_RL_doFMV_W_X ;
  // rule RL_doFMV_X_W
  assign CAN_FIRE_RL_doFMV_X_W =
	     requestR[214] && stateR == 2'd0 &&
	     requestR[213:207] == 7'b1010011 &&
	     requestR[206:200] == 7'h70 &&
	     requestR[194:192] == 3'h0 ;
  assign WILL_FIRE_RL_doFMV_X_W = CAN_FIRE_RL_doFMV_X_W ;
  // rule RL_doFEQ_S
  assign CAN_FIRE_RL_doFEQ_S =
	     requestR[214] && stateR == 2'd0 &&
	     requestR[213:207] == 7'b1010011 &&
	     requestR[206:200] == 7'h50 &&
	     requestR[194:192] == 3'h2 ;
  assign WILL_FIRE_RL_doFEQ_S = CAN_FIRE_RL_doFEQ_S ;
  // rule RL_doFLT_S
  assign CAN_FIRE_RL_doFLT_S =
	     requestR[214] && stateR == 2'd0 &&
	     requestR[213:207] == 7'b1010011 &&
	     requestR[206:200] == 7'h50 &&
	     requestR[194:192] == 3'h1 ;
  assign WILL_FIRE_RL_doFLT_S = CAN_FIRE_RL_doFLT_S ;
  // rule RL_doFLE_S
  assign CAN_FIRE_RL_doFLE_S =
	     requestR[214] && stateR == 2'd0 &&
	     requestR[213:207] == 7'b1010011 &&
	     requestR[206:200] == 7'h50 &&
	     requestR[194:192] == 3'h0 ;
  assign WILL_FIRE_RL_doFLE_S = CAN_FIRE_RL_doFLE_S ;
  // rule RL_doFCLASS_S
  assign CAN_FIRE_RL_doFCLASS_S =
	     requestR[214] && stateR == 2'd0 &&
	     requestR[213:207] == 7'b1010011 &&
	     requestR[206:200] == 7'h70 &&
	     requestR[194:192] == 3'h1 ;
  assign WILL_FIRE_RL_doFCLASS_S = CAN_FIRE_RL_doFCLASS_S ;
  // rule RL_doFADD_D
  assign CAN_FIRE_RL_doFADD_D =
	     fpu$RDY_request_put && requestR[214] && stateR == 2'd0 &&
	     requestR[213:207] == 7'b1010011 &&
	     requestR[206:200] == 7'h01 ;
  assign WILL_FIRE_RL_doFADD_D = CAN_FIRE_RL_doFADD_D ;
  // rule RL_doFSUB_D
  assign CAN_FIRE_RL_doFSUB_D =
	     fpu$RDY_request_put && requestR[214] && stateR == 2'd0 &&
	     requestR[213:207] == 7'b1010011 &&
	     requestR[206:200] == 7'h05 ;
  assign WILL_FIRE_RL_doFSUB_D = CAN_FIRE_RL_doFSUB_D ;
  // rule RL_doFMUL_D
  assign CAN_FIRE_RL_doFMUL_D =
	     fpu$RDY_request_put && requestR[214] && stateR == 2'd0 &&
	     requestR[213:207] == 7'b1010011 &&
	     requestR[206:200] == 7'h09 ;
  assign WILL_FIRE_RL_doFMUL_D = CAN_FIRE_RL_doFMUL_D ;
  // rule RL_doFMADD_D
  assign CAN_FIRE_RL_doFMADD_D =
	     fpu$RDY_request_put && requestR[214] && stateR == 2'd0 &&
	     requestR[213:207] == 7'b1000011 &&
	     requestR[201:200] == 2'd1 ;
  assign WILL_FIRE_RL_doFMADD_D = CAN_FIRE_RL_doFMADD_D ;
  // rule RL_doFMSUB_D
  assign CAN_FIRE_RL_doFMSUB_D =
	     fpu$RDY_request_put && requestR[214] && stateR == 2'd0 &&
	     requestR[213:207] == 7'b1000111 &&
	     requestR[201:200] == 2'd1 ;
  assign WILL_FIRE_RL_doFMSUB_D = CAN_FIRE_RL_doFMSUB_D ;
  // rule RL_doFNMADD_D
  assign CAN_FIRE_RL_doFNMADD_D =
	     fpu$RDY_request_put && requestR[214] && stateR == 2'd0 &&
	     requestR[213:207] == 7'b1001111 &&
	     requestR[201:200] == 2'd1 ;
  assign WILL_FIRE_RL_doFNMADD_D = CAN_FIRE_RL_doFNMADD_D ;
  // rule RL_doFNMSUB_D
  assign CAN_FIRE_RL_doFNMSUB_D =
	     fpu$RDY_request_put && requestR[214] && stateR == 2'd0 &&
	     requestR[213:207] == 7'b1001011 &&
	     requestR[201:200] == 2'd1 ;
  assign WILL_FIRE_RL_doFNMSUB_D = CAN_FIRE_RL_doFNMSUB_D ;
  // rule RL_doFSGNJ_D
  assign CAN_FIRE_RL_doFSGNJ_D =
	     requestR[214] && stateR == 2'd0 &&
	     requestR[213:207] == 7'b1010011 &&
	     requestR[206:200] == 7'h11 &&
	     requestR[194:192] == 3'h0 ;
  assign WILL_FIRE_RL_doFSGNJ_D = CAN_FIRE_RL_doFSGNJ_D ;
  // rule RL_doFSGNJN_D
  assign CAN_FIRE_RL_doFSGNJN_D =
	     requestR[214] && stateR == 2'd0 &&
	     requestR[213:207] == 7'b1010011 &&
	     requestR[206:200] == 7'h11 &&
	     requestR[194:192] == 3'h1 ;
  assign WILL_FIRE_RL_doFSGNJN_D = CAN_FIRE_RL_doFSGNJN_D ;
  // rule RL_doFSGNJX_D
  assign CAN_FIRE_RL_doFSGNJX_D =
	     requestR[214] && stateR == 2'd0 &&
	     requestR[213:207] == 7'b1010011 &&
	     requestR[206:200] == 7'h11 &&
	     requestR[194:192] == 3'h2 ;
  assign WILL_FIRE_RL_doFSGNJX_D = CAN_FIRE_RL_doFSGNJX_D ;
  // rule RL_doFCVT_D_W
  assign CAN_FIRE_RL_doFCVT_D_W =
	     requestR[214] && stateR == 2'd0 &&
	     requestR[213:207] == 7'b1010011 &&
	     requestR[206:200] == 7'h69 &&
	     requestR[199:195] == 5'd0 ;
  assign WILL_FIRE_RL_doFCVT_D_W = CAN_FIRE_RL_doFCVT_D_W ;
  // rule RL_doFCVT_D_WU
  assign CAN_FIRE_RL_doFCVT_D_WU =
	     requestR[214] && stateR == 2'd0 &&
	     requestR[213:207] == 7'b1010011 &&
	     requestR[206:200] == 7'h69 &&
	     requestR[199:195] == 5'd1 ;
  assign WILL_FIRE_RL_doFCVT_D_WU = CAN_FIRE_RL_doFCVT_D_WU ;
  // rule RL_doFCVT_W_D
  assign CAN_FIRE_RL_doFCVT_W_D =
	     requestR[214] && stateR == 2'd0 &&
	     requestR[213:207] == 7'b1010011 &&
	     requestR[206:200] == 7'h61 &&
	     requestR[199:195] == 5'd0 ;
  assign WILL_FIRE_RL_doFCVT_W_D = CAN_FIRE_RL_doFCVT_W_D ;
  // rule RL_doFCVT_WU_D
  assign CAN_FIRE_RL_doFCVT_WU_D =
	     requestR[214] && stateR == 2'd0 &&
	     requestR[213:207] == 7'b1010011 &&
	     requestR[206:200] == 7'h61 &&
	     requestR[199:195] == 5'd1 ;
  assign WILL_FIRE_RL_doFCVT_WU_D = CAN_FIRE_RL_doFCVT_WU_D ;
  // rule RL_doFCVT_D_L
  assign CAN_FIRE_RL_doFCVT_D_L =
	     requestR[214] && stateR == 2'd0 &&
	     requestR[213:207] == 7'b1010011 &&
	     requestR[206:200] == 7'h69 &&
	     requestR[199:195] == 5'd2 ;
  assign WILL_FIRE_RL_doFCVT_D_L = CAN_FIRE_RL_doFCVT_D_L ;
  // rule RL_doFCVT_D_LU
  assign CAN_FIRE_RL_doFCVT_D_LU =
	     requestR[214] && stateR == 2'd0 &&
	     requestR[213:207] == 7'b1010011 &&
	     requestR[206:200] == 7'h69 &&
	     requestR[199:195] == 5'd3 ;
  assign WILL_FIRE_RL_doFCVT_D_LU = CAN_FIRE_RL_doFCVT_D_LU ;
  // rule RL_doFCVT_L_D
  assign CAN_FIRE_RL_doFCVT_L_D =
	     requestR[214] && stateR == 2'd0 &&
	     requestR[213:207] == 7'b1010011 &&
	     requestR[206:200] == 7'h61 &&
	     requestR[199:195] == 5'd2 ;
  assign WILL_FIRE_RL_doFCVT_L_D = CAN_FIRE_RL_doFCVT_L_D ;
  // rule RL_doFCVT_LU_D
  assign CAN_FIRE_RL_doFCVT_LU_D =
	     requestR[214] && stateR == 2'd0 &&
	     requestR[213:207] == 7'b1010011 &&
	     requestR[206:200] == 7'h61 &&
	     requestR[199:195] == 5'd3 ;
  assign WILL_FIRE_RL_doFCVT_LU_D = CAN_FIRE_RL_doFCVT_LU_D ;
  // rule RL_doFCVT_S_D
  assign CAN_FIRE_RL_doFCVT_S_D =
	     requestR[214] && stateR == 2'd0 &&
	     requestR[213:207] == 7'b1010011 &&
	     requestR[206:200] == 7'h20 &&
	     requestR[199:195] == 5'd1 ;
  assign WILL_FIRE_RL_doFCVT_S_D = CAN_FIRE_RL_doFCVT_S_D ;
  // rule RL_doFCVT_D_S
  assign CAN_FIRE_RL_doFCVT_D_S =
	     requestR[214] && stateR == 2'd0 &&
	     requestR[213:207] == 7'b1010011 &&
	     requestR[206:200] == 7'h21 &&
	     requestR[199:195] == 5'd0 ;
  assign WILL_FIRE_RL_doFCVT_D_S = CAN_FIRE_RL_doFCVT_D_S ;
  // rule RL_doFMIN_D
  assign CAN_FIRE_RL_doFMIN_D =
	     requestR[214] && stateR == 2'd0 &&
	     requestR[213:207] == 7'b1010011 &&
	     requestR[206:200] == 7'h15 &&
	     requestR[194:192] == 3'h0 ;
  assign WILL_FIRE_RL_doFMIN_D = CAN_FIRE_RL_doFMIN_D ;
  // rule RL_doFMAX_D
  assign CAN_FIRE_RL_doFMAX_D =
	     requestR[214] && stateR == 2'd0 &&
	     requestR[213:207] == 7'b1010011 &&
	     requestR[206:200] == 7'h15 &&
	     requestR[194:192] == 3'h1 ;
  assign WILL_FIRE_RL_doFMAX_D = CAN_FIRE_RL_doFMAX_D ;
  // rule RL_doFEQ_D
  assign CAN_FIRE_RL_doFEQ_D =
	     requestR[214] && stateR == 2'd0 &&
	     requestR[213:207] == 7'b1010011 &&
	     requestR[206:200] == 7'h51 &&
	     requestR[194:192] == 3'h2 ;
  assign WILL_FIRE_RL_doFEQ_D = CAN_FIRE_RL_doFEQ_D ;
  // rule RL_doFLT_D
  assign CAN_FIRE_RL_doFLT_D =
	     requestR[214] && stateR == 2'd0 &&
	     requestR[213:207] == 7'b1010011 &&
	     requestR[206:200] == 7'h51 &&
	     requestR[194:192] == 3'h1 ;
  assign WILL_FIRE_RL_doFLT_D = CAN_FIRE_RL_doFLT_D ;
  // rule RL_doFLE_D
  assign CAN_FIRE_RL_doFLE_D =
	     requestR[214] && stateR == 2'd0 &&
	     requestR[213:207] == 7'b1010011 &&
	     requestR[206:200] == 7'h51 &&
	     requestR[194:192] == 3'h0 ;
  assign WILL_FIRE_RL_doFLE_D = CAN_FIRE_RL_doFLE_D ;
  // rule RL_doFMV_D_X
  assign CAN_FIRE_RL_doFMV_D_X =
	     requestR[214] && stateR == 2'd0 &&
	     requestR[213:207] == 7'b1010011 &&
	     requestR[206:200] == 7'h79 &&
	     requestR[194:192] == 3'h0 ;
  assign WILL_FIRE_RL_doFMV_D_X = CAN_FIRE_RL_doFMV_D_X ;
  // rule RL_doFMV_X_D
  assign CAN_FIRE_RL_doFMV_X_D =
	     requestR[214] && stateR == 2'd0 &&
	     requestR[213:207] == 7'b1010011 &&
	     requestR[206:200] == 7'h71 &&
	     requestR[194:192] == 3'h0 ;
  assign WILL_FIRE_RL_doFMV_X_D = CAN_FIRE_RL_doFMV_X_D ;
  // rule RL_doFCLASS_D
  assign CAN_FIRE_RL_doFCLASS_D =
	     requestR[214] && stateR == 2'd0 &&
	     requestR[213:207] == 7'b1010011 &&
	     requestR[206:200] == 7'h71 &&
	     requestR[194:192] == 3'h1 ;
  assign WILL_FIRE_RL_doFCLASS_D = CAN_FIRE_RL_doFCLASS_D ;
  // rule RL_rl_get_fpu_result
  assign CAN_FIRE_RL_rl_get_fpu_result =
	     fpu$RDY_response_get && stateR == 2'd1 ;
  assign WILL_FIRE_RL_rl_get_fpu_result = CAN_FIRE_RL_rl_get_fpu_result ;
  // rule RL_rl_drive_fpu_result
  assign CAN_FIRE_RL_rl_drive_fpu_result = stateR == 2'd2 ;
  assign WILL_FIRE_RL_rl_drive_fpu_result = stateR == 2'd2 ;
  // inputs to muxes for submodule ports
  assign MUX_dw_result$wset_1__SEL_1 =
	     requestR[214] && stateR == 2'd0 &&
	     requestR[213:207] == 7'b1010011 &&
	     requestR[206:200] == 7'h10 &&
	     requestR[194:192] == 3'h1 ;
  assign MUX_dw_result$wset_1__SEL_2 =
	     requestR[214] && stateR == 2'd0 &&
	     requestR[213:207] == 7'b1010011 &&
	     requestR[206:200] == 7'h10 &&
	     requestR[194:192] == 3'h0 ;
  assign MUX_dw_result$wset_1__SEL_38 =
	     WILL_FIRE_RL_doFMV_X_D || WILL_FIRE_RL_doFMV_D_X ;
  assign MUX_dw_result$wset_1__VAL_1 = { x__h1927, 5'd0 } ;
  assign MUX_dw_result$wset_1__VAL_2 = { x__h1781, 5'd0 } ;
  assign MUX_dw_result$wset_1__VAL_3 = { x__h2061, 5'd0 } ;
  assign MUX_dw_result$wset_1__VAL_4 = { x__h2209, x__h13083 } ;
  assign MUX_dw_result$wset_1__VAL_5 = { x__h13371, x__h23674 } ;
  assign MUX_dw_result$wset_1__VAL_6 = { x__h23959, x__h30129 } ;
  assign MUX_dw_result$wset_1__VAL_7 = { x__h30414, x__h36272 } ;
  assign MUX_dw_result$wset_1__VAL_8 = { x__h36556, x__h38337 } ;
  assign MUX_dw_result$wset_1__VAL_9 = { x__h38594, x__h39093 } ;
  assign MUX_dw_result$wset_1__VAL_10 = { x__h39336, x__h40655 } ;
  assign MUX_dw_result$wset_1__VAL_11 = { x__h40912, x__h41414 } ;
  assign MUX_dw_result$wset_1__VAL_12 = { x__h41662, x__h43701 } ;
  assign MUX_dw_result$wset_1__VAL_13 = { x__h44296, x__h43701 } ;
  assign MUX_dw_result$wset_1__VAL_14 = { x__h46821, 5'd0 } ;
  assign MUX_dw_result$wset_1__VAL_15 = { x__h46942, 5'd0 } ;
  assign MUX_dw_result$wset_1__VAL_16 = { x__h47080, x__h43701 } ;
  assign MUX_dw_result$wset_1__VAL_17 = { x__h48563, x__h49451 } ;
  assign MUX_dw_result$wset_1__VAL_18 = { x__h49632, x__h49451 } ;
  assign MUX_dw_result$wset_1__VAL_19 = { x__h50718, 5'd0 } ;
  assign MUX_dw_result$wset_1__VAL_20 = { x__h51885, 5'd0 } ;
  assign MUX_dw_result$wset_1__VAL_21 = { x__h52007, 5'd0 } ;
  assign MUX_dw_result$wset_1__VAL_22 = { x__h52131, 5'd0 } ;
  assign MUX_dw_result$wset_1__VAL_23 = { x__h52261, x__h61924 } ;
  assign MUX_dw_result$wset_1__VAL_24 = { x__h62209, x__h71592 } ;
  assign MUX_dw_result$wset_1__VAL_25 = { x__h71876, x__h73195 } ;
  assign MUX_dw_result$wset_1__VAL_26 = { x__h73452, x__h73954 } ;
  assign MUX_dw_result$wset_1__VAL_27 = { x__h74198, x__h85465 } ;
  assign MUX_dw_result$wset_1__VAL_28 = { x__h85750, x__h96449 } ;
  assign MUX_dw_result$wset_1__VAL_29 = { x__h96733, x__h98497 } ;
  assign MUX_dw_result$wset_1__VAL_30 = { x__h98754, x__h99253 } ;
  assign MUX_dw_result$wset_1__VAL_31 = { x__h99497, x__h147219 } ;
  assign MUX_dw_result$wset_1__VAL_32 = { x__h148202, x__h189005 } ;
  assign MUX_dw_result$wset_1__VAL_33 = { x__h189928, x__h193477 } ;
  assign MUX_dw_result$wset_1__VAL_34 = { x__h194476, x__h193477 } ;
  assign MUX_dw_result$wset_1__VAL_35 = { x__h198920, x__h193477 } ;
  assign MUX_dw_result$wset_1__VAL_36 = { x__h201615, x__h203311 } ;
  assign MUX_dw_result$wset_1__VAL_37 = { x__h203492, x__h203311 } ;
  assign MUX_dw_result$wset_1__VAL_38 = { requestR[191:128], 5'd0 } ;
  assign MUX_dw_result$wset_1__VAL_39 = { x__h205619, 5'd0 } ;
  assign MUX_dw_result$wset_1__VAL_40 =
	     { x__h206269, fpu$response_get[4:0] } ;
  assign MUX_fpu$request_put_1__VAL_1 =
	     { 33'h1AAAAAAAA,
	       requestR[191:160] == 32'hFFFFFFFF && requestR[159],
	       IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d19,
	       33'h1AAAAAAAA,
	       requestR_BITS_127_TO_96_2_EQ_0xFFFFFFFF_3_AND__ETC___d28,
	       65'h0AAAAAAAAAAAAAAAA,
	       IF_requestR_BITS_194_TO_192_0_EQ_0x0_1_THEN_re_ETC___d40,
	       4'd0 } ;
  assign MUX_fpu$request_put_1__VAL_2 =
	     { 33'h1AAAAAAAA,
	       requestR[191:160] == 32'hFFFFFFFF && requestR[159],
	       IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d19,
	       33'h1AAAAAAAA,
	       requestR_BITS_127_TO_96_2_EQ_0xFFFFFFFF_3_AND__ETC___d28,
	       65'h0AAAAAAAAAAAAAAAA,
	       IF_requestR_BITS_194_TO_192_0_EQ_0x0_1_THEN_re_ETC___d40,
	       4'd1 } ;
  assign MUX_fpu$request_put_1__VAL_3 =
	     { 33'h1AAAAAAAA,
	       requestR[191:160] == 32'hFFFFFFFF && requestR[159],
	       IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d19,
	       33'h1AAAAAAAA,
	       requestR_BITS_127_TO_96_2_EQ_0xFFFFFFFF_3_AND__ETC___d28,
	       65'h0AAAAAAAAAAAAAAAA,
	       IF_requestR_BITS_194_TO_192_0_EQ_0x0_1_THEN_re_ETC___d40,
	       4'd2 } ;
  assign MUX_fpu$request_put_1__VAL_4 =
	     { 33'h1AAAAAAAA,
	       requestR[191:160] == 32'hFFFFFFFF && requestR[159],
	       IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d19,
	       33'h1AAAAAAAA,
	       requestR_BITS_127_TO_96_2_EQ_0xFFFFFFFF_3_AND__ETC___d28,
	       _1_CONCAT_DONTCARE_CONCAT_requestR_BITS_63_TO_3_ETC___d68,
	       IF_requestR_BITS_194_TO_192_0_EQ_0x0_1_THEN_re_ETC___d40,
	       4'd5 } ;
  assign MUX_fpu$request_put_1__VAL_5 =
	     { 33'h1AAAAAAAA,
	       requestR[191:160] == 32'hFFFFFFFF && requestR[159],
	       IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d19,
	       33'h1AAAAAAAA,
	       requestR_BITS_127_TO_96_2_EQ_0xFFFFFFFF_3_AND__ETC___d28,
	       _1_CONCAT_DONTCARE_CONCAT_requestR_BITS_63_TO_3_ETC___d68,
	       IF_requestR_BITS_194_TO_192_0_EQ_0x0_1_THEN_re_ETC___d40,
	       4'd6 } ;
  assign MUX_fpu$request_put_1__VAL_6 =
	     { 33'h1AAAAAAAA,
	       requestR[191:160] == 32'hFFFFFFFF && requestR[159],
	       IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d19,
	       33'h1AAAAAAAA,
	       requestR_BITS_127_TO_96_2_EQ_0xFFFFFFFF_3_AND__ETC___d28,
	       _1_CONCAT_DONTCARE_CONCAT_requestR_BITS_63_TO_3_ETC___d68,
	       IF_requestR_BITS_194_TO_192_0_EQ_0x0_1_THEN_re_ETC___d40,
	       4'd7 } ;
  assign MUX_fpu$request_put_1__VAL_7 =
	     { 33'h1AAAAAAAA,
	       requestR[191:160] == 32'hFFFFFFFF && requestR[159],
	       IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d19,
	       33'h1AAAAAAAA,
	       requestR_BITS_127_TO_96_2_EQ_0xFFFFFFFF_3_AND__ETC___d28,
	       _1_CONCAT_DONTCARE_CONCAT_requestR_BITS_63_TO_3_ETC___d68,
	       IF_requestR_BITS_194_TO_192_0_EQ_0x0_1_THEN_re_ETC___d40,
	       4'd8 } ;
  assign MUX_fpu$request_put_1__VAL_8 =
	     { 1'd0,
	       requestR[191:128],
	       1'd0,
	       requestR[127:64],
	       65'h0AAAAAAAAAAAAAAAA,
	       IF_requestR_BITS_194_TO_192_0_EQ_0x0_1_THEN_re_ETC___d40,
	       4'd0 } ;
  assign MUX_fpu$request_put_1__VAL_9 =
	     { 1'd0,
	       requestR[191:128],
	       1'd0,
	       requestR[127:64],
	       65'h0AAAAAAAAAAAAAAAA,
	       IF_requestR_BITS_194_TO_192_0_EQ_0x0_1_THEN_re_ETC___d40,
	       4'd1 } ;
  assign MUX_fpu$request_put_1__VAL_10 =
	     { 1'd0,
	       requestR[191:128],
	       1'd0,
	       requestR[127:64],
	       65'h0AAAAAAAAAAAAAAAA,
	       IF_requestR_BITS_194_TO_192_0_EQ_0x0_1_THEN_re_ETC___d40,
	       4'd2 } ;
  assign MUX_fpu$request_put_1__VAL_11 =
	     { 1'd0,
	       requestR[191:128],
	       1'd0,
	       requestR[127:64],
	       1'd0,
	       requestR[63:0],
	       IF_requestR_BITS_194_TO_192_0_EQ_0x0_1_THEN_re_ETC___d40,
	       4'd5 } ;
  assign MUX_fpu$request_put_1__VAL_12 =
	     { 1'd0,
	       requestR[191:128],
	       1'd0,
	       requestR[127:64],
	       1'd0,
	       requestR[63:0],
	       IF_requestR_BITS_194_TO_192_0_EQ_0x0_1_THEN_re_ETC___d40,
	       4'd6 } ;
  assign MUX_fpu$request_put_1__VAL_13 =
	     { 1'd0,
	       requestR[191:128],
	       1'd0,
	       requestR[127:64],
	       1'd0,
	       requestR[63:0],
	       IF_requestR_BITS_194_TO_192_0_EQ_0x0_1_THEN_re_ETC___d40,
	       4'd7 } ;
  assign MUX_fpu$request_put_1__VAL_14 =
	     { 1'd0,
	       requestR[191:128],
	       1'd0,
	       requestR[127:64],
	       1'd0,
	       requestR[63:0],
	       IF_requestR_BITS_194_TO_192_0_EQ_0x0_1_THEN_re_ETC___d40,
	       4'd8 } ;
  assign MUX_resultR$write_1__VAL_2 =
	     { 1'd1, x__h206269, fpu$response_get[4:0] } ;
  assign MUX_resultR$write_1__VAL_3 = { 1'd1, x__h205619, 5'd0 } ;
  assign MUX_resultR$write_1__VAL_4 = { 1'd1, requestR[191:128], 5'd0 } ;
  assign MUX_resultR$write_1__VAL_6 = { 1'd1, x__h203492, x__h203311 } ;
  assign MUX_resultR$write_1__VAL_7 = { 1'd1, x__h201615, x__h203311 } ;
  assign MUX_resultR$write_1__VAL_8 = { 1'd1, x__h198920, x__h193477 } ;
  assign MUX_resultR$write_1__VAL_9 = { 1'd1, x__h194476, x__h193477 } ;
  assign MUX_resultR$write_1__VAL_10 = { 1'd1, x__h189928, x__h193477 } ;
  assign MUX_resultR$write_1__VAL_11 = { 1'd1, x__h148202, x__h189005 } ;
  assign MUX_resultR$write_1__VAL_12 = { 1'd1, x__h99497, x__h147219 } ;
  assign MUX_resultR$write_1__VAL_13 = { 1'd1, x__h98754, x__h99253 } ;
  assign MUX_resultR$write_1__VAL_14 = { 1'd1, x__h96733, x__h98497 } ;
  assign MUX_resultR$write_1__VAL_15 = { 1'd1, x__h85750, x__h96449 } ;
  assign MUX_resultR$write_1__VAL_16 = { 1'd1, x__h74198, x__h85465 } ;
  assign MUX_resultR$write_1__VAL_17 = { 1'd1, x__h73452, x__h73954 } ;
  assign MUX_resultR$write_1__VAL_18 = { 1'd1, x__h71876, x__h73195 } ;
  assign MUX_resultR$write_1__VAL_19 = { 1'd1, x__h62209, x__h71592 } ;
  assign MUX_resultR$write_1__VAL_20 = { 1'd1, x__h52261, x__h61924 } ;
  assign MUX_resultR$write_1__VAL_21 = { 1'd1, x__h52131, 5'd0 } ;
  assign MUX_resultR$write_1__VAL_22 = { 1'd1, x__h52007, 5'd0 } ;
  assign MUX_resultR$write_1__VAL_23 = { 1'd1, x__h51885, 5'd0 } ;
  assign MUX_resultR$write_1__VAL_24 = { 1'd1, x__h50718, 5'd0 } ;
  assign MUX_resultR$write_1__VAL_25 = { 1'd1, x__h49632, x__h49451 } ;
  assign MUX_resultR$write_1__VAL_26 = { 1'd1, x__h48563, x__h49451 } ;
  assign MUX_resultR$write_1__VAL_27 = { 1'd1, x__h47080, x__h43701 } ;
  assign MUX_resultR$write_1__VAL_28 = { 1'd1, x__h46942, 5'd0 } ;
  assign MUX_resultR$write_1__VAL_29 = { 1'd1, x__h46821, 5'd0 } ;
  assign MUX_resultR$write_1__VAL_30 = { 1'd1, x__h44296, x__h43701 } ;
  assign MUX_resultR$write_1__VAL_31 = { 1'd1, x__h41662, x__h43701 } ;
  assign MUX_resultR$write_1__VAL_32 = { 1'd1, x__h40912, x__h41414 } ;
  assign MUX_resultR$write_1__VAL_33 = { 1'd1, x__h39336, x__h40655 } ;
  assign MUX_resultR$write_1__VAL_34 = { 1'd1, x__h38594, x__h39093 } ;
  assign MUX_resultR$write_1__VAL_35 = { 1'd1, x__h36556, x__h38337 } ;
  assign MUX_resultR$write_1__VAL_36 = { 1'd1, x__h30414, x__h36272 } ;
  assign MUX_resultR$write_1__VAL_37 = { 1'd1, x__h23959, x__h30129 } ;
  assign MUX_resultR$write_1__VAL_38 = { 1'd1, x__h13371, x__h23674 } ;
  assign MUX_resultR$write_1__VAL_39 = { 1'd1, x__h2209, x__h13083 } ;
  assign MUX_resultR$write_1__VAL_40 = { 1'd1, x__h2061, 5'd0 } ;
  assign MUX_resultR$write_1__VAL_41 = { 1'd1, x__h1927, 5'd0 } ;
  assign MUX_resultR$write_1__VAL_42 = { 1'd1, x__h1781, 5'd0 } ;
  // inlined wires
  assign dw_valid$wget = !WILL_FIRE_RL_rl_drive_fpu_result || resultR[69] ;
  assign dw_valid$whas =
	     WILL_FIRE_RL_rl_drive_fpu_result ||
	     WILL_FIRE_RL_rl_get_fpu_result ||
	     WILL_FIRE_RL_doFCLASS_D ||
	     WILL_FIRE_RL_doFMV_X_D ||
	     WILL_FIRE_RL_doFMV_D_X ||
	     WILL_FIRE_RL_doFLE_D ||
	     WILL_FIRE_RL_doFLT_D ||
	     WILL_FIRE_RL_doFEQ_D ||
	     WILL_FIRE_RL_doFMAX_D ||
	     WILL_FIRE_RL_doFMIN_D ||
	     WILL_FIRE_RL_doFCVT_D_S ||
	     WILL_FIRE_RL_doFCVT_S_D ||
	     WILL_FIRE_RL_doFCVT_LU_D ||
	     WILL_FIRE_RL_doFCVT_L_D ||
	     WILL_FIRE_RL_doFCVT_D_LU ||
	     WILL_FIRE_RL_doFCVT_D_L ||
	     WILL_FIRE_RL_doFCVT_WU_D ||
	     WILL_FIRE_RL_doFCVT_W_D ||
	     WILL_FIRE_RL_doFCVT_D_WU ||
	     WILL_FIRE_RL_doFCVT_D_W ||
	     WILL_FIRE_RL_doFSGNJX_D ||
	     WILL_FIRE_RL_doFSGNJN_D ||
	     WILL_FIRE_RL_doFSGNJ_D ||
	     WILL_FIRE_RL_doFCLASS_S ||
	     WILL_FIRE_RL_doFLE_S ||
	     WILL_FIRE_RL_doFLT_S ||
	     WILL_FIRE_RL_doFEQ_S ||
	     WILL_FIRE_RL_doFMV_X_W ||
	     WILL_FIRE_RL_doFMV_W_X ||
	     WILL_FIRE_RL_doFMAX_S ||
	     WILL_FIRE_RL_doFMIN_S ||
	     WILL_FIRE_RL_doFCVT_WU_S ||
	     WILL_FIRE_RL_doFCVT_W_S ||
	     WILL_FIRE_RL_doFCVT_LU_S ||
	     WILL_FIRE_RL_doFCVT_L_S ||
	     WILL_FIRE_RL_doFCVT_S_WU ||
	     WILL_FIRE_RL_doFCVT_S_W ||
	     WILL_FIRE_RL_doFCVT_S_LU ||
	     WILL_FIRE_RL_doFCVT_S_L ||
	     WILL_FIRE_RL_doFSGNJX_S ||
	     WILL_FIRE_RL_doFSGNJN_S ||
	     WILL_FIRE_RL_doFSGNJ_S ;
  always@(WILL_FIRE_RL_doFSGNJN_S or
	  MUX_dw_result$wset_1__VAL_1 or
	  WILL_FIRE_RL_doFSGNJ_S or
	  MUX_dw_result$wset_1__VAL_2 or
	  WILL_FIRE_RL_doFSGNJX_S or
	  MUX_dw_result$wset_1__VAL_3 or
	  WILL_FIRE_RL_doFCVT_S_L or
	  MUX_dw_result$wset_1__VAL_4 or
	  WILL_FIRE_RL_doFCVT_S_LU or
	  MUX_dw_result$wset_1__VAL_5 or
	  WILL_FIRE_RL_doFCVT_S_W or
	  MUX_dw_result$wset_1__VAL_6 or
	  WILL_FIRE_RL_doFCVT_S_WU or
	  MUX_dw_result$wset_1__VAL_7 or
	  WILL_FIRE_RL_doFCVT_L_S or
	  MUX_dw_result$wset_1__VAL_8 or
	  WILL_FIRE_RL_doFCVT_LU_S or
	  MUX_dw_result$wset_1__VAL_9 or
	  WILL_FIRE_RL_doFCVT_W_S or
	  MUX_dw_result$wset_1__VAL_10 or
	  WILL_FIRE_RL_doFCVT_WU_S or
	  MUX_dw_result$wset_1__VAL_11 or
	  WILL_FIRE_RL_doFMIN_S or
	  MUX_dw_result$wset_1__VAL_12 or
	  WILL_FIRE_RL_doFMAX_S or
	  MUX_dw_result$wset_1__VAL_13 or
	  WILL_FIRE_RL_doFMV_W_X or
	  MUX_dw_result$wset_1__VAL_14 or
	  WILL_FIRE_RL_doFMV_X_W or
	  MUX_dw_result$wset_1__VAL_15 or
	  WILL_FIRE_RL_doFEQ_S or
	  MUX_dw_result$wset_1__VAL_16 or
	  WILL_FIRE_RL_doFLT_S or
	  MUX_dw_result$wset_1__VAL_17 or
	  WILL_FIRE_RL_doFLE_S or
	  MUX_dw_result$wset_1__VAL_18 or
	  WILL_FIRE_RL_doFCLASS_S or
	  MUX_dw_result$wset_1__VAL_19 or
	  WILL_FIRE_RL_doFSGNJ_D or
	  MUX_dw_result$wset_1__VAL_20 or
	  WILL_FIRE_RL_doFSGNJN_D or
	  MUX_dw_result$wset_1__VAL_21 or
	  WILL_FIRE_RL_doFSGNJX_D or
	  MUX_dw_result$wset_1__VAL_22 or
	  WILL_FIRE_RL_doFCVT_D_W or
	  MUX_dw_result$wset_1__VAL_23 or
	  WILL_FIRE_RL_doFCVT_D_WU or
	  MUX_dw_result$wset_1__VAL_24 or
	  WILL_FIRE_RL_doFCVT_W_D or
	  MUX_dw_result$wset_1__VAL_25 or
	  WILL_FIRE_RL_doFCVT_WU_D or
	  MUX_dw_result$wset_1__VAL_26 or
	  WILL_FIRE_RL_doFCVT_D_L or
	  MUX_dw_result$wset_1__VAL_27 or
	  WILL_FIRE_RL_doFCVT_D_LU or
	  MUX_dw_result$wset_1__VAL_28 or
	  WILL_FIRE_RL_doFCVT_L_D or
	  MUX_dw_result$wset_1__VAL_29 or
	  WILL_FIRE_RL_doFCVT_LU_D or
	  MUX_dw_result$wset_1__VAL_30 or
	  WILL_FIRE_RL_doFCVT_S_D or
	  MUX_dw_result$wset_1__VAL_31 or
	  WILL_FIRE_RL_doFCVT_D_S or
	  MUX_dw_result$wset_1__VAL_32 or
	  WILL_FIRE_RL_doFMIN_D or
	  MUX_dw_result$wset_1__VAL_33 or
	  WILL_FIRE_RL_doFMAX_D or
	  MUX_dw_result$wset_1__VAL_34 or
	  WILL_FIRE_RL_doFEQ_D or
	  MUX_dw_result$wset_1__VAL_35 or
	  WILL_FIRE_RL_doFLT_D or
	  MUX_dw_result$wset_1__VAL_36 or
	  WILL_FIRE_RL_doFLE_D or
	  MUX_dw_result$wset_1__VAL_37 or
	  MUX_dw_result$wset_1__SEL_38 or
	  MUX_dw_result$wset_1__VAL_38 or
	  WILL_FIRE_RL_doFCLASS_D or
	  MUX_dw_result$wset_1__VAL_39 or
	  WILL_FIRE_RL_rl_get_fpu_result or
	  MUX_dw_result$wset_1__VAL_40 or
	  WILL_FIRE_RL_rl_drive_fpu_result or resultR)
  begin
    case (1'b1) // synopsys parallel_case
      WILL_FIRE_RL_doFSGNJN_S: dw_result$wget = MUX_dw_result$wset_1__VAL_1;
      WILL_FIRE_RL_doFSGNJ_S: dw_result$wget = MUX_dw_result$wset_1__VAL_2;
      WILL_FIRE_RL_doFSGNJX_S: dw_result$wget = MUX_dw_result$wset_1__VAL_3;
      WILL_FIRE_RL_doFCVT_S_L: dw_result$wget = MUX_dw_result$wset_1__VAL_4;
      WILL_FIRE_RL_doFCVT_S_LU: dw_result$wget = MUX_dw_result$wset_1__VAL_5;
      WILL_FIRE_RL_doFCVT_S_W: dw_result$wget = MUX_dw_result$wset_1__VAL_6;
      WILL_FIRE_RL_doFCVT_S_WU: dw_result$wget = MUX_dw_result$wset_1__VAL_7;
      WILL_FIRE_RL_doFCVT_L_S: dw_result$wget = MUX_dw_result$wset_1__VAL_8;
      WILL_FIRE_RL_doFCVT_LU_S: dw_result$wget = MUX_dw_result$wset_1__VAL_9;
      WILL_FIRE_RL_doFCVT_W_S: dw_result$wget = MUX_dw_result$wset_1__VAL_10;
      WILL_FIRE_RL_doFCVT_WU_S: dw_result$wget = MUX_dw_result$wset_1__VAL_11;
      WILL_FIRE_RL_doFMIN_S: dw_result$wget = MUX_dw_result$wset_1__VAL_12;
      WILL_FIRE_RL_doFMAX_S: dw_result$wget = MUX_dw_result$wset_1__VAL_13;
      WILL_FIRE_RL_doFMV_W_X: dw_result$wget = MUX_dw_result$wset_1__VAL_14;
      WILL_FIRE_RL_doFMV_X_W: dw_result$wget = MUX_dw_result$wset_1__VAL_15;
      WILL_FIRE_RL_doFEQ_S: dw_result$wget = MUX_dw_result$wset_1__VAL_16;
      WILL_FIRE_RL_doFLT_S: dw_result$wget = MUX_dw_result$wset_1__VAL_17;
      WILL_FIRE_RL_doFLE_S: dw_result$wget = MUX_dw_result$wset_1__VAL_18;
      WILL_FIRE_RL_doFCLASS_S: dw_result$wget = MUX_dw_result$wset_1__VAL_19;
      WILL_FIRE_RL_doFSGNJ_D: dw_result$wget = MUX_dw_result$wset_1__VAL_20;
      WILL_FIRE_RL_doFSGNJN_D: dw_result$wget = MUX_dw_result$wset_1__VAL_21;
      WILL_FIRE_RL_doFSGNJX_D: dw_result$wget = MUX_dw_result$wset_1__VAL_22;
      WILL_FIRE_RL_doFCVT_D_W: dw_result$wget = MUX_dw_result$wset_1__VAL_23;
      WILL_FIRE_RL_doFCVT_D_WU: dw_result$wget = MUX_dw_result$wset_1__VAL_24;
      WILL_FIRE_RL_doFCVT_W_D: dw_result$wget = MUX_dw_result$wset_1__VAL_25;
      WILL_FIRE_RL_doFCVT_WU_D: dw_result$wget = MUX_dw_result$wset_1__VAL_26;
      WILL_FIRE_RL_doFCVT_D_L: dw_result$wget = MUX_dw_result$wset_1__VAL_27;
      WILL_FIRE_RL_doFCVT_D_LU: dw_result$wget = MUX_dw_result$wset_1__VAL_28;
      WILL_FIRE_RL_doFCVT_L_D: dw_result$wget = MUX_dw_result$wset_1__VAL_29;
      WILL_FIRE_RL_doFCVT_LU_D: dw_result$wget = MUX_dw_result$wset_1__VAL_30;
      WILL_FIRE_RL_doFCVT_S_D: dw_result$wget = MUX_dw_result$wset_1__VAL_31;
      WILL_FIRE_RL_doFCVT_D_S: dw_result$wget = MUX_dw_result$wset_1__VAL_32;
      WILL_FIRE_RL_doFMIN_D: dw_result$wget = MUX_dw_result$wset_1__VAL_33;
      WILL_FIRE_RL_doFMAX_D: dw_result$wget = MUX_dw_result$wset_1__VAL_34;
      WILL_FIRE_RL_doFEQ_D: dw_result$wget = MUX_dw_result$wset_1__VAL_35;
      WILL_FIRE_RL_doFLT_D: dw_result$wget = MUX_dw_result$wset_1__VAL_36;
      WILL_FIRE_RL_doFLE_D: dw_result$wget = MUX_dw_result$wset_1__VAL_37;
      MUX_dw_result$wset_1__SEL_38:
	  dw_result$wget = MUX_dw_result$wset_1__VAL_38;
      WILL_FIRE_RL_doFCLASS_D: dw_result$wget = MUX_dw_result$wset_1__VAL_39;
      WILL_FIRE_RL_rl_get_fpu_result:
	  dw_result$wget = MUX_dw_result$wset_1__VAL_40;
      WILL_FIRE_RL_rl_drive_fpu_result: dw_result$wget = resultR[68:0];
      default: dw_result$wget =
		   69'h0AAAAAAAAAAAAAAAAA /* unspecified value */ ;
    endcase
  end
  // register cfg_verbosity
  assign cfg_verbosity$D_IN = set_verbosity_verbosity ;
  assign cfg_verbosity$EN = EN_set_verbosity ;
  // register requestR
  assign requestR$D_IN =
	     { 1'd1,
	       req_opcode,
	       req_f7,
	       req_rs2,
	       req_rm,
	       req_v1,
	       req_v2,
	       req_v3 } ;
  assign requestR$EN = EN_req ;
  // register resultR
  always@(EN_req or
	  WILL_FIRE_RL_rl_get_fpu_result or
	  MUX_resultR$write_1__VAL_2 or
	  WILL_FIRE_RL_doFCLASS_D or
	  MUX_resultR$write_1__VAL_3 or
	  WILL_FIRE_RL_doFMV_X_D or
	  MUX_resultR$write_1__VAL_4 or
	  WILL_FIRE_RL_doFMV_D_X or
	  WILL_FIRE_RL_doFLE_D or
	  MUX_resultR$write_1__VAL_6 or
	  WILL_FIRE_RL_doFLT_D or
	  MUX_resultR$write_1__VAL_7 or
	  WILL_FIRE_RL_doFEQ_D or
	  MUX_resultR$write_1__VAL_8 or
	  WILL_FIRE_RL_doFMAX_D or
	  MUX_resultR$write_1__VAL_9 or
	  WILL_FIRE_RL_doFMIN_D or
	  MUX_resultR$write_1__VAL_10 or
	  WILL_FIRE_RL_doFCVT_D_S or
	  MUX_resultR$write_1__VAL_11 or
	  WILL_FIRE_RL_doFCVT_S_D or
	  MUX_resultR$write_1__VAL_12 or
	  WILL_FIRE_RL_doFCVT_LU_D or
	  MUX_resultR$write_1__VAL_13 or
	  WILL_FIRE_RL_doFCVT_L_D or
	  MUX_resultR$write_1__VAL_14 or
	  WILL_FIRE_RL_doFCVT_D_LU or
	  MUX_resultR$write_1__VAL_15 or
	  WILL_FIRE_RL_doFCVT_D_L or
	  MUX_resultR$write_1__VAL_16 or
	  WILL_FIRE_RL_doFCVT_WU_D or
	  MUX_resultR$write_1__VAL_17 or
	  WILL_FIRE_RL_doFCVT_W_D or
	  MUX_resultR$write_1__VAL_18 or
	  WILL_FIRE_RL_doFCVT_D_WU or
	  MUX_resultR$write_1__VAL_19 or
	  WILL_FIRE_RL_doFCVT_D_W or
	  MUX_resultR$write_1__VAL_20 or
	  WILL_FIRE_RL_doFSGNJX_D or
	  MUX_resultR$write_1__VAL_21 or
	  WILL_FIRE_RL_doFSGNJN_D or
	  MUX_resultR$write_1__VAL_22 or
	  WILL_FIRE_RL_doFSGNJ_D or
	  MUX_resultR$write_1__VAL_23 or
	  WILL_FIRE_RL_doFCLASS_S or
	  MUX_resultR$write_1__VAL_24 or
	  WILL_FIRE_RL_doFLE_S or
	  MUX_resultR$write_1__VAL_25 or
	  WILL_FIRE_RL_doFLT_S or
	  MUX_resultR$write_1__VAL_26 or
	  WILL_FIRE_RL_doFEQ_S or
	  MUX_resultR$write_1__VAL_27 or
	  WILL_FIRE_RL_doFMV_X_W or
	  MUX_resultR$write_1__VAL_28 or
	  WILL_FIRE_RL_doFMV_W_X or
	  MUX_resultR$write_1__VAL_29 or
	  WILL_FIRE_RL_doFMAX_S or
	  MUX_resultR$write_1__VAL_30 or
	  WILL_FIRE_RL_doFMIN_S or
	  MUX_resultR$write_1__VAL_31 or
	  WILL_FIRE_RL_doFCVT_WU_S or
	  MUX_resultR$write_1__VAL_32 or
	  WILL_FIRE_RL_doFCVT_W_S or
	  MUX_resultR$write_1__VAL_33 or
	  WILL_FIRE_RL_doFCVT_LU_S or
	  MUX_resultR$write_1__VAL_34 or
	  WILL_FIRE_RL_doFCVT_L_S or
	  MUX_resultR$write_1__VAL_35 or
	  WILL_FIRE_RL_doFCVT_S_WU or
	  MUX_resultR$write_1__VAL_36 or
	  WILL_FIRE_RL_doFCVT_S_W or
	  MUX_resultR$write_1__VAL_37 or
	  WILL_FIRE_RL_doFCVT_S_LU or
	  MUX_resultR$write_1__VAL_38 or
	  WILL_FIRE_RL_doFCVT_S_L or
	  MUX_resultR$write_1__VAL_39 or
	  WILL_FIRE_RL_doFSGNJX_S or
	  MUX_resultR$write_1__VAL_40 or
	  WILL_FIRE_RL_doFSGNJN_S or
	  MUX_resultR$write_1__VAL_41 or
	  WILL_FIRE_RL_doFSGNJ_S or MUX_resultR$write_1__VAL_42)
  case (1'b1)
    EN_req: resultR$D_IN = 70'h0AAAAAAAAAAAAAAAAA;
    WILL_FIRE_RL_rl_get_fpu_result: resultR$D_IN = MUX_resultR$write_1__VAL_2;
    WILL_FIRE_RL_doFCLASS_D: resultR$D_IN = MUX_resultR$write_1__VAL_3;
    WILL_FIRE_RL_doFMV_X_D: resultR$D_IN = MUX_resultR$write_1__VAL_4;
    WILL_FIRE_RL_doFMV_D_X: resultR$D_IN = MUX_resultR$write_1__VAL_4;
    WILL_FIRE_RL_doFLE_D: resultR$D_IN = MUX_resultR$write_1__VAL_6;
    WILL_FIRE_RL_doFLT_D: resultR$D_IN = MUX_resultR$write_1__VAL_7;
    WILL_FIRE_RL_doFEQ_D: resultR$D_IN = MUX_resultR$write_1__VAL_8;
    WILL_FIRE_RL_doFMAX_D: resultR$D_IN = MUX_resultR$write_1__VAL_9;
    WILL_FIRE_RL_doFMIN_D: resultR$D_IN = MUX_resultR$write_1__VAL_10;
    WILL_FIRE_RL_doFCVT_D_S: resultR$D_IN = MUX_resultR$write_1__VAL_11;
    WILL_FIRE_RL_doFCVT_S_D: resultR$D_IN = MUX_resultR$write_1__VAL_12;
    WILL_FIRE_RL_doFCVT_LU_D: resultR$D_IN = MUX_resultR$write_1__VAL_13;
    WILL_FIRE_RL_doFCVT_L_D: resultR$D_IN = MUX_resultR$write_1__VAL_14;
    WILL_FIRE_RL_doFCVT_D_LU: resultR$D_IN = MUX_resultR$write_1__VAL_15;
    WILL_FIRE_RL_doFCVT_D_L: resultR$D_IN = MUX_resultR$write_1__VAL_16;
    WILL_FIRE_RL_doFCVT_WU_D: resultR$D_IN = MUX_resultR$write_1__VAL_17;
    WILL_FIRE_RL_doFCVT_W_D: resultR$D_IN = MUX_resultR$write_1__VAL_18;
    WILL_FIRE_RL_doFCVT_D_WU: resultR$D_IN = MUX_resultR$write_1__VAL_19;
    WILL_FIRE_RL_doFCVT_D_W: resultR$D_IN = MUX_resultR$write_1__VAL_20;
    WILL_FIRE_RL_doFSGNJX_D: resultR$D_IN = MUX_resultR$write_1__VAL_21;
    WILL_FIRE_RL_doFSGNJN_D: resultR$D_IN = MUX_resultR$write_1__VAL_22;
    WILL_FIRE_RL_doFSGNJ_D: resultR$D_IN = MUX_resultR$write_1__VAL_23;
    WILL_FIRE_RL_doFCLASS_S: resultR$D_IN = MUX_resultR$write_1__VAL_24;
    WILL_FIRE_RL_doFLE_S: resultR$D_IN = MUX_resultR$write_1__VAL_25;
    WILL_FIRE_RL_doFLT_S: resultR$D_IN = MUX_resultR$write_1__VAL_26;
    WILL_FIRE_RL_doFEQ_S: resultR$D_IN = MUX_resultR$write_1__VAL_27;
    WILL_FIRE_RL_doFMV_X_W: resultR$D_IN = MUX_resultR$write_1__VAL_28;
    WILL_FIRE_RL_doFMV_W_X: resultR$D_IN = MUX_resultR$write_1__VAL_29;
    WILL_FIRE_RL_doFMAX_S: resultR$D_IN = MUX_resultR$write_1__VAL_30;
    WILL_FIRE_RL_doFMIN_S: resultR$D_IN = MUX_resultR$write_1__VAL_31;
    WILL_FIRE_RL_doFCVT_WU_S: resultR$D_IN = MUX_resultR$write_1__VAL_32;
    WILL_FIRE_RL_doFCVT_W_S: resultR$D_IN = MUX_resultR$write_1__VAL_33;
    WILL_FIRE_RL_doFCVT_LU_S: resultR$D_IN = MUX_resultR$write_1__VAL_34;
    WILL_FIRE_RL_doFCVT_L_S: resultR$D_IN = MUX_resultR$write_1__VAL_35;
    WILL_FIRE_RL_doFCVT_S_WU: resultR$D_IN = MUX_resultR$write_1__VAL_36;
    WILL_FIRE_RL_doFCVT_S_W: resultR$D_IN = MUX_resultR$write_1__VAL_37;
    WILL_FIRE_RL_doFCVT_S_LU: resultR$D_IN = MUX_resultR$write_1__VAL_38;
    WILL_FIRE_RL_doFCVT_S_L: resultR$D_IN = MUX_resultR$write_1__VAL_39;
    WILL_FIRE_RL_doFSGNJX_S: resultR$D_IN = MUX_resultR$write_1__VAL_40;
    WILL_FIRE_RL_doFSGNJN_S: resultR$D_IN = MUX_resultR$write_1__VAL_41;
    WILL_FIRE_RL_doFSGNJ_S: resultR$D_IN = MUX_resultR$write_1__VAL_42;
    default: resultR$D_IN = 70'h2AAAAAAAAAAAAAAAAA /* unspecified value */ ;
  endcase
  assign resultR$EN =
	     EN_req || WILL_FIRE_RL_doFMV_X_D || WILL_FIRE_RL_doFMV_D_X ||
	     WILL_FIRE_RL_doFSGNJ_S ||
	     WILL_FIRE_RL_doFSGNJN_S ||
	     WILL_FIRE_RL_doFSGNJX_S ||
	     WILL_FIRE_RL_doFCVT_S_L ||
	     WILL_FIRE_RL_doFCVT_S_LU ||
	     WILL_FIRE_RL_doFCVT_S_W ||
	     WILL_FIRE_RL_doFCVT_S_WU ||
	     WILL_FIRE_RL_doFCVT_L_S ||
	     WILL_FIRE_RL_doFCVT_LU_S ||
	     WILL_FIRE_RL_doFCVT_W_S ||
	     WILL_FIRE_RL_doFCVT_WU_S ||
	     WILL_FIRE_RL_doFMIN_S ||
	     WILL_FIRE_RL_doFMAX_S ||
	     WILL_FIRE_RL_doFMV_W_X ||
	     WILL_FIRE_RL_doFMV_X_W ||
	     WILL_FIRE_RL_doFEQ_S ||
	     WILL_FIRE_RL_doFLT_S ||
	     WILL_FIRE_RL_doFLE_S ||
	     WILL_FIRE_RL_doFCLASS_S ||
	     WILL_FIRE_RL_doFSGNJ_D ||
	     WILL_FIRE_RL_doFSGNJN_D ||
	     WILL_FIRE_RL_doFSGNJX_D ||
	     WILL_FIRE_RL_doFCVT_D_W ||
	     WILL_FIRE_RL_doFCVT_D_WU ||
	     WILL_FIRE_RL_doFCVT_W_D ||
	     WILL_FIRE_RL_doFCVT_WU_D ||
	     WILL_FIRE_RL_doFCVT_D_L ||
	     WILL_FIRE_RL_doFCVT_D_LU ||
	     WILL_FIRE_RL_doFCVT_L_D ||
	     WILL_FIRE_RL_doFCVT_LU_D ||
	     WILL_FIRE_RL_doFCVT_S_D ||
	     WILL_FIRE_RL_doFCVT_D_S ||
	     WILL_FIRE_RL_doFMIN_D ||
	     WILL_FIRE_RL_doFMAX_D ||
	     WILL_FIRE_RL_doFEQ_D ||
	     WILL_FIRE_RL_doFLT_D ||
	     WILL_FIRE_RL_doFLE_D ||
	     WILL_FIRE_RL_doFCLASS_D ||
	     WILL_FIRE_RL_rl_get_fpu_result ;
  // register stateR
  always@(EN_req or
	  WILL_FIRE_RL_rl_get_fpu_result or
	  WILL_FIRE_RL_doFCLASS_D or
	  WILL_FIRE_RL_doFMV_X_D or
	  WILL_FIRE_RL_doFMV_D_X or
	  WILL_FIRE_RL_doFLE_D or
	  WILL_FIRE_RL_doFLT_D or
	  WILL_FIRE_RL_doFEQ_D or
	  WILL_FIRE_RL_doFMAX_D or
	  WILL_FIRE_RL_doFMIN_D or
	  WILL_FIRE_RL_doFCVT_D_S or
	  WILL_FIRE_RL_doFCVT_S_D or
	  WILL_FIRE_RL_doFCVT_LU_D or
	  WILL_FIRE_RL_doFCVT_L_D or
	  WILL_FIRE_RL_doFCVT_D_LU or
	  WILL_FIRE_RL_doFCVT_D_L or
	  WILL_FIRE_RL_doFCVT_WU_D or
	  WILL_FIRE_RL_doFCVT_W_D or
	  WILL_FIRE_RL_doFCVT_D_WU or
	  WILL_FIRE_RL_doFCVT_D_W or
	  WILL_FIRE_RL_doFSGNJX_D or
	  WILL_FIRE_RL_doFSGNJN_D or
	  WILL_FIRE_RL_doFSGNJ_D or
	  WILL_FIRE_RL_doFNMSUB_D or
	  WILL_FIRE_RL_doFNMADD_D or
	  WILL_FIRE_RL_doFMSUB_D or
	  WILL_FIRE_RL_doFMADD_D or
	  WILL_FIRE_RL_doFMUL_D or
	  WILL_FIRE_RL_doFSUB_D or
	  WILL_FIRE_RL_doFADD_D or
	  WILL_FIRE_RL_doFCLASS_S or
	  WILL_FIRE_RL_doFLE_S or
	  WILL_FIRE_RL_doFLT_S or
	  WILL_FIRE_RL_doFEQ_S or
	  WILL_FIRE_RL_doFMV_X_W or
	  WILL_FIRE_RL_doFMV_W_X or
	  WILL_FIRE_RL_doFMAX_S or
	  WILL_FIRE_RL_doFMIN_S or
	  WILL_FIRE_RL_doFCVT_WU_S or
	  WILL_FIRE_RL_doFCVT_W_S or
	  WILL_FIRE_RL_doFCVT_LU_S or
	  WILL_FIRE_RL_doFCVT_L_S or
	  WILL_FIRE_RL_doFCVT_S_WU or
	  WILL_FIRE_RL_doFCVT_S_W or
	  WILL_FIRE_RL_doFCVT_S_LU or
	  WILL_FIRE_RL_doFCVT_S_L or
	  WILL_FIRE_RL_doFSGNJX_S or
	  WILL_FIRE_RL_doFSGNJN_S or
	  WILL_FIRE_RL_doFSGNJ_S or
	  WILL_FIRE_RL_doFNMSUB_S or
	  WILL_FIRE_RL_doFNMADD_S or
	  WILL_FIRE_RL_doFMSUB_S or
	  WILL_FIRE_RL_doFMADD_S or
	  WILL_FIRE_RL_doFMUL_S or
	  WILL_FIRE_RL_doFSUB_S or WILL_FIRE_RL_doFADD_S)
  case (1'b1)
    EN_req: stateR$D_IN = 2'd0;
    WILL_FIRE_RL_rl_get_fpu_result || WILL_FIRE_RL_doFCLASS_D ||
    WILL_FIRE_RL_doFMV_X_D ||
    WILL_FIRE_RL_doFMV_D_X ||
    WILL_FIRE_RL_doFLE_D ||
    WILL_FIRE_RL_doFLT_D ||
    WILL_FIRE_RL_doFEQ_D ||
    WILL_FIRE_RL_doFMAX_D ||
    WILL_FIRE_RL_doFMIN_D ||
    WILL_FIRE_RL_doFCVT_D_S ||
    WILL_FIRE_RL_doFCVT_S_D ||
    WILL_FIRE_RL_doFCVT_LU_D ||
    WILL_FIRE_RL_doFCVT_L_D ||
    WILL_FIRE_RL_doFCVT_D_LU ||
    WILL_FIRE_RL_doFCVT_D_L ||
    WILL_FIRE_RL_doFCVT_WU_D ||
    WILL_FIRE_RL_doFCVT_W_D ||
    WILL_FIRE_RL_doFCVT_D_WU ||
    WILL_FIRE_RL_doFCVT_D_W ||
    WILL_FIRE_RL_doFSGNJX_D ||
    WILL_FIRE_RL_doFSGNJN_D ||
    WILL_FIRE_RL_doFSGNJ_D:
	stateR$D_IN = 2'd2;
    WILL_FIRE_RL_doFNMSUB_D || WILL_FIRE_RL_doFNMADD_D ||
    WILL_FIRE_RL_doFMSUB_D ||
    WILL_FIRE_RL_doFMADD_D ||
    WILL_FIRE_RL_doFMUL_D ||
    WILL_FIRE_RL_doFSUB_D ||
    WILL_FIRE_RL_doFADD_D:
	stateR$D_IN = 2'd1;
    WILL_FIRE_RL_doFCLASS_S || WILL_FIRE_RL_doFLE_S || WILL_FIRE_RL_doFLT_S ||
    WILL_FIRE_RL_doFEQ_S ||
    WILL_FIRE_RL_doFMV_X_W ||
    WILL_FIRE_RL_doFMV_W_X ||
    WILL_FIRE_RL_doFMAX_S ||
    WILL_FIRE_RL_doFMIN_S ||
    WILL_FIRE_RL_doFCVT_WU_S ||
    WILL_FIRE_RL_doFCVT_W_S ||
    WILL_FIRE_RL_doFCVT_LU_S ||
    WILL_FIRE_RL_doFCVT_L_S ||
    WILL_FIRE_RL_doFCVT_S_WU ||
    WILL_FIRE_RL_doFCVT_S_W ||
    WILL_FIRE_RL_doFCVT_S_LU ||
    WILL_FIRE_RL_doFCVT_S_L ||
    WILL_FIRE_RL_doFSGNJX_S ||
    WILL_FIRE_RL_doFSGNJN_S ||
    WILL_FIRE_RL_doFSGNJ_S:
	stateR$D_IN = 2'd2;
    WILL_FIRE_RL_doFNMSUB_S || WILL_FIRE_RL_doFNMADD_S ||
    WILL_FIRE_RL_doFMSUB_S ||
    WILL_FIRE_RL_doFMADD_S ||
    WILL_FIRE_RL_doFMUL_S ||
    WILL_FIRE_RL_doFSUB_S ||
    WILL_FIRE_RL_doFADD_S:
	stateR$D_IN = 2'd1;
    default: stateR$D_IN = 2'b10 /* unspecified value */ ;
  endcase
  assign stateR$EN =
	     EN_req || WILL_FIRE_RL_doFNMSUB_D || WILL_FIRE_RL_doFNMADD_D ||
	     WILL_FIRE_RL_doFMSUB_D ||
	     WILL_FIRE_RL_doFMADD_D ||
	     WILL_FIRE_RL_doFMUL_D ||
	     WILL_FIRE_RL_doFSUB_D ||
	     WILL_FIRE_RL_doFADD_D ||
	     WILL_FIRE_RL_doFNMSUB_S ||
	     WILL_FIRE_RL_doFNMADD_S ||
	     WILL_FIRE_RL_doFMSUB_S ||
	     WILL_FIRE_RL_doFMADD_S ||
	     WILL_FIRE_RL_doFMUL_S ||
	     WILL_FIRE_RL_doFSUB_S ||
	     WILL_FIRE_RL_doFADD_S ||
	     WILL_FIRE_RL_rl_get_fpu_result ||
	     WILL_FIRE_RL_doFCLASS_D ||
	     WILL_FIRE_RL_doFMV_X_D ||
	     WILL_FIRE_RL_doFMV_D_X ||
	     WILL_FIRE_RL_doFLE_D ||
	     WILL_FIRE_RL_doFLT_D ||
	     WILL_FIRE_RL_doFEQ_D ||
	     WILL_FIRE_RL_doFMAX_D ||
	     WILL_FIRE_RL_doFMIN_D ||
	     WILL_FIRE_RL_doFCVT_D_S ||
	     WILL_FIRE_RL_doFCVT_S_D ||
	     WILL_FIRE_RL_doFCVT_LU_D ||
	     WILL_FIRE_RL_doFCVT_L_D ||
	     WILL_FIRE_RL_doFCVT_D_LU ||
	     WILL_FIRE_RL_doFCVT_D_L ||
	     WILL_FIRE_RL_doFCVT_WU_D ||
	     WILL_FIRE_RL_doFCVT_W_D ||
	     WILL_FIRE_RL_doFCVT_D_WU ||
	     WILL_FIRE_RL_doFCVT_D_W ||
	     WILL_FIRE_RL_doFSGNJX_D ||
	     WILL_FIRE_RL_doFSGNJN_D ||
	     WILL_FIRE_RL_doFSGNJ_D ||
	     WILL_FIRE_RL_doFCLASS_S ||
	     WILL_FIRE_RL_doFLE_S ||
	     WILL_FIRE_RL_doFLT_S ||
	     WILL_FIRE_RL_doFEQ_S ||
	     WILL_FIRE_RL_doFMV_X_W ||
	     WILL_FIRE_RL_doFMV_W_X ||
	     WILL_FIRE_RL_doFMAX_S ||
	     WILL_FIRE_RL_doFMIN_S ||
	     WILL_FIRE_RL_doFCVT_WU_S ||
	     WILL_FIRE_RL_doFCVT_W_S ||
	     WILL_FIRE_RL_doFCVT_LU_S ||
	     WILL_FIRE_RL_doFCVT_L_S ||
	     WILL_FIRE_RL_doFCVT_S_WU ||
	     WILL_FIRE_RL_doFCVT_S_W ||
	     WILL_FIRE_RL_doFCVT_S_LU ||
	     WILL_FIRE_RL_doFCVT_S_L ||
	     WILL_FIRE_RL_doFSGNJX_S ||
	     WILL_FIRE_RL_doFSGNJN_S ||
	     WILL_FIRE_RL_doFSGNJ_S ;
  // submodule fpu
  always@(WILL_FIRE_RL_doFADD_S or
	  MUX_fpu$request_put_1__VAL_1 or
	  WILL_FIRE_RL_doFSUB_S or
	  MUX_fpu$request_put_1__VAL_2 or
	  WILL_FIRE_RL_doFMUL_S or
	  MUX_fpu$request_put_1__VAL_3 or
	  WILL_FIRE_RL_doFMADD_S or
	  MUX_fpu$request_put_1__VAL_4 or
	  WILL_FIRE_RL_doFMSUB_S or
	  MUX_fpu$request_put_1__VAL_5 or
	  WILL_FIRE_RL_doFNMADD_S or
	  MUX_fpu$request_put_1__VAL_6 or
	  WILL_FIRE_RL_doFNMSUB_S or
	  MUX_fpu$request_put_1__VAL_7 or
	  WILL_FIRE_RL_doFADD_D or
	  MUX_fpu$request_put_1__VAL_8 or
	  WILL_FIRE_RL_doFSUB_D or
	  MUX_fpu$request_put_1__VAL_9 or
	  WILL_FIRE_RL_doFMUL_D or
	  MUX_fpu$request_put_1__VAL_10 or
	  WILL_FIRE_RL_doFMADD_D or
	  MUX_fpu$request_put_1__VAL_11 or
	  WILL_FIRE_RL_doFMSUB_D or
	  MUX_fpu$request_put_1__VAL_12 or
	  WILL_FIRE_RL_doFNMADD_D or
	  MUX_fpu$request_put_1__VAL_13 or
	  WILL_FIRE_RL_doFNMSUB_D or MUX_fpu$request_put_1__VAL_14)
  begin
    case (1'b1) // synopsys parallel_case
      WILL_FIRE_RL_doFADD_S: fpu$request_put = MUX_fpu$request_put_1__VAL_1;
      WILL_FIRE_RL_doFSUB_S: fpu$request_put = MUX_fpu$request_put_1__VAL_2;
      WILL_FIRE_RL_doFMUL_S: fpu$request_put = MUX_fpu$request_put_1__VAL_3;
      WILL_FIRE_RL_doFMADD_S: fpu$request_put = MUX_fpu$request_put_1__VAL_4;
      WILL_FIRE_RL_doFMSUB_S: fpu$request_put = MUX_fpu$request_put_1__VAL_5;
      WILL_FIRE_RL_doFNMADD_S: fpu$request_put = MUX_fpu$request_put_1__VAL_6;
      WILL_FIRE_RL_doFNMSUB_S: fpu$request_put = MUX_fpu$request_put_1__VAL_7;
      WILL_FIRE_RL_doFADD_D: fpu$request_put = MUX_fpu$request_put_1__VAL_8;
      WILL_FIRE_RL_doFSUB_D: fpu$request_put = MUX_fpu$request_put_1__VAL_9;
      WILL_FIRE_RL_doFMUL_D: fpu$request_put = MUX_fpu$request_put_1__VAL_10;
      WILL_FIRE_RL_doFMADD_D: fpu$request_put = MUX_fpu$request_put_1__VAL_11;
      WILL_FIRE_RL_doFMSUB_D: fpu$request_put = MUX_fpu$request_put_1__VAL_12;
      WILL_FIRE_RL_doFNMADD_D:
	  fpu$request_put = MUX_fpu$request_put_1__VAL_13;
      WILL_FIRE_RL_doFNMSUB_D:
	  fpu$request_put = MUX_fpu$request_put_1__VAL_14;
      default: fpu$request_put =
		   202'h2AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA /* unspecified value */ ;
    endcase
  end
  assign fpu$EN_request_put =
	     WILL_FIRE_RL_doFADD_S || WILL_FIRE_RL_doFSUB_S ||
	     WILL_FIRE_RL_doFMUL_S ||
	     WILL_FIRE_RL_doFMADD_S ||
	     WILL_FIRE_RL_doFMSUB_S ||
	     WILL_FIRE_RL_doFNMADD_S ||
	     WILL_FIRE_RL_doFNMSUB_S ||
	     WILL_FIRE_RL_doFADD_D ||
	     WILL_FIRE_RL_doFSUB_D ||
	     WILL_FIRE_RL_doFMUL_D ||
	     WILL_FIRE_RL_doFMADD_D ||
	     WILL_FIRE_RL_doFMSUB_D ||
	     WILL_FIRE_RL_doFNMADD_D ||
	     WILL_FIRE_RL_doFNMSUB_D ;
  assign fpu$EN_response_get = CAN_FIRE_RL_rl_get_fpu_result ;
  // submodule frmFpuF
  assign frmFpuF$D_IN = 1'b0 ;
  assign frmFpuF$ENQ = 1'b0 ;
  assign frmFpuF$DEQ = 1'b0 ;
  assign frmFpuF$CLR = 1'b0 ;
  // remaining internal signals
  assign IF_0_CONCAT_IF_IF_0b0_CONCAT_NOT_requestR_BITS_ETC__q114 =
	     _0_CONCAT_IF_IF_0b0_CONCAT_NOT_requestR_BITS_19_ETC___d3539 ?
	       _theResult___snd__h119527 :
	       _theResult____h111357 ;
  assign IF_0_CONCAT_IF_IF_3074_MINUS_SEXT_IF_requestR__ETC__q151 =
	     _0_CONCAT_IF_IF_3074_MINUS_SEXT_IF_requestR_BIT_ETC___d4817 ?
	       _theResult___snd__h178715 :
	       _theResult____h170416 ;
  assign IF_0_CONCAT_IF_IF_3970_MINUS_SEXT_requestR_BIT_ETC__q119 =
	     _0_CONCAT_IF_IF_3970_MINUS_SEXT_requestR_BITS_1_ETC___d3983 ?
	       _theResult___snd__h137380 :
	       _theResult____h129081 ;
  assign IF_0_CONCAT_IF_IF_requestR_BITS_191_TO_160_4_E_ETC__q148 =
	     _0_CONCAT_IF_IF_requestR_BITS_191_TO_160_4_EQ_0_ETC___d4497 ?
	       _theResult___snd__h169068 :
	       57'd0 ;
  assign IF_0_CONCAT_IF_IF_requestR_BITS_191_TO_160_4_E_ETC__q154 =
	     _0_CONCAT_IF_IF_requestR_BITS_191_TO_160_4_EQ_0_ETC___d4890 ?
	       _theResult___snd__h169068 :
	       _theResult___snd__h187467 ;
  assign IF_0_CONCAT_IF_requestR_BITS_190_TO_180_599_EQ_ETC__q116 =
	     _0_CONCAT_IF_requestR_BITS_190_TO_180_599_EQ_0__ETC___d3661 ?
	       _theResult___snd__h128139 :
	       57'd0 ;
  assign IF_0_CONCAT_IF_requestR_BITS_190_TO_180_599_EQ_ETC__q122 =
	     _0_CONCAT_IF_requestR_BITS_190_TO_180_599_EQ_0__ETC___d4056 ?
	       _theResult___snd__h128139 :
	       _theResult___snd__h146016 ;
  assign IF_3074_MINUS_0_CONCAT_IF_requestR_BIT_179_71__ETC___d4241 =
	     _3074_MINUS_0_CONCAT_IF_requestR_BIT_179_71_THE_ETC___d3305 ?
	       ((_theResult___fst_exp__h119464 == 8'd255) ?
		  requestR[191] :
		  ((requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
		    requestR[194:192] != 3'h3 &&
		    requestR[194:192] != 3'h4) ?
		     CASE_guard11367_0b0_requestR_BIT_191_0b1_reque_ETC__q140 :
		     CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q141)) :
	       ((_theResult___fst_exp__h128150 == 8'd255) ?
		  requestR[191] :
		  ((requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
		    requestR[194:192] != 3'h3 &&
		    requestR[194:192] != 3'h4) ?
		     CASE_guard20102_0b0_requestR_BIT_191_0b1_reque_ETC__q142 :
		     CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q143)) ;
  assign IF_32_MINUS_0_CONCAT_IF_IF_requestR_BIT_159_6__ETC___d1313 =
	     _32_MINUS_0_CONCAT_IF_IF_requestR_BIT_159_6_THE_ETC___d1261 ?
	       ((requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
		 requestR[194:192] != 3'h3 &&
		 requestR[194:192] != 3'h4) ?
		  CASE_guard8894_0b0_requestR_BIT_159_0b1_reques_ETC__q40 :
		  CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q41) :
	       ((x__h29436[7:0] == 8'd255) ?
		  requestR[159] :
		  ((requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
		    requestR[194:192] != 3'h3 &&
		    requestR[194:192] != 3'h4) ?
		     CASE_guard9421_0b0_requestR_BIT_159_0b1_reques_ETC__q42 :
		     CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q43)) ;
  assign IF_32_MINUS_0_CONCAT_IF_IF_requestR_BIT_159_6__ETC___d1463 =
	     _32_MINUS_0_CONCAT_IF_IF_requestR_BIT_159_6_THE_ETC___d1261 ?
	       guard__h28894 != 2'b0 :
	       x__h29436[7:0] != 8'd255 && guard__h29421 != 2'b0 ;
  assign IF_32_MINUS_0_CONCAT_IF_IF_requestR_BIT_159_6__ETC___d2289 =
	     _32_MINUS_0_CONCAT_IF_IF_requestR_BIT_159_6_THE_ETC___d2238 ?
	       ((requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
		 requestR[194:192] != 3'h3 &&
		 requestR[194:192] != 3'h4) ?
		  CASE_guard0287_0b0_requestR_BIT_159_0b1_reques_ETC__q69 :
		  CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q70) :
	       ((x__h61032[10:0] == 11'd2047) ?
		  requestR[159] :
		  ((requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
		    requestR[194:192] != 3'h3 &&
		    requestR[194:192] != 3'h4) ?
		     CASE_guard1017_0b0_requestR_BIT_159_0b1_reques_ETC__q71 :
		     CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q72)) ;
  assign IF_32_MINUS_0_CONCAT_IF_IF_requestR_BIT_159_6__ETC___d2404 =
	     _32_MINUS_0_CONCAT_IF_IF_requestR_BIT_159_6_THE_ETC___d2238 ?
	       guard__h60287 != 2'b0 :
	       x__h61032[10:0] != 11'd2047 && guard__h61017 != 2'b0 ;
  assign IF_32_MINUS_0_CONCAT_IF_requestR_BIT_159_6_THE_ETC___d1651 =
	     _32_MINUS_0_CONCAT_IF_requestR_BIT_159_6_THEN_0_ETC___d1513 ?
	       guard__h35065 != 2'b0 :
	       x__h35606[7:0] != 8'd255 && guard__h35591 != 2'b0 ;
  assign IF_32_MINUS_0_CONCAT_IF_requestR_BIT_159_6_THE_ETC___d2587 =
	     _32_MINUS_0_CONCAT_IF_requestR_BIT_159_6_THEN_0_ETC___d2451 ?
	       guard__h69983 != 2'b0 :
	       x__h70727[10:0] != 11'd2047 && guard__h70712 != 2'b0 ;
  assign IF_64_MINUS_0_CONCAT_IF_IF_requestR_BIT_191_27_ETC___d2824 =
	     _64_MINUS_0_CONCAT_IF_IF_requestR_BIT_191_27_TH_ETC___d2775 ?
	       ((requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
		 requestR[194:192] != 3'h3 &&
		 requestR[194:192] != 3'h4) ?
		  CASE_guard3828_0b0_requestR_BIT_191_0b1_reques_ETC__q94 :
		  CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q95) :
	       ((x__h84573[10:0] == 11'd2047) ?
		  requestR[191] :
		  ((requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
		    requestR[194:192] != 3'h3 &&
		    requestR[194:192] != 3'h4) ?
		     CASE_guard4558_0b0_requestR_BIT_191_0b1_reques_ETC__q96 :
		     CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q97)) ;
  assign IF_64_MINUS_0_CONCAT_IF_IF_requestR_BIT_191_27_ETC___d2941 =
	     _64_MINUS_0_CONCAT_IF_IF_requestR_BIT_191_27_TH_ETC___d2775 ?
	       guard__h83828 != 2'b0 :
	       x__h84573[10:0] != 11'd2047 && guard__h84558 != 2'b0 ;
  assign IF_64_MINUS_0_CONCAT_IF_IF_requestR_BIT_191_27_ETC___d454 =
	     _64_MINUS_0_CONCAT_IF_IF_requestR_BIT_191_27_TH_ETC___d393 ?
	       ((requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
		 requestR[194:192] != 3'h3 &&
		 requestR[194:192] != 3'h4) ?
		  CASE_guard1845_0b0_requestR_BIT_191_0b1_reques_ETC__q10 :
		  CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q11) :
	       ((x__h12390[7:0] == 8'd255) ?
		  requestR[191] :
		  ((requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
		    requestR[194:192] != 3'h3 &&
		    requestR[194:192] != 3'h4) ?
		     CASE_guard2375_0b0_requestR_BIT_191_0b1_reques_ETC__q12 :
		     CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q13)) ;
  assign IF_64_MINUS_0_CONCAT_IF_IF_requestR_BIT_191_27_ETC___d636 =
	     _64_MINUS_0_CONCAT_IF_IF_requestR_BIT_191_27_TH_ETC___d393 ?
	       guard__h11845 != 2'b0 :
	       x__h12390[7:0] != 8'd255 && guard__h12375 != 2'b0 ;
  assign IF_64_MINUS_0_CONCAT_IF_requestR_BIT_191_27_TH_ETC___d1109 =
	     _64_MINUS_0_CONCAT_IF_requestR_BIT_191_27_THEN__ETC___d907 ?
	       guard__h22467 != 2'b0 :
	       x__h23008[7:0] != 8'd255 && guard__h22993 != 2'b0 ;
  assign IF_64_MINUS_0_CONCAT_IF_requestR_BIT_191_27_TH_ETC___d3094 =
	     _64_MINUS_0_CONCAT_IF_requestR_BIT_191_27_THEN__ETC___d2957 ?
	       guard__h94840 != 2'b0 :
	       x__h95584[10:0] != 11'd2047 && guard__h95569 != 2'b0 ;
  assign IF_IF_0b0_CONCAT_NOT_requestR_BITS_190_TO_180__ETC___d3537 =
	     (_theResult____h111357[56] ?
		6'd0 :
		(_theResult____h111357[55] ?
		   6'd1 :
		   (_theResult____h111357[54] ?
		      6'd2 :
		      (_theResult____h111357[53] ?
			 6'd3 :
			 (_theResult____h111357[52] ?
			    6'd4 :
			    (_theResult____h111357[51] ?
			       6'd5 :
			       (_theResult____h111357[50] ?
				  6'd6 :
				  (_theResult____h111357[49] ?
				     6'd7 :
				     (_theResult____h111357[48] ?
					6'd8 :
					(_theResult____h111357[47] ?
					   6'd9 :
					   (_theResult____h111357[46] ?
					      6'd10 :
					      (_theResult____h111357[45] ?
						 6'd11 :
						 (_theResult____h111357[44] ?
						    6'd12 :
						    (_theResult____h111357[43] ?
						       6'd13 :
						       (_theResult____h111357[42] ?
							  6'd14 :
							  (_theResult____h111357[41] ?
							     6'd15 :
							     (_theResult____h111357[40] ?
								6'd16 :
								(_theResult____h111357[39] ?
								   6'd17 :
								   (_theResult____h111357[38] ?
								      6'd18 :
								      (_theResult____h111357[37] ?
									 6'd19 :
									 (_theResult____h111357[36] ?
									    6'd20 :
									    (_theResult____h111357[35] ?
									       6'd21 :
									       (_theResult____h111357[34] ?
										  6'd22 :
										  (_theResult____h111357[33] ?
										     6'd23 :
										     (_theResult____h111357[32] ?
											6'd24 :
											(_theResult____h111357[31] ?
											   6'd25 :
											   (_theResult____h111357[30] ?
											      6'd26 :
											      (_theResult____h111357[29] ?
												 6'd27 :
												 (_theResult____h111357[28] ?
												    6'd28 :
												    (_theResult____h111357[27] ?
												       6'd29 :
												       (_theResult____h111357[26] ?
													  6'd30 :
													  (_theResult____h111357[25] ?
													     6'd31 :
													     (_theResult____h111357[24] ?
														6'd32 :
														(_theResult____h111357[23] ?
														   6'd33 :
														   (_theResult____h111357[22] ?
														      6'd34 :
														      (_theResult____h111357[21] ?
															 6'd35 :
															 (_theResult____h111357[20] ?
															    6'd36 :
															    (_theResult____h111357[19] ?
															       6'd37 :
															       (_theResult____h111357[18] ?
																  6'd38 :
																  (_theResult____h111357[17] ?
																     6'd39 :
																     (_theResult____h111357[16] ?
																	6'd40 :
																	(_theResult____h111357[15] ?
																	   6'd41 :
																	   (_theResult____h111357[14] ?
																	      6'd42 :
																	      (_theResult____h111357[13] ?
																		 6'd43 :
																		 (_theResult____h111357[12] ?
																		    6'd44 :
																		    (_theResult____h111357[11] ?
																		       6'd45 :
																		       (_theResult____h111357[10] ?
																			  6'd46 :
																			  (_theResult____h111357[9] ?
																			     6'd47 :
																			     (_theResult____h111357[8] ?
																				6'd48 :
																				(_theResult____h111357[7] ?
																				   6'd49 :
																				   (_theResult____h111357[6] ?
																				      6'd50 :
																				      (_theResult____h111357[5] ?
																					 6'd51 :
																					 (_theResult____h111357[4] ?
																					    6'd52 :
																					    (_theResult____h111357[3] ?
																					       6'd53 :
																					       (_theResult____h111357[2] ?
																						  6'd54 :
																						  (_theResult____h111357[1] ?
																						     6'd55 :
																						     (_theResult____h111357[0] ?
																							6'd56 :
																							6'd57))))))))))))))))))))))))))))))))))))))))))))))))))))))))) -
	     6'd1 ;
  assign IF_IF_3074_MINUS_SEXT_IF_requestR_BITS_191_TO__ETC___d4815 =
	     (_theResult____h170416[56] ?
		6'd0 :
		(_theResult____h170416[55] ?
		   6'd1 :
		   (_theResult____h170416[54] ?
		      6'd2 :
		      (_theResult____h170416[53] ?
			 6'd3 :
			 (_theResult____h170416[52] ?
			    6'd4 :
			    (_theResult____h170416[51] ?
			       6'd5 :
			       (_theResult____h170416[50] ?
				  6'd6 :
				  (_theResult____h170416[49] ?
				     6'd7 :
				     (_theResult____h170416[48] ?
					6'd8 :
					(_theResult____h170416[47] ?
					   6'd9 :
					   (_theResult____h170416[46] ?
					      6'd10 :
					      (_theResult____h170416[45] ?
						 6'd11 :
						 (_theResult____h170416[44] ?
						    6'd12 :
						    (_theResult____h170416[43] ?
						       6'd13 :
						       (_theResult____h170416[42] ?
							  6'd14 :
							  (_theResult____h170416[41] ?
							     6'd15 :
							     (_theResult____h170416[40] ?
								6'd16 :
								(_theResult____h170416[39] ?
								   6'd17 :
								   (_theResult____h170416[38] ?
								      6'd18 :
								      (_theResult____h170416[37] ?
									 6'd19 :
									 (_theResult____h170416[36] ?
									    6'd20 :
									    (_theResult____h170416[35] ?
									       6'd21 :
									       (_theResult____h170416[34] ?
										  6'd22 :
										  (_theResult____h170416[33] ?
										     6'd23 :
										     (_theResult____h170416[32] ?
											6'd24 :
											(_theResult____h170416[31] ?
											   6'd25 :
											   (_theResult____h170416[30] ?
											      6'd26 :
											      (_theResult____h170416[29] ?
												 6'd27 :
												 (_theResult____h170416[28] ?
												    6'd28 :
												    (_theResult____h170416[27] ?
												       6'd29 :
												       (_theResult____h170416[26] ?
													  6'd30 :
													  (_theResult____h170416[25] ?
													     6'd31 :
													     (_theResult____h170416[24] ?
														6'd32 :
														(_theResult____h170416[23] ?
														   6'd33 :
														   (_theResult____h170416[22] ?
														      6'd34 :
														      (_theResult____h170416[21] ?
															 6'd35 :
															 (_theResult____h170416[20] ?
															    6'd36 :
															    (_theResult____h170416[19] ?
															       6'd37 :
															       (_theResult____h170416[18] ?
																  6'd38 :
																  (_theResult____h170416[17] ?
																     6'd39 :
																     (_theResult____h170416[16] ?
																	6'd40 :
																	(_theResult____h170416[15] ?
																	   6'd41 :
																	   (_theResult____h170416[14] ?
																	      6'd42 :
																	      (_theResult____h170416[13] ?
																		 6'd43 :
																		 (_theResult____h170416[12] ?
																		    6'd44 :
																		    (_theResult____h170416[11] ?
																		       6'd45 :
																		       (_theResult____h170416[10] ?
																			  6'd46 :
																			  (_theResult____h170416[9] ?
																			     6'd47 :
																			     (_theResult____h170416[8] ?
																				6'd48 :
																				(_theResult____h170416[7] ?
																				   6'd49 :
																				   (_theResult____h170416[6] ?
																				      6'd50 :
																				      (_theResult____h170416[5] ?
																					 6'd51 :
																					 (_theResult____h170416[4] ?
																					    6'd52 :
																					    (_theResult____h170416[3] ?
																					       6'd53 :
																					       (_theResult____h170416[2] ?
																						  6'd54 :
																						  (_theResult____h170416[1] ?
																						     6'd55 :
																						     (_theResult____h170416[0] ?
																							6'd56 :
																							6'd57))))))))))))))))))))))))))))))))))))))))))))))))))))))))) -
	     6'd1 ;
  assign IF_IF_3970_MINUS_SEXT_requestR_BITS_190_TO_180_ETC___d3981 =
	     (_theResult____h129081[56] ?
		6'd0 :
		(_theResult____h129081[55] ?
		   6'd1 :
		   (_theResult____h129081[54] ?
		      6'd2 :
		      (_theResult____h129081[53] ?
			 6'd3 :
			 (_theResult____h129081[52] ?
			    6'd4 :
			    (_theResult____h129081[51] ?
			       6'd5 :
			       (_theResult____h129081[50] ?
				  6'd6 :
				  (_theResult____h129081[49] ?
				     6'd7 :
				     (_theResult____h129081[48] ?
					6'd8 :
					(_theResult____h129081[47] ?
					   6'd9 :
					   (_theResult____h129081[46] ?
					      6'd10 :
					      (_theResult____h129081[45] ?
						 6'd11 :
						 (_theResult____h129081[44] ?
						    6'd12 :
						    (_theResult____h129081[43] ?
						       6'd13 :
						       (_theResult____h129081[42] ?
							  6'd14 :
							  (_theResult____h129081[41] ?
							     6'd15 :
							     (_theResult____h129081[40] ?
								6'd16 :
								(_theResult____h129081[39] ?
								   6'd17 :
								   (_theResult____h129081[38] ?
								      6'd18 :
								      (_theResult____h129081[37] ?
									 6'd19 :
									 (_theResult____h129081[36] ?
									    6'd20 :
									    (_theResult____h129081[35] ?
									       6'd21 :
									       (_theResult____h129081[34] ?
										  6'd22 :
										  (_theResult____h129081[33] ?
										     6'd23 :
										     (_theResult____h129081[32] ?
											6'd24 :
											(_theResult____h129081[31] ?
											   6'd25 :
											   (_theResult____h129081[30] ?
											      6'd26 :
											      (_theResult____h129081[29] ?
												 6'd27 :
												 (_theResult____h129081[28] ?
												    6'd28 :
												    (_theResult____h129081[27] ?
												       6'd29 :
												       (_theResult____h129081[26] ?
													  6'd30 :
													  (_theResult____h129081[25] ?
													     6'd31 :
													     (_theResult____h129081[24] ?
														6'd32 :
														(_theResult____h129081[23] ?
														   6'd33 :
														   (_theResult____h129081[22] ?
														      6'd34 :
														      (_theResult____h129081[21] ?
															 6'd35 :
															 (_theResult____h129081[20] ?
															    6'd36 :
															    (_theResult____h129081[19] ?
															       6'd37 :
															       (_theResult____h129081[18] ?
																  6'd38 :
																  (_theResult____h129081[17] ?
																     6'd39 :
																     (_theResult____h129081[16] ?
																	6'd40 :
																	(_theResult____h129081[15] ?
																	   6'd41 :
																	   (_theResult____h129081[14] ?
																	      6'd42 :
																	      (_theResult____h129081[13] ?
																		 6'd43 :
																		 (_theResult____h129081[12] ?
																		    6'd44 :
																		    (_theResult____h129081[11] ?
																		       6'd45 :
																		       (_theResult____h129081[10] ?
																			  6'd46 :
																			  (_theResult____h129081[9] ?
																			     6'd47 :
																			     (_theResult____h129081[8] ?
																				6'd48 :
																				(_theResult____h129081[7] ?
																				   6'd49 :
																				   (_theResult____h129081[6] ?
																				      6'd50 :
																				      (_theResult____h129081[5] ?
																					 6'd51 :
																					 (_theResult____h129081[4] ?
																					    6'd52 :
																					    (_theResult____h129081[3] ?
																					       6'd53 :
																					       (_theResult____h129081[2] ?
																						  6'd54 :
																						  (_theResult____h129081[1] ?
																						     6'd55 :
																						     (_theResult____h129081[0] ?
																							6'd56 :
																							6'd57))))))))))))))))))))))))))))))))))))))))))))))))))))))))) -
	     6'd1 ;
  assign IF_IF_IF_3074_MINUS_SEXT_IF_requestR_BITS_191__ETC___d5059 =
	     (_theResult___fst_exp__h178652 == 11'd2047) ?
	       requestR[191:160] == 32'hFFFFFFFF && requestR[159] :
	       ((requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
		 requestR[194:192] != 3'h3 &&
		 requestR[194:192] != 3'h4) ?
		  CASE_guard70426_0b0_requestR_BITS_191_TO_160_E_ETC__q164 :
		  CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q165) ;
  assign IF_IF_IF_IF_0b0_CONCAT_NOT_requestR_BITS_190_T_ETC___d3596 =
	     (guard__h111367 == 2'b0 || requestR[191]) ?
	       _theResult___fst_exp__h119464 :
	       _theResult___exp__h119990 ;
  assign IF_IF_IF_IF_0b0_CONCAT_NOT_requestR_BITS_190_T_ETC___d3598 =
	     (guard__h111367 == 2'b0) ?
	       _theResult___fst_exp__h119464 :
	       (requestR[191] ?
		  _theResult___exp__h119990 :
		  _theResult___fst_exp__h119464) ;
  assign IF_IF_IF_IF_0b0_CONCAT_NOT_requestR_BITS_190_T_ETC___d4143 =
	     (guard__h111367 == 2'b0 || requestR[191]) ?
	       sfdin__h119458[56:34] :
	       _theResult___sfd__h119991 ;
  assign IF_IF_IF_IF_0b0_CONCAT_NOT_requestR_BITS_190_T_ETC___d4145 =
	     (guard__h111367 == 2'b0) ?
	       sfdin__h119458[56:34] :
	       (requestR[191] ?
		  _theResult___sfd__h119991 :
		  sfdin__h119458[56:34]) ;
  assign IF_IF_IF_IF_3074_MINUS_SEXT_IF_requestR_BITS_1_ETC___d4874 =
	     (guard__h170426 == 2'b0 ||
	      requestR[191:160] == 32'hFFFFFFFF && requestR[159]) ?
	       _theResult___fst_exp__h178652 :
	       _theResult___exp__h179381 ;
  assign IF_IF_IF_IF_3074_MINUS_SEXT_IF_requestR_BITS_1_ETC___d4876 =
	     (guard__h170426 == 2'b0) ?
	       _theResult___fst_exp__h178652 :
	       ((requestR[191:160] == 32'hFFFFFFFF && requestR[159]) ?
		  _theResult___exp__h179381 :
		  _theResult___fst_exp__h178652) ;
  assign IF_IF_IF_IF_3074_MINUS_SEXT_IF_requestR_BITS_1_ETC___d5003 =
	     (guard__h170426 == 2'b0 ||
	      requestR[191:160] == 32'hFFFFFFFF && requestR[159]) ?
	       sfdin__h178646[56:5] :
	       _theResult___sfd__h179382 ;
  assign IF_IF_IF_IF_3074_MINUS_SEXT_IF_requestR_BITS_1_ETC___d5005 =
	     (guard__h170426 == 2'b0) ?
	       sfdin__h178646[56:5] :
	       ((requestR[191:160] == 32'hFFFFFFFF && requestR[159]) ?
		  _theResult___sfd__h179382 :
		  sfdin__h178646[56:5]) ;
  assign IF_IF_IF_IF_3970_MINUS_SEXT_requestR_BITS_190__ETC___d4040 =
	     (guard__h129091 == 2'b0 || requestR[191]) ?
	       _theResult___fst_exp__h137317 :
	       _theResult___exp__h137843 ;
  assign IF_IF_IF_IF_3970_MINUS_SEXT_requestR_BITS_190__ETC___d4042 =
	     (guard__h129091 == 2'b0) ?
	       _theResult___fst_exp__h137317 :
	       (requestR[191] ?
		  _theResult___exp__h137843 :
		  _theResult___fst_exp__h137317) ;
  assign IF_IF_IF_IF_3970_MINUS_SEXT_requestR_BITS_190__ETC___d4189 =
	     (guard__h129091 == 2'b0 || requestR[191]) ?
	       sfdin__h137311[56:34] :
	       _theResult___sfd__h137844 ;
  assign IF_IF_IF_IF_3970_MINUS_SEXT_requestR_BITS_190__ETC___d4191 =
	     (guard__h129091 == 2'b0) ?
	       sfdin__h137311[56:34] :
	       (requestR[191] ?
		  _theResult___sfd__h137844 :
		  sfdin__h137311[56:34]) ;
  assign IF_IF_IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFF_ETC___d4549 =
	     (guard__h161118 == 2'b0 ||
	      requestR[191:160] == 32'hFFFFFFFF && requestR[159]) ?
	       _theResult___fst_exp__h169079 :
	       _theResult___exp__h169734 ;
  assign IF_IF_IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFF_ETC___d4551 =
	     (guard__h161118 == 2'b0) ?
	       _theResult___fst_exp__h169079 :
	       ((requestR[191:160] == 32'hFFFFFFFF && requestR[159]) ?
		  _theResult___exp__h169734 :
		  _theResult___fst_exp__h169079) ;
  assign IF_IF_IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFF_ETC___d4943 =
	     (guard__h179493 == 2'b0 ||
	      requestR[191:160] == 32'hFFFFFFFF && requestR[159]) ?
	       _theResult___fst_exp__h187483 :
	       _theResult___exp__h188163 ;
  assign IF_IF_IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFF_ETC___d4945 =
	     (guard__h179493 == 2'b0) ?
	       _theResult___fst_exp__h187483 :
	       ((requestR[191:160] == 32'hFFFFFFFF && requestR[159]) ?
		  _theResult___exp__h188163 :
		  _theResult___fst_exp__h187483) ;
  assign IF_IF_IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFF_ETC___d4976 =
	     (guard__h161118 == 2'b0 ||
	      requestR[191:160] == 32'hFFFFFFFF && requestR[159]) ?
	       _theResult___snd__h169030[56:5] :
	       _theResult___sfd__h169735 ;
  assign IF_IF_IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFF_ETC___d4978 =
	     (guard__h161118 == 2'b0) ?
	       _theResult___snd__h169030[56:5] :
	       ((requestR[191:160] == 32'hFFFFFFFF && requestR[159]) ?
		  _theResult___sfd__h169735 :
		  _theResult___snd__h169030[56:5]) ;
  assign IF_IF_IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFF_ETC___d5022 =
	     (guard__h179493 == 2'b0 ||
	      requestR[191:160] == 32'hFFFFFFFF && requestR[159]) ?
	       _theResult___snd__h187429[56:5] :
	       _theResult___sfd__h188164 ;
  assign IF_IF_IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFF_ETC___d5024 =
	     (guard__h179493 == 2'b0) ?
	       _theResult___snd__h187429[56:5] :
	       ((requestR[191:160] == 32'hFFFFFFFF && requestR[159]) ?
		  _theResult___sfd__h188164 :
		  _theResult___snd__h187429[56:5]) ;
  assign IF_IF_IF_requestR_BITS_190_TO_180_599_EQ_0_609_ETC___d3713 =
	     (guard__h120102 == 2'b0 || requestR[191]) ?
	       _theResult___fst_exp__h128150 :
	       _theResult___exp__h128602 ;
  assign IF_IF_IF_requestR_BITS_190_TO_180_599_EQ_0_609_ETC___d3715 =
	     (guard__h120102 == 2'b0) ?
	       _theResult___fst_exp__h128150 :
	       (requestR[191] ?
		  _theResult___exp__h128602 :
		  _theResult___fst_exp__h128150) ;
  assign IF_IF_IF_requestR_BITS_190_TO_180_599_EQ_0_609_ETC___d4109 =
	     (guard__h137955 == 2'b0 || requestR[191]) ?
	       _theResult___fst_exp__h146032 :
	       _theResult___exp__h146509 ;
  assign IF_IF_IF_requestR_BITS_190_TO_180_599_EQ_0_609_ETC___d4111 =
	     (guard__h137955 == 2'b0) ?
	       _theResult___fst_exp__h146032 :
	       (requestR[191] ?
		  _theResult___exp__h146509 :
		  _theResult___fst_exp__h146032) ;
  assign IF_IF_IF_requestR_BITS_190_TO_180_599_EQ_0_609_ETC___d4162 =
	     (guard__h120102 == 2'b0 || requestR[191]) ?
	       _theResult___snd__h128101[56:34] :
	       _theResult___sfd__h128603 ;
  assign IF_IF_IF_requestR_BITS_190_TO_180_599_EQ_0_609_ETC___d4164 =
	     (guard__h120102 == 2'b0) ?
	       _theResult___snd__h128101[56:34] :
	       (requestR[191] ?
		  _theResult___sfd__h128603 :
		  _theResult___snd__h128101[56:34]) ;
  assign IF_IF_IF_requestR_BITS_190_TO_180_599_EQ_0_609_ETC___d4208 =
	     (guard__h137955 == 2'b0 || requestR[191]) ?
	       _theResult___snd__h145978[56:34] :
	       _theResult___sfd__h146510 ;
  assign IF_IF_IF_requestR_BITS_190_TO_180_599_EQ_0_609_ETC___d4210 =
	     (guard__h137955 == 2'b0) ?
	       _theResult___snd__h145978[56:34] :
	       (requestR[191] ?
		  _theResult___sfd__h146510 :
		  _theResult___snd__h145978[56:34]) ;
  assign IF_IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFF_ETC___d5067 =
	     (_theResult___fst_exp__h187483 == 11'd2047) ?
	       requestR[191:160] == 32'hFFFFFFFF && requestR[159] :
	       ((requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
		 requestR[194:192] != 3'h3 &&
		 requestR[194:192] != 3'h4) ?
		  CASE_guard79493_0b0_requestR_BITS_191_TO_160_E_ETC__q166 :
		  CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q167) ;
  assign IF_IF_IF_requestR_BIT_159_6_THEN_NEG_requestR__ETC___d1335 =
	     (guard__h28894 == 2'b0) ?
	       8'd0 :
	       (requestR[159] ? _theResult___exp__h29307 : 8'd0) ;
  assign IF_IF_IF_requestR_BIT_159_6_THEN_NEG_requestR__ETC___d1361 =
	     (guard__h29421 == 2'b0 || requestR[159]) ?
	       x__h29436[7:0] :
	       _theResult___exp__h29860 ;
  assign IF_IF_IF_requestR_BIT_159_6_THEN_NEG_requestR__ETC___d1363 =
	     (guard__h29421 == 2'b0) ?
	       x__h29436[7:0] :
	       (requestR[159] ? _theResult___exp__h29860 : x__h29436[7:0]) ;
  assign IF_IF_IF_requestR_BIT_159_6_THEN_NEG_requestR__ETC___d1384 =
	     (guard__h28894 == 2'b0 || requestR[159]) ?
	       sfd___3__h28884[31:9] :
	       _theResult___sfd__h29308 ;
  assign IF_IF_IF_requestR_BIT_159_6_THEN_NEG_requestR__ETC___d1386 =
	     (guard__h28894 == 2'b0) ?
	       sfd___3__h28884[31:9] :
	       (requestR[159] ?
		  _theResult___sfd__h29308 :
		  sfd___3__h28884[31:9]) ;
  assign IF_IF_IF_requestR_BIT_159_6_THEN_NEG_requestR__ETC___d1402 =
	     (guard__h29421 == 2'b0 || requestR[159]) ?
	       sfd___3__h28884[30:8] :
	       _theResult___sfd__h29861 ;
  assign IF_IF_IF_requestR_BIT_159_6_THEN_NEG_requestR__ETC___d1404 =
	     (guard__h29421 == 2'b0) ?
	       sfd___3__h28884[30:8] :
	       (requestR[159] ?
		  _theResult___sfd__h29861 :
		  sfd___3__h28884[30:8]) ;
  assign IF_IF_IF_requestR_BIT_159_6_THEN_NEG_requestR__ETC___d2310 =
	     (guard__h60287 == 2'b0) ?
	       11'd0 :
	       (requestR[159] ? _theResult___exp__h60903 : 11'd0) ;
  assign IF_IF_IF_requestR_BIT_159_6_THEN_NEG_requestR__ETC___d2336 =
	     (guard__h61017 == 2'b0 || requestR[159]) ?
	       x__h61032[10:0] :
	       _theResult___exp__h61659 ;
  assign IF_IF_IF_requestR_BIT_159_6_THEN_NEG_requestR__ETC___d2338 =
	     (guard__h61017 == 2'b0) ?
	       x__h61032[10:0] :
	       (requestR[159] ? _theResult___exp__h61659 : x__h61032[10:0]) ;
  assign IF_IF_IF_requestR_BIT_159_6_THEN_NEG_requestR__ETC___d2359 =
	     (guard__h60287 == 2'b0 || requestR[159]) ?
	       sfd___3__h60277[54:3] :
	       _theResult___sfd__h60904 ;
  assign IF_IF_IF_requestR_BIT_159_6_THEN_NEG_requestR__ETC___d2361 =
	     (guard__h60287 == 2'b0) ?
	       sfd___3__h60277[54:3] :
	       (requestR[159] ?
		  _theResult___sfd__h60904 :
		  sfd___3__h60277[54:3]) ;
  assign IF_IF_IF_requestR_BIT_159_6_THEN_NEG_requestR__ETC___d2377 =
	     (guard__h61017 == 2'b0 || requestR[159]) ?
	       sfd___3__h60277[53:2] :
	       _theResult___sfd__h61660 ;
  assign IF_IF_IF_requestR_BIT_159_6_THEN_NEG_requestR__ETC___d2379 =
	     (guard__h61017 == 2'b0) ?
	       sfd___3__h60277[53:2] :
	       (requestR[159] ?
		  _theResult___sfd__h61660 :
		  sfd___3__h60277[53:2]) ;
  assign IF_IF_IF_requestR_BIT_191_27_THEN_NEG_requestR_ETC___d2845 =
	     (guard__h83828 == 2'b0) ?
	       11'd0 :
	       (requestR[191] ? _theResult___exp__h84444 : 11'd0) ;
  assign IF_IF_IF_requestR_BIT_191_27_THEN_NEG_requestR_ETC___d2871 =
	     (guard__h84558 == 2'b0 || requestR[191]) ?
	       x__h84573[10:0] :
	       _theResult___exp__h85200 ;
  assign IF_IF_IF_requestR_BIT_191_27_THEN_NEG_requestR_ETC___d2873 =
	     (guard__h84558 == 2'b0) ?
	       x__h84573[10:0] :
	       (requestR[191] ? _theResult___exp__h85200 : x__h84573[10:0]) ;
  assign IF_IF_IF_requestR_BIT_191_27_THEN_NEG_requestR_ETC___d2894 =
	     (guard__h83828 == 2'b0 || requestR[191]) ?
	       sfd___3__h11835[63:12] :
	       _theResult___sfd__h84445 ;
  assign IF_IF_IF_requestR_BIT_191_27_THEN_NEG_requestR_ETC___d2896 =
	     (guard__h83828 == 2'b0) ?
	       sfd___3__h11835[63:12] :
	       (requestR[191] ?
		  _theResult___sfd__h84445 :
		  sfd___3__h11835[63:12]) ;
  assign IF_IF_IF_requestR_BIT_191_27_THEN_NEG_requestR_ETC___d2912 =
	     (guard__h84558 == 2'b0 || requestR[191]) ?
	       sfd___3__h11835[62:11] :
	       _theResult___sfd__h85201 ;
  assign IF_IF_IF_requestR_BIT_191_27_THEN_NEG_requestR_ETC___d2914 =
	     (guard__h84558 == 2'b0) ?
	       sfd___3__h11835[62:11] :
	       (requestR[191] ?
		  _theResult___sfd__h85201 :
		  sfd___3__h11835[62:11]) ;
  assign IF_IF_IF_requestR_BIT_191_27_THEN_NEG_requestR_ETC___d476 =
	     (guard__h11845 == 2'b0) ?
	       8'd0 :
	       (requestR[191] ? _theResult___exp__h12261 : 8'd0) ;
  assign IF_IF_IF_requestR_BIT_191_27_THEN_NEG_requestR_ETC___d502 =
	     (guard__h12375 == 2'b0 || requestR[191]) ?
	       x__h12390[7:0] :
	       _theResult___exp__h12814 ;
  assign IF_IF_IF_requestR_BIT_191_27_THEN_NEG_requestR_ETC___d504 =
	     (guard__h12375 == 2'b0) ?
	       x__h12390[7:0] :
	       (requestR[191] ? _theResult___exp__h12814 : x__h12390[7:0]) ;
  assign IF_IF_IF_requestR_BIT_191_27_THEN_NEG_requestR_ETC___d525 =
	     (guard__h11845 == 2'b0 || requestR[191]) ?
	       sfd___3__h11835[63:41] :
	       _theResult___sfd__h12262 ;
  assign IF_IF_IF_requestR_BIT_191_27_THEN_NEG_requestR_ETC___d527 =
	     (guard__h11845 == 2'b0) ?
	       sfd___3__h11835[63:41] :
	       (requestR[191] ?
		  _theResult___sfd__h12262 :
		  sfd___3__h11835[63:41]) ;
  assign IF_IF_IF_requestR_BIT_191_27_THEN_NEG_requestR_ETC___d543 =
	     (guard__h12375 == 2'b0 || requestR[191]) ?
	       sfd___3__h11835[62:40] :
	       _theResult___sfd__h12815 ;
  assign IF_IF_IF_requestR_BIT_191_27_THEN_NEG_requestR_ETC___d545 =
	     (guard__h12375 == 2'b0) ?
	       sfd___3__h11835[62:40] :
	       (requestR[191] ?
		  _theResult___sfd__h12815 :
		  sfd___3__h11835[62:40]) ;
  assign IF_IF_requestR_BITS_127_TO_96_2_EQ_0xFFFFFFFF__ETC___d2036 =
	     (sV2_exp__h926 == 8'd255 && sV2_sfd__h927[22] ||
	      IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d2005) ?
	       { requestR[191:160] == 32'hFFFFFFFF && requestR[159],
		 IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d19 } :
	       (IF_requestR_BITS_127_TO_96_2_EQ_0xFFFFFFFF_3_T_ETC___d2009 ?
		  requestR_BITS_127_TO_96_2_EQ_0xFFFFFFFF_3_AND__ETC___d28 :
		  IF_NOT_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFF_ETC___d2034) ;
  assign IF_IF_requestR_BITS_127_TO_96_2_EQ_0xFFFFFFFF__ETC___d2040 =
	     (sV2_exp__h926 == 8'd255 && sV2_sfd__h927 != 23'd0 &&
	      !sV2_sfd__h927[22]) ?
	       res__h42577 :
	       IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_ETC___d2039 ;
  assign IF_IF_requestR_BITS_127_TO_96_2_EQ_0xFFFFFFFF__ETC___d2050 =
	     IF_requestR_BITS_127_TO_96_2_EQ_0xFFFFFFFF_3_T_ETC___d2009 ?
	       { requestR[191:160] == 32'hFFFFFFFF && requestR[159],
		 IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d19 } :
	       IF_NOT_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFF_ETC___d2049 ;
  assign IF_IF_requestR_BITS_127_TO_96_2_EQ_0xFFFFFFFF__ETC___d2052 =
	     (sV2_exp__h926 == 8'd255 && sV2_sfd__h927[22]) ?
	       { requestR[191:160] == 32'hFFFFFFFF && requestR[159],
		 IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d19 } :
	       (IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d2005 ?
		  requestR_BITS_127_TO_96_2_EQ_0xFFFFFFFF_3_AND__ETC___d28 :
		  IF_IF_requestR_BITS_127_TO_96_2_EQ_0xFFFFFFFF__ETC___d2050) ;
  assign IF_IF_requestR_BITS_127_TO_96_2_EQ_0xFFFFFFFF__ETC___d2056 =
	     (sV2_exp__h926 == 8'd255 && sV2_sfd__h927 != 23'd0 &&
	      !sV2_sfd__h927[22]) ?
	       res__h42577 :
	       IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_ETC___d2055 ;
  assign IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_ETC___d1748 =
	     (sV1_exp__h823 == 8'd255 && sV1_sfd__h824 == 23'd0) ?
	       IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d1677 :
	       ((sV1_exp__h823 == 8'd0 && sV1_sfd__h824 == 23'd0) ?
		  64'd0 :
		  IF_NEG_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0_ETC___d1746) ;
  assign IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_ETC___d1807 =
	     (sV1_exp__h823 == 8'd0 && sV1_sfd__h824 == 23'd0) ?
	       64'd0 :
	       (NEG_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFF_ETC___d1778[19] ?
		  64'hFFFFFFFFFFFFFFFF :
		  IF_NEG_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0_ETC___d1805) ;
  assign IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_ETC___d1897 =
	     (sV1_exp__h823 == 8'd255 && sV1_sfd__h824 == 23'd0) ?
	       IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d1834 :
	       ((sV1_exp__h823 == 8'd0 && sV1_sfd__h824 == 23'd0) ?
		  32'd0 :
		  IF_NEG_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0_ETC___d1895) ;
  assign IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_ETC___d1951 =
	     (sV1_exp__h823 == 8'd0 && sV1_sfd__h824 == 23'd0) ?
	       32'd0 :
	       (NEG_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFF_ETC___d1922[19] ?
		  32'hFFFFFFFF :
		  IF_NEG_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0_ETC___d1949) ;
  assign IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_ETC___d2037 =
	     (sV1_exp__h823 == 8'd255 && sV1_sfd__h824[22]) ?
	       requestR_BITS_127_TO_96_2_EQ_0xFFFFFFFF_3_AND__ETC___d28 :
	       IF_IF_requestR_BITS_127_TO_96_2_EQ_0xFFFFFFFF__ETC___d2036 ;
  assign IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_ETC___d2039 =
	     (sV1_exp__h823 == 8'd255 && sV1_sfd__h824[22] &&
	      sV2_exp__h926 == 8'd255 &&
	      sV2_sfd__h927[22]) ?
	       64'hFFFFFFFF7FC00000 :
	       { 32'hFFFFFFFF,
		 IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_ETC___d2037 } ;
  assign IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_ETC___d2041 =
	     (sV1_exp__h823 == 8'd255 && sV1_sfd__h824 != 23'd0 &&
	      !sV1_sfd__h824[22]) ?
	       res__h42340 :
	       IF_IF_requestR_BITS_127_TO_96_2_EQ_0xFFFFFFFF__ETC___d2040 ;
  assign IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_ETC___d2053 =
	     (sV1_exp__h823 == 8'd255 && sV1_sfd__h824[22]) ?
	       requestR_BITS_127_TO_96_2_EQ_0xFFFFFFFF_3_AND__ETC___d28 :
	       IF_IF_requestR_BITS_127_TO_96_2_EQ_0xFFFFFFFF__ETC___d2052 ;
  assign IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_ETC___d2055 =
	     (sV1_exp__h823 == 8'd255 && sV1_sfd__h824[22] &&
	      sV2_exp__h926 == 8'd255 &&
	      sV2_sfd__h927[22]) ?
	       64'hFFFFFFFF7FC00000 :
	       { 32'hFFFFFFFF,
		 IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_ETC___d2053 } ;
  assign IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_ETC___d2057 =
	     (sV1_exp__h823 == 8'd255 && sV1_sfd__h824 != 23'd0 &&
	      !sV1_sfd__h824[22]) ?
	       res__h42340 :
	       IF_IF_requestR_BITS_127_TO_96_2_EQ_0xFFFFFFFF__ETC___d2056 ;
  assign IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_ETC___d2127 =
	     (sV1_exp__h823 == 8'd0 && sV1_sfd__h824 == 23'd0) ?
	       res___1__h50982 :
	       ((sV1_exp__h823 == 8'd0) ? res___1__h51001 : res__h51017) ;
  assign IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_ETC___d2128 =
	     (sV1_exp__h823 == 8'd255 && sV1_sfd__h824 == 23'd0) ?
	       res___1__h50972 :
	       IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_ETC___d2127 ;
  assign IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_ETC___d4495 =
	     ((sV1_exp__h823 == 8'd0) ?
		(sV1_sfd__h824[22] ?
		   6'd2 :
		   (sV1_sfd__h824[21] ?
		      6'd3 :
		      (sV1_sfd__h824[20] ?
			 6'd4 :
			 (sV1_sfd__h824[19] ?
			    6'd5 :
			    (sV1_sfd__h824[18] ?
			       6'd6 :
			       (sV1_sfd__h824[17] ?
				  6'd7 :
				  (sV1_sfd__h824[16] ?
				     6'd8 :
				     (sV1_sfd__h824[15] ?
					6'd9 :
					(sV1_sfd__h824[14] ?
					   6'd10 :
					   (sV1_sfd__h824[13] ?
					      6'd11 :
					      (sV1_sfd__h824[12] ?
						 6'd12 :
						 (sV1_sfd__h824[11] ?
						    6'd13 :
						    (sV1_sfd__h824[10] ?
						       6'd14 :
						       (sV1_sfd__h824[9] ?
							  6'd15 :
							  (sV1_sfd__h824[8] ?
							     6'd16 :
							     (sV1_sfd__h824[7] ?
								6'd17 :
								(sV1_sfd__h824[6] ?
								   6'd18 :
								   (sV1_sfd__h824[5] ?
								      6'd19 :
								      (sV1_sfd__h824[4] ?
									 6'd20 :
									 (sV1_sfd__h824[3] ?
									    6'd21 :
									    (sV1_sfd__h824[2] ?
									       6'd22 :
									       (sV1_sfd__h824[1] ?
										  6'd23 :
										  (sV1_sfd__h824[0] ?
										     6'd24 :
										     6'd57))))))))))))))))))))))) :
		6'd1) -
	     6'd1 ;
  assign IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_ETC___d5035 =
	     (sV1_exp__h823 == 8'd255 && sV1_sfd__h824 != 23'd0) ?
	       _theResult___snd_fst_sfd__h150153 :
	       _theResult___fst_sfd__h188280 ;
  assign IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_ETC___d5071 =
	     (sV1_exp__h823 == 8'd255 && sV1_sfd__h824 != 23'd0 ||
	      (sV1_exp__h823 == 8'd255 || sV1_exp__h823 == 8'd0) &&
	      sV1_sfd__h824 == 23'd0) ?
	       requestR[191:160] == 32'hFFFFFFFF && requestR[159] :
	       ((sV1_exp__h823 == 8'd0) ?
		  IF_NOT_3970_MINUS_0_CONCAT_IF_IF_requestR_BITS_ETC___d5051 :
		  IF_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFFF_ETC___d5069) ;
  assign IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_ETC___d5106 =
	     (sV1_exp__h823 == 8'd0) ?
	       _3970_MINUS_0_CONCAT_IF_IF_requestR_BITS_191_TO_ETC___d4424 &&
	       !_3970_MINUS_0_CONCAT_IF_IF_requestR_BITS_191_TO_ETC___d4425 &&
	       _0_CONCAT_IF_IF_requestR_BITS_191_TO_160_4_EQ_0_ETC___d5085[4] :
	       SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFF_ETC___d4567 &&
	       SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFF_ETC___d4568 &&
	       _0_CONCAT_IF_IF_3074_MINUS_SEXT_IF_requestR_BIT_ETC___d5102[4] ;
  assign IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_ETC___d5109 =
	     (sV1_exp__h823 == 8'd255 && sV1_sfd__h824 != 23'd0) ?
	       sV1_exp__h823 == 8'd255 && sV1_sfd__h824 != 23'd0 &&
	       !sV1_sfd__h824[22] :
	       (sV1_exp__h823 != 8'd255 || sV1_sfd__h824 != 23'd0) &&
	       (value_BIT_23___h161776 || sV1_sfd__h824 != 23'd0) &&
	       IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_ETC___d5106 ;
  assign IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_ETC___d5116 =
	     (sV1_exp__h823 == 8'd0) ?
	       _3970_MINUS_0_CONCAT_IF_IF_requestR_BITS_191_TO_ETC___d4424 &&
	       !_3970_MINUS_0_CONCAT_IF_IF_requestR_BITS_191_TO_ETC___d4425 &&
	       _0_CONCAT_IF_IF_requestR_BITS_191_TO_160_4_EQ_0_ETC___d5085[3] :
	       SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFF_ETC___d4567 &&
	       SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFF_ETC___d4568 &&
	       _0_CONCAT_IF_IF_3074_MINUS_SEXT_IF_requestR_BIT_ETC___d5102[3] ;
  assign IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_ETC___d5130 =
	     (sV1_exp__h823 == 8'd0) ?
	       !_3970_MINUS_0_CONCAT_IF_IF_requestR_BITS_191_TO_ETC___d4424 ||
	       !_3970_MINUS_0_CONCAT_IF_IF_requestR_BITS_191_TO_ETC___d4425 &&
	       _0_CONCAT_IF_IF_requestR_BITS_191_TO_160_4_EQ_0_ETC___d5085[2] :
	       !SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFF_ETC___d4567 ||
	       IF_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFFF_ETC___d5128 ;
  assign IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_ETC___d5142 =
	     (sV1_exp__h823 == 8'd0) ?
	       _3970_MINUS_0_CONCAT_IF_IF_requestR_BITS_191_TO_ETC___d4424 &&
	       (_3970_MINUS_0_CONCAT_IF_IF_requestR_BITS_191_TO_ETC___d4425 ||
		_0_CONCAT_IF_IF_requestR_BITS_191_TO_160_4_EQ_0_ETC___d5085[1]) :
	       SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFF_ETC___d4567 &&
	       IF_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFFF_ETC___d5140 ;
  assign IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_ETC___d5154 =
	     (sV1_exp__h823 == 8'd0) ?
	       !_3970_MINUS_0_CONCAT_IF_IF_requestR_BITS_191_TO_ETC___d4424 ||
	       !_3970_MINUS_0_CONCAT_IF_IF_requestR_BITS_191_TO_ETC___d4425 &&
	       _0_CONCAT_IF_IF_requestR_BITS_191_TO_160_4_EQ_0_ETC___d5085[0] :
	       !SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFF_ETC___d4567 ||
	       IF_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFFF_ETC___d5152 ;
  assign IF_IF_requestR_BIT_159_6_THEN_NEG_requestR_BIT_ETC___d1252 =
	     sfd__h23980[31] ?
	       6'd0 :
	       (sfd__h23980[30] ?
		  6'd1 :
		  (sfd__h23980[29] ?
		     6'd2 :
		     (sfd__h23980[28] ?
			6'd3 :
			(sfd__h23980[27] ?
			   6'd4 :
			   (sfd__h23980[26] ?
			      6'd5 :
			      (sfd__h23980[25] ?
				 6'd6 :
				 (sfd__h23980[24] ?
				    6'd7 :
				    (sfd__h23980[23] ?
				       6'd8 :
				       (sfd__h23980[22] ?
					  6'd9 :
					  (sfd__h23980[21] ?
					     6'd10 :
					     (sfd__h23980[20] ?
						6'd11 :
						(sfd__h23980[19] ?
						   6'd12 :
						   (sfd__h23980[18] ?
						      6'd13 :
						      (sfd__h23980[17] ?
							 6'd14 :
							 (sfd__h23980[16] ?
							    6'd15 :
							    (sfd__h23980[15] ?
							       6'd16 :
							       (sfd__h23980[14] ?
								  6'd17 :
								  (sfd__h23980[13] ?
								     6'd18 :
								     (sfd__h23980[12] ?
									6'd19 :
									(sfd__h23980[11] ?
									   6'd20 :
									   (sfd__h23980[10] ?
									      6'd21 :
									      (sfd__h23980[9] ?
										 6'd22 :
										 (sfd__h23980[8] ?
										    6'd23 :
										    (sfd__h23980[7] ?
										       6'd24 :
										       (sfd__h23980[6] ?
											  6'd25 :
											  (sfd__h23980[5] ?
											     6'd26 :
											     (sfd__h23980[4] ?
												6'd27 :
												(sfd__h23980[3] ?
												   6'd28 :
												   (sfd__h23980[2] ?
												      6'd29 :
												      (sfd__h23980[1] ?
													 6'd30 :
													 (sfd__h23980[0] ?
													    6'd31 :
													    6'd32))))))))))))))))))))))))))))))) ;
  assign IF_IF_requestR_BIT_159_6_THEN_NEG_requestR_BIT_ETC___d2230 =
	     sfd__h23980[31] ?
	       6'd0 :
	       (sfd__h23980[30] ?
		  6'd1 :
		  (sfd__h23980[29] ?
		     6'd2 :
		     (sfd__h23980[28] ?
			6'd3 :
			(sfd__h23980[27] ?
			   6'd4 :
			   (sfd__h23980[26] ?
			      6'd5 :
			      (sfd__h23980[25] ?
				 6'd6 :
				 (sfd__h23980[24] ?
				    6'd7 :
				    (sfd__h23980[23] ?
				       6'd8 :
				       (sfd__h23980[22] ?
					  6'd9 :
					  (sfd__h23980[21] ?
					     6'd10 :
					     (sfd__h23980[20] ?
						6'd11 :
						(sfd__h23980[19] ?
						   6'd12 :
						   (sfd__h23980[18] ?
						      6'd13 :
						      (sfd__h23980[17] ?
							 6'd14 :
							 (sfd__h23980[16] ?
							    6'd15 :
							    (sfd__h23980[15] ?
							       6'd16 :
							       (sfd__h23980[14] ?
								  6'd17 :
								  (sfd__h23980[13] ?
								     6'd18 :
								     (sfd__h23980[12] ?
									6'd19 :
									(sfd__h23980[11] ?
									   6'd20 :
									   (sfd__h23980[10] ?
									      6'd21 :
									      (sfd__h23980[9] ?
										 6'd22 :
										 (sfd__h23980[8] ?
										    6'd23 :
										    (sfd__h23980[7] ?
										       6'd24 :
										       (sfd__h23980[6] ?
											  6'd25 :
											  (sfd__h23980[5] ?
											     6'd26 :
											     (sfd__h23980[4] ?
												6'd27 :
												(sfd__h23980[3] ?
												   6'd28 :
												   (sfd__h23980[2] ?
												      6'd29 :
												      (sfd__h23980[1] ?
													 6'd30 :
													 (sfd__h23980[0] ?
													    6'd31 :
													    6'd55))))))))))))))))))))))))))))))) ;
  assign IF_IF_requestR_BIT_191_27_THEN_NEG_requestR_BI_ETC___d384 =
	     sfd__h2230[63] ?
	       7'd0 :
	       (sfd__h2230[62] ?
		  7'd1 :
		  (sfd__h2230[61] ?
		     7'd2 :
		     (sfd__h2230[60] ?
			7'd3 :
			(sfd__h2230[59] ?
			   7'd4 :
			   (sfd__h2230[58] ?
			      7'd5 :
			      (sfd__h2230[57] ?
				 7'd6 :
				 (sfd__h2230[56] ?
				    7'd7 :
				    (sfd__h2230[55] ?
				       7'd8 :
				       (sfd__h2230[54] ?
					  7'd9 :
					  (sfd__h2230[53] ?
					     7'd10 :
					     (sfd__h2230[52] ?
						7'd11 :
						(sfd__h2230[51] ?
						   7'd12 :
						   (sfd__h2230[50] ?
						      7'd13 :
						      (sfd__h2230[49] ?
							 7'd14 :
							 (sfd__h2230[48] ?
							    7'd15 :
							    (sfd__h2230[47] ?
							       7'd16 :
							       (sfd__h2230[46] ?
								  7'd17 :
								  (sfd__h2230[45] ?
								     7'd18 :
								     (sfd__h2230[44] ?
									7'd19 :
									(sfd__h2230[43] ?
									   7'd20 :
									   (sfd__h2230[42] ?
									      7'd21 :
									      (sfd__h2230[41] ?
										 7'd22 :
										 (sfd__h2230[40] ?
										    7'd23 :
										    (sfd__h2230[39] ?
										       7'd24 :
										       (sfd__h2230[38] ?
											  7'd25 :
											  (sfd__h2230[37] ?
											     7'd26 :
											     (sfd__h2230[36] ?
												7'd27 :
												(sfd__h2230[35] ?
												   7'd28 :
												   (sfd__h2230[34] ?
												      7'd29 :
												      (sfd__h2230[33] ?
													 7'd30 :
													 (sfd__h2230[32] ?
													    7'd31 :
													    (sfd__h2230[31] ?
													       7'd32 :
													       (sfd__h2230[30] ?
														  7'd33 :
														  (sfd__h2230[29] ?
														     7'd34 :
														     (sfd__h2230[28] ?
															7'd35 :
															(sfd__h2230[27] ?
															   7'd36 :
															   (sfd__h2230[26] ?
															      7'd37 :
															      (sfd__h2230[25] ?
																 7'd38 :
																 (sfd__h2230[24] ?
																    7'd39 :
																    (sfd__h2230[23] ?
																       7'd40 :
																       (sfd__h2230[22] ?
																	  7'd41 :
																	  (sfd__h2230[21] ?
																	     7'd42 :
																	     (sfd__h2230[20] ?
																		7'd43 :
																		(sfd__h2230[19] ?
																		   7'd44 :
																		   (sfd__h2230[18] ?
																		      7'd45 :
																		      (sfd__h2230[17] ?
																			 7'd46 :
																			 (sfd__h2230[16] ?
																			    7'd47 :
																			    (sfd__h2230[15] ?
																			       7'd48 :
																			       (sfd__h2230[14] ?
																				  7'd49 :
																				  (sfd__h2230[13] ?
																				     7'd50 :
																				     (sfd__h2230[12] ?
																					7'd51 :
																					(sfd__h2230[11] ?
																					   7'd52 :
																					   (sfd__h2230[10] ?
																					      7'd53 :
																					      (sfd__h2230[9] ?
																						 7'd54 :
																						 (sfd__h2230[8] ?
																						    7'd55 :
																						    (sfd__h2230[7] ?
																						       7'd56 :
																						       (sfd__h2230[6] ?
																							  7'd57 :
																							  (sfd__h2230[5] ?
																							     7'd58 :
																							     (sfd__h2230[4] ?
																								7'd59 :
																								(sfd__h2230[3] ?
																								   7'd60 :
																								   (sfd__h2230[2] ?
																								      7'd61 :
																								      (sfd__h2230[1] ?
																									 7'd62 :
																									 (sfd__h2230[0] ?
																									    7'd63 :
																									    7'd64))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) ;
  assign IF_NEG_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0_ETC___d1744 =
	     NEG_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFF_ETC___d1717 ?
	       (IF_requestR_BITS_194_TO_192_0_EQ_0x0_1_OR_NOT__ETC___d1738 ?
		  ((x__h37699[88:25] == 64'h7FFFFFFFFFFFFFFF) ?
		     x__h37699[88:25] :
		     x__h37699[88:25] + 64'd1) :
		  x__h37699[88:25]) :
	       64'd0 ;
  assign IF_NEG_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0_ETC___d1746 =
	     (NEG_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFF_ETC___d1682 ==
	      20'd1048513) ?
	       ((_theResult_____2__h36734[64:63] == 2'b11) ?
		  _theResult_____2__h36734[63:0] :
		  IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d1677) :
	       (NEG_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFF_ETC___d1715[19] ?
		  IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d1677 :
		  IF_NEG_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0_ETC___d1744) ;
  assign IF_NEG_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0_ETC___d1769 =
	     (NEG_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFF_ETC___d1682 ==
	      20'd1048513) ?
	       _theResult_____2__h36734[64:63] == 2'b11 &&
	       guard__h36732 != 2'd0 :
	       !NEG_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFF_ETC___d1715[19] &&
	       (!NEG_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFF_ETC___d1717 ||
		guard__h37510 != 2'd0) ;
  assign IF_NEG_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0_ETC___d1805 =
	     NEG_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFF_ETC___d1780 ?
	       (IF_requestR_BITS_194_TO_192_0_EQ_0x0_1_OR_NOT__ETC___d1799 ?
		  ((x__h39015[88:25] == 64'hFFFFFFFFFFFFFFFF) ?
		     x__h39015[88:25] :
		     x__h39015[88:25] + 64'd1) :
		  x__h39015[88:25]) :
	       64'd0 ;
  assign IF_NEG_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0_ETC___d1893 =
	     NEG_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFF_ETC___d1866 ?
	       (IF_requestR_BITS_194_TO_192_0_EQ_0x0_1_OR_NOT__ETC___d1887 ?
		  ((x__h40258[56:25] == 32'h7FFFFFFF) ?
		     x__h40258[56:25] :
		     x__h40258[56:25] + 32'd1) :
		  x__h40258[56:25]) :
	       32'd0 ;
  assign IF_NEG_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0_ETC___d1895 =
	     (NEG_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFF_ETC___d1682 ==
	      20'd1048545) ?
	       ((_theResult_____2__h39517[32:31] == 2'b11) ?
		  _theResult_____2__h39517[31:0] :
		  IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d1834) :
	       (NEG_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFF_ETC___d1864[19] ?
		  IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d1834 :
		  IF_NEG_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0_ETC___d1893) ;
  assign IF_NEG_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0_ETC___d1913 =
	     (NEG_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFF_ETC___d1682 ==
	      20'd1048545) ?
	       _theResult_____2__h39517[32:31] == 2'b11 &&
	       guard__h39515 != 2'd0 :
	       !NEG_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFF_ETC___d1864[19] &&
	       (!NEG_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFF_ETC___d1866 ||
		guard__h40069 != 2'd0) ;
  assign IF_NEG_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0_ETC___d1949 =
	     NEG_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFF_ETC___d1924 ?
	       (IF_requestR_BITS_194_TO_192_0_EQ_0x0_1_OR_NOT__ETC___d1943 ?
		  ((x__h41336[56:25] == 32'hFFFFFFFF) ?
		     x__h41336[56:25] :
		     x__h41336[56:25] + 32'd1) :
		  x__h41336[56:25]) :
	       32'd0 ;
  assign IF_NEG_SEXT_requestR_BITS_190_TO_180_599_MINUS_ETC___d2675 =
	     NEG_SEXT_requestR_BITS_190_TO_180_599_MINUS_10_ETC___d2648 ?
	       (IF_requestR_BITS_194_TO_192_0_EQ_0x0_1_OR_NOT__ETC___d2669 ?
		  ((x__h72798[85:54] == 32'h7FFFFFFF) ?
		     x__h72798[85:54] :
		     x__h72798[85:54] + 32'd1) :
		  x__h72798[85:54]) :
	       32'd0 ;
  assign IF_NEG_SEXT_requestR_BITS_190_TO_180_599_MINUS_ETC___d2677 =
	     (NEG_SEXT_requestR_BITS_190_TO_180_599_MINUS_10_ETC___d2613 ==
	      24'd16777185) ?
	       ((_theResult_____2__h72057[32:31] == 2'b11) ?
		  _theResult_____2__h72057[31:0] :
		  IF_requestR_BIT_191_27_THEN_2147483648_ELSE_21_ETC___d2608) :
	       (NEG_SEXT_requestR_BITS_190_TO_180_599_MINUS_10_ETC___d2646[23] ?
		  IF_requestR_BIT_191_27_THEN_2147483648_ELSE_21_ETC___d2608 :
		  IF_NEG_SEXT_requestR_BITS_190_TO_180_599_MINUS_ETC___d2675) ;
  assign IF_NEG_SEXT_requestR_BITS_190_TO_180_599_MINUS_ETC___d2701 =
	     (NEG_SEXT_requestR_BITS_190_TO_180_599_MINUS_10_ETC___d2613 ==
	      24'd16777185) ?
	       _theResult_____2__h72057[32:31] == 2'b11 &&
	       guard__h72055 != 2'd0 :
	       !NEG_SEXT_requestR_BITS_190_TO_180_599_MINUS_10_ETC___d2646[23] &&
	       (!NEG_SEXT_requestR_BITS_190_TO_180_599_MINUS_10_ETC___d2648 ||
		guard__h72609 != 2'd0) ;
  assign IF_NEG_SEXT_requestR_BITS_190_TO_180_599_MINUS_ETC___d2737 =
	     NEG_SEXT_requestR_BITS_190_TO_180_599_MINUS_10_ETC___d2712 ?
	       (IF_requestR_BITS_194_TO_192_0_EQ_0x0_1_OR_NOT__ETC___d2731 ?
		  ((x__h73876[85:54] == 32'hFFFFFFFF) ?
		     x__h73876[85:54] :
		     x__h73876[85:54] + 32'd1) :
		  x__h73876[85:54]) :
	       32'd0 ;
  assign IF_NEG_SEXT_requestR_BITS_190_TO_180_599_MINUS_ETC___d3164 =
	     NEG_SEXT_requestR_BITS_190_TO_180_599_MINUS_10_ETC___d3137 ?
	       (IF_requestR_BITS_194_TO_192_0_EQ_0x0_1_OR_NOT__ETC___d3158 ?
		  ((x__h97876[117:54] == 64'h7FFFFFFFFFFFFFFF) ?
		     x__h97876[117:54] :
		     x__h97876[117:54] + 64'd1) :
		  x__h97876[117:54]) :
	       64'd0 ;
  assign IF_NEG_SEXT_requestR_BITS_190_TO_180_599_MINUS_ETC___d3166 =
	     (NEG_SEXT_requestR_BITS_190_TO_180_599_MINUS_10_ETC___d2613 ==
	      24'd16777153) ?
	       ((_theResult_____2__h96911[64:63] == 2'b11) ?
		  _theResult_____2__h96911[63:0] :
		  IF_requestR_BIT_191_27_THEN_922337203685477580_ETC___d3105) :
	       (NEG_SEXT_requestR_BITS_190_TO_180_599_MINUS_10_ETC___d3135[23] ?
		  IF_requestR_BIT_191_27_THEN_922337203685477580_ETC___d3105 :
		  IF_NEG_SEXT_requestR_BITS_190_TO_180_599_MINUS_ETC___d3164) ;
  assign IF_NEG_SEXT_requestR_BITS_190_TO_180_599_MINUS_ETC___d3183 =
	     (NEG_SEXT_requestR_BITS_190_TO_180_599_MINUS_10_ETC___d2613 ==
	      24'd16777153) ?
	       _theResult_____2__h96911[64:63] == 2'b11 &&
	       guard__h96909 != 2'd0 :
	       !NEG_SEXT_requestR_BITS_190_TO_180_599_MINUS_10_ETC___d3135[23] &&
	       (!NEG_SEXT_requestR_BITS_190_TO_180_599_MINUS_10_ETC___d3137 ||
		guard__h97687 != 2'd0) ;
  assign IF_NEG_SEXT_requestR_BITS_190_TO_180_599_MINUS_ETC___d3219 =
	     NEG_SEXT_requestR_BITS_190_TO_180_599_MINUS_10_ETC___d3194 ?
	       (IF_requestR_BITS_194_TO_192_0_EQ_0x0_1_OR_NOT__ETC___d3213 ?
		  ((x__h99175[117:54] == 64'hFFFFFFFFFFFFFFFF) ?
		     x__h99175[117:54] :
		     x__h99175[117:54] + 64'd1) :
		  x__h99175[117:54]) :
	       64'd0 ;
  assign IF_NOT_32_MINUS_0_CONCAT_IF_IF_requestR_BIT_15_ETC___d2290 =
	     (!_32_MINUS_0_CONCAT_IF_IF_requestR_BIT_159_6_THE_ETC___d2234 ||
	      _32_MINUS_0_CONCAT_IF_IF_requestR_BIT_159_6_THE_ETC___d2236) ?
	       requestR[159] :
	       IF_32_MINUS_0_CONCAT_IF_IF_requestR_BIT_159_6__ETC___d2289 ;
  assign IF_NOT_3970_MINUS_0_CONCAT_IF_IF_requestR_BITS_ETC___d5051 =
	     (!_3970_MINUS_0_CONCAT_IF_IF_requestR_BITS_191_TO_ETC___d4424 ||
	      _3970_MINUS_0_CONCAT_IF_IF_requestR_BITS_191_TO_ETC___d4425 ||
	      _theResult___fst_exp__h169079 == 11'd2047) ?
	       requestR[191:160] == 32'hFFFFFFFF && requestR[159] :
	       ((requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
		 requestR[194:192] != 3'h3 &&
		 requestR[194:192] != 3'h4) ?
		  CASE_guard61118_0b0_requestR_BITS_191_TO_160_E_ETC__q162 :
		  CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q163) ;
  assign IF_NOT_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFF_ETC___d2034 =
	     NOT_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFF_ETC___d2033 ?
	       { requestR[191:160] == 32'hFFFFFFFF && requestR[159],
		 IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d19 } :
	       requestR_BITS_127_TO_96_2_EQ_0xFFFFFFFF_3_AND__ETC___d28 ;
  assign IF_NOT_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFF_ETC___d2049 =
	     NOT_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFF_ETC___d2033 ?
	       requestR_BITS_127_TO_96_2_EQ_0xFFFFFFFF_3_AND__ETC___d28 :
	       { requestR[191:160] == 32'hFFFFFFFF && requestR[159],
		 IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d19 } ;
  assign IF_NOT_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFF_ETC___d2029 =
	     (requestR[191:160] != 32'hFFFFFFFF || !requestR[159]) ?
	       IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d2018 ||
	       IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d2019 &&
	       IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d2020 :
	       !IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d2023 ||
	       IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d2019 &&
	       !IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d2025 ;
  assign IF_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFFF_ETC___d4889 =
	     ((SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFF_ETC__q150[10:0] ==
	       11'd0) ?
		12'd3074 :
		{ SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFF_ETC__q153[10],
		  SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFF_ETC__q153 }) -
	     12'd3074 ;
  assign IF_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFFF_ETC___d5069 =
	     SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFF_ETC___d4567 ?
	       (SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFF_ETC___d4568 ?
		  IF_IF_IF_3074_MINUS_SEXT_IF_requestR_BITS_191__ETC___d5059 :
		  IF_IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFF_ETC___d5067) :
	       requestR[191:160] == 32'hFFFFFFFF && requestR[159] ;
  assign IF_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFFF_ETC___d5128 =
	     SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFF_ETC___d4568 ?
	       _0_CONCAT_IF_IF_3074_MINUS_SEXT_IF_requestR_BIT_ETC___d5102[2] :
	       _theResult___fst_exp__h188264 == 11'd2047 &&
	       _theResult___fst_sfd__h188265 == 52'd0 ;
  assign IF_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFFF_ETC___d5140 =
	     SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFF_ETC___d4568 ?
	       _0_CONCAT_IF_IF_3074_MINUS_SEXT_IF_requestR_BIT_ETC___d5102[1] :
	       _theResult___fst_exp__h187483 == 11'd0 &&
	       guard__h179493 != 2'b0 ;
  assign IF_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFFF_ETC___d5152 =
	     SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFF_ETC___d4568 ?
	       _0_CONCAT_IF_IF_3074_MINUS_SEXT_IF_requestR_BIT_ETC___d5102[0] :
	       _theResult___fst_exp__h187483 != 11'd2047 &&
	       guard__h179493 != 2'b0 ;
  assign IF_SEXT_requestR_BITS_190_TO_180_599_MINUS_102_ETC___d4055 =
	     ((SEXT_requestR_BITS_190_TO_180_599_MINUS_1023_6_ETC__q118[7:0] ==
	       8'd0) ?
		9'd386 :
		{ SEXT_requestR_BITS_190_TO_180_599_MINUS_1023_6_ETC__q121[7],
		  SEXT_requestR_BITS_190_TO_180_599_MINUS_1023_6_ETC__q121 }) -
	     9'd386 ;
  assign IF_SEXT_requestR_BITS_190_TO_180_599_MINUS_102_ETC___d4259 =
	     SEXT_requestR_BITS_190_TO_180_599_MINUS_1023_6_ETC___d3736 ?
	       ((_theResult___fst_exp__h137317 == 8'd255) ?
		  requestR[191] :
		  ((requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
		    requestR[194:192] != 3'h3 &&
		    requestR[194:192] != 3'h4) ?
		     CASE_guard29091_0b0_requestR_BIT_191_0b1_reque_ETC__q144 :
		     CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q145)) :
	       ((_theResult___fst_exp__h146032 == 8'd255) ?
		  requestR[191] :
		  ((requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
		    requestR[194:192] != 3'h3 &&
		    requestR[194:192] != 3'h4) ?
		     CASE_guard37955_0b0_requestR_BIT_191_0b1_reque_ETC__q146 :
		     CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q147)) ;
  assign IF_SEXT_requestR_BITS_190_TO_180_599_MINUS_102_ETC___d4337 =
	     SEXT_requestR_BITS_190_TO_180_599_MINUS_1023_6_ETC___d3736 ?
	       _0_CONCAT_IF_IF_3970_MINUS_SEXT_requestR_BITS_1_ETC___d4308[2] :
	       _theResult___fst_exp__h146610 == 8'd255 &&
	       _theResult___fst_sfd__h146611 == 23'd0 ;
  assign IF_SEXT_requestR_BITS_190_TO_180_599_MINUS_102_ETC___d4350 =
	     SEXT_requestR_BITS_190_TO_180_599_MINUS_1023_6_ETC___d3736 ?
	       _0_CONCAT_IF_IF_3970_MINUS_SEXT_requestR_BITS_1_ETC___d4308[1] :
	       _theResult___fst_exp__h146032 == 8'd0 &&
	       guard__h137955 != 2'b0 ;
  assign IF_SEXT_requestR_BITS_190_TO_180_599_MINUS_102_ETC___d4363 =
	     SEXT_requestR_BITS_190_TO_180_599_MINUS_1023_6_ETC___d3736 ?
	       _0_CONCAT_IF_IF_3970_MINUS_SEXT_requestR_BITS_1_ETC___d4308[0] :
	       _theResult___fst_exp__h146032 != 8'd255 &&
	       guard__h137955 != 2'b0 ;
  assign IF_requestR_BITS_126_TO_116_166_EQ_2047_167_AN_ETC___d5214 =
	     (requestR[126:116] == 11'd2047 && requestR[115] ||
	      requestR_BITS_190_TO_180_599_EQ_0_609_AND_requ_ETC___d5183) ?
	       requestR[191:128] :
	       (requestR_BITS_126_TO_116_166_EQ_0_180_AND_requ_ETC___d5187 ?
		  requestR[127:64] :
		  res__h193345) ;
  assign IF_requestR_BITS_127_TO_96_2_EQ_0xFFFFFFFF_3_T_ETC___d2009 =
	     sV2_exp__h926 == 8'd0 && sV2_sfd__h927 == 23'd0 &&
	     requestR[127:96] == 32'hFFFFFFFF &&
	     requestR[95] &&
	     sV1_exp__h823 == 8'd0 &&
	     sV1_sfd__h824 == 23'd0 &&
	     (requestR[191:160] != 32'hFFFFFFFF || !requestR[159]) ;
  assign IF_requestR_BITS_159_TO_128_121_EQ_0_122_OR_NO_ETC___d1373 =
	     (requestR[159:128] == 32'd0 ||
	      !sfd__h23980[31] && !sfd__h23980[30] && !sfd__h23980[29] &&
	      !sfd__h23980[28] &&
	      !sfd__h23980[27] &&
	      !sfd__h23980[26] &&
	      !sfd__h23980[25] &&
	      !sfd__h23980[24] &&
	      !sfd__h23980[23] &&
	      !sfd__h23980[22] &&
	      !sfd__h23980[21] &&
	      !sfd__h23980[20] &&
	      !sfd__h23980[19] &&
	      !sfd__h23980[18] &&
	      !sfd__h23980[17] &&
	      !sfd__h23980[16] &&
	      !sfd__h23980[15] &&
	      !sfd__h23980[14] &&
	      !sfd__h23980[13] &&
	      !sfd__h23980[12] &&
	      !sfd__h23980[11] &&
	      !sfd__h23980[10] &&
	      !sfd__h23980[9] &&
	      !sfd__h23980[8] &&
	      !sfd__h23980[7] &&
	      !sfd__h23980[6] &&
	      !sfd__h23980[5] &&
	      !sfd__h23980[4] &&
	      !sfd__h23980[3] &&
	      !sfd__h23980[2] &&
	      !sfd__h23980[1] &&
	      !sfd__h23980[0]) ?
	       8'd0 :
	       _theResult___snd_fst_exp__h29969 ;
  assign IF_requestR_BITS_159_TO_128_121_EQ_0_122_OR_NO_ETC___d1596 =
	     (requestR[159:128] == 32'd0 ||
	      !requestR[159] &&
	      NOT_requestR_BIT_158_12_13_AND_NOT_requestR_BI_ETC___d803) ?
	       8'd0 :
	       _theResult___snd_fst_exp__h36138 ;
  assign IF_requestR_BITS_159_TO_128_121_EQ_0_122_OR_NO_ETC___d2387 =
	     (requestR[159:128] == 32'd0 ||
	      !_32_MINUS_0_CONCAT_IF_IF_requestR_BIT_159_6_THE_ETC___d2234 ||
	      _32_MINUS_0_CONCAT_IF_IF_requestR_BIT_159_6_THE_ETC___d2236) ?
	       52'd0 :
	       _theResult___snd_fst_sfd__h61763 ;
  assign IF_requestR_BITS_159_TO_128_121_EQ_0_122_OR_NO_ETC___d2570 =
	     (requestR[159:128] == 32'd0 ||
	      !_32_MINUS_0_CONCAT_IF_requestR_BIT_159_6_THEN_0_ETC___d2449 ||
	      _32_MINUS_0_CONCAT_IF_requestR_BIT_159_6_THEN_0_ETC___d2450) ?
	       52'd0 :
	       _theResult___snd_fst_sfd__h71457 ;
  assign IF_requestR_BITS_190_TO_180_599_EQ_0_609_AND_r_ETC___d2739 =
	     (requestR[190:180] == 11'd0 && requestR[179:128] == 52'd0) ?
	       32'd0 :
	       (NEG_SEXT_requestR_BITS_190_TO_180_599_MINUS_10_ETC___d2710[23] ?
		  32'hFFFFFFFF :
		  IF_NEG_SEXT_requestR_BITS_190_TO_180_599_MINUS_ETC___d2737) ;
  assign IF_requestR_BITS_190_TO_180_599_EQ_0_609_AND_r_ETC___d3221 =
	     (requestR[190:180] == 11'd0 && requestR[179:128] == 52'd0) ?
	       64'd0 :
	       (NEG_SEXT_requestR_BITS_190_TO_180_599_MINUS_10_ETC___d3192[23] ?
		  64'hFFFFFFFFFFFFFFFF :
		  IF_NEG_SEXT_requestR_BITS_190_TO_180_599_MINUS_ETC___d3219) ;
  assign IF_requestR_BITS_190_TO_180_599_EQ_0_609_AND_r_ETC___d5228 =
	     requestR_BITS_190_TO_180_599_EQ_0_609_AND_requ_ETC___d5183 ?
	       requestR[127:64] :
	       (requestR_BITS_126_TO_116_166_EQ_0_180_AND_requ_ETC___d5187 ?
		  requestR[191:128] :
		  res__h197893) ;
  assign IF_requestR_BITS_190_TO_180_599_EQ_0_609_AND_r_ETC___d5299 =
	     (requestR[190:180] == 11'd0 && requestR[179:128] == 52'd0) ?
	       res___1__h206085 :
	       ((requestR[190:180] == 11'd0) ?
		  res___1__h206104 :
		  res__h206120) ;
  assign IF_requestR_BITS_190_TO_180_599_EQ_0_609_THEN__ETC___d3659 =
	     ((requestR[190:180] == 11'd0) ?
		(requestR[179] ?
		   6'd2 :
		   (requestR[178] ?
		      6'd3 :
		      (requestR[177] ?
			 6'd4 :
			 (requestR[176] ?
			    6'd5 :
			    (requestR[175] ?
			       6'd6 :
			       (requestR[174] ?
				  6'd7 :
				  (requestR[173] ?
				     6'd8 :
				     (requestR[172] ?
					6'd9 :
					(requestR[171] ?
					   6'd10 :
					   (requestR[170] ?
					      6'd11 :
					      (requestR[169] ?
						 6'd12 :
						 (requestR[168] ?
						    6'd13 :
						    (requestR[167] ?
						       6'd14 :
						       (requestR[166] ?
							  6'd15 :
							  (requestR[165] ?
							     6'd16 :
							     (requestR[164] ?
								6'd17 :
								(requestR[163] ?
								   6'd18 :
								   (requestR[162] ?
								      6'd19 :
								      (requestR[161] ?
									 6'd20 :
									 (requestR[160] ?
									    6'd21 :
									    (requestR[159] ?
									       6'd22 :
									       (requestR[158] ?
										  6'd23 :
										  (requestR[157] ?
										     6'd24 :
										     (requestR[156] ?
											6'd25 :
											(requestR[155] ?
											   6'd26 :
											   (requestR[154] ?
											      6'd27 :
											      (requestR[153] ?
												 6'd28 :
												 (requestR[152] ?
												    6'd29 :
												    (requestR[151] ?
												       6'd30 :
												       (requestR[150] ?
													  6'd31 :
													  (requestR[149] ?
													     6'd32 :
													     (requestR[148] ?
														6'd33 :
														(requestR[147] ?
														   6'd34 :
														   (requestR[146] ?
														      6'd35 :
														      (requestR[145] ?
															 6'd36 :
															 (requestR[144] ?
															    6'd37 :
															    (requestR[143] ?
															       6'd38 :
															       (requestR[142] ?
																  6'd39 :
																  (requestR[141] ?
																     6'd40 :
																     (requestR[140] ?
																	6'd41 :
																	(requestR[139] ?
																	   6'd42 :
																	   (requestR[138] ?
																	      6'd43 :
																	      (requestR[137] ?
																		 6'd44 :
																		 (requestR[136] ?
																		    6'd45 :
																		    (requestR[135] ?
																		       6'd46 :
																		       (requestR[134] ?
																			  6'd47 :
																			  (requestR[133] ?
																			     6'd48 :
																			     (requestR[132] ?
																				6'd49 :
																				(requestR[131] ?
																				   6'd50 :
																				   (requestR[130] ?
																				      6'd51 :
																				      (requestR[129] ?
																					 6'd52 :
																					 (requestR[128] ?
																					    6'd53 :
																					    6'd57)))))))))))))))))))))))))))))))))))))))))))))))))))) :
		6'd1) -
	     6'd1 ;
  assign IF_requestR_BITS_190_TO_180_599_EQ_0_609_THEN__ETC___d4261 =
	     (requestR[190:180] == 11'd0) ?
	       (_3074_MINUS_0_CONCAT_IF_requestR_BIT_179_71_THE_ETC___d3304 ?
		  IF_3074_MINUS_0_CONCAT_IF_requestR_BIT_179_71__ETC___d4241 :
		  requestR[191]) :
	       (SEXT_requestR_BITS_190_TO_180_599_MINUS_1023_6_ETC___d3735 ?
		  IF_SEXT_requestR_BITS_190_TO_180_599_MINUS_102_ETC___d4259 :
		  requestR[191]) ;
  assign IF_requestR_BITS_190_TO_180_599_EQ_0_609_THEN__ETC___d4312 =
	     (requestR[190:180] == 11'd0) ?
	       _3074_MINUS_0_CONCAT_IF_requestR_BIT_179_71_THE_ETC___d4294 :
	       SEXT_requestR_BITS_190_TO_180_599_MINUS_1023_6_ETC___d3735 &&
	       SEXT_requestR_BITS_190_TO_180_599_MINUS_1023_6_ETC___d3736 &&
	       _0_CONCAT_IF_IF_3970_MINUS_SEXT_requestR_BITS_1_ETC___d4308[4] ;
  assign IF_requestR_BITS_190_TO_180_599_EQ_0_609_THEN__ETC___d4323 =
	     (requestR[190:180] == 11'd0) ?
	       _3074_MINUS_0_CONCAT_IF_requestR_BIT_179_71_THE_ETC___d4319 :
	       SEXT_requestR_BITS_190_TO_180_599_MINUS_1023_6_ETC___d3735 &&
	       SEXT_requestR_BITS_190_TO_180_599_MINUS_1023_6_ETC___d3736 &&
	       _0_CONCAT_IF_IF_3970_MINUS_SEXT_requestR_BITS_1_ETC___d4308[3] ;
  assign IF_requestR_BITS_190_TO_180_599_EQ_0_609_THEN__ETC___d4339 =
	     (requestR[190:180] == 11'd0) ?
	       NOT_3074_MINUS_0_CONCAT_IF_requestR_BIT_179_71_ETC___d4331 :
	       !SEXT_requestR_BITS_190_TO_180_599_MINUS_1023_6_ETC___d3735 ||
	       IF_SEXT_requestR_BITS_190_TO_180_599_MINUS_102_ETC___d4337 ;
  assign IF_requestR_BITS_190_TO_180_599_EQ_0_609_THEN__ETC___d4352 =
	     (requestR[190:180] == 11'd0) ?
	       _3074_MINUS_0_CONCAT_IF_requestR_BIT_179_71_THE_ETC___d4346 :
	       SEXT_requestR_BITS_190_TO_180_599_MINUS_1023_6_ETC___d3735 &&
	       IF_SEXT_requestR_BITS_190_TO_180_599_MINUS_102_ETC___d4350 ;
  assign IF_requestR_BITS_190_TO_180_599_EQ_0_609_THEN__ETC___d4365 =
	     (requestR[190:180] == 11'd0) ?
	       NOT_3074_MINUS_0_CONCAT_IF_requestR_BIT_179_71_ETC___d4359 :
	       !SEXT_requestR_BITS_190_TO_180_599_MINUS_1023_6_ETC___d3735 ||
	       IF_SEXT_requestR_BITS_190_TO_180_599_MINUS_102_ETC___d4363 ;
  assign IF_requestR_BITS_190_TO_180_599_EQ_2047_600_AN_ETC___d2679 =
	     (requestR[190:180] == 11'd2047 && requestR[179:128] == 52'd0) ?
	       IF_requestR_BIT_191_27_THEN_2147483648_ELSE_21_ETC___d2608 :
	       ((requestR[190:180] == 11'd0 && requestR[179:128] == 52'd0) ?
		  32'd0 :
		  IF_NEG_SEXT_requestR_BITS_190_TO_180_599_MINUS_ETC___d2677) ;
  assign IF_requestR_BITS_190_TO_180_599_EQ_2047_600_AN_ETC___d3168 =
	     (requestR[190:180] == 11'd2047 && requestR[179:128] == 52'd0) ?
	       IF_requestR_BIT_191_27_THEN_922337203685477580_ETC___d3105 :
	       ((requestR[190:180] == 11'd0 && requestR[179:128] == 52'd0) ?
		  64'd0 :
		  IF_NEG_SEXT_requestR_BITS_190_TO_180_599_MINUS_ETC___d3166) ;
  assign IF_requestR_BITS_190_TO_180_599_EQ_2047_600_AN_ETC___d4221 =
	     (requestR[190:180] == 11'd2047 && requestR[179:128] != 52'd0) ?
	       _theResult___snd_fst_sfd__h103681 :
	       _theResult___fst_sfd__h146626 ;
  assign IF_requestR_BITS_191_TO_128_24_EQ_0_25_OR_NOT__ETC___d2883 =
	     (requestR[191:128] == 64'd0 ||
	      !sfd__h2230[63] && !sfd__h2230[62] && !sfd__h2230[61] &&
	      !sfd__h2230[60] &&
	      !sfd__h2230[59] &&
	      !sfd__h2230[58] &&
	      !sfd__h2230[57] &&
	      !sfd__h2230[56] &&
	      !sfd__h2230[55] &&
	      !sfd__h2230[54] &&
	      !sfd__h2230[53] &&
	      !sfd__h2230[52] &&
	      !sfd__h2230[51] &&
	      !sfd__h2230[50] &&
	      !sfd__h2230[49] &&
	      !sfd__h2230[48] &&
	      !sfd__h2230[47] &&
	      !sfd__h2230[46] &&
	      !sfd__h2230[45] &&
	      !sfd__h2230[44] &&
	      !sfd__h2230[43] &&
	      !sfd__h2230[42] &&
	      !sfd__h2230[41] &&
	      !sfd__h2230[40] &&
	      !sfd__h2230[39] &&
	      !sfd__h2230[38] &&
	      !sfd__h2230[37] &&
	      !sfd__h2230[36] &&
	      !sfd__h2230[35] &&
	      !sfd__h2230[34] &&
	      !sfd__h2230[33] &&
	      !sfd__h2230[32] &&
	      !sfd__h2230[31] &&
	      !sfd__h2230[30] &&
	      !sfd__h2230[29] &&
	      !sfd__h2230[28] &&
	      !sfd__h2230[27] &&
	      !sfd__h2230[26] &&
	      !sfd__h2230[25] &&
	      !sfd__h2230[24] &&
	      !sfd__h2230[23] &&
	      !sfd__h2230[22] &&
	      !sfd__h2230[21] &&
	      !sfd__h2230[20] &&
	      !sfd__h2230[19] &&
	      !sfd__h2230[18] &&
	      !sfd__h2230[17] &&
	      !sfd__h2230[16] &&
	      !sfd__h2230[15] &&
	      !sfd__h2230[14] &&
	      !sfd__h2230[13] &&
	      !sfd__h2230[12] &&
	      !sfd__h2230[11] &&
	      !sfd__h2230[10] &&
	      !sfd__h2230[9] &&
	      !sfd__h2230[8] &&
	      !sfd__h2230[7] &&
	      !sfd__h2230[6] &&
	      !sfd__h2230[5] &&
	      !sfd__h2230[4] &&
	      !sfd__h2230[3] &&
	      !sfd__h2230[2] &&
	      !sfd__h2230[1] &&
	      !sfd__h2230[0]) ?
	       11'd0 :
	       _theResult___snd_fst_exp__h85309 ;
  assign IF_requestR_BITS_191_TO_128_24_EQ_0_25_OR_NOT__ETC___d514 =
	     (requestR[191:128] == 64'd0 ||
	      !sfd__h2230[63] && !sfd__h2230[62] && !sfd__h2230[61] &&
	      !sfd__h2230[60] &&
	      !sfd__h2230[59] &&
	      !sfd__h2230[58] &&
	      !sfd__h2230[57] &&
	      !sfd__h2230[56] &&
	      !sfd__h2230[55] &&
	      !sfd__h2230[54] &&
	      !sfd__h2230[53] &&
	      !sfd__h2230[52] &&
	      !sfd__h2230[51] &&
	      !sfd__h2230[50] &&
	      !sfd__h2230[49] &&
	      !sfd__h2230[48] &&
	      !sfd__h2230[47] &&
	      !sfd__h2230[46] &&
	      !sfd__h2230[45] &&
	      !sfd__h2230[44] &&
	      !sfd__h2230[43] &&
	      !sfd__h2230[42] &&
	      !sfd__h2230[41] &&
	      !sfd__h2230[40] &&
	      !sfd__h2230[39] &&
	      !sfd__h2230[38] &&
	      !sfd__h2230[37] &&
	      !sfd__h2230[36] &&
	      !sfd__h2230[35] &&
	      !sfd__h2230[34] &&
	      !sfd__h2230[33] &&
	      !sfd__h2230[32] &&
	      !sfd__h2230[31] &&
	      !sfd__h2230[30] &&
	      !sfd__h2230[29] &&
	      !sfd__h2230[28] &&
	      !sfd__h2230[27] &&
	      !sfd__h2230[26] &&
	      !sfd__h2230[25] &&
	      !sfd__h2230[24] &&
	      !sfd__h2230[23] &&
	      !sfd__h2230[22] &&
	      !sfd__h2230[21] &&
	      !sfd__h2230[20] &&
	      !sfd__h2230[19] &&
	      !sfd__h2230[18] &&
	      !sfd__h2230[17] &&
	      !sfd__h2230[16] &&
	      !sfd__h2230[15] &&
	      !sfd__h2230[14] &&
	      !sfd__h2230[13] &&
	      !sfd__h2230[12] &&
	      !sfd__h2230[11] &&
	      !sfd__h2230[10] &&
	      !sfd__h2230[9] &&
	      !sfd__h2230[8] &&
	      !sfd__h2230[7] &&
	      !sfd__h2230[6] &&
	      !sfd__h2230[5] &&
	      !sfd__h2230[4] &&
	      !sfd__h2230[3] &&
	      !sfd__h2230[2] &&
	      !sfd__h2230[1] &&
	      !sfd__h2230[0]) ?
	       8'd0 :
	       _theResult___snd_fst_exp__h12923 ;
  assign IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d1676 =
	     sV1_exp__h823 == 8'd255 && sV1_sfd__h824 != 23'd0 ||
	     (requestR[191:160] != 32'hFFFFFFFF || !requestR[159]) &&
	     sV1_exp__h823 == 8'd255 &&
	     sV1_sfd__h824 == 23'd0 ;
  assign IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d1677 =
	     (requestR[191:160] == 32'hFFFFFFFF && requestR[159]) ?
	       64'h8000000000000000 :
	       64'h7FFFFFFFFFFFFFFF ;
  assign IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d1680 =
	     sV1_exp__h823 - 8'd127 ;
  assign IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d1689 =
	     (requestR[191:160] == 32'hFFFFFFFF && requestR[159]) ?
	       -b__h36799 :
	       b__h36799 ;
  assign IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d1809 =
	     (requestR[191:160] == 32'hFFFFFFFF && requestR[159]) ?
	       64'd0 :
	       ((sV1_exp__h823 == 8'd255 && sV1_sfd__h824 == 23'd0) ?
		  64'hFFFFFFFFFFFFFFFF :
		  IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_ETC___d1807) ;
  assign IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d1815 =
	     sV1_exp__h823 == 8'd255 && sV1_sfd__h824 == 23'd0 ||
	     (value_BIT_23___h161776 || sV1_sfd__h824 != 23'd0) &&
	     (NEG_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFF_ETC___d1778[19] ||
	      NEG_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFF_ETC___d1780 &&
	      IF_requestR_BITS_194_TO_192_0_EQ_0x0_1_OR_NOT__ETC___d1799 &&
	      x__h39015[88:25] == 64'hFFFFFFFFFFFFFFFF) ;
  assign IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d1827 =
	     { sV1_exp__h823 == 8'd255 && sV1_sfd__h824 != 23'd0 ||
	       IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d1815,
	       3'd0,
	       (sV1_exp__h823 != 8'd255 || sV1_sfd__h824 == 23'd0) &&
	       (sV1_exp__h823 != 8'd255 || sV1_sfd__h824 != 23'd0) &&
	       NOT_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFF_ETC___d1821 } ==
	     5'd0 ||
	     sV1_exp__h823 == 8'd255 && sV1_sfd__h824 != 23'd0 ||
	     IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d1815 ;
  assign IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d1828 =
	     (requestR[191:160] == 32'hFFFFFFFF && requestR[159]) ?
	       IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d1827 :
	       sV1_exp__h823 == 8'd255 && sV1_sfd__h824 != 23'd0 ||
	       IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d1815 ;
  assign IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d1834 =
	     (requestR[191:160] == 32'hFFFFFFFF && requestR[159]) ?
	       32'h80000000 :
	       32'h7FFFFFFF ;
  assign IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d1838 =
	     (requestR[191:160] == 32'hFFFFFFFF && requestR[159]) ?
	       -b__h39582 :
	       b__h39582 ;
  assign IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d19 =
	     (requestR[191:160] == 32'hFFFFFFFF) ?
	       requestR[158:128] :
	       31'h7FC00000 ;
  assign IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d1953 =
	     (requestR[191:160] == 32'hFFFFFFFF && requestR[159]) ?
	       32'd0 :
	       ((sV1_exp__h823 == 8'd255 && sV1_sfd__h824 == 23'd0) ?
		  32'hFFFFFFFF :
		  IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_ETC___d1951) ;
  assign IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d1960 =
	     sV1_exp__h823 == 8'd255 && sV1_sfd__h824 == 23'd0 ||
	     (value_BIT_23___h161776 || sV1_sfd__h824 != 23'd0) &&
	     (NEG_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFF_ETC___d1922[19] ||
	      NEG_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFF_ETC___d1924 &&
	      IF_requestR_BITS_194_TO_192_0_EQ_0x0_1_OR_NOT__ETC___d1943 &&
	      x__h41336[56:25] == 32'hFFFFFFFF) ;
  assign IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d1972 =
	     { sV1_exp__h823 == 8'd255 && sV1_sfd__h824 != 23'd0 ||
	       IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d1960,
	       3'd0,
	       (sV1_exp__h823 != 8'd255 || sV1_sfd__h824 == 23'd0) &&
	       (sV1_exp__h823 != 8'd255 || sV1_sfd__h824 != 23'd0) &&
	       NOT_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFF_ETC___d1966 } ==
	     5'd0 ||
	     sV1_exp__h823 == 8'd255 && sV1_sfd__h824 != 23'd0 ||
	     IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d1960 ;
  assign IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d1973 =
	     (requestR[191:160] == 32'hFFFFFFFF && requestR[159]) ?
	       IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d1972 :
	       sV1_exp__h823 == 8'd255 && sV1_sfd__h824 != 23'd0 ||
	       IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d1960 ;
  assign IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d1995 =
	     sV1_exp__h823 == 8'd255 && sV1_sfd__h824 != 23'd0 &&
	     !sV1_sfd__h824[22] &&
	     sV2_exp__h926 == 8'd255 &&
	     sV2_sfd__h927 != 23'd0 &&
	     !sV2_sfd__h927[22] ;
  assign IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d2005 =
	     sV1_exp__h823 == 8'd0 && sV1_sfd__h824 == 23'd0 &&
	     requestR[191:160] == 32'hFFFFFFFF &&
	     requestR[159] &&
	     sV2_exp__h926 == 8'd0 &&
	     sV2_sfd__h927 == 23'd0 &&
	     (requestR[127:96] != 32'hFFFFFFFF || !requestR[95]) ;
  assign IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d2018 =
	     sV1_exp__h823 < sV2_exp__h926 ;
  assign IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d2019 =
	     sV1_exp__h823 == sV2_exp__h926 ;
  assign IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d2020 =
	     sV1_sfd__h824 < sV2_sfd__h927 ;
  assign IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d2023 =
	     sV1_exp__h823 <= sV2_exp__h926 ;
  assign IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d2025 =
	     sV1_sfd__h824 <= sV2_sfd__h927 ;
  assign IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d2043 =
	     sV1_exp__h823 == 8'd255 && sV1_sfd__h824 != 23'd0 &&
	     !sV1_sfd__h824[22] ||
	     sV2_exp__h926 == 8'd255 && sV2_sfd__h927 != 23'd0 &&
	     !sV2_sfd__h927[22] ;
  assign IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d2080 =
	     IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d2043 ||
	     sV1_exp__h823 == 8'd255 && sV1_sfd__h824[22] ||
	     sV2_exp__h926 == 8'd255 && sV2_sfd__h927[22] ;
  assign IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d2091 =
	     IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d2023 &&
	     (!IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d2019 ||
	      IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d2025) &&
	     !IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d2018 &&
	     (!IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d2019 ||
	      !IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d2020) ;
  assign IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d2095 =
	     sV1_exp__h823 == 8'd0 && sV1_sfd__h824 == 23'd0 &&
	     sV2_exp__h926 == 8'd0 &&
	     sV2_sfd__h927 == 23'd0 ||
	     NOT_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5_ETC___d2094 ;
  assign IF_requestR_BITS_194_TO_192_0_EQ_0x0_1_OR_NOT__ETC___d1706 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       ((guard__h36732 == 2'b10) ?
		  IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d1689[24] :
		  guard__h36732 == 2'b11) :
	       ((requestR[194:192] == 3'h3) ?
		  guard__h36732 != 2'd0 :
		  requestR[194:192] == 3'h1 &&
		  IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d1689[88] &&
		  guard__h36732 != 2'd0) ;
  assign IF_requestR_BITS_194_TO_192_0_EQ_0x0_1_OR_NOT__ETC___d1738 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       ((guard__h37510 == 2'b10) ?
		  x__h37699[25] :
		  guard__h37510 == 2'b11) :
	       ((requestR[194:192] == 3'h3) ?
		  guard__h37510 != 2'd0 :
		  requestR[194:192] == 3'h1 && x__h37699[88] &&
		  guard__h37510 != 2'd0) ;
  assign IF_requestR_BITS_194_TO_192_0_EQ_0x0_1_OR_NOT__ETC___d1799 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       ((guard__h38794 == 2'b10) ?
		  x__h39015[25] :
		  guard__h38794 == 2'b11) :
	       requestR[194:192] == 3'h3 && guard__h38794 != 2'd0 ;
  assign IF_requestR_BITS_194_TO_192_0_EQ_0x0_1_OR_NOT__ETC___d1855 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       ((guard__h39515 == 2'b10) ?
		  IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d1838[24] :
		  guard__h39515 == 2'b11) :
	       ((requestR[194:192] == 3'h3) ?
		  guard__h39515 != 2'd0 :
		  requestR[194:192] == 3'h1 &&
		  IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d1838[56] &&
		  guard__h39515 != 2'd0) ;
  assign IF_requestR_BITS_194_TO_192_0_EQ_0x0_1_OR_NOT__ETC___d1887 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       ((guard__h40069 == 2'b10) ?
		  x__h40258[25] :
		  guard__h40069 == 2'b11) :
	       ((requestR[194:192] == 3'h3) ?
		  guard__h40069 != 2'd0 :
		  requestR[194:192] == 3'h1 && x__h40258[56] &&
		  guard__h40069 != 2'd0) ;
  assign IF_requestR_BITS_194_TO_192_0_EQ_0x0_1_OR_NOT__ETC___d1943 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       ((guard__h41115 == 2'b10) ?
		  x__h41336[25] :
		  guard__h41115 == 2'b11) :
	       requestR[194:192] == 3'h3 && guard__h41115 != 2'd0 ;
  assign IF_requestR_BITS_194_TO_192_0_EQ_0x0_1_OR_NOT__ETC___d2637 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       ((guard__h72055 == 2'b10) ?
		  IF_requestR_BIT_191_27_THEN_NEG_0b0_CONCAT_NOT_ETC___d2620[53] :
		  guard__h72055 == 2'b11) :
	       ((requestR[194:192] == 3'h3) ?
		  guard__h72055 != 2'd0 :
		  requestR[194:192] == 3'h1 &&
		  IF_requestR_BIT_191_27_THEN_NEG_0b0_CONCAT_NOT_ETC___d2620[85] &&
		  guard__h72055 != 2'd0) ;
  assign IF_requestR_BITS_194_TO_192_0_EQ_0x0_1_OR_NOT__ETC___d2669 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       ((guard__h72609 == 2'b10) ?
		  x__h72798[54] :
		  guard__h72609 == 2'b11) :
	       ((requestR[194:192] == 3'h3) ?
		  guard__h72609 != 2'd0 :
		  requestR[194:192] == 3'h1 && x__h72798[85] &&
		  guard__h72609 != 2'd0) ;
  assign IF_requestR_BITS_194_TO_192_0_EQ_0x0_1_OR_NOT__ETC___d2731 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       ((guard__h73655 == 2'b10) ?
		  x__h73876[54] :
		  guard__h73655 == 2'b11) :
	       requestR[194:192] == 3'h3 && guard__h73655 != 2'd0 ;
  assign IF_requestR_BITS_194_TO_192_0_EQ_0x0_1_OR_NOT__ETC___d3126 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       ((guard__h96909 == 2'b10) ?
		  IF_requestR_BIT_191_27_THEN_NEG_0b0_CONCAT_NOT_ETC___d3109[53] :
		  guard__h96909 == 2'b11) :
	       ((requestR[194:192] == 3'h3) ?
		  guard__h96909 != 2'd0 :
		  requestR[194:192] == 3'h1 &&
		  IF_requestR_BIT_191_27_THEN_NEG_0b0_CONCAT_NOT_ETC___d3109[117] &&
		  guard__h96909 != 2'd0) ;
  assign IF_requestR_BITS_194_TO_192_0_EQ_0x0_1_OR_NOT__ETC___d3158 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       ((guard__h97687 == 2'b10) ?
		  x__h97876[54] :
		  guard__h97687 == 2'b11) :
	       ((requestR[194:192] == 3'h3) ?
		  guard__h97687 != 2'd0 :
		  requestR[194:192] == 3'h1 && x__h97876[117] &&
		  guard__h97687 != 2'd0) ;
  assign IF_requestR_BITS_194_TO_192_0_EQ_0x0_1_OR_NOT__ETC___d3213 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       ((guard__h98954 == 2'b10) ?
		  x__h99175[54] :
		  guard__h98954 == 2'b11) :
	       requestR[194:192] == 3'h3 && guard__h98954 != 2'd0 ;
  assign IF_requestR_BIT_159_6_THEN_0_ELSE_IF_requestR__ETC___d1507 =
	     requestR[159] ?
	       6'd0 :
	       (requestR[158] ?
		  6'd1 :
		  (requestR[157] ?
		     6'd2 :
		     (requestR[156] ?
			6'd3 :
			(requestR[155] ?
			   6'd4 :
			   (requestR[154] ?
			      6'd5 :
			      (requestR[153] ?
				 6'd6 :
				 (requestR[152] ?
				    6'd7 :
				    (requestR[151] ?
				       6'd8 :
				       (requestR[150] ?
					  6'd9 :
					  (requestR[149] ?
					     6'd10 :
					     (requestR[148] ?
						6'd11 :
						(requestR[147] ?
						   6'd12 :
						   (requestR[146] ?
						      6'd13 :
						      (requestR[145] ?
							 6'd14 :
							 (requestR[144] ?
							    6'd15 :
							    (requestR[143] ?
							       6'd16 :
							       (requestR[142] ?
								  6'd17 :
								  (requestR[141] ?
								     6'd18 :
								     (requestR[140] ?
									6'd19 :
									(requestR[139] ?
									   6'd20 :
									   (requestR[138] ?
									      6'd21 :
									      (requestR[137] ?
										 6'd22 :
										 (requestR[136] ?
										    6'd23 :
										    (requestR[135] ?
										       6'd24 :
										       (requestR[134] ?
											  6'd25 :
											  (requestR[133] ?
											     6'd26 :
											     (requestR[132] ?
												6'd27 :
												(requestR[131] ?
												   6'd28 :
												   (requestR[130] ?
												      6'd29 :
												      (requestR[129] ?
													 6'd30 :
													 (requestR[128] ?
													    6'd31 :
													    6'd32))))))))))))))))))))))))))))))) ;
  assign IF_requestR_BIT_159_6_THEN_0_ELSE_IF_requestR__ETC___d2445 =
	     requestR[159] ?
	       6'd0 :
	       (requestR[158] ?
		  6'd1 :
		  (requestR[157] ?
		     6'd2 :
		     (requestR[156] ?
			6'd3 :
			(requestR[155] ?
			   6'd4 :
			   (requestR[154] ?
			      6'd5 :
			      (requestR[153] ?
				 6'd6 :
				 (requestR[152] ?
				    6'd7 :
				    (requestR[151] ?
				       6'd8 :
				       (requestR[150] ?
					  6'd9 :
					  (requestR[149] ?
					     6'd10 :
					     (requestR[148] ?
						6'd11 :
						(requestR[147] ?
						   6'd12 :
						   (requestR[146] ?
						      6'd13 :
						      (requestR[145] ?
							 6'd14 :
							 (requestR[144] ?
							    6'd15 :
							    (requestR[143] ?
							       6'd16 :
							       (requestR[142] ?
								  6'd17 :
								  (requestR[141] ?
								     6'd18 :
								     (requestR[140] ?
									6'd19 :
									(requestR[139] ?
									   6'd20 :
									   (requestR[138] ?
									      6'd21 :
									      (requestR[137] ?
										 6'd22 :
										 (requestR[136] ?
										    6'd23 :
										    (requestR[135] ?
										       6'd24 :
										       (requestR[134] ?
											  6'd25 :
											  (requestR[133] ?
											     6'd26 :
											     (requestR[132] ?
												6'd27 :
												(requestR[131] ?
												   6'd28 :
												   (requestR[130] ?
												      6'd29 :
												      (requestR[129] ?
													 6'd30 :
													 (requestR[128] ?
													    6'd31 :
													    6'd55))))))))))))))))))))))))))))))) ;
  assign IF_requestR_BIT_159_6_THEN_NEG_requestR_BITS_1_ETC___d1454 =
	     (sfd__h23980[31] || sfd__h23980[30] || sfd__h23980[29] ||
	      sfd__h23980[28] ||
	      sfd__h23980[27] ||
	      sfd__h23980[26] ||
	      sfd__h23980[25] ||
	      sfd__h23980[24] ||
	      sfd__h23980[23] ||
	      sfd__h23980[22] ||
	      sfd__h23980[21] ||
	      sfd__h23980[20] ||
	      sfd__h23980[19] ||
	      sfd__h23980[18] ||
	      sfd__h23980[17] ||
	      sfd__h23980[16] ||
	      sfd__h23980[15] ||
	      sfd__h23980[14] ||
	      sfd__h23980[13] ||
	      sfd__h23980[12] ||
	      sfd__h23980[11] ||
	      sfd__h23980[10] ||
	      sfd__h23980[9] ||
	      sfd__h23980[8] ||
	      sfd__h23980[7] ||
	      sfd__h23980[6] ||
	      sfd__h23980[5] ||
	      sfd__h23980[4] ||
	      sfd__h23980[3] ||
	      sfd__h23980[2] ||
	      sfd__h23980[1] ||
	      sfd__h23980[0]) &&
	     (!_32_MINUS_0_CONCAT_IF_IF_requestR_BIT_159_6_THE_ETC___d1256 ||
	      !_32_MINUS_0_CONCAT_IF_IF_requestR_BIT_159_6_THE_ETC___d1258 &&
	      !_32_MINUS_0_CONCAT_IF_IF_requestR_BIT_159_6_THE_ETC___d1261 &&
	      _theResult___fst_exp__h29960 == 8'd255 &&
	      _theResult___fst_sfd__h29961 == 23'd0) ;
  assign IF_requestR_BIT_159_6_THEN_NEG_requestR_BITS_1_ETC___d1457 =
	     (sfd__h23980[31] || sfd__h23980[30] || sfd__h23980[29] ||
	      sfd__h23980[28] ||
	      sfd__h23980[27] ||
	      sfd__h23980[26] ||
	      sfd__h23980[25] ||
	      sfd__h23980[24] ||
	      sfd__h23980[23] ||
	      sfd__h23980[22] ||
	      sfd__h23980[21] ||
	      sfd__h23980[20] ||
	      sfd__h23980[19] ||
	      sfd__h23980[18] ||
	      sfd__h23980[17] ||
	      sfd__h23980[16] ||
	      sfd__h23980[15] ||
	      sfd__h23980[14] ||
	      sfd__h23980[13] ||
	      sfd__h23980[12] ||
	      sfd__h23980[11] ||
	      sfd__h23980[10] ||
	      sfd__h23980[9] ||
	      sfd__h23980[8] ||
	      sfd__h23980[7] ||
	      sfd__h23980[6] ||
	      sfd__h23980[5] ||
	      sfd__h23980[4] ||
	      sfd__h23980[3] ||
	      sfd__h23980[2] ||
	      sfd__h23980[1] ||
	      sfd__h23980[0]) &&
	     _32_MINUS_0_CONCAT_IF_IF_requestR_BIT_159_6_THE_ETC___d1256 &&
	     _32_MINUS_0_CONCAT_IF_IF_requestR_BIT_159_6_THE_ETC___d1258 ;
  assign IF_requestR_BIT_159_6_THEN_NEG_requestR_BITS_1_ETC___d1466 =
	     (sfd__h23980[31] || sfd__h23980[30] || sfd__h23980[29] ||
	      sfd__h23980[28] ||
	      sfd__h23980[27] ||
	      sfd__h23980[26] ||
	      sfd__h23980[25] ||
	      sfd__h23980[24] ||
	      sfd__h23980[23] ||
	      sfd__h23980[22] ||
	      sfd__h23980[21] ||
	      sfd__h23980[20] ||
	      sfd__h23980[19] ||
	      sfd__h23980[18] ||
	      sfd__h23980[17] ||
	      sfd__h23980[16] ||
	      sfd__h23980[15] ||
	      sfd__h23980[14] ||
	      sfd__h23980[13] ||
	      sfd__h23980[12] ||
	      sfd__h23980[11] ||
	      sfd__h23980[10] ||
	      sfd__h23980[9] ||
	      sfd__h23980[8] ||
	      sfd__h23980[7] ||
	      sfd__h23980[6] ||
	      sfd__h23980[5] ||
	      sfd__h23980[4] ||
	      sfd__h23980[3] ||
	      sfd__h23980[2] ||
	      sfd__h23980[1] ||
	      sfd__h23980[0]) &&
	     _32_MINUS_0_CONCAT_IF_IF_requestR_BIT_159_6_THE_ETC___d1256 &&
	     !_32_MINUS_0_CONCAT_IF_IF_requestR_BIT_159_6_THE_ETC___d1258 &&
	     IF_32_MINUS_0_CONCAT_IF_IF_requestR_BIT_159_6__ETC___d1463 ;
  assign IF_requestR_BIT_191_27_THEN_0_ELSE_IF_requestR_ETC___d901 =
	     requestR[191] ?
	       7'd0 :
	       (requestR[190] ?
		  7'd1 :
		  (requestR[189] ?
		     7'd2 :
		     (requestR[188] ?
			7'd3 :
			(requestR[187] ?
			   7'd4 :
			   (requestR[186] ?
			      7'd5 :
			      (requestR[185] ?
				 7'd6 :
				 (requestR[184] ?
				    7'd7 :
				    (requestR[183] ?
				       7'd8 :
				       (requestR[182] ?
					  7'd9 :
					  (requestR[181] ?
					     7'd10 :
					     (requestR[180] ?
						7'd11 :
						(requestR[179] ?
						   7'd12 :
						   (requestR[178] ?
						      7'd13 :
						      (requestR[177] ?
							 7'd14 :
							 (requestR[176] ?
							    7'd15 :
							    (requestR[175] ?
							       7'd16 :
							       (requestR[174] ?
								  7'd17 :
								  (requestR[173] ?
								     7'd18 :
								     (requestR[172] ?
									7'd19 :
									(requestR[171] ?
									   7'd20 :
									   (requestR[170] ?
									      7'd21 :
									      (requestR[169] ?
										 7'd22 :
										 (requestR[168] ?
										    7'd23 :
										    (requestR[167] ?
										       7'd24 :
										       (requestR[166] ?
											  7'd25 :
											  (requestR[165] ?
											     7'd26 :
											     (requestR[164] ?
												7'd27 :
												(requestR[163] ?
												   7'd28 :
												   (requestR[162] ?
												      7'd29 :
												      (requestR[161] ?
													 7'd30 :
													 (requestR[160] ?
													    7'd31 :
													    (requestR[159] ?
													       7'd32 :
													       (requestR[158] ?
														  7'd33 :
														  (requestR[157] ?
														     7'd34 :
														     (requestR[156] ?
															7'd35 :
															(requestR[155] ?
															   7'd36 :
															   (requestR[154] ?
															      7'd37 :
															      (requestR[153] ?
																 7'd38 :
																 (requestR[152] ?
																    7'd39 :
																    (requestR[151] ?
																       7'd40 :
																       (requestR[150] ?
																	  7'd41 :
																	  (requestR[149] ?
																	     7'd42 :
																	     (requestR[148] ?
																		7'd43 :
																		(requestR[147] ?
																		   7'd44 :
																		   (requestR[146] ?
																		      7'd45 :
																		      (requestR[145] ?
																			 7'd46 :
																			 (requestR[144] ?
																			    7'd47 :
																			    (requestR[143] ?
																			       7'd48 :
																			       (requestR[142] ?
																				  7'd49 :
																				  (requestR[141] ?
																				     7'd50 :
																				     (requestR[140] ?
																					7'd51 :
																					(requestR[139] ?
																					   7'd52 :
																					   (requestR[138] ?
																					      7'd53 :
																					      (requestR[137] ?
																						 7'd54 :
																						 (requestR[136] ?
																						    7'd55 :
																						    (requestR[135] ?
																						       7'd56 :
																						       (requestR[134] ?
																							  7'd57 :
																							  (requestR[133] ?
																							     7'd58 :
																							     (requestR[132] ?
																								7'd59 :
																								(requestR[131] ?
																								   7'd60 :
																								   (requestR[130] ?
																								      7'd61 :
																								      (requestR[129] ?
																									 7'd62 :
																									 (requestR[128] ?
																									    7'd63 :
																									    7'd64))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) ;
  assign IF_requestR_BIT_191_27_THEN_2147483648_ELSE_21_ETC___d2608 =
	     requestR[191] ? 32'h80000000 : 32'h7FFFFFFF ;
  assign IF_requestR_BIT_191_27_THEN_922337203685477580_ETC___d3105 =
	     requestR[191] ? 64'h8000000000000000 : 64'h7FFFFFFFFFFFFFFF ;
  assign IF_requestR_BIT_191_27_THEN_NEG_0b0_CONCAT_NOT_ETC___d2620 =
	     requestR[191] ? -b__h72122 : b__h72122 ;
  assign IF_requestR_BIT_191_27_THEN_NEG_0b0_CONCAT_NOT_ETC___d3109 =
	     requestR[191] ? -b__h96976 : b__h96976 ;
  assign IF_requestR_BIT_191_27_THEN_NEG_requestR_BITS__ETC___d2932 =
	     (sfd__h2230[63] || sfd__h2230[62] || sfd__h2230[61] ||
	      sfd__h2230[60] ||
	      sfd__h2230[59] ||
	      sfd__h2230[58] ||
	      sfd__h2230[57] ||
	      sfd__h2230[56] ||
	      sfd__h2230[55] ||
	      sfd__h2230[54] ||
	      sfd__h2230[53] ||
	      sfd__h2230[52] ||
	      sfd__h2230[51] ||
	      sfd__h2230[50] ||
	      sfd__h2230[49] ||
	      sfd__h2230[48] ||
	      sfd__h2230[47] ||
	      sfd__h2230[46] ||
	      sfd__h2230[45] ||
	      sfd__h2230[44] ||
	      sfd__h2230[43] ||
	      sfd__h2230[42] ||
	      sfd__h2230[41] ||
	      sfd__h2230[40] ||
	      sfd__h2230[39] ||
	      sfd__h2230[38] ||
	      sfd__h2230[37] ||
	      sfd__h2230[36] ||
	      sfd__h2230[35] ||
	      sfd__h2230[34] ||
	      sfd__h2230[33] ||
	      sfd__h2230[32] ||
	      sfd__h2230[31] ||
	      sfd__h2230[30] ||
	      sfd__h2230[29] ||
	      sfd__h2230[28] ||
	      sfd__h2230[27] ||
	      sfd__h2230[26] ||
	      sfd__h2230[25] ||
	      sfd__h2230[24] ||
	      sfd__h2230[23] ||
	      sfd__h2230[22] ||
	      sfd__h2230[21] ||
	      sfd__h2230[20] ||
	      sfd__h2230[19] ||
	      sfd__h2230[18] ||
	      sfd__h2230[17] ||
	      sfd__h2230[16] ||
	      sfd__h2230[15] ||
	      sfd__h2230[14] ||
	      sfd__h2230[13] ||
	      sfd__h2230[12] ||
	      sfd__h2230[11] ||
	      sfd__h2230[10] ||
	      sfd__h2230[9] ||
	      sfd__h2230[8] ||
	      sfd__h2230[7] ||
	      sfd__h2230[6] ||
	      sfd__h2230[5] ||
	      sfd__h2230[4] ||
	      sfd__h2230[3] ||
	      sfd__h2230[2] ||
	      sfd__h2230[1] ||
	      sfd__h2230[0]) &&
	     (!_64_MINUS_0_CONCAT_IF_IF_requestR_BIT_191_27_TH_ETC___d2770 ||
	      !_64_MINUS_0_CONCAT_IF_IF_requestR_BIT_191_27_TH_ETC___d2772 &&
	      !_64_MINUS_0_CONCAT_IF_IF_requestR_BIT_191_27_TH_ETC___d2775 &&
	      _theResult___fst_exp__h85300 == 11'd2047 &&
	      _theResult___fst_sfd__h85301 == 52'd0) ;
  assign IF_requestR_BIT_191_27_THEN_NEG_requestR_BITS__ETC___d2935 =
	     (sfd__h2230[63] || sfd__h2230[62] || sfd__h2230[61] ||
	      sfd__h2230[60] ||
	      sfd__h2230[59] ||
	      sfd__h2230[58] ||
	      sfd__h2230[57] ||
	      sfd__h2230[56] ||
	      sfd__h2230[55] ||
	      sfd__h2230[54] ||
	      sfd__h2230[53] ||
	      sfd__h2230[52] ||
	      sfd__h2230[51] ||
	      sfd__h2230[50] ||
	      sfd__h2230[49] ||
	      sfd__h2230[48] ||
	      sfd__h2230[47] ||
	      sfd__h2230[46] ||
	      sfd__h2230[45] ||
	      sfd__h2230[44] ||
	      sfd__h2230[43] ||
	      sfd__h2230[42] ||
	      sfd__h2230[41] ||
	      sfd__h2230[40] ||
	      sfd__h2230[39] ||
	      sfd__h2230[38] ||
	      sfd__h2230[37] ||
	      sfd__h2230[36] ||
	      sfd__h2230[35] ||
	      sfd__h2230[34] ||
	      sfd__h2230[33] ||
	      sfd__h2230[32] ||
	      sfd__h2230[31] ||
	      sfd__h2230[30] ||
	      sfd__h2230[29] ||
	      sfd__h2230[28] ||
	      sfd__h2230[27] ||
	      sfd__h2230[26] ||
	      sfd__h2230[25] ||
	      sfd__h2230[24] ||
	      sfd__h2230[23] ||
	      sfd__h2230[22] ||
	      sfd__h2230[21] ||
	      sfd__h2230[20] ||
	      sfd__h2230[19] ||
	      sfd__h2230[18] ||
	      sfd__h2230[17] ||
	      sfd__h2230[16] ||
	      sfd__h2230[15] ||
	      sfd__h2230[14] ||
	      sfd__h2230[13] ||
	      sfd__h2230[12] ||
	      sfd__h2230[11] ||
	      sfd__h2230[10] ||
	      sfd__h2230[9] ||
	      sfd__h2230[8] ||
	      sfd__h2230[7] ||
	      sfd__h2230[6] ||
	      sfd__h2230[5] ||
	      sfd__h2230[4] ||
	      sfd__h2230[3] ||
	      sfd__h2230[2] ||
	      sfd__h2230[1] ||
	      sfd__h2230[0]) &&
	     _64_MINUS_0_CONCAT_IF_IF_requestR_BIT_191_27_TH_ETC___d2770 &&
	     _64_MINUS_0_CONCAT_IF_IF_requestR_BIT_191_27_TH_ETC___d2772 ;
  assign IF_requestR_BIT_191_27_THEN_NEG_requestR_BITS__ETC___d2944 =
	     (sfd__h2230[63] || sfd__h2230[62] || sfd__h2230[61] ||
	      sfd__h2230[60] ||
	      sfd__h2230[59] ||
	      sfd__h2230[58] ||
	      sfd__h2230[57] ||
	      sfd__h2230[56] ||
	      sfd__h2230[55] ||
	      sfd__h2230[54] ||
	      sfd__h2230[53] ||
	      sfd__h2230[52] ||
	      sfd__h2230[51] ||
	      sfd__h2230[50] ||
	      sfd__h2230[49] ||
	      sfd__h2230[48] ||
	      sfd__h2230[47] ||
	      sfd__h2230[46] ||
	      sfd__h2230[45] ||
	      sfd__h2230[44] ||
	      sfd__h2230[43] ||
	      sfd__h2230[42] ||
	      sfd__h2230[41] ||
	      sfd__h2230[40] ||
	      sfd__h2230[39] ||
	      sfd__h2230[38] ||
	      sfd__h2230[37] ||
	      sfd__h2230[36] ||
	      sfd__h2230[35] ||
	      sfd__h2230[34] ||
	      sfd__h2230[33] ||
	      sfd__h2230[32] ||
	      sfd__h2230[31] ||
	      sfd__h2230[30] ||
	      sfd__h2230[29] ||
	      sfd__h2230[28] ||
	      sfd__h2230[27] ||
	      sfd__h2230[26] ||
	      sfd__h2230[25] ||
	      sfd__h2230[24] ||
	      sfd__h2230[23] ||
	      sfd__h2230[22] ||
	      sfd__h2230[21] ||
	      sfd__h2230[20] ||
	      sfd__h2230[19] ||
	      sfd__h2230[18] ||
	      sfd__h2230[17] ||
	      sfd__h2230[16] ||
	      sfd__h2230[15] ||
	      sfd__h2230[14] ||
	      sfd__h2230[13] ||
	      sfd__h2230[12] ||
	      sfd__h2230[11] ||
	      sfd__h2230[10] ||
	      sfd__h2230[9] ||
	      sfd__h2230[8] ||
	      sfd__h2230[7] ||
	      sfd__h2230[6] ||
	      sfd__h2230[5] ||
	      sfd__h2230[4] ||
	      sfd__h2230[3] ||
	      sfd__h2230[2] ||
	      sfd__h2230[1] ||
	      sfd__h2230[0]) &&
	     _64_MINUS_0_CONCAT_IF_IF_requestR_BIT_191_27_TH_ETC___d2770 &&
	     !_64_MINUS_0_CONCAT_IF_IF_requestR_BIT_191_27_TH_ETC___d2772 &&
	     IF_64_MINUS_0_CONCAT_IF_IF_requestR_BIT_191_27_ETC___d2941 ;
  assign IF_requestR_BIT_191_27_THEN_NEG_requestR_BITS__ETC___d627 =
	     (sfd__h2230[63] || sfd__h2230[62] || sfd__h2230[61] ||
	      sfd__h2230[60] ||
	      sfd__h2230[59] ||
	      sfd__h2230[58] ||
	      sfd__h2230[57] ||
	      sfd__h2230[56] ||
	      sfd__h2230[55] ||
	      sfd__h2230[54] ||
	      sfd__h2230[53] ||
	      sfd__h2230[52] ||
	      sfd__h2230[51] ||
	      sfd__h2230[50] ||
	      sfd__h2230[49] ||
	      sfd__h2230[48] ||
	      sfd__h2230[47] ||
	      sfd__h2230[46] ||
	      sfd__h2230[45] ||
	      sfd__h2230[44] ||
	      sfd__h2230[43] ||
	      sfd__h2230[42] ||
	      sfd__h2230[41] ||
	      sfd__h2230[40] ||
	      sfd__h2230[39] ||
	      sfd__h2230[38] ||
	      sfd__h2230[37] ||
	      sfd__h2230[36] ||
	      sfd__h2230[35] ||
	      sfd__h2230[34] ||
	      sfd__h2230[33] ||
	      sfd__h2230[32] ||
	      sfd__h2230[31] ||
	      sfd__h2230[30] ||
	      sfd__h2230[29] ||
	      sfd__h2230[28] ||
	      sfd__h2230[27] ||
	      sfd__h2230[26] ||
	      sfd__h2230[25] ||
	      sfd__h2230[24] ||
	      sfd__h2230[23] ||
	      sfd__h2230[22] ||
	      sfd__h2230[21] ||
	      sfd__h2230[20] ||
	      sfd__h2230[19] ||
	      sfd__h2230[18] ||
	      sfd__h2230[17] ||
	      sfd__h2230[16] ||
	      sfd__h2230[15] ||
	      sfd__h2230[14] ||
	      sfd__h2230[13] ||
	      sfd__h2230[12] ||
	      sfd__h2230[11] ||
	      sfd__h2230[10] ||
	      sfd__h2230[9] ||
	      sfd__h2230[8] ||
	      sfd__h2230[7] ||
	      sfd__h2230[6] ||
	      sfd__h2230[5] ||
	      sfd__h2230[4] ||
	      sfd__h2230[3] ||
	      sfd__h2230[2] ||
	      sfd__h2230[1] ||
	      sfd__h2230[0]) &&
	     (!_64_MINUS_0_CONCAT_IF_IF_requestR_BIT_191_27_TH_ETC___d388 ||
	      !_64_MINUS_0_CONCAT_IF_IF_requestR_BIT_191_27_TH_ETC___d390 &&
	      !_64_MINUS_0_CONCAT_IF_IF_requestR_BIT_191_27_TH_ETC___d393 &&
	      _theResult___fst_exp__h12914 == 8'd255 &&
	      _theResult___fst_sfd__h12915 == 23'd0) ;
  assign IF_requestR_BIT_191_27_THEN_NEG_requestR_BITS__ETC___d630 =
	     (sfd__h2230[63] || sfd__h2230[62] || sfd__h2230[61] ||
	      sfd__h2230[60] ||
	      sfd__h2230[59] ||
	      sfd__h2230[58] ||
	      sfd__h2230[57] ||
	      sfd__h2230[56] ||
	      sfd__h2230[55] ||
	      sfd__h2230[54] ||
	      sfd__h2230[53] ||
	      sfd__h2230[52] ||
	      sfd__h2230[51] ||
	      sfd__h2230[50] ||
	      sfd__h2230[49] ||
	      sfd__h2230[48] ||
	      sfd__h2230[47] ||
	      sfd__h2230[46] ||
	      sfd__h2230[45] ||
	      sfd__h2230[44] ||
	      sfd__h2230[43] ||
	      sfd__h2230[42] ||
	      sfd__h2230[41] ||
	      sfd__h2230[40] ||
	      sfd__h2230[39] ||
	      sfd__h2230[38] ||
	      sfd__h2230[37] ||
	      sfd__h2230[36] ||
	      sfd__h2230[35] ||
	      sfd__h2230[34] ||
	      sfd__h2230[33] ||
	      sfd__h2230[32] ||
	      sfd__h2230[31] ||
	      sfd__h2230[30] ||
	      sfd__h2230[29] ||
	      sfd__h2230[28] ||
	      sfd__h2230[27] ||
	      sfd__h2230[26] ||
	      sfd__h2230[25] ||
	      sfd__h2230[24] ||
	      sfd__h2230[23] ||
	      sfd__h2230[22] ||
	      sfd__h2230[21] ||
	      sfd__h2230[20] ||
	      sfd__h2230[19] ||
	      sfd__h2230[18] ||
	      sfd__h2230[17] ||
	      sfd__h2230[16] ||
	      sfd__h2230[15] ||
	      sfd__h2230[14] ||
	      sfd__h2230[13] ||
	      sfd__h2230[12] ||
	      sfd__h2230[11] ||
	      sfd__h2230[10] ||
	      sfd__h2230[9] ||
	      sfd__h2230[8] ||
	      sfd__h2230[7] ||
	      sfd__h2230[6] ||
	      sfd__h2230[5] ||
	      sfd__h2230[4] ||
	      sfd__h2230[3] ||
	      sfd__h2230[2] ||
	      sfd__h2230[1] ||
	      sfd__h2230[0]) &&
	     _64_MINUS_0_CONCAT_IF_IF_requestR_BIT_191_27_TH_ETC___d388 &&
	     _64_MINUS_0_CONCAT_IF_IF_requestR_BIT_191_27_TH_ETC___d390 ;
  assign IF_requestR_BIT_191_27_THEN_NEG_requestR_BITS__ETC___d639 =
	     (sfd__h2230[63] || sfd__h2230[62] || sfd__h2230[61] ||
	      sfd__h2230[60] ||
	      sfd__h2230[59] ||
	      sfd__h2230[58] ||
	      sfd__h2230[57] ||
	      sfd__h2230[56] ||
	      sfd__h2230[55] ||
	      sfd__h2230[54] ||
	      sfd__h2230[53] ||
	      sfd__h2230[52] ||
	      sfd__h2230[51] ||
	      sfd__h2230[50] ||
	      sfd__h2230[49] ||
	      sfd__h2230[48] ||
	      sfd__h2230[47] ||
	      sfd__h2230[46] ||
	      sfd__h2230[45] ||
	      sfd__h2230[44] ||
	      sfd__h2230[43] ||
	      sfd__h2230[42] ||
	      sfd__h2230[41] ||
	      sfd__h2230[40] ||
	      sfd__h2230[39] ||
	      sfd__h2230[38] ||
	      sfd__h2230[37] ||
	      sfd__h2230[36] ||
	      sfd__h2230[35] ||
	      sfd__h2230[34] ||
	      sfd__h2230[33] ||
	      sfd__h2230[32] ||
	      sfd__h2230[31] ||
	      sfd__h2230[30] ||
	      sfd__h2230[29] ||
	      sfd__h2230[28] ||
	      sfd__h2230[27] ||
	      sfd__h2230[26] ||
	      sfd__h2230[25] ||
	      sfd__h2230[24] ||
	      sfd__h2230[23] ||
	      sfd__h2230[22] ||
	      sfd__h2230[21] ||
	      sfd__h2230[20] ||
	      sfd__h2230[19] ||
	      sfd__h2230[18] ||
	      sfd__h2230[17] ||
	      sfd__h2230[16] ||
	      sfd__h2230[15] ||
	      sfd__h2230[14] ||
	      sfd__h2230[13] ||
	      sfd__h2230[12] ||
	      sfd__h2230[11] ||
	      sfd__h2230[10] ||
	      sfd__h2230[9] ||
	      sfd__h2230[8] ||
	      sfd__h2230[7] ||
	      sfd__h2230[6] ||
	      sfd__h2230[5] ||
	      sfd__h2230[4] ||
	      sfd__h2230[3] ||
	      sfd__h2230[2] ||
	      sfd__h2230[1] ||
	      sfd__h2230[0]) &&
	     _64_MINUS_0_CONCAT_IF_IF_requestR_BIT_191_27_TH_ETC___d388 &&
	     !_64_MINUS_0_CONCAT_IF_IF_requestR_BIT_191_27_TH_ETC___d390 &&
	     IF_64_MINUS_0_CONCAT_IF_IF_requestR_BIT_191_27_ETC___d636 ;
  assign IF_requestR_BIT_191_27_THEN_NOT_requestR_BITS__ETC___d5207 =
	     requestR[191] ?
	       !requestR_BITS_190_TO_180_599_ULE_requestR_BITS_ETC___d5196 ||
	       requestR_BITS_190_TO_180_599_EQ_requestR_BITS__ETC___d5198 &&
	       !requestR_BITS_179_TO_128_601_ULE_requestR_BITS_ETC___d5199 :
	       requestR_BITS_190_TO_180_599_ULT_requestR_BITS_ETC___d5203 ||
	       requestR_BITS_190_TO_180_599_EQ_requestR_BITS__ETC___d5198 &&
	       requestR_BITS_179_TO_128_601_ULT_requestR_BITS_ETC___d5204 ;
  assign IF_sfd___30277_BIT_1_THEN_2_ELSE_0__q68 =
	     sfd___3__h60277[1] ? 2'd2 : 2'd0 ;
  assign IF_sfd___30277_BIT_2_THEN_2_ELSE_0__q67 =
	     sfd___3__h60277[2] ? 2'd2 : 2'd0 ;
  assign IF_sfd___31835_BIT_10_THEN_2_ELSE_0__q9 =
	     sfd___3__h11835[10] ? 2'd2 : 2'd0 ;
  assign IF_sfd___31835_BIT_11_THEN_2_ELSE_0__q8 =
	     sfd___3__h11835[11] ? 2'd2 : 2'd0 ;
  assign IF_sfd___31835_BIT_39_THEN_2_ELSE_0__q7 =
	     sfd___3__h11835[39] ? 2'd2 : 2'd0 ;
  assign IF_sfd___31835_BIT_40_THEN_2_ELSE_0__q6 =
	     sfd___3__h11835[40] ? 2'd2 : 2'd0 ;
  assign IF_sfd___32457_BIT_10_THEN_2_ELSE_0__q25 =
	     sfd___3__h22457[10] ? 2'd2 : 2'd0 ;
  assign IF_sfd___32457_BIT_11_THEN_2_ELSE_0__q24 =
	     sfd___3__h22457[11] ? 2'd2 : 2'd0 ;
  assign IF_sfd___32457_BIT_39_THEN_2_ELSE_0__q23 =
	     sfd___3__h22457[39] ? 2'd2 : 2'd0 ;
  assign IF_sfd___32457_BIT_40_THEN_2_ELSE_0__q22 =
	     sfd___3__h22457[40] ? 2'd2 : 2'd0 ;
  assign IF_sfd___35055_BIT_7_THEN_2_ELSE_0__q53 =
	     sfd___3__h35055[7] ? 2'd2 : 2'd0 ;
  assign IF_sfd___35055_BIT_8_THEN_2_ELSE_0__q52 =
	     sfd___3__h35055[8] ? 2'd2 : 2'd0 ;
  assign IF_sfd___38884_BIT_7_THEN_2_ELSE_0__q39 =
	     sfd___3__h28884[7] ? 2'd2 : 2'd0 ;
  assign IF_sfd___38884_BIT_8_THEN_2_ELSE_0__q38 =
	     sfd___3__h28884[8] ? 2'd2 : 2'd0 ;
  assign IF_sfd___39973_BIT_1_THEN_2_ELSE_0__q82 =
	     sfd___3__h69973[1] ? 2'd2 : 2'd0 ;
  assign IF_sfd___39973_BIT_2_THEN_2_ELSE_0__q81 =
	     sfd___3__h69973[2] ? 2'd2 : 2'd0 ;
  assign IF_sfdin19458_BIT_33_THEN_2_ELSE_0__q115 =
	     sfdin__h119458[33] ? 2'd2 : 2'd0 ;
  assign IF_sfdin37311_BIT_33_THEN_2_ELSE_0__q120 =
	     sfdin__h137311[33] ? 2'd2 : 2'd0 ;
  assign IF_sfdin78646_BIT_4_THEN_2_ELSE_0__q152 =
	     sfdin__h178646[4] ? 2'd2 : 2'd0 ;
  assign IF_theResult___snd28101_BIT_33_THEN_2_ELSE_0__q117 =
	     _theResult___snd__h128101[33] ? 2'd2 : 2'd0 ;
  assign IF_theResult___snd45978_BIT_33_THEN_2_ELSE_0__q123 =
	     _theResult___snd__h145978[33] ? 2'd2 : 2'd0 ;
  assign IF_theResult___snd69030_BIT_4_THEN_2_ELSE_0__q149 =
	     _theResult___snd__h169030[4] ? 2'd2 : 2'd0 ;
  assign IF_theResult___snd87429_BIT_4_THEN_2_ELSE_0__q155 =
	     _theResult___snd__h187429[4] ? 2'd2 : 2'd0 ;
  assign IF_x0258_BIT_24_THEN_2_ELSE_0__q65 = x__h40258[24] ? 2'd2 : 2'd0 ;
  assign IF_x1336_BIT_24_THEN_2_ELSE_0__q66 = x__h41336[24] ? 2'd2 : 2'd0 ;
  assign IF_x2798_BIT_53_THEN_2_ELSE_0__q92 = x__h72798[53] ? 2'd2 : 2'd0 ;
  assign IF_x3876_BIT_53_THEN_2_ELSE_0__q93 = x__h73876[53] ? 2'd2 : 2'd0 ;
  assign IF_x7699_BIT_24_THEN_2_ELSE_0__q63 = x__h37699[24] ? 2'd2 : 2'd0 ;
  assign IF_x7876_BIT_53_THEN_2_ELSE_0__q112 = x__h97876[53] ? 2'd2 : 2'd0 ;
  assign IF_x9015_BIT_24_THEN_2_ELSE_0__q64 = x__h39015[24] ? 2'd2 : 2'd0 ;
  assign IF_x9175_BIT_53_THEN_2_ELSE_0__q113 = x__h99175[53] ? 2'd2 : 2'd0 ;
  assign NEG_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFF_ETC___d1682 =
	     -{ {12{IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d1680[7]}},
		IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d1680 } ;
  assign NEG_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFF_ETC___d1714 =
	     NEG_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFF_ETC___d1682 +
	     20'd64 ;
  assign NEG_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFF_ETC___d1715 =
	     NEG_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFF_ETC___d1714 -
	     20'd2 ;
  assign NEG_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFF_ETC___d1717 =
	     (NEG_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFF_ETC___d1715 ^
	      20'h80000) <=
	     20'd524352 ;
  assign NEG_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFF_ETC___d1778 =
	     NEG_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFF_ETC___d1714 -
	     20'd1 ;
  assign NEG_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFF_ETC___d1780 =
	     (NEG_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFF_ETC___d1778 ^
	      20'h80000) <=
	     20'd524352 ;
  assign NEG_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFF_ETC___d1863 =
	     NEG_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFF_ETC___d1682 +
	     20'd32 ;
  assign NEG_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFF_ETC___d1864 =
	     NEG_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFF_ETC___d1863 -
	     20'd2 ;
  assign NEG_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFF_ETC___d1866 =
	     (NEG_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFF_ETC___d1864 ^
	      20'h80000) <=
	     20'd524320 ;
  assign NEG_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFF_ETC___d1922 =
	     NEG_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFF_ETC___d1863 -
	     20'd1 ;
  assign NEG_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFF_ETC___d1924 =
	     (NEG_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFF_ETC___d1922 ^
	      20'h80000) <=
	     20'd524320 ;
  assign NEG_SEXT_requestR_BITS_190_TO_180_599_MINUS_10_ETC___d2613 =
	     -{ {13{requestR_BITS_190_TO_180_599_MINUS_1023___d2611[10]}},
		requestR_BITS_190_TO_180_599_MINUS_1023___d2611 } ;
  assign NEG_SEXT_requestR_BITS_190_TO_180_599_MINUS_10_ETC___d2645 =
	     NEG_SEXT_requestR_BITS_190_TO_180_599_MINUS_10_ETC___d2613 +
	     24'd32 ;
  assign NEG_SEXT_requestR_BITS_190_TO_180_599_MINUS_10_ETC___d2646 =
	     NEG_SEXT_requestR_BITS_190_TO_180_599_MINUS_10_ETC___d2645 -
	     24'd2 ;
  assign NEG_SEXT_requestR_BITS_190_TO_180_599_MINUS_10_ETC___d2648 =
	     (NEG_SEXT_requestR_BITS_190_TO_180_599_MINUS_10_ETC___d2646 ^
	      24'h800000) <=
	     24'd8388640 ;
  assign NEG_SEXT_requestR_BITS_190_TO_180_599_MINUS_10_ETC___d2710 =
	     NEG_SEXT_requestR_BITS_190_TO_180_599_MINUS_10_ETC___d2645 -
	     24'd1 ;
  assign NEG_SEXT_requestR_BITS_190_TO_180_599_MINUS_10_ETC___d2712 =
	     (NEG_SEXT_requestR_BITS_190_TO_180_599_MINUS_10_ETC___d2710 ^
	      24'h800000) <=
	     24'd8388640 ;
  assign NEG_SEXT_requestR_BITS_190_TO_180_599_MINUS_10_ETC___d3134 =
	     NEG_SEXT_requestR_BITS_190_TO_180_599_MINUS_10_ETC___d2613 +
	     24'd64 ;
  assign NEG_SEXT_requestR_BITS_190_TO_180_599_MINUS_10_ETC___d3135 =
	     NEG_SEXT_requestR_BITS_190_TO_180_599_MINUS_10_ETC___d3134 -
	     24'd2 ;
  assign NEG_SEXT_requestR_BITS_190_TO_180_599_MINUS_10_ETC___d3137 =
	     (NEG_SEXT_requestR_BITS_190_TO_180_599_MINUS_10_ETC___d3135 ^
	      24'h800000) <=
	     24'd8388672 ;
  assign NEG_SEXT_requestR_BITS_190_TO_180_599_MINUS_10_ETC___d3192 =
	     NEG_SEXT_requestR_BITS_190_TO_180_599_MINUS_10_ETC___d3134 -
	     24'd1 ;
  assign NEG_SEXT_requestR_BITS_190_TO_180_599_MINUS_10_ETC___d3194 =
	     (NEG_SEXT_requestR_BITS_190_TO_180_599_MINUS_10_ETC___d3192 ^
	      24'h800000) <=
	     24'd8388672 ;
  assign NOT_3074_MINUS_0_CONCAT_IF_requestR_BIT_179_71_ETC___d4331 =
	     !_3074_MINUS_0_CONCAT_IF_requestR_BIT_179_71_THE_ETC___d3304 ||
	     (_3074_MINUS_0_CONCAT_IF_requestR_BIT_179_71_THE_ETC___d3305 ?
		_0_CONCAT_IF_IF_0b0_CONCAT_NOT_requestR_BITS_19_ETC___d4279[2] :
		_0_CONCAT_IF_requestR_BITS_190_TO_180_599_EQ_0__ETC___d4291[2]) ;
  assign NOT_3074_MINUS_0_CONCAT_IF_requestR_BIT_179_71_ETC___d4359 =
	     !_3074_MINUS_0_CONCAT_IF_requestR_BIT_179_71_THE_ETC___d3304 ||
	     (_3074_MINUS_0_CONCAT_IF_requestR_BIT_179_71_THE_ETC___d3305 ?
		_0_CONCAT_IF_IF_0b0_CONCAT_NOT_requestR_BITS_19_ETC___d4279[0] :
		_0_CONCAT_IF_requestR_BITS_190_TO_180_599_EQ_0__ETC___d4291[0]) ;
  assign NOT_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFF_ETC___d1758 =
	     (value_BIT_23___h161776 || sV1_sfd__h824 != 23'd0) &&
	     ((NEG_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFF_ETC___d1682 ==
	       20'd1048513) ?
		_theResult_____2__h36734[64:63] != 2'b11 :
		NEG_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFF_ETC___d1715[19] ||
		NEG_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFF_ETC___d1717 &&
		IF_requestR_BITS_194_TO_192_0_EQ_0x0_1_OR_NOT__ETC___d1738 &&
		x__h37699[88:25] == 64'h7FFFFFFFFFFFFFFF) ;
  assign NOT_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFF_ETC___d1821 =
	     (value_BIT_23___h161776 || sV1_sfd__h824 != 23'd0) &&
	     !NEG_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFF_ETC___d1778[19] &&
	     (!NEG_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFF_ETC___d1780 ||
	      guard__h38794 != 2'd0) ;
  assign NOT_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFF_ETC___d1905 =
	     (value_BIT_23___h161776 || sV1_sfd__h824 != 23'd0) &&
	     ((NEG_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFF_ETC___d1682 ==
	       20'd1048545) ?
		_theResult_____2__h39517[32:31] != 2'b11 :
		NEG_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFF_ETC___d1864[19] ||
		NEG_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFF_ETC___d1866 &&
		IF_requestR_BITS_194_TO_192_0_EQ_0x0_1_OR_NOT__ETC___d1887 &&
		x__h40258[56:25] == 32'h7FFFFFFF) ;
  assign NOT_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFF_ETC___d1966 =
	     (value_BIT_23___h161776 || sV1_sfd__h824 != 23'd0) &&
	     !NEG_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFF_ETC___d1922[19] &&
	     (!NEG_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFF_ETC___d1924 ||
	      guard__h41115 != 2'd0) ;
  assign NOT_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFF_ETC___d2032 =
	     (value_BIT_23___h161776 || sV1_sfd__h824 != 23'd0 ||
	      sV2_exp__h926 != 8'd0 ||
	      sV2_sfd__h927 != 23'd0) &&
	     requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5_AND_ETC___d2031 ;
  assign NOT_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFF_ETC___d2033 =
	     (sV1_exp__h823 != 8'd255 || sV1_sfd__h824 == 23'd0) &&
	     (sV2_exp__h926 != 8'd255 || sV2_sfd__h927 == 23'd0) &&
	     NOT_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFF_ETC___d2032 ;
  assign NOT_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFF_ETC___d2090 =
	     !IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d2018 &&
	     (!IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d2019 ||
	      !IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d2020) &&
	     IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d2023 &&
	     (!IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d2019 ||
	      IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d2025) ;
  assign NOT_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFF_ETC___d2096 =
	     (sV1_exp__h823 != 8'd255 || sV1_sfd__h824 == 23'd0) &&
	     (sV2_exp__h926 != 8'd255 || sV2_sfd__h927 == 23'd0) &&
	     IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d2095 ;
  assign NOT_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFF_ETC___d2114 =
	     (sV1_exp__h823 != 8'd255 || sV1_sfd__h824 == 23'd0) &&
	     (sV2_exp__h926 != 8'd255 || sV2_sfd__h927 == 23'd0) &&
	     (requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5_AND_ETC___d2031 ||
	      IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d2095) ;
  assign NOT_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFF_ETC___d4468 =
	     !sV1_sfd__h824[21] && !sV1_sfd__h824[20] && !sV1_sfd__h824[19] &&
	     !sV1_sfd__h824[18] &&
	     !sV1_sfd__h824[17] &&
	     !sV1_sfd__h824[16] &&
	     !sV1_sfd__h824[15] &&
	     !sV1_sfd__h824[14] &&
	     !sV1_sfd__h824[13] &&
	     !sV1_sfd__h824[12] &&
	     !sV1_sfd__h824[11] &&
	     !sV1_sfd__h824[10] &&
	     !sV1_sfd__h824[9] &&
	     !sV1_sfd__h824[8] &&
	     !sV1_sfd__h824[7] &&
	     !sV1_sfd__h824[6] &&
	     !sV1_sfd__h824[5] &&
	     !sV1_sfd__h824[4] &&
	     !sV1_sfd__h824[3] &&
	     !sV1_sfd__h824[2] &&
	     !sV1_sfd__h824[1] &&
	     !sV1_sfd__h824[0] ;
  assign NOT_IF_requestR_BIT_159_6_THEN_NEG_requestR_BI_ETC___d1260 =
	     !sfd__h23980[31] && !sfd__h23980[30] && !sfd__h23980[29] &&
	     !sfd__h23980[28] &&
	     !sfd__h23980[27] &&
	     !sfd__h23980[26] &&
	     !sfd__h23980[25] &&
	     !sfd__h23980[24] &&
	     !sfd__h23980[23] &&
	     !sfd__h23980[22] &&
	     !sfd__h23980[21] &&
	     !sfd__h23980[20] &&
	     !sfd__h23980[19] &&
	     !sfd__h23980[18] &&
	     !sfd__h23980[17] &&
	     !sfd__h23980[16] &&
	     !sfd__h23980[15] &&
	     !sfd__h23980[14] &&
	     !sfd__h23980[13] &&
	     !sfd__h23980[12] &&
	     !sfd__h23980[11] &&
	     !sfd__h23980[10] &&
	     !sfd__h23980[9] &&
	     !sfd__h23980[8] &&
	     !sfd__h23980[7] &&
	     !sfd__h23980[6] &&
	     !sfd__h23980[5] &&
	     !sfd__h23980[4] &&
	     !sfd__h23980[3] &&
	     !sfd__h23980[2] &&
	     !sfd__h23980[1] &&
	     !sfd__h23980[0] ||
	     !_32_MINUS_0_CONCAT_IF_IF_requestR_BIT_159_6_THE_ETC___d1256 ||
	     _32_MINUS_0_CONCAT_IF_IF_requestR_BIT_159_6_THE_ETC___d1258 ;
  assign NOT_IF_requestR_BIT_191_27_THEN_NEG_requestR_B_ETC___d2774 =
	     !sfd__h2230[63] && !sfd__h2230[62] && !sfd__h2230[61] &&
	     !sfd__h2230[60] &&
	     !sfd__h2230[59] &&
	     !sfd__h2230[58] &&
	     !sfd__h2230[57] &&
	     !sfd__h2230[56] &&
	     !sfd__h2230[55] &&
	     !sfd__h2230[54] &&
	     !sfd__h2230[53] &&
	     !sfd__h2230[52] &&
	     !sfd__h2230[51] &&
	     !sfd__h2230[50] &&
	     !sfd__h2230[49] &&
	     !sfd__h2230[48] &&
	     !sfd__h2230[47] &&
	     !sfd__h2230[46] &&
	     !sfd__h2230[45] &&
	     !sfd__h2230[44] &&
	     !sfd__h2230[43] &&
	     !sfd__h2230[42] &&
	     !sfd__h2230[41] &&
	     !sfd__h2230[40] &&
	     !sfd__h2230[39] &&
	     !sfd__h2230[38] &&
	     !sfd__h2230[37] &&
	     !sfd__h2230[36] &&
	     !sfd__h2230[35] &&
	     !sfd__h2230[34] &&
	     !sfd__h2230[33] &&
	     !sfd__h2230[32] &&
	     !sfd__h2230[31] &&
	     !sfd__h2230[30] &&
	     !sfd__h2230[29] &&
	     !sfd__h2230[28] &&
	     !sfd__h2230[27] &&
	     !sfd__h2230[26] &&
	     !sfd__h2230[25] &&
	     !sfd__h2230[24] &&
	     !sfd__h2230[23] &&
	     !sfd__h2230[22] &&
	     !sfd__h2230[21] &&
	     !sfd__h2230[20] &&
	     !sfd__h2230[19] &&
	     !sfd__h2230[18] &&
	     !sfd__h2230[17] &&
	     !sfd__h2230[16] &&
	     !sfd__h2230[15] &&
	     !sfd__h2230[14] &&
	     !sfd__h2230[13] &&
	     !sfd__h2230[12] &&
	     !sfd__h2230[11] &&
	     !sfd__h2230[10] &&
	     !sfd__h2230[9] &&
	     !sfd__h2230[8] &&
	     !sfd__h2230[7] &&
	     !sfd__h2230[6] &&
	     !sfd__h2230[5] &&
	     !sfd__h2230[4] &&
	     !sfd__h2230[3] &&
	     !sfd__h2230[2] &&
	     !sfd__h2230[1] &&
	     !sfd__h2230[0] ||
	     !_64_MINUS_0_CONCAT_IF_IF_requestR_BIT_191_27_TH_ETC___d2770 ||
	     _64_MINUS_0_CONCAT_IF_IF_requestR_BIT_191_27_TH_ETC___d2772 ;
  assign NOT_IF_requestR_BIT_191_27_THEN_NEG_requestR_B_ETC___d392 =
	     !sfd__h2230[63] && !sfd__h2230[62] && !sfd__h2230[61] &&
	     !sfd__h2230[60] &&
	     !sfd__h2230[59] &&
	     !sfd__h2230[58] &&
	     !sfd__h2230[57] &&
	     !sfd__h2230[56] &&
	     !sfd__h2230[55] &&
	     !sfd__h2230[54] &&
	     !sfd__h2230[53] &&
	     !sfd__h2230[52] &&
	     !sfd__h2230[51] &&
	     !sfd__h2230[50] &&
	     !sfd__h2230[49] &&
	     !sfd__h2230[48] &&
	     !sfd__h2230[47] &&
	     !sfd__h2230[46] &&
	     !sfd__h2230[45] &&
	     !sfd__h2230[44] &&
	     !sfd__h2230[43] &&
	     !sfd__h2230[42] &&
	     !sfd__h2230[41] &&
	     !sfd__h2230[40] &&
	     !sfd__h2230[39] &&
	     !sfd__h2230[38] &&
	     !sfd__h2230[37] &&
	     !sfd__h2230[36] &&
	     !sfd__h2230[35] &&
	     !sfd__h2230[34] &&
	     !sfd__h2230[33] &&
	     !sfd__h2230[32] &&
	     !sfd__h2230[31] &&
	     !sfd__h2230[30] &&
	     !sfd__h2230[29] &&
	     !sfd__h2230[28] &&
	     !sfd__h2230[27] &&
	     !sfd__h2230[26] &&
	     !sfd__h2230[25] &&
	     !sfd__h2230[24] &&
	     !sfd__h2230[23] &&
	     !sfd__h2230[22] &&
	     !sfd__h2230[21] &&
	     !sfd__h2230[20] &&
	     !sfd__h2230[19] &&
	     !sfd__h2230[18] &&
	     !sfd__h2230[17] &&
	     !sfd__h2230[16] &&
	     !sfd__h2230[15] &&
	     !sfd__h2230[14] &&
	     !sfd__h2230[13] &&
	     !sfd__h2230[12] &&
	     !sfd__h2230[11] &&
	     !sfd__h2230[10] &&
	     !sfd__h2230[9] &&
	     !sfd__h2230[8] &&
	     !sfd__h2230[7] &&
	     !sfd__h2230[6] &&
	     !sfd__h2230[5] &&
	     !sfd__h2230[4] &&
	     !sfd__h2230[3] &&
	     !sfd__h2230[2] &&
	     !sfd__h2230[1] &&
	     !sfd__h2230[0] ||
	     !_64_MINUS_0_CONCAT_IF_IF_requestR_BIT_191_27_TH_ETC___d388 ||
	     _64_MINUS_0_CONCAT_IF_IF_requestR_BIT_191_27_TH_ETC___d390 ;
  assign NOT_requestR_BITS_159_TO_128_121_EQ_0_122_123__ETC___d1643 =
	     requestR[159:128] != 32'd0 &&
	     (requestR[159] ||
	      requestR_BIT_158_12_OR_requestR_BIT_157_14_OR__ETC___d1058) &&
	     (!_32_MINUS_0_CONCAT_IF_requestR_BIT_159_6_THEN_0_ETC___d1511 ||
	      !_32_MINUS_0_CONCAT_IF_requestR_BIT_159_6_THEN_0_ETC___d1512 &&
	      !_32_MINUS_0_CONCAT_IF_requestR_BIT_159_6_THEN_0_ETC___d1513 &&
	      _theResult___fst_exp__h36129 == 8'd255 &&
	      _theResult___fst_sfd__h36130 == 23'd0) ;
  assign NOT_requestR_BITS_190_TO_180_599_EQ_0_609_615__ETC___d2690 =
	     (requestR[190:180] != 11'd0 || requestR[179:128] != 52'd0) &&
	     ((NEG_SEXT_requestR_BITS_190_TO_180_599_MINUS_10_ETC___d2613 ==
	       24'd16777185) ?
		_theResult_____2__h72057[32:31] != 2'b11 :
		NEG_SEXT_requestR_BITS_190_TO_180_599_MINUS_10_ETC___d2646[23] ||
		NEG_SEXT_requestR_BITS_190_TO_180_599_MINUS_10_ETC___d2648 &&
		IF_requestR_BITS_194_TO_192_0_EQ_0x0_1_OR_NOT__ETC___d2669 &&
		x__h72798[85:54] == 32'h7FFFFFFF) ;
  assign NOT_requestR_BITS_190_TO_180_599_EQ_0_609_615__ETC___d2754 =
	     (requestR[190:180] != 11'd0 || requestR[179:128] != 52'd0) &&
	     !NEG_SEXT_requestR_BITS_190_TO_180_599_MINUS_10_ETC___d2710[23] &&
	     (!NEG_SEXT_requestR_BITS_190_TO_180_599_MINUS_10_ETC___d2712 ||
	      guard__h73655 != 2'd0) ;
  assign NOT_requestR_BITS_190_TO_180_599_EQ_0_609_615__ETC___d3175 =
	     (requestR[190:180] != 11'd0 || requestR[179:128] != 52'd0) &&
	     ((NEG_SEXT_requestR_BITS_190_TO_180_599_MINUS_10_ETC___d2613 ==
	       24'd16777153) ?
		_theResult_____2__h96911[64:63] != 2'b11 :
		NEG_SEXT_requestR_BITS_190_TO_180_599_MINUS_10_ETC___d3135[23] ||
		NEG_SEXT_requestR_BITS_190_TO_180_599_MINUS_10_ETC___d3137 &&
		IF_requestR_BITS_194_TO_192_0_EQ_0x0_1_OR_NOT__ETC___d3158 &&
		x__h97876[117:54] == 64'h7FFFFFFFFFFFFFFF) ;
  assign NOT_requestR_BITS_190_TO_180_599_EQ_0_609_615__ETC___d3235 =
	     (requestR[190:180] != 11'd0 || requestR[179:128] != 52'd0) &&
	     !NEG_SEXT_requestR_BITS_190_TO_180_599_MINUS_10_ETC___d3192[23] &&
	     (!NEG_SEXT_requestR_BITS_190_TO_180_599_MINUS_10_ETC___d3194 ||
	      guard__h98954 != 2'd0) ;
  assign NOT_requestR_BITS_190_TO_180_599_EQ_2047_600_6_ETC___d5211 =
	     (requestR[190:180] != 11'd2047 || requestR[179:128] == 52'd0) &&
	     (requestR[126:116] != 11'd2047 || requestR[115:64] == 52'd0) &&
	     (requestR[190:180] != 11'd0 || requestR[179:128] != 52'd0 ||
	      requestR[126:116] != 11'd0 ||
	      requestR[115:64] != 52'd0) &&
	     (requestR[191] && !requestR[127] ||
	      (requestR[191] || !requestR[127]) &&
	      IF_requestR_BIT_191_27_THEN_NOT_requestR_BITS__ETC___d5207) ;
  assign NOT_requestR_BITS_190_TO_180_599_EQ_2047_600_6_ETC___d5276 =
	     (requestR[190:180] != 11'd2047 || requestR[179:128] == 52'd0) &&
	     (requestR[126:116] != 11'd2047 || requestR[115:64] == 52'd0) &&
	     (requestR[191] && !requestR[127] ||
	      (requestR[191] || !requestR[127]) &&
	      IF_requestR_BIT_191_27_THEN_NOT_requestR_BITS__ETC___d5207 ||
	      requestR_BITS_190_TO_180_599_EQ_0_609_AND_requ_ETC___d5257) ;
  assign NOT_requestR_BITS_190_TO_180_599_ULT_requestR__ETC___d5253 =
	     !requestR_BITS_190_TO_180_599_ULT_requestR_BITS_ETC___d5203 &&
	     (!requestR_BITS_190_TO_180_599_EQ_requestR_BITS__ETC___d5198 ||
	      !requestR_BITS_179_TO_128_601_ULT_requestR_BITS_ETC___d5204) &&
	     requestR_BITS_190_TO_180_599_ULE_requestR_BITS_ETC___d5196 &&
	     (!requestR_BITS_190_TO_180_599_EQ_requestR_BITS__ETC___d5198 ||
	      requestR_BITS_179_TO_128_601_ULE_requestR_BITS_ETC___d5199) ;
  assign NOT_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5_ETC___d2094 =
	     (requestR[191:160] != 32'hFFFFFFFF || !requestR[159] ||
	      requestR[127:96] == 32'hFFFFFFFF && requestR[95]) &&
	     (requestR[191:160] == 32'hFFFFFFFF && requestR[159] ||
	      requestR[127:96] != 32'hFFFFFFFF ||
	      !requestR[95]) &&
	     ((requestR[191:160] != 32'hFFFFFFFF || !requestR[159]) ?
		NOT_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFF_ETC___d2090 :
		IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d2091) ;
  assign NOT_requestR_BIT_158_12_13_AND_NOT_requestR_BI_ETC___d803 =
	     !requestR[158] && !requestR[157] && !requestR[156] &&
	     !requestR[155] &&
	     !requestR[154] &&
	     !requestR[153] &&
	     !requestR[152] &&
	     !requestR[151] &&
	     !requestR[150] &&
	     !requestR[149] &&
	     !requestR[148] &&
	     !requestR[147] &&
	     !requestR[146] &&
	     !requestR[145] &&
	     !requestR[144] &&
	     !requestR[143] &&
	     !requestR[142] &&
	     !requestR[141] &&
	     !requestR[140] &&
	     !requestR[139] &&
	     !requestR[138] &&
	     !requestR[137] &&
	     !requestR[136] &&
	     !requestR[135] &&
	     !requestR[134] &&
	     !requestR[133] &&
	     !requestR[132] &&
	     !requestR[131] &&
	     !requestR[130] &&
	     !requestR[129] &&
	     !requestR[128] ;
  assign NOT_requestR_BIT_179_71_72_AND_NOT_requestR_BI_ETC___d824 =
	     !requestR[179] && !requestR[178] && !requestR[177] &&
	     !requestR[176] &&
	     !requestR[175] &&
	     !requestR[174] &&
	     !requestR[173] &&
	     !requestR[172] &&
	     !requestR[171] &&
	     !requestR[170] &&
	     !requestR[169] &&
	     !requestR[168] &&
	     !requestR[167] &&
	     !requestR[166] &&
	     !requestR[165] &&
	     !requestR[164] &&
	     !requestR[163] &&
	     !requestR[162] &&
	     !requestR[161] &&
	     !requestR[160] &&
	     !requestR[159] &&
	     NOT_requestR_BIT_158_12_13_AND_NOT_requestR_BI_ETC___d803 ;
  assign NOT_requestR_BIT_191_27_48_AND_NOT_requestR_BI_ETC___d3042 =
	     !requestR[191] && !requestR[190] && !requestR[189] &&
	     !requestR[188] &&
	     !requestR[187] &&
	     !requestR[186] &&
	     !requestR[185] &&
	     !requestR[184] &&
	     !requestR[183] &&
	     !requestR[182] &&
	     !requestR[181] &&
	     !requestR[180] &&
	     NOT_requestR_BIT_179_71_72_AND_NOT_requestR_BI_ETC___d824 ||
	     !_64_MINUS_0_CONCAT_IF_requestR_BIT_191_27_THEN__ETC___d2955 ||
	     _64_MINUS_0_CONCAT_IF_requestR_BIT_191_27_THEN__ETC___d2956 ;
  assign NOT_requestR_BIT_191_27_48_AND_NOT_requestR_BI_ETC___d994 =
	     !requestR[191] && !requestR[190] && !requestR[189] &&
	     !requestR[188] &&
	     !requestR[187] &&
	     !requestR[186] &&
	     !requestR[185] &&
	     !requestR[184] &&
	     !requestR[183] &&
	     !requestR[182] &&
	     !requestR[181] &&
	     !requestR[180] &&
	     NOT_requestR_BIT_179_71_72_AND_NOT_requestR_BI_ETC___d824 ||
	     !_64_MINUS_0_CONCAT_IF_requestR_BIT_191_27_THEN__ETC___d905 ||
	     _64_MINUS_0_CONCAT_IF_requestR_BIT_191_27_THEN__ETC___d906 ;
  assign SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFF_ETC___d4566 =
	     { {4{IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d1680[7]}},
	       IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d1680 } ;
  assign SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFF_ETC___d4567 =
	     (SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFF_ETC___d4566 ^
	      12'h800) <=
	     12'd3071 ;
  assign SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFF_ETC___d4568 =
	     (SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFF_ETC___d4566 ^
	      12'h800) <
	     12'd1026 ;
  assign SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFF_ETC__q150 =
	     SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFF_ETC___d4566 +
	     12'd1023 ;
  assign SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFF_ETC__q153 =
	     SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFF_ETC__q150[10:0] -
	     11'd1023 ;
  assign SEXT_requestR_BITS_190_TO_180_599_MINUS_1023_611___d3734 =
	     { requestR_BITS_190_TO_180_599_MINUS_1023___d2611[10],
	       requestR_BITS_190_TO_180_599_MINUS_1023___d2611 } ;
  assign SEXT_requestR_BITS_190_TO_180_599_MINUS_1023_6_ETC___d3735 =
	     (SEXT_requestR_BITS_190_TO_180_599_MINUS_1023_611___d3734 ^
	      12'h800) <=
	     12'd2175 ;
  assign SEXT_requestR_BITS_190_TO_180_599_MINUS_1023_6_ETC___d3736 =
	     (SEXT_requestR_BITS_190_TO_180_599_MINUS_1023_611___d3734 ^
	      12'h800) <
	     12'd1922 ;
  assign SEXT_requestR_BITS_190_TO_180_599_MINUS_1023_6_ETC__q118 =
	     SEXT_requestR_BITS_190_TO_180_599_MINUS_1023_611___d3734 +
	     12'd127 ;
  assign SEXT_requestR_BITS_190_TO_180_599_MINUS_1023_6_ETC__q121 =
	     SEXT_requestR_BITS_190_TO_180_599_MINUS_1023_6_ETC__q118[7:0] -
	     8'd127 ;
  assign _0_CONCAT_IF_IF_0b0_CONCAT_NOT_requestR_BITS_19_ETC___d3539 =
	     ({ 3'd0,
		IF_IF_0b0_CONCAT_NOT_requestR_BITS_190_TO_180__ETC___d3537 } ^
	      9'h100) <=
	     9'd256 ;
  assign _0_CONCAT_IF_IF_0b0_CONCAT_NOT_requestR_BITS_19_ETC___d4279 =
	     { 3'd0,
	       _theResult___fst_exp__h119464 == 8'd0 &&
	       (sfdin__h119458[56:34] == 23'd0 || guard__h111367 != 2'b0),
	       1'd0 } |
	     { 2'd0,
	       _theResult___fst_exp__h120091 == 8'd255 &&
	       _theResult___fst_sfd__h120092 == 23'd0,
	       1'd0,
	       _theResult___fst_exp__h119464 != 8'd255 &&
	       guard__h111367 != 2'b0 } ;
  assign _0_CONCAT_IF_IF_3074_MINUS_SEXT_IF_requestR_BIT_ETC___d4817 =
	     ({ 6'd0,
		IF_IF_3074_MINUS_SEXT_IF_requestR_BITS_191_TO__ETC___d4815 } ^
	      12'h800) <=
	     12'd2048 ;
  assign _0_CONCAT_IF_IF_3074_MINUS_SEXT_IF_requestR_BIT_ETC___d5102 =
	     { 3'd0,
	       _theResult___fst_exp__h178652 == 11'd0 &&
	       (sfdin__h178646[56:5] == 52'd0 || guard__h170426 != 2'b0),
	       1'd0 } |
	     { 2'd0,
	       _theResult___fst_exp__h179482 == 11'd2047 &&
	       _theResult___fst_sfd__h179483 == 52'd0,
	       1'd0,
	       _theResult___fst_exp__h178652 != 11'd2047 &&
	       guard__h170426 != 2'b0 } ;
  assign _0_CONCAT_IF_IF_3970_MINUS_SEXT_requestR_BITS_1_ETC___d3983 =
	     ({ 3'd0,
		IF_IF_3970_MINUS_SEXT_requestR_BITS_190_TO_180_ETC___d3981 } ^
	      9'h100) <=
	     9'd256 ;
  assign _0_CONCAT_IF_IF_3970_MINUS_SEXT_requestR_BITS_1_ETC___d4308 =
	     { 3'd0,
	       _theResult___fst_exp__h137317 == 8'd0 &&
	       (sfdin__h137311[56:34] == 23'd0 || guard__h129091 != 2'b0),
	       1'd0 } |
	     { 2'd0,
	       _theResult___fst_exp__h137944 == 8'd255 &&
	       _theResult___fst_sfd__h137945 == 23'd0,
	       1'd0,
	       _theResult___fst_exp__h137317 != 8'd255 &&
	       guard__h129091 != 2'b0 } ;
  assign _0_CONCAT_IF_IF_requestR_BITS_191_TO_160_4_EQ_0_ETC___d4497 =
	     ({ 6'd0,
		IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_ETC___d4495 } ^
	      12'h800) <=
	     12'd2944 ;
  assign _0_CONCAT_IF_IF_requestR_BITS_191_TO_160_4_EQ_0_ETC___d4890 =
	     ({ 6'd0,
		IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_ETC___d4495 } ^
	      12'h800) <=
	     (IF_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFFF_ETC___d4889 ^
	      12'h800) ;
  assign _0_CONCAT_IF_IF_requestR_BITS_191_TO_160_4_EQ_0_ETC___d5085 =
	     { 3'd0,
	       _theResult___fst_exp__h169079 == 11'd0 &&
	       guard__h161118 != 2'b0,
	       1'd0 } |
	     { 2'd0,
	       _theResult___fst_exp__h169835 == 11'd2047 &&
	       _theResult___fst_sfd__h169836 == 52'd0,
	       1'd0,
	       _theResult___fst_exp__h169079 != 11'd2047 &&
	       guard__h161118 != 2'b0 } ;
  assign _0_CONCAT_IF_requestR_BITS_190_TO_180_599_EQ_0__ETC___d3661 =
	     ({ 3'd0,
		IF_requestR_BITS_190_TO_180_599_EQ_0_609_THEN__ETC___d3659 } ^
	      9'h100) <=
	     9'd384 ;
  assign _0_CONCAT_IF_requestR_BITS_190_TO_180_599_EQ_0__ETC___d4056 =
	     ({ 3'd0,
		IF_requestR_BITS_190_TO_180_599_EQ_0_609_THEN__ETC___d3659 } ^
	      9'h100) <=
	     (IF_SEXT_requestR_BITS_190_TO_180_599_MINUS_102_ETC___d4055 ^
	      9'h100) ;
  assign _0_CONCAT_IF_requestR_BITS_190_TO_180_599_EQ_0__ETC___d4291 =
	     { 3'd0,
	       _theResult___fst_exp__h128150 == 8'd0 &&
	       guard__h120102 != 2'b0,
	       1'd0 } |
	     { 2'd0,
	       _theResult___fst_exp__h128703 == 8'd255 &&
	       _theResult___fst_sfd__h128704 == 23'd0,
	       1'd0,
	       _theResult___fst_exp__h128150 != 8'd255 &&
	       guard__h120102 != 2'b0 } ;
  assign _0b0_CONCAT_NOT_IF_requestR_BITS_191_TO_160_4_E_ETC___d4573 =
	     b__h39582 >>
	     _3074_MINUS_SEXT_IF_requestR_BITS_191_TO_160_4__ETC___d4569 ;
  assign _0b0_CONCAT_NOT_requestR_BITS_190_TO_180_599_EQ_ETC___d3741 =
	     sfd__h103727 >>
	     _3970_MINUS_SEXT_requestR_BITS_190_TO_180_599_M_ETC___d3737 ;
  assign _1_CONCAT_DONTCARE_CONCAT_requestR_BITS_63_TO_3_ETC___d68 =
	     { 33'h1AAAAAAAA,
	       requestR[63:32] == 32'hFFFFFFFF && requestR[31],
	       (requestR[63:32] == 32'hFFFFFFFF) ?
		 requestR[30:0] :
		 31'h7FC00000 } ;
  assign _3074_MINUS_0_CONCAT_IF_requestR_BIT_179_71_THE_ETC___d3303 =
	     12'd3074 -
	     { 6'd0,
	       requestR[179] ?
		 6'd0 :
		 (requestR[178] ?
		    6'd1 :
		    (requestR[177] ?
		       6'd2 :
		       (requestR[176] ?
			  6'd3 :
			  (requestR[175] ?
			     6'd4 :
			     (requestR[174] ?
				6'd5 :
				(requestR[173] ?
				   6'd6 :
				   (requestR[172] ?
				      6'd7 :
				      (requestR[171] ?
					 6'd8 :
					 (requestR[170] ?
					    6'd9 :
					    (requestR[169] ?
					       6'd10 :
					       (requestR[168] ?
						  6'd11 :
						  (requestR[167] ?
						     6'd12 :
						     (requestR[166] ?
							6'd13 :
							(requestR[165] ?
							   6'd14 :
							   (requestR[164] ?
							      6'd15 :
							      (requestR[163] ?
								 6'd16 :
								 (requestR[162] ?
								    6'd17 :
								    (requestR[161] ?
								       6'd18 :
								       (requestR[160] ?
									  6'd19 :
									  (requestR[159] ?
									     6'd20 :
									     (requestR[158] ?
										6'd21 :
										(requestR[157] ?
										   6'd22 :
										   (requestR[156] ?
										      6'd23 :
										      (requestR[155] ?
											 6'd24 :
											 (requestR[154] ?
											    6'd25 :
											    (requestR[153] ?
											       6'd26 :
											       (requestR[152] ?
												  6'd27 :
												  (requestR[151] ?
												     6'd28 :
												     (requestR[150] ?
													6'd29 :
													(requestR[149] ?
													   6'd30 :
													   (requestR[148] ?
													      6'd31 :
													      (requestR[147] ?
														 6'd32 :
														 (requestR[146] ?
														    6'd33 :
														    (requestR[145] ?
														       6'd34 :
														       (requestR[144] ?
															  6'd35 :
															  (requestR[143] ?
															     6'd36 :
															     (requestR[142] ?
																6'd37 :
																(requestR[141] ?
																   6'd38 :
																   (requestR[140] ?
																      6'd39 :
																      (requestR[139] ?
																	 6'd40 :
																	 (requestR[138] ?
																	    6'd41 :
																	    (requestR[137] ?
																	       6'd42 :
																	       (requestR[136] ?
																		  6'd43 :
																		  (requestR[135] ?
																		     6'd44 :
																		     (requestR[134] ?
																			6'd45 :
																			(requestR[133] ?
																			   6'd46 :
																			   (requestR[132] ?
																			      6'd47 :
																			      (requestR[131] ?
																				 6'd48 :
																				 (requestR[130] ?
																				    6'd49 :
																				    (requestR[129] ?
																				       6'd50 :
																				       (requestR[128] ?
																					  6'd51 :
																					  6'd52))))))))))))))))))))))))))))))))))))))))))))))))))) } ;
  assign _3074_MINUS_0_CONCAT_IF_requestR_BIT_179_71_THE_ETC___d3304 =
	     (_3074_MINUS_0_CONCAT_IF_requestR_BIT_179_71_THE_ETC___d3303 ^
	      12'h800) <=
	     12'd2175 ;
  assign _3074_MINUS_0_CONCAT_IF_requestR_BIT_179_71_THE_ETC___d3305 =
	     (_3074_MINUS_0_CONCAT_IF_requestR_BIT_179_71_THE_ETC___d3303 ^
	      12'h800) <
	     12'd1922 ;
  assign _3074_MINUS_0_CONCAT_IF_requestR_BIT_179_71_THE_ETC___d4294 =
	     _3074_MINUS_0_CONCAT_IF_requestR_BIT_179_71_THE_ETC___d3304 &&
	     (_3074_MINUS_0_CONCAT_IF_requestR_BIT_179_71_THE_ETC___d3305 ?
		_0_CONCAT_IF_IF_0b0_CONCAT_NOT_requestR_BITS_19_ETC___d4279[4] :
		_0_CONCAT_IF_requestR_BITS_190_TO_180_599_EQ_0__ETC___d4291[4]) ;
  assign _3074_MINUS_0_CONCAT_IF_requestR_BIT_179_71_THE_ETC___d4319 =
	     _3074_MINUS_0_CONCAT_IF_requestR_BIT_179_71_THE_ETC___d3304 &&
	     (_3074_MINUS_0_CONCAT_IF_requestR_BIT_179_71_THE_ETC___d3305 ?
		_0_CONCAT_IF_IF_0b0_CONCAT_NOT_requestR_BITS_19_ETC___d4279[3] :
		_0_CONCAT_IF_requestR_BITS_190_TO_180_599_EQ_0__ETC___d4291[3]) ;
  assign _3074_MINUS_0_CONCAT_IF_requestR_BIT_179_71_THE_ETC___d4346 =
	     _3074_MINUS_0_CONCAT_IF_requestR_BIT_179_71_THE_ETC___d3304 &&
	     (_3074_MINUS_0_CONCAT_IF_requestR_BIT_179_71_THE_ETC___d3305 ?
		_0_CONCAT_IF_IF_0b0_CONCAT_NOT_requestR_BITS_19_ETC___d4279[1] :
		_0_CONCAT_IF_requestR_BITS_190_TO_180_599_EQ_0__ETC___d4291[1]) ;
  assign _3074_MINUS_SEXT_IF_requestR_BITS_191_TO_160_4__ETC___d4569 =
	     12'd3074 -
	     SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFF_ETC___d4566 ;
  assign _32_MINUS_0_CONCAT_IF_IF_requestR_BIT_159_6_THE_ETC___d1255 =
	     (9'd32 -
	      { 3'd0,
		IF_IF_requestR_BIT_159_6_THEN_NEG_requestR_BIT_ETC___d1252 }) -
	     9'd1 ;
  assign _32_MINUS_0_CONCAT_IF_IF_requestR_BIT_159_6_THE_ETC___d1256 =
	     (_32_MINUS_0_CONCAT_IF_IF_requestR_BIT_159_6_THE_ETC___d1255 ^
	      9'h100) <=
	     9'd383 ;
  assign _32_MINUS_0_CONCAT_IF_IF_requestR_BIT_159_6_THE_ETC___d1258 =
	     (_32_MINUS_0_CONCAT_IF_IF_requestR_BIT_159_6_THE_ETC___d1255 ^
	      9'h100) <
	     9'd107 ;
  assign _32_MINUS_0_CONCAT_IF_IF_requestR_BIT_159_6_THE_ETC___d1261 =
	     (_32_MINUS_0_CONCAT_IF_IF_requestR_BIT_159_6_THE_ETC___d1255 ^
	      9'h100) <
	     9'd130 ;
  assign _32_MINUS_0_CONCAT_IF_IF_requestR_BIT_159_6_THE_ETC___d2233 =
	     (12'd32 -
	      { 6'd0,
		IF_IF_requestR_BIT_159_6_THEN_NEG_requestR_BIT_ETC___d2230 }) -
	     12'd1 ;
  assign _32_MINUS_0_CONCAT_IF_IF_requestR_BIT_159_6_THE_ETC___d2234 =
	     (_32_MINUS_0_CONCAT_IF_IF_requestR_BIT_159_6_THE_ETC___d2233 ^
	      12'h800) <=
	     12'd3071 ;
  assign _32_MINUS_0_CONCAT_IF_IF_requestR_BIT_159_6_THE_ETC___d2236 =
	     (_32_MINUS_0_CONCAT_IF_IF_requestR_BIT_159_6_THE_ETC___d2233 ^
	      12'h800) <
	     12'd974 ;
  assign _32_MINUS_0_CONCAT_IF_IF_requestR_BIT_159_6_THE_ETC___d2238 =
	     (_32_MINUS_0_CONCAT_IF_IF_requestR_BIT_159_6_THE_ETC___d2233 ^
	      12'h800) <
	     12'd1026 ;
  assign _32_MINUS_0_CONCAT_IF_requestR_BIT_159_6_THEN_0_ETC___d1510 =
	     (9'd32 -
	      { 3'd0,
		IF_requestR_BIT_159_6_THEN_0_ELSE_IF_requestR__ETC___d1507 }) -
	     9'd1 ;
  assign _32_MINUS_0_CONCAT_IF_requestR_BIT_159_6_THEN_0_ETC___d1511 =
	     (_32_MINUS_0_CONCAT_IF_requestR_BIT_159_6_THEN_0_ETC___d1510 ^
	      9'h100) <=
	     9'd383 ;
  assign _32_MINUS_0_CONCAT_IF_requestR_BIT_159_6_THEN_0_ETC___d1512 =
	     (_32_MINUS_0_CONCAT_IF_requestR_BIT_159_6_THEN_0_ETC___d1510 ^
	      9'h100) <
	     9'd107 ;
  assign _32_MINUS_0_CONCAT_IF_requestR_BIT_159_6_THEN_0_ETC___d1513 =
	     (_32_MINUS_0_CONCAT_IF_requestR_BIT_159_6_THEN_0_ETC___d1510 ^
	      9'h100) <
	     9'd130 ;
  assign _32_MINUS_0_CONCAT_IF_requestR_BIT_159_6_THEN_0_ETC___d2448 =
	     (12'd32 -
	      { 6'd0,
		IF_requestR_BIT_159_6_THEN_0_ELSE_IF_requestR__ETC___d2445 }) -
	     12'd1 ;
  assign _32_MINUS_0_CONCAT_IF_requestR_BIT_159_6_THEN_0_ETC___d2449 =
	     (_32_MINUS_0_CONCAT_IF_requestR_BIT_159_6_THEN_0_ETC___d2448 ^
	      12'h800) <=
	     12'd3071 ;
  assign _32_MINUS_0_CONCAT_IF_requestR_BIT_159_6_THEN_0_ETC___d2450 =
	     (_32_MINUS_0_CONCAT_IF_requestR_BIT_159_6_THEN_0_ETC___d2448 ^
	      12'h800) <
	     12'd974 ;
  assign _32_MINUS_0_CONCAT_IF_requestR_BIT_159_6_THEN_0_ETC___d2451 =
	     (_32_MINUS_0_CONCAT_IF_requestR_BIT_159_6_THEN_0_ETC___d2448 ^
	      12'h800) <
	     12'd1026 ;
  assign _3970_MINUS_0_CONCAT_IF_IF_requestR_BITS_191_TO_ETC___d4423 =
	     12'd3970 -
	     { 7'd0,
	       sV1_sfd__h824[22] ?
		 5'd0 :
		 (sV1_sfd__h824[21] ?
		    5'd1 :
		    (sV1_sfd__h824[20] ?
		       5'd2 :
		       (sV1_sfd__h824[19] ?
			  5'd3 :
			  (sV1_sfd__h824[18] ?
			     5'd4 :
			     (sV1_sfd__h824[17] ?
				5'd5 :
				(sV1_sfd__h824[16] ?
				   5'd6 :
				   (sV1_sfd__h824[15] ?
				      5'd7 :
				      (sV1_sfd__h824[14] ?
					 5'd8 :
					 (sV1_sfd__h824[13] ?
					    5'd9 :
					    (sV1_sfd__h824[12] ?
					       5'd10 :
					       (sV1_sfd__h824[11] ?
						  5'd11 :
						  (sV1_sfd__h824[10] ?
						     5'd12 :
						     (sV1_sfd__h824[9] ?
							5'd13 :
							(sV1_sfd__h824[8] ?
							   5'd14 :
							   (sV1_sfd__h824[7] ?
							      5'd15 :
							      (sV1_sfd__h824[6] ?
								 5'd16 :
								 (sV1_sfd__h824[5] ?
								    5'd17 :
								    (sV1_sfd__h824[4] ?
								       5'd18 :
								       (sV1_sfd__h824[3] ?
									  5'd19 :
									  (sV1_sfd__h824[2] ?
									     5'd20 :
									     (sV1_sfd__h824[1] ?
										5'd21 :
										(sV1_sfd__h824[0] ?
										   5'd22 :
										   5'd23)))))))))))))))))))))) } ;
  assign _3970_MINUS_0_CONCAT_IF_IF_requestR_BITS_191_TO_ETC___d4424 =
	     (_3970_MINUS_0_CONCAT_IF_IF_requestR_BITS_191_TO_ETC___d4423 ^
	      12'h800) <=
	     12'd3071 ;
  assign _3970_MINUS_0_CONCAT_IF_IF_requestR_BITS_191_TO_ETC___d4425 =
	     (_3970_MINUS_0_CONCAT_IF_IF_requestR_BITS_191_TO_ETC___d4423 ^
	      12'h800) <
	     12'd1026 ;
  assign _3970_MINUS_SEXT_requestR_BITS_190_TO_180_599_M_ETC___d3737 =
	     12'd3970 -
	     SEXT_requestR_BITS_190_TO_180_599_MINUS_1023_611___d3734 ;
  assign _64_MINUS_0_CONCAT_IF_IF_requestR_BIT_191_27_TH_ETC___d2769 =
	     (12'd64 -
	      { 5'd0,
		IF_IF_requestR_BIT_191_27_THEN_NEG_requestR_BI_ETC___d384 }) -
	     12'd1 ;
  assign _64_MINUS_0_CONCAT_IF_IF_requestR_BIT_191_27_TH_ETC___d2770 =
	     (_64_MINUS_0_CONCAT_IF_IF_requestR_BIT_191_27_TH_ETC___d2769 ^
	      12'h800) <=
	     12'd3071 ;
  assign _64_MINUS_0_CONCAT_IF_IF_requestR_BIT_191_27_TH_ETC___d2772 =
	     (_64_MINUS_0_CONCAT_IF_IF_requestR_BIT_191_27_TH_ETC___d2769 ^
	      12'h800) <
	     12'd974 ;
  assign _64_MINUS_0_CONCAT_IF_IF_requestR_BIT_191_27_TH_ETC___d2775 =
	     (_64_MINUS_0_CONCAT_IF_IF_requestR_BIT_191_27_TH_ETC___d2769 ^
	      12'h800) <
	     12'd1026 ;
  assign _64_MINUS_0_CONCAT_IF_IF_requestR_BIT_191_27_TH_ETC___d387 =
	     (9'd64 -
	      { 2'd0,
		IF_IF_requestR_BIT_191_27_THEN_NEG_requestR_BI_ETC___d384 }) -
	     9'd1 ;
  assign _64_MINUS_0_CONCAT_IF_IF_requestR_BIT_191_27_TH_ETC___d388 =
	     (_64_MINUS_0_CONCAT_IF_IF_requestR_BIT_191_27_TH_ETC___d387 ^
	      9'h100) <=
	     9'd383 ;
  assign _64_MINUS_0_CONCAT_IF_IF_requestR_BIT_191_27_TH_ETC___d390 =
	     (_64_MINUS_0_CONCAT_IF_IF_requestR_BIT_191_27_TH_ETC___d387 ^
	      9'h100) <
	     9'd107 ;
  assign _64_MINUS_0_CONCAT_IF_IF_requestR_BIT_191_27_TH_ETC___d393 =
	     (_64_MINUS_0_CONCAT_IF_IF_requestR_BIT_191_27_TH_ETC___d387 ^
	      9'h100) <
	     9'd130 ;
  assign _64_MINUS_0_CONCAT_IF_requestR_BIT_191_27_THEN__ETC___d2954 =
	     (12'd64 -
	      { 5'd0,
		IF_requestR_BIT_191_27_THEN_0_ELSE_IF_requestR_ETC___d901 }) -
	     12'd1 ;
  assign _64_MINUS_0_CONCAT_IF_requestR_BIT_191_27_THEN__ETC___d2955 =
	     (_64_MINUS_0_CONCAT_IF_requestR_BIT_191_27_THEN__ETC___d2954 ^
	      12'h800) <=
	     12'd3071 ;
  assign _64_MINUS_0_CONCAT_IF_requestR_BIT_191_27_THEN__ETC___d2956 =
	     (_64_MINUS_0_CONCAT_IF_requestR_BIT_191_27_THEN__ETC___d2954 ^
	      12'h800) <
	     12'd974 ;
  assign _64_MINUS_0_CONCAT_IF_requestR_BIT_191_27_THEN__ETC___d2957 =
	     (_64_MINUS_0_CONCAT_IF_requestR_BIT_191_27_THEN__ETC___d2954 ^
	      12'h800) <
	     12'd1026 ;
  assign _64_MINUS_0_CONCAT_IF_requestR_BIT_191_27_THEN__ETC___d904 =
	     (9'd64 -
	      { 2'd0,
		IF_requestR_BIT_191_27_THEN_0_ELSE_IF_requestR_ETC___d901 }) -
	     9'd1 ;
  assign _64_MINUS_0_CONCAT_IF_requestR_BIT_191_27_THEN__ETC___d905 =
	     (_64_MINUS_0_CONCAT_IF_requestR_BIT_191_27_THEN__ETC___d904 ^
	      9'h100) <=
	     9'd383 ;
  assign _64_MINUS_0_CONCAT_IF_requestR_BIT_191_27_THEN__ETC___d906 =
	     (_64_MINUS_0_CONCAT_IF_requestR_BIT_191_27_THEN__ETC___d904 ^
	      9'h100) <
	     9'd107 ;
  assign _64_MINUS_0_CONCAT_IF_requestR_BIT_191_27_THEN__ETC___d907 =
	     (_64_MINUS_0_CONCAT_IF_requestR_BIT_191_27_THEN__ETC___d904 ^
	      9'h100) <
	     9'd130 ;
  assign _theResult_____2__h36734 =
	     IF_requestR_BITS_194_TO_192_0_EQ_0x0_1_OR_NOT__ETC___d1706 ?
	       out1___1__h37450 :
	       IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d1689[88:24] ;
  assign _theResult_____2__h39517 =
	     IF_requestR_BITS_194_TO_192_0_EQ_0x0_1_OR_NOT__ETC___d1855 ?
	       out1___1__h40009 :
	       IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d1838[56:24] ;
  assign _theResult_____2__h72057 =
	     IF_requestR_BITS_194_TO_192_0_EQ_0x0_1_OR_NOT__ETC___d2637 ?
	       out1___1__h72549 :
	       IF_requestR_BIT_191_27_THEN_NEG_0b0_CONCAT_NOT_ETC___d2620[85:53] ;
  assign _theResult_____2__h96911 =
	     IF_requestR_BITS_194_TO_192_0_EQ_0x0_1_OR_NOT__ETC___d3126 ?
	       out1___1__h97627 :
	       IF_requestR_BIT_191_27_THEN_NEG_0b0_CONCAT_NOT_ETC___d3109[117:53] ;
  assign _theResult____h111357 =
	     (value__h72124 == 54'd0) ? sfd__h103727 : 57'd1 ;
  assign _theResult____h129081 =
	     ((_3970_MINUS_SEXT_requestR_BITS_190_TO_180_599_M_ETC___d3737 ^
	       12'h800) <
	      12'd2105) ?
	       result__h129694 :
	       _theResult____h111357 ;
  assign _theResult____h170416 =
	     ((_3074_MINUS_SEXT_IF_requestR_BITS_191_TO_160_4__ETC___d4569 ^
	       12'h800) <
	      12'd2105) ?
	       result__h171029 :
	       ((value__h36801 == 25'd0) ? b__h39582 : 57'd1) ;
  assign _theResult___exp__h119990 =
	     sfd__h119556[24] ?
	       ((_theResult___fst_exp__h119464 == 8'd254) ?
		  8'd255 :
		  din_inc___2_exp__h146641) :
	       ((_theResult___fst_exp__h119464 == 8'd0 &&
		 sfd__h119556[24:23] == 2'b01) ?
		  8'd1 :
		  _theResult___fst_exp__h119464) ;
  assign _theResult___exp__h12261 =
	     (sfd__h11862[24] || sfd__h11862[24:23] == 2'b01) ? 8'd1 : 8'd0 ;
  assign _theResult___exp__h12814 =
	     sfd__h12405[24] ?
	       ((x__h12390[7:0] == 8'd254) ?
		  8'd255 :
		  din_inc___2_exp__h12957) :
	       ((x__h12390[7:0] == 8'd0 && sfd__h12405[24:23] == 2'b01) ?
		  8'd1 :
		  x__h12390[7:0]) ;
  assign _theResult___exp__h128602 =
	     sfd__h128168[24] ?
	       ((_theResult___fst_exp__h128150 == 8'd254) ?
		  8'd255 :
		  din_inc___2_exp__h146665) :
	       ((_theResult___fst_exp__h128150 == 8'd0 &&
		 sfd__h128168[24:23] == 2'b01) ?
		  8'd1 :
		  _theResult___fst_exp__h128150) ;
  assign _theResult___exp__h137843 =
	     sfd__h137409[24] ?
	       ((_theResult___fst_exp__h137317 == 8'd254) ?
		  8'd255 :
		  din_inc___2_exp__h146695) :
	       ((_theResult___fst_exp__h137317 == 8'd0 &&
		 sfd__h137409[24:23] == 2'b01) ?
		  8'd1 :
		  _theResult___fst_exp__h137317) ;
  assign _theResult___exp__h146509 =
	     sfd__h146051[24] ?
	       ((_theResult___fst_exp__h146032 == 8'd254) ?
		  8'd255 :
		  din_inc___2_exp__h146719) :
	       ((_theResult___fst_exp__h146032 == 8'd0 &&
		 sfd__h146051[24:23] == 2'b01) ?
		  8'd1 :
		  _theResult___fst_exp__h146032) ;
  assign _theResult___exp__h169734 =
	     sfd__h169097[53] ?
	       ((_theResult___fst_exp__h169079 == 11'd2046) ?
		  11'd2047 :
		  din_inc___2_exp__h188299) :
	       ((_theResult___fst_exp__h169079 == 11'd0 &&
		 sfd__h169097[53:52] == 2'b01) ?
		  11'd1 :
		  _theResult___fst_exp__h169079) ;
  assign _theResult___exp__h179381 =
	     sfd__h178744[53] ?
	       ((_theResult___fst_exp__h178652 == 11'd2046) ?
		  11'd2047 :
		  din_inc___2_exp__h188329) :
	       ((_theResult___fst_exp__h178652 == 11'd0 &&
		 sfd__h178744[53:52] == 2'b01) ?
		  11'd1 :
		  _theResult___fst_exp__h178652) ;
  assign _theResult___exp__h188163 =
	     sfd__h187502[53] ?
	       ((_theResult___fst_exp__h187483 == 11'd2046) ?
		  11'd2047 :
		  din_inc___2_exp__h188353) :
	       ((_theResult___fst_exp__h187483 == 11'd0 &&
		 sfd__h187502[53:52] == 2'b01) ?
		  11'd1 :
		  _theResult___fst_exp__h187483) ;
  assign _theResult___exp__h22880 =
	     (sfd__h22484[24] || sfd__h22484[24:23] == 2'b01) ? 8'd1 : 8'd0 ;
  assign _theResult___exp__h23432 =
	     sfd__h23023[24] ?
	       ((x__h23008[7:0] == 8'd254) ?
		  8'd255 :
		  din_inc___2_exp__h23570) :
	       ((x__h23008[7:0] == 8'd0 && sfd__h23023[24:23] == 2'b01) ?
		  8'd1 :
		  x__h23008[7:0]) ;
  assign _theResult___exp__h29307 =
	     (sfd__h28911[24] || sfd__h28911[24:23] == 2'b01) ? 8'd1 : 8'd0 ;
  assign _theResult___exp__h29860 =
	     sfd__h29451[24] ?
	       ((x__h29436[7:0] == 8'd254) ?
		  8'd255 :
		  din_inc___2_exp__h30003) :
	       ((x__h29436[7:0] == 8'd0 && sfd__h29451[24:23] == 2'b01) ?
		  8'd1 :
		  x__h29436[7:0]) ;
  assign _theResult___exp__h35478 =
	     (sfd__h35082[24] || sfd__h35082[24:23] == 2'b01) ? 8'd1 : 8'd0 ;
  assign _theResult___exp__h36030 =
	     sfd__h35621[24] ?
	       ((x__h35606[7:0] == 8'd254) ?
		  8'd255 :
		  din_inc___2_exp__h36168) :
	       ((x__h35606[7:0] == 8'd0 && sfd__h35621[24:23] == 2'b01) ?
		  8'd1 :
		  x__h35606[7:0]) ;
  assign _theResult___exp__h60903 =
	     (sfd__h60304[53] || sfd__h60304[53:52] == 2'b01) ?
	       11'd1 :
	       11'd0 ;
  assign _theResult___exp__h61659 =
	     sfd__h61047[53] ?
	       ((x__h61032[10:0] == 11'd2046) ?
		  11'd2047 :
		  din_inc___2_exp__h61802) :
	       ((x__h61032[10:0] == 11'd0 && sfd__h61047[53:52] == 2'b01) ?
		  11'd1 :
		  x__h61032[10:0]) ;
  assign _theResult___exp__h70599 =
	     (sfd__h70000[53] || sfd__h70000[53:52] == 2'b01) ?
	       11'd1 :
	       11'd0 ;
  assign _theResult___exp__h71354 =
	     sfd__h70742[53] ?
	       ((x__h70727[10:0] == 11'd2046) ?
		  11'd2047 :
		  din_inc___2_exp__h71492) :
	       ((x__h70727[10:0] == 11'd0 && sfd__h70742[53:52] == 2'b01) ?
		  11'd1 :
		  x__h70727[10:0]) ;
  assign _theResult___exp__h84444 =
	     (sfd__h83845[53] || sfd__h83845[53:52] == 2'b01) ?
	       11'd1 :
	       11'd0 ;
  assign _theResult___exp__h85200 =
	     sfd__h84588[53] ?
	       ((x__h84573[10:0] == 11'd2046) ?
		  11'd2047 :
		  din_inc___2_exp__h85343) :
	       ((x__h84573[10:0] == 11'd0 && sfd__h84588[53:52] == 2'b01) ?
		  11'd1 :
		  x__h84573[10:0]) ;
  assign _theResult___exp__h95456 =
	     (sfd__h94857[53] || sfd__h94857[53:52] == 2'b01) ?
	       11'd1 :
	       11'd0 ;
  assign _theResult___exp__h96211 =
	     sfd__h95599[53] ?
	       ((x__h95584[10:0] == 11'd2046) ?
		  11'd2047 :
		  din_inc___2_exp__h96349) :
	       ((x__h95584[10:0] == 11'd0 && sfd__h95599[53:52] == 2'b01) ?
		  11'd1 :
		  x__h95584[10:0]) ;
  assign _theResult___fst_exp__h111339 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3) ?
	       8'd255 :
	       CASE_requestR_BITS_194_TO_192_0x1_254_0x2_IF_r_ETC__q2 ;
  assign _theResult___fst_exp__h119464 =
	     _theResult____h111357[56] ?
	       8'd2 :
	       _theResult___fst_exp__h119538 ;
  assign _theResult___fst_exp__h119529 =
	     8'd0 -
	     { 2'd0,
	       IF_IF_0b0_CONCAT_NOT_requestR_BITS_190_TO_180__ETC___d3537 } ;
  assign _theResult___fst_exp__h119535 =
	     (!_theResult____h111357[56] && !_theResult____h111357[55] &&
	      !_theResult____h111357[54] &&
	      !_theResult____h111357[53] &&
	      !_theResult____h111357[52] &&
	      !_theResult____h111357[51] &&
	      !_theResult____h111357[50] &&
	      !_theResult____h111357[49] &&
	      !_theResult____h111357[48] &&
	      !_theResult____h111357[47] &&
	      !_theResult____h111357[46] &&
	      !_theResult____h111357[45] &&
	      !_theResult____h111357[44] &&
	      !_theResult____h111357[43] &&
	      !_theResult____h111357[42] &&
	      !_theResult____h111357[41] &&
	      !_theResult____h111357[40] &&
	      !_theResult____h111357[39] &&
	      !_theResult____h111357[38] &&
	      !_theResult____h111357[37] &&
	      !_theResult____h111357[36] &&
	      !_theResult____h111357[35] &&
	      !_theResult____h111357[34] &&
	      !_theResult____h111357[33] &&
	      !_theResult____h111357[32] &&
	      !_theResult____h111357[31] &&
	      !_theResult____h111357[30] &&
	      !_theResult____h111357[29] &&
	      !_theResult____h111357[28] &&
	      !_theResult____h111357[27] &&
	      !_theResult____h111357[26] &&
	      !_theResult____h111357[25] &&
	      !_theResult____h111357[24] &&
	      !_theResult____h111357[23] &&
	      !_theResult____h111357[22] &&
	      !_theResult____h111357[21] &&
	      !_theResult____h111357[20] &&
	      !_theResult____h111357[19] &&
	      !_theResult____h111357[18] &&
	      !_theResult____h111357[17] &&
	      !_theResult____h111357[16] &&
	      !_theResult____h111357[15] &&
	      !_theResult____h111357[14] &&
	      !_theResult____h111357[13] &&
	      !_theResult____h111357[12] &&
	      !_theResult____h111357[11] &&
	      !_theResult____h111357[10] &&
	      !_theResult____h111357[9] &&
	      !_theResult____h111357[8] &&
	      !_theResult____h111357[7] &&
	      !_theResult____h111357[6] &&
	      !_theResult____h111357[5] &&
	      !_theResult____h111357[4] &&
	      !_theResult____h111357[3] &&
	      !_theResult____h111357[2] &&
	      !_theResult____h111357[1] &&
	      !_theResult____h111357[0] ||
	      !_0_CONCAT_IF_IF_0b0_CONCAT_NOT_requestR_BITS_19_ETC___d3539) ?
	       8'd0 :
	       _theResult___fst_exp__h119529 ;
  assign _theResult___fst_exp__h119538 =
	     (!_theResult____h111357[56] && _theResult____h111357[55]) ?
	       8'd1 :
	       _theResult___fst_exp__h119535 ;
  assign _theResult___fst_exp__h120088 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       CASE_guard11367_0b0_theResult___fst_exp19464_0_ETC__q125 :
	       IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d3602 ;
  assign _theResult___fst_exp__h120091 =
	     (_theResult___fst_exp__h119464 == 8'd255) ?
	       _theResult___fst_exp__h119464 :
	       _theResult___fst_exp__h120088 ;
  assign _theResult___fst_exp__h12358 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       CASE_guard1845_0b0_0_0b1_0_0b10_out_exp2264_0b_ETC__q15 :
	       IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d479 ;
  assign _theResult___fst_exp__h128141 =
	     8'd129 -
	     { 2'd0,
	       IF_requestR_BITS_190_TO_180_599_EQ_0_609_THEN__ETC___d3659 } ;
  assign _theResult___fst_exp__h128147 =
	     (requestR[190:180] == 11'd0 &&
	      NOT_requestR_BIT_179_71_72_AND_NOT_requestR_BI_ETC___d824 ||
	      !_0_CONCAT_IF_requestR_BITS_190_TO_180_599_EQ_0__ETC___d3661) ?
	       8'd0 :
	       _theResult___fst_exp__h128141 ;
  assign _theResult___fst_exp__h128150 =
	     (requestR[190:180] == 11'd0) ?
	       _theResult___fst_exp__h128147 :
	       8'd129 ;
  assign _theResult___fst_exp__h128700 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       CASE_guard20102_0b0_theResult___fst_exp28150_0_ETC__q127 :
	       IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d3719 ;
  assign _theResult___fst_exp__h128703 =
	     (_theResult___fst_exp__h128150 == 8'd255) ?
	       _theResult___fst_exp__h128150 :
	       _theResult___fst_exp__h128700 ;
  assign _theResult___fst_exp__h12911 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       CASE_guard2375_0b0_x2390_BITS_7_TO_0_0b1_x2390_ETC__q17 :
	       IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d508 ;
  assign _theResult___fst_exp__h12914 =
	     (x__h12390[7:0] == 8'd255) ?
	       x__h12390[7:0] :
	       _theResult___fst_exp__h12911 ;
  assign _theResult___fst_exp__h137317 =
	     _theResult____h129081[56] ?
	       8'd2 :
	       _theResult___fst_exp__h137391 ;
  assign _theResult___fst_exp__h137382 =
	     8'd0 -
	     { 2'd0,
	       IF_IF_3970_MINUS_SEXT_requestR_BITS_190_TO_180_ETC___d3981 } ;
  assign _theResult___fst_exp__h137388 =
	     (!_theResult____h129081[56] && !_theResult____h129081[55] &&
	      !_theResult____h129081[54] &&
	      !_theResult____h129081[53] &&
	      !_theResult____h129081[52] &&
	      !_theResult____h129081[51] &&
	      !_theResult____h129081[50] &&
	      !_theResult____h129081[49] &&
	      !_theResult____h129081[48] &&
	      !_theResult____h129081[47] &&
	      !_theResult____h129081[46] &&
	      !_theResult____h129081[45] &&
	      !_theResult____h129081[44] &&
	      !_theResult____h129081[43] &&
	      !_theResult____h129081[42] &&
	      !_theResult____h129081[41] &&
	      !_theResult____h129081[40] &&
	      !_theResult____h129081[39] &&
	      !_theResult____h129081[38] &&
	      !_theResult____h129081[37] &&
	      !_theResult____h129081[36] &&
	      !_theResult____h129081[35] &&
	      !_theResult____h129081[34] &&
	      !_theResult____h129081[33] &&
	      !_theResult____h129081[32] &&
	      !_theResult____h129081[31] &&
	      !_theResult____h129081[30] &&
	      !_theResult____h129081[29] &&
	      !_theResult____h129081[28] &&
	      !_theResult____h129081[27] &&
	      !_theResult____h129081[26] &&
	      !_theResult____h129081[25] &&
	      !_theResult____h129081[24] &&
	      !_theResult____h129081[23] &&
	      !_theResult____h129081[22] &&
	      !_theResult____h129081[21] &&
	      !_theResult____h129081[20] &&
	      !_theResult____h129081[19] &&
	      !_theResult____h129081[18] &&
	      !_theResult____h129081[17] &&
	      !_theResult____h129081[16] &&
	      !_theResult____h129081[15] &&
	      !_theResult____h129081[14] &&
	      !_theResult____h129081[13] &&
	      !_theResult____h129081[12] &&
	      !_theResult____h129081[11] &&
	      !_theResult____h129081[10] &&
	      !_theResult____h129081[9] &&
	      !_theResult____h129081[8] &&
	      !_theResult____h129081[7] &&
	      !_theResult____h129081[6] &&
	      !_theResult____h129081[5] &&
	      !_theResult____h129081[4] &&
	      !_theResult____h129081[3] &&
	      !_theResult____h129081[2] &&
	      !_theResult____h129081[1] &&
	      !_theResult____h129081[0] ||
	      !_0_CONCAT_IF_IF_3970_MINUS_SEXT_requestR_BITS_1_ETC___d3983) ?
	       8'd0 :
	       _theResult___fst_exp__h137382 ;
  assign _theResult___fst_exp__h137391 =
	     (!_theResult____h129081[56] && _theResult____h129081[55]) ?
	       8'd1 :
	       _theResult___fst_exp__h137388 ;
  assign _theResult___fst_exp__h137941 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       CASE_guard29091_0b0_theResult___fst_exp37317_0_ETC__q129 :
	       IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d4046 ;
  assign _theResult___fst_exp__h137944 =
	     (_theResult___fst_exp__h137317 == 8'd255) ?
	       _theResult___fst_exp__h137317 :
	       _theResult___fst_exp__h137941 ;
  assign _theResult___fst_exp__h145984 =
	     (SEXT_requestR_BITS_190_TO_180_599_MINUS_1023_6_ETC__q118[7:0] ==
	      8'd0) ?
	       8'd1 :
	       SEXT_requestR_BITS_190_TO_180_599_MINUS_1023_6_ETC__q118[7:0] ;
  assign _theResult___fst_exp__h146023 =
	     SEXT_requestR_BITS_190_TO_180_599_MINUS_1023_6_ETC__q118[7:0] -
	     { 2'd0,
	       IF_requestR_BITS_190_TO_180_599_EQ_0_609_THEN__ETC___d3659 } ;
  assign _theResult___fst_exp__h146029 =
	     (requestR[190:180] == 11'd0 &&
	      NOT_requestR_BIT_179_71_72_AND_NOT_requestR_BI_ETC___d824 ||
	      !_0_CONCAT_IF_requestR_BITS_190_TO_180_599_EQ_0__ETC___d4056) ?
	       8'd0 :
	       _theResult___fst_exp__h146023 ;
  assign _theResult___fst_exp__h146032 =
	     (requestR[190:180] == 11'd0) ?
	       _theResult___fst_exp__h146029 :
	       _theResult___fst_exp__h145984 ;
  assign _theResult___fst_exp__h146607 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       CASE_guard37955_0b0_theResult___fst_exp46032_0_ETC__q131 :
	       IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d4115 ;
  assign _theResult___fst_exp__h146610 =
	     (_theResult___fst_exp__h146032 == 8'd255) ?
	       _theResult___fst_exp__h146032 :
	       _theResult___fst_exp__h146607 ;
  assign _theResult___fst_exp__h146619 =
	     (requestR[190:180] == 11'd0) ?
	       (_3074_MINUS_0_CONCAT_IF_requestR_BIT_179_71_THE_ETC___d3304 ?
		  _theResult___snd_fst_exp__h128706 :
		  _theResult___fst_exp__h111339) :
	       (SEXT_requestR_BITS_190_TO_180_599_MINUS_1023_6_ETC___d3735 ?
		  _theResult___snd_fst_exp__h146613 :
		  _theResult___fst_exp__h111339) ;
  assign _theResult___fst_exp__h146622 =
	     (requestR[190:180] == 11'd0 && requestR[179:128] == 52'd0) ?
	       8'd0 :
	       _theResult___fst_exp__h146619 ;
  assign _theResult___fst_exp__h154006 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3) ?
	       11'd2047 :
	       CASE_requestR_BITS_194_TO_192_0x1_2046_0x2_IF__ETC__q4 ;
  assign _theResult___fst_exp__h169070 =
	     11'd897 -
	     { 5'd0,
	       IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_ETC___d4495 } ;
  assign _theResult___fst_exp__h169076 =
	     (sV1_exp__h823 == 8'd0 && !sV1_sfd__h824[22] &&
	      NOT_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFF_ETC___d4468 ||
	      !_0_CONCAT_IF_IF_requestR_BITS_191_TO_160_4_EQ_0_ETC___d4497) ?
	       11'd0 :
	       _theResult___fst_exp__h169070 ;
  assign _theResult___fst_exp__h169079 =
	     (sV1_exp__h823 == 8'd0) ?
	       _theResult___fst_exp__h169076 :
	       11'd897 ;
  assign _theResult___fst_exp__h169832 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       CASE_guard61118_0b0_theResult___fst_exp69079_0_ETC__q157 :
	       IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d4555 ;
  assign _theResult___fst_exp__h169835 =
	     (_theResult___fst_exp__h169079 == 11'd2047) ?
	       _theResult___fst_exp__h169079 :
	       _theResult___fst_exp__h169832 ;
  assign _theResult___fst_exp__h178652 =
	     _theResult____h170416[56] ?
	       11'd2 :
	       _theResult___fst_exp__h178726 ;
  assign _theResult___fst_exp__h178717 =
	     11'd0 -
	     { 5'd0,
	       IF_IF_3074_MINUS_SEXT_IF_requestR_BITS_191_TO__ETC___d4815 } ;
  assign _theResult___fst_exp__h178723 =
	     (!_theResult____h170416[56] && !_theResult____h170416[55] &&
	      !_theResult____h170416[54] &&
	      !_theResult____h170416[53] &&
	      !_theResult____h170416[52] &&
	      !_theResult____h170416[51] &&
	      !_theResult____h170416[50] &&
	      !_theResult____h170416[49] &&
	      !_theResult____h170416[48] &&
	      !_theResult____h170416[47] &&
	      !_theResult____h170416[46] &&
	      !_theResult____h170416[45] &&
	      !_theResult____h170416[44] &&
	      !_theResult____h170416[43] &&
	      !_theResult____h170416[42] &&
	      !_theResult____h170416[41] &&
	      !_theResult____h170416[40] &&
	      !_theResult____h170416[39] &&
	      !_theResult____h170416[38] &&
	      !_theResult____h170416[37] &&
	      !_theResult____h170416[36] &&
	      !_theResult____h170416[35] &&
	      !_theResult____h170416[34] &&
	      !_theResult____h170416[33] &&
	      !_theResult____h170416[32] &&
	      !_theResult____h170416[31] &&
	      !_theResult____h170416[30] &&
	      !_theResult____h170416[29] &&
	      !_theResult____h170416[28] &&
	      !_theResult____h170416[27] &&
	      !_theResult____h170416[26] &&
	      !_theResult____h170416[25] &&
	      !_theResult____h170416[24] &&
	      !_theResult____h170416[23] &&
	      !_theResult____h170416[22] &&
	      !_theResult____h170416[21] &&
	      !_theResult____h170416[20] &&
	      !_theResult____h170416[19] &&
	      !_theResult____h170416[18] &&
	      !_theResult____h170416[17] &&
	      !_theResult____h170416[16] &&
	      !_theResult____h170416[15] &&
	      !_theResult____h170416[14] &&
	      !_theResult____h170416[13] &&
	      !_theResult____h170416[12] &&
	      !_theResult____h170416[11] &&
	      !_theResult____h170416[10] &&
	      !_theResult____h170416[9] &&
	      !_theResult____h170416[8] &&
	      !_theResult____h170416[7] &&
	      !_theResult____h170416[6] &&
	      !_theResult____h170416[5] &&
	      !_theResult____h170416[4] &&
	      !_theResult____h170416[3] &&
	      !_theResult____h170416[2] &&
	      !_theResult____h170416[1] &&
	      !_theResult____h170416[0] ||
	      !_0_CONCAT_IF_IF_3074_MINUS_SEXT_IF_requestR_BIT_ETC___d4817) ?
	       11'd0 :
	       _theResult___fst_exp__h178717 ;
  assign _theResult___fst_exp__h178726 =
	     (!_theResult____h170416[56] && _theResult____h170416[55]) ?
	       11'd1 :
	       _theResult___fst_exp__h178723 ;
  assign _theResult___fst_exp__h179479 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       CASE_guard70426_0b0_theResult___fst_exp78652_0_ETC__q159 :
	       IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d4880 ;
  assign _theResult___fst_exp__h179482 =
	     (_theResult___fst_exp__h178652 == 11'd2047) ?
	       _theResult___fst_exp__h178652 :
	       _theResult___fst_exp__h179479 ;
  assign _theResult___fst_exp__h187435 =
	     (SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFF_ETC__q150[10:0] ==
	      11'd0) ?
	       11'd1 :
	       SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFF_ETC__q150[10:0] ;
  assign _theResult___fst_exp__h187474 =
	     SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFF_ETC__q150[10:0] -
	     { 5'd0,
	       IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_ETC___d4495 } ;
  assign _theResult___fst_exp__h187480 =
	     (sV1_exp__h823 == 8'd0 && !sV1_sfd__h824[22] &&
	      NOT_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFF_ETC___d4468 ||
	      !_0_CONCAT_IF_IF_requestR_BITS_191_TO_160_4_EQ_0_ETC___d4890) ?
	       11'd0 :
	       _theResult___fst_exp__h187474 ;
  assign _theResult___fst_exp__h187483 =
	     (sV1_exp__h823 == 8'd0) ?
	       _theResult___fst_exp__h187480 :
	       _theResult___fst_exp__h187435 ;
  assign _theResult___fst_exp__h188261 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       CASE_guard79493_0b0_theResult___fst_exp87483_0_ETC__q161 :
	       IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d4949 ;
  assign _theResult___fst_exp__h188264 =
	     (_theResult___fst_exp__h187483 == 11'd2047) ?
	       _theResult___fst_exp__h187483 :
	       _theResult___fst_exp__h188261 ;
  assign _theResult___fst_exp__h188273 =
	     (sV1_exp__h823 == 8'd0) ?
	       (_3970_MINUS_0_CONCAT_IF_IF_requestR_BITS_191_TO_ETC___d4424 ?
		  _theResult___snd_fst_exp__h169838 :
		  _theResult___fst_exp__h154006) :
	       (SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFF_ETC___d4567 ?
		  _theResult___snd_fst_exp__h188267 :
		  _theResult___fst_exp__h154006) ;
  assign _theResult___fst_exp__h188276 =
	     (sV1_exp__h823 == 8'd0 && sV1_sfd__h824 == 23'd0) ?
	       11'd0 :
	       _theResult___fst_exp__h188273 ;
  assign _theResult___fst_exp__h22976 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       CASE_guard2467_0b0_0_0b1_0_0b10_out_exp2883_0b_ETC__q26 :
	       CASE_requestR_BITS_194_TO_192_0x3_IF_guard2467_ETC__q28 ;
  assign _theResult___fst_exp__h23528 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       CASE_guard2993_0b0_x3008_BITS_7_TO_0_0b1_x3008_ETC__q33 :
	       IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d985 ;
  assign _theResult___fst_exp__h23531 =
	     (x__h23008[7:0] == 8'd255) ?
	       x__h23008[7:0] :
	       _theResult___fst_exp__h23528 ;
  assign _theResult___fst_exp__h29404 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       CASE_guard8894_0b0_0_0b1_0_0b10_out_exp9310_0b_ETC__q45 :
	       IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d1338 ;
  assign _theResult___fst_exp__h29957 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       CASE_guard9421_0b0_x9436_BITS_7_TO_0_0b1_x9436_ETC__q47 :
	       IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d1367 ;
  assign _theResult___fst_exp__h29960 =
	     (x__h29436[7:0] == 8'd255) ?
	       x__h29436[7:0] :
	       _theResult___fst_exp__h29957 ;
  assign _theResult___fst_exp__h35574 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       CASE_guard5065_0b0_0_0b1_0_0b10_out_exp5481_0b_ETC__q54 :
	       CASE_requestR_BITS_194_TO_192_0x3_IF_guard5065_ETC__q56 ;
  assign _theResult___fst_exp__h36126 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       CASE_guard5591_0b0_x5606_BITS_7_TO_0_0b1_x5606_ETC__q58 :
	       IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d1590 ;
  assign _theResult___fst_exp__h36129 =
	     (x__h35606[7:0] == 8'd255) ?
	       x__h35606[7:0] :
	       _theResult___fst_exp__h36126 ;
  assign _theResult___fst_exp__h61000 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       CASE_guard0287_0b0_0_0b1_0_0b10_out_exp0906_0b_ETC__q78 :
	       IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d2313 ;
  assign _theResult___fst_exp__h61756 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       CASE_guard1017_0b0_x1032_BITS_10_TO_0_0b1_x103_ETC__q74 :
	       IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d2342 ;
  assign _theResult___fst_exp__h61759 =
	     (x__h61032[10:0] == 11'd2047) ?
	       x__h61032[10:0] :
	       _theResult___fst_exp__h61756 ;
  assign _theResult___fst_exp__h70695 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       CASE_guard9983_0b0_0_0b1_0_0b10_out_exp0602_0b_ETC__q83 :
	       CASE_requestR_BITS_194_TO_192_0x3_IF_guard9983_ETC__q85 ;
  assign _theResult___fst_exp__h71450 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       CASE_guard0712_0b0_x0727_BITS_10_TO_0_0b1_x072_ETC__q87 :
	       IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d2529 ;
  assign _theResult___fst_exp__h71453 =
	     (x__h70727[10:0] == 11'd2047) ?
	       x__h70727[10:0] :
	       _theResult___fst_exp__h71450 ;
  assign _theResult___fst_exp__h84541 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       CASE_guard3828_0b0_0_0b1_0_0b10_out_exp4447_0b_ETC__q103 :
	       IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d2848 ;
  assign _theResult___fst_exp__h85297 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       CASE_guard4558_0b0_x4573_BITS_10_TO_0_0b1_x457_ETC__q99 :
	       IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d2877 ;
  assign _theResult___fst_exp__h85300 =
	     (x__h84573[10:0] == 11'd2047) ?
	       x__h84573[10:0] :
	       _theResult___fst_exp__h85297 ;
  assign _theResult___fst_exp__h95552 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       CASE_guard4840_0b0_0_0b1_0_0b10_out_exp5459_0b_ETC__q29 :
	       CASE_requestR_BITS_194_TO_192_0x3_IF_guard4840_ETC__q31 ;
  assign _theResult___fst_exp__h96307 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       CASE_guard5569_0b0_x5584_BITS_10_TO_0_0b1_x558_ETC__q107 :
	       IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d3033 ;
  assign _theResult___fst_exp__h96310 =
	     (x__h95584[10:0] == 11'd2047) ?
	       x__h95584[10:0] :
	       _theResult___fst_exp__h96307 ;
  assign _theResult___fst_sfd__h100023 = { 1'd1, requestR[178:128] } ;
  assign _theResult___fst_sfd__h111340 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3) ?
	       23'd0 :
	       CASE_requestR_BITS_194_TO_192_0x1_8388607_0x2__ETC__q3 ;
  assign _theResult___fst_sfd__h120089 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       CASE_guard11367_0b0_sfdin19458_BITS_56_TO_34_0_ETC__q135 :
	       IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d4149 ;
  assign _theResult___fst_sfd__h120092 =
	     (_theResult___fst_exp__h119464 == 8'd255) ?
	       sfdin__h119458[56:34] :
	       _theResult___fst_sfd__h120089 ;
  assign _theResult___fst_sfd__h12359 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       CASE_guard1845_0b0_sfd___31835_BITS_63_TO_41_0_ETC__q19 :
	       IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d531 ;
  assign _theResult___fst_sfd__h128701 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       CASE_guard20102_0b0_theResult___snd28101_BITS__ETC__q133 :
	       IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d4168 ;
  assign _theResult___fst_sfd__h128704 =
	     (_theResult___fst_exp__h128150 == 8'd255) ?
	       _theResult___snd__h128101[56:34] :
	       _theResult___fst_sfd__h128701 ;
  assign _theResult___fst_sfd__h12912 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       CASE_guard2375_0b0_sfd___31835_BITS_62_TO_40_0_ETC__q21 :
	       IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d549 ;
  assign _theResult___fst_sfd__h12915 =
	     (x__h12390[7:0] == 8'd255) ?
	       sfd___3__h11835[62:40] :
	       _theResult___fst_sfd__h12912 ;
  assign _theResult___fst_sfd__h137942 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       CASE_guard29091_0b0_sfdin37311_BITS_56_TO_34_0_ETC__q137 :
	       IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d4195 ;
  assign _theResult___fst_sfd__h137945 =
	     (_theResult___fst_exp__h137317 == 8'd255) ?
	       sfdin__h137311[56:34] :
	       _theResult___fst_sfd__h137942 ;
  assign _theResult___fst_sfd__h146608 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       CASE_guard37955_0b0_theResult___snd45978_BITS__ETC__q139 :
	       IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d4214 ;
  assign _theResult___fst_sfd__h146611 =
	     (_theResult___fst_exp__h146032 == 8'd255) ?
	       _theResult___snd__h145978[56:34] :
	       _theResult___fst_sfd__h146608 ;
  assign _theResult___fst_sfd__h146620 =
	     (requestR[190:180] == 11'd0) ?
	       (_3074_MINUS_0_CONCAT_IF_requestR_BIT_179_71_THE_ETC___d3304 ?
		  _theResult___snd_fst_sfd__h128707 :
		  _theResult___fst_sfd__h111340) :
	       (SEXT_requestR_BITS_190_TO_180_599_MINUS_1023_6_ETC___d3735 ?
		  _theResult___snd_fst_sfd__h146614 :
		  _theResult___fst_sfd__h111340) ;
  assign _theResult___fst_sfd__h146626 =
	     ((requestR[190:180] == 11'd2047 || requestR[190:180] == 11'd0) &&
	      requestR[179:128] == 52'd0) ?
	       23'd0 :
	       _theResult___fst_sfd__h146620 ;
  assign _theResult___fst_sfd__h148525 = { 1'd1, sV1_sfd__h824[21:0] } ;
  assign _theResult___fst_sfd__h154007 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3) ?
	       52'd0 :
	       CASE_requestR_BITS_194_TO_192_0x1_450359962737_ETC__q5 ;
  assign _theResult___fst_sfd__h169833 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       CASE_guard61118_0b0_theResult___snd69030_BITS__ETC__q169 :
	       IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d4982 ;
  assign _theResult___fst_sfd__h169836 =
	     (_theResult___fst_exp__h169079 == 11'd2047) ?
	       _theResult___snd__h169030[56:5] :
	       _theResult___fst_sfd__h169833 ;
  assign _theResult___fst_sfd__h179480 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       CASE_guard70426_0b0_sfdin78646_BITS_56_TO_5_0b_ETC__q171 :
	       IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d5009 ;
  assign _theResult___fst_sfd__h179483 =
	     (_theResult___fst_exp__h178652 == 11'd2047) ?
	       sfdin__h178646[56:5] :
	       _theResult___fst_sfd__h179480 ;
  assign _theResult___fst_sfd__h188262 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       CASE_guard79493_0b0_theResult___snd87429_BITS__ETC__q173 :
	       IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d5028 ;
  assign _theResult___fst_sfd__h188265 =
	     (_theResult___fst_exp__h187483 == 11'd2047) ?
	       _theResult___snd__h187429[56:5] :
	       _theResult___fst_sfd__h188262 ;
  assign _theResult___fst_sfd__h188274 =
	     (sV1_exp__h823 == 8'd0) ?
	       (_3970_MINUS_0_CONCAT_IF_IF_requestR_BITS_191_TO_ETC___d4424 ?
		  _theResult___snd_fst_sfd__h169839 :
		  _theResult___fst_sfd__h154007) :
	       (SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFF_ETC___d4567 ?
		  _theResult___snd_fst_sfd__h188268 :
		  _theResult___fst_sfd__h154007) ;
  assign _theResult___fst_sfd__h188280 =
	     ((sV1_exp__h823 == 8'd255 || sV1_exp__h823 == 8'd0) &&
	      sV1_sfd__h824 == 23'd0) ?
	       52'd0 :
	       _theResult___fst_sfd__h188274 ;
  assign _theResult___fst_sfd__h22977 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       CASE_guard2467_0b0_sfd___32457_BITS_63_TO_41_0_ETC__q37 :
	       IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d1008 ;
  assign _theResult___fst_sfd__h23529 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       CASE_guard2993_0b0_sfd___32457_BITS_62_TO_40_0_ETC__q35 :
	       IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d1023 ;
  assign _theResult___fst_sfd__h23532 =
	     (x__h23008[7:0] == 8'd255) ?
	       sfd___3__h22457[62:40] :
	       _theResult___fst_sfd__h23529 ;
  assign _theResult___fst_sfd__h29405 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       CASE_guard8894_0b0_sfd___38884_BITS_31_TO_9_0b_ETC__q49 :
	       IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d1390 ;
  assign _theResult___fst_sfd__h29958 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       CASE_guard9421_0b0_sfd___38884_BITS_30_TO_8_0b_ETC__q51 :
	       IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d1408 ;
  assign _theResult___fst_sfd__h29961 =
	     (x__h29436[7:0] == 8'd255) ?
	       sfd___3__h28884[30:8] :
	       _theResult___fst_sfd__h29958 ;
  assign _theResult___fst_sfd__h35575 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       CASE_guard5065_0b0_sfd___35055_BITS_31_TO_9_0b_ETC__q62 :
	       IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d1613 ;
  assign _theResult___fst_sfd__h36127 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       CASE_guard5591_0b0_sfd___35055_BITS_30_TO_8_0b_ETC__q60 :
	       IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d1628 ;
  assign _theResult___fst_sfd__h36130 =
	     (x__h35606[7:0] == 8'd255) ?
	       sfd___3__h35055[30:8] :
	       _theResult___fst_sfd__h36127 ;
  assign _theResult___fst_sfd__h61001 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       CASE_guard0287_0b0_sfd___30277_BITS_54_TO_3_0b_ETC__q80 :
	       IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d2365 ;
  assign _theResult___fst_sfd__h61757 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       CASE_guard1017_0b0_sfd___30277_BITS_53_TO_2_0b_ETC__q76 :
	       IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d2383 ;
  assign _theResult___fst_sfd__h61760 =
	     (x__h61032[10:0] == 11'd2047) ?
	       sfd___3__h60277[53:2] :
	       _theResult___fst_sfd__h61757 ;
  assign _theResult___fst_sfd__h70696 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       CASE_guard9983_0b0_sfd___39973_BITS_54_TO_3_0b_ETC__q91 :
	       IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d2551 ;
  assign _theResult___fst_sfd__h71451 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       CASE_guard0712_0b0_sfd___39973_BITS_53_TO_2_0b_ETC__q89 :
	       IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d2566 ;
  assign _theResult___fst_sfd__h71454 =
	     (x__h70727[10:0] == 11'd2047) ?
	       sfd___3__h69973[53:2] :
	       _theResult___fst_sfd__h71451 ;
  assign _theResult___fst_sfd__h84542 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       CASE_guard3828_0b0_sfd___31835_BITS_63_TO_12_0_ETC__q105 :
	       IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d2900 ;
  assign _theResult___fst_sfd__h85298 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       CASE_guard4558_0b0_sfd___31835_BITS_62_TO_11_0_ETC__q101 :
	       IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d2918 ;
  assign _theResult___fst_sfd__h85301 =
	     (x__h84573[10:0] == 11'd2047) ?
	       sfd___3__h11835[62:11] :
	       _theResult___fst_sfd__h85298 ;
  assign _theResult___fst_sfd__h95553 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       CASE_guard4840_0b0_sfd___32457_BITS_63_TO_12_0_ETC__q111 :
	       IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d3056 ;
  assign _theResult___fst_sfd__h96308 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       CASE_guard5569_0b0_sfd___32457_BITS_62_TO_11_0_ETC__q109 :
	       IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d3071 ;
  assign _theResult___fst_sfd__h96311 =
	     (x__h95584[10:0] == 11'd2047) ?
	       sfd___3__h22457[62:11] :
	       _theResult___fst_sfd__h96308 ;
  assign _theResult___sfd__h119991 =
	     sfd__h119556[24] ?
	       ((_theResult___fst_exp__h119464 == 8'd254) ?
		  23'd0 :
		  sfd__h119556[23:1]) :
	       sfd__h119556[22:0] ;
  assign _theResult___sfd__h12262 =
	     sfd__h11862[24] ? sfd__h11862[23:1] : sfd__h11862[22:0] ;
  assign _theResult___sfd__h12815 =
	     sfd__h12405[24] ?
	       ((x__h12390[7:0] == 8'd254) ? 23'd0 : sfd__h12405[23:1]) :
	       sfd__h12405[22:0] ;
  assign _theResult___sfd__h128603 =
	     sfd__h128168[24] ?
	       ((_theResult___fst_exp__h128150 == 8'd254) ?
		  23'd0 :
		  sfd__h128168[23:1]) :
	       sfd__h128168[22:0] ;
  assign _theResult___sfd__h137844 =
	     sfd__h137409[24] ?
	       ((_theResult___fst_exp__h137317 == 8'd254) ?
		  23'd0 :
		  sfd__h137409[23:1]) :
	       sfd__h137409[22:0] ;
  assign _theResult___sfd__h146510 =
	     sfd__h146051[24] ?
	       ((_theResult___fst_exp__h146032 == 8'd254) ?
		  23'd0 :
		  sfd__h146051[23:1]) :
	       sfd__h146051[22:0] ;
  assign _theResult___sfd__h169735 =
	     sfd__h169097[53] ?
	       ((_theResult___fst_exp__h169079 == 11'd2046) ?
		  52'd0 :
		  sfd__h169097[52:1]) :
	       sfd__h169097[51:0] ;
  assign _theResult___sfd__h179382 =
	     sfd__h178744[53] ?
	       ((_theResult___fst_exp__h178652 == 11'd2046) ?
		  52'd0 :
		  sfd__h178744[52:1]) :
	       sfd__h178744[51:0] ;
  assign _theResult___sfd__h188164 =
	     sfd__h187502[53] ?
	       ((_theResult___fst_exp__h187483 == 11'd2046) ?
		  52'd0 :
		  sfd__h187502[52:1]) :
	       sfd__h187502[51:0] ;
  assign _theResult___sfd__h22881 =
	     sfd__h22484[24] ? sfd__h22484[23:1] : sfd__h22484[22:0] ;
  assign _theResult___sfd__h23433 =
	     sfd__h23023[24] ?
	       ((x__h23008[7:0] == 8'd254) ? 23'd0 : sfd__h23023[23:1]) :
	       sfd__h23023[22:0] ;
  assign _theResult___sfd__h29308 =
	     sfd__h28911[24] ? sfd__h28911[23:1] : sfd__h28911[22:0] ;
  assign _theResult___sfd__h29861 =
	     sfd__h29451[24] ?
	       ((x__h29436[7:0] == 8'd254) ? 23'd0 : sfd__h29451[23:1]) :
	       sfd__h29451[22:0] ;
  assign _theResult___sfd__h35479 =
	     sfd__h35082[24] ? sfd__h35082[23:1] : sfd__h35082[22:0] ;
  assign _theResult___sfd__h36031 =
	     sfd__h35621[24] ?
	       ((x__h35606[7:0] == 8'd254) ? 23'd0 : sfd__h35621[23:1]) :
	       sfd__h35621[22:0] ;
  assign _theResult___sfd__h60904 =
	     sfd__h60304[53] ? sfd__h60304[52:1] : sfd__h60304[51:0] ;
  assign _theResult___sfd__h61660 =
	     sfd__h61047[53] ?
	       ((x__h61032[10:0] == 11'd2046) ? 52'd0 : sfd__h61047[52:1]) :
	       sfd__h61047[51:0] ;
  assign _theResult___sfd__h70600 =
	     sfd__h70000[53] ? sfd__h70000[52:1] : sfd__h70000[51:0] ;
  assign _theResult___sfd__h71355 =
	     sfd__h70742[53] ?
	       ((x__h70727[10:0] == 11'd2046) ? 52'd0 : sfd__h70742[52:1]) :
	       sfd__h70742[51:0] ;
  assign _theResult___sfd__h84445 =
	     sfd__h83845[53] ? sfd__h83845[52:1] : sfd__h83845[51:0] ;
  assign _theResult___sfd__h85201 =
	     sfd__h84588[53] ?
	       ((x__h84573[10:0] == 11'd2046) ? 52'd0 : sfd__h84588[52:1]) :
	       sfd__h84588[51:0] ;
  assign _theResult___sfd__h95457 =
	     sfd__h94857[53] ? sfd__h94857[52:1] : sfd__h94857[51:0] ;
  assign _theResult___sfd__h96212 =
	     sfd__h95599[53] ?
	       ((x__h95584[10:0] == 11'd2046) ? 52'd0 : sfd__h95599[52:1]) :
	       sfd__h95599[51:0] ;
  assign _theResult___snd__h119475 = { _theResult____h111357[55:0], 1'd0 } ;
  assign _theResult___snd__h119486 =
	     (!_theResult____h111357[56] && _theResult____h111357[55]) ?
	       _theResult___snd__h119488 :
	       _theResult___snd__h119498 ;
  assign _theResult___snd__h119488 = { _theResult____h111357[54:0], 2'd0 } ;
  assign _theResult___snd__h119498 =
	     (!_theResult____h111357[56] && !_theResult____h111357[55] &&
	      !_theResult____h111357[54] &&
	      !_theResult____h111357[53] &&
	      !_theResult____h111357[52] &&
	      !_theResult____h111357[51] &&
	      !_theResult____h111357[50] &&
	      !_theResult____h111357[49] &&
	      !_theResult____h111357[48] &&
	      !_theResult____h111357[47] &&
	      !_theResult____h111357[46] &&
	      !_theResult____h111357[45] &&
	      !_theResult____h111357[44] &&
	      !_theResult____h111357[43] &&
	      !_theResult____h111357[42] &&
	      !_theResult____h111357[41] &&
	      !_theResult____h111357[40] &&
	      !_theResult____h111357[39] &&
	      !_theResult____h111357[38] &&
	      !_theResult____h111357[37] &&
	      !_theResult____h111357[36] &&
	      !_theResult____h111357[35] &&
	      !_theResult____h111357[34] &&
	      !_theResult____h111357[33] &&
	      !_theResult____h111357[32] &&
	      !_theResult____h111357[31] &&
	      !_theResult____h111357[30] &&
	      !_theResult____h111357[29] &&
	      !_theResult____h111357[28] &&
	      !_theResult____h111357[27] &&
	      !_theResult____h111357[26] &&
	      !_theResult____h111357[25] &&
	      !_theResult____h111357[24] &&
	      !_theResult____h111357[23] &&
	      !_theResult____h111357[22] &&
	      !_theResult____h111357[21] &&
	      !_theResult____h111357[20] &&
	      !_theResult____h111357[19] &&
	      !_theResult____h111357[18] &&
	      !_theResult____h111357[17] &&
	      !_theResult____h111357[16] &&
	      !_theResult____h111357[15] &&
	      !_theResult____h111357[14] &&
	      !_theResult____h111357[13] &&
	      !_theResult____h111357[12] &&
	      !_theResult____h111357[11] &&
	      !_theResult____h111357[10] &&
	      !_theResult____h111357[9] &&
	      !_theResult____h111357[8] &&
	      !_theResult____h111357[7] &&
	      !_theResult____h111357[6] &&
	      !_theResult____h111357[5] &&
	      !_theResult____h111357[4] &&
	      !_theResult____h111357[3] &&
	      !_theResult____h111357[2] &&
	      !_theResult____h111357[1] &&
	      !_theResult____h111357[0]) ?
	       _theResult____h111357 :
	       _theResult___snd__h119504 ;
  assign _theResult___snd__h119504 =
	     { IF_0_CONCAT_IF_IF_0b0_CONCAT_NOT_requestR_BITS_ETC__q114[54:0],
	       2'd0 } ;
  assign _theResult___snd__h119527 =
	     _theResult____h111357 <<
	     IF_IF_0b0_CONCAT_NOT_requestR_BITS_190_TO_180__ETC___d3537 ;
  assign _theResult___snd__h128101 =
	     (requestR[190:180] == 11'd0) ?
	       _theResult___snd__h128110 :
	       _theResult___snd__h128103 ;
  assign _theResult___snd__h128103 = { requestR[179:128], 5'd0 } ;
  assign _theResult___snd__h128110 =
	     (requestR[190:180] == 11'd0 &&
	      NOT_requestR_BIT_179_71_72_AND_NOT_requestR_BI_ETC___d824) ?
	       sfd__h103727 :
	       _theResult___snd__h128116 ;
  assign _theResult___snd__h128116 =
	     { IF_0_CONCAT_IF_requestR_BITS_190_TO_180_599_EQ_ETC__q116[54:0],
	       2'd0 } ;
  assign _theResult___snd__h128139 =
	     sfd__h103727 <<
	     IF_requestR_BITS_190_TO_180_599_EQ_0_609_THEN__ETC___d3659 ;
  assign _theResult___snd__h137328 = { _theResult____h129081[55:0], 1'd0 } ;
  assign _theResult___snd__h137339 =
	     (!_theResult____h129081[56] && _theResult____h129081[55]) ?
	       _theResult___snd__h137341 :
	       _theResult___snd__h137351 ;
  assign _theResult___snd__h137341 = { _theResult____h129081[54:0], 2'd0 } ;
  assign _theResult___snd__h137351 =
	     (!_theResult____h129081[56] && !_theResult____h129081[55] &&
	      !_theResult____h129081[54] &&
	      !_theResult____h129081[53] &&
	      !_theResult____h129081[52] &&
	      !_theResult____h129081[51] &&
	      !_theResult____h129081[50] &&
	      !_theResult____h129081[49] &&
	      !_theResult____h129081[48] &&
	      !_theResult____h129081[47] &&
	      !_theResult____h129081[46] &&
	      !_theResult____h129081[45] &&
	      !_theResult____h129081[44] &&
	      !_theResult____h129081[43] &&
	      !_theResult____h129081[42] &&
	      !_theResult____h129081[41] &&
	      !_theResult____h129081[40] &&
	      !_theResult____h129081[39] &&
	      !_theResult____h129081[38] &&
	      !_theResult____h129081[37] &&
	      !_theResult____h129081[36] &&
	      !_theResult____h129081[35] &&
	      !_theResult____h129081[34] &&
	      !_theResult____h129081[33] &&
	      !_theResult____h129081[32] &&
	      !_theResult____h129081[31] &&
	      !_theResult____h129081[30] &&
	      !_theResult____h129081[29] &&
	      !_theResult____h129081[28] &&
	      !_theResult____h129081[27] &&
	      !_theResult____h129081[26] &&
	      !_theResult____h129081[25] &&
	      !_theResult____h129081[24] &&
	      !_theResult____h129081[23] &&
	      !_theResult____h129081[22] &&
	      !_theResult____h129081[21] &&
	      !_theResult____h129081[20] &&
	      !_theResult____h129081[19] &&
	      !_theResult____h129081[18] &&
	      !_theResult____h129081[17] &&
	      !_theResult____h129081[16] &&
	      !_theResult____h129081[15] &&
	      !_theResult____h129081[14] &&
	      !_theResult____h129081[13] &&
	      !_theResult____h129081[12] &&
	      !_theResult____h129081[11] &&
	      !_theResult____h129081[10] &&
	      !_theResult____h129081[9] &&
	      !_theResult____h129081[8] &&
	      !_theResult____h129081[7] &&
	      !_theResult____h129081[6] &&
	      !_theResult____h129081[5] &&
	      !_theResult____h129081[4] &&
	      !_theResult____h129081[3] &&
	      !_theResult____h129081[2] &&
	      !_theResult____h129081[1] &&
	      !_theResult____h129081[0]) ?
	       _theResult____h129081 :
	       _theResult___snd__h137357 ;
  assign _theResult___snd__h137357 =
	     { IF_0_CONCAT_IF_IF_3970_MINUS_SEXT_requestR_BIT_ETC__q119[54:0],
	       2'd0 } ;
  assign _theResult___snd__h137380 =
	     _theResult____h129081 <<
	     IF_IF_3970_MINUS_SEXT_requestR_BITS_190_TO_180_ETC___d3981 ;
  assign _theResult___snd__h145978 =
	     (requestR[190:180] == 11'd0) ?
	       _theResult___snd__h145992 :
	       _theResult___snd__h128103 ;
  assign _theResult___snd__h145992 =
	     (requestR[190:180] == 11'd0 &&
	      NOT_requestR_BIT_179_71_72_AND_NOT_requestR_BI_ETC___d824) ?
	       sfd__h103727 :
	       _theResult___snd__h145998 ;
  assign _theResult___snd__h145998 =
	     { IF_0_CONCAT_IF_requestR_BITS_190_TO_180_599_EQ_ETC__q122[54:0],
	       2'd0 } ;
  assign _theResult___snd__h146016 =
	     sfd__h103727 <<
	     IF_SEXT_requestR_BITS_190_TO_180_599_MINUS_102_ETC___d4055 ;
  assign _theResult___snd__h169030 =
	     (sV1_exp__h823 == 8'd0) ?
	       _theResult___snd__h169039 :
	       _theResult___snd__h169032 ;
  assign _theResult___snd__h169032 = { sV1_sfd__h824, 34'd0 } ;
  assign _theResult___snd__h169039 =
	     (sV1_exp__h823 == 8'd0 && !sV1_sfd__h824[22] &&
	      NOT_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFF_ETC___d4468) ?
	       b__h39582 :
	       _theResult___snd__h169045 ;
  assign _theResult___snd__h169045 =
	     { IF_0_CONCAT_IF_IF_requestR_BITS_191_TO_160_4_E_ETC__q148[54:0],
	       2'd0 } ;
  assign _theResult___snd__h169068 =
	     b__h39582 <<
	     IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_ETC___d4495 ;
  assign _theResult___snd__h178663 = { _theResult____h170416[55:0], 1'd0 } ;
  assign _theResult___snd__h178674 =
	     (!_theResult____h170416[56] && _theResult____h170416[55]) ?
	       _theResult___snd__h178676 :
	       _theResult___snd__h178686 ;
  assign _theResult___snd__h178676 = { _theResult____h170416[54:0], 2'd0 } ;
  assign _theResult___snd__h178686 =
	     (!_theResult____h170416[56] && !_theResult____h170416[55] &&
	      !_theResult____h170416[54] &&
	      !_theResult____h170416[53] &&
	      !_theResult____h170416[52] &&
	      !_theResult____h170416[51] &&
	      !_theResult____h170416[50] &&
	      !_theResult____h170416[49] &&
	      !_theResult____h170416[48] &&
	      !_theResult____h170416[47] &&
	      !_theResult____h170416[46] &&
	      !_theResult____h170416[45] &&
	      !_theResult____h170416[44] &&
	      !_theResult____h170416[43] &&
	      !_theResult____h170416[42] &&
	      !_theResult____h170416[41] &&
	      !_theResult____h170416[40] &&
	      !_theResult____h170416[39] &&
	      !_theResult____h170416[38] &&
	      !_theResult____h170416[37] &&
	      !_theResult____h170416[36] &&
	      !_theResult____h170416[35] &&
	      !_theResult____h170416[34] &&
	      !_theResult____h170416[33] &&
	      !_theResult____h170416[32] &&
	      !_theResult____h170416[31] &&
	      !_theResult____h170416[30] &&
	      !_theResult____h170416[29] &&
	      !_theResult____h170416[28] &&
	      !_theResult____h170416[27] &&
	      !_theResult____h170416[26] &&
	      !_theResult____h170416[25] &&
	      !_theResult____h170416[24] &&
	      !_theResult____h170416[23] &&
	      !_theResult____h170416[22] &&
	      !_theResult____h170416[21] &&
	      !_theResult____h170416[20] &&
	      !_theResult____h170416[19] &&
	      !_theResult____h170416[18] &&
	      !_theResult____h170416[17] &&
	      !_theResult____h170416[16] &&
	      !_theResult____h170416[15] &&
	      !_theResult____h170416[14] &&
	      !_theResult____h170416[13] &&
	      !_theResult____h170416[12] &&
	      !_theResult____h170416[11] &&
	      !_theResult____h170416[10] &&
	      !_theResult____h170416[9] &&
	      !_theResult____h170416[8] &&
	      !_theResult____h170416[7] &&
	      !_theResult____h170416[6] &&
	      !_theResult____h170416[5] &&
	      !_theResult____h170416[4] &&
	      !_theResult____h170416[3] &&
	      !_theResult____h170416[2] &&
	      !_theResult____h170416[1] &&
	      !_theResult____h170416[0]) ?
	       _theResult____h170416 :
	       _theResult___snd__h178692 ;
  assign _theResult___snd__h178692 =
	     { IF_0_CONCAT_IF_IF_3074_MINUS_SEXT_IF_requestR__ETC__q151[54:0],
	       2'd0 } ;
  assign _theResult___snd__h178715 =
	     _theResult____h170416 <<
	     IF_IF_3074_MINUS_SEXT_IF_requestR_BITS_191_TO__ETC___d4815 ;
  assign _theResult___snd__h187429 =
	     (sV1_exp__h823 == 8'd0) ?
	       _theResult___snd__h187443 :
	       _theResult___snd__h169032 ;
  assign _theResult___snd__h187443 =
	     (sV1_exp__h823 == 8'd0 && !sV1_sfd__h824[22] &&
	      NOT_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFF_ETC___d4468) ?
	       b__h39582 :
	       _theResult___snd__h187449 ;
  assign _theResult___snd__h187449 =
	     { IF_0_CONCAT_IF_IF_requestR_BITS_191_TO_160_4_E_ETC__q154[54:0],
	       2'd0 } ;
  assign _theResult___snd__h187467 =
	     b__h39582 <<
	     IF_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFFF_ETC___d4889 ;
  assign _theResult___snd_fst_exp__h128706 =
	     _3074_MINUS_0_CONCAT_IF_requestR_BIT_179_71_THE_ETC___d3305 ?
	       _theResult___fst_exp__h120091 :
	       _theResult___fst_exp__h128703 ;
  assign _theResult___snd_fst_exp__h12917 =
	     _64_MINUS_0_CONCAT_IF_IF_requestR_BIT_191_27_TH_ETC___d393 ?
	       _theResult___fst_exp__h12358 :
	       _theResult___fst_exp__h12914 ;
  assign _theResult___snd_fst_exp__h12920 =
	     _64_MINUS_0_CONCAT_IF_IF_requestR_BIT_191_27_TH_ETC___d390 ?
	       8'd0 :
	       _theResult___snd_fst_exp__h12917 ;
  assign _theResult___snd_fst_exp__h12923 =
	     _64_MINUS_0_CONCAT_IF_IF_requestR_BIT_191_27_TH_ETC___d388 ?
	       _theResult___snd_fst_exp__h12920 :
	       8'd255 ;
  assign _theResult___snd_fst_exp__h146613 =
	     SEXT_requestR_BITS_190_TO_180_599_MINUS_1023_6_ETC___d3736 ?
	       _theResult___fst_exp__h137944 :
	       _theResult___fst_exp__h146610 ;
  assign _theResult___snd_fst_exp__h169838 =
	     _3970_MINUS_0_CONCAT_IF_IF_requestR_BITS_191_TO_ETC___d4425 ?
	       11'd0 :
	       _theResult___fst_exp__h169835 ;
  assign _theResult___snd_fst_exp__h188267 =
	     SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFF_ETC___d4568 ?
	       _theResult___fst_exp__h179482 :
	       _theResult___fst_exp__h188264 ;
  assign _theResult___snd_fst_exp__h23534 =
	     _64_MINUS_0_CONCAT_IF_requestR_BIT_191_27_THEN__ETC___d907 ?
	       _theResult___fst_exp__h22976 :
	       _theResult___fst_exp__h23531 ;
  assign _theResult___snd_fst_exp__h23537 =
	     _64_MINUS_0_CONCAT_IF_requestR_BIT_191_27_THEN__ETC___d906 ?
	       8'd0 :
	       _theResult___snd_fst_exp__h23534 ;
  assign _theResult___snd_fst_exp__h23540 =
	     _64_MINUS_0_CONCAT_IF_requestR_BIT_191_27_THEN__ETC___d905 ?
	       _theResult___snd_fst_exp__h23537 :
	       8'd255 ;
  assign _theResult___snd_fst_exp__h29963 =
	     _32_MINUS_0_CONCAT_IF_IF_requestR_BIT_159_6_THE_ETC___d1261 ?
	       _theResult___fst_exp__h29404 :
	       _theResult___fst_exp__h29960 ;
  assign _theResult___snd_fst_exp__h29966 =
	     _32_MINUS_0_CONCAT_IF_IF_requestR_BIT_159_6_THE_ETC___d1258 ?
	       8'd0 :
	       _theResult___snd_fst_exp__h29963 ;
  assign _theResult___snd_fst_exp__h29969 =
	     _32_MINUS_0_CONCAT_IF_IF_requestR_BIT_159_6_THE_ETC___d1256 ?
	       _theResult___snd_fst_exp__h29966 :
	       8'd255 ;
  assign _theResult___snd_fst_exp__h36132 =
	     _32_MINUS_0_CONCAT_IF_requestR_BIT_159_6_THEN_0_ETC___d1513 ?
	       _theResult___fst_exp__h35574 :
	       _theResult___fst_exp__h36129 ;
  assign _theResult___snd_fst_exp__h36135 =
	     _32_MINUS_0_CONCAT_IF_requestR_BIT_159_6_THEN_0_ETC___d1512 ?
	       8'd0 :
	       _theResult___snd_fst_exp__h36132 ;
  assign _theResult___snd_fst_exp__h36138 =
	     _32_MINUS_0_CONCAT_IF_requestR_BIT_159_6_THEN_0_ETC___d1511 ?
	       _theResult___snd_fst_exp__h36135 :
	       8'd255 ;
  assign _theResult___snd_fst_exp__h61762 =
	     _32_MINUS_0_CONCAT_IF_IF_requestR_BIT_159_6_THE_ETC___d2238 ?
	       _theResult___fst_exp__h61000 :
	       _theResult___fst_exp__h61759 ;
  assign _theResult___snd_fst_exp__h61765 =
	     _32_MINUS_0_CONCAT_IF_IF_requestR_BIT_159_6_THE_ETC___d2236 ?
	       11'd0 :
	       _theResult___snd_fst_exp__h61762 ;
  assign _theResult___snd_fst_exp__h61768 =
	     _32_MINUS_0_CONCAT_IF_IF_requestR_BIT_159_6_THE_ETC___d2234 ?
	       _theResult___snd_fst_exp__h61765 :
	       11'd2047 ;
  assign _theResult___snd_fst_exp__h71456 =
	     _32_MINUS_0_CONCAT_IF_requestR_BIT_159_6_THEN_0_ETC___d2451 ?
	       _theResult___fst_exp__h70695 :
	       _theResult___fst_exp__h71453 ;
  assign _theResult___snd_fst_exp__h71459 =
	     _32_MINUS_0_CONCAT_IF_requestR_BIT_159_6_THEN_0_ETC___d2450 ?
	       11'd0 :
	       _theResult___snd_fst_exp__h71456 ;
  assign _theResult___snd_fst_exp__h71462 =
	     _32_MINUS_0_CONCAT_IF_requestR_BIT_159_6_THEN_0_ETC___d2449 ?
	       _theResult___snd_fst_exp__h71459 :
	       11'd2047 ;
  assign _theResult___snd_fst_exp__h85303 =
	     _64_MINUS_0_CONCAT_IF_IF_requestR_BIT_191_27_TH_ETC___d2775 ?
	       _theResult___fst_exp__h84541 :
	       _theResult___fst_exp__h85300 ;
  assign _theResult___snd_fst_exp__h85306 =
	     _64_MINUS_0_CONCAT_IF_IF_requestR_BIT_191_27_TH_ETC___d2772 ?
	       11'd0 :
	       _theResult___snd_fst_exp__h85303 ;
  assign _theResult___snd_fst_exp__h85309 =
	     _64_MINUS_0_CONCAT_IF_IF_requestR_BIT_191_27_TH_ETC___d2770 ?
	       _theResult___snd_fst_exp__h85306 :
	       11'd2047 ;
  assign _theResult___snd_fst_exp__h96313 =
	     _64_MINUS_0_CONCAT_IF_requestR_BIT_191_27_THEN__ETC___d2957 ?
	       _theResult___fst_exp__h95552 :
	       _theResult___fst_exp__h96310 ;
  assign _theResult___snd_fst_exp__h96316 =
	     _64_MINUS_0_CONCAT_IF_requestR_BIT_191_27_THEN__ETC___d2956 ?
	       11'd0 :
	       _theResult___snd_fst_exp__h96313 ;
  assign _theResult___snd_fst_exp__h96319 =
	     _64_MINUS_0_CONCAT_IF_requestR_BIT_191_27_THEN__ETC___d2955 ?
	       _theResult___snd_fst_exp__h96316 :
	       11'd2047 ;
  assign _theResult___snd_fst_sfd__h103681 =
	     (value__h99566[51:29] == 23'd0) ?
	       23'd2097152 :
	       value__h99566[51:29] ;
  assign _theResult___snd_fst_sfd__h128707 =
	     _3074_MINUS_0_CONCAT_IF_requestR_BIT_179_71_THE_ETC___d3305 ?
	       _theResult___fst_sfd__h120092 :
	       _theResult___fst_sfd__h128704 ;
  assign _theResult___snd_fst_sfd__h12918 =
	     _64_MINUS_0_CONCAT_IF_IF_requestR_BIT_191_27_TH_ETC___d393 ?
	       _theResult___fst_sfd__h12359 :
	       _theResult___fst_sfd__h12915 ;
  assign _theResult___snd_fst_sfd__h146614 =
	     SEXT_requestR_BITS_190_TO_180_599_MINUS_1023_6_ETC___d3736 ?
	       _theResult___fst_sfd__h137945 :
	       _theResult___fst_sfd__h146611 ;
  assign _theResult___snd_fst_sfd__h150153 =
	     (value__h148270 == 23'd0) ?
	       52'h4000000000000 :
	       out___1_sfd__h148267 ;
  assign _theResult___snd_fst_sfd__h169839 =
	     _3970_MINUS_0_CONCAT_IF_IF_requestR_BITS_191_TO_ETC___d4425 ?
	       52'd0 :
	       _theResult___fst_sfd__h169836 ;
  assign _theResult___snd_fst_sfd__h188268 =
	     SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFF_ETC___d4568 ?
	       _theResult___fst_sfd__h179483 :
	       _theResult___fst_sfd__h188265 ;
  assign _theResult___snd_fst_sfd__h23535 =
	     _64_MINUS_0_CONCAT_IF_requestR_BIT_191_27_THEN__ETC___d907 ?
	       _theResult___fst_sfd__h22977 :
	       _theResult___fst_sfd__h23532 ;
  assign _theResult___snd_fst_sfd__h29964 =
	     _32_MINUS_0_CONCAT_IF_IF_requestR_BIT_159_6_THE_ETC___d1261 ?
	       _theResult___fst_sfd__h29405 :
	       _theResult___fst_sfd__h29961 ;
  assign _theResult___snd_fst_sfd__h36133 =
	     _32_MINUS_0_CONCAT_IF_requestR_BIT_159_6_THEN_0_ETC___d1513 ?
	       _theResult___fst_sfd__h35575 :
	       _theResult___fst_sfd__h36130 ;
  assign _theResult___snd_fst_sfd__h61763 =
	     _32_MINUS_0_CONCAT_IF_IF_requestR_BIT_159_6_THE_ETC___d2238 ?
	       _theResult___fst_sfd__h61001 :
	       _theResult___fst_sfd__h61760 ;
  assign _theResult___snd_fst_sfd__h71457 =
	     _32_MINUS_0_CONCAT_IF_requestR_BIT_159_6_THEN_0_ETC___d2451 ?
	       _theResult___fst_sfd__h70696 :
	       _theResult___fst_sfd__h71454 ;
  assign _theResult___snd_fst_sfd__h85304 =
	     _64_MINUS_0_CONCAT_IF_IF_requestR_BIT_191_27_TH_ETC___d2775 ?
	       _theResult___fst_sfd__h84542 :
	       _theResult___fst_sfd__h85301 ;
  assign _theResult___snd_fst_sfd__h96314 =
	     _64_MINUS_0_CONCAT_IF_requestR_BIT_191_27_THEN__ETC___d2957 ?
	       _theResult___fst_sfd__h95553 :
	       _theResult___fst_sfd__h96311 ;
  assign ab__h206728 = dw_result$wget ;
  assign b__h36799 = { value__h36801, 64'd0 } ;
  assign b__h39582 = { value__h36801, 32'd0 } ;
  assign b__h72122 = { value__h72124, 32'd0 } ;
  assign b__h96976 = { value__h72124, 64'd0 } ;
  assign din_inc___2_exp__h12957 = x__h12390[7:0] + 8'd1 ;
  assign din_inc___2_exp__h146641 = _theResult___fst_exp__h119464 + 8'd1 ;
  assign din_inc___2_exp__h146665 = _theResult___fst_exp__h128150 + 8'd1 ;
  assign din_inc___2_exp__h146695 = _theResult___fst_exp__h137317 + 8'd1 ;
  assign din_inc___2_exp__h146719 = _theResult___fst_exp__h146032 + 8'd1 ;
  assign din_inc___2_exp__h188299 = _theResult___fst_exp__h169079 + 11'd1 ;
  assign din_inc___2_exp__h188329 = _theResult___fst_exp__h178652 + 11'd1 ;
  assign din_inc___2_exp__h188353 = _theResult___fst_exp__h187483 + 11'd1 ;
  assign din_inc___2_exp__h23570 = x__h23008[7:0] + 8'd1 ;
  assign din_inc___2_exp__h30003 = x__h29436[7:0] + 8'd1 ;
  assign din_inc___2_exp__h36168 = x__h35606[7:0] + 8'd1 ;
  assign din_inc___2_exp__h61802 = x__h61032[10:0] + 11'd1 ;
  assign din_inc___2_exp__h71492 = x__h70727[10:0] + 11'd1 ;
  assign din_inc___2_exp__h85343 = x__h84573[10:0] + 11'd1 ;
  assign din_inc___2_exp__h96349 = x__h95584[10:0] + 11'd1 ;
  assign guard__h111367 =
	     { IF_sfdin19458_BIT_33_THEN_2_ELSE_0__q115[1],
	       { sfdin__h119458[32:0], 23'd0 } != 56'd0 } ;
  assign guard__h11845 =
	     { IF_sfd___31835_BIT_40_THEN_2_ELSE_0__q6[1],
	       { sfd___3__h11835[39:0], 23'd0 } != 63'd0 } ;
  assign guard__h120102 =
	     { IF_theResult___snd28101_BIT_33_THEN_2_ELSE_0__q117[1],
	       { _theResult___snd__h128101[32:0], 23'd0 } != 56'd0 } ;
  assign guard__h12375 =
	     { IF_sfd___31835_BIT_39_THEN_2_ELSE_0__q7[1],
	       { sfd___3__h11835[38:0], 24'd0 } != 63'd0 } ;
  assign guard__h129091 =
	     { IF_sfdin37311_BIT_33_THEN_2_ELSE_0__q120[1],
	       { sfdin__h137311[32:0], 23'd0 } != 56'd0 } ;
  assign guard__h129689 = x__h129789 != 57'd0 ;
  assign guard__h137955 =
	     { IF_theResult___snd45978_BIT_33_THEN_2_ELSE_0__q123[1],
	       { _theResult___snd__h145978[32:0], 23'd0 } != 56'd0 } ;
  assign guard__h161118 =
	     { IF_theResult___snd69030_BIT_4_THEN_2_ELSE_0__q149[1],
	       { _theResult___snd__h169030[3:0], 52'd0 } != 56'd0 } ;
  assign guard__h170426 =
	     { IF_sfdin78646_BIT_4_THEN_2_ELSE_0__q152[1],
	       { sfdin__h178646[3:0], 52'd0 } != 56'd0 } ;
  assign guard__h171024 = x__h171124 != 57'd0 ;
  assign guard__h179493 =
	     { IF_theResult___snd87429_BIT_4_THEN_2_ELSE_0__q155[1],
	       { _theResult___snd__h187429[3:0], 52'd0 } != 56'd0 } ;
  assign guard__h22467 =
	     { IF_sfd___32457_BIT_40_THEN_2_ELSE_0__q22[1],
	       { sfd___3__h22457[39:0], 23'd0 } != 63'd0 } ;
  assign guard__h22993 =
	     { IF_sfd___32457_BIT_39_THEN_2_ELSE_0__q23[1],
	       { sfd___3__h22457[38:0], 24'd0 } != 63'd0 } ;
  assign guard__h28894 =
	     { IF_sfd___38884_BIT_8_THEN_2_ELSE_0__q38[1],
	       { sfd___3__h28884[7:0], 23'd0 } != 31'd0 } ;
  assign guard__h29421 =
	     { IF_sfd___38884_BIT_7_THEN_2_ELSE_0__q39[1],
	       { sfd___3__h28884[6:0], 24'd0 } != 31'd0 } ;
  assign guard__h35065 =
	     { IF_sfd___35055_BIT_8_THEN_2_ELSE_0__q52[1],
	       { sfd___3__h35055[7:0], 23'd0 } != 31'd0 } ;
  assign guard__h35591 =
	     { IF_sfd___35055_BIT_7_THEN_2_ELSE_0__q53[1],
	       { sfd___3__h35055[6:0], 24'd0 } != 31'd0 } ;
  assign guard__h36732 =
	     { IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d1689[23],
	       { IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d1689[22:0],
		 65'd0 } !=
	       88'd0 } ;
  assign guard__h37510 =
	     { IF_x7699_BIT_24_THEN_2_ELSE_0__q63[1],
	       { x__h37699[23:0], 64'd0 } != 88'd0 } ;
  assign guard__h38794 =
	     { IF_x9015_BIT_24_THEN_2_ELSE_0__q64[1],
	       { x__h39015[23:0], 64'd0 } != 88'd0 } ;
  assign guard__h39515 =
	     { IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d1838[23],
	       { IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d1838[22:0],
		 33'd0 } !=
	       56'd0 } ;
  assign guard__h40069 =
	     { IF_x0258_BIT_24_THEN_2_ELSE_0__q65[1],
	       { x__h40258[23:0], 32'd0 } != 56'd0 } ;
  assign guard__h41115 =
	     { IF_x1336_BIT_24_THEN_2_ELSE_0__q66[1],
	       { x__h41336[23:0], 32'd0 } != 56'd0 } ;
  assign guard__h60287 =
	     { IF_sfd___30277_BIT_2_THEN_2_ELSE_0__q67[1],
	       { sfd___3__h60277[1:0], 52'd0 } != 54'd0 } ;
  assign guard__h61017 =
	     { IF_sfd___30277_BIT_1_THEN_2_ELSE_0__q68[1],
	       { sfd___3__h60277[0], 53'd0 } != 54'd0 } ;
  assign guard__h69983 =
	     { IF_sfd___39973_BIT_2_THEN_2_ELSE_0__q81[1],
	       { sfd___3__h69973[1:0], 52'd0 } != 54'd0 } ;
  assign guard__h70712 =
	     { IF_sfd___39973_BIT_1_THEN_2_ELSE_0__q82[1],
	       { sfd___3__h69973[0], 53'd0 } != 54'd0 } ;
  assign guard__h72055 =
	     { IF_requestR_BIT_191_27_THEN_NEG_0b0_CONCAT_NOT_ETC___d2620[52],
	       { IF_requestR_BIT_191_27_THEN_NEG_0b0_CONCAT_NOT_ETC___d2620[51:0],
		 33'd0 } !=
	       85'd0 } ;
  assign guard__h72609 =
	     { IF_x2798_BIT_53_THEN_2_ELSE_0__q92[1],
	       { x__h72798[52:0], 32'd0 } != 85'd0 } ;
  assign guard__h73655 =
	     { IF_x3876_BIT_53_THEN_2_ELSE_0__q93[1],
	       { x__h73876[52:0], 32'd0 } != 85'd0 } ;
  assign guard__h83828 =
	     { IF_sfd___31835_BIT_11_THEN_2_ELSE_0__q8[1],
	       { sfd___3__h11835[10:0], 52'd0 } != 63'd0 } ;
  assign guard__h84558 =
	     { IF_sfd___31835_BIT_10_THEN_2_ELSE_0__q9[1],
	       { sfd___3__h11835[9:0], 53'd0 } != 63'd0 } ;
  assign guard__h94840 =
	     { IF_sfd___32457_BIT_11_THEN_2_ELSE_0__q24[1],
	       { sfd___3__h22457[10:0], 52'd0 } != 63'd0 } ;
  assign guard__h95569 =
	     { IF_sfd___32457_BIT_10_THEN_2_ELSE_0__q25[1],
	       { sfd___3__h22457[9:0], 53'd0 } != 63'd0 } ;
  assign guard__h96909 =
	     { IF_requestR_BIT_191_27_THEN_NEG_0b0_CONCAT_NOT_ETC___d3109[52],
	       { IF_requestR_BIT_191_27_THEN_NEG_0b0_CONCAT_NOT_ETC___d3109[51:0],
		 65'd0 } !=
	       117'd0 } ;
  assign guard__h97687 =
	     { IF_x7876_BIT_53_THEN_2_ELSE_0__q112[1],
	       { x__h97876[52:0], 64'd0 } != 117'd0 } ;
  assign guard__h98954 =
	     { IF_x9175_BIT_53_THEN_2_ELSE_0__q113[1],
	       { x__h99175[52:0], 64'd0 } != 117'd0 } ;
  assign out1___1__h37450 =
	     IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d1689[88:24] +
	     65'd1 ;
  assign out1___1__h40009 =
	     IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d1838[56:24] +
	     33'd1 ;
  assign out1___1__h72549 =
	     IF_requestR_BIT_191_27_THEN_NEG_0b0_CONCAT_NOT_ETC___d2620[85:53] +
	     33'd1 ;
  assign out1___1__h97627 =
	     IF_requestR_BIT_191_27_THEN_NEG_0b0_CONCAT_NOT_ETC___d3109[117:53] +
	     65'd1 ;
  assign out___1_sfd__h148267 = { value__h148270, 29'd0 } ;
  assign out_exp__h119993 =
	     sfdin__h119458[34] ?
	       _theResult___exp__h119990 :
	       _theResult___fst_exp__h119464 ;
  assign out_exp__h12264 =
	     sfd___3__h11835[41] ? _theResult___exp__h12261 : 8'd0 ;
  assign out_exp__h12817 =
	     sfd___3__h11835[40] ? _theResult___exp__h12814 : x__h12390[7:0] ;
  assign out_exp__h128605 =
	     _theResult___snd__h128101[34] ?
	       _theResult___exp__h128602 :
	       _theResult___fst_exp__h128150 ;
  assign out_exp__h137846 =
	     sfdin__h137311[34] ?
	       _theResult___exp__h137843 :
	       _theResult___fst_exp__h137317 ;
  assign out_exp__h146512 =
	     _theResult___snd__h145978[34] ?
	       _theResult___exp__h146509 :
	       _theResult___fst_exp__h146032 ;
  assign out_exp__h169737 =
	     _theResult___snd__h169030[5] ?
	       _theResult___exp__h169734 :
	       _theResult___fst_exp__h169079 ;
  assign out_exp__h179384 =
	     sfdin__h178646[5] ?
	       _theResult___exp__h179381 :
	       _theResult___fst_exp__h178652 ;
  assign out_exp__h188166 =
	     _theResult___snd__h187429[5] ?
	       _theResult___exp__h188163 :
	       _theResult___fst_exp__h187483 ;
  assign out_exp__h22883 =
	     sfd___3__h22457[41] ? _theResult___exp__h22880 : 8'd0 ;
  assign out_exp__h23435 =
	     sfd___3__h22457[40] ? _theResult___exp__h23432 : x__h23008[7:0] ;
  assign out_exp__h29310 =
	     sfd___3__h28884[9] ? _theResult___exp__h29307 : 8'd0 ;
  assign out_exp__h29863 =
	     sfd___3__h28884[8] ? _theResult___exp__h29860 : x__h29436[7:0] ;
  assign out_exp__h35481 =
	     sfd___3__h35055[9] ? _theResult___exp__h35478 : 8'd0 ;
  assign out_exp__h36033 =
	     sfd___3__h35055[8] ? _theResult___exp__h36030 : x__h35606[7:0] ;
  assign out_exp__h60906 =
	     sfd___3__h60277[3] ? _theResult___exp__h60903 : 11'd0 ;
  assign out_exp__h61662 =
	     sfd___3__h60277[2] ? _theResult___exp__h61659 : x__h61032[10:0] ;
  assign out_exp__h70602 =
	     sfd___3__h69973[3] ? _theResult___exp__h70599 : 11'd0 ;
  assign out_exp__h71357 =
	     sfd___3__h69973[2] ? _theResult___exp__h71354 : x__h70727[10:0] ;
  assign out_exp__h84447 =
	     sfd___3__h11835[12] ? _theResult___exp__h84444 : 11'd0 ;
  assign out_exp__h85203 =
	     sfd___3__h11835[11] ?
	       _theResult___exp__h85200 :
	       x__h84573[10:0] ;
  assign out_exp__h95459 =
	     sfd___3__h22457[12] ? _theResult___exp__h95456 : 11'd0 ;
  assign out_exp__h96214 =
	     sfd___3__h22457[11] ?
	       _theResult___exp__h96211 :
	       x__h95584[10:0] ;
  assign out_sfd__h119994 =
	     sfdin__h119458[34] ?
	       _theResult___sfd__h119991 :
	       sfdin__h119458[56:34] ;
  assign out_sfd__h12265 =
	     sfd___3__h11835[41] ?
	       _theResult___sfd__h12262 :
	       sfd___3__h11835[63:41] ;
  assign out_sfd__h12818 =
	     sfd___3__h11835[40] ?
	       _theResult___sfd__h12815 :
	       sfd___3__h11835[62:40] ;
  assign out_sfd__h128606 =
	     _theResult___snd__h128101[34] ?
	       _theResult___sfd__h128603 :
	       _theResult___snd__h128101[56:34] ;
  assign out_sfd__h137847 =
	     sfdin__h137311[34] ?
	       _theResult___sfd__h137844 :
	       sfdin__h137311[56:34] ;
  assign out_sfd__h146513 =
	     _theResult___snd__h145978[34] ?
	       _theResult___sfd__h146510 :
	       _theResult___snd__h145978[56:34] ;
  assign out_sfd__h169738 =
	     _theResult___snd__h169030[5] ?
	       _theResult___sfd__h169735 :
	       _theResult___snd__h169030[56:5] ;
  assign out_sfd__h179385 =
	     sfdin__h178646[5] ?
	       _theResult___sfd__h179382 :
	       sfdin__h178646[56:5] ;
  assign out_sfd__h188167 =
	     _theResult___snd__h187429[5] ?
	       _theResult___sfd__h188164 :
	       _theResult___snd__h187429[56:5] ;
  assign out_sfd__h22884 =
	     sfd___3__h22457[41] ?
	       _theResult___sfd__h22881 :
	       sfd___3__h22457[63:41] ;
  assign out_sfd__h23436 =
	     sfd___3__h22457[40] ?
	       _theResult___sfd__h23433 :
	       sfd___3__h22457[62:40] ;
  assign out_sfd__h29311 =
	     sfd___3__h28884[9] ?
	       _theResult___sfd__h29308 :
	       sfd___3__h28884[31:9] ;
  assign out_sfd__h29864 =
	     sfd___3__h28884[8] ?
	       _theResult___sfd__h29861 :
	       sfd___3__h28884[30:8] ;
  assign out_sfd__h35482 =
	     sfd___3__h35055[9] ?
	       _theResult___sfd__h35479 :
	       sfd___3__h35055[31:9] ;
  assign out_sfd__h36034 =
	     sfd___3__h35055[8] ?
	       _theResult___sfd__h36031 :
	       sfd___3__h35055[30:8] ;
  assign out_sfd__h60907 =
	     sfd___3__h60277[3] ?
	       _theResult___sfd__h60904 :
	       sfd___3__h60277[54:3] ;
  assign out_sfd__h61663 =
	     sfd___3__h60277[2] ?
	       _theResult___sfd__h61660 :
	       sfd___3__h60277[53:2] ;
  assign out_sfd__h70603 =
	     sfd___3__h69973[3] ?
	       _theResult___sfd__h70600 :
	       sfd___3__h69973[54:3] ;
  assign out_sfd__h71358 =
	     sfd___3__h69973[2] ?
	       _theResult___sfd__h71355 :
	       sfd___3__h69973[53:2] ;
  assign out_sfd__h84448 =
	     sfd___3__h11835[12] ?
	       _theResult___sfd__h84445 :
	       sfd___3__h11835[63:12] ;
  assign out_sfd__h85204 =
	     sfd___3__h11835[11] ?
	       _theResult___sfd__h85201 :
	       sfd___3__h11835[62:11] ;
  assign out_sfd__h95460 =
	     sfd___3__h22457[12] ?
	       _theResult___sfd__h95457 :
	       sfd___3__h22457[63:12] ;
  assign out_sfd__h96215 =
	     sfd___3__h22457[11] ?
	       _theResult___sfd__h96212 :
	       sfd___3__h22457[62:11] ;
  assign requestR_BITS_126_TO_116_166_EQ_0_180_AND_requ_ETC___d5187 =
	     requestR[126:116] == 11'd0 && requestR[115:64] == 52'd0 &&
	     requestR[127] &&
	     requestR[190:180] == 11'd0 &&
	     requestR[179:128] == 52'd0 &&
	     !requestR[191] ;
  assign requestR_BITS_127_TO_96_2_EQ_0xFFFFFFFF_3_AND__ETC___d28 =
	     { requestR[127:96] == 32'hFFFFFFFF && requestR[95],
	       (requestR[127:96] == 32'hFFFFFFFF) ?
		 requestR[94:64] :
		 31'h7FC00000 } ;
  assign requestR_BITS_159_TO_128__q1 = requestR[159:128] ;
  assign requestR_BITS_179_TO_128_601_ULE_requestR_BITS_ETC___d5199 =
	     requestR[179:128] <= requestR[115:64] ;
  assign requestR_BITS_179_TO_128_601_ULT_requestR_BITS_ETC___d5204 =
	     requestR[179:128] < requestR[115:64] ;
  assign requestR_BITS_190_TO_180_599_EQ_0_609_AND_requ_ETC___d5183 =
	     requestR[190:180] == 11'd0 && requestR[179:128] == 52'd0 &&
	     requestR[191] &&
	     requestR[126:116] == 11'd0 &&
	     requestR[115:64] == 52'd0 &&
	     !requestR[127] ;
  assign requestR_BITS_190_TO_180_599_EQ_0_609_AND_requ_ETC___d5257 =
	     requestR[190:180] == 11'd0 && requestR[179:128] == 52'd0 &&
	     requestR[126:116] == 11'd0 &&
	     requestR[115:64] == 52'd0 ||
	     (!requestR[191] || requestR[127]) &&
	     (requestR[191] || !requestR[127]) &&
	     (requestR[191] ?
		requestR_BITS_190_TO_180_599_ULE_requestR_BITS_ETC___d5252 :
		NOT_requestR_BITS_190_TO_180_599_ULT_requestR__ETC___d5253) ;
  assign requestR_BITS_190_TO_180_599_EQ_2047_600_AND_0_ETC___d2749 =
	     requestR[190:180] == 11'd2047 && requestR[179:128] != 52'd0 ||
	     requestR[190:180] == 11'd2047 && requestR[179:128] == 52'd0 ||
	     (requestR[190:180] != 11'd0 || requestR[179:128] != 52'd0) &&
	     (NEG_SEXT_requestR_BITS_190_TO_180_599_MINUS_10_ETC___d2710[23] ||
	      NEG_SEXT_requestR_BITS_190_TO_180_599_MINUS_10_ETC___d2712 &&
	      IF_requestR_BITS_194_TO_192_0_EQ_0x0_1_OR_NOT__ETC___d2731 &&
	      x__h73876[85:54] == 32'hFFFFFFFF) ;
  assign requestR_BITS_190_TO_180_599_EQ_2047_600_AND_0_ETC___d2760 =
	     { requestR_BITS_190_TO_180_599_EQ_2047_600_AND_0_ETC___d2749,
	       3'd0,
	       (requestR[190:180] != 11'd2047 ||
		requestR[179:128] == 52'd0) &&
	       (requestR[190:180] != 11'd2047 ||
		requestR[179:128] != 52'd0) &&
	       NOT_requestR_BITS_190_TO_180_599_EQ_0_609_615__ETC___d2754 } ==
	     5'd0 ||
	     requestR_BITS_190_TO_180_599_EQ_2047_600_AND_0_ETC___d2749 ;
  assign requestR_BITS_190_TO_180_599_EQ_2047_600_AND_0_ETC___d3230 =
	     requestR[190:180] == 11'd2047 && requestR[179:128] != 52'd0 ||
	     requestR[190:180] == 11'd2047 && requestR[179:128] == 52'd0 ||
	     (requestR[190:180] != 11'd0 || requestR[179:128] != 52'd0) &&
	     (NEG_SEXT_requestR_BITS_190_TO_180_599_MINUS_10_ETC___d3192[23] ||
	      NEG_SEXT_requestR_BITS_190_TO_180_599_MINUS_10_ETC___d3194 &&
	      IF_requestR_BITS_194_TO_192_0_EQ_0x0_1_OR_NOT__ETC___d3213 &&
	      x__h99175[117:54] == 64'hFFFFFFFFFFFFFFFF) ;
  assign requestR_BITS_190_TO_180_599_EQ_2047_600_AND_0_ETC___d3241 =
	     { requestR_BITS_190_TO_180_599_EQ_2047_600_AND_0_ETC___d3230,
	       3'd0,
	       (requestR[190:180] != 11'd2047 ||
		requestR[179:128] == 52'd0) &&
	       (requestR[190:180] != 11'd2047 ||
		requestR[179:128] != 52'd0) &&
	       NOT_requestR_BITS_190_TO_180_599_EQ_0_609_615__ETC___d3235 } ==
	     5'd0 ||
	     requestR_BITS_190_TO_180_599_EQ_2047_600_AND_0_ETC___d3230 ;
  assign requestR_BITS_190_TO_180_599_EQ_2047_600_AND_N_ETC___d5175 =
	     requestR[190:180] == 11'd2047 && requestR[179:128] != 52'd0 &&
	     !requestR[179] &&
	     requestR[126:116] == 11'd2047 &&
	     requestR[115:64] != 52'd0 &&
	     !requestR[115] ;
  assign requestR_BITS_190_TO_180_599_EQ_2047_600_AND_N_ETC___d5220 =
	     requestR[190:180] == 11'd2047 && requestR[179:128] != 52'd0 &&
	     !requestR[179] ||
	     requestR[126:116] == 11'd2047 && requestR[115:64] != 52'd0 &&
	     !requestR[115] ;
  assign requestR_BITS_190_TO_180_599_EQ_2047_600_AND_N_ETC___d5242 =
	     requestR_BITS_190_TO_180_599_EQ_2047_600_AND_N_ETC___d5220 ||
	     requestR[190:180] == 11'd2047 && requestR[179] ||
	     requestR[126:116] == 11'd2047 && requestR[115] ;
  assign requestR_BITS_190_TO_180_599_EQ_requestR_BITS__ETC___d5198 =
	     requestR[190:180] == requestR[126:116] ;
  assign requestR_BITS_190_TO_180_599_MINUS_1023___d2611 =
	     requestR[190:180] - 11'd1023 ;
  assign requestR_BITS_190_TO_180_599_ULE_requestR_BITS_ETC___d5196 =
	     requestR[190:180] <= requestR[126:116] ;
  assign requestR_BITS_190_TO_180_599_ULE_requestR_BITS_ETC___d5252 =
	     requestR_BITS_190_TO_180_599_ULE_requestR_BITS_ETC___d5196 &&
	     (!requestR_BITS_190_TO_180_599_EQ_requestR_BITS__ETC___d5198 ||
	      requestR_BITS_179_TO_128_601_ULE_requestR_BITS_ETC___d5199) &&
	     !requestR_BITS_190_TO_180_599_ULT_requestR_BITS_ETC___d5203 &&
	     (!requestR_BITS_190_TO_180_599_EQ_requestR_BITS__ETC___d5198 ||
	      !requestR_BITS_179_TO_128_601_ULT_requestR_BITS_ETC___d5204) ;
  assign requestR_BITS_190_TO_180_599_ULT_requestR_BITS_ETC___d5203 =
	     requestR[190:180] < requestR[126:116] ;
  assign requestR_BITS_191_TO_128_24_EQ_0_25_OR_NOT_req_ETC___d837 =
	     requestR[191:128] == 64'd0 ||
	     !requestR[191] && !requestR[190] && !requestR[189] &&
	     !requestR[188] &&
	     !requestR[187] &&
	     !requestR[186] &&
	     !requestR[185] &&
	     !requestR[184] &&
	     !requestR[183] &&
	     !requestR[182] &&
	     !requestR[181] &&
	     !requestR[180] &&
	     NOT_requestR_BIT_179_71_72_AND_NOT_requestR_BI_ETC___d824 ;
  assign requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5_AND_ETC___d2031 =
	     requestR[191:160] == 32'hFFFFFFFF && requestR[159] &&
	     (requestR[127:96] != 32'hFFFFFFFF || !requestR[95]) ||
	     (requestR[191:160] == 32'hFFFFFFFF && requestR[159] ||
	      requestR[127:96] != 32'hFFFFFFFF ||
	      !requestR[95]) &&
	     IF_NOT_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFF_ETC___d2029 ;
  assign requestR_BIT_158_12_OR_requestR_BIT_157_14_OR__ETC___d1058 =
	     requestR[158] || requestR[157] || requestR[156] ||
	     requestR[155] ||
	     requestR[154] ||
	     requestR[153] ||
	     requestR[152] ||
	     requestR[151] ||
	     requestR[150] ||
	     requestR[149] ||
	     requestR[148] ||
	     requestR[147] ||
	     requestR[146] ||
	     requestR[145] ||
	     requestR[144] ||
	     requestR[143] ||
	     requestR[142] ||
	     requestR[141] ||
	     requestR[140] ||
	     requestR[139] ||
	     requestR[138] ||
	     requestR[137] ||
	     requestR[136] ||
	     requestR[135] ||
	     requestR[134] ||
	     requestR[133] ||
	     requestR[132] ||
	     requestR[131] ||
	     requestR[130] ||
	     requestR[129] ||
	     requestR[128] ;
  assign requestR_BIT_159_6_OR_requestR_BIT_158_12_OR_r_ETC___d1654 =
	     (requestR[159] ||
	      requestR_BIT_158_12_OR_requestR_BIT_157_14_OR__ETC___d1058) &&
	     _32_MINUS_0_CONCAT_IF_requestR_BIT_159_6_THEN_0_ETC___d1511 &&
	     !_32_MINUS_0_CONCAT_IF_requestR_BIT_159_6_THEN_0_ETC___d1512 &&
	     IF_32_MINUS_0_CONCAT_IF_requestR_BIT_159_6_THE_ETC___d1651 ;
  assign requestR_BIT_179_71_OR_requestR_BIT_178_73_OR__ETC___d1079 =
	     requestR[179] || requestR[178] || requestR[177] ||
	     requestR[176] ||
	     requestR[175] ||
	     requestR[174] ||
	     requestR[173] ||
	     requestR[172] ||
	     requestR[171] ||
	     requestR[170] ||
	     requestR[169] ||
	     requestR[168] ||
	     requestR[167] ||
	     requestR[166] ||
	     requestR[165] ||
	     requestR[164] ||
	     requestR[163] ||
	     requestR[162] ||
	     requestR[161] ||
	     requestR[160] ||
	     requestR[159] ||
	     requestR_BIT_158_12_OR_requestR_BIT_157_14_OR__ETC___d1058 ;
  assign requestR_BIT_191_27_OR_requestR_BIT_190_49_OR__ETC___d1100 =
	     (requestR[191] || requestR[190] || requestR[189] ||
	      requestR[188] ||
	      requestR[187] ||
	      requestR[186] ||
	      requestR[185] ||
	      requestR[184] ||
	      requestR[183] ||
	      requestR[182] ||
	      requestR[181] ||
	      requestR[180] ||
	      requestR_BIT_179_71_OR_requestR_BIT_178_73_OR__ETC___d1079) &&
	     (!_64_MINUS_0_CONCAT_IF_requestR_BIT_191_27_THEN__ETC___d905 ||
	      !_64_MINUS_0_CONCAT_IF_requestR_BIT_191_27_THEN__ETC___d906 &&
	      !_64_MINUS_0_CONCAT_IF_requestR_BIT_191_27_THEN__ETC___d907 &&
	      _theResult___fst_exp__h23531 == 8'd255 &&
	      _theResult___fst_sfd__h23532 == 23'd0) ;
  assign requestR_BIT_191_27_OR_requestR_BIT_190_49_OR__ETC___d1103 =
	     (requestR[191] || requestR[190] || requestR[189] ||
	      requestR[188] ||
	      requestR[187] ||
	      requestR[186] ||
	      requestR[185] ||
	      requestR[184] ||
	      requestR[183] ||
	      requestR[182] ||
	      requestR[181] ||
	      requestR[180] ||
	      requestR_BIT_179_71_OR_requestR_BIT_178_73_OR__ETC___d1079) &&
	     _64_MINUS_0_CONCAT_IF_requestR_BIT_191_27_THEN__ETC___d905 &&
	     _64_MINUS_0_CONCAT_IF_requestR_BIT_191_27_THEN__ETC___d906 ;
  assign requestR_BIT_191_27_OR_requestR_BIT_190_49_OR__ETC___d1112 =
	     (requestR[191] || requestR[190] || requestR[189] ||
	      requestR[188] ||
	      requestR[187] ||
	      requestR[186] ||
	      requestR[185] ||
	      requestR[184] ||
	      requestR[183] ||
	      requestR[182] ||
	      requestR[181] ||
	      requestR[180] ||
	      requestR_BIT_179_71_OR_requestR_BIT_178_73_OR__ETC___d1079) &&
	     _64_MINUS_0_CONCAT_IF_requestR_BIT_191_27_THEN__ETC___d905 &&
	     !_64_MINUS_0_CONCAT_IF_requestR_BIT_191_27_THEN__ETC___d906 &&
	     IF_64_MINUS_0_CONCAT_IF_requestR_BIT_191_27_TH_ETC___d1109 ;
  assign requestR_BIT_191_27_OR_requestR_BIT_190_49_OR__ETC___d3085 =
	     (requestR[191] || requestR[190] || requestR[189] ||
	      requestR[188] ||
	      requestR[187] ||
	      requestR[186] ||
	      requestR[185] ||
	      requestR[184] ||
	      requestR[183] ||
	      requestR[182] ||
	      requestR[181] ||
	      requestR[180] ||
	      requestR_BIT_179_71_OR_requestR_BIT_178_73_OR__ETC___d1079) &&
	     (!_64_MINUS_0_CONCAT_IF_requestR_BIT_191_27_THEN__ETC___d2955 ||
	      !_64_MINUS_0_CONCAT_IF_requestR_BIT_191_27_THEN__ETC___d2956 &&
	      !_64_MINUS_0_CONCAT_IF_requestR_BIT_191_27_THEN__ETC___d2957 &&
	      _theResult___fst_exp__h96310 == 11'd2047 &&
	      _theResult___fst_sfd__h96311 == 52'd0) ;
  assign requestR_BIT_191_27_OR_requestR_BIT_190_49_OR__ETC___d3088 =
	     (requestR[191] || requestR[190] || requestR[189] ||
	      requestR[188] ||
	      requestR[187] ||
	      requestR[186] ||
	      requestR[185] ||
	      requestR[184] ||
	      requestR[183] ||
	      requestR[182] ||
	      requestR[181] ||
	      requestR[180] ||
	      requestR_BIT_179_71_OR_requestR_BIT_178_73_OR__ETC___d1079) &&
	     _64_MINUS_0_CONCAT_IF_requestR_BIT_191_27_THEN__ETC___d2955 &&
	     _64_MINUS_0_CONCAT_IF_requestR_BIT_191_27_THEN__ETC___d2956 ;
  assign requestR_BIT_191_27_OR_requestR_BIT_190_49_OR__ETC___d3097 =
	     (requestR[191] || requestR[190] || requestR[189] ||
	      requestR[188] ||
	      requestR[187] ||
	      requestR[186] ||
	      requestR[185] ||
	      requestR[184] ||
	      requestR[183] ||
	      requestR[182] ||
	      requestR[181] ||
	      requestR[180] ||
	      requestR_BIT_179_71_OR_requestR_BIT_178_73_OR__ETC___d1079) &&
	     _64_MINUS_0_CONCAT_IF_requestR_BIT_191_27_THEN__ETC___d2955 &&
	     !_64_MINUS_0_CONCAT_IF_requestR_BIT_191_27_THEN__ETC___d2956 &&
	     IF_64_MINUS_0_CONCAT_IF_requestR_BIT_191_27_TH_ETC___d3094 ;
  assign res___1__h205637 =
	     (requestR[190:180] == 11'd2047 && requestR[179]) ?
	       64'd512 :
	       64'd256 ;
  assign res___1__h206075 = requestR[191] ? 64'd1 : 64'd128 ;
  assign res___1__h206085 = requestR[191] ? 64'd8 : 64'd16 ;
  assign res___1__h206104 = requestR[191] ? 64'd4 : 64'd32 ;
  assign res___1__h50736 =
	     (sV1_exp__h823 == 8'd255 && sV1_sfd__h824[22]) ?
	       64'd512 :
	       64'd256 ;
  assign res___1__h50972 =
	     (requestR[191:160] == 32'hFFFFFFFF && requestR[159]) ?
	       64'd1 :
	       64'd128 ;
  assign res___1__h50982 =
	     (requestR[191:160] == 32'hFFFFFFFF && requestR[159]) ?
	       64'd8 :
	       64'd16 ;
  assign res___1__h51001 =
	     (requestR[191:160] == 32'hFFFFFFFF && requestR[159]) ?
	       64'd4 :
	       64'd32 ;
  assign res__h147098 = { 32'hFFFFFFFF, x__h147104 } ;
  assign res__h188903 =
	     { IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_ETC___d5071,
	       x__h148211,
	       IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_ETC___d5035 } ;
  assign res__h193345 =
	     NOT_requestR_BITS_190_TO_180_599_EQ_2047_600_6_ETC___d5211 ?
	       requestR[191:128] :
	       requestR[127:64] ;
  assign res__h197893 =
	     NOT_requestR_BITS_190_TO_180_599_EQ_2047_600_6_ETC___d5211 ?
	       requestR[127:64] :
	       requestR[191:128] ;
  assign res__h200597 =
	     ((requestR[190:180] != 11'd2047 || requestR[179:128] == 52'd0) &&
	      (requestR[126:116] != 11'd2047 || requestR[115:64] == 52'd0) &&
	      requestR_BITS_190_TO_180_599_EQ_0_609_AND_requ_ETC___d5257) ?
	       64'd1 :
	       64'd0 ;
  assign res__h203292 =
	     NOT_requestR_BITS_190_TO_180_599_EQ_2047_600_6_ETC___d5211 ?
	       64'd1 :
	       64'd0 ;
  assign res__h205169 =
	     NOT_requestR_BITS_190_TO_180_599_EQ_2047_600_6_ETC___d5276 ?
	       64'd1 :
	       64'd0 ;
  assign res__h206120 = requestR[191] ? 64'd2 : 64'd64 ;
  assign res__h206301 = { 32'hFFFFFFFF, fpu$response_get[36:5] } ;
  assign res__h42340 =
	     { 32'hFFFFFFFF,
	       requestR_BITS_127_TO_96_2_EQ_0xFFFFFFFF_3_AND__ETC___d28 } ;
  assign res__h42577 =
	     { 32'hFFFFFFFF,
	       requestR[191:160] == 32'hFFFFFFFF && requestR[159],
	       IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d19 } ;
  assign res__h47949 =
	     NOT_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFF_ETC___d2096 ?
	       64'd1 :
	       64'd0 ;
  assign res__h49432 =
	     NOT_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFF_ETC___d2033 ?
	       64'd1 :
	       64'd0 ;
  assign res__h50501 =
	     NOT_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFF_ETC___d2114 ?
	       64'd1 :
	       64'd0 ;
  assign res__h51017 =
	     (requestR[191:160] == 32'hFFFFFFFF && requestR[159]) ?
	       64'd2 :
	       64'd64 ;
  assign result__h129694 =
	     { _0b0_CONCAT_NOT_requestR_BITS_190_TO_180_599_EQ_ETC___d3741[56:1],
	       _0b0_CONCAT_NOT_requestR_BITS_190_TO_180_599_EQ_ETC___d3741[0] |
	       guard__h129689 } ;
  assign result__h171029 =
	     { _0b0_CONCAT_NOT_IF_requestR_BITS_191_TO_160_4_E_ETC___d4573[56:1],
	       _0b0_CONCAT_NOT_IF_requestR_BITS_191_TO_160_4_E_ETC___d4573[0] |
	       guard__h171024 } ;
  assign sV1_exp__h823 =
	     (requestR[191:160] == 32'hFFFFFFFF) ?
	       requestR[158:151] :
	       8'd255 ;
  assign sV1_sfd__h824 =
	     (requestR[191:160] == 32'hFFFFFFFF) ?
	       requestR[150:128] :
	       23'd4194304 ;
  assign sV2_exp__h926 =
	     (requestR[127:96] == 32'hFFFFFFFF) ? requestR[94:87] : 8'd255 ;
  assign sV2_sfd__h927 =
	     (requestR[127:96] == 32'hFFFFFFFF) ?
	       requestR[86:64] :
	       23'd4194304 ;
  assign sfd___3__h11835 =
	     sfd__h2230 <<
	     IF_IF_requestR_BIT_191_27_THEN_NEG_requestR_BI_ETC___d384 ;
  assign sfd___3__h22457 =
	     requestR[191:128] <<
	     IF_requestR_BIT_191_27_THEN_0_ELSE_IF_requestR_ETC___d901 ;
  assign sfd___3__h28884 =
	     sfd__h23980 <<
	     IF_IF_requestR_BIT_159_6_THEN_NEG_requestR_BIT_ETC___d1252 ;
  assign sfd___3__h35055 =
	     requestR[159:128] <<
	     IF_requestR_BIT_159_6_THEN_0_ELSE_IF_requestR__ETC___d1507 ;
  assign sfd___3__h60277 =
	     sfd__h52276 <<
	     IF_IF_requestR_BIT_159_6_THEN_NEG_requestR_BIT_ETC___d2230 ;
  assign sfd___3__h69973 =
	     sfd__h62221 <<
	     IF_requestR_BIT_159_6_THEN_0_ELSE_IF_requestR__ETC___d2445 ;
  assign sfd__h103727 = { value__h72124, 3'd0 } ;
  assign sfd__h11862 = { 2'd0, sfd___3__h11835[63:41] } + 25'd1 ;
  assign sfd__h119556 =
	     { 1'b0,
	       _theResult___fst_exp__h119464 != 8'd0,
	       sfdin__h119458[56:34] } +
	     25'd1 ;
  assign sfd__h12405 =
	     { 1'b0, x__h12390[7:0] != 8'd0, sfd___3__h11835[62:40] } +
	     25'd1 ;
  assign sfd__h128168 =
	     { 1'b0,
	       _theResult___fst_exp__h128150 != 8'd0,
	       _theResult___snd__h128101[56:34] } +
	     25'd1 ;
  assign sfd__h137409 =
	     { 1'b0,
	       _theResult___fst_exp__h137317 != 8'd0,
	       sfdin__h137311[56:34] } +
	     25'd1 ;
  assign sfd__h146051 =
	     { 1'b0,
	       _theResult___fst_exp__h146032 != 8'd0,
	       _theResult___snd__h145978[56:34] } +
	     25'd1 ;
  assign sfd__h169097 =
	     { 1'b0,
	       _theResult___fst_exp__h169079 != 11'd0,
	       _theResult___snd__h169030[56:5] } +
	     54'd1 ;
  assign sfd__h178744 =
	     { 1'b0,
	       _theResult___fst_exp__h178652 != 11'd0,
	       sfdin__h178646[56:5] } +
	     54'd1 ;
  assign sfd__h187502 =
	     { 1'b0,
	       _theResult___fst_exp__h187483 != 11'd0,
	       _theResult___snd__h187429[56:5] } +
	     54'd1 ;
  assign sfd__h2230 = requestR[191] ? -requestR[191:128] : requestR[191:128] ;
  assign sfd__h22484 = { 2'd0, sfd___3__h22457[63:41] } + 25'd1 ;
  assign sfd__h23023 =
	     { 1'b0, x__h23008[7:0] != 8'd0, sfd___3__h22457[62:40] } +
	     25'd1 ;
  assign sfd__h23980 =
	     requestR[159] ? -requestR[159:128] : requestR[159:128] ;
  assign sfd__h28911 = { 2'd0, sfd___3__h28884[31:9] } + 25'd1 ;
  assign sfd__h29451 =
	     { 1'b0, x__h29436[7:0] != 8'd0, sfd___3__h28884[30:8] } + 25'd1 ;
  assign sfd__h35082 = { 2'd0, sfd___3__h35055[31:9] } + 25'd1 ;
  assign sfd__h35621 =
	     { 1'b0, x__h35606[7:0] != 8'd0, sfd___3__h35055[30:8] } + 25'd1 ;
  assign sfd__h52276 = { sfd__h23980, 23'd0 } ;
  assign sfd__h60304 = { 2'd0, sfd___3__h60277[54:3] } + 54'd1 ;
  assign sfd__h61047 =
	     { 1'b0, x__h61032[10:0] != 11'd0, sfd___3__h60277[53:2] } +
	     54'd1 ;
  assign sfd__h62221 = { requestR[159:128], 23'd0 } ;
  assign sfd__h70000 = { 2'd0, sfd___3__h69973[54:3] } + 54'd1 ;
  assign sfd__h70742 =
	     { 1'b0, x__h70727[10:0] != 11'd0, sfd___3__h69973[53:2] } +
	     54'd1 ;
  assign sfd__h83845 = { 2'd0, sfd___3__h11835[63:12] } + 54'd1 ;
  assign sfd__h84588 =
	     { 1'b0, x__h84573[10:0] != 11'd0, sfd___3__h11835[62:11] } +
	     54'd1 ;
  assign sfd__h94857 = { 2'd0, sfd___3__h22457[63:12] } + 54'd1 ;
  assign sfd__h95599 =
	     { 1'b0, x__h95584[10:0] != 11'd0, sfd___3__h22457[62:11] } +
	     54'd1 ;
  assign sfdin__h119458 =
	     _theResult____h111357[56] ?
	       _theResult___snd__h119475 :
	       _theResult___snd__h119486 ;
  assign sfdin__h137311 =
	     _theResult____h129081[56] ?
	       _theResult___snd__h137328 :
	       _theResult___snd__h137339 ;
  assign sfdin__h178646 =
	     _theResult____h170416[56] ?
	       _theResult___snd__h178663 :
	       _theResult___snd__h178674 ;
  assign value_BIT_23___h161776 = sV1_exp__h823 != 8'd0 ;
  assign value__h148270 =
	     (sV1_exp__h823 == 8'd255 && sV1_sfd__h824 != 23'd0 &&
	      !sV1_sfd__h824[22]) ?
	       _theResult___fst_sfd__h148525 :
	       sV1_sfd__h824 ;
  assign value__h36801 = { 1'b0, value_BIT_23___h161776, sV1_sfd__h824 } ;
  assign value__h72124 =
	     { 1'b0, requestR[190:180] != 11'd0, requestR[179:128] } ;
  assign value__h99566 =
	     (requestR[190:180] == 11'd2047 && requestR[179:128] != 52'd0 &&
	      !requestR[179]) ?
	       _theResult___fst_sfd__h100023 :
	       requestR[179:128] ;
  assign x__h12390 =
	     _64_MINUS_0_CONCAT_IF_IF_requestR_BIT_191_27_TH_ETC___d387 +
	     9'd127 ;
  assign x__h129789 = sfd__h103727 << x__h129822 ;
  assign x__h129822 =
	     12'd57 -
	     _3970_MINUS_SEXT_requestR_BITS_190_TO_180_599_M_ETC___d3737 ;
  assign x__h13083 =
	     { 2'd0,
	       requestR[191:128] != 64'd0 &&
	       IF_requestR_BIT_191_27_THEN_NEG_requestR_BITS__ETC___d627,
	       requestR[191:128] != 64'd0 &&
	       IF_requestR_BIT_191_27_THEN_NEG_requestR_BITS__ETC___d630,
	       requestR[191:128] != 64'd0 &&
	       IF_requestR_BIT_191_27_THEN_NEG_requestR_BITS__ETC___d639 } ;
  assign x__h13371 =
	     { 33'h1FFFFFFFE,
	       requestR_BITS_191_TO_128_24_EQ_0_25_OR_NOT_req_ETC___d837 ?
		 8'd0 :
		 _theResult___snd_fst_exp__h23540,
	       (requestR[191:128] == 64'd0 ||
		NOT_requestR_BIT_191_27_48_AND_NOT_requestR_BI_ETC___d994) ?
		 23'd0 :
		 _theResult___snd_fst_sfd__h23535 } ;
  assign x__h147104 =
	     { (requestR[190:180] == 11'd2047 && requestR[179:128] != 52'd0 ||
		(requestR[190:180] == 11'd2047 ||
		 requestR[190:180] == 11'd0) &&
		requestR[179:128] == 52'd0) ?
		 requestR[191] :
		 IF_requestR_BITS_190_TO_180_599_EQ_0_609_THEN__ETC___d4261,
	       x__h99506,
	       IF_requestR_BITS_190_TO_180_599_EQ_2047_600_AN_ETC___d4221 } ;
  assign x__h147219 =
	     { (requestR[190:180] == 11'd2047 && requestR[179:128] != 52'd0) ?
		 requestR[190:180] == 11'd2047 &&
		 requestR[179:128] != 52'd0 &&
		 !requestR[179] :
		 (requestR[190:180] != 11'd2047 ||
		  requestR[179:128] != 52'd0) &&
		 (requestR[190:180] != 11'd0 || requestR[179:128] != 52'd0) &&
		 IF_requestR_BITS_190_TO_180_599_EQ_0_609_THEN__ETC___d4312,
	       (requestR[190:180] != 11'd2047 ||
		requestR[179:128] == 52'd0) &&
	       (requestR[190:180] != 11'd2047 ||
		requestR[179:128] != 52'd0) &&
	       (requestR[190:180] != 11'd0 || requestR[179:128] != 52'd0) &&
	       IF_requestR_BITS_190_TO_180_599_EQ_0_609_THEN__ETC___d4323,
	       (requestR[190:180] != 11'd2047 ||
		requestR[179:128] == 52'd0) &&
	       (requestR[190:180] != 11'd2047 ||
		requestR[179:128] != 52'd0) &&
	       (requestR[190:180] != 11'd0 || requestR[179:128] != 52'd0) &&
	       IF_requestR_BITS_190_TO_180_599_EQ_0_609_THEN__ETC___d4339,
	       (requestR[190:180] != 11'd2047 ||
		requestR[179:128] == 52'd0) &&
	       (requestR[190:180] != 11'd2047 ||
		requestR[179:128] != 52'd0) &&
	       (requestR[190:180] != 11'd0 || requestR[179:128] != 52'd0) &&
	       IF_requestR_BITS_190_TO_180_599_EQ_0_609_THEN__ETC___d4352,
	       (requestR[190:180] != 11'd2047 ||
		requestR[179:128] == 52'd0) &&
	       (requestR[190:180] != 11'd2047 ||
		requestR[179:128] != 52'd0) &&
	       (requestR[190:180] != 11'd0 || requestR[179:128] != 52'd0) &&
	       IF_requestR_BITS_190_TO_180_599_EQ_0_609_THEN__ETC___d4365 } ;
  assign x__h148202 =
	     (x__h148211 == 11'd2047 &&
	      IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_ETC___d5035[51]) ?
	       64'h7FF8000000000000 :
	       res__h188903 ;
  assign x__h148211 =
	     (sV1_exp__h823 == 8'd255) ?
	       11'd2047 :
	       _theResult___fst_exp__h188276 ;
  assign x__h171124 = b__h39582 << x__h171157 ;
  assign x__h171157 =
	     12'd57 -
	     _3074_MINUS_SEXT_IF_requestR_BITS_191_TO_160_4__ETC___d4569 ;
  assign x__h1781 = { 32'hFFFFFFFF, x__h1787 } ;
  assign x__h1787 =
	     { requestR[127:96] == 32'hFFFFFFFF && requestR[95],
	       IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d19 } ;
  assign x__h189005 =
	     { IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_ETC___d5109,
	       (sV1_exp__h823 != 8'd255 || sV1_sfd__h824 == 23'd0) &&
	       (sV1_exp__h823 != 8'd255 || sV1_sfd__h824 != 23'd0) &&
	       (value_BIT_23___h161776 || sV1_sfd__h824 != 23'd0) &&
	       IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_ETC___d5116,
	       (sV1_exp__h823 != 8'd255 || sV1_sfd__h824 == 23'd0) &&
	       (sV1_exp__h823 != 8'd255 || sV1_sfd__h824 != 23'd0) &&
	       (value_BIT_23___h161776 || sV1_sfd__h824 != 23'd0) &&
	       IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_ETC___d5130,
	       (sV1_exp__h823 != 8'd255 || sV1_sfd__h824 == 23'd0) &&
	       (sV1_exp__h823 != 8'd255 || sV1_sfd__h824 != 23'd0) &&
	       (value_BIT_23___h161776 || sV1_sfd__h824 != 23'd0) &&
	       IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_ETC___d5142,
	       (sV1_exp__h823 != 8'd255 || sV1_sfd__h824 == 23'd0) &&
	       (sV1_exp__h823 != 8'd255 || sV1_sfd__h824 != 23'd0) &&
	       (value_BIT_23___h161776 || sV1_sfd__h824 != 23'd0) &&
	       IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_ETC___d5154 } ;
  assign x__h189928 =
	     requestR_BITS_190_TO_180_599_EQ_2047_600_AND_N_ETC___d5175 ?
	       64'h7FF8000000000000 :
	       ((requestR[190:180] == 11'd2047 &&
		 requestR[179:128] != 52'd0 &&
		 !requestR[179]) ?
		  requestR[127:64] :
		  ((requestR[126:116] == 11'd2047 &&
		    requestR[115:64] != 52'd0 &&
		    !requestR[115]) ?
		     requestR[191:128] :
		     ((requestR[190:180] == 11'd2047 && requestR[179] &&
		       requestR[126:116] == 11'd2047 &&
		       requestR[115]) ?
			64'h7FF8000000000000 :
			((requestR[190:180] == 11'd2047 && requestR[179]) ?
			   requestR[127:64] :
			   IF_requestR_BITS_126_TO_116_166_EQ_2047_167_AN_ETC___d5214)))) ;
  assign x__h1927 = { 32'hFFFFFFFF, x__h1933 } ;
  assign x__h1933 =
	     { requestR[127:96] != 32'hFFFFFFFF || !requestR[95],
	       IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d19 } ;
  assign x__h193477 =
	     { requestR_BITS_190_TO_180_599_EQ_2047_600_AND_N_ETC___d5220,
	       4'd0 } ;
  assign x__h194476 =
	     requestR_BITS_190_TO_180_599_EQ_2047_600_AND_N_ETC___d5175 ?
	       64'h7FF8000000000000 :
	       ((requestR[190:180] == 11'd2047 &&
		 requestR[179:128] != 52'd0 &&
		 !requestR[179]) ?
		  requestR[127:64] :
		  ((requestR[126:116] == 11'd2047 &&
		    requestR[115:64] != 52'd0 &&
		    !requestR[115]) ?
		     requestR[191:128] :
		     ((requestR[190:180] == 11'd2047 && requestR[179] &&
		       requestR[126:116] == 11'd2047 &&
		       requestR[115]) ?
			64'h7FF8000000000000 :
			((requestR[190:180] == 11'd2047 && requestR[179]) ?
			   requestR[127:64] :
			   ((requestR[126:116] == 11'd2047 && requestR[115]) ?
			      requestR[191:128] :
			      IF_requestR_BITS_190_TO_180_599_EQ_0_609_AND_r_ETC___d5228))))) ;
  assign x__h198920 =
	     requestR_BITS_190_TO_180_599_EQ_2047_600_AND_N_ETC___d5242 ?
	       64'd0 :
	       res__h200597 ;
  assign x__h201615 =
	     requestR_BITS_190_TO_180_599_EQ_2047_600_AND_N_ETC___d5242 ?
	       64'd0 :
	       res__h203292 ;
  assign x__h203311 =
	     { requestR[190:180] == 11'd2047 && requestR[179:128] != 52'd0 ||
	       requestR[126:116] == 11'd2047 && requestR[115:64] != 52'd0,
	       4'd0 } ;
  assign x__h203492 =
	     requestR_BITS_190_TO_180_599_EQ_2047_600_AND_N_ETC___d5242 ?
	       64'd0 :
	       res__h205169 ;
  assign x__h205619 =
	     (requestR[190:180] == 11'd2047 && requestR[179:128] != 52'd0) ?
	       res___1__h205637 :
	       ((requestR[190:180] == 11'd2047 &&
		 requestR[179:128] == 52'd0) ?
		  res___1__h206075 :
		  IF_requestR_BITS_190_TO_180_599_EQ_0_609_AND_r_ETC___d5299) ;
  assign x__h2061 = { 32'hFFFFFFFF, x__h2067 } ;
  assign x__h206269 =
	     fpu$response_get[69] ? res__h206301 : fpu$response_get[68:5] ;
  assign x__h2067 =
	     { (requestR[191:160] == 32'hFFFFFFFF && requestR[159]) !=
	       (requestR[127:96] == 32'hFFFFFFFF && requestR[95]),
	       IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d19 } ;
  assign x__h2209 = { 32'hFFFFFFFF, x__h2215 } ;
  assign x__h2215 =
	     { requestR[191:128] != 64'd0 &&
	       (NOT_IF_requestR_BIT_191_27_THEN_NEG_requestR_B_ETC___d392 ?
		  requestR[191] :
		  IF_64_MINUS_0_CONCAT_IF_IF_requestR_BIT_191_27_ETC___d454),
	       IF_requestR_BITS_191_TO_128_24_EQ_0_25_OR_NOT__ETC___d514,
	       (requestR[191:128] == 64'd0 ||
		NOT_IF_requestR_BIT_191_27_THEN_NEG_requestR_B_ETC___d392) ?
		 23'd0 :
		 _theResult___snd_fst_sfd__h12918 } ;
  assign x__h23008 =
	     _64_MINUS_0_CONCAT_IF_requestR_BIT_191_27_THEN__ETC___d904 +
	     9'd127 ;
  assign x__h23674 =
	     { 2'd0,
	       requestR[191:128] != 64'd0 &&
	       requestR_BIT_191_27_OR_requestR_BIT_190_49_OR__ETC___d1100,
	       requestR[191:128] != 64'd0 &&
	       requestR_BIT_191_27_OR_requestR_BIT_190_49_OR__ETC___d1103,
	       requestR[191:128] != 64'd0 &&
	       requestR_BIT_191_27_OR_requestR_BIT_190_49_OR__ETC___d1112 } ;
  assign x__h23959 = { 32'hFFFFFFFF, x__h23965 } ;
  assign x__h23965 =
	     { requestR[159:128] != 32'd0 &&
	       (NOT_IF_requestR_BIT_159_6_THEN_NEG_requestR_BI_ETC___d1260 ?
		  requestR[159] :
		  IF_32_MINUS_0_CONCAT_IF_IF_requestR_BIT_159_6__ETC___d1313),
	       IF_requestR_BITS_159_TO_128_121_EQ_0_122_OR_NO_ETC___d1373,
	       (requestR[159:128] == 32'd0 ||
		NOT_IF_requestR_BIT_159_6_THEN_NEG_requestR_BI_ETC___d1260) ?
		 23'd0 :
		 _theResult___snd_fst_sfd__h29964 } ;
  assign x__h29436 =
	     _32_MINUS_0_CONCAT_IF_IF_requestR_BIT_159_6_THE_ETC___d1255 +
	     9'd127 ;
  assign x__h30129 =
	     { 2'd0,
	       requestR[159:128] != 32'd0 &&
	       IF_requestR_BIT_159_6_THEN_NEG_requestR_BITS_1_ETC___d1454,
	       requestR[159:128] != 32'd0 &&
	       IF_requestR_BIT_159_6_THEN_NEG_requestR_BITS_1_ETC___d1457,
	       requestR[159:128] != 32'd0 &&
	       IF_requestR_BIT_159_6_THEN_NEG_requestR_BITS_1_ETC___d1466 } ;
  assign x__h30414 =
	     { 33'h1FFFFFFFE,
	       IF_requestR_BITS_159_TO_128_121_EQ_0_122_OR_NO_ETC___d1596,
	       (requestR[159:128] == 32'd0 ||
		!requestR[159] &&
		NOT_requestR_BIT_158_12_13_AND_NOT_requestR_BI_ETC___d803 ||
		!_32_MINUS_0_CONCAT_IF_requestR_BIT_159_6_THEN_0_ETC___d1511 ||
		_32_MINUS_0_CONCAT_IF_requestR_BIT_159_6_THEN_0_ETC___d1512) ?
		 23'd0 :
		 _theResult___snd_fst_sfd__h36133 } ;
  assign x__h35606 =
	     _32_MINUS_0_CONCAT_IF_requestR_BIT_159_6_THEN_0_ETC___d1510 +
	     9'd127 ;
  assign x__h36272 =
	     { 2'd0,
	       NOT_requestR_BITS_159_TO_128_121_EQ_0_122_123__ETC___d1643,
	       requestR[159:128] != 32'd0 &&
	       (requestR[159] ||
		requestR_BIT_158_12_OR_requestR_BIT_157_14_OR__ETC___d1058) &&
	       _32_MINUS_0_CONCAT_IF_requestR_BIT_159_6_THEN_0_ETC___d1511 &&
	       _32_MINUS_0_CONCAT_IF_requestR_BIT_159_6_THEN_0_ETC___d1512,
	       requestR[159:128] != 32'd0 &&
	       requestR_BIT_159_6_OR_requestR_BIT_158_12_OR_r_ETC___d1654 } ;
  assign x__h36556 =
	     IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d1676 ?
	       64'h7FFFFFFFFFFFFFFF :
	       IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_ETC___d1748 ;
  assign x__h37699 =
	     IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d1689 >>
	     NEG_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFF_ETC___d1715 |
	     ~(89'h1FFFFFFFFFFFFFFFFFFFFFF >>
	       NEG_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFF_ETC___d1715) &
	     {89{IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d1689[88]}} ;
  assign x__h38337 =
	     { sV1_exp__h823 == 8'd255 && sV1_sfd__h824 != 23'd0 ||
	       sV1_exp__h823 == 8'd255 && sV1_sfd__h824 == 23'd0 ||
	       NOT_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFF_ETC___d1758,
	       3'd0,
	       (sV1_exp__h823 != 8'd255 || sV1_sfd__h824 == 23'd0) &&
	       (sV1_exp__h823 != 8'd255 || sV1_sfd__h824 != 23'd0) &&
	       (value_BIT_23___h161776 || sV1_sfd__h824 != 23'd0) &&
	       IF_NEG_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0_ETC___d1769 } ;
  assign x__h38594 =
	     IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d1676 ?
	       64'hFFFFFFFFFFFFFFFF :
	       IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d1809 ;
  assign x__h39015 =
	     { value_BIT_23___h161776, sV1_sfd__h824, 65'd0 } >>
	     NEG_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFF_ETC___d1778 ;
  assign x__h39093 =
	     { IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d1828,
	       3'd0,
	       (sV1_exp__h823 != 8'd255 || sV1_sfd__h824 == 23'd0) &&
	       (sV1_exp__h823 != 8'd255 || sV1_sfd__h824 != 23'd0) &&
	       NOT_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFF_ETC___d1821 } ;
  assign x__h39336 = { {32{x__h39339[31]}}, x__h39339 } ;
  assign x__h39339 =
	     IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d1676 ?
	       32'h7FFFFFFF :
	       IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_ETC___d1897 ;
  assign x__h40258 =
	     IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d1838 >>
	     NEG_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFF_ETC___d1864 |
	     ~(57'h1FFFFFFFFFFFFFF >>
	       NEG_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFF_ETC___d1864) &
	     {57{IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d1838[56]}} ;
  assign x__h40655 =
	     { sV1_exp__h823 == 8'd255 && sV1_sfd__h824 != 23'd0 ||
	       sV1_exp__h823 == 8'd255 && sV1_sfd__h824 == 23'd0 ||
	       NOT_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFF_ETC___d1905,
	       3'd0,
	       (sV1_exp__h823 != 8'd255 || sV1_sfd__h824 == 23'd0) &&
	       (sV1_exp__h823 != 8'd255 || sV1_sfd__h824 != 23'd0) &&
	       (value_BIT_23___h161776 || sV1_sfd__h824 != 23'd0) &&
	       IF_NEG_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0_ETC___d1913 } ;
  assign x__h40912 = { {32{x__h40915[31]}}, x__h40915 } ;
  assign x__h40915 =
	     IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d1676 ?
	       32'hFFFFFFFF :
	       IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d1953 ;
  assign x__h41336 =
	     { value_BIT_23___h161776, sV1_sfd__h824, 33'd0 } >>
	     NEG_SEXT_IF_requestR_BITS_191_TO_160_4_EQ_0xFF_ETC___d1922 ;
  assign x__h41414 =
	     { IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d1973,
	       3'd0,
	       (sV1_exp__h823 != 8'd255 || sV1_sfd__h824 == 23'd0) &&
	       (sV1_exp__h823 != 8'd255 || sV1_sfd__h824 != 23'd0) &&
	       NOT_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFF_ETC___d1966 } ;
  assign x__h41662 =
	     IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d1995 ?
	       64'hFFFFFFFF7FC00000 :
	       IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_ETC___d2041 ;
  assign x__h43701 =
	     { IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d2043,
	       4'd0 } ;
  assign x__h44296 =
	     IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d1995 ?
	       64'hFFFFFFFF7FC00000 :
	       IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_ETC___d2057 ;
  assign x__h46821 = { 32'hFFFFFFFF, requestR[159:128] } ;
  assign x__h46942 =
	     { {32{requestR_BITS_159_TO_128__q1[31]}},
	       requestR_BITS_159_TO_128__q1 } ;
  assign x__h47080 =
	     IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d2080 ?
	       64'd0 :
	       res__h47949 ;
  assign x__h48563 =
	     IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d2080 ?
	       64'd0 :
	       res__h49432 ;
  assign x__h49451 =
	     { sV1_exp__h823 == 8'd255 && sV1_sfd__h824 != 23'd0 ||
	       sV2_exp__h926 == 8'd255 && sV2_sfd__h927 != 23'd0,
	       4'd0 } ;
  assign x__h49632 =
	     IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_5__ETC___d2080 ?
	       64'd0 :
	       res__h50501 ;
  assign x__h50718 =
	     (sV1_exp__h823 == 8'd255 && sV1_sfd__h824 != 23'd0) ?
	       res___1__h50736 :
	       IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFFFFFFFF_ETC___d2128 ;
  assign x__h51885 = { requestR[127], requestR[190:128] } ;
  assign x__h52007 = { !requestR[127], requestR[190:128] } ;
  assign x__h52131 = { requestR[191] != requestR[127], requestR[190:128] } ;
  assign x__h52261 =
	     { requestR[159:128] != 32'd0 &&
	       IF_NOT_32_MINUS_0_CONCAT_IF_IF_requestR_BIT_15_ETC___d2290,
	       (requestR[159:128] == 32'd0) ?
		 11'd0 :
		 _theResult___snd_fst_exp__h61768,
	       IF_requestR_BITS_159_TO_128_121_EQ_0_122_OR_NO_ETC___d2387 } ;
  assign x__h61032 =
	     _32_MINUS_0_CONCAT_IF_IF_requestR_BIT_159_6_THE_ETC___d2233 +
	     12'd1023 ;
  assign x__h61924 =
	     { 2'd0,
	       requestR[159:128] != 32'd0 &&
	       (!_32_MINUS_0_CONCAT_IF_IF_requestR_BIT_159_6_THE_ETC___d2234 ||
		!_32_MINUS_0_CONCAT_IF_IF_requestR_BIT_159_6_THE_ETC___d2236 &&
		!_32_MINUS_0_CONCAT_IF_IF_requestR_BIT_159_6_THE_ETC___d2238 &&
		_theResult___fst_exp__h61759 == 11'd2047 &&
		_theResult___fst_sfd__h61760 == 52'd0),
	       requestR[159:128] != 32'd0 &&
	       _32_MINUS_0_CONCAT_IF_IF_requestR_BIT_159_6_THE_ETC___d2234 &&
	       _32_MINUS_0_CONCAT_IF_IF_requestR_BIT_159_6_THE_ETC___d2236,
	       requestR[159:128] != 32'd0 &&
	       _32_MINUS_0_CONCAT_IF_IF_requestR_BIT_159_6_THE_ETC___d2234 &&
	       !_32_MINUS_0_CONCAT_IF_IF_requestR_BIT_159_6_THE_ETC___d2236 &&
	       IF_32_MINUS_0_CONCAT_IF_IF_requestR_BIT_159_6__ETC___d2404 } ;
  assign x__h62209 =
	     { 1'd0,
	       (requestR[159:128] == 32'd0) ?
		 11'd0 :
		 _theResult___snd_fst_exp__h71462,
	       IF_requestR_BITS_159_TO_128_121_EQ_0_122_OR_NO_ETC___d2570 } ;
  assign x__h70727 =
	     _32_MINUS_0_CONCAT_IF_requestR_BIT_159_6_THEN_0_ETC___d2448 +
	     12'd1023 ;
  assign x__h71592 =
	     { 2'd0,
	       requestR[159:128] != 32'd0 &&
	       (!_32_MINUS_0_CONCAT_IF_requestR_BIT_159_6_THEN_0_ETC___d2449 ||
		!_32_MINUS_0_CONCAT_IF_requestR_BIT_159_6_THEN_0_ETC___d2450 &&
		!_32_MINUS_0_CONCAT_IF_requestR_BIT_159_6_THEN_0_ETC___d2451 &&
		_theResult___fst_exp__h71453 == 11'd2047 &&
		_theResult___fst_sfd__h71454 == 52'd0),
	       requestR[159:128] != 32'd0 &&
	       _32_MINUS_0_CONCAT_IF_requestR_BIT_159_6_THEN_0_ETC___d2449 &&
	       _32_MINUS_0_CONCAT_IF_requestR_BIT_159_6_THEN_0_ETC___d2450,
	       requestR[159:128] != 32'd0 &&
	       _32_MINUS_0_CONCAT_IF_requestR_BIT_159_6_THEN_0_ETC___d2449 &&
	       !_32_MINUS_0_CONCAT_IF_requestR_BIT_159_6_THEN_0_ETC___d2450 &&
	       IF_32_MINUS_0_CONCAT_IF_requestR_BIT_159_6_THE_ETC___d2587 } ;
  assign x__h71876 = { {32{x__h71879[31]}}, x__h71879 } ;
  assign x__h71879 =
	     (requestR[190:180] == 11'd2047 && requestR[179:128] != 52'd0 ||
	      !requestR[191] && requestR[190:180] == 11'd2047 &&
	      requestR[179:128] == 52'd0) ?
	       32'h7FFFFFFF :
	       IF_requestR_BITS_190_TO_180_599_EQ_2047_600_AN_ETC___d2679 ;
  assign x__h72798 =
	     IF_requestR_BIT_191_27_THEN_NEG_0b0_CONCAT_NOT_ETC___d2620 >>
	     NEG_SEXT_requestR_BITS_190_TO_180_599_MINUS_10_ETC___d2646 |
	     ~(86'h3FFFFFFFFFFFFFFFFFFFFF >>
	       NEG_SEXT_requestR_BITS_190_TO_180_599_MINUS_10_ETC___d2646) &
	     {86{IF_requestR_BIT_191_27_THEN_NEG_0b0_CONCAT_NOT_ETC___d2620[85]}} ;
  assign x__h73195 =
	     { requestR[190:180] == 11'd2047 && requestR[179:128] != 52'd0 ||
	       requestR[190:180] == 11'd2047 && requestR[179:128] == 52'd0 ||
	       NOT_requestR_BITS_190_TO_180_599_EQ_0_609_615__ETC___d2690,
	       3'd0,
	       (requestR[190:180] != 11'd2047 ||
		requestR[179:128] == 52'd0) &&
	       (requestR[190:180] != 11'd2047 ||
		requestR[179:128] != 52'd0) &&
	       (requestR[190:180] != 11'd0 || requestR[179:128] != 52'd0) &&
	       IF_NEG_SEXT_requestR_BITS_190_TO_180_599_MINUS_ETC___d2701 } ;
  assign x__h73452 = { {32{x__h73455[31]}}, x__h73455 } ;
  assign x__h73455 =
	     (requestR[190:180] == 11'd2047 && requestR[179:128] != 52'd0 ||
	      !requestR[191] && requestR[190:180] == 11'd2047 &&
	      requestR[179:128] == 52'd0) ?
	       32'hFFFFFFFF :
	       (requestR[191] ?
		  32'd0 :
		  ((requestR[190:180] == 11'd2047 &&
		    requestR[179:128] == 52'd0) ?
		     32'hFFFFFFFF :
		     IF_requestR_BITS_190_TO_180_599_EQ_0_609_AND_r_ETC___d2739)) ;
  assign x__h73876 =
	     { requestR[190:180] != 11'd0, requestR[179:128], 33'd0 } >>
	     NEG_SEXT_requestR_BITS_190_TO_180_599_MINUS_10_ETC___d2710 ;
  assign x__h73954 =
	     { requestR[191] ?
		 requestR_BITS_190_TO_180_599_EQ_2047_600_AND_0_ETC___d2760 :
		 requestR_BITS_190_TO_180_599_EQ_2047_600_AND_0_ETC___d2749,
	       3'd0,
	       (requestR[190:180] != 11'd2047 ||
		requestR[179:128] == 52'd0) &&
	       (requestR[190:180] != 11'd2047 ||
		requestR[179:128] != 52'd0) &&
	       NOT_requestR_BITS_190_TO_180_599_EQ_0_609_615__ETC___d2754 } ;
  assign x__h74198 =
	     { requestR[191:128] != 64'd0 &&
	       (NOT_IF_requestR_BIT_191_27_THEN_NEG_requestR_B_ETC___d2774 ?
		  requestR[191] :
		  IF_64_MINUS_0_CONCAT_IF_IF_requestR_BIT_191_27_ETC___d2824),
	       IF_requestR_BITS_191_TO_128_24_EQ_0_25_OR_NOT__ETC___d2883,
	       (requestR[191:128] == 64'd0 ||
		NOT_IF_requestR_BIT_191_27_THEN_NEG_requestR_B_ETC___d2774) ?
		 52'd0 :
		 _theResult___snd_fst_sfd__h85304 } ;
  assign x__h84573 =
	     _64_MINUS_0_CONCAT_IF_IF_requestR_BIT_191_27_TH_ETC___d2769 +
	     12'd1023 ;
  assign x__h85465 =
	     { 2'd0,
	       requestR[191:128] != 64'd0 &&
	       IF_requestR_BIT_191_27_THEN_NEG_requestR_BITS__ETC___d2932,
	       requestR[191:128] != 64'd0 &&
	       IF_requestR_BIT_191_27_THEN_NEG_requestR_BITS__ETC___d2935,
	       requestR[191:128] != 64'd0 &&
	       IF_requestR_BIT_191_27_THEN_NEG_requestR_BITS__ETC___d2944 } ;
  assign x__h85750 =
	     { 1'd0,
	       requestR_BITS_191_TO_128_24_EQ_0_25_OR_NOT_req_ETC___d837 ?
		 11'd0 :
		 _theResult___snd_fst_exp__h96319,
	       (requestR[191:128] == 64'd0 ||
		NOT_requestR_BIT_191_27_48_AND_NOT_requestR_BI_ETC___d3042) ?
		 52'd0 :
		 _theResult___snd_fst_sfd__h96314 } ;
  assign x__h95584 =
	     _64_MINUS_0_CONCAT_IF_requestR_BIT_191_27_THEN__ETC___d2954 +
	     12'd1023 ;
  assign x__h96449 =
	     { 2'd0,
	       requestR[191:128] != 64'd0 &&
	       requestR_BIT_191_27_OR_requestR_BIT_190_49_OR__ETC___d3085,
	       requestR[191:128] != 64'd0 &&
	       requestR_BIT_191_27_OR_requestR_BIT_190_49_OR__ETC___d3088,
	       requestR[191:128] != 64'd0 &&
	       requestR_BIT_191_27_OR_requestR_BIT_190_49_OR__ETC___d3097 } ;
  assign x__h96733 =
	     (requestR[190:180] == 11'd2047 && requestR[179:128] != 52'd0 ||
	      !requestR[191] && requestR[190:180] == 11'd2047 &&
	      requestR[179:128] == 52'd0) ?
	       64'h7FFFFFFFFFFFFFFF :
	       IF_requestR_BITS_190_TO_180_599_EQ_2047_600_AN_ETC___d3168 ;
  assign x__h97876 =
	     IF_requestR_BIT_191_27_THEN_NEG_0b0_CONCAT_NOT_ETC___d3109 >>
	     NEG_SEXT_requestR_BITS_190_TO_180_599_MINUS_10_ETC___d3135 |
	     ~(118'h3FFFFFFFFFFFFFFFFFFFFFFFFFFFFF >>
	       NEG_SEXT_requestR_BITS_190_TO_180_599_MINUS_10_ETC___d3135) &
	     {118{IF_requestR_BIT_191_27_THEN_NEG_0b0_CONCAT_NOT_ETC___d3109[117]}} ;
  assign x__h98497 =
	     { requestR[190:180] == 11'd2047 && requestR[179:128] != 52'd0 ||
	       requestR[190:180] == 11'd2047 && requestR[179:128] == 52'd0 ||
	       NOT_requestR_BITS_190_TO_180_599_EQ_0_609_615__ETC___d3175,
	       3'd0,
	       (requestR[190:180] != 11'd2047 ||
		requestR[179:128] == 52'd0) &&
	       (requestR[190:180] != 11'd2047 ||
		requestR[179:128] != 52'd0) &&
	       (requestR[190:180] != 11'd0 || requestR[179:128] != 52'd0) &&
	       IF_NEG_SEXT_requestR_BITS_190_TO_180_599_MINUS_ETC___d3183 } ;
  assign x__h98754 =
	     (requestR[190:180] == 11'd2047 && requestR[179:128] != 52'd0 ||
	      !requestR[191] && requestR[190:180] == 11'd2047 &&
	      requestR[179:128] == 52'd0) ?
	       64'hFFFFFFFFFFFFFFFF :
	       (requestR[191] ?
		  64'd0 :
		  ((requestR[190:180] == 11'd2047 &&
		    requestR[179:128] == 52'd0) ?
		     64'hFFFFFFFFFFFFFFFF :
		     IF_requestR_BITS_190_TO_180_599_EQ_0_609_AND_r_ETC___d3221)) ;
  assign x__h99175 =
	     { requestR[190:180] != 11'd0, requestR[179:128], 65'd0 } >>
	     NEG_SEXT_requestR_BITS_190_TO_180_599_MINUS_10_ETC___d3192 ;
  assign x__h99253 =
	     { requestR[191] ?
		 requestR_BITS_190_TO_180_599_EQ_2047_600_AND_0_ETC___d3241 :
		 requestR_BITS_190_TO_180_599_EQ_2047_600_AND_0_ETC___d3230,
	       3'd0,
	       (requestR[190:180] != 11'd2047 ||
		requestR[179:128] == 52'd0) &&
	       (requestR[190:180] != 11'd2047 ||
		requestR[179:128] != 52'd0) &&
	       NOT_requestR_BITS_190_TO_180_599_EQ_0_609_615__ETC___d3235 } ;
  assign x__h99497 =
	     (x__h99506 == 8'd255 &&
	      IF_requestR_BITS_190_TO_180_599_EQ_2047_600_AN_ETC___d4221[22]) ?
	       64'hFFFFFFFF7FC00000 :
	       res__h147098 ;
  assign x__h99506 =
	     (requestR[190:180] == 11'd2047) ?
	       8'd255 :
	       _theResult___fst_exp__h146622 ;
  always@(requestR)
  begin
    case (requestR[194:192])
      3'h1: CASE_requestR_BITS_194_TO_192_0x1_254_0x2_IF_r_ETC__q2 = 8'd254;
      3'h2:
	  CASE_requestR_BITS_194_TO_192_0x1_254_0x2_IF_r_ETC__q2 =
	      requestR[191] ? 8'd255 : 8'd254;
      3'h3:
	  CASE_requestR_BITS_194_TO_192_0x1_254_0x2_IF_r_ETC__q2 =
	      requestR[191] ? 8'd254 : 8'd255;
      default: CASE_requestR_BITS_194_TO_192_0x1_254_0x2_IF_r_ETC__q2 = 8'd0;
    endcase
  end
  always@(requestR)
  begin
    case (requestR[194:192])
      3'h1:
	  CASE_requestR_BITS_194_TO_192_0x1_8388607_0x2__ETC__q3 =
	      23'd8388607;
      3'h2:
	  CASE_requestR_BITS_194_TO_192_0x1_8388607_0x2__ETC__q3 =
	      requestR[191] ? 23'd0 : 23'd8388607;
      3'h3:
	  CASE_requestR_BITS_194_TO_192_0x1_8388607_0x2__ETC__q3 =
	      requestR[191] ? 23'd8388607 : 23'd0;
      default: CASE_requestR_BITS_194_TO_192_0x1_8388607_0x2__ETC__q3 = 23'd0;
    endcase
  end
  always@(requestR)
  begin
    case (requestR[194:192])
      3'h1: CASE_requestR_BITS_194_TO_192_0x1_2046_0x2_IF__ETC__q4 = 11'd2046;
      3'h2:
	  CASE_requestR_BITS_194_TO_192_0x1_2046_0x2_IF__ETC__q4 =
	      (requestR[191:160] == 32'hFFFFFFFF && requestR[159]) ?
		11'd2047 :
		11'd2046;
      3'h3:
	  CASE_requestR_BITS_194_TO_192_0x1_2046_0x2_IF__ETC__q4 =
	      (requestR[191:160] == 32'hFFFFFFFF && requestR[159]) ?
		11'd2046 :
		11'd2047;
      default: CASE_requestR_BITS_194_TO_192_0x1_2046_0x2_IF__ETC__q4 = 11'd0;
    endcase
  end
  always@(requestR)
  begin
    case (requestR[194:192])
      3'h1:
	  CASE_requestR_BITS_194_TO_192_0x1_450359962737_ETC__q5 =
	      52'hFFFFFFFFFFFFF;
      3'h2:
	  CASE_requestR_BITS_194_TO_192_0x1_450359962737_ETC__q5 =
	      (requestR[191:160] == 32'hFFFFFFFF && requestR[159]) ?
		52'd0 :
		52'hFFFFFFFFFFFFF;
      3'h3:
	  CASE_requestR_BITS_194_TO_192_0x1_450359962737_ETC__q5 =
	      (requestR[191:160] == 32'hFFFFFFFF && requestR[159]) ?
		52'hFFFFFFFFFFFFF :
		52'd0;
      default: CASE_requestR_BITS_194_TO_192_0x1_450359962737_ETC__q5 = 52'd0;
    endcase
  end
  always@(requestR)
  begin
    case (requestR[194:192])
      3'h0:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x0_1_THEN_re_ETC___d40 =
	      requestR[194:192];
      3'h1: IF_requestR_BITS_194_TO_192_0_EQ_0x0_1_THEN_re_ETC___d40 = 3'd4;
      3'h2: IF_requestR_BITS_194_TO_192_0_EQ_0x0_1_THEN_re_ETC___d40 = 3'd3;
      3'h3: IF_requestR_BITS_194_TO_192_0_EQ_0x0_1_THEN_re_ETC___d40 = 3'd2;
      3'h4: IF_requestR_BITS_194_TO_192_0_EQ_0x0_1_THEN_re_ETC___d40 = 3'd1;
      default: IF_requestR_BITS_194_TO_192_0_EQ_0x0_1_THEN_re_ETC___d40 =
		   3'd0;
    endcase
  end
  always@(guard__h11845 or requestR)
  begin
    case (guard__h11845)
      2'b0, 2'b01, 2'b10:
	  CASE_guard1845_0b0_requestR_BIT_191_0b1_reques_ETC__q10 =
	      requestR[191];
      2'd3:
	  CASE_guard1845_0b0_requestR_BIT_191_0b1_reques_ETC__q10 =
	      guard__h11845 == 2'b11 && requestR[191];
    endcase
  end
  always@(requestR or guard__h11845)
  begin
    case (requestR[194:192])
      3'h2, 3'h3:
	  CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q11 =
	      requestR[191];
      3'h4:
	  CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q11 =
	      (guard__h11845 == 2'b0) ?
		requestR[191] :
		(guard__h11845 == 2'b01 || guard__h11845 == 2'b10 ||
		 guard__h11845 == 2'b11) &&
		requestR[191];
      default: CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q11 =
		   requestR[194:192] == 3'h1 && requestR[191];
    endcase
  end
  always@(guard__h12375 or requestR)
  begin
    case (guard__h12375)
      2'b0, 2'b01, 2'b10:
	  CASE_guard2375_0b0_requestR_BIT_191_0b1_reques_ETC__q12 =
	      requestR[191];
      2'd3:
	  CASE_guard2375_0b0_requestR_BIT_191_0b1_reques_ETC__q12 =
	      guard__h12375 == 2'b11 && requestR[191];
    endcase
  end
  always@(requestR or guard__h12375)
  begin
    case (requestR[194:192])
      3'h2, 3'h3:
	  CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q13 =
	      requestR[191];
      3'h4:
	  CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q13 =
	      (guard__h12375 == 2'b0) ?
		requestR[191] :
		(guard__h12375 == 2'b01 || guard__h12375 == 2'b10 ||
		 guard__h12375 == 2'b11) &&
		requestR[191];
      default: CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q13 =
		   requestR[194:192] == 3'h1 && requestR[191];
    endcase
  end
  always@(guard__h11845 or _theResult___exp__h12261)
  begin
    case (guard__h11845)
      2'b0: CASE_guard1845_0b0_0_0b1_theResult___exp2261_0_ETC__q14 = 8'd0;
      2'b01, 2'b10, 2'b11:
	  CASE_guard1845_0b0_0_0b1_theResult___exp2261_0_ETC__q14 =
	      _theResult___exp__h12261;
    endcase
  end
  always@(requestR or
	  IF_IF_IF_requestR_BIT_191_27_THEN_NEG_requestR_ETC___d476 or
	  guard__h11845 or
	  _theResult___exp__h12261 or
	  CASE_guard1845_0b0_0_0b1_theResult___exp2261_0_ETC__q14)
  begin
    case (requestR[194:192])
      3'h2:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d479 =
	      IF_IF_IF_requestR_BIT_191_27_THEN_NEG_requestR_ETC___d476;
      3'h3:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d479 =
	      (guard__h11845 == 2'b0 || requestR[191]) ?
		8'd0 :
		_theResult___exp__h12261;
      3'h4:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d479 =
	      CASE_guard1845_0b0_0_0b1_theResult___exp2261_0_ETC__q14;
      default: IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d479 =
		   8'd0;
    endcase
  end
  always@(guard__h11845 or out_exp__h12264 or _theResult___exp__h12261)
  begin
    case (guard__h11845)
      2'b0, 2'b01:
	  CASE_guard1845_0b0_0_0b1_0_0b10_out_exp2264_0b_ETC__q15 = 8'd0;
      2'b10:
	  CASE_guard1845_0b0_0_0b1_0_0b10_out_exp2264_0b_ETC__q15 =
	      out_exp__h12264;
      2'b11:
	  CASE_guard1845_0b0_0_0b1_0_0b10_out_exp2264_0b_ETC__q15 =
	      _theResult___exp__h12261;
    endcase
  end
  always@(guard__h12375 or x__h12390 or _theResult___exp__h12814)
  begin
    case (guard__h12375)
      2'b0:
	  CASE_guard2375_0b0_x2390_BITS_7_TO_0_0b1_theRe_ETC__q16 =
	      x__h12390[7:0];
      2'b01, 2'b10, 2'b11:
	  CASE_guard2375_0b0_x2390_BITS_7_TO_0_0b1_theRe_ETC__q16 =
	      _theResult___exp__h12814;
    endcase
  end
  always@(requestR or
	  x__h12390 or
	  IF_IF_IF_requestR_BIT_191_27_THEN_NEG_requestR_ETC___d504 or
	  IF_IF_IF_requestR_BIT_191_27_THEN_NEG_requestR_ETC___d502 or
	  CASE_guard2375_0b0_x2390_BITS_7_TO_0_0b1_theRe_ETC__q16)
  begin
    case (requestR[194:192])
      3'h1:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d508 =
	      x__h12390[7:0];
      3'h2:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d508 =
	      IF_IF_IF_requestR_BIT_191_27_THEN_NEG_requestR_ETC___d504;
      3'h3:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d508 =
	      IF_IF_IF_requestR_BIT_191_27_THEN_NEG_requestR_ETC___d502;
      3'h4:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d508 =
	      CASE_guard2375_0b0_x2390_BITS_7_TO_0_0b1_theRe_ETC__q16;
      default: IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d508 =
		   8'd0;
    endcase
  end
  always@(guard__h12375 or
	  x__h12390 or out_exp__h12817 or _theResult___exp__h12814)
  begin
    case (guard__h12375)
      2'b0, 2'b01:
	  CASE_guard2375_0b0_x2390_BITS_7_TO_0_0b1_x2390_ETC__q17 =
	      x__h12390[7:0];
      2'b10:
	  CASE_guard2375_0b0_x2390_BITS_7_TO_0_0b1_x2390_ETC__q17 =
	      out_exp__h12817;
      2'b11:
	  CASE_guard2375_0b0_x2390_BITS_7_TO_0_0b1_x2390_ETC__q17 =
	      _theResult___exp__h12814;
    endcase
  end
  always@(guard__h11845 or sfd___3__h11835 or _theResult___sfd__h12262)
  begin
    case (guard__h11845)
      2'b0:
	  CASE_guard1845_0b0_sfd___31835_BITS_63_TO_41_0_ETC__q18 =
	      sfd___3__h11835[63:41];
      2'b01, 2'b10, 2'b11:
	  CASE_guard1845_0b0_sfd___31835_BITS_63_TO_41_0_ETC__q18 =
	      _theResult___sfd__h12262;
    endcase
  end
  always@(requestR or
	  sfd___3__h11835 or
	  IF_IF_IF_requestR_BIT_191_27_THEN_NEG_requestR_ETC___d527 or
	  IF_IF_IF_requestR_BIT_191_27_THEN_NEG_requestR_ETC___d525 or
	  CASE_guard1845_0b0_sfd___31835_BITS_63_TO_41_0_ETC__q18)
  begin
    case (requestR[194:192])
      3'h1:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d531 =
	      sfd___3__h11835[63:41];
      3'h2:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d531 =
	      IF_IF_IF_requestR_BIT_191_27_THEN_NEG_requestR_ETC___d527;
      3'h3:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d531 =
	      IF_IF_IF_requestR_BIT_191_27_THEN_NEG_requestR_ETC___d525;
      3'h4:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d531 =
	      CASE_guard1845_0b0_sfd___31835_BITS_63_TO_41_0_ETC__q18;
      default: IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d531 =
		   23'd0;
    endcase
  end
  always@(guard__h11845 or
	  sfd___3__h11835 or out_sfd__h12265 or _theResult___sfd__h12262)
  begin
    case (guard__h11845)
      2'b0, 2'b01:
	  CASE_guard1845_0b0_sfd___31835_BITS_63_TO_41_0_ETC__q19 =
	      sfd___3__h11835[63:41];
      2'b10:
	  CASE_guard1845_0b0_sfd___31835_BITS_63_TO_41_0_ETC__q19 =
	      out_sfd__h12265;
      2'b11:
	  CASE_guard1845_0b0_sfd___31835_BITS_63_TO_41_0_ETC__q19 =
	      _theResult___sfd__h12262;
    endcase
  end
  always@(guard__h12375 or sfd___3__h11835 or _theResult___sfd__h12815)
  begin
    case (guard__h12375)
      2'b0:
	  CASE_guard2375_0b0_sfd___31835_BITS_62_TO_40_0_ETC__q20 =
	      sfd___3__h11835[62:40];
      2'b01, 2'b10, 2'b11:
	  CASE_guard2375_0b0_sfd___31835_BITS_62_TO_40_0_ETC__q20 =
	      _theResult___sfd__h12815;
    endcase
  end
  always@(requestR or
	  sfd___3__h11835 or
	  IF_IF_IF_requestR_BIT_191_27_THEN_NEG_requestR_ETC___d545 or
	  IF_IF_IF_requestR_BIT_191_27_THEN_NEG_requestR_ETC___d543 or
	  CASE_guard2375_0b0_sfd___31835_BITS_62_TO_40_0_ETC__q20)
  begin
    case (requestR[194:192])
      3'h1:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d549 =
	      sfd___3__h11835[62:40];
      3'h2:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d549 =
	      IF_IF_IF_requestR_BIT_191_27_THEN_NEG_requestR_ETC___d545;
      3'h3:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d549 =
	      IF_IF_IF_requestR_BIT_191_27_THEN_NEG_requestR_ETC___d543;
      3'h4:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d549 =
	      CASE_guard2375_0b0_sfd___31835_BITS_62_TO_40_0_ETC__q20;
      default: IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d549 =
		   23'd0;
    endcase
  end
  always@(guard__h12375 or
	  sfd___3__h11835 or out_sfd__h12818 or _theResult___sfd__h12815)
  begin
    case (guard__h12375)
      2'b0, 2'b01:
	  CASE_guard2375_0b0_sfd___31835_BITS_62_TO_40_0_ETC__q21 =
	      sfd___3__h11835[62:40];
      2'b10:
	  CASE_guard2375_0b0_sfd___31835_BITS_62_TO_40_0_ETC__q21 =
	      out_sfd__h12818;
      2'b11:
	  CASE_guard2375_0b0_sfd___31835_BITS_62_TO_40_0_ETC__q21 =
	      _theResult___sfd__h12815;
    endcase
  end
  always@(guard__h22467 or out_exp__h22883 or _theResult___exp__h22880)
  begin
    case (guard__h22467)
      2'b0, 2'b01:
	  CASE_guard2467_0b0_0_0b1_0_0b10_out_exp2883_0b_ETC__q26 = 8'd0;
      2'b10:
	  CASE_guard2467_0b0_0_0b1_0_0b10_out_exp2883_0b_ETC__q26 =
	      out_exp__h22883;
      2'b11:
	  CASE_guard2467_0b0_0_0b1_0_0b10_out_exp2883_0b_ETC__q26 =
	      _theResult___exp__h22880;
    endcase
  end
  always@(guard__h22467 or _theResult___exp__h22880)
  begin
    case (guard__h22467)
      2'b0: CASE_guard2467_0b0_0_0b1_theResult___exp2880_0_ETC__q27 = 8'd0;
      2'b01, 2'b10, 2'b11:
	  CASE_guard2467_0b0_0_0b1_theResult___exp2880_0_ETC__q27 =
	      _theResult___exp__h22880;
    endcase
  end
  always@(requestR or
	  guard__h22467 or
	  _theResult___exp__h22880 or
	  CASE_guard2467_0b0_0_0b1_theResult___exp2880_0_ETC__q27)
  begin
    case (requestR[194:192])
      3'h3:
	  CASE_requestR_BITS_194_TO_192_0x3_IF_guard2467_ETC__q28 =
	      (guard__h22467 == 2'b0) ? 8'd0 : _theResult___exp__h22880;
      3'h4:
	  CASE_requestR_BITS_194_TO_192_0x3_IF_guard2467_ETC__q28 =
	      CASE_guard2467_0b0_0_0b1_theResult___exp2880_0_ETC__q27;
      default: CASE_requestR_BITS_194_TO_192_0x3_IF_guard2467_ETC__q28 = 8'd0;
    endcase
  end
  always@(guard__h94840 or out_exp__h95459 or _theResult___exp__h95456)
  begin
    case (guard__h94840)
      2'b0, 2'b01:
	  CASE_guard4840_0b0_0_0b1_0_0b10_out_exp5459_0b_ETC__q29 = 11'd0;
      2'b10:
	  CASE_guard4840_0b0_0_0b1_0_0b10_out_exp5459_0b_ETC__q29 =
	      out_exp__h95459;
      2'b11:
	  CASE_guard4840_0b0_0_0b1_0_0b10_out_exp5459_0b_ETC__q29 =
	      _theResult___exp__h95456;
    endcase
  end
  always@(guard__h94840 or _theResult___exp__h95456)
  begin
    case (guard__h94840)
      2'b0: CASE_guard4840_0b0_0_0b1_theResult___exp5456_0_ETC__q30 = 11'd0;
      2'b01, 2'b10, 2'b11:
	  CASE_guard4840_0b0_0_0b1_theResult___exp5456_0_ETC__q30 =
	      _theResult___exp__h95456;
    endcase
  end
  always@(requestR or
	  guard__h94840 or
	  _theResult___exp__h95456 or
	  CASE_guard4840_0b0_0_0b1_theResult___exp5456_0_ETC__q30)
  begin
    case (requestR[194:192])
      3'h3:
	  CASE_requestR_BITS_194_TO_192_0x3_IF_guard4840_ETC__q31 =
	      (guard__h94840 == 2'b0) ? 11'd0 : _theResult___exp__h95456;
      3'h4:
	  CASE_requestR_BITS_194_TO_192_0x3_IF_guard4840_ETC__q31 =
	      CASE_guard4840_0b0_0_0b1_theResult___exp5456_0_ETC__q30;
      default: CASE_requestR_BITS_194_TO_192_0x3_IF_guard4840_ETC__q31 =
		   11'd0;
    endcase
  end
  always@(guard__h22993 or x__h23008 or _theResult___exp__h23432)
  begin
    case (guard__h22993)
      2'b0:
	  CASE_guard2993_0b0_x3008_BITS_7_TO_0_0b1_theRe_ETC__q32 =
	      x__h23008[7:0];
      2'b01, 2'b10, 2'b11:
	  CASE_guard2993_0b0_x3008_BITS_7_TO_0_0b1_theRe_ETC__q32 =
	      _theResult___exp__h23432;
    endcase
  end
  always@(requestR or
	  x__h23008 or
	  guard__h22993 or
	  _theResult___exp__h23432 or
	  CASE_guard2993_0b0_x3008_BITS_7_TO_0_0b1_theRe_ETC__q32)
  begin
    case (requestR[194:192])
      3'h1, 3'h2:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d985 =
	      x__h23008[7:0];
      3'h3:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d985 =
	      (guard__h22993 == 2'b0) ?
		x__h23008[7:0] :
		_theResult___exp__h23432;
      3'h4:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d985 =
	      CASE_guard2993_0b0_x3008_BITS_7_TO_0_0b1_theRe_ETC__q32;
      default: IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d985 =
		   8'd0;
    endcase
  end
  always@(guard__h22993 or
	  x__h23008 or out_exp__h23435 or _theResult___exp__h23432)
  begin
    case (guard__h22993)
      2'b0, 2'b01:
	  CASE_guard2993_0b0_x3008_BITS_7_TO_0_0b1_x3008_ETC__q33 =
	      x__h23008[7:0];
      2'b10:
	  CASE_guard2993_0b0_x3008_BITS_7_TO_0_0b1_x3008_ETC__q33 =
	      out_exp__h23435;
      2'b11:
	  CASE_guard2993_0b0_x3008_BITS_7_TO_0_0b1_x3008_ETC__q33 =
	      _theResult___exp__h23432;
    endcase
  end
  always@(guard__h22993 or sfd___3__h22457 or _theResult___sfd__h23433)
  begin
    case (guard__h22993)
      2'b0:
	  CASE_guard2993_0b0_sfd___32457_BITS_62_TO_40_0_ETC__q34 =
	      sfd___3__h22457[62:40];
      2'b01, 2'b10, 2'b11:
	  CASE_guard2993_0b0_sfd___32457_BITS_62_TO_40_0_ETC__q34 =
	      _theResult___sfd__h23433;
    endcase
  end
  always@(requestR or
	  sfd___3__h22457 or
	  guard__h22993 or
	  _theResult___sfd__h23433 or
	  CASE_guard2993_0b0_sfd___32457_BITS_62_TO_40_0_ETC__q34)
  begin
    case (requestR[194:192])
      3'h1, 3'h2:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d1023 =
	      sfd___3__h22457[62:40];
      3'h3:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d1023 =
	      (guard__h22993 == 2'b0) ?
		sfd___3__h22457[62:40] :
		_theResult___sfd__h23433;
      3'h4:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d1023 =
	      CASE_guard2993_0b0_sfd___32457_BITS_62_TO_40_0_ETC__q34;
      default: IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d1023 =
		   23'd0;
    endcase
  end
  always@(guard__h22993 or
	  sfd___3__h22457 or out_sfd__h23436 or _theResult___sfd__h23433)
  begin
    case (guard__h22993)
      2'b0, 2'b01:
	  CASE_guard2993_0b0_sfd___32457_BITS_62_TO_40_0_ETC__q35 =
	      sfd___3__h22457[62:40];
      2'b10:
	  CASE_guard2993_0b0_sfd___32457_BITS_62_TO_40_0_ETC__q35 =
	      out_sfd__h23436;
      2'b11:
	  CASE_guard2993_0b0_sfd___32457_BITS_62_TO_40_0_ETC__q35 =
	      _theResult___sfd__h23433;
    endcase
  end
  always@(guard__h22467 or sfd___3__h22457 or _theResult___sfd__h22881)
  begin
    case (guard__h22467)
      2'b0:
	  CASE_guard2467_0b0_sfd___32457_BITS_63_TO_41_0_ETC__q36 =
	      sfd___3__h22457[63:41];
      2'b01, 2'b10, 2'b11:
	  CASE_guard2467_0b0_sfd___32457_BITS_63_TO_41_0_ETC__q36 =
	      _theResult___sfd__h22881;
    endcase
  end
  always@(requestR or
	  sfd___3__h22457 or
	  guard__h22467 or
	  _theResult___sfd__h22881 or
	  CASE_guard2467_0b0_sfd___32457_BITS_63_TO_41_0_ETC__q36)
  begin
    case (requestR[194:192])
      3'h1, 3'h2:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d1008 =
	      sfd___3__h22457[63:41];
      3'h3:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d1008 =
	      (guard__h22467 == 2'b0) ?
		sfd___3__h22457[63:41] :
		_theResult___sfd__h22881;
      3'h4:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d1008 =
	      CASE_guard2467_0b0_sfd___32457_BITS_63_TO_41_0_ETC__q36;
      default: IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d1008 =
		   23'd0;
    endcase
  end
  always@(guard__h22467 or
	  sfd___3__h22457 or out_sfd__h22884 or _theResult___sfd__h22881)
  begin
    case (guard__h22467)
      2'b0, 2'b01:
	  CASE_guard2467_0b0_sfd___32457_BITS_63_TO_41_0_ETC__q37 =
	      sfd___3__h22457[63:41];
      2'b10:
	  CASE_guard2467_0b0_sfd___32457_BITS_63_TO_41_0_ETC__q37 =
	      out_sfd__h22884;
      2'b11:
	  CASE_guard2467_0b0_sfd___32457_BITS_63_TO_41_0_ETC__q37 =
	      _theResult___sfd__h22881;
    endcase
  end
  always@(guard__h28894 or requestR)
  begin
    case (guard__h28894)
      2'b0, 2'b01, 2'b10:
	  CASE_guard8894_0b0_requestR_BIT_159_0b1_reques_ETC__q40 =
	      requestR[159];
      2'd3:
	  CASE_guard8894_0b0_requestR_BIT_159_0b1_reques_ETC__q40 =
	      guard__h28894 == 2'b11 && requestR[159];
    endcase
  end
  always@(requestR or guard__h28894)
  begin
    case (requestR[194:192])
      3'h2, 3'h3:
	  CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q41 =
	      requestR[159];
      3'h4:
	  CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q41 =
	      (guard__h28894 == 2'b0) ?
		requestR[159] :
		(guard__h28894 == 2'b01 || guard__h28894 == 2'b10 ||
		 guard__h28894 == 2'b11) &&
		requestR[159];
      default: CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q41 =
		   requestR[194:192] == 3'h1 && requestR[159];
    endcase
  end
  always@(guard__h29421 or requestR)
  begin
    case (guard__h29421)
      2'b0, 2'b01, 2'b10:
	  CASE_guard9421_0b0_requestR_BIT_159_0b1_reques_ETC__q42 =
	      requestR[159];
      2'd3:
	  CASE_guard9421_0b0_requestR_BIT_159_0b1_reques_ETC__q42 =
	      guard__h29421 == 2'b11 && requestR[159];
    endcase
  end
  always@(requestR or guard__h29421)
  begin
    case (requestR[194:192])
      3'h2, 3'h3:
	  CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q43 =
	      requestR[159];
      3'h4:
	  CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q43 =
	      (guard__h29421 == 2'b0) ?
		requestR[159] :
		(guard__h29421 == 2'b01 || guard__h29421 == 2'b10 ||
		 guard__h29421 == 2'b11) &&
		requestR[159];
      default: CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q43 =
		   requestR[194:192] == 3'h1 && requestR[159];
    endcase
  end
  always@(guard__h28894 or _theResult___exp__h29307)
  begin
    case (guard__h28894)
      2'b0: CASE_guard8894_0b0_0_0b1_theResult___exp9307_0_ETC__q44 = 8'd0;
      2'b01, 2'b10, 2'b11:
	  CASE_guard8894_0b0_0_0b1_theResult___exp9307_0_ETC__q44 =
	      _theResult___exp__h29307;
    endcase
  end
  always@(requestR or
	  IF_IF_IF_requestR_BIT_159_6_THEN_NEG_requestR__ETC___d1335 or
	  guard__h28894 or
	  _theResult___exp__h29307 or
	  CASE_guard8894_0b0_0_0b1_theResult___exp9307_0_ETC__q44)
  begin
    case (requestR[194:192])
      3'h2:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d1338 =
	      IF_IF_IF_requestR_BIT_159_6_THEN_NEG_requestR__ETC___d1335;
      3'h3:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d1338 =
	      (guard__h28894 == 2'b0 || requestR[159]) ?
		8'd0 :
		_theResult___exp__h29307;
      3'h4:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d1338 =
	      CASE_guard8894_0b0_0_0b1_theResult___exp9307_0_ETC__q44;
      default: IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d1338 =
		   8'd0;
    endcase
  end
  always@(guard__h28894 or out_exp__h29310 or _theResult___exp__h29307)
  begin
    case (guard__h28894)
      2'b0, 2'b01:
	  CASE_guard8894_0b0_0_0b1_0_0b10_out_exp9310_0b_ETC__q45 = 8'd0;
      2'b10:
	  CASE_guard8894_0b0_0_0b1_0_0b10_out_exp9310_0b_ETC__q45 =
	      out_exp__h29310;
      2'b11:
	  CASE_guard8894_0b0_0_0b1_0_0b10_out_exp9310_0b_ETC__q45 =
	      _theResult___exp__h29307;
    endcase
  end
  always@(guard__h29421 or x__h29436 or _theResult___exp__h29860)
  begin
    case (guard__h29421)
      2'b0:
	  CASE_guard9421_0b0_x9436_BITS_7_TO_0_0b1_theRe_ETC__q46 =
	      x__h29436[7:0];
      2'b01, 2'b10, 2'b11:
	  CASE_guard9421_0b0_x9436_BITS_7_TO_0_0b1_theRe_ETC__q46 =
	      _theResult___exp__h29860;
    endcase
  end
  always@(requestR or
	  x__h29436 or
	  IF_IF_IF_requestR_BIT_159_6_THEN_NEG_requestR__ETC___d1363 or
	  IF_IF_IF_requestR_BIT_159_6_THEN_NEG_requestR__ETC___d1361 or
	  CASE_guard9421_0b0_x9436_BITS_7_TO_0_0b1_theRe_ETC__q46)
  begin
    case (requestR[194:192])
      3'h1:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d1367 =
	      x__h29436[7:0];
      3'h2:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d1367 =
	      IF_IF_IF_requestR_BIT_159_6_THEN_NEG_requestR__ETC___d1363;
      3'h3:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d1367 =
	      IF_IF_IF_requestR_BIT_159_6_THEN_NEG_requestR__ETC___d1361;
      3'h4:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d1367 =
	      CASE_guard9421_0b0_x9436_BITS_7_TO_0_0b1_theRe_ETC__q46;
      default: IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d1367 =
		   8'd0;
    endcase
  end
  always@(guard__h29421 or
	  x__h29436 or out_exp__h29863 or _theResult___exp__h29860)
  begin
    case (guard__h29421)
      2'b0, 2'b01:
	  CASE_guard9421_0b0_x9436_BITS_7_TO_0_0b1_x9436_ETC__q47 =
	      x__h29436[7:0];
      2'b10:
	  CASE_guard9421_0b0_x9436_BITS_7_TO_0_0b1_x9436_ETC__q47 =
	      out_exp__h29863;
      2'b11:
	  CASE_guard9421_0b0_x9436_BITS_7_TO_0_0b1_x9436_ETC__q47 =
	      _theResult___exp__h29860;
    endcase
  end
  always@(guard__h28894 or sfd___3__h28884 or _theResult___sfd__h29308)
  begin
    case (guard__h28894)
      2'b0:
	  CASE_guard8894_0b0_sfd___38884_BITS_31_TO_9_0b_ETC__q48 =
	      sfd___3__h28884[31:9];
      2'b01, 2'b10, 2'b11:
	  CASE_guard8894_0b0_sfd___38884_BITS_31_TO_9_0b_ETC__q48 =
	      _theResult___sfd__h29308;
    endcase
  end
  always@(requestR or
	  sfd___3__h28884 or
	  IF_IF_IF_requestR_BIT_159_6_THEN_NEG_requestR__ETC___d1386 or
	  IF_IF_IF_requestR_BIT_159_6_THEN_NEG_requestR__ETC___d1384 or
	  CASE_guard8894_0b0_sfd___38884_BITS_31_TO_9_0b_ETC__q48)
  begin
    case (requestR[194:192])
      3'h1:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d1390 =
	      sfd___3__h28884[31:9];
      3'h2:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d1390 =
	      IF_IF_IF_requestR_BIT_159_6_THEN_NEG_requestR__ETC___d1386;
      3'h3:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d1390 =
	      IF_IF_IF_requestR_BIT_159_6_THEN_NEG_requestR__ETC___d1384;
      3'h4:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d1390 =
	      CASE_guard8894_0b0_sfd___38884_BITS_31_TO_9_0b_ETC__q48;
      default: IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d1390 =
		   23'd0;
    endcase
  end
  always@(guard__h28894 or
	  sfd___3__h28884 or out_sfd__h29311 or _theResult___sfd__h29308)
  begin
    case (guard__h28894)
      2'b0, 2'b01:
	  CASE_guard8894_0b0_sfd___38884_BITS_31_TO_9_0b_ETC__q49 =
	      sfd___3__h28884[31:9];
      2'b10:
	  CASE_guard8894_0b0_sfd___38884_BITS_31_TO_9_0b_ETC__q49 =
	      out_sfd__h29311;
      2'b11:
	  CASE_guard8894_0b0_sfd___38884_BITS_31_TO_9_0b_ETC__q49 =
	      _theResult___sfd__h29308;
    endcase
  end
  always@(guard__h29421 or sfd___3__h28884 or _theResult___sfd__h29861)
  begin
    case (guard__h29421)
      2'b0:
	  CASE_guard9421_0b0_sfd___38884_BITS_30_TO_8_0b_ETC__q50 =
	      sfd___3__h28884[30:8];
      2'b01, 2'b10, 2'b11:
	  CASE_guard9421_0b0_sfd___38884_BITS_30_TO_8_0b_ETC__q50 =
	      _theResult___sfd__h29861;
    endcase
  end
  always@(requestR or
	  sfd___3__h28884 or
	  IF_IF_IF_requestR_BIT_159_6_THEN_NEG_requestR__ETC___d1404 or
	  IF_IF_IF_requestR_BIT_159_6_THEN_NEG_requestR__ETC___d1402 or
	  CASE_guard9421_0b0_sfd___38884_BITS_30_TO_8_0b_ETC__q50)
  begin
    case (requestR[194:192])
      3'h1:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d1408 =
	      sfd___3__h28884[30:8];
      3'h2:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d1408 =
	      IF_IF_IF_requestR_BIT_159_6_THEN_NEG_requestR__ETC___d1404;
      3'h3:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d1408 =
	      IF_IF_IF_requestR_BIT_159_6_THEN_NEG_requestR__ETC___d1402;
      3'h4:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d1408 =
	      CASE_guard9421_0b0_sfd___38884_BITS_30_TO_8_0b_ETC__q50;
      default: IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d1408 =
		   23'd0;
    endcase
  end
  always@(guard__h29421 or
	  sfd___3__h28884 or out_sfd__h29864 or _theResult___sfd__h29861)
  begin
    case (guard__h29421)
      2'b0, 2'b01:
	  CASE_guard9421_0b0_sfd___38884_BITS_30_TO_8_0b_ETC__q51 =
	      sfd___3__h28884[30:8];
      2'b10:
	  CASE_guard9421_0b0_sfd___38884_BITS_30_TO_8_0b_ETC__q51 =
	      out_sfd__h29864;
      2'b11:
	  CASE_guard9421_0b0_sfd___38884_BITS_30_TO_8_0b_ETC__q51 =
	      _theResult___sfd__h29861;
    endcase
  end
  always@(guard__h35065 or out_exp__h35481 or _theResult___exp__h35478)
  begin
    case (guard__h35065)
      2'b0, 2'b01:
	  CASE_guard5065_0b0_0_0b1_0_0b10_out_exp5481_0b_ETC__q54 = 8'd0;
      2'b10:
	  CASE_guard5065_0b0_0_0b1_0_0b10_out_exp5481_0b_ETC__q54 =
	      out_exp__h35481;
      2'b11:
	  CASE_guard5065_0b0_0_0b1_0_0b10_out_exp5481_0b_ETC__q54 =
	      _theResult___exp__h35478;
    endcase
  end
  always@(guard__h35065 or _theResult___exp__h35478)
  begin
    case (guard__h35065)
      2'b0: CASE_guard5065_0b0_0_0b1_theResult___exp5478_0_ETC__q55 = 8'd0;
      2'b01, 2'b10, 2'b11:
	  CASE_guard5065_0b0_0_0b1_theResult___exp5478_0_ETC__q55 =
	      _theResult___exp__h35478;
    endcase
  end
  always@(requestR or
	  guard__h35065 or
	  _theResult___exp__h35478 or
	  CASE_guard5065_0b0_0_0b1_theResult___exp5478_0_ETC__q55)
  begin
    case (requestR[194:192])
      3'h3:
	  CASE_requestR_BITS_194_TO_192_0x3_IF_guard5065_ETC__q56 =
	      (guard__h35065 == 2'b0) ? 8'd0 : _theResult___exp__h35478;
      3'h4:
	  CASE_requestR_BITS_194_TO_192_0x3_IF_guard5065_ETC__q56 =
	      CASE_guard5065_0b0_0_0b1_theResult___exp5478_0_ETC__q55;
      default: CASE_requestR_BITS_194_TO_192_0x3_IF_guard5065_ETC__q56 = 8'd0;
    endcase
  end
  always@(guard__h35591 or x__h35606 or _theResult___exp__h36030)
  begin
    case (guard__h35591)
      2'b0:
	  CASE_guard5591_0b0_x5606_BITS_7_TO_0_0b1_theRe_ETC__q57 =
	      x__h35606[7:0];
      2'b01, 2'b10, 2'b11:
	  CASE_guard5591_0b0_x5606_BITS_7_TO_0_0b1_theRe_ETC__q57 =
	      _theResult___exp__h36030;
    endcase
  end
  always@(requestR or
	  x__h35606 or
	  guard__h35591 or
	  _theResult___exp__h36030 or
	  CASE_guard5591_0b0_x5606_BITS_7_TO_0_0b1_theRe_ETC__q57)
  begin
    case (requestR[194:192])
      3'h1, 3'h2:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d1590 =
	      x__h35606[7:0];
      3'h3:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d1590 =
	      (guard__h35591 == 2'b0) ?
		x__h35606[7:0] :
		_theResult___exp__h36030;
      3'h4:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d1590 =
	      CASE_guard5591_0b0_x5606_BITS_7_TO_0_0b1_theRe_ETC__q57;
      default: IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d1590 =
		   8'd0;
    endcase
  end
  always@(guard__h35591 or
	  x__h35606 or out_exp__h36033 or _theResult___exp__h36030)
  begin
    case (guard__h35591)
      2'b0, 2'b01:
	  CASE_guard5591_0b0_x5606_BITS_7_TO_0_0b1_x5606_ETC__q58 =
	      x__h35606[7:0];
      2'b10:
	  CASE_guard5591_0b0_x5606_BITS_7_TO_0_0b1_x5606_ETC__q58 =
	      out_exp__h36033;
      2'b11:
	  CASE_guard5591_0b0_x5606_BITS_7_TO_0_0b1_x5606_ETC__q58 =
	      _theResult___exp__h36030;
    endcase
  end
  always@(guard__h35591 or sfd___3__h35055 or _theResult___sfd__h36031)
  begin
    case (guard__h35591)
      2'b0:
	  CASE_guard5591_0b0_sfd___35055_BITS_30_TO_8_0b_ETC__q59 =
	      sfd___3__h35055[30:8];
      2'b01, 2'b10, 2'b11:
	  CASE_guard5591_0b0_sfd___35055_BITS_30_TO_8_0b_ETC__q59 =
	      _theResult___sfd__h36031;
    endcase
  end
  always@(requestR or
	  sfd___3__h35055 or
	  guard__h35591 or
	  _theResult___sfd__h36031 or
	  CASE_guard5591_0b0_sfd___35055_BITS_30_TO_8_0b_ETC__q59)
  begin
    case (requestR[194:192])
      3'h1, 3'h2:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d1628 =
	      sfd___3__h35055[30:8];
      3'h3:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d1628 =
	      (guard__h35591 == 2'b0) ?
		sfd___3__h35055[30:8] :
		_theResult___sfd__h36031;
      3'h4:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d1628 =
	      CASE_guard5591_0b0_sfd___35055_BITS_30_TO_8_0b_ETC__q59;
      default: IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d1628 =
		   23'd0;
    endcase
  end
  always@(guard__h35591 or
	  sfd___3__h35055 or out_sfd__h36034 or _theResult___sfd__h36031)
  begin
    case (guard__h35591)
      2'b0, 2'b01:
	  CASE_guard5591_0b0_sfd___35055_BITS_30_TO_8_0b_ETC__q60 =
	      sfd___3__h35055[30:8];
      2'b10:
	  CASE_guard5591_0b0_sfd___35055_BITS_30_TO_8_0b_ETC__q60 =
	      out_sfd__h36034;
      2'b11:
	  CASE_guard5591_0b0_sfd___35055_BITS_30_TO_8_0b_ETC__q60 =
	      _theResult___sfd__h36031;
    endcase
  end
  always@(guard__h35065 or sfd___3__h35055 or _theResult___sfd__h35479)
  begin
    case (guard__h35065)
      2'b0:
	  CASE_guard5065_0b0_sfd___35055_BITS_31_TO_9_0b_ETC__q61 =
	      sfd___3__h35055[31:9];
      2'b01, 2'b10, 2'b11:
	  CASE_guard5065_0b0_sfd___35055_BITS_31_TO_9_0b_ETC__q61 =
	      _theResult___sfd__h35479;
    endcase
  end
  always@(requestR or
	  sfd___3__h35055 or
	  guard__h35065 or
	  _theResult___sfd__h35479 or
	  CASE_guard5065_0b0_sfd___35055_BITS_31_TO_9_0b_ETC__q61)
  begin
    case (requestR[194:192])
      3'h1, 3'h2:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d1613 =
	      sfd___3__h35055[31:9];
      3'h3:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d1613 =
	      (guard__h35065 == 2'b0) ?
		sfd___3__h35055[31:9] :
		_theResult___sfd__h35479;
      3'h4:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d1613 =
	      CASE_guard5065_0b0_sfd___35055_BITS_31_TO_9_0b_ETC__q61;
      default: IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d1613 =
		   23'd0;
    endcase
  end
  always@(guard__h35065 or
	  sfd___3__h35055 or out_sfd__h35482 or _theResult___sfd__h35479)
  begin
    case (guard__h35065)
      2'b0, 2'b01:
	  CASE_guard5065_0b0_sfd___35055_BITS_31_TO_9_0b_ETC__q62 =
	      sfd___3__h35055[31:9];
      2'b10:
	  CASE_guard5065_0b0_sfd___35055_BITS_31_TO_9_0b_ETC__q62 =
	      out_sfd__h35482;
      2'b11:
	  CASE_guard5065_0b0_sfd___35055_BITS_31_TO_9_0b_ETC__q62 =
	      _theResult___sfd__h35479;
    endcase
  end
  always@(guard__h60287 or requestR)
  begin
    case (guard__h60287)
      2'b0, 2'b01, 2'b10:
	  CASE_guard0287_0b0_requestR_BIT_159_0b1_reques_ETC__q69 =
	      requestR[159];
      2'd3:
	  CASE_guard0287_0b0_requestR_BIT_159_0b1_reques_ETC__q69 =
	      guard__h60287 == 2'b11 && requestR[159];
    endcase
  end
  always@(requestR or guard__h60287)
  begin
    case (requestR[194:192])
      3'h2, 3'h3:
	  CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q70 =
	      requestR[159];
      3'h4:
	  CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q70 =
	      (guard__h60287 == 2'b0) ?
		requestR[159] :
		(guard__h60287 == 2'b01 || guard__h60287 == 2'b10 ||
		 guard__h60287 == 2'b11) &&
		requestR[159];
      default: CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q70 =
		   requestR[194:192] == 3'h1 && requestR[159];
    endcase
  end
  always@(guard__h61017 or requestR)
  begin
    case (guard__h61017)
      2'b0, 2'b01, 2'b10:
	  CASE_guard1017_0b0_requestR_BIT_159_0b1_reques_ETC__q71 =
	      requestR[159];
      2'd3:
	  CASE_guard1017_0b0_requestR_BIT_159_0b1_reques_ETC__q71 =
	      guard__h61017 == 2'b11 && requestR[159];
    endcase
  end
  always@(requestR or guard__h61017)
  begin
    case (requestR[194:192])
      3'h2, 3'h3:
	  CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q72 =
	      requestR[159];
      3'h4:
	  CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q72 =
	      (guard__h61017 == 2'b0) ?
		requestR[159] :
		(guard__h61017 == 2'b01 || guard__h61017 == 2'b10 ||
		 guard__h61017 == 2'b11) &&
		requestR[159];
      default: CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q72 =
		   requestR[194:192] == 3'h1 && requestR[159];
    endcase
  end
  always@(guard__h61017 or x__h61032 or _theResult___exp__h61659)
  begin
    case (guard__h61017)
      2'b0:
	  CASE_guard1017_0b0_x1032_BITS_10_TO_0_0b1_theR_ETC__q73 =
	      x__h61032[10:0];
      2'b01, 2'b10, 2'b11:
	  CASE_guard1017_0b0_x1032_BITS_10_TO_0_0b1_theR_ETC__q73 =
	      _theResult___exp__h61659;
    endcase
  end
  always@(requestR or
	  x__h61032 or
	  IF_IF_IF_requestR_BIT_159_6_THEN_NEG_requestR__ETC___d2338 or
	  IF_IF_IF_requestR_BIT_159_6_THEN_NEG_requestR__ETC___d2336 or
	  CASE_guard1017_0b0_x1032_BITS_10_TO_0_0b1_theR_ETC__q73)
  begin
    case (requestR[194:192])
      3'h1:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d2342 =
	      x__h61032[10:0];
      3'h2:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d2342 =
	      IF_IF_IF_requestR_BIT_159_6_THEN_NEG_requestR__ETC___d2338;
      3'h3:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d2342 =
	      IF_IF_IF_requestR_BIT_159_6_THEN_NEG_requestR__ETC___d2336;
      3'h4:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d2342 =
	      CASE_guard1017_0b0_x1032_BITS_10_TO_0_0b1_theR_ETC__q73;
      default: IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d2342 =
		   11'd0;
    endcase
  end
  always@(guard__h61017 or
	  x__h61032 or out_exp__h61662 or _theResult___exp__h61659)
  begin
    case (guard__h61017)
      2'b0, 2'b01:
	  CASE_guard1017_0b0_x1032_BITS_10_TO_0_0b1_x103_ETC__q74 =
	      x__h61032[10:0];
      2'b10:
	  CASE_guard1017_0b0_x1032_BITS_10_TO_0_0b1_x103_ETC__q74 =
	      out_exp__h61662;
      2'b11:
	  CASE_guard1017_0b0_x1032_BITS_10_TO_0_0b1_x103_ETC__q74 =
	      _theResult___exp__h61659;
    endcase
  end
  always@(guard__h61017 or sfd___3__h60277 or _theResult___sfd__h61660)
  begin
    case (guard__h61017)
      2'b0:
	  CASE_guard1017_0b0_sfd___30277_BITS_53_TO_2_0b_ETC__q75 =
	      sfd___3__h60277[53:2];
      2'b01, 2'b10, 2'b11:
	  CASE_guard1017_0b0_sfd___30277_BITS_53_TO_2_0b_ETC__q75 =
	      _theResult___sfd__h61660;
    endcase
  end
  always@(requestR or
	  sfd___3__h60277 or
	  IF_IF_IF_requestR_BIT_159_6_THEN_NEG_requestR__ETC___d2379 or
	  IF_IF_IF_requestR_BIT_159_6_THEN_NEG_requestR__ETC___d2377 or
	  CASE_guard1017_0b0_sfd___30277_BITS_53_TO_2_0b_ETC__q75)
  begin
    case (requestR[194:192])
      3'h1:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d2383 =
	      sfd___3__h60277[53:2];
      3'h2:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d2383 =
	      IF_IF_IF_requestR_BIT_159_6_THEN_NEG_requestR__ETC___d2379;
      3'h3:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d2383 =
	      IF_IF_IF_requestR_BIT_159_6_THEN_NEG_requestR__ETC___d2377;
      3'h4:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d2383 =
	      CASE_guard1017_0b0_sfd___30277_BITS_53_TO_2_0b_ETC__q75;
      default: IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d2383 =
		   52'd0;
    endcase
  end
  always@(guard__h61017 or
	  sfd___3__h60277 or out_sfd__h61663 or _theResult___sfd__h61660)
  begin
    case (guard__h61017)
      2'b0, 2'b01:
	  CASE_guard1017_0b0_sfd___30277_BITS_53_TO_2_0b_ETC__q76 =
	      sfd___3__h60277[53:2];
      2'b10:
	  CASE_guard1017_0b0_sfd___30277_BITS_53_TO_2_0b_ETC__q76 =
	      out_sfd__h61663;
      2'b11:
	  CASE_guard1017_0b0_sfd___30277_BITS_53_TO_2_0b_ETC__q76 =
	      _theResult___sfd__h61660;
    endcase
  end
  always@(guard__h60287 or _theResult___exp__h60903)
  begin
    case (guard__h60287)
      2'b0: CASE_guard0287_0b0_0_0b1_theResult___exp0903_0_ETC__q77 = 11'd0;
      2'b01, 2'b10, 2'b11:
	  CASE_guard0287_0b0_0_0b1_theResult___exp0903_0_ETC__q77 =
	      _theResult___exp__h60903;
    endcase
  end
  always@(requestR or
	  IF_IF_IF_requestR_BIT_159_6_THEN_NEG_requestR__ETC___d2310 or
	  guard__h60287 or
	  _theResult___exp__h60903 or
	  CASE_guard0287_0b0_0_0b1_theResult___exp0903_0_ETC__q77)
  begin
    case (requestR[194:192])
      3'h2:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d2313 =
	      IF_IF_IF_requestR_BIT_159_6_THEN_NEG_requestR__ETC___d2310;
      3'h3:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d2313 =
	      (guard__h60287 == 2'b0 || requestR[159]) ?
		11'd0 :
		_theResult___exp__h60903;
      3'h4:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d2313 =
	      CASE_guard0287_0b0_0_0b1_theResult___exp0903_0_ETC__q77;
      default: IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d2313 =
		   11'd0;
    endcase
  end
  always@(guard__h60287 or out_exp__h60906 or _theResult___exp__h60903)
  begin
    case (guard__h60287)
      2'b0, 2'b01:
	  CASE_guard0287_0b0_0_0b1_0_0b10_out_exp0906_0b_ETC__q78 = 11'd0;
      2'b10:
	  CASE_guard0287_0b0_0_0b1_0_0b10_out_exp0906_0b_ETC__q78 =
	      out_exp__h60906;
      2'b11:
	  CASE_guard0287_0b0_0_0b1_0_0b10_out_exp0906_0b_ETC__q78 =
	      _theResult___exp__h60903;
    endcase
  end
  always@(guard__h60287 or sfd___3__h60277 or _theResult___sfd__h60904)
  begin
    case (guard__h60287)
      2'b0:
	  CASE_guard0287_0b0_sfd___30277_BITS_54_TO_3_0b_ETC__q79 =
	      sfd___3__h60277[54:3];
      2'b01, 2'b10, 2'b11:
	  CASE_guard0287_0b0_sfd___30277_BITS_54_TO_3_0b_ETC__q79 =
	      _theResult___sfd__h60904;
    endcase
  end
  always@(requestR or
	  sfd___3__h60277 or
	  IF_IF_IF_requestR_BIT_159_6_THEN_NEG_requestR__ETC___d2361 or
	  IF_IF_IF_requestR_BIT_159_6_THEN_NEG_requestR__ETC___d2359 or
	  CASE_guard0287_0b0_sfd___30277_BITS_54_TO_3_0b_ETC__q79)
  begin
    case (requestR[194:192])
      3'h1:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d2365 =
	      sfd___3__h60277[54:3];
      3'h2:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d2365 =
	      IF_IF_IF_requestR_BIT_159_6_THEN_NEG_requestR__ETC___d2361;
      3'h3:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d2365 =
	      IF_IF_IF_requestR_BIT_159_6_THEN_NEG_requestR__ETC___d2359;
      3'h4:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d2365 =
	      CASE_guard0287_0b0_sfd___30277_BITS_54_TO_3_0b_ETC__q79;
      default: IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d2365 =
		   52'd0;
    endcase
  end
  always@(guard__h60287 or
	  sfd___3__h60277 or out_sfd__h60907 or _theResult___sfd__h60904)
  begin
    case (guard__h60287)
      2'b0, 2'b01:
	  CASE_guard0287_0b0_sfd___30277_BITS_54_TO_3_0b_ETC__q80 =
	      sfd___3__h60277[54:3];
      2'b10:
	  CASE_guard0287_0b0_sfd___30277_BITS_54_TO_3_0b_ETC__q80 =
	      out_sfd__h60907;
      2'b11:
	  CASE_guard0287_0b0_sfd___30277_BITS_54_TO_3_0b_ETC__q80 =
	      _theResult___sfd__h60904;
    endcase
  end
  always@(guard__h69983 or out_exp__h70602 or _theResult___exp__h70599)
  begin
    case (guard__h69983)
      2'b0, 2'b01:
	  CASE_guard9983_0b0_0_0b1_0_0b10_out_exp0602_0b_ETC__q83 = 11'd0;
      2'b10:
	  CASE_guard9983_0b0_0_0b1_0_0b10_out_exp0602_0b_ETC__q83 =
	      out_exp__h70602;
      2'b11:
	  CASE_guard9983_0b0_0_0b1_0_0b10_out_exp0602_0b_ETC__q83 =
	      _theResult___exp__h70599;
    endcase
  end
  always@(guard__h69983 or _theResult___exp__h70599)
  begin
    case (guard__h69983)
      2'b0: CASE_guard9983_0b0_0_0b1_theResult___exp0599_0_ETC__q84 = 11'd0;
      2'b01, 2'b10, 2'b11:
	  CASE_guard9983_0b0_0_0b1_theResult___exp0599_0_ETC__q84 =
	      _theResult___exp__h70599;
    endcase
  end
  always@(requestR or
	  guard__h69983 or
	  _theResult___exp__h70599 or
	  CASE_guard9983_0b0_0_0b1_theResult___exp0599_0_ETC__q84)
  begin
    case (requestR[194:192])
      3'h3:
	  CASE_requestR_BITS_194_TO_192_0x3_IF_guard9983_ETC__q85 =
	      (guard__h69983 == 2'b0) ? 11'd0 : _theResult___exp__h70599;
      3'h4:
	  CASE_requestR_BITS_194_TO_192_0x3_IF_guard9983_ETC__q85 =
	      CASE_guard9983_0b0_0_0b1_theResult___exp0599_0_ETC__q84;
      default: CASE_requestR_BITS_194_TO_192_0x3_IF_guard9983_ETC__q85 =
		   11'd0;
    endcase
  end
  always@(guard__h70712 or x__h70727 or _theResult___exp__h71354)
  begin
    case (guard__h70712)
      2'b0:
	  CASE_guard0712_0b0_x0727_BITS_10_TO_0_0b1_theR_ETC__q86 =
	      x__h70727[10:0];
      2'b01, 2'b10, 2'b11:
	  CASE_guard0712_0b0_x0727_BITS_10_TO_0_0b1_theR_ETC__q86 =
	      _theResult___exp__h71354;
    endcase
  end
  always@(requestR or
	  x__h70727 or
	  guard__h70712 or
	  _theResult___exp__h71354 or
	  CASE_guard0712_0b0_x0727_BITS_10_TO_0_0b1_theR_ETC__q86)
  begin
    case (requestR[194:192])
      3'h1, 3'h2:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d2529 =
	      x__h70727[10:0];
      3'h3:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d2529 =
	      (guard__h70712 == 2'b0) ?
		x__h70727[10:0] :
		_theResult___exp__h71354;
      3'h4:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d2529 =
	      CASE_guard0712_0b0_x0727_BITS_10_TO_0_0b1_theR_ETC__q86;
      default: IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d2529 =
		   11'd0;
    endcase
  end
  always@(guard__h70712 or
	  x__h70727 or out_exp__h71357 or _theResult___exp__h71354)
  begin
    case (guard__h70712)
      2'b0, 2'b01:
	  CASE_guard0712_0b0_x0727_BITS_10_TO_0_0b1_x072_ETC__q87 =
	      x__h70727[10:0];
      2'b10:
	  CASE_guard0712_0b0_x0727_BITS_10_TO_0_0b1_x072_ETC__q87 =
	      out_exp__h71357;
      2'b11:
	  CASE_guard0712_0b0_x0727_BITS_10_TO_0_0b1_x072_ETC__q87 =
	      _theResult___exp__h71354;
    endcase
  end
  always@(guard__h70712 or sfd___3__h69973 or _theResult___sfd__h71355)
  begin
    case (guard__h70712)
      2'b0:
	  CASE_guard0712_0b0_sfd___39973_BITS_53_TO_2_0b_ETC__q88 =
	      sfd___3__h69973[53:2];
      2'b01, 2'b10, 2'b11:
	  CASE_guard0712_0b0_sfd___39973_BITS_53_TO_2_0b_ETC__q88 =
	      _theResult___sfd__h71355;
    endcase
  end
  always@(requestR or
	  sfd___3__h69973 or
	  guard__h70712 or
	  _theResult___sfd__h71355 or
	  CASE_guard0712_0b0_sfd___39973_BITS_53_TO_2_0b_ETC__q88)
  begin
    case (requestR[194:192])
      3'h1, 3'h2:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d2566 =
	      sfd___3__h69973[53:2];
      3'h3:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d2566 =
	      (guard__h70712 == 2'b0) ?
		sfd___3__h69973[53:2] :
		_theResult___sfd__h71355;
      3'h4:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d2566 =
	      CASE_guard0712_0b0_sfd___39973_BITS_53_TO_2_0b_ETC__q88;
      default: IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d2566 =
		   52'd0;
    endcase
  end
  always@(guard__h70712 or
	  sfd___3__h69973 or out_sfd__h71358 or _theResult___sfd__h71355)
  begin
    case (guard__h70712)
      2'b0, 2'b01:
	  CASE_guard0712_0b0_sfd___39973_BITS_53_TO_2_0b_ETC__q89 =
	      sfd___3__h69973[53:2];
      2'b10:
	  CASE_guard0712_0b0_sfd___39973_BITS_53_TO_2_0b_ETC__q89 =
	      out_sfd__h71358;
      2'b11:
	  CASE_guard0712_0b0_sfd___39973_BITS_53_TO_2_0b_ETC__q89 =
	      _theResult___sfd__h71355;
    endcase
  end
  always@(guard__h69983 or sfd___3__h69973 or _theResult___sfd__h70600)
  begin
    case (guard__h69983)
      2'b0:
	  CASE_guard9983_0b0_sfd___39973_BITS_54_TO_3_0b_ETC__q90 =
	      sfd___3__h69973[54:3];
      2'b01, 2'b10, 2'b11:
	  CASE_guard9983_0b0_sfd___39973_BITS_54_TO_3_0b_ETC__q90 =
	      _theResult___sfd__h70600;
    endcase
  end
  always@(requestR or
	  sfd___3__h69973 or
	  guard__h69983 or
	  _theResult___sfd__h70600 or
	  CASE_guard9983_0b0_sfd___39973_BITS_54_TO_3_0b_ETC__q90)
  begin
    case (requestR[194:192])
      3'h1, 3'h2:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d2551 =
	      sfd___3__h69973[54:3];
      3'h3:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d2551 =
	      (guard__h69983 == 2'b0) ?
		sfd___3__h69973[54:3] :
		_theResult___sfd__h70600;
      3'h4:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d2551 =
	      CASE_guard9983_0b0_sfd___39973_BITS_54_TO_3_0b_ETC__q90;
      default: IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d2551 =
		   52'd0;
    endcase
  end
  always@(guard__h69983 or
	  sfd___3__h69973 or out_sfd__h70603 or _theResult___sfd__h70600)
  begin
    case (guard__h69983)
      2'b0, 2'b01:
	  CASE_guard9983_0b0_sfd___39973_BITS_54_TO_3_0b_ETC__q91 =
	      sfd___3__h69973[54:3];
      2'b10:
	  CASE_guard9983_0b0_sfd___39973_BITS_54_TO_3_0b_ETC__q91 =
	      out_sfd__h70603;
      2'b11:
	  CASE_guard9983_0b0_sfd___39973_BITS_54_TO_3_0b_ETC__q91 =
	      _theResult___sfd__h70600;
    endcase
  end
  always@(guard__h83828 or requestR)
  begin
    case (guard__h83828)
      2'b0, 2'b01, 2'b10:
	  CASE_guard3828_0b0_requestR_BIT_191_0b1_reques_ETC__q94 =
	      requestR[191];
      2'd3:
	  CASE_guard3828_0b0_requestR_BIT_191_0b1_reques_ETC__q94 =
	      guard__h83828 == 2'b11 && requestR[191];
    endcase
  end
  always@(requestR or guard__h83828)
  begin
    case (requestR[194:192])
      3'h2, 3'h3:
	  CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q95 =
	      requestR[191];
      3'h4:
	  CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q95 =
	      (guard__h83828 == 2'b0) ?
		requestR[191] :
		(guard__h83828 == 2'b01 || guard__h83828 == 2'b10 ||
		 guard__h83828 == 2'b11) &&
		requestR[191];
      default: CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q95 =
		   requestR[194:192] == 3'h1 && requestR[191];
    endcase
  end
  always@(guard__h84558 or requestR)
  begin
    case (guard__h84558)
      2'b0, 2'b01, 2'b10:
	  CASE_guard4558_0b0_requestR_BIT_191_0b1_reques_ETC__q96 =
	      requestR[191];
      2'd3:
	  CASE_guard4558_0b0_requestR_BIT_191_0b1_reques_ETC__q96 =
	      guard__h84558 == 2'b11 && requestR[191];
    endcase
  end
  always@(requestR or guard__h84558)
  begin
    case (requestR[194:192])
      3'h2, 3'h3:
	  CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q97 =
	      requestR[191];
      3'h4:
	  CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q97 =
	      (guard__h84558 == 2'b0) ?
		requestR[191] :
		(guard__h84558 == 2'b01 || guard__h84558 == 2'b10 ||
		 guard__h84558 == 2'b11) &&
		requestR[191];
      default: CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q97 =
		   requestR[194:192] == 3'h1 && requestR[191];
    endcase
  end
  always@(guard__h84558 or x__h84573 or _theResult___exp__h85200)
  begin
    case (guard__h84558)
      2'b0:
	  CASE_guard4558_0b0_x4573_BITS_10_TO_0_0b1_theR_ETC__q98 =
	      x__h84573[10:0];
      2'b01, 2'b10, 2'b11:
	  CASE_guard4558_0b0_x4573_BITS_10_TO_0_0b1_theR_ETC__q98 =
	      _theResult___exp__h85200;
    endcase
  end
  always@(requestR or
	  x__h84573 or
	  IF_IF_IF_requestR_BIT_191_27_THEN_NEG_requestR_ETC___d2873 or
	  IF_IF_IF_requestR_BIT_191_27_THEN_NEG_requestR_ETC___d2871 or
	  CASE_guard4558_0b0_x4573_BITS_10_TO_0_0b1_theR_ETC__q98)
  begin
    case (requestR[194:192])
      3'h1:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d2877 =
	      x__h84573[10:0];
      3'h2:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d2877 =
	      IF_IF_IF_requestR_BIT_191_27_THEN_NEG_requestR_ETC___d2873;
      3'h3:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d2877 =
	      IF_IF_IF_requestR_BIT_191_27_THEN_NEG_requestR_ETC___d2871;
      3'h4:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d2877 =
	      CASE_guard4558_0b0_x4573_BITS_10_TO_0_0b1_theR_ETC__q98;
      default: IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d2877 =
		   11'd0;
    endcase
  end
  always@(guard__h84558 or
	  x__h84573 or out_exp__h85203 or _theResult___exp__h85200)
  begin
    case (guard__h84558)
      2'b0, 2'b01:
	  CASE_guard4558_0b0_x4573_BITS_10_TO_0_0b1_x457_ETC__q99 =
	      x__h84573[10:0];
      2'b10:
	  CASE_guard4558_0b0_x4573_BITS_10_TO_0_0b1_x457_ETC__q99 =
	      out_exp__h85203;
      2'b11:
	  CASE_guard4558_0b0_x4573_BITS_10_TO_0_0b1_x457_ETC__q99 =
	      _theResult___exp__h85200;
    endcase
  end
  always@(guard__h84558 or sfd___3__h11835 or _theResult___sfd__h85201)
  begin
    case (guard__h84558)
      2'b0:
	  CASE_guard4558_0b0_sfd___31835_BITS_62_TO_11_0_ETC__q100 =
	      sfd___3__h11835[62:11];
      2'b01, 2'b10, 2'b11:
	  CASE_guard4558_0b0_sfd___31835_BITS_62_TO_11_0_ETC__q100 =
	      _theResult___sfd__h85201;
    endcase
  end
  always@(requestR or
	  sfd___3__h11835 or
	  IF_IF_IF_requestR_BIT_191_27_THEN_NEG_requestR_ETC___d2914 or
	  IF_IF_IF_requestR_BIT_191_27_THEN_NEG_requestR_ETC___d2912 or
	  CASE_guard4558_0b0_sfd___31835_BITS_62_TO_11_0_ETC__q100)
  begin
    case (requestR[194:192])
      3'h1:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d2918 =
	      sfd___3__h11835[62:11];
      3'h2:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d2918 =
	      IF_IF_IF_requestR_BIT_191_27_THEN_NEG_requestR_ETC___d2914;
      3'h3:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d2918 =
	      IF_IF_IF_requestR_BIT_191_27_THEN_NEG_requestR_ETC___d2912;
      3'h4:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d2918 =
	      CASE_guard4558_0b0_sfd___31835_BITS_62_TO_11_0_ETC__q100;
      default: IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d2918 =
		   52'd0;
    endcase
  end
  always@(guard__h84558 or
	  sfd___3__h11835 or out_sfd__h85204 or _theResult___sfd__h85201)
  begin
    case (guard__h84558)
      2'b0, 2'b01:
	  CASE_guard4558_0b0_sfd___31835_BITS_62_TO_11_0_ETC__q101 =
	      sfd___3__h11835[62:11];
      2'b10:
	  CASE_guard4558_0b0_sfd___31835_BITS_62_TO_11_0_ETC__q101 =
	      out_sfd__h85204;
      2'b11:
	  CASE_guard4558_0b0_sfd___31835_BITS_62_TO_11_0_ETC__q101 =
	      _theResult___sfd__h85201;
    endcase
  end
  always@(guard__h83828 or _theResult___exp__h84444)
  begin
    case (guard__h83828)
      2'b0: CASE_guard3828_0b0_0_0b1_theResult___exp4444_0_ETC__q102 = 11'd0;
      2'b01, 2'b10, 2'b11:
	  CASE_guard3828_0b0_0_0b1_theResult___exp4444_0_ETC__q102 =
	      _theResult___exp__h84444;
    endcase
  end
  always@(requestR or
	  IF_IF_IF_requestR_BIT_191_27_THEN_NEG_requestR_ETC___d2845 or
	  guard__h83828 or
	  _theResult___exp__h84444 or
	  CASE_guard3828_0b0_0_0b1_theResult___exp4444_0_ETC__q102)
  begin
    case (requestR[194:192])
      3'h2:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d2848 =
	      IF_IF_IF_requestR_BIT_191_27_THEN_NEG_requestR_ETC___d2845;
      3'h3:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d2848 =
	      (guard__h83828 == 2'b0 || requestR[191]) ?
		11'd0 :
		_theResult___exp__h84444;
      3'h4:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d2848 =
	      CASE_guard3828_0b0_0_0b1_theResult___exp4444_0_ETC__q102;
      default: IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d2848 =
		   11'd0;
    endcase
  end
  always@(guard__h83828 or out_exp__h84447 or _theResult___exp__h84444)
  begin
    case (guard__h83828)
      2'b0, 2'b01:
	  CASE_guard3828_0b0_0_0b1_0_0b10_out_exp4447_0b_ETC__q103 = 11'd0;
      2'b10:
	  CASE_guard3828_0b0_0_0b1_0_0b10_out_exp4447_0b_ETC__q103 =
	      out_exp__h84447;
      2'b11:
	  CASE_guard3828_0b0_0_0b1_0_0b10_out_exp4447_0b_ETC__q103 =
	      _theResult___exp__h84444;
    endcase
  end
  always@(guard__h83828 or sfd___3__h11835 or _theResult___sfd__h84445)
  begin
    case (guard__h83828)
      2'b0:
	  CASE_guard3828_0b0_sfd___31835_BITS_63_TO_12_0_ETC__q104 =
	      sfd___3__h11835[63:12];
      2'b01, 2'b10, 2'b11:
	  CASE_guard3828_0b0_sfd___31835_BITS_63_TO_12_0_ETC__q104 =
	      _theResult___sfd__h84445;
    endcase
  end
  always@(requestR or
	  sfd___3__h11835 or
	  IF_IF_IF_requestR_BIT_191_27_THEN_NEG_requestR_ETC___d2896 or
	  IF_IF_IF_requestR_BIT_191_27_THEN_NEG_requestR_ETC___d2894 or
	  CASE_guard3828_0b0_sfd___31835_BITS_63_TO_12_0_ETC__q104)
  begin
    case (requestR[194:192])
      3'h1:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d2900 =
	      sfd___3__h11835[63:12];
      3'h2:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d2900 =
	      IF_IF_IF_requestR_BIT_191_27_THEN_NEG_requestR_ETC___d2896;
      3'h3:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d2900 =
	      IF_IF_IF_requestR_BIT_191_27_THEN_NEG_requestR_ETC___d2894;
      3'h4:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d2900 =
	      CASE_guard3828_0b0_sfd___31835_BITS_63_TO_12_0_ETC__q104;
      default: IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d2900 =
		   52'd0;
    endcase
  end
  always@(guard__h83828 or
	  sfd___3__h11835 or out_sfd__h84448 or _theResult___sfd__h84445)
  begin
    case (guard__h83828)
      2'b0, 2'b01:
	  CASE_guard3828_0b0_sfd___31835_BITS_63_TO_12_0_ETC__q105 =
	      sfd___3__h11835[63:12];
      2'b10:
	  CASE_guard3828_0b0_sfd___31835_BITS_63_TO_12_0_ETC__q105 =
	      out_sfd__h84448;
      2'b11:
	  CASE_guard3828_0b0_sfd___31835_BITS_63_TO_12_0_ETC__q105 =
	      _theResult___sfd__h84445;
    endcase
  end
  always@(guard__h95569 or x__h95584 or _theResult___exp__h96211)
  begin
    case (guard__h95569)
      2'b0:
	  CASE_guard5569_0b0_x5584_BITS_10_TO_0_0b1_theR_ETC__q106 =
	      x__h95584[10:0];
      2'b01, 2'b10, 2'b11:
	  CASE_guard5569_0b0_x5584_BITS_10_TO_0_0b1_theR_ETC__q106 =
	      _theResult___exp__h96211;
    endcase
  end
  always@(requestR or
	  x__h95584 or
	  guard__h95569 or
	  _theResult___exp__h96211 or
	  CASE_guard5569_0b0_x5584_BITS_10_TO_0_0b1_theR_ETC__q106)
  begin
    case (requestR[194:192])
      3'h1, 3'h2:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d3033 =
	      x__h95584[10:0];
      3'h3:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d3033 =
	      (guard__h95569 == 2'b0) ?
		x__h95584[10:0] :
		_theResult___exp__h96211;
      3'h4:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d3033 =
	      CASE_guard5569_0b0_x5584_BITS_10_TO_0_0b1_theR_ETC__q106;
      default: IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d3033 =
		   11'd0;
    endcase
  end
  always@(guard__h95569 or
	  x__h95584 or out_exp__h96214 or _theResult___exp__h96211)
  begin
    case (guard__h95569)
      2'b0, 2'b01:
	  CASE_guard5569_0b0_x5584_BITS_10_TO_0_0b1_x558_ETC__q107 =
	      x__h95584[10:0];
      2'b10:
	  CASE_guard5569_0b0_x5584_BITS_10_TO_0_0b1_x558_ETC__q107 =
	      out_exp__h96214;
      2'b11:
	  CASE_guard5569_0b0_x5584_BITS_10_TO_0_0b1_x558_ETC__q107 =
	      _theResult___exp__h96211;
    endcase
  end
  always@(guard__h95569 or sfd___3__h22457 or _theResult___sfd__h96212)
  begin
    case (guard__h95569)
      2'b0:
	  CASE_guard5569_0b0_sfd___32457_BITS_62_TO_11_0_ETC__q108 =
	      sfd___3__h22457[62:11];
      2'b01, 2'b10, 2'b11:
	  CASE_guard5569_0b0_sfd___32457_BITS_62_TO_11_0_ETC__q108 =
	      _theResult___sfd__h96212;
    endcase
  end
  always@(requestR or
	  sfd___3__h22457 or
	  guard__h95569 or
	  _theResult___sfd__h96212 or
	  CASE_guard5569_0b0_sfd___32457_BITS_62_TO_11_0_ETC__q108)
  begin
    case (requestR[194:192])
      3'h1, 3'h2:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d3071 =
	      sfd___3__h22457[62:11];
      3'h3:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d3071 =
	      (guard__h95569 == 2'b0) ?
		sfd___3__h22457[62:11] :
		_theResult___sfd__h96212;
      3'h4:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d3071 =
	      CASE_guard5569_0b0_sfd___32457_BITS_62_TO_11_0_ETC__q108;
      default: IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d3071 =
		   52'd0;
    endcase
  end
  always@(guard__h95569 or
	  sfd___3__h22457 or out_sfd__h96215 or _theResult___sfd__h96212)
  begin
    case (guard__h95569)
      2'b0, 2'b01:
	  CASE_guard5569_0b0_sfd___32457_BITS_62_TO_11_0_ETC__q109 =
	      sfd___3__h22457[62:11];
      2'b10:
	  CASE_guard5569_0b0_sfd___32457_BITS_62_TO_11_0_ETC__q109 =
	      out_sfd__h96215;
      2'b11:
	  CASE_guard5569_0b0_sfd___32457_BITS_62_TO_11_0_ETC__q109 =
	      _theResult___sfd__h96212;
    endcase
  end
  always@(guard__h94840 or sfd___3__h22457 or _theResult___sfd__h95457)
  begin
    case (guard__h94840)
      2'b0:
	  CASE_guard4840_0b0_sfd___32457_BITS_63_TO_12_0_ETC__q110 =
	      sfd___3__h22457[63:12];
      2'b01, 2'b10, 2'b11:
	  CASE_guard4840_0b0_sfd___32457_BITS_63_TO_12_0_ETC__q110 =
	      _theResult___sfd__h95457;
    endcase
  end
  always@(requestR or
	  sfd___3__h22457 or
	  guard__h94840 or
	  _theResult___sfd__h95457 or
	  CASE_guard4840_0b0_sfd___32457_BITS_63_TO_12_0_ETC__q110)
  begin
    case (requestR[194:192])
      3'h1, 3'h2:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d3056 =
	      sfd___3__h22457[63:12];
      3'h3:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d3056 =
	      (guard__h94840 == 2'b0) ?
		sfd___3__h22457[63:12] :
		_theResult___sfd__h95457;
      3'h4:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d3056 =
	      CASE_guard4840_0b0_sfd___32457_BITS_63_TO_12_0_ETC__q110;
      default: IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d3056 =
		   52'd0;
    endcase
  end
  always@(guard__h94840 or
	  sfd___3__h22457 or out_sfd__h95460 or _theResult___sfd__h95457)
  begin
    case (guard__h94840)
      2'b0, 2'b01:
	  CASE_guard4840_0b0_sfd___32457_BITS_63_TO_12_0_ETC__q111 =
	      sfd___3__h22457[63:12];
      2'b10:
	  CASE_guard4840_0b0_sfd___32457_BITS_63_TO_12_0_ETC__q111 =
	      out_sfd__h95460;
      2'b11:
	  CASE_guard4840_0b0_sfd___32457_BITS_63_TO_12_0_ETC__q111 =
	      _theResult___sfd__h95457;
    endcase
  end
  always@(guard__h111367 or
	  _theResult___fst_exp__h119464 or _theResult___exp__h119990)
  begin
    case (guard__h111367)
      2'b0:
	  CASE_guard11367_0b0_theResult___fst_exp19464_0_ETC__q124 =
	      _theResult___fst_exp__h119464;
      2'b01, 2'b10, 2'b11:
	  CASE_guard11367_0b0_theResult___fst_exp19464_0_ETC__q124 =
	      _theResult___exp__h119990;
    endcase
  end
  always@(requestR or
	  _theResult___fst_exp__h119464 or
	  IF_IF_IF_IF_0b0_CONCAT_NOT_requestR_BITS_190_T_ETC___d3598 or
	  IF_IF_IF_IF_0b0_CONCAT_NOT_requestR_BITS_190_T_ETC___d3596 or
	  CASE_guard11367_0b0_theResult___fst_exp19464_0_ETC__q124)
  begin
    case (requestR[194:192])
      3'h1:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d3602 =
	      _theResult___fst_exp__h119464;
      3'h2:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d3602 =
	      IF_IF_IF_IF_0b0_CONCAT_NOT_requestR_BITS_190_T_ETC___d3598;
      3'h3:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d3602 =
	      IF_IF_IF_IF_0b0_CONCAT_NOT_requestR_BITS_190_T_ETC___d3596;
      3'h4:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d3602 =
	      CASE_guard11367_0b0_theResult___fst_exp19464_0_ETC__q124;
      default: IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d3602 =
		   8'd0;
    endcase
  end
  always@(guard__h111367 or
	  _theResult___fst_exp__h119464 or
	  out_exp__h119993 or _theResult___exp__h119990)
  begin
    case (guard__h111367)
      2'b0, 2'b01:
	  CASE_guard11367_0b0_theResult___fst_exp19464_0_ETC__q125 =
	      _theResult___fst_exp__h119464;
      2'b10:
	  CASE_guard11367_0b0_theResult___fst_exp19464_0_ETC__q125 =
	      out_exp__h119993;
      2'b11:
	  CASE_guard11367_0b0_theResult___fst_exp19464_0_ETC__q125 =
	      _theResult___exp__h119990;
    endcase
  end
  always@(guard__h120102 or
	  _theResult___fst_exp__h128150 or _theResult___exp__h128602)
  begin
    case (guard__h120102)
      2'b0:
	  CASE_guard20102_0b0_theResult___fst_exp28150_0_ETC__q126 =
	      _theResult___fst_exp__h128150;
      2'b01, 2'b10, 2'b11:
	  CASE_guard20102_0b0_theResult___fst_exp28150_0_ETC__q126 =
	      _theResult___exp__h128602;
    endcase
  end
  always@(requestR or
	  _theResult___fst_exp__h128150 or
	  IF_IF_IF_requestR_BITS_190_TO_180_599_EQ_0_609_ETC___d3715 or
	  IF_IF_IF_requestR_BITS_190_TO_180_599_EQ_0_609_ETC___d3713 or
	  CASE_guard20102_0b0_theResult___fst_exp28150_0_ETC__q126)
  begin
    case (requestR[194:192])
      3'h1:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d3719 =
	      _theResult___fst_exp__h128150;
      3'h2:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d3719 =
	      IF_IF_IF_requestR_BITS_190_TO_180_599_EQ_0_609_ETC___d3715;
      3'h3:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d3719 =
	      IF_IF_IF_requestR_BITS_190_TO_180_599_EQ_0_609_ETC___d3713;
      3'h4:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d3719 =
	      CASE_guard20102_0b0_theResult___fst_exp28150_0_ETC__q126;
      default: IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d3719 =
		   8'd0;
    endcase
  end
  always@(guard__h120102 or
	  _theResult___fst_exp__h128150 or
	  out_exp__h128605 or _theResult___exp__h128602)
  begin
    case (guard__h120102)
      2'b0, 2'b01:
	  CASE_guard20102_0b0_theResult___fst_exp28150_0_ETC__q127 =
	      _theResult___fst_exp__h128150;
      2'b10:
	  CASE_guard20102_0b0_theResult___fst_exp28150_0_ETC__q127 =
	      out_exp__h128605;
      2'b11:
	  CASE_guard20102_0b0_theResult___fst_exp28150_0_ETC__q127 =
	      _theResult___exp__h128602;
    endcase
  end
  always@(guard__h129091 or
	  _theResult___fst_exp__h137317 or _theResult___exp__h137843)
  begin
    case (guard__h129091)
      2'b0:
	  CASE_guard29091_0b0_theResult___fst_exp37317_0_ETC__q128 =
	      _theResult___fst_exp__h137317;
      2'b01, 2'b10, 2'b11:
	  CASE_guard29091_0b0_theResult___fst_exp37317_0_ETC__q128 =
	      _theResult___exp__h137843;
    endcase
  end
  always@(requestR or
	  _theResult___fst_exp__h137317 or
	  IF_IF_IF_IF_3970_MINUS_SEXT_requestR_BITS_190__ETC___d4042 or
	  IF_IF_IF_IF_3970_MINUS_SEXT_requestR_BITS_190__ETC___d4040 or
	  CASE_guard29091_0b0_theResult___fst_exp37317_0_ETC__q128)
  begin
    case (requestR[194:192])
      3'h1:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d4046 =
	      _theResult___fst_exp__h137317;
      3'h2:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d4046 =
	      IF_IF_IF_IF_3970_MINUS_SEXT_requestR_BITS_190__ETC___d4042;
      3'h3:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d4046 =
	      IF_IF_IF_IF_3970_MINUS_SEXT_requestR_BITS_190__ETC___d4040;
      3'h4:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d4046 =
	      CASE_guard29091_0b0_theResult___fst_exp37317_0_ETC__q128;
      default: IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d4046 =
		   8'd0;
    endcase
  end
  always@(guard__h129091 or
	  _theResult___fst_exp__h137317 or
	  out_exp__h137846 or _theResult___exp__h137843)
  begin
    case (guard__h129091)
      2'b0, 2'b01:
	  CASE_guard29091_0b0_theResult___fst_exp37317_0_ETC__q129 =
	      _theResult___fst_exp__h137317;
      2'b10:
	  CASE_guard29091_0b0_theResult___fst_exp37317_0_ETC__q129 =
	      out_exp__h137846;
      2'b11:
	  CASE_guard29091_0b0_theResult___fst_exp37317_0_ETC__q129 =
	      _theResult___exp__h137843;
    endcase
  end
  always@(guard__h137955 or
	  _theResult___fst_exp__h146032 or _theResult___exp__h146509)
  begin
    case (guard__h137955)
      2'b0:
	  CASE_guard37955_0b0_theResult___fst_exp46032_0_ETC__q130 =
	      _theResult___fst_exp__h146032;
      2'b01, 2'b10, 2'b11:
	  CASE_guard37955_0b0_theResult___fst_exp46032_0_ETC__q130 =
	      _theResult___exp__h146509;
    endcase
  end
  always@(requestR or
	  _theResult___fst_exp__h146032 or
	  IF_IF_IF_requestR_BITS_190_TO_180_599_EQ_0_609_ETC___d4111 or
	  IF_IF_IF_requestR_BITS_190_TO_180_599_EQ_0_609_ETC___d4109 or
	  CASE_guard37955_0b0_theResult___fst_exp46032_0_ETC__q130)
  begin
    case (requestR[194:192])
      3'h1:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d4115 =
	      _theResult___fst_exp__h146032;
      3'h2:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d4115 =
	      IF_IF_IF_requestR_BITS_190_TO_180_599_EQ_0_609_ETC___d4111;
      3'h3:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d4115 =
	      IF_IF_IF_requestR_BITS_190_TO_180_599_EQ_0_609_ETC___d4109;
      3'h4:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d4115 =
	      CASE_guard37955_0b0_theResult___fst_exp46032_0_ETC__q130;
      default: IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d4115 =
		   8'd0;
    endcase
  end
  always@(guard__h137955 or
	  _theResult___fst_exp__h146032 or
	  out_exp__h146512 or _theResult___exp__h146509)
  begin
    case (guard__h137955)
      2'b0, 2'b01:
	  CASE_guard37955_0b0_theResult___fst_exp46032_0_ETC__q131 =
	      _theResult___fst_exp__h146032;
      2'b10:
	  CASE_guard37955_0b0_theResult___fst_exp46032_0_ETC__q131 =
	      out_exp__h146512;
      2'b11:
	  CASE_guard37955_0b0_theResult___fst_exp46032_0_ETC__q131 =
	      _theResult___exp__h146509;
    endcase
  end
  always@(guard__h120102 or
	  _theResult___snd__h128101 or _theResult___sfd__h128603)
  begin
    case (guard__h120102)
      2'b0:
	  CASE_guard20102_0b0_theResult___snd28101_BITS__ETC__q132 =
	      _theResult___snd__h128101[56:34];
      2'b01, 2'b10, 2'b11:
	  CASE_guard20102_0b0_theResult___snd28101_BITS__ETC__q132 =
	      _theResult___sfd__h128603;
    endcase
  end
  always@(requestR or
	  _theResult___snd__h128101 or
	  IF_IF_IF_requestR_BITS_190_TO_180_599_EQ_0_609_ETC___d4164 or
	  IF_IF_IF_requestR_BITS_190_TO_180_599_EQ_0_609_ETC___d4162 or
	  CASE_guard20102_0b0_theResult___snd28101_BITS__ETC__q132)
  begin
    case (requestR[194:192])
      3'h1:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d4168 =
	      _theResult___snd__h128101[56:34];
      3'h2:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d4168 =
	      IF_IF_IF_requestR_BITS_190_TO_180_599_EQ_0_609_ETC___d4164;
      3'h3:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d4168 =
	      IF_IF_IF_requestR_BITS_190_TO_180_599_EQ_0_609_ETC___d4162;
      3'h4:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d4168 =
	      CASE_guard20102_0b0_theResult___snd28101_BITS__ETC__q132;
      default: IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d4168 =
		   23'd0;
    endcase
  end
  always@(guard__h120102 or
	  _theResult___snd__h128101 or
	  out_sfd__h128606 or _theResult___sfd__h128603)
  begin
    case (guard__h120102)
      2'b0, 2'b01:
	  CASE_guard20102_0b0_theResult___snd28101_BITS__ETC__q133 =
	      _theResult___snd__h128101[56:34];
      2'b10:
	  CASE_guard20102_0b0_theResult___snd28101_BITS__ETC__q133 =
	      out_sfd__h128606;
      2'b11:
	  CASE_guard20102_0b0_theResult___snd28101_BITS__ETC__q133 =
	      _theResult___sfd__h128603;
    endcase
  end
  always@(guard__h111367 or sfdin__h119458 or _theResult___sfd__h119991)
  begin
    case (guard__h111367)
      2'b0:
	  CASE_guard11367_0b0_sfdin19458_BITS_56_TO_34_0_ETC__q134 =
	      sfdin__h119458[56:34];
      2'b01, 2'b10, 2'b11:
	  CASE_guard11367_0b0_sfdin19458_BITS_56_TO_34_0_ETC__q134 =
	      _theResult___sfd__h119991;
    endcase
  end
  always@(requestR or
	  sfdin__h119458 or
	  IF_IF_IF_IF_0b0_CONCAT_NOT_requestR_BITS_190_T_ETC___d4145 or
	  IF_IF_IF_IF_0b0_CONCAT_NOT_requestR_BITS_190_T_ETC___d4143 or
	  CASE_guard11367_0b0_sfdin19458_BITS_56_TO_34_0_ETC__q134)
  begin
    case (requestR[194:192])
      3'h1:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d4149 =
	      sfdin__h119458[56:34];
      3'h2:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d4149 =
	      IF_IF_IF_IF_0b0_CONCAT_NOT_requestR_BITS_190_T_ETC___d4145;
      3'h3:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d4149 =
	      IF_IF_IF_IF_0b0_CONCAT_NOT_requestR_BITS_190_T_ETC___d4143;
      3'h4:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d4149 =
	      CASE_guard11367_0b0_sfdin19458_BITS_56_TO_34_0_ETC__q134;
      default: IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d4149 =
		   23'd0;
    endcase
  end
  always@(guard__h111367 or
	  sfdin__h119458 or out_sfd__h119994 or _theResult___sfd__h119991)
  begin
    case (guard__h111367)
      2'b0, 2'b01:
	  CASE_guard11367_0b0_sfdin19458_BITS_56_TO_34_0_ETC__q135 =
	      sfdin__h119458[56:34];
      2'b10:
	  CASE_guard11367_0b0_sfdin19458_BITS_56_TO_34_0_ETC__q135 =
	      out_sfd__h119994;
      2'b11:
	  CASE_guard11367_0b0_sfdin19458_BITS_56_TO_34_0_ETC__q135 =
	      _theResult___sfd__h119991;
    endcase
  end
  always@(guard__h129091 or sfdin__h137311 or _theResult___sfd__h137844)
  begin
    case (guard__h129091)
      2'b0:
	  CASE_guard29091_0b0_sfdin37311_BITS_56_TO_34_0_ETC__q136 =
	      sfdin__h137311[56:34];
      2'b01, 2'b10, 2'b11:
	  CASE_guard29091_0b0_sfdin37311_BITS_56_TO_34_0_ETC__q136 =
	      _theResult___sfd__h137844;
    endcase
  end
  always@(requestR or
	  sfdin__h137311 or
	  IF_IF_IF_IF_3970_MINUS_SEXT_requestR_BITS_190__ETC___d4191 or
	  IF_IF_IF_IF_3970_MINUS_SEXT_requestR_BITS_190__ETC___d4189 or
	  CASE_guard29091_0b0_sfdin37311_BITS_56_TO_34_0_ETC__q136)
  begin
    case (requestR[194:192])
      3'h1:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d4195 =
	      sfdin__h137311[56:34];
      3'h2:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d4195 =
	      IF_IF_IF_IF_3970_MINUS_SEXT_requestR_BITS_190__ETC___d4191;
      3'h3:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d4195 =
	      IF_IF_IF_IF_3970_MINUS_SEXT_requestR_BITS_190__ETC___d4189;
      3'h4:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d4195 =
	      CASE_guard29091_0b0_sfdin37311_BITS_56_TO_34_0_ETC__q136;
      default: IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d4195 =
		   23'd0;
    endcase
  end
  always@(guard__h129091 or
	  sfdin__h137311 or out_sfd__h137847 or _theResult___sfd__h137844)
  begin
    case (guard__h129091)
      2'b0, 2'b01:
	  CASE_guard29091_0b0_sfdin37311_BITS_56_TO_34_0_ETC__q137 =
	      sfdin__h137311[56:34];
      2'b10:
	  CASE_guard29091_0b0_sfdin37311_BITS_56_TO_34_0_ETC__q137 =
	      out_sfd__h137847;
      2'b11:
	  CASE_guard29091_0b0_sfdin37311_BITS_56_TO_34_0_ETC__q137 =
	      _theResult___sfd__h137844;
    endcase
  end
  always@(guard__h137955 or
	  _theResult___snd__h145978 or _theResult___sfd__h146510)
  begin
    case (guard__h137955)
      2'b0:
	  CASE_guard37955_0b0_theResult___snd45978_BITS__ETC__q138 =
	      _theResult___snd__h145978[56:34];
      2'b01, 2'b10, 2'b11:
	  CASE_guard37955_0b0_theResult___snd45978_BITS__ETC__q138 =
	      _theResult___sfd__h146510;
    endcase
  end
  always@(requestR or
	  _theResult___snd__h145978 or
	  IF_IF_IF_requestR_BITS_190_TO_180_599_EQ_0_609_ETC___d4210 or
	  IF_IF_IF_requestR_BITS_190_TO_180_599_EQ_0_609_ETC___d4208 or
	  CASE_guard37955_0b0_theResult___snd45978_BITS__ETC__q138)
  begin
    case (requestR[194:192])
      3'h1:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d4214 =
	      _theResult___snd__h145978[56:34];
      3'h2:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d4214 =
	      IF_IF_IF_requestR_BITS_190_TO_180_599_EQ_0_609_ETC___d4210;
      3'h3:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d4214 =
	      IF_IF_IF_requestR_BITS_190_TO_180_599_EQ_0_609_ETC___d4208;
      3'h4:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d4214 =
	      CASE_guard37955_0b0_theResult___snd45978_BITS__ETC__q138;
      default: IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d4214 =
		   23'd0;
    endcase
  end
  always@(guard__h137955 or
	  _theResult___snd__h145978 or
	  out_sfd__h146513 or _theResult___sfd__h146510)
  begin
    case (guard__h137955)
      2'b0, 2'b01:
	  CASE_guard37955_0b0_theResult___snd45978_BITS__ETC__q139 =
	      _theResult___snd__h145978[56:34];
      2'b10:
	  CASE_guard37955_0b0_theResult___snd45978_BITS__ETC__q139 =
	      out_sfd__h146513;
      2'b11:
	  CASE_guard37955_0b0_theResult___snd45978_BITS__ETC__q139 =
	      _theResult___sfd__h146510;
    endcase
  end
  always@(guard__h111367 or requestR)
  begin
    case (guard__h111367)
      2'b0, 2'b01, 2'b10:
	  CASE_guard11367_0b0_requestR_BIT_191_0b1_reque_ETC__q140 =
	      requestR[191];
      2'd3:
	  CASE_guard11367_0b0_requestR_BIT_191_0b1_reque_ETC__q140 =
	      guard__h111367 == 2'b11 && requestR[191];
    endcase
  end
  always@(requestR or guard__h111367)
  begin
    case (requestR[194:192])
      3'h2, 3'h3:
	  CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q141 =
	      requestR[191];
      3'h4:
	  CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q141 =
	      (guard__h111367 == 2'b0) ?
		requestR[191] :
		(guard__h111367 == 2'b01 || guard__h111367 == 2'b10 ||
		 guard__h111367 == 2'b11) &&
		requestR[191];
      default: CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q141 =
		   requestR[194:192] == 3'h1 && requestR[191];
    endcase
  end
  always@(guard__h120102 or requestR)
  begin
    case (guard__h120102)
      2'b0, 2'b01, 2'b10:
	  CASE_guard20102_0b0_requestR_BIT_191_0b1_reque_ETC__q142 =
	      requestR[191];
      2'd3:
	  CASE_guard20102_0b0_requestR_BIT_191_0b1_reque_ETC__q142 =
	      guard__h120102 == 2'b11 && requestR[191];
    endcase
  end
  always@(requestR or guard__h120102)
  begin
    case (requestR[194:192])
      3'h2, 3'h3:
	  CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q143 =
	      requestR[191];
      3'h4:
	  CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q143 =
	      (guard__h120102 == 2'b0) ?
		requestR[191] :
		(guard__h120102 == 2'b01 || guard__h120102 == 2'b10 ||
		 guard__h120102 == 2'b11) &&
		requestR[191];
      default: CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q143 =
		   requestR[194:192] == 3'h1 && requestR[191];
    endcase
  end
  always@(guard__h129091 or requestR)
  begin
    case (guard__h129091)
      2'b0, 2'b01, 2'b10:
	  CASE_guard29091_0b0_requestR_BIT_191_0b1_reque_ETC__q144 =
	      requestR[191];
      2'd3:
	  CASE_guard29091_0b0_requestR_BIT_191_0b1_reque_ETC__q144 =
	      guard__h129091 == 2'b11 && requestR[191];
    endcase
  end
  always@(requestR or guard__h129091)
  begin
    case (requestR[194:192])
      3'h2, 3'h3:
	  CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q145 =
	      requestR[191];
      3'h4:
	  CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q145 =
	      (guard__h129091 == 2'b0) ?
		requestR[191] :
		(guard__h129091 == 2'b01 || guard__h129091 == 2'b10 ||
		 guard__h129091 == 2'b11) &&
		requestR[191];
      default: CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q145 =
		   requestR[194:192] == 3'h1 && requestR[191];
    endcase
  end
  always@(guard__h137955 or requestR)
  begin
    case (guard__h137955)
      2'b0, 2'b01, 2'b10:
	  CASE_guard37955_0b0_requestR_BIT_191_0b1_reque_ETC__q146 =
	      requestR[191];
      2'd3:
	  CASE_guard37955_0b0_requestR_BIT_191_0b1_reque_ETC__q146 =
	      guard__h137955 == 2'b11 && requestR[191];
    endcase
  end
  always@(requestR or guard__h137955)
  begin
    case (requestR[194:192])
      3'h2, 3'h3:
	  CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q147 =
	      requestR[191];
      3'h4:
	  CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q147 =
	      (guard__h137955 == 2'b0) ?
		requestR[191] :
		(guard__h137955 == 2'b01 || guard__h137955 == 2'b10 ||
		 guard__h137955 == 2'b11) &&
		requestR[191];
      default: CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q147 =
		   requestR[194:192] == 3'h1 && requestR[191];
    endcase
  end
  always@(guard__h161118 or
	  _theResult___fst_exp__h169079 or _theResult___exp__h169734)
  begin
    case (guard__h161118)
      2'b0:
	  CASE_guard61118_0b0_theResult___fst_exp69079_0_ETC__q156 =
	      _theResult___fst_exp__h169079;
      2'b01, 2'b10, 2'b11:
	  CASE_guard61118_0b0_theResult___fst_exp69079_0_ETC__q156 =
	      _theResult___exp__h169734;
    endcase
  end
  always@(requestR or
	  _theResult___fst_exp__h169079 or
	  IF_IF_IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFF_ETC___d4551 or
	  IF_IF_IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFF_ETC___d4549 or
	  CASE_guard61118_0b0_theResult___fst_exp69079_0_ETC__q156)
  begin
    case (requestR[194:192])
      3'h1:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d4555 =
	      _theResult___fst_exp__h169079;
      3'h2:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d4555 =
	      IF_IF_IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFF_ETC___d4551;
      3'h3:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d4555 =
	      IF_IF_IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFF_ETC___d4549;
      3'h4:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d4555 =
	      CASE_guard61118_0b0_theResult___fst_exp69079_0_ETC__q156;
      default: IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d4555 =
		   11'd0;
    endcase
  end
  always@(guard__h161118 or
	  _theResult___fst_exp__h169079 or
	  out_exp__h169737 or _theResult___exp__h169734)
  begin
    case (guard__h161118)
      2'b0, 2'b01:
	  CASE_guard61118_0b0_theResult___fst_exp69079_0_ETC__q157 =
	      _theResult___fst_exp__h169079;
      2'b10:
	  CASE_guard61118_0b0_theResult___fst_exp69079_0_ETC__q157 =
	      out_exp__h169737;
      2'b11:
	  CASE_guard61118_0b0_theResult___fst_exp69079_0_ETC__q157 =
	      _theResult___exp__h169734;
    endcase
  end
  always@(guard__h170426 or
	  _theResult___fst_exp__h178652 or _theResult___exp__h179381)
  begin
    case (guard__h170426)
      2'b0:
	  CASE_guard70426_0b0_theResult___fst_exp78652_0_ETC__q158 =
	      _theResult___fst_exp__h178652;
      2'b01, 2'b10, 2'b11:
	  CASE_guard70426_0b0_theResult___fst_exp78652_0_ETC__q158 =
	      _theResult___exp__h179381;
    endcase
  end
  always@(requestR or
	  _theResult___fst_exp__h178652 or
	  IF_IF_IF_IF_3074_MINUS_SEXT_IF_requestR_BITS_1_ETC___d4876 or
	  IF_IF_IF_IF_3074_MINUS_SEXT_IF_requestR_BITS_1_ETC___d4874 or
	  CASE_guard70426_0b0_theResult___fst_exp78652_0_ETC__q158)
  begin
    case (requestR[194:192])
      3'h1:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d4880 =
	      _theResult___fst_exp__h178652;
      3'h2:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d4880 =
	      IF_IF_IF_IF_3074_MINUS_SEXT_IF_requestR_BITS_1_ETC___d4876;
      3'h3:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d4880 =
	      IF_IF_IF_IF_3074_MINUS_SEXT_IF_requestR_BITS_1_ETC___d4874;
      3'h4:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d4880 =
	      CASE_guard70426_0b0_theResult___fst_exp78652_0_ETC__q158;
      default: IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d4880 =
		   11'd0;
    endcase
  end
  always@(guard__h170426 or
	  _theResult___fst_exp__h178652 or
	  out_exp__h179384 or _theResult___exp__h179381)
  begin
    case (guard__h170426)
      2'b0, 2'b01:
	  CASE_guard70426_0b0_theResult___fst_exp78652_0_ETC__q159 =
	      _theResult___fst_exp__h178652;
      2'b10:
	  CASE_guard70426_0b0_theResult___fst_exp78652_0_ETC__q159 =
	      out_exp__h179384;
      2'b11:
	  CASE_guard70426_0b0_theResult___fst_exp78652_0_ETC__q159 =
	      _theResult___exp__h179381;
    endcase
  end
  always@(guard__h179493 or
	  _theResult___fst_exp__h187483 or _theResult___exp__h188163)
  begin
    case (guard__h179493)
      2'b0:
	  CASE_guard79493_0b0_theResult___fst_exp87483_0_ETC__q160 =
	      _theResult___fst_exp__h187483;
      2'b01, 2'b10, 2'b11:
	  CASE_guard79493_0b0_theResult___fst_exp87483_0_ETC__q160 =
	      _theResult___exp__h188163;
    endcase
  end
  always@(requestR or
	  _theResult___fst_exp__h187483 or
	  IF_IF_IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFF_ETC___d4945 or
	  IF_IF_IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFF_ETC___d4943 or
	  CASE_guard79493_0b0_theResult___fst_exp87483_0_ETC__q160)
  begin
    case (requestR[194:192])
      3'h1:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d4949 =
	      _theResult___fst_exp__h187483;
      3'h2:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d4949 =
	      IF_IF_IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFF_ETC___d4945;
      3'h3:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d4949 =
	      IF_IF_IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFF_ETC___d4943;
      3'h4:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d4949 =
	      CASE_guard79493_0b0_theResult___fst_exp87483_0_ETC__q160;
      default: IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d4949 =
		   11'd0;
    endcase
  end
  always@(guard__h179493 or
	  _theResult___fst_exp__h187483 or
	  out_exp__h188166 or _theResult___exp__h188163)
  begin
    case (guard__h179493)
      2'b0, 2'b01:
	  CASE_guard79493_0b0_theResult___fst_exp87483_0_ETC__q161 =
	      _theResult___fst_exp__h187483;
      2'b10:
	  CASE_guard79493_0b0_theResult___fst_exp87483_0_ETC__q161 =
	      out_exp__h188166;
      2'b11:
	  CASE_guard79493_0b0_theResult___fst_exp87483_0_ETC__q161 =
	      _theResult___exp__h188163;
    endcase
  end
  always@(guard__h161118 or requestR)
  begin
    case (guard__h161118)
      2'b0, 2'b01, 2'b10:
	  CASE_guard61118_0b0_requestR_BITS_191_TO_160_E_ETC__q162 =
	      requestR[191:160] == 32'hFFFFFFFF && requestR[159];
      2'd3:
	  CASE_guard61118_0b0_requestR_BITS_191_TO_160_E_ETC__q162 =
	      guard__h161118 == 2'b11 && requestR[191:160] == 32'hFFFFFFFF &&
	      requestR[159];
    endcase
  end
  always@(requestR or guard__h161118)
  begin
    case (requestR[194:192])
      3'h2, 3'h3:
	  CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q163 =
	      requestR[191:160] == 32'hFFFFFFFF && requestR[159];
      3'h4:
	  CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q163 =
	      (guard__h161118 == 2'b0) ?
		requestR[191:160] == 32'hFFFFFFFF && requestR[159] :
		(guard__h161118 == 2'b01 || guard__h161118 == 2'b10 ||
		 guard__h161118 == 2'b11) &&
		requestR[191:160] == 32'hFFFFFFFF &&
		requestR[159];
      default: CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q163 =
		   requestR[194:192] == 3'h1 &&
		   requestR[191:160] == 32'hFFFFFFFF &&
		   requestR[159];
    endcase
  end
  always@(guard__h170426 or requestR)
  begin
    case (guard__h170426)
      2'b0, 2'b01, 2'b10:
	  CASE_guard70426_0b0_requestR_BITS_191_TO_160_E_ETC__q164 =
	      requestR[191:160] == 32'hFFFFFFFF && requestR[159];
      2'd3:
	  CASE_guard70426_0b0_requestR_BITS_191_TO_160_E_ETC__q164 =
	      guard__h170426 == 2'b11 && requestR[191:160] == 32'hFFFFFFFF &&
	      requestR[159];
    endcase
  end
  always@(requestR or guard__h170426)
  begin
    case (requestR[194:192])
      3'h2, 3'h3:
	  CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q165 =
	      requestR[191:160] == 32'hFFFFFFFF && requestR[159];
      3'h4:
	  CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q165 =
	      (guard__h170426 == 2'b0) ?
		requestR[191:160] == 32'hFFFFFFFF && requestR[159] :
		(guard__h170426 == 2'b01 || guard__h170426 == 2'b10 ||
		 guard__h170426 == 2'b11) &&
		requestR[191:160] == 32'hFFFFFFFF &&
		requestR[159];
      default: CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q165 =
		   requestR[194:192] == 3'h1 &&
		   requestR[191:160] == 32'hFFFFFFFF &&
		   requestR[159];
    endcase
  end
  always@(guard__h179493 or requestR)
  begin
    case (guard__h179493)
      2'b0, 2'b01, 2'b10:
	  CASE_guard79493_0b0_requestR_BITS_191_TO_160_E_ETC__q166 =
	      requestR[191:160] == 32'hFFFFFFFF && requestR[159];
      2'd3:
	  CASE_guard79493_0b0_requestR_BITS_191_TO_160_E_ETC__q166 =
	      guard__h179493 == 2'b11 && requestR[191:160] == 32'hFFFFFFFF &&
	      requestR[159];
    endcase
  end
  always@(requestR or guard__h179493)
  begin
    case (requestR[194:192])
      3'h2, 3'h3:
	  CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q167 =
	      requestR[191:160] == 32'hFFFFFFFF && requestR[159];
      3'h4:
	  CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q167 =
	      (guard__h179493 == 2'b0) ?
		requestR[191:160] == 32'hFFFFFFFF && requestR[159] :
		(guard__h179493 == 2'b01 || guard__h179493 == 2'b10 ||
		 guard__h179493 == 2'b11) &&
		requestR[191:160] == 32'hFFFFFFFF &&
		requestR[159];
      default: CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q167 =
		   requestR[194:192] == 3'h1 &&
		   requestR[191:160] == 32'hFFFFFFFF &&
		   requestR[159];
    endcase
  end
  always@(guard__h161118 or
	  _theResult___snd__h169030 or _theResult___sfd__h169735)
  begin
    case (guard__h161118)
      2'b0:
	  CASE_guard61118_0b0_theResult___snd69030_BITS__ETC__q168 =
	      _theResult___snd__h169030[56:5];
      2'b01, 2'b10, 2'b11:
	  CASE_guard61118_0b0_theResult___snd69030_BITS__ETC__q168 =
	      _theResult___sfd__h169735;
    endcase
  end
  always@(requestR or
	  _theResult___snd__h169030 or
	  IF_IF_IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFF_ETC___d4978 or
	  IF_IF_IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFF_ETC___d4976 or
	  CASE_guard61118_0b0_theResult___snd69030_BITS__ETC__q168)
  begin
    case (requestR[194:192])
      3'h1:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d4982 =
	      _theResult___snd__h169030[56:5];
      3'h2:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d4982 =
	      IF_IF_IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFF_ETC___d4978;
      3'h3:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d4982 =
	      IF_IF_IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFF_ETC___d4976;
      3'h4:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d4982 =
	      CASE_guard61118_0b0_theResult___snd69030_BITS__ETC__q168;
      default: IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d4982 =
		   52'd0;
    endcase
  end
  always@(guard__h161118 or
	  _theResult___snd__h169030 or
	  out_sfd__h169738 or _theResult___sfd__h169735)
  begin
    case (guard__h161118)
      2'b0, 2'b01:
	  CASE_guard61118_0b0_theResult___snd69030_BITS__ETC__q169 =
	      _theResult___snd__h169030[56:5];
      2'b10:
	  CASE_guard61118_0b0_theResult___snd69030_BITS__ETC__q169 =
	      out_sfd__h169738;
      2'b11:
	  CASE_guard61118_0b0_theResult___snd69030_BITS__ETC__q169 =
	      _theResult___sfd__h169735;
    endcase
  end
  always@(guard__h170426 or sfdin__h178646 or _theResult___sfd__h179382)
  begin
    case (guard__h170426)
      2'b0:
	  CASE_guard70426_0b0_sfdin78646_BITS_56_TO_5_0b_ETC__q170 =
	      sfdin__h178646[56:5];
      2'b01, 2'b10, 2'b11:
	  CASE_guard70426_0b0_sfdin78646_BITS_56_TO_5_0b_ETC__q170 =
	      _theResult___sfd__h179382;
    endcase
  end
  always@(requestR or
	  sfdin__h178646 or
	  IF_IF_IF_IF_3074_MINUS_SEXT_IF_requestR_BITS_1_ETC___d5005 or
	  IF_IF_IF_IF_3074_MINUS_SEXT_IF_requestR_BITS_1_ETC___d5003 or
	  CASE_guard70426_0b0_sfdin78646_BITS_56_TO_5_0b_ETC__q170)
  begin
    case (requestR[194:192])
      3'h1:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d5009 =
	      sfdin__h178646[56:5];
      3'h2:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d5009 =
	      IF_IF_IF_IF_3074_MINUS_SEXT_IF_requestR_BITS_1_ETC___d5005;
      3'h3:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d5009 =
	      IF_IF_IF_IF_3074_MINUS_SEXT_IF_requestR_BITS_1_ETC___d5003;
      3'h4:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d5009 =
	      CASE_guard70426_0b0_sfdin78646_BITS_56_TO_5_0b_ETC__q170;
      default: IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d5009 =
		   52'd0;
    endcase
  end
  always@(guard__h170426 or
	  sfdin__h178646 or out_sfd__h179385 or _theResult___sfd__h179382)
  begin
    case (guard__h170426)
      2'b0, 2'b01:
	  CASE_guard70426_0b0_sfdin78646_BITS_56_TO_5_0b_ETC__q171 =
	      sfdin__h178646[56:5];
      2'b10:
	  CASE_guard70426_0b0_sfdin78646_BITS_56_TO_5_0b_ETC__q171 =
	      out_sfd__h179385;
      2'b11:
	  CASE_guard70426_0b0_sfdin78646_BITS_56_TO_5_0b_ETC__q171 =
	      _theResult___sfd__h179382;
    endcase
  end
  always@(guard__h179493 or
	  _theResult___snd__h187429 or _theResult___sfd__h188164)
  begin
    case (guard__h179493)
      2'b0:
	  CASE_guard79493_0b0_theResult___snd87429_BITS__ETC__q172 =
	      _theResult___snd__h187429[56:5];
      2'b01, 2'b10, 2'b11:
	  CASE_guard79493_0b0_theResult___snd87429_BITS__ETC__q172 =
	      _theResult___sfd__h188164;
    endcase
  end
  always@(requestR or
	  _theResult___snd__h187429 or
	  IF_IF_IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFF_ETC___d5024 or
	  IF_IF_IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFF_ETC___d5022 or
	  CASE_guard79493_0b0_theResult___snd87429_BITS__ETC__q172)
  begin
    case (requestR[194:192])
      3'h1:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d5028 =
	      _theResult___snd__h187429[56:5];
      3'h2:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d5028 =
	      IF_IF_IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFF_ETC___d5024;
      3'h3:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d5028 =
	      IF_IF_IF_IF_requestR_BITS_191_TO_160_4_EQ_0xFF_ETC___d5022;
      3'h4:
	  IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d5028 =
	      CASE_guard79493_0b0_theResult___snd87429_BITS__ETC__q172;
      default: IF_requestR_BITS_194_TO_192_0_EQ_0x4_5_THEN_IF_ETC___d5028 =
		   52'd0;
    endcase
  end
  always@(guard__h179493 or
	  _theResult___snd__h187429 or
	  out_sfd__h188167 or _theResult___sfd__h188164)
  begin
    case (guard__h179493)
      2'b0, 2'b01:
	  CASE_guard79493_0b0_theResult___snd87429_BITS__ETC__q173 =
	      _theResult___snd__h187429[56:5];
      2'b10:
	  CASE_guard79493_0b0_theResult___snd87429_BITS__ETC__q173 =
	      out_sfd__h188167;
      2'b11:
	  CASE_guard79493_0b0_theResult___snd87429_BITS__ETC__q173 =
	      _theResult___sfd__h188164;
    endcase
  end
  // handling of inlined registers
  always@(posedge CLK)
  begin
    if (RST_N == `BSV_RESET_VALUE)
      begin
        cfg_verbosity <= `BSV_ASSIGNMENT_DELAY 4'd0;
	requestR <= `BSV_ASSIGNMENT_DELAY
	    215'h2AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
	resultR <= `BSV_ASSIGNMENT_DELAY 70'h0AAAAAAAAAAAAAAAAA;
	stateR <= `BSV_ASSIGNMENT_DELAY 2'd0;
      end
    else
      begin
        if (cfg_verbosity$EN)
	  cfg_verbosity <= `BSV_ASSIGNMENT_DELAY cfg_verbosity$D_IN;
	if (requestR$EN) requestR <= `BSV_ASSIGNMENT_DELAY requestR$D_IN;
	if (resultR$EN) resultR <= `BSV_ASSIGNMENT_DELAY resultR$D_IN;
	if (stateR$EN) stateR <= `BSV_ASSIGNMENT_DELAY stateR$D_IN;
      end
  end
  // synopsys translate_off
  `ifdef BSV_NO_INITIAL_BLOCKS
  `else // not BSV_NO_INITIAL_BLOCKS
  initial
  begin
    cfg_verbosity = 4'hA;
    requestR = 215'h2AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
    resultR = 70'h2AAAAAAAAAAAAAAAAA;
    stateR = 2'h2;
  end
  `endif // BSV_NO_INITIAL_BLOCKS
  // synopsys translate_on
endmodule