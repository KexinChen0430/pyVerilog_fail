module outputs
  wire [4 : 0] output_arbs_0_select,
	       output_arbs_1_select,
	       output_arbs_2_select,
	       output_arbs_3_select,
	       output_arbs_4_select;
  // register oas_0_token
  reg [4 : 0] oas_0_token;
  wire [4 : 0] oas_0_token$D_IN;
  wire oas_0_token$EN;
  // register oas_1_token
  reg [4 : 0] oas_1_token;
  wire [4 : 0] oas_1_token$D_IN;
  wire oas_1_token$EN;
  // register oas_2_token
  reg [4 : 0] oas_2_token;
  wire [4 : 0] oas_2_token$D_IN;
  wire oas_2_token$EN;
  // register oas_3_token
  reg [4 : 0] oas_3_token;
  wire [4 : 0] oas_3_token$D_IN;
  wire oas_3_token$EN;
  // register oas_4_token
  reg [4 : 0] oas_4_token;
  wire [4 : 0] oas_4_token$D_IN;
  wire oas_4_token$EN;
  // remaining internal signals
  wire [1 : 0] ab__h12572,
	       ab__h12587,
	       ab__h12602,
	       ab__h12617,
	       ab__h12632,
	       ab__h14013,
	       ab__h14460,
	       ab__h14853,
	       ab__h15197,
	       ab__h15492,
	       ab__h19612,
	       ab__h19627,
	       ab__h19642,
	       ab__h19657,
	       ab__h19672,
	       ab__h21053,
	       ab__h21500,
	       ab__h21893,
	       ab__h22237,
	       ab__h22532,
	       ab__h26652,
	       ab__h26667,
	       ab__h26682,
	       ab__h26697,
	       ab__h26712,
	       ab__h28093,
	       ab__h28540,
	       ab__h28933,
	       ab__h29277,
	       ab__h29572,
	       ab__h33692,
	       ab__h33707,
	       ab__h33722,
	       ab__h33737,
	       ab__h33752,
	       ab__h35133,
	       ab__h35580,
	       ab__h35973,
	       ab__h36317,
	       ab__h36612,
	       ab__h5532,
	       ab__h5547,
	       ab__h5562,
	       ab__h5577,
	       ab__h5592,
	       ab__h6973,
	       ab__h7420,
	       ab__h7813,
	       ab__h8157,
	       ab__h8452;
  wire NOT_gen_grant_carry_00_BIT_1_01_14_AND_NOT_gen_ETC___d328,
       NOT_gen_grant_carry_00_BIT_1_01_14_AND_NOT_gen_ETC___d348,
       NOT_gen_grant_carry_0_BIT_1_1_04_AND_NOT_gen_g_ETC___d118,
       NOT_gen_grant_carry_0_BIT_1_1_04_AND_NOT_gen_g_ETC___d138,
       NOT_gen_grant_carry_0_BIT_1_1_4_AND_NOT_gen_gr_ETC___d48,
       NOT_gen_grant_carry_0_BIT_1_1_4_AND_NOT_gen_gr_ETC___d68,
       NOT_gen_grant_carry_22_BIT_1_54_60_AND_NOT_gen_ETC___d276,
       NOT_gen_grant_carry_26_BIT_1_47_51_AND_NOT_gen_ETC___d267,
       NOT_gen_grant_carry_2_BIT_1_14_20_AND_NOT_gen__ETC___d136,
       NOT_gen_grant_carry_2_BIT_1_4_0_AND_NOT_gen_gr_ETC___d66,
       NOT_gen_grant_carry_30_BIT_1_31_44_AND_NOT_gen_ETC___d258,
       NOT_gen_grant_carry_30_BIT_1_31_44_AND_NOT_gen_ETC___d278,
       NOT_gen_grant_carry_52_BIT_1_84_90_AND_NOT_gen_ETC___d206,
       NOT_gen_grant_carry_56_BIT_1_77_81_AND_NOT_gen_ETC___d197,
       NOT_gen_grant_carry_60_BIT_1_61_74_AND_NOT_gen_ETC___d188,
       NOT_gen_grant_carry_60_BIT_1_61_74_AND_NOT_gen_ETC___d208,
       NOT_gen_grant_carry_6_BIT_1_07_11_AND_NOT_gen__ETC___d127,
       NOT_gen_grant_carry_6_BIT_1_7_1_AND_NOT_gen_gr_ETC___d57,
       NOT_gen_grant_carry_92_BIT_1_24_30_AND_NOT_gen_ETC___d346,
       NOT_gen_grant_carry_96_BIT_1_17_21_AND_NOT_gen_ETC___d337,
       ab_BIT_0___h13184,
       ab_BIT_0___h13291,
       ab_BIT_0___h13398,
       ab_BIT_0___h13505,
       ab_BIT_0___h14084,
       ab_BIT_0___h14220,
       ab_BIT_0___h14613,
       ab_BIT_0___h14957,
       ab_BIT_0___h15252,
       ab_BIT_0___h20224,
       ab_BIT_0___h20331,
       ab_BIT_0___h20438,
       ab_BIT_0___h20545,
       ab_BIT_0___h21124,
       ab_BIT_0___h21260,
       ab_BIT_0___h21653,
       ab_BIT_0___h21997,
       ab_BIT_0___h22292,
       ab_BIT_0___h27264,
       ab_BIT_0___h27371,
       ab_BIT_0___h27478,
       ab_BIT_0___h27585,
       ab_BIT_0___h28164,
       ab_BIT_0___h28300,
       ab_BIT_0___h28693,
       ab_BIT_0___h29037,
       ab_BIT_0___h29332,
       ab_BIT_0___h34304,
       ab_BIT_0___h34411,
       ab_BIT_0___h34518,
       ab_BIT_0___h34625,
       ab_BIT_0___h35204,
       ab_BIT_0___h35340,
       ab_BIT_0___h35733,
       ab_BIT_0___h36077,
       ab_BIT_0___h36372,
       ab_BIT_0___h6144,
       ab_BIT_0___h6251,
       ab_BIT_0___h6358,
       ab_BIT_0___h6465,
       ab_BIT_0___h7044,
       ab_BIT_0___h7180,
       ab_BIT_0___h7573,
       ab_BIT_0___h7917,
       ab_BIT_0___h8212,
       oas_0_token_BIT_0___h6142,
       oas_0_token_BIT_1___h6249,
       oas_0_token_BIT_2___h6356,
       oas_0_token_BIT_3___h6463,
       oas_0_token_BIT_4___h6570,
       oas_1_token_BIT_0___h13182,
       oas_1_token_BIT_1___h13289,
       oas_1_token_BIT_2___h13396,
       oas_1_token_BIT_3___h13503,
       oas_1_token_BIT_4___h13610,
       oas_2_token_BIT_0___h20222,
       oas_2_token_BIT_1___h20329,
       oas_2_token_BIT_2___h20436,
       oas_2_token_BIT_3___h20543,
       oas_2_token_BIT_4___h20650,
       oas_3_token_BIT_0___h27262,
       oas_3_token_BIT_1___h27369,
       oas_3_token_BIT_2___h27476,
       oas_3_token_BIT_3___h27583,
       oas_3_token_BIT_4___h27690,
       oas_4_token_BIT_0___h34302,
       oas_4_token_BIT_1___h34409,
       oas_4_token_BIT_2___h34516,
       oas_4_token_BIT_3___h34623,
       oas_4_token_BIT_4___h34730;
  // value method output_arbs_0_select
  assign output_arbs_0_select =
	     { ab__h5532[1] || ab__h6973[1],
	       !ab__h5532[1] && !ab__h6973[1] &&
	       (ab__h5547[1] || ab__h7420[1]),
	       NOT_gen_grant_carry_0_BIT_1_1_4_AND_NOT_gen_gr_ETC___d48,
	       !ab__h5532[1] && !ab__h6973[1] &&
	       NOT_gen_grant_carry_6_BIT_1_7_1_AND_NOT_gen_gr_ETC___d57,
	       NOT_gen_grant_carry_0_BIT_1_1_4_AND_NOT_gen_gr_ETC___d68 } ;
  // value method output_arbs_1_select
  assign output_arbs_1_select =
	     { ab__h12572[1] || ab__h14013[1],
	       !ab__h12572[1] && !ab__h14013[1] &&
	       (ab__h12587[1] || ab__h14460[1]),
	       NOT_gen_grant_carry_0_BIT_1_1_04_AND_NOT_gen_g_ETC___d118,
	       !ab__h12572[1] && !ab__h14013[1] &&
	       NOT_gen_grant_carry_6_BIT_1_07_11_AND_NOT_gen__ETC___d127,
	       NOT_gen_grant_carry_0_BIT_1_1_04_AND_NOT_gen_g_ETC___d138 } ;
  // value method output_arbs_2_select
  assign output_arbs_2_select =
	     { ab__h19612[1] || ab__h21053[1],
	       !ab__h19612[1] && !ab__h21053[1] &&
	       (ab__h19627[1] || ab__h21500[1]),
	       NOT_gen_grant_carry_60_BIT_1_61_74_AND_NOT_gen_ETC___d188,
	       !ab__h19612[1] && !ab__h21053[1] &&
	       NOT_gen_grant_carry_56_BIT_1_77_81_AND_NOT_gen_ETC___d197,
	       NOT_gen_grant_carry_60_BIT_1_61_74_AND_NOT_gen_ETC___d208 } ;
  // value method output_arbs_3_select
  assign output_arbs_3_select =
	     { ab__h26652[1] || ab__h28093[1],
	       !ab__h26652[1] && !ab__h28093[1] &&
	       (ab__h26667[1] || ab__h28540[1]),
	       NOT_gen_grant_carry_30_BIT_1_31_44_AND_NOT_gen_ETC___d258,
	       !ab__h26652[1] && !ab__h28093[1] &&
	       NOT_gen_grant_carry_26_BIT_1_47_51_AND_NOT_gen_ETC___d267,
	       NOT_gen_grant_carry_30_BIT_1_31_44_AND_NOT_gen_ETC___d278 } ;
  // value method output_arbs_4_select
  assign output_arbs_4_select =
	     { ab__h33692[1] || ab__h35133[1],
	       !ab__h33692[1] && !ab__h35133[1] &&
	       (ab__h33707[1] || ab__h35580[1]),
	       NOT_gen_grant_carry_00_BIT_1_01_14_AND_NOT_gen_ETC___d328,
	       !ab__h33692[1] && !ab__h35133[1] &&
	       NOT_gen_grant_carry_96_BIT_1_17_21_AND_NOT_gen_ETC___d337,
	       NOT_gen_grant_carry_00_BIT_1_01_14_AND_NOT_gen_ETC___d348 } ;
  // register oas_0_token
  assign oas_0_token$D_IN = { oas_0_token[0], oas_0_token[4:1] } ;
  assign oas_0_token$EN = EN_output_arbs_0_next ;
  // register oas_1_token
  assign oas_1_token$D_IN = { oas_1_token[0], oas_1_token[4:1] } ;
  assign oas_1_token$EN = EN_output_arbs_1_next ;
  // register oas_2_token
  assign oas_2_token$D_IN = { oas_2_token[0], oas_2_token[4:1] } ;
  assign oas_2_token$EN = EN_output_arbs_2_next ;
  // register oas_3_token
  assign oas_3_token$D_IN = { oas_3_token[0], oas_3_token[4:1] } ;
  assign oas_3_token$EN = EN_output_arbs_3_next ;
  // register oas_4_token
  assign oas_4_token$D_IN = { oas_4_token[0], oas_4_token[4:1] } ;
  assign oas_4_token$EN = EN_output_arbs_4_next ;
  // remaining internal signals
  module_gen_grant_carry instance_gen_grant_carry_45(.gen_grant_carry_c(1'd0),
						     .gen_grant_carry_r(output_arbs_0_select_requests[0]),
						     .gen_grant_carry_p(oas_0_token_BIT_0___h6142),
						     .gen_grant_carry(ab__h5592));
  module_gen_grant_carry instance_gen_grant_carry_1(.gen_grant_carry_c(ab_BIT_0___h6144),
						    .gen_grant_carry_r(output_arbs_0_select_requests[1]),
						    .gen_grant_carry_p(oas_0_token_BIT_1___h6249),
						    .gen_grant_carry(ab__h5577));
  module_gen_grant_carry instance_gen_grant_carry_0(.gen_grant_carry_c(ab_BIT_0___h6251),
						    .gen_grant_carry_r(output_arbs_0_select_requests[2]),
						    .gen_grant_carry_p(oas_0_token_BIT_2___h6356),
						    .gen_grant_carry(ab__h5562));
  module_gen_grant_carry instance_gen_grant_carry_2(.gen_grant_carry_c(ab_BIT_0___h6358),
						    .gen_grant_carry_r(output_arbs_0_select_requests[3]),
						    .gen_grant_carry_p(oas_0_token_BIT_3___h6463),
						    .gen_grant_carry(ab__h5547));
  module_gen_grant_carry instance_gen_grant_carry_3(.gen_grant_carry_c(ab_BIT_0___h6465),
						    .gen_grant_carry_r(output_arbs_0_select_requests[4]),
						    .gen_grant_carry_p(oas_0_token_BIT_4___h6570),
						    .gen_grant_carry(ab__h5532));
  module_gen_grant_carry instance_gen_grant_carry_4(.gen_grant_carry_c(ab_BIT_0___h7044),
						    .gen_grant_carry_r(output_arbs_0_select_requests[0]),
						    .gen_grant_carry_p(oas_0_token_BIT_0___h6142),
						    .gen_grant_carry(ab__h8452));
  module_gen_grant_carry instance_gen_grant_carry_5(.gen_grant_carry_c(ab_BIT_0___h8212),
						    .gen_grant_carry_r(output_arbs_0_select_requests[1]),
						    .gen_grant_carry_p(oas_0_token_BIT_1___h6249),
						    .gen_grant_carry(ab__h8157));
  module_gen_grant_carry instance_gen_grant_carry_6(.gen_grant_carry_c(ab_BIT_0___h7917),
						    .gen_grant_carry_r(output_arbs_0_select_requests[2]),
						    .gen_grant_carry_p(oas_0_token_BIT_2___h6356),
						    .gen_grant_carry(ab__h7813));
  module_gen_grant_carry instance_gen_grant_carry_7(.gen_grant_carry_c(ab_BIT_0___h7573),
						    .gen_grant_carry_r(output_arbs_0_select_requests[3]),
						    .gen_grant_carry_p(oas_0_token_BIT_3___h6463),
						    .gen_grant_carry(ab__h7420));
  module_gen_grant_carry instance_gen_grant_carry_8(.gen_grant_carry_c(ab_BIT_0___h7180),
						    .gen_grant_carry_r(output_arbs_0_select_requests[4]),
						    .gen_grant_carry_p(oas_0_token_BIT_4___h6570),
						    .gen_grant_carry(ab__h6973));
  module_gen_grant_carry instance_gen_grant_carry_46(.gen_grant_carry_c(1'd0),
						     .gen_grant_carry_r(output_arbs_1_select_requests[0]),
						     .gen_grant_carry_p(oas_1_token_BIT_0___h13182),
						     .gen_grant_carry(ab__h12632));
  module_gen_grant_carry instance_gen_grant_carry_9(.gen_grant_carry_c(ab_BIT_0___h13184),
						    .gen_grant_carry_r(output_arbs_1_select_requests[1]),
						    .gen_grant_carry_p(oas_1_token_BIT_1___h13289),
						    .gen_grant_carry(ab__h12617));
  module_gen_grant_carry instance_gen_grant_carry_10(.gen_grant_carry_c(ab_BIT_0___h13291),
						     .gen_grant_carry_r(output_arbs_1_select_requests[2]),
						     .gen_grant_carry_p(oas_1_token_BIT_2___h13396),
						     .gen_grant_carry(ab__h12602));
  module_gen_grant_carry instance_gen_grant_carry_11(.gen_grant_carry_c(ab_BIT_0___h13398),
						     .gen_grant_carry_r(output_arbs_1_select_requests[3]),
						     .gen_grant_carry_p(oas_1_token_BIT_3___h13503),
						     .gen_grant_carry(ab__h12587));
  module_gen_grant_carry instance_gen_grant_carry_12(.gen_grant_carry_c(ab_BIT_0___h13505),
						     .gen_grant_carry_r(output_arbs_1_select_requests[4]),
						     .gen_grant_carry_p(oas_1_token_BIT_4___h13610),
						     .gen_grant_carry(ab__h12572));
  module_gen_grant_carry instance_gen_grant_carry_13(.gen_grant_carry_c(ab_BIT_0___h14084),
						     .gen_grant_carry_r(output_arbs_1_select_requests[0]),
						     .gen_grant_carry_p(oas_1_token_BIT_0___h13182),
						     .gen_grant_carry(ab__h15492));
  module_gen_grant_carry instance_gen_grant_carry_14(.gen_grant_carry_c(ab_BIT_0___h15252),
						     .gen_grant_carry_r(output_arbs_1_select_requests[1]),
						     .gen_grant_carry_p(oas_1_token_BIT_1___h13289),
						     .gen_grant_carry(ab__h15197));
  module_gen_grant_carry instance_gen_grant_carry_15(.gen_grant_carry_c(ab_BIT_0___h14957),
						     .gen_grant_carry_r(output_arbs_1_select_requests[2]),
						     .gen_grant_carry_p(oas_1_token_BIT_2___h13396),
						     .gen_grant_carry(ab__h14853));
  module_gen_grant_carry instance_gen_grant_carry_16(.gen_grant_carry_c(ab_BIT_0___h14613),
						     .gen_grant_carry_r(output_arbs_1_select_requests[3]),
						     .gen_grant_carry_p(oas_1_token_BIT_3___h13503),
						     .gen_grant_carry(ab__h14460));
  module_gen_grant_carry instance_gen_grant_carry_17(.gen_grant_carry_c(ab_BIT_0___h14220),
						     .gen_grant_carry_r(output_arbs_1_select_requests[4]),
						     .gen_grant_carry_p(oas_1_token_BIT_4___h13610),
						     .gen_grant_carry(ab__h14013));
  module_gen_grant_carry instance_gen_grant_carry_47(.gen_grant_carry_c(1'd0),
						     .gen_grant_carry_r(output_arbs_2_select_requests[0]),
						     .gen_grant_carry_p(oas_2_token_BIT_0___h20222),
						     .gen_grant_carry(ab__h19672));
  module_gen_grant_carry instance_gen_grant_carry_18(.gen_grant_carry_c(ab_BIT_0___h20224),
						     .gen_grant_carry_r(output_arbs_2_select_requests[1]),
						     .gen_grant_carry_p(oas_2_token_BIT_1___h20329),
						     .gen_grant_carry(ab__h19657));
  module_gen_grant_carry instance_gen_grant_carry_19(.gen_grant_carry_c(ab_BIT_0___h20331),
						     .gen_grant_carry_r(output_arbs_2_select_requests[2]),
						     .gen_grant_carry_p(oas_2_token_BIT_2___h20436),
						     .gen_grant_carry(ab__h19642));
  module_gen_grant_carry instance_gen_grant_carry_20(.gen_grant_carry_c(ab_BIT_0___h20438),
						     .gen_grant_carry_r(output_arbs_2_select_requests[3]),
						     .gen_grant_carry_p(oas_2_token_BIT_3___h20543),
						     .gen_grant_carry(ab__h19627));
  module_gen_grant_carry instance_gen_grant_carry_21(.gen_grant_carry_c(ab_BIT_0___h20545),
						     .gen_grant_carry_r(output_arbs_2_select_requests[4]),
						     .gen_grant_carry_p(oas_2_token_BIT_4___h20650),
						     .gen_grant_carry(ab__h19612));
  module_gen_grant_carry instance_gen_grant_carry_22(.gen_grant_carry_c(ab_BIT_0___h21124),
						     .gen_grant_carry_r(output_arbs_2_select_requests[0]),
						     .gen_grant_carry_p(oas_2_token_BIT_0___h20222),
						     .gen_grant_carry(ab__h22532));
  module_gen_grant_carry instance_gen_grant_carry_23(.gen_grant_carry_c(ab_BIT_0___h22292),
						     .gen_grant_carry_r(output_arbs_2_select_requests[1]),
						     .gen_grant_carry_p(oas_2_token_BIT_1___h20329),
						     .gen_grant_carry(ab__h22237));
  module_gen_grant_carry instance_gen_grant_carry_24(.gen_grant_carry_c(ab_BIT_0___h21997),
						     .gen_grant_carry_r(output_arbs_2_select_requests[2]),
						     .gen_grant_carry_p(oas_2_token_BIT_2___h20436),
						     .gen_grant_carry(ab__h21893));
  module_gen_grant_carry instance_gen_grant_carry_25(.gen_grant_carry_c(ab_BIT_0___h21653),
						     .gen_grant_carry_r(output_arbs_2_select_requests[3]),
						     .gen_grant_carry_p(oas_2_token_BIT_3___h20543),
						     .gen_grant_carry(ab__h21500));
  module_gen_grant_carry instance_gen_grant_carry_26(.gen_grant_carry_c(ab_BIT_0___h21260),
						     .gen_grant_carry_r(output_arbs_2_select_requests[4]),
						     .gen_grant_carry_p(oas_2_token_BIT_4___h20650),
						     .gen_grant_carry(ab__h21053));
  module_gen_grant_carry instance_gen_grant_carry_48(.gen_grant_carry_c(1'd0),
						     .gen_grant_carry_r(output_arbs_3_select_requests[0]),
						     .gen_grant_carry_p(oas_3_token_BIT_0___h27262),
						     .gen_grant_carry(ab__h26712));
  module_gen_grant_carry instance_gen_grant_carry_27(.gen_grant_carry_c(ab_BIT_0___h27264),
						     .gen_grant_carry_r(output_arbs_3_select_requests[1]),
						     .gen_grant_carry_p(oas_3_token_BIT_1___h27369),
						     .gen_grant_carry(ab__h26697));
  module_gen_grant_carry instance_gen_grant_carry_28(.gen_grant_carry_c(ab_BIT_0___h27371),
						     .gen_grant_carry_r(output_arbs_3_select_requests[2]),
						     .gen_grant_carry_p(oas_3_token_BIT_2___h27476),
						     .gen_grant_carry(ab__h26682));
  module_gen_grant_carry instance_gen_grant_carry_29(.gen_grant_carry_c(ab_BIT_0___h27478),
						     .gen_grant_carry_r(output_arbs_3_select_requests[3]),
						     .gen_grant_carry_p(oas_3_token_BIT_3___h27583),
						     .gen_grant_carry(ab__h26667));
  module_gen_grant_carry instance_gen_grant_carry_30(.gen_grant_carry_c(ab_BIT_0___h27585),
						     .gen_grant_carry_r(output_arbs_3_select_requests[4]),
						     .gen_grant_carry_p(oas_3_token_BIT_4___h27690),
						     .gen_grant_carry(ab__h26652));
  module_gen_grant_carry instance_gen_grant_carry_31(.gen_grant_carry_c(ab_BIT_0___h28164),
						     .gen_grant_carry_r(output_arbs_3_select_requests[0]),
						     .gen_grant_carry_p(oas_3_token_BIT_0___h27262),
						     .gen_grant_carry(ab__h29572));
  module_gen_grant_carry instance_gen_grant_carry_32(.gen_grant_carry_c(ab_BIT_0___h29332),
						     .gen_grant_carry_r(output_arbs_3_select_requests[1]),
						     .gen_grant_carry_p(oas_3_token_BIT_1___h27369),
						     .gen_grant_carry(ab__h29277));
  module_gen_grant_carry instance_gen_grant_carry_33(.gen_grant_carry_c(ab_BIT_0___h29037),
						     .gen_grant_carry_r(output_arbs_3_select_requests[2]),
						     .gen_grant_carry_p(oas_3_token_BIT_2___h27476),
						     .gen_grant_carry(ab__h28933));
  module_gen_grant_carry instance_gen_grant_carry_34(.gen_grant_carry_c(ab_BIT_0___h28693),
						     .gen_grant_carry_r(output_arbs_3_select_requests[3]),
						     .gen_grant_carry_p(oas_3_token_BIT_3___h27583),
						     .gen_grant_carry(ab__h28540));
  module_gen_grant_carry instance_gen_grant_carry_35(.gen_grant_carry_c(ab_BIT_0___h28300),
						     .gen_grant_carry_r(output_arbs_3_select_requests[4]),
						     .gen_grant_carry_p(oas_3_token_BIT_4___h27690),
						     .gen_grant_carry(ab__h28093));
  module_gen_grant_carry instance_gen_grant_carry_49(.gen_grant_carry_c(1'd0),
						     .gen_grant_carry_r(output_arbs_4_select_requests[0]),
						     .gen_grant_carry_p(oas_4_token_BIT_0___h34302),
						     .gen_grant_carry(ab__h33752));
  module_gen_grant_carry instance_gen_grant_carry_36(.gen_grant_carry_c(ab_BIT_0___h34304),
						     .gen_grant_carry_r(output_arbs_4_select_requests[1]),
						     .gen_grant_carry_p(oas_4_token_BIT_1___h34409),
						     .gen_grant_carry(ab__h33737));
  module_gen_grant_carry instance_gen_grant_carry_37(.gen_grant_carry_c(ab_BIT_0___h34411),
						     .gen_grant_carry_r(output_arbs_4_select_requests[2]),
						     .gen_grant_carry_p(oas_4_token_BIT_2___h34516),
						     .gen_grant_carry(ab__h33722));
  module_gen_grant_carry instance_gen_grant_carry_38(.gen_grant_carry_c(ab_BIT_0___h34518),
						     .gen_grant_carry_r(output_arbs_4_select_requests[3]),
						     .gen_grant_carry_p(oas_4_token_BIT_3___h34623),
						     .gen_grant_carry(ab__h33707));
  module_gen_grant_carry instance_gen_grant_carry_39(.gen_grant_carry_c(ab_BIT_0___h34625),
						     .gen_grant_carry_r(output_arbs_4_select_requests[4]),
						     .gen_grant_carry_p(oas_4_token_BIT_4___h34730),
						     .gen_grant_carry(ab__h33692));
  module_gen_grant_carry instance_gen_grant_carry_40(.gen_grant_carry_c(ab_BIT_0___h35204),
						     .gen_grant_carry_r(output_arbs_4_select_requests[0]),
						     .gen_grant_carry_p(oas_4_token_BIT_0___h34302),
						     .gen_grant_carry(ab__h36612));
  module_gen_grant_carry instance_gen_grant_carry_41(.gen_grant_carry_c(ab_BIT_0___h36372),
						     .gen_grant_carry_r(output_arbs_4_select_requests[1]),
						     .gen_grant_carry_p(oas_4_token_BIT_1___h34409),
						     .gen_grant_carry(ab__h36317));
  module_gen_grant_carry instance_gen_grant_carry_42(.gen_grant_carry_c(ab_BIT_0___h36077),
						     .gen_grant_carry_r(output_arbs_4_select_requests[2]),
						     .gen_grant_carry_p(oas_4_token_BIT_2___h34516),
						     .gen_grant_carry(ab__h35973));
  module_gen_grant_carry instance_gen_grant_carry_43(.gen_grant_carry_c(ab_BIT_0___h35733),
						     .gen_grant_carry_r(output_arbs_4_select_requests[3]),
						     .gen_grant_carry_p(oas_4_token_BIT_3___h34623),
						     .gen_grant_carry(ab__h35580));
  module_gen_grant_carry instance_gen_grant_carry_44(.gen_grant_carry_c(ab_BIT_0___h35340),
						     .gen_grant_carry_r(output_arbs_4_select_requests[4]),
						     .gen_grant_carry_p(oas_4_token_BIT_4___h34730),
						     .gen_grant_carry(ab__h35133));
  assign NOT_gen_grant_carry_00_BIT_1_01_14_AND_NOT_gen_ETC___d328 =
	     !ab__h33692[1] && !ab__h35133[1] && !ab__h33707[1] &&
	     !ab__h35580[1] &&
	     (ab__h33722[1] || ab__h35973[1]) ;
  assign NOT_gen_grant_carry_00_BIT_1_01_14_AND_NOT_gen_ETC___d348 =
	     !ab__h33692[1] && !ab__h35133[1] && !ab__h33707[1] &&
	     !ab__h35580[1] &&
	     NOT_gen_grant_carry_92_BIT_1_24_30_AND_NOT_gen_ETC___d346 ;
  assign NOT_gen_grant_carry_0_BIT_1_1_04_AND_NOT_gen_g_ETC___d118 =
	     !ab__h12572[1] && !ab__h14013[1] && !ab__h12587[1] &&
	     !ab__h14460[1] &&
	     (ab__h12602[1] || ab__h14853[1]) ;
  assign NOT_gen_grant_carry_0_BIT_1_1_04_AND_NOT_gen_g_ETC___d138 =
	     !ab__h12572[1] && !ab__h14013[1] && !ab__h12587[1] &&
	     !ab__h14460[1] &&
	     NOT_gen_grant_carry_2_BIT_1_14_20_AND_NOT_gen__ETC___d136 ;
  assign NOT_gen_grant_carry_0_BIT_1_1_4_AND_NOT_gen_gr_ETC___d48 =
	     !ab__h5532[1] && !ab__h6973[1] && !ab__h5547[1] &&
	     !ab__h7420[1] &&
	     (ab__h5562[1] || ab__h7813[1]) ;
  assign NOT_gen_grant_carry_0_BIT_1_1_4_AND_NOT_gen_gr_ETC___d68 =
	     !ab__h5532[1] && !ab__h6973[1] && !ab__h5547[1] &&
	     !ab__h7420[1] &&
	     NOT_gen_grant_carry_2_BIT_1_4_0_AND_NOT_gen_gr_ETC___d66 ;
  assign NOT_gen_grant_carry_22_BIT_1_54_60_AND_NOT_gen_ETC___d276 =
	     !ab__h26682[1] && !ab__h28933[1] && !ab__h26697[1] &&
	     !ab__h29277[1] &&
	     (ab__h26712[1] || ab__h29572[1]) ;
  assign NOT_gen_grant_carry_26_BIT_1_47_51_AND_NOT_gen_ETC___d267 =
	     !ab__h26667[1] && !ab__h28540[1] && !ab__h26682[1] &&
	     !ab__h28933[1] &&
	     (ab__h26697[1] || ab__h29277[1]) ;
  assign NOT_gen_grant_carry_2_BIT_1_14_20_AND_NOT_gen__ETC___d136 =
	     !ab__h12602[1] && !ab__h14853[1] && !ab__h12617[1] &&
	     !ab__h15197[1] &&
	     (ab__h12632[1] || ab__h15492[1]) ;
  assign NOT_gen_grant_carry_2_BIT_1_4_0_AND_NOT_gen_gr_ETC___d66 =
	     !ab__h5562[1] && !ab__h7813[1] && !ab__h5577[1] &&
	     !ab__h8157[1] &&
	     (ab__h5592[1] || ab__h8452[1]) ;
  assign NOT_gen_grant_carry_30_BIT_1_31_44_AND_NOT_gen_ETC___d258 =
	     !ab__h26652[1] && !ab__h28093[1] && !ab__h26667[1] &&
	     !ab__h28540[1] &&
	     (ab__h26682[1] || ab__h28933[1]) ;
  assign NOT_gen_grant_carry_30_BIT_1_31_44_AND_NOT_gen_ETC___d278 =
	     !ab__h26652[1] && !ab__h28093[1] && !ab__h26667[1] &&
	     !ab__h28540[1] &&
	     NOT_gen_grant_carry_22_BIT_1_54_60_AND_NOT_gen_ETC___d276 ;
  assign NOT_gen_grant_carry_52_BIT_1_84_90_AND_NOT_gen_ETC___d206 =
	     !ab__h19642[1] && !ab__h21893[1] && !ab__h19657[1] &&
	     !ab__h22237[1] &&
	     (ab__h19672[1] || ab__h22532[1]) ;
  assign NOT_gen_grant_carry_56_BIT_1_77_81_AND_NOT_gen_ETC___d197 =
	     !ab__h19627[1] && !ab__h21500[1] && !ab__h19642[1] &&
	     !ab__h21893[1] &&
	     (ab__h19657[1] || ab__h22237[1]) ;
  assign NOT_gen_grant_carry_60_BIT_1_61_74_AND_NOT_gen_ETC___d188 =
	     !ab__h19612[1] && !ab__h21053[1] && !ab__h19627[1] &&
	     !ab__h21500[1] &&
	     (ab__h19642[1] || ab__h21893[1]) ;
  assign NOT_gen_grant_carry_60_BIT_1_61_74_AND_NOT_gen_ETC___d208 =
	     !ab__h19612[1] && !ab__h21053[1] && !ab__h19627[1] &&
	     !ab__h21500[1] &&
	     NOT_gen_grant_carry_52_BIT_1_84_90_AND_NOT_gen_ETC___d206 ;
  assign NOT_gen_grant_carry_6_BIT_1_07_11_AND_NOT_gen__ETC___d127 =
	     !ab__h12587[1] && !ab__h14460[1] && !ab__h12602[1] &&
	     !ab__h14853[1] &&
	     (ab__h12617[1] || ab__h15197[1]) ;
  assign NOT_gen_grant_carry_6_BIT_1_7_1_AND_NOT_gen_gr_ETC___d57 =
	     !ab__h5547[1] && !ab__h7420[1] && !ab__h5562[1] &&
	     !ab__h7813[1] &&
	     (ab__h5577[1] || ab__h8157[1]) ;
  assign NOT_gen_grant_carry_92_BIT_1_24_30_AND_NOT_gen_ETC___d346 =
	     !ab__h33722[1] && !ab__h35973[1] && !ab__h33737[1] &&
	     !ab__h36317[1] &&
	     (ab__h33752[1] || ab__h36612[1]) ;
  assign NOT_gen_grant_carry_96_BIT_1_17_21_AND_NOT_gen_ETC___d337 =
	     !ab__h33707[1] && !ab__h35580[1] && !ab__h33722[1] &&
	     !ab__h35973[1] &&
	     (ab__h33737[1] || ab__h36317[1]) ;
  assign ab_BIT_0___h13184 = ab__h12632[0] ;
  assign ab_BIT_0___h13291 = ab__h12617[0] ;
  assign ab_BIT_0___h13398 = ab__h12602[0] ;
  assign ab_BIT_0___h13505 = ab__h12587[0] ;
  assign ab_BIT_0___h14084 = ab__h12572[0] ;
  assign ab_BIT_0___h14220 = ab__h14460[0] ;
  assign ab_BIT_0___h14613 = ab__h14853[0] ;
  assign ab_BIT_0___h14957 = ab__h15197[0] ;
  assign ab_BIT_0___h15252 = ab__h15492[0] ;
  assign ab_BIT_0___h20224 = ab__h19672[0] ;
  assign ab_BIT_0___h20331 = ab__h19657[0] ;
  assign ab_BIT_0___h20438 = ab__h19642[0] ;
  assign ab_BIT_0___h20545 = ab__h19627[0] ;
  assign ab_BIT_0___h21124 = ab__h19612[0] ;
  assign ab_BIT_0___h21260 = ab__h21500[0] ;
  assign ab_BIT_0___h21653 = ab__h21893[0] ;
  assign ab_BIT_0___h21997 = ab__h22237[0] ;
  assign ab_BIT_0___h22292 = ab__h22532[0] ;
  assign ab_BIT_0___h27264 = ab__h26712[0] ;
  assign ab_BIT_0___h27371 = ab__h26697[0] ;
  assign ab_BIT_0___h27478 = ab__h26682[0] ;
  assign ab_BIT_0___h27585 = ab__h26667[0] ;
  assign ab_BIT_0___h28164 = ab__h26652[0] ;
  assign ab_BIT_0___h28300 = ab__h28540[0] ;
  assign ab_BIT_0___h28693 = ab__h28933[0] ;
  assign ab_BIT_0___h29037 = ab__h29277[0] ;
  assign ab_BIT_0___h29332 = ab__h29572[0] ;
  assign ab_BIT_0___h34304 = ab__h33752[0] ;
  assign ab_BIT_0___h34411 = ab__h33737[0] ;
  assign ab_BIT_0___h34518 = ab__h33722[0] ;
  assign ab_BIT_0___h34625 = ab__h33707[0] ;
  assign ab_BIT_0___h35204 = ab__h33692[0] ;
  assign ab_BIT_0___h35340 = ab__h35580[0] ;
  assign ab_BIT_0___h35733 = ab__h35973[0] ;
  assign ab_BIT_0___h36077 = ab__h36317[0] ;
  assign ab_BIT_0___h36372 = ab__h36612[0] ;
  assign ab_BIT_0___h6144 = ab__h5592[0] ;
  assign ab_BIT_0___h6251 = ab__h5577[0] ;
  assign ab_BIT_0___h6358 = ab__h5562[0] ;
  assign ab_BIT_0___h6465 = ab__h5547[0] ;
  assign ab_BIT_0___h7044 = ab__h5532[0] ;
  assign ab_BIT_0___h7180 = ab__h7420[0] ;
  assign ab_BIT_0___h7573 = ab__h7813[0] ;
  assign ab_BIT_0___h7917 = ab__h8157[0] ;
  assign ab_BIT_0___h8212 = ab__h8452[0] ;
  assign oas_0_token_BIT_0___h6142 = oas_0_token[0] ;
  assign oas_0_token_BIT_1___h6249 = oas_0_token[1] ;
  assign oas_0_token_BIT_2___h6356 = oas_0_token[2] ;
  assign oas_0_token_BIT_3___h6463 = oas_0_token[3] ;
  assign oas_0_token_BIT_4___h6570 = oas_0_token[4] ;
  assign oas_1_token_BIT_0___h13182 = oas_1_token[0] ;
  assign oas_1_token_BIT_1___h13289 = oas_1_token[1] ;
  assign oas_1_token_BIT_2___h13396 = oas_1_token[2] ;
  assign oas_1_token_BIT_3___h13503 = oas_1_token[3] ;
  assign oas_1_token_BIT_4___h13610 = oas_1_token[4] ;
  assign oas_2_token_BIT_0___h20222 = oas_2_token[0] ;
  assign oas_2_token_BIT_1___h20329 = oas_2_token[1] ;
  assign oas_2_token_BIT_2___h20436 = oas_2_token[2] ;
  assign oas_2_token_BIT_3___h20543 = oas_2_token[3] ;
  assign oas_2_token_BIT_4___h20650 = oas_2_token[4] ;
  assign oas_3_token_BIT_0___h27262 = oas_3_token[0] ;
  assign oas_3_token_BIT_1___h27369 = oas_3_token[1] ;
  assign oas_3_token_BIT_2___h27476 = oas_3_token[2] ;
  assign oas_3_token_BIT_3___h27583 = oas_3_token[3] ;
  assign oas_3_token_BIT_4___h27690 = oas_3_token[4] ;
  assign oas_4_token_BIT_0___h34302 = oas_4_token[0] ;
  assign oas_4_token_BIT_1___h34409 = oas_4_token[1] ;
  assign oas_4_token_BIT_2___h34516 = oas_4_token[2] ;
  assign oas_4_token_BIT_3___h34623 = oas_4_token[3] ;
  assign oas_4_token_BIT_4___h34730 = oas_4_token[4] ;
  // handling of inlined registers
  always@(posedge CLK)
  begin
    if (!RST_N)
      begin
        oas_0_token <= `BSV_ASSIGNMENT_DELAY 5'd1;
	oas_1_token <= `BSV_ASSIGNMENT_DELAY 5'd2;
	oas_2_token <= `BSV_ASSIGNMENT_DELAY 5'd4;
	oas_3_token <= `BSV_ASSIGNMENT_DELAY 5'd8;
	oas_4_token <= `BSV_ASSIGNMENT_DELAY 5'd16;
      end
    else
      begin
        if (oas_0_token$EN)
	  oas_0_token <= `BSV_ASSIGNMENT_DELAY oas_0_token$D_IN;
	if (oas_1_token$EN)
	  oas_1_token <= `BSV_ASSIGNMENT_DELAY oas_1_token$D_IN;
	if (oas_2_token$EN)
	  oas_2_token <= `BSV_ASSIGNMENT_DELAY oas_2_token$D_IN;
	if (oas_3_token$EN)
	  oas_3_token <= `BSV_ASSIGNMENT_DELAY oas_3_token$D_IN;
	if (oas_4_token$EN)
	  oas_4_token <= `BSV_ASSIGNMENT_DELAY oas_4_token$D_IN;
      end
  end
  // synopsys translate_off
  `ifdef BSV_NO_INITIAL_BLOCKS
  `else // not BSV_NO_INITIAL_BLOCKS
  initial
  begin
    oas_0_token = 5'h0A;
    oas_1_token = 5'h0A;
    oas_2_token = 5'h0A;
    oas_3_token = 5'h0A;
    oas_4_token = 5'h0A;
  end
  `endif // BSV_NO_INITIAL_BLOCKS
  // synopsys translate_on
endmodule