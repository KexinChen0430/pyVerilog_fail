module float32_to_int (
                         CLK, ce, inp, out
);
   parameter INSTANCE_NAME="INST";
  input wire CLK;
  input wire ce;
  input [31 : 0] inp;
  output [31 : 0] out;
   wire           clk;
   assign clk=CLK;
   wire [31:0]    a;
   assign a=inp;
   wire [31:0]    result;
   assign out=result;
  wire sig00000001;
  wire sig00000002;
  wire sig00000003;
  wire sig00000004;
  wire sig00000005;
  wire sig00000006;
  wire sig00000007;
  wire sig00000008;
  wire sig00000009;
  wire sig0000000a;
  wire sig0000000b;
  wire sig0000000c;
  wire sig0000000d;
  wire sig0000000e;
  wire sig0000000f;
  wire sig00000010;
  wire sig00000011;
  wire sig00000012;
  wire sig00000013;
  wire sig00000014;
  wire sig00000015;
  wire sig00000016;
  wire sig00000017;
  wire sig00000018;
  wire sig00000019;
  wire sig0000001a;
  wire sig0000001b;
  wire sig0000001c;
  wire sig0000001d;
  wire sig0000001e;
  wire sig0000001f;
  wire sig00000020;
  wire sig00000021;
  wire sig00000022;
  wire sig00000023;
  wire sig00000024;
  wire sig00000025;
  wire sig00000026;
  wire sig00000027;
  wire sig00000028;
  wire sig00000029;
  wire sig0000002a;
  wire sig0000002b;
  wire sig0000002c;
  wire sig0000002d;
  wire sig0000002e;
  wire sig0000002f;
  wire sig00000030;
  wire sig00000031;
  wire sig00000032;
  wire sig00000033;
  wire sig00000034;
  wire sig00000035;
  wire sig00000036;
  wire sig00000037;
  wire sig00000038;
  wire sig00000039;
  wire sig0000003a;
  wire sig0000003b;
  wire sig0000003c;
  wire sig0000003d;
  wire sig0000003e;
  wire sig0000003f;
  wire sig00000040;
  wire sig00000041;
  wire sig00000042;
  wire sig00000043;
  wire sig00000044;
  wire sig00000045;
  wire sig00000046;
  wire sig00000047;
  wire sig00000048;
  wire sig00000049;
  wire sig0000004a;
  wire sig0000004b;
  wire sig0000004c;
  wire sig0000004d;
  wire sig0000004e;
  wire sig0000004f;
  wire sig00000050;
  wire sig00000051;
  wire sig00000052;
  wire sig00000053;
  wire sig00000054;
  wire sig00000055;
  wire sig00000056;
  wire sig00000057;
  wire sig00000058;
  wire sig00000059;
  wire sig0000005a;
  wire sig0000005b;
  wire sig0000005c;
  wire sig0000005d;
  wire sig0000005e;
  wire sig0000005f;
  wire sig00000060;
  wire sig00000061;
  wire sig00000062;
  wire sig00000063;
  wire sig00000064;
  wire sig00000065;
  wire sig00000066;
  wire sig00000067;
  wire sig00000068;
  wire sig00000069;
  wire sig0000006a;
  wire sig0000006b;
  wire sig0000006c;
  wire sig0000006d;
  wire sig0000006e;
  wire sig0000006f;
  wire sig00000070;
  wire sig00000071;
  wire sig00000072;
  wire sig00000073;
  wire sig00000074;
  wire sig00000075;
  wire sig00000076;
  wire sig00000077;
  wire sig00000078;
  wire sig00000079;
  wire sig0000007a;
  wire sig0000007b;
  wire sig0000007c;
  wire sig0000007d;
  wire sig0000007e;
  wire sig0000007f;
  wire sig00000080;
  wire sig00000081;
  wire sig00000082;
  wire sig00000083;
  wire sig00000084;
  wire sig00000085;
  wire sig00000086;
  wire sig00000087;
  wire sig00000088;
  wire sig00000089;
  wire sig0000008a;
  wire sig0000008b;
  wire sig0000008c;
  wire sig0000008d;
  wire sig0000008e;
  wire sig0000008f;
  wire sig00000090;
  wire sig00000091;
  wire sig00000092;
  wire sig00000093;
  wire sig00000094;
  wire sig00000095;
  wire sig00000096;
  wire sig00000097;
  wire sig00000098;
  wire sig00000099;
  wire sig0000009a;
  wire sig0000009b;
  wire sig0000009c;
  wire sig0000009d;
  wire sig0000009e;
  wire sig0000009f;
  wire sig000000a0;
  wire sig000000a1;
  wire sig000000a2;
  wire sig000000a3;
  wire sig000000a4;
  wire sig000000a5;
  wire sig000000a6;
  wire sig000000a7;
  wire sig000000a8;
  wire sig000000a9;
  wire sig000000aa;
  wire sig000000ab;
  wire sig000000ac;
  wire sig000000ad;
  wire sig000000ae;
  wire sig000000af;
  wire sig000000b0;
  wire sig000000b1;
  wire sig000000b2;
  wire sig000000b3;
  wire sig000000b4;
  wire sig000000b5;
  wire sig000000b6;
  wire sig000000b7;
  wire sig000000b8;
  wire sig000000b9;
  wire sig000000ba;
  wire sig000000bb;
  wire sig000000bc;
  wire sig000000bd;
  wire sig000000be;
  wire sig000000bf;
  wire sig000000c0;
  wire sig000000c1;
  wire sig000000c2;
  wire sig000000c3;
  wire sig000000c4;
  wire sig000000c5;
  wire sig000000c6;
  wire sig000000c7;
  wire sig000000c8;
  wire sig000000c9;
  wire sig000000ca;
  wire sig000000cb;
  wire sig000000cc;
  wire sig000000cd;
  wire sig000000ce;
  wire sig000000cf;
  wire sig000000d0;
  wire sig000000d1;
  wire sig000000d2;
  wire sig000000d3;
  wire sig000000d4;
  wire sig000000d5;
  wire sig000000d6;
  wire sig000000d7;
  wire sig000000d8;
  wire sig000000d9;
  wire sig000000da;
  wire sig000000db;
  wire sig000000dc;
  wire sig000000dd;
  wire sig000000de;
  wire sig000000df;
  wire sig000000e0;
  wire sig000000e1;
  wire sig000000e2;
  wire sig000000e3;
  wire sig000000e4;
  wire sig000000e5;
  wire sig000000e6;
  wire sig000000e7;
  wire sig000000e8;
  wire sig000000e9;
  wire sig000000ea;
  wire sig000000eb;
  wire sig000000ec;
  wire sig000000ed;
  wire sig000000ee;
  wire sig000000ef;
  wire sig000000f0;
  wire sig000000f1;
  wire sig000000f2;
  wire sig000000f3;
  wire sig000000f4;
  wire sig000000f5;
  wire sig000000f6;
  wire sig000000f7;
  wire sig000000f8;
  wire sig000000f9;
  wire sig000000fa;
  wire sig000000fb;
  wire sig000000fc;
  wire sig000000fd;
  wire sig000000fe;
  wire sig000000ff;
  wire sig00000100;
  wire sig00000101;
  wire sig00000102;
  wire sig00000103;
  wire sig00000104;
  wire sig00000105;
  wire sig00000106;
  wire sig00000107;
  wire sig00000108;
  wire sig00000109;
  wire sig0000010a;
  wire sig0000010b;
  wire sig0000010c;
  wire sig0000010d;
  wire sig0000010e;
  wire sig0000010f;
  wire sig00000110;
  wire sig00000111;
  wire sig00000112;
  wire sig00000113;
  wire sig00000114;
  wire sig00000115;
  wire sig00000116;
  wire sig00000117;
  wire sig00000118;
  wire sig00000119;
  wire sig0000011a;
  wire sig0000011b;
  wire sig0000011c;
  wire sig0000011d;
  wire sig0000011e;
  wire sig0000011f;
  wire sig00000120;
  wire sig00000121;
  wire sig00000122;
  wire sig00000123;
  wire sig00000124;
  wire sig00000125;
  wire sig00000126;
  wire sig00000127;
  wire sig00000128;
  wire sig00000129;
  wire sig0000012a;
  wire sig0000012b;
  wire sig0000012c;
  wire sig0000012d;
  wire sig0000012e;
  wire sig0000012f;
  wire sig00000130;
  wire sig00000131;
  wire sig00000132;
  wire sig00000133;
  wire sig00000134;
  wire sig00000135;
  wire sig00000136;
  wire sig00000137;
  wire sig00000138;
  wire sig00000139;
  wire sig0000013a;
  wire sig0000013b;
  wire sig0000013c;
  wire sig0000013d;
  wire sig0000013e;
  wire sig0000013f;
  wire sig00000140;
  wire sig00000141;
  wire sig00000142;
  wire sig00000143;
  wire sig00000144;
  wire sig00000145;
  wire sig00000146;
  wire sig00000147;
  wire sig00000148;
  wire sig00000149;
  wire sig0000014a;
  wire sig0000014b;
  wire sig0000014c;
  wire sig0000014d;
  wire sig0000014e;
  wire sig0000014f;
  wire sig00000150;
  wire sig00000151;
  wire sig00000152;
  wire sig00000153;
  wire sig00000154;
  wire sig00000155;
  wire sig00000156;
  wire sig00000157;
  wire sig00000158;
  wire sig00000159;
  wire sig0000015a;
  wire sig0000015b;
  wire sig0000015c;
  wire sig0000015d;
  wire sig0000015e;
  wire sig0000015f;
  wire sig00000160;
  wire sig00000161;
  wire sig00000162;
  wire sig00000163;
  wire sig00000164;
  wire sig00000165;
  wire sig00000166;
  wire sig00000167;
  wire sig00000168;
  wire sig00000169;
  wire sig0000016a;
  wire sig0000016b;
  wire sig0000016c;
  wire sig0000016d;
  wire sig0000016e;
  wire sig0000016f;
  wire sig00000170;
  wire sig00000171;
  wire sig00000172;
  wire sig00000173;
  wire sig00000174;
  wire sig00000175;
  wire sig00000176;
  wire sig00000177;
  wire sig00000178;
  wire sig00000179;
  wire sig0000017a;
  wire sig0000017b;
  wire sig0000017c;
  wire sig0000017d;
  wire sig0000017e;
  wire sig0000017f;
  wire sig00000180;
  wire sig00000181;
  wire sig00000182;
  wire sig00000183;
  wire sig00000184;
  wire sig00000185;
  wire sig00000186;
  wire sig00000187;
  wire sig00000188;
  wire sig00000189;
  wire sig0000018a;
  wire sig0000018b;
  wire sig0000018c;
  wire sig0000018d;
  wire sig0000018e;
  wire sig0000018f;
  wire sig00000190;
  wire sig00000191;
  wire sig00000192;
  wire sig00000193;
  wire sig00000194;
  wire sig00000195;
  wire sig00000196;
  wire sig00000197;
  wire sig00000198;
  wire sig00000199;
  wire sig0000019a;
  wire sig0000019b;
  wire sig0000019c;
  wire sig0000019d;
  wire sig0000019e;
  wire sig0000019f;
  wire sig000001a0;
  wire sig000001a1;
  wire sig000001a2;
  wire sig000001a3;
  wire sig000001a4;
  wire sig000001a5;
  wire sig000001a6;
  wire sig000001a7;
  wire sig000001a8;
  wire sig000001a9;
  wire sig000001aa;
  wire sig000001ab;
  wire sig000001ac;
  wire sig000001ad;
  wire sig000001ae;
  wire sig000001af;
  wire sig000001b0;
  wire sig000001b1;
  wire sig000001b2;
  wire sig000001b3;
  wire sig000001b4;
  wire sig000001b5;
  wire sig000001b6;
  wire sig000001b7;
  wire sig000001b8;
  wire sig000001b9;
  wire sig000001ba;
  wire sig000001bb;
  wire sig000001bc;
  wire sig000001bd;
  wire sig000001be;
  wire sig000001bf;
  wire sig000001c0;
  wire sig000001c1;
  wire sig000001c2;
  wire sig000001c3;
  wire sig000001c4;
  wire sig000001c5;
  wire sig000001c6;
  wire sig000001c7;
  wire sig000001c8;
  wire sig000001c9;
  wire sig000001ca;
  wire sig000001cb;
  wire sig000001cc;
  wire sig000001cd;
  wire sig000001ce;
  wire sig000001cf;
  wire sig000001d0;
  wire sig000001d1;
  wire sig000001d2;
  wire sig000001d3;
  wire sig000001d4;
  wire sig000001d5;
  wire sig000001d6;
  wire sig000001d7;
  wire sig000001d8;
  wire sig000001d9;
  wire sig000001da;
  wire sig000001db;
  wire sig000001dc;
  wire sig000001dd;
  wire sig000001de;
  wire sig000001df;
  wire sig000001e0;
  wire sig000001e1;
  wire sig000001e2;
  wire sig000001e3;
  wire sig000001e4;
  wire sig000001e5;
  wire sig000001e6;
  wire sig000001e7;
  wire sig000001e8;
  wire sig000001e9;
  wire sig000001ea;
  wire sig000001eb;
  wire sig000001ec;
  wire sig000001ed;
  wire sig000001ee;
  wire NLW_blk00000008_O_UNCONNECTED;
  wire NLW_blk000000d2_O_UNCONNECTED;
  wire NLW_blk00000113_O_UNCONNECTED;
  wire NLW_blk00000206_Q15_UNCONNECTED;
  wire NLW_blk00000208_Q15_UNCONNECTED;
  wire NLW_blk0000020a_Q15_UNCONNECTED;
  wire NLW_blk0000020c_Q15_UNCONNECTED;
  wire NLW_blk0000020e_Q15_UNCONNECTED;
  wire NLW_blk00000210_Q15_UNCONNECTED;
  wire [31 : 0] \U0/op_inst/FLT_PT_OP/FLT_TO_FIX_OP.SPD.OP/RESULT ;
  assign
    result[31] = \U0/op_inst/FLT_PT_OP/FLT_TO_FIX_OP.SPD.OP/RESULT [31],
    result[30] = \U0/op_inst/FLT_PT_OP/FLT_TO_FIX_OP.SPD.OP/RESULT [30],
    result[29] = \U0/op_inst/FLT_PT_OP/FLT_TO_FIX_OP.SPD.OP/RESULT [29],
    result[28] = \U0/op_inst/FLT_PT_OP/FLT_TO_FIX_OP.SPD.OP/RESULT [28],
    result[27] = \U0/op_inst/FLT_PT_OP/FLT_TO_FIX_OP.SPD.OP/RESULT [27],
    result[26] = \U0/op_inst/FLT_PT_OP/FLT_TO_FIX_OP.SPD.OP/RESULT [26],
    result[25] = \U0/op_inst/FLT_PT_OP/FLT_TO_FIX_OP.SPD.OP/RESULT [25],
    result[24] = \U0/op_inst/FLT_PT_OP/FLT_TO_FIX_OP.SPD.OP/RESULT [24],
    result[23] = \U0/op_inst/FLT_PT_OP/FLT_TO_FIX_OP.SPD.OP/RESULT [23],
    result[22] = \U0/op_inst/FLT_PT_OP/FLT_TO_FIX_OP.SPD.OP/RESULT [22],
    result[21] = \U0/op_inst/FLT_PT_OP/FLT_TO_FIX_OP.SPD.OP/RESULT [21],
    result[20] = \U0/op_inst/FLT_PT_OP/FLT_TO_FIX_OP.SPD.OP/RESULT [20],
    result[19] = \U0/op_inst/FLT_PT_OP/FLT_TO_FIX_OP.SPD.OP/RESULT [19],
    result[18] = \U0/op_inst/FLT_PT_OP/FLT_TO_FIX_OP.SPD.OP/RESULT [18],
    result[17] = \U0/op_inst/FLT_PT_OP/FLT_TO_FIX_OP.SPD.OP/RESULT [17],
    result[16] = \U0/op_inst/FLT_PT_OP/FLT_TO_FIX_OP.SPD.OP/RESULT [16],
    result[15] = \U0/op_inst/FLT_PT_OP/FLT_TO_FIX_OP.SPD.OP/RESULT [15],
    result[14] = \U0/op_inst/FLT_PT_OP/FLT_TO_FIX_OP.SPD.OP/RESULT [14],
    result[13] = \U0/op_inst/FLT_PT_OP/FLT_TO_FIX_OP.SPD.OP/RESULT [13],
    result[12] = \U0/op_inst/FLT_PT_OP/FLT_TO_FIX_OP.SPD.OP/RESULT [12],
    result[11] = \U0/op_inst/FLT_PT_OP/FLT_TO_FIX_OP.SPD.OP/RESULT [11],
    result[10] = \U0/op_inst/FLT_PT_OP/FLT_TO_FIX_OP.SPD.OP/RESULT [10],
    result[9] = \U0/op_inst/FLT_PT_OP/FLT_TO_FIX_OP.SPD.OP/RESULT [9],
    result[8] = \U0/op_inst/FLT_PT_OP/FLT_TO_FIX_OP.SPD.OP/RESULT [8],
    result[7] = \U0/op_inst/FLT_PT_OP/FLT_TO_FIX_OP.SPD.OP/RESULT [7],
    result[6] = \U0/op_inst/FLT_PT_OP/FLT_TO_FIX_OP.SPD.OP/RESULT [6],
    result[5] = \U0/op_inst/FLT_PT_OP/FLT_TO_FIX_OP.SPD.OP/RESULT [5],
    result[4] = \U0/op_inst/FLT_PT_OP/FLT_TO_FIX_OP.SPD.OP/RESULT [4],
    result[3] = \U0/op_inst/FLT_PT_OP/FLT_TO_FIX_OP.SPD.OP/RESULT [3],
    result[2] = \U0/op_inst/FLT_PT_OP/FLT_TO_FIX_OP.SPD.OP/RESULT [2],
    result[1] = \U0/op_inst/FLT_PT_OP/FLT_TO_FIX_OP.SPD.OP/RESULT [1],
    result[0] = \U0/op_inst/FLT_PT_OP/FLT_TO_FIX_OP.SPD.OP/RESULT [0];
  VCC   blk00000001 (
    .P(sig00000001)
  );
  GND   blk00000002 (
    .G(sig00000002)
  );
  MUXCY   blk00000003 (
    .CI(sig00000001),
    .DI(sig00000002),
    .S(sig0000000a),
    .O(sig00000004)
  );
  MUXCY   blk00000004 (
    .CI(sig00000004),
    .DI(sig00000002),
    .S(sig0000000b),
    .O(sig00000005)
  );
  MUXCY   blk00000005 (
    .CI(sig00000005),
    .DI(sig00000002),
    .S(sig0000000c),
    .O(sig00000006)
  );
  MUXCY   blk00000006 (
    .CI(sig00000006),
    .DI(sig00000002),
    .S(sig0000000d),
    .O(sig00000007)
  );
  MUXCY   blk00000007 (
    .CI(sig00000007),
    .DI(sig00000002),
    .S(sig0000000e),
    .O(sig00000008)
  );
  MUXCY   blk00000008 (
    .CI(sig00000008),
    .DI(sig00000002),
    .S(sig00000009),
    .O(NLW_blk00000008_O_UNCONNECTED)
  );
  MUXCY   blk00000009 (
    .CI(sig00000013),
    .DI(sig00000002),
    .S(sig00000011),
    .O(sig00000012)
  );
  MUXCY   blk0000000a (
    .CI(sig00000001),
    .DI(sig00000002),
    .S(sig00000010),
    .O(sig00000013)
  );
  MUXCY   blk0000000b (
    .CI(sig00000001),
    .DI(sig00000002),
    .S(sig00000017),
    .O(sig00000015)
  );
  MUXCY   blk0000000c (
    .CI(sig00000015),
    .DI(sig00000002),
    .S(sig00000018),
    .O(sig00000016)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000000d (
    .C(clk),
    .CE(ce),
    .D(a[31]),
    .Q(sig000000cd)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000000e (
    .C(clk),
    .CE(ce),
    .D(sig0000001d),
    .Q(sig000000aa)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000000f (
    .C(clk),
    .CE(ce),
    .D(sig00000086),
    .Q(sig00000065)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000010 (
    .C(clk),
    .CE(ce),
    .D(sig00000012),
    .Q(sig000000ce)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000011 (
    .C(clk),
    .CE(ce),
    .D(sig00000016),
    .Q(sig00000014)
  );
  FDE   blk00000012 (
    .C(clk),
    .CE(ce),
    .D(sig00000019),
    .Q(\U0/op_inst/FLT_PT_OP/FLT_TO_FIX_OP.SPD.OP/RESULT [31])
  );
  FDE   blk00000013 (
    .C(clk),
    .CE(ce),
    .D(sig00000045),
    .Q(\U0/op_inst/FLT_PT_OP/FLT_TO_FIX_OP.SPD.OP/RESULT [30])
  );
  FDE   blk00000014 (
    .C(clk),
    .CE(ce),
    .D(sig00000044),
    .Q(\U0/op_inst/FLT_PT_OP/FLT_TO_FIX_OP.SPD.OP/RESULT [29])
  );
  FDE   blk00000015 (
    .C(clk),
    .CE(ce),
    .D(sig00000043),
    .Q(\U0/op_inst/FLT_PT_OP/FLT_TO_FIX_OP.SPD.OP/RESULT [28])
  );
  FDE   blk00000016 (
    .C(clk),
    .CE(ce),
    .D(sig00000042),
    .Q(\U0/op_inst/FLT_PT_OP/FLT_TO_FIX_OP.SPD.OP/RESULT [27])
  );
  FDE   blk00000017 (
    .C(clk),
    .CE(ce),
    .D(sig00000041),
    .Q(\U0/op_inst/FLT_PT_OP/FLT_TO_FIX_OP.SPD.OP/RESULT [26])
  );
  FDE   blk00000018 (
    .C(clk),
    .CE(ce),
    .D(sig00000040),
    .Q(\U0/op_inst/FLT_PT_OP/FLT_TO_FIX_OP.SPD.OP/RESULT [25])
  );
  FDE   blk00000019 (
    .C(clk),
    .CE(ce),
    .D(sig0000003f),
    .Q(\U0/op_inst/FLT_PT_OP/FLT_TO_FIX_OP.SPD.OP/RESULT [24])
  );
  FDE   blk0000001a (
    .C(clk),
    .CE(ce),
    .D(sig0000003e),
    .Q(\U0/op_inst/FLT_PT_OP/FLT_TO_FIX_OP.SPD.OP/RESULT [23])
  );
  FDE   blk0000001b (
    .C(clk),
    .CE(ce),
    .D(sig0000003d),
    .Q(\U0/op_inst/FLT_PT_OP/FLT_TO_FIX_OP.SPD.OP/RESULT [22])
  );
  FDE   blk0000001c (
    .C(clk),
    .CE(ce),
    .D(sig0000003c),
    .Q(\U0/op_inst/FLT_PT_OP/FLT_TO_FIX_OP.SPD.OP/RESULT [21])
  );
  FDE   blk0000001d (
    .C(clk),
    .CE(ce),
    .D(sig0000003b),
    .Q(\U0/op_inst/FLT_PT_OP/FLT_TO_FIX_OP.SPD.OP/RESULT [20])
  );
  FDE   blk0000001e (
    .C(clk),
    .CE(ce),
    .D(sig0000003a),
    .Q(\U0/op_inst/FLT_PT_OP/FLT_TO_FIX_OP.SPD.OP/RESULT [19])
  );
  FDE   blk0000001f (
    .C(clk),
    .CE(ce),
    .D(sig00000039),
    .Q(\U0/op_inst/FLT_PT_OP/FLT_TO_FIX_OP.SPD.OP/RESULT [18])
  );
  FDE   blk00000020 (
    .C(clk),
    .CE(ce),
    .D(sig00000038),
    .Q(\U0/op_inst/FLT_PT_OP/FLT_TO_FIX_OP.SPD.OP/RESULT [17])
  );
  FDE   blk00000021 (
    .C(clk),
    .CE(ce),
    .D(sig00000037),
    .Q(\U0/op_inst/FLT_PT_OP/FLT_TO_FIX_OP.SPD.OP/RESULT [16])
  );
  FDE   blk00000022 (
    .C(clk),
    .CE(ce),
    .D(sig00000036),
    .Q(\U0/op_inst/FLT_PT_OP/FLT_TO_FIX_OP.SPD.OP/RESULT [15])
  );
  FDE   blk00000023 (
    .C(clk),
    .CE(ce),
    .D(sig00000035),
    .Q(\U0/op_inst/FLT_PT_OP/FLT_TO_FIX_OP.SPD.OP/RESULT [14])
  );
  FDE   blk00000024 (
    .C(clk),
    .CE(ce),
    .D(sig00000034),
    .Q(\U0/op_inst/FLT_PT_OP/FLT_TO_FIX_OP.SPD.OP/RESULT [13])
  );
  FDE   blk00000025 (
    .C(clk),
    .CE(ce),
    .D(sig00000033),
    .Q(\U0/op_inst/FLT_PT_OP/FLT_TO_FIX_OP.SPD.OP/RESULT [12])
  );
  FDE   blk00000026 (
    .C(clk),
    .CE(ce),
    .D(sig00000032),
    .Q(\U0/op_inst/FLT_PT_OP/FLT_TO_FIX_OP.SPD.OP/RESULT [11])
  );
  FDE   blk00000027 (
    .C(clk),
    .CE(ce),
    .D(sig00000031),
    .Q(\U0/op_inst/FLT_PT_OP/FLT_TO_FIX_OP.SPD.OP/RESULT [10])
  );
  FDE   blk00000028 (
    .C(clk),
    .CE(ce),
    .D(sig00000030),
    .Q(\U0/op_inst/FLT_PT_OP/FLT_TO_FIX_OP.SPD.OP/RESULT [9])
  );
  FDE   blk00000029 (
    .C(clk),
    .CE(ce),
    .D(sig0000002f),
    .Q(\U0/op_inst/FLT_PT_OP/FLT_TO_FIX_OP.SPD.OP/RESULT [8])
  );
  FDE   blk0000002a (
    .C(clk),
    .CE(ce),
    .D(sig0000002e),
    .Q(\U0/op_inst/FLT_PT_OP/FLT_TO_FIX_OP.SPD.OP/RESULT [7])
  );
  FDE   blk0000002b (
    .C(clk),
    .CE(ce),
    .D(sig0000002d),
    .Q(\U0/op_inst/FLT_PT_OP/FLT_TO_FIX_OP.SPD.OP/RESULT [6])
  );
  FDE   blk0000002c (
    .C(clk),
    .CE(ce),
    .D(sig0000002c),
    .Q(\U0/op_inst/FLT_PT_OP/FLT_TO_FIX_OP.SPD.OP/RESULT [5])
  );
  FDE   blk0000002d (
    .C(clk),
    .CE(ce),
    .D(sig0000002b),
    .Q(\U0/op_inst/FLT_PT_OP/FLT_TO_FIX_OP.SPD.OP/RESULT [4])
  );
  FDE   blk0000002e (
    .C(clk),
    .CE(ce),
    .D(sig0000002a),
    .Q(\U0/op_inst/FLT_PT_OP/FLT_TO_FIX_OP.SPD.OP/RESULT [3])
  );
  FDE   blk0000002f (
    .C(clk),
    .CE(ce),
    .D(sig00000029),
    .Q(\U0/op_inst/FLT_PT_OP/FLT_TO_FIX_OP.SPD.OP/RESULT [2])
  );
  FDE   blk00000030 (
    .C(clk),
    .CE(ce),
    .D(sig00000028),
    .Q(\U0/op_inst/FLT_PT_OP/FLT_TO_FIX_OP.SPD.OP/RESULT [1])
  );
  FDE   blk00000031 (
    .C(clk),
    .CE(ce),
    .D(sig00000027),
    .Q(\U0/op_inst/FLT_PT_OP/FLT_TO_FIX_OP.SPD.OP/RESULT [0])
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000032 (
    .C(clk),
    .CE(ce),
    .D(a[22]),
    .Q(sig000000cc)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000033 (
    .C(clk),
    .CE(ce),
    .D(a[21]),
    .Q(sig000000cb)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000034 (
    .C(clk),
    .CE(ce),
    .D(a[20]),
    .Q(sig000000ca)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000035 (
    .C(clk),
    .CE(ce),
    .D(a[19]),
    .Q(sig000000c9)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000036 (
    .C(clk),
    .CE(ce),
    .D(a[18]),
    .Q(sig000000c8)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000037 (
    .C(clk),
    .CE(ce),
    .D(a[17]),
    .Q(sig000000c7)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000038 (
    .C(clk),
    .CE(ce),
    .D(a[16]),
    .Q(sig000000c6)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000039 (
    .C(clk),
    .CE(ce),
    .D(a[15]),
    .Q(sig000000c5)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000003a (
    .C(clk),
    .CE(ce),
    .D(a[14]),
    .Q(sig000000c4)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000003b (
    .C(clk),
    .CE(ce),
    .D(a[13]),
    .Q(sig000000c3)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000003c (
    .C(clk),
    .CE(ce),
    .D(a[12]),
    .Q(sig000000c2)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000003d (
    .C(clk),
    .CE(ce),
    .D(a[11]),
    .Q(sig000000c1)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000003e (
    .C(clk),
    .CE(ce),
    .D(a[10]),
    .Q(sig000000c0)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000003f (
    .C(clk),
    .CE(ce),
    .D(a[9]),
    .Q(sig000000bf)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000040 (
    .C(clk),
    .CE(ce),
    .D(a[8]),
    .Q(sig000000be)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000041 (
    .C(clk),
    .CE(ce),
    .D(a[7]),
    .Q(sig000000bd)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000042 (
    .C(clk),
    .CE(ce),
    .D(a[6]),
    .Q(sig000000bc)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000043 (
    .C(clk),
    .CE(ce),
    .D(a[5]),
    .Q(sig000000bb)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000044 (
    .C(clk),
    .CE(ce),
    .D(a[4]),
    .Q(sig000000ba)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000045 (
    .C(clk),
    .CE(ce),
    .D(a[3]),
    .Q(sig000000b9)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000046 (
    .C(clk),
    .CE(ce),
    .D(a[2]),
    .Q(sig000000b8)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000047 (
    .C(clk),
    .CE(ce),
    .D(a[1]),
    .Q(sig000000b7)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000048 (
    .C(clk),
    .CE(ce),
    .D(a[0]),
    .Q(sig000000b6)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000049 (
    .C(clk),
    .CE(ce),
    .D(sig00000026),
    .Q(sig000000b5)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000004a (
    .C(clk),
    .CE(ce),
    .D(sig00000025),
    .Q(sig000000b4)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000004b (
    .C(clk),
    .CE(ce),
    .D(sig00000024),
    .Q(sig000000b3)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000004c (
    .C(clk),
    .CE(ce),
    .D(sig00000023),
    .Q(sig000000b2)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000004d (
    .C(clk),
    .CE(ce),
    .D(sig00000022),
    .Q(sig000000b1)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000004e (
    .C(clk),
    .CE(ce),
    .D(sig00000021),
    .Q(sig000000b0)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000004f (
    .C(clk),
    .CE(ce),
    .D(sig00000020),
    .Q(sig000000af)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000050 (
    .C(clk),
    .CE(ce),
    .D(a[24]),
    .Q(sig000000ae)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000051 (
    .C(clk),
    .CE(ce),
    .D(sig0000000f),
    .Q(sig000000ad)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000052 (
    .C(clk),
    .CE(ce),
    .D(sig0000001f),
    .Q(sig000000ac)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000053 (
    .C(clk),
    .CE(ce),
    .D(sig0000001e),
    .Q(sig000000ab)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000054 (
    .C(clk),
    .CE(ce),
    .D(sig0000001c),
    .Q(sig000000d0)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000055 (
    .C(clk),
    .CE(ce),
    .D(sig0000001b),
    .Q(sig000000cf)
  );
  MUXF8   blk00000056 (
    .I0(sig000000d8),
    .I1(sig000000d7),
    .S(sig00000002),
    .O(sig000000d6)
  );
  MUXF7   blk00000057 (
    .I0(sig000001e5),
    .I1(sig000001e6),
    .S(sig000000e1),
    .O(sig000000d7)
  );
  MUXF7   blk00000058 (
    .I0(sig000001e7),
    .I1(sig000001e8),
    .S(sig000000e1),
    .O(sig000000d8)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000059 (
    .C(clk),
    .CE(ce),
    .D(sig000000af),
    .Q(sig0000017a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000005a (
    .C(clk),
    .CE(ce),
    .D(sig000000ab),
    .Q(sig000000e4)
  );
  MUXCY   blk0000005b (
    .CI(sig000000f3),
    .DI(sig00000002),
    .S(sig00000002),
    .O(sig000000f2)
  );
  MUXCY   blk0000005c (
    .CI(sig000000f4),
    .DI(sig00000002),
    .S(sig000000d5),
    .O(sig000000f3)
  );
  MUXCY   blk0000005d (
    .CI(sig000000f5),
    .DI(sig00000002),
    .S(sig000000d4),
    .O(sig000000f4)
  );
  MUXCY   blk0000005e (
    .CI(sig000000f6),
    .DI(sig00000002),
    .S(sig000000d3),
    .O(sig000000f5)
  );
  MUXCY   blk0000005f (
    .CI(sig000000f7),
    .DI(sig00000002),
    .S(sig000000d2),
    .O(sig000000f6)
  );
  MUXCY   blk00000060 (
    .CI(sig00000001),
    .DI(sig00000002),
    .S(sig000000d1),
    .O(sig000000f7)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000061 (
    .C(clk),
    .CE(ce),
    .D(sig000000f2),
    .Q(sig000000ed)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000062 (
    .C(clk),
    .CE(ce),
    .D(sig000000f3),
    .Q(sig000000ee)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000063 (
    .C(clk),
    .CE(ce),
    .D(sig000000f4),
    .Q(sig000000ec)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000064 (
    .C(clk),
    .CE(ce),
    .D(sig000000f5),
    .Q(sig000000ef)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000065 (
    .C(clk),
    .CE(ce),
    .D(sig000000f6),
    .Q(sig000000f0)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000066 (
    .C(clk),
    .CE(ce),
    .D(sig000000f7),
    .Q(sig000000f1)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000067 (
    .C(clk),
    .CE(ce),
    .D(sig000000d6),
    .Q(sig000000a7)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000068 (
    .C(clk),
    .CE(ce),
    .D(sig00000001),
    .Q(sig000000e6)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000069 (
    .C(clk),
    .CE(ce),
    .D(sig000000d9),
    .Q(sig000000e2)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000006a (
    .C(clk),
    .CE(ce),
    .D(sig000000da),
    .Q(sig000000e3)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000006b (
    .C(clk),
    .CE(ce),
    .D(sig000000db),
    .Q(sig000000e7)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000006c (
    .C(clk),
    .CE(ce),
    .D(sig000000dc),
    .Q(sig000000e5)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000006d (
    .C(clk),
    .CE(ce),
    .D(sig000000dd),
    .Q(sig000000e9)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000006e (
    .C(clk),
    .CE(ce),
    .D(sig000000de),
    .Q(sig000000ea)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000006f (
    .C(clk),
    .CE(ce),
    .D(sig000000df),
    .Q(sig000000eb)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000070 (
    .C(clk),
    .CE(ce),
    .D(sig000000e0),
    .Q(sig000000e8)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000071 (
    .C(clk),
    .CE(ce),
    .D(sig000000b0),
    .Q(sig0000017b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000072 (
    .C(clk),
    .CE(ce),
    .D(sig00000117),
    .Q(sig000000a6)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000073 (
    .C(clk),
    .CE(ce),
    .D(sig00000116),
    .Q(sig000000a5)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000074 (
    .C(clk),
    .CE(ce),
    .D(sig00000115),
    .Q(sig000000a4)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000075 (
    .C(clk),
    .CE(ce),
    .D(sig00000114),
    .Q(sig000000a3)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000076 (
    .C(clk),
    .CE(ce),
    .D(sig00000113),
    .Q(sig000000a2)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000077 (
    .C(clk),
    .CE(ce),
    .D(sig00000112),
    .Q(sig000000a1)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000078 (
    .C(clk),
    .CE(ce),
    .D(sig00000111),
    .Q(sig000000a0)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000079 (
    .C(clk),
    .CE(ce),
    .D(sig00000110),
    .Q(sig0000009f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000007a (
    .C(clk),
    .CE(ce),
    .D(sig0000010f),
    .Q(sig0000009e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000007b (
    .C(clk),
    .CE(ce),
    .D(sig0000010e),
    .Q(sig0000009d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000007c (
    .C(clk),
    .CE(ce),
    .D(sig0000010d),
    .Q(sig0000009c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000007d (
    .C(clk),
    .CE(ce),
    .D(sig0000010c),
    .Q(sig0000009b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000007e (
    .C(clk),
    .CE(ce),
    .D(sig0000010b),
    .Q(sig0000009a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000007f (
    .C(clk),
    .CE(ce),
    .D(sig0000010a),
    .Q(sig00000099)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000080 (
    .C(clk),
    .CE(ce),
    .D(sig00000109),
    .Q(sig00000098)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000081 (
    .C(clk),
    .CE(ce),
    .D(sig00000108),
    .Q(sig00000097)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000082 (
    .C(clk),
    .CE(ce),
    .D(sig00000107),
    .Q(sig00000096)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000083 (
    .C(clk),
    .CE(ce),
    .D(sig00000106),
    .Q(sig00000095)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000084 (
    .C(clk),
    .CE(ce),
    .D(sig00000105),
    .Q(sig00000094)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000085 (
    .C(clk),
    .CE(ce),
    .D(sig00000104),
    .Q(sig00000093)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000086 (
    .C(clk),
    .CE(ce),
    .D(sig00000103),
    .Q(sig00000092)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000087 (
    .C(clk),
    .CE(ce),
    .D(sig00000102),
    .Q(sig00000091)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000088 (
    .C(clk),
    .CE(ce),
    .D(sig00000101),
    .Q(sig00000090)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000089 (
    .C(clk),
    .CE(ce),
    .D(sig00000100),
    .Q(sig0000008f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000008a (
    .C(clk),
    .CE(ce),
    .D(sig000000ff),
    .Q(sig0000008e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000008b (
    .C(clk),
    .CE(ce),
    .D(sig000000fe),
    .Q(sig0000008d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000008c (
    .C(clk),
    .CE(ce),
    .D(sig000000fd),
    .Q(sig0000008c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000008d (
    .C(clk),
    .CE(ce),
    .D(sig000000fc),
    .Q(sig0000008b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000008e (
    .C(clk),
    .CE(ce),
    .D(sig000000fb),
    .Q(sig0000008a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000008f (
    .C(clk),
    .CE(ce),
    .D(sig000000fa),
    .Q(sig00000089)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000090 (
    .C(clk),
    .CE(ce),
    .D(sig000000f9),
    .Q(sig00000088)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000091 (
    .C(clk),
    .CE(ce),
    .D(sig000000f8),
    .Q(sig00000087)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000092 (
    .C(clk),
    .CE(ce),
    .D(sig00000137),
    .Q(sig00000179)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000093 (
    .C(clk),
    .CE(ce),
    .D(sig00000136),
    .Q(sig00000178)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000094 (
    .C(clk),
    .CE(ce),
    .D(sig00000135),
    .Q(sig00000177)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000095 (
    .C(clk),
    .CE(ce),
    .D(sig00000134),
    .Q(sig00000176)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000096 (
    .C(clk),
    .CE(ce),
    .D(sig00000133),
    .Q(sig00000175)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000097 (
    .C(clk),
    .CE(ce),
    .D(sig00000132),
    .Q(sig00000174)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000098 (
    .C(clk),
    .CE(ce),
    .D(sig00000131),
    .Q(sig00000173)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000099 (
    .C(clk),
    .CE(ce),
    .D(sig00000130),
    .Q(sig00000172)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000009a (
    .C(clk),
    .CE(ce),
    .D(sig0000012f),
    .Q(sig00000171)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000009b (
    .C(clk),
    .CE(ce),
    .D(sig0000012e),
    .Q(sig00000170)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000009c (
    .C(clk),
    .CE(ce),
    .D(sig0000012d),
    .Q(sig0000016f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000009d (
    .C(clk),
    .CE(ce),
    .D(sig0000012c),
    .Q(sig0000016e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000009e (
    .C(clk),
    .CE(ce),
    .D(sig0000012b),
    .Q(sig0000016d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000009f (
    .C(clk),
    .CE(ce),
    .D(sig0000012a),
    .Q(sig0000016c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000a0 (
    .C(clk),
    .CE(ce),
    .D(sig00000129),
    .Q(sig0000016b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000a1 (
    .C(clk),
    .CE(ce),
    .D(sig00000128),
    .Q(sig0000016a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000a2 (
    .C(clk),
    .CE(ce),
    .D(sig00000127),
    .Q(sig00000169)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000a3 (
    .C(clk),
    .CE(ce),
    .D(sig00000126),
    .Q(sig00000168)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000a4 (
    .C(clk),
    .CE(ce),
    .D(sig00000125),
    .Q(sig00000167)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000a5 (
    .C(clk),
    .CE(ce),
    .D(sig00000124),
    .Q(sig00000166)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000a6 (
    .C(clk),
    .CE(ce),
    .D(sig00000123),
    .Q(sig00000165)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000a7 (
    .C(clk),
    .CE(ce),
    .D(sig00000122),
    .Q(sig00000164)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000a8 (
    .C(clk),
    .CE(ce),
    .D(sig00000121),
    .Q(sig00000163)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000a9 (
    .C(clk),
    .CE(ce),
    .D(sig00000120),
    .Q(sig00000162)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000aa (
    .C(clk),
    .CE(ce),
    .D(sig0000011f),
    .Q(sig00000161)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000ab (
    .C(clk),
    .CE(ce),
    .D(sig0000011e),
    .Q(sig00000160)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000ac (
    .C(clk),
    .CE(ce),
    .D(sig0000011d),
    .Q(sig0000015f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000ad (
    .C(clk),
    .CE(ce),
    .D(sig0000011c),
    .Q(sig0000015e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000ae (
    .C(clk),
    .CE(ce),
    .D(sig0000011b),
    .Q(sig0000015d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000af (
    .C(clk),
    .CE(ce),
    .D(sig0000011a),
    .Q(sig0000015c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000b0 (
    .C(clk),
    .CE(ce),
    .D(sig00000119),
    .Q(sig0000015b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000b1 (
    .C(clk),
    .CE(ce),
    .D(sig00000118),
    .Q(sig0000015a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000b2 (
    .C(clk),
    .CE(ce),
    .D(sig00000157),
    .Q(sig0000019b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000b3 (
    .C(clk),
    .CE(ce),
    .D(sig00000156),
    .Q(sig0000019a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000b4 (
    .C(clk),
    .CE(ce),
    .D(sig00000155),
    .Q(sig00000199)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000b5 (
    .C(clk),
    .CE(ce),
    .D(sig00000154),
    .Q(sig00000198)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000b6 (
    .C(clk),
    .CE(ce),
    .D(sig00000153),
    .Q(sig00000197)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000b7 (
    .C(clk),
    .CE(ce),
    .D(sig00000152),
    .Q(sig00000196)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000b8 (
    .C(clk),
    .CE(ce),
    .D(sig00000151),
    .Q(sig00000195)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000b9 (
    .C(clk),
    .CE(ce),
    .D(sig00000150),
    .Q(sig00000194)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000ba (
    .C(clk),
    .CE(ce),
    .D(sig0000014f),
    .Q(sig00000193)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000bb (
    .C(clk),
    .CE(ce),
    .D(sig0000014e),
    .Q(sig00000192)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000bc (
    .C(clk),
    .CE(ce),
    .D(sig0000014d),
    .Q(sig00000191)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000bd (
    .C(clk),
    .CE(ce),
    .D(sig0000014c),
    .Q(sig00000190)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000be (
    .C(clk),
    .CE(ce),
    .D(sig0000014b),
    .Q(sig0000018f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000bf (
    .C(clk),
    .CE(ce),
    .D(sig0000014a),
    .Q(sig0000018e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000c0 (
    .C(clk),
    .CE(ce),
    .D(sig00000149),
    .Q(sig0000018d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000c1 (
    .C(clk),
    .CE(ce),
    .D(sig00000148),
    .Q(sig0000018c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000c2 (
    .C(clk),
    .CE(ce),
    .D(sig00000147),
    .Q(sig0000018b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000c3 (
    .C(clk),
    .CE(ce),
    .D(sig00000146),
    .Q(sig0000018a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000c4 (
    .C(clk),
    .CE(ce),
    .D(sig00000145),
    .Q(sig00000189)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000c5 (
    .C(clk),
    .CE(ce),
    .D(sig00000144),
    .Q(sig00000188)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000c6 (
    .C(clk),
    .CE(ce),
    .D(sig00000143),
    .Q(sig00000187)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000c7 (
    .C(clk),
    .CE(ce),
    .D(sig00000142),
    .Q(sig00000186)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000c8 (
    .C(clk),
    .CE(ce),
    .D(sig00000141),
    .Q(sig00000185)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000c9 (
    .C(clk),
    .CE(ce),
    .D(sig00000140),
    .Q(sig00000184)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000ca (
    .C(clk),
    .CE(ce),
    .D(sig0000013f),
    .Q(sig00000183)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000cb (
    .C(clk),
    .CE(ce),
    .D(sig0000013e),
    .Q(sig00000182)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000cc (
    .C(clk),
    .CE(ce),
    .D(sig0000013d),
    .Q(sig00000181)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000cd (
    .C(clk),
    .CE(ce),
    .D(sig0000013c),
    .Q(sig00000180)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000ce (
    .C(clk),
    .CE(ce),
    .D(sig0000013b),
    .Q(sig0000017f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000cf (
    .C(clk),
    .CE(ce),
    .D(sig0000013a),
    .Q(sig0000017e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000d0 (
    .C(clk),
    .CE(ce),
    .D(sig00000139),
    .Q(sig0000017d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000d1 (
    .C(clk),
    .CE(ce),
    .D(sig00000138),
    .Q(sig0000017c)
  );
  XORCY   blk000000d2 (
    .CI(sig0000019d),
    .LI(sig00000002),
    .O(NLW_blk000000d2_O_UNCONNECTED)
  );
  XORCY   blk000000d3 (
    .CI(sig0000019f),
    .LI(sig000001e4),
    .O(sig0000019c)
  );
  MUXCY   blk000000d4 (
    .CI(sig0000019f),
    .DI(sig00000002),
    .S(sig000001e4),
    .O(sig0000019d)
  );
  XORCY   blk000000d5 (
    .CI(sig000001a1),
    .LI(sig00000064),
    .O(sig0000019e)
  );
  MUXCY   blk000000d6 (
    .CI(sig000001a1),
    .DI(sig00000002),
    .S(sig00000064),
    .O(sig0000019f)
  );
  XORCY   blk000000d7 (
    .CI(sig000001a3),
    .LI(sig00000063),
    .O(sig000001a0)
  );
  MUXCY   blk000000d8 (
    .CI(sig000001a3),
    .DI(sig00000002),
    .S(sig00000063),
    .O(sig000001a1)
  );
  XORCY   blk000000d9 (
    .CI(sig000001a5),
    .LI(sig00000062),
    .O(sig000001a2)
  );
  MUXCY   blk000000da (
    .CI(sig000001a5),
    .DI(sig00000002),
    .S(sig00000062),
    .O(sig000001a3)
  );
  XORCY   blk000000db (
    .CI(sig000001a7),
    .LI(sig00000061),
    .O(sig000001a4)
  );
  MUXCY   blk000000dc (
    .CI(sig000001a7),
    .DI(sig00000002),
    .S(sig00000061),
    .O(sig000001a5)
  );
  XORCY   blk000000dd (
    .CI(sig000001a9),
    .LI(sig00000060),
    .O(sig000001a6)
  );
  MUXCY   blk000000de (
    .CI(sig000001a9),
    .DI(sig00000002),
    .S(sig00000060),
    .O(sig000001a7)
  );
  XORCY   blk000000df (
    .CI(sig000001ab),
    .LI(sig0000005f),
    .O(sig000001a8)
  );
  MUXCY   blk000000e0 (
    .CI(sig000001ab),
    .DI(sig00000002),
    .S(sig0000005f),
    .O(sig000001a9)
  );
  XORCY   blk000000e1 (
    .CI(sig000001ad),
    .LI(sig0000005e),
    .O(sig000001aa)
  );
  MUXCY   blk000000e2 (
    .CI(sig000001ad),
    .DI(sig00000002),
    .S(sig0000005e),
    .O(sig000001ab)
  );
  XORCY   blk000000e3 (
    .CI(sig000001af),
    .LI(sig0000005d),
    .O(sig000001ac)
  );
  MUXCY   blk000000e4 (
    .CI(sig000001af),
    .DI(sig00000002),
    .S(sig0000005d),
    .O(sig000001ad)
  );
  XORCY   blk000000e5 (
    .CI(sig000001b1),
    .LI(sig0000005c),
    .O(sig000001ae)
  );
  MUXCY   blk000000e6 (
    .CI(sig000001b1),
    .DI(sig00000002),
    .S(sig0000005c),
    .O(sig000001af)
  );
  XORCY   blk000000e7 (
    .CI(sig000001b3),
    .LI(sig0000005b),
    .O(sig000001b0)
  );
  MUXCY   blk000000e8 (
    .CI(sig000001b3),
    .DI(sig00000002),
    .S(sig0000005b),
    .O(sig000001b1)
  );
  XORCY   blk000000e9 (
    .CI(sig000001b5),
    .LI(sig0000005a),
    .O(sig000001b2)
  );
  MUXCY   blk000000ea (
    .CI(sig000001b5),
    .DI(sig00000002),
    .S(sig0000005a),
    .O(sig000001b3)
  );
  XORCY   blk000000eb (
    .CI(sig000001b7),
    .LI(sig00000059),
    .O(sig000001b4)
  );
  MUXCY   blk000000ec (
    .CI(sig000001b7),
    .DI(sig00000002),
    .S(sig00000059),
    .O(sig000001b5)
  );
  XORCY   blk000000ed (
    .CI(sig000001b9),
    .LI(sig00000058),
    .O(sig000001b6)
  );
  MUXCY   blk000000ee (
    .CI(sig000001b9),
    .DI(sig00000002),
    .S(sig00000058),
    .O(sig000001b7)
  );
  XORCY   blk000000ef (
    .CI(sig000001bb),
    .LI(sig00000057),
    .O(sig000001b8)
  );
  MUXCY   blk000000f0 (
    .CI(sig000001bb),
    .DI(sig00000002),
    .S(sig00000057),
    .O(sig000001b9)
  );
  XORCY   blk000000f1 (
    .CI(sig000001bd),
    .LI(sig00000056),
    .O(sig000001ba)
  );
  MUXCY   blk000000f2 (
    .CI(sig000001bd),
    .DI(sig00000002),
    .S(sig00000056),
    .O(sig000001bb)
  );
  XORCY   blk000000f3 (
    .CI(sig000001bf),
    .LI(sig00000055),
    .O(sig000001bc)
  );
  MUXCY   blk000000f4 (
    .CI(sig000001bf),
    .DI(sig00000002),
    .S(sig00000055),
    .O(sig000001bd)
  );
  XORCY   blk000000f5 (
    .CI(sig000001c1),
    .LI(sig00000054),
    .O(sig000001be)
  );
  MUXCY   blk000000f6 (
    .CI(sig000001c1),
    .DI(sig00000002),
    .S(sig00000054),
    .O(sig000001bf)
  );
  XORCY   blk000000f7 (
    .CI(sig000001c3),
    .LI(sig00000053),
    .O(sig000001c0)
  );
  MUXCY   blk000000f8 (
    .CI(sig000001c3),
    .DI(sig00000002),
    .S(sig00000053),
    .O(sig000001c1)
  );
  XORCY   blk000000f9 (
    .CI(sig000001c5),
    .LI(sig00000052),
    .O(sig000001c2)
  );
  MUXCY   blk000000fa (
    .CI(sig000001c5),
    .DI(sig00000002),
    .S(sig00000052),
    .O(sig000001c3)
  );
  XORCY   blk000000fb (
    .CI(sig000001c7),
    .LI(sig00000051),
    .O(sig000001c4)
  );
  MUXCY   blk000000fc (
    .CI(sig000001c7),
    .DI(sig00000002),
    .S(sig00000051),
    .O(sig000001c5)
  );
  XORCY   blk000000fd (
    .CI(sig000001c9),
    .LI(sig00000050),
    .O(sig000001c6)
  );
  MUXCY   blk000000fe (
    .CI(sig000001c9),
    .DI(sig00000002),
    .S(sig00000050),
    .O(sig000001c7)
  );
  XORCY   blk000000ff (
    .CI(sig000001cb),
    .LI(sig0000004f),
    .O(sig000001c8)
  );
  MUXCY   blk00000100 (
    .CI(sig000001cb),
    .DI(sig00000002),
    .S(sig0000004f),
    .O(sig000001c9)
  );
  XORCY   blk00000101 (
    .CI(sig000001cd),
    .LI(sig0000004e),
    .O(sig000001ca)
  );
  MUXCY   blk00000102 (
    .CI(sig000001cd),
    .DI(sig00000002),
    .S(sig0000004e),
    .O(sig000001cb)
  );
  XORCY   blk00000103 (
    .CI(sig000001cf),
    .LI(sig0000004d),
    .O(sig000001cc)
  );
  MUXCY   blk00000104 (
    .CI(sig000001cf),
    .DI(sig00000002),
    .S(sig0000004d),
    .O(sig000001cd)
  );
  XORCY   blk00000105 (
    .CI(sig000001d1),
    .LI(sig0000004c),
    .O(sig000001ce)
  );
  MUXCY   blk00000106 (
    .CI(sig000001d1),
    .DI(sig00000002),
    .S(sig0000004c),
    .O(sig000001cf)
  );
  XORCY   blk00000107 (
    .CI(sig000001d3),
    .LI(sig0000004b),
    .O(sig000001d0)
  );
  MUXCY   blk00000108 (
    .CI(sig000001d3),
    .DI(sig00000002),
    .S(sig0000004b),
    .O(sig000001d1)
  );
  XORCY   blk00000109 (
    .CI(sig000001d5),
    .LI(sig0000004a),
    .O(sig000001d2)
  );
  MUXCY   blk0000010a (
    .CI(sig000001d5),
    .DI(sig00000002),
    .S(sig0000004a),
    .O(sig000001d3)
  );
  XORCY   blk0000010b (
    .CI(sig000001d7),
    .LI(sig00000049),
    .O(sig000001d4)
  );
  MUXCY   blk0000010c (
    .CI(sig000001d7),
    .DI(sig00000002),
    .S(sig00000049),
    .O(sig000001d5)
  );
  XORCY   blk0000010d (
    .CI(sig000001d9),
    .LI(sig00000048),
    .O(sig000001d6)
  );
  MUXCY   blk0000010e (
    .CI(sig000001d9),
    .DI(sig00000002),
    .S(sig00000048),
    .O(sig000001d7)
  );
  XORCY   blk0000010f (
    .CI(sig000001db),
    .LI(sig00000047),
    .O(sig000001d8)
  );
  MUXCY   blk00000110 (
    .CI(sig000001db),
    .DI(sig00000002),
    .S(sig00000047),
    .O(sig000001d9)
  );
  XORCY   blk00000111 (
    .CI(sig000001dc),
    .LI(sig00000046),
    .O(sig000001da)
  );
  MUXCY   blk00000112 (
    .CI(sig000001dc),
    .DI(sig00000002),
    .S(sig00000046),
    .O(sig000001db)
  );
  XORCY   blk00000113 (
    .CI(sig00000001),
    .LI(sig0000001a),
    .O(NLW_blk00000113_O_UNCONNECTED)
  );
  MUXCY   blk00000114 (
    .CI(sig00000001),
    .DI(sig00000002),
    .S(sig0000001a),
    .O(sig000001dc)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000115 (
    .C(clk),
    .CE(ce),
    .D(sig0000019c),
    .Q(sig00000085)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000116 (
    .C(clk),
    .CE(ce),
    .D(sig0000019e),
    .Q(sig00000084)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000117 (
    .C(clk),
    .CE(ce),
    .D(sig000001a0),
    .Q(sig00000083)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000118 (
    .C(clk),
    .CE(ce),
    .D(sig000001a2),
    .Q(sig00000082)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000119 (
    .C(clk),
    .CE(ce),
    .D(sig000001a4),
    .Q(sig00000081)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000011a (
    .C(clk),
    .CE(ce),
    .D(sig000001a6),
    .Q(sig00000080)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000011b (
    .C(clk),
    .CE(ce),
    .D(sig000001a8),
    .Q(sig0000007f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000011c (
    .C(clk),
    .CE(ce),
    .D(sig000001aa),
    .Q(sig0000007e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000011d (
    .C(clk),
    .CE(ce),
    .D(sig000001ac),
    .Q(sig0000007d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000011e (
    .C(clk),
    .CE(ce),
    .D(sig000001ae),
    .Q(sig0000007c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000011f (
    .C(clk),
    .CE(ce),
    .D(sig000001b0),
    .Q(sig0000007b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000120 (
    .C(clk),
    .CE(ce),
    .D(sig000001b2),
    .Q(sig0000007a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000121 (
    .C(clk),
    .CE(ce),
    .D(sig000001b4),
    .Q(sig00000079)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000122 (
    .C(clk),
    .CE(ce),
    .D(sig000001b6),
    .Q(sig00000078)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000123 (
    .C(clk),
    .CE(ce),
    .D(sig000001b8),
    .Q(sig00000077)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000124 (
    .C(clk),
    .CE(ce),
    .D(sig000001ba),
    .Q(sig00000076)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000125 (
    .C(clk),
    .CE(ce),
    .D(sig000001bc),
    .Q(sig00000075)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000126 (
    .C(clk),
    .CE(ce),
    .D(sig000001be),
    .Q(sig00000074)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000127 (
    .C(clk),
    .CE(ce),
    .D(sig000001c0),
    .Q(sig00000073)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000128 (
    .C(clk),
    .CE(ce),
    .D(sig000001c2),
    .Q(sig00000072)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000129 (
    .C(clk),
    .CE(ce),
    .D(sig000001c4),
    .Q(sig00000071)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000012a (
    .C(clk),
    .CE(ce),
    .D(sig000001c6),
    .Q(sig00000070)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000012b (
    .C(clk),
    .CE(ce),
    .D(sig000001c8),
    .Q(sig0000006f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000012c (
    .C(clk),
    .CE(ce),
    .D(sig000001ca),
    .Q(sig0000006e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000012d (
    .C(clk),
    .CE(ce),
    .D(sig000001cc),
    .Q(sig0000006d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000012e (
    .C(clk),
    .CE(ce),
    .D(sig000001ce),
    .Q(sig0000006c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000012f (
    .C(clk),
    .CE(ce),
    .D(sig000001d0),
    .Q(sig0000006b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000130 (
    .C(clk),
    .CE(ce),
    .D(sig000001d2),
    .Q(sig0000006a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000131 (
    .C(clk),
    .CE(ce),
    .D(sig000001d4),
    .Q(sig00000069)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000132 (
    .C(clk),
    .CE(ce),
    .D(sig000001d6),
    .Q(sig00000068)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000133 (
    .C(clk),
    .CE(ce),
    .D(sig000001d8),
    .Q(sig00000067)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000134 (
    .C(clk),
    .CE(ce),
    .D(sig000001da),
    .Q(sig00000066)
  );
  LUT4 #(
    .INIT ( 16'h0001 ))
  blk00000135 (
    .I0(a[27]),
    .I1(a[28]),
    .I2(a[29]),
    .I3(a[30]),
    .O(sig00000018)
  );
  LUT5 #(
    .INIT ( 32'hAAAA88A8 ))
  blk00000136 (
    .I0(a[30]),
    .I1(a[28]),
    .I2(a[27]),
    .I3(sig00000003),
    .I4(a[29]),
    .O(sig00000026)
  );
  LUT5 #(
    .INIT ( 32'hA9AAA9A9 ))
  blk00000137 (
    .I0(a[30]),
    .I1(a[28]),
    .I2(a[29]),
    .I3(sig00000003),
    .I4(a[27]),
    .O(sig00000025)
  );
  LUT3 #(
    .INIT ( 8'h95 ))
  blk00000138 (
    .I0(a[26]),
    .I1(a[25]),
    .I2(a[24]),
    .O(sig00000021)
  );
  LUT4 #(
    .INIT ( 16'hC999 ))
  blk00000139 (
    .I0(a[26]),
    .I1(a[27]),
    .I2(a[24]),
    .I3(a[25]),
    .O(sig0000001f)
  );
  LUT4 #(
    .INIT ( 16'h0001 ))
  blk0000013a (
    .I0(a[15]),
    .I1(a[14]),
    .I2(a[12]),
    .I3(a[13]),
    .O(sig0000000d)
  );
  LUT4 #(
    .INIT ( 16'h3BC4 ))
  blk0000013b (
    .I0(sig000000a7),
    .I1(sig00000087),
    .I2(sig00000088),
    .I3(sig00000086),
    .O(sig0000001a)
  );
  LUT3 #(
    .INIT ( 8'h7F ))
  blk0000013c (
    .I0(a[24]),
    .I1(a[25]),
    .I2(a[26]),
    .O(sig00000003)
  );
  LUT5 #(
    .INIT ( 32'hF8080888 ))
  blk0000013d (
    .I0(sig00000085),
    .I1(sig00000065),
    .I2(ce),
    .I3(sig000000a8),
    .I4(sig000000a9),
    .O(sig00000019)
  );
  LUT4 #(
    .INIT ( 16'h0001 ))
  blk0000013e (
    .I0(a[19]),
    .I1(a[18]),
    .I2(a[17]),
    .I3(a[16]),
    .O(sig0000000e)
  );
  LUT3 #(
    .INIT ( 8'h01 ))
  blk0000013f (
    .I0(a[20]),
    .I1(a[21]),
    .I2(a[22]),
    .O(sig00000009)
  );
  LUT4 #(
    .INIT ( 16'h0001 ))
  blk00000140 (
    .I0(a[0]),
    .I1(a[1]),
    .I2(a[2]),
    .I3(a[3]),
    .O(sig0000000a)
  );
  LUT4 #(
    .INIT ( 16'h0001 ))
  blk00000141 (
    .I0(a[4]),
    .I1(a[5]),
    .I2(a[6]),
    .I3(a[7]),
    .O(sig0000000b)
  );
  LUT4 #(
    .INIT ( 16'h0001 ))
  blk00000142 (
    .I0(a[8]),
    .I1(a[9]),
    .I2(a[10]),
    .I3(a[11]),
    .O(sig0000000c)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000143 (
    .I0(sig00000088),
    .I1(sig00000086),
    .O(sig00000046)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000144 (
    .I0(sig00000092),
    .I1(sig00000086),
    .O(sig00000050)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000145 (
    .I0(sig00000093),
    .I1(sig00000086),
    .O(sig00000051)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000146 (
    .I0(sig00000094),
    .I1(sig00000086),
    .O(sig00000052)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000147 (
    .I0(sig00000095),
    .I1(sig00000086),
    .O(sig00000053)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000148 (
    .I0(sig00000096),
    .I1(sig00000086),
    .O(sig00000054)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000149 (
    .I0(sig00000097),
    .I1(sig00000086),
    .O(sig00000055)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk0000014a (
    .I0(sig00000098),
    .I1(sig00000086),
    .O(sig00000056)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk0000014b (
    .I0(sig00000099),
    .I1(sig00000086),
    .O(sig00000057)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk0000014c (
    .I0(sig0000009a),
    .I1(sig00000086),
    .O(sig00000058)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk0000014d (
    .I0(sig0000009b),
    .I1(sig00000086),
    .O(sig00000059)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk0000014e (
    .I0(sig00000089),
    .I1(sig00000086),
    .O(sig00000047)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk0000014f (
    .I0(sig0000009c),
    .I1(sig00000086),
    .O(sig0000005a)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000150 (
    .I0(sig0000009d),
    .I1(sig00000086),
    .O(sig0000005b)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000151 (
    .I0(sig0000009e),
    .I1(sig00000086),
    .O(sig0000005c)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000152 (
    .I0(sig0000009f),
    .I1(sig00000086),
    .O(sig0000005d)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000153 (
    .I0(sig000000a0),
    .I1(sig00000086),
    .O(sig0000005e)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000154 (
    .I0(sig000000a1),
    .I1(sig00000086),
    .O(sig0000005f)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000155 (
    .I0(sig000000a2),
    .I1(sig00000086),
    .O(sig00000060)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000156 (
    .I0(sig000000a3),
    .I1(sig00000086),
    .O(sig00000061)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000157 (
    .I0(sig000000a4),
    .I1(sig00000086),
    .O(sig00000062)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000158 (
    .I0(sig000000a5),
    .I1(sig00000086),
    .O(sig00000063)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000159 (
    .I0(sig0000008a),
    .I1(sig00000086),
    .O(sig00000048)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk0000015a (
    .I0(sig000000a6),
    .I1(sig00000086),
    .O(sig00000064)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk0000015b (
    .I0(sig0000008b),
    .I1(sig00000086),
    .O(sig00000049)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk0000015c (
    .I0(sig0000008c),
    .I1(sig00000086),
    .O(sig0000004a)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk0000015d (
    .I0(sig0000008d),
    .I1(sig00000086),
    .O(sig0000004b)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk0000015e (
    .I0(sig0000008e),
    .I1(sig00000086),
    .O(sig0000004c)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk0000015f (
    .I0(sig0000008f),
    .I1(sig00000086),
    .O(sig0000004d)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000160 (
    .I0(sig00000090),
    .I1(sig00000086),
    .O(sig0000004e)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000161 (
    .I0(sig00000091),
    .I1(sig00000086),
    .O(sig0000004f)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000162 (
    .I0(a[25]),
    .I1(a[24]),
    .O(sig00000020)
  );
  LUT4 #(
    .INIT ( 16'h8000 ))
  blk00000163 (
    .I0(a[27]),
    .I1(a[28]),
    .I2(a[29]),
    .I3(a[30]),
    .O(sig00000011)
  );
  LUT4 #(
    .INIT ( 16'h0001 ))
  blk00000164 (
    .I0(a[23]),
    .I1(a[24]),
    .I2(a[25]),
    .I3(a[26]),
    .O(sig00000017)
  );
  LUT5 #(
    .INIT ( 32'h011155FF ))
  blk00000165 (
    .I0(sig000000ca),
    .I1(sig000000cb),
    .I2(sig000000cc),
    .I3(sig000000ad),
    .I4(sig000000ae),
    .O(sig000000db)
  );
  LUT5 #(
    .INIT ( 32'h011155FF ))
  blk00000166 (
    .I0(sig000000c6),
    .I1(sig000000c7),
    .I2(sig000000c8),
    .I3(sig000000ad),
    .I4(sig000000ae),
    .O(sig000000dc)
  );
  LUT5 #(
    .INIT ( 32'h011155FF ))
  blk00000167 (
    .I0(sig000000c2),
    .I1(sig000000c3),
    .I2(sig000000c4),
    .I3(sig000000ad),
    .I4(sig000000ae),
    .O(sig000000dd)
  );
  LUT5 #(
    .INIT ( 32'h011155FF ))
  blk00000168 (
    .I0(sig000000be),
    .I1(sig000000bf),
    .I2(sig000000c0),
    .I3(sig000000ad),
    .I4(sig000000ae),
    .O(sig000000de)
  );
  LUT5 #(
    .INIT ( 32'h011155FF ))
  blk00000169 (
    .I0(sig000000ba),
    .I1(sig000000bb),
    .I2(sig000000bc),
    .I3(sig000000ad),
    .I4(sig000000ae),
    .O(sig000000df)
  );
  LUT5 #(
    .INIT ( 32'h011155FF ))
  blk0000016a (
    .I0(sig000000b6),
    .I1(sig000000b7),
    .I2(sig000000b8),
    .I3(sig000000ad),
    .I4(sig000000ae),
    .O(sig000000e0)
  );
  LUT4 #(
    .INIT ( 16'h0001 ))
  blk0000016b (
    .I0(sig000000b6),
    .I1(sig000000b7),
    .I2(sig000000b8),
    .I3(sig000000b9),
    .O(sig000000d1)
  );
  LUT4 #(
    .INIT ( 16'h0001 ))
  blk0000016c (
    .I0(sig000000ba),
    .I1(sig000000bb),
    .I2(sig000000bc),
    .I3(sig000000bd),
    .O(sig000000d2)
  );
  LUT4 #(
    .INIT ( 16'h0001 ))
  blk0000016d (
    .I0(sig000000be),
    .I1(sig000000bf),
    .I2(sig000000c0),
    .I3(sig000000c1),
    .O(sig000000d3)
  );
  LUT4 #(
    .INIT ( 16'h0001 ))
  blk0000016e (
    .I0(sig000000c2),
    .I1(sig000000c3),
    .I2(sig000000c4),
    .I3(sig000000c5),
    .O(sig000000d4)
  );
  LUT4 #(
    .INIT ( 16'h0001 ))
  blk0000016f (
    .I0(sig000000c6),
    .I1(sig000000c7),
    .I2(sig000000c8),
    .I3(sig000000c9),
    .O(sig000000d5)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk00000170 (
    .I0(sig00000158),
    .I1(sig00000159),
    .I2(sig0000016d),
    .I3(sig0000016f),
    .I4(sig0000016e),
    .I5(sig0000016c),
    .O(sig0000010a)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk00000171 (
    .I0(sig00000158),
    .I1(sig00000159),
    .I2(sig0000016f),
    .I3(sig00000171),
    .I4(sig00000170),
    .I5(sig0000016e),
    .O(sig0000010c)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk00000172 (
    .I0(sig00000158),
    .I1(sig00000159),
    .I2(sig0000016c),
    .I3(sig0000016e),
    .I4(sig0000016d),
    .I5(sig0000016b),
    .O(sig00000109)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk00000173 (
    .I0(sig00000158),
    .I1(sig00000159),
    .I2(sig0000016e),
    .I3(sig00000170),
    .I4(sig0000016f),
    .I5(sig0000016d),
    .O(sig0000010b)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk00000174 (
    .I0(sig00000158),
    .I1(sig00000159),
    .I2(sig0000016b),
    .I3(sig0000016d),
    .I4(sig0000016c),
    .I5(sig0000016a),
    .O(sig00000108)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk00000175 (
    .I0(sig00000158),
    .I1(sig00000159),
    .I2(sig0000016a),
    .I3(sig0000016c),
    .I4(sig0000016b),
    .I5(sig00000169),
    .O(sig00000107)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk00000176 (
    .I0(sig00000158),
    .I1(sig00000159),
    .I2(sig00000169),
    .I3(sig0000016b),
    .I4(sig0000016a),
    .I5(sig00000168),
    .O(sig00000106)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk00000177 (
    .I0(sig00000158),
    .I1(sig00000159),
    .I2(sig00000168),
    .I3(sig0000016a),
    .I4(sig00000169),
    .I5(sig00000167),
    .O(sig00000105)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk00000178 (
    .I0(sig00000158),
    .I1(sig00000159),
    .I2(sig00000167),
    .I3(sig00000169),
    .I4(sig00000168),
    .I5(sig00000166),
    .O(sig00000104)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk00000179 (
    .I0(sig00000158),
    .I1(sig00000159),
    .I2(sig00000166),
    .I3(sig00000168),
    .I4(sig00000167),
    .I5(sig00000165),
    .O(sig00000103)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk0000017a (
    .I0(sig00000158),
    .I1(sig00000159),
    .I2(sig00000165),
    .I3(sig00000167),
    .I4(sig00000166),
    .I5(sig00000164),
    .O(sig00000102)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk0000017b (
    .I0(sig00000158),
    .I1(sig00000159),
    .I2(sig00000164),
    .I3(sig00000166),
    .I4(sig00000165),
    .I5(sig00000163),
    .O(sig00000101)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk0000017c (
    .I0(sig00000158),
    .I1(sig00000159),
    .I2(sig00000163),
    .I3(sig00000165),
    .I4(sig00000164),
    .I5(sig00000162),
    .O(sig00000100)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk0000017d (
    .I0(sig00000158),
    .I1(sig00000159),
    .I2(sig00000162),
    .I3(sig00000164),
    .I4(sig00000163),
    .I5(sig00000161),
    .O(sig000000ff)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk0000017e (
    .I0(sig00000158),
    .I1(sig00000159),
    .I2(sig00000161),
    .I3(sig00000163),
    .I4(sig00000162),
    .I5(sig00000160),
    .O(sig000000fe)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk0000017f (
    .I0(sig00000158),
    .I1(sig00000159),
    .I2(sig00000160),
    .I3(sig00000162),
    .I4(sig00000161),
    .I5(sig0000015f),
    .O(sig000000fd)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk00000180 (
    .I0(sig00000158),
    .I1(sig00000159),
    .I2(sig00000177),
    .I3(sig00000179),
    .I4(sig00000178),
    .I5(sig00000176),
    .O(sig00000114)
  );
  LUT4 #(
    .INIT ( 16'h5410 ))
  blk00000181 (
    .I0(sig00000159),
    .I1(sig00000158),
    .I2(sig00000178),
    .I3(sig00000179),
    .O(sig00000116)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk00000182 (
    .I0(sig00000158),
    .I1(sig00000159),
    .I2(sig0000015e),
    .I3(sig00000160),
    .I4(sig0000015f),
    .I5(sig0000015d),
    .O(sig000000fb)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk00000183 (
    .I0(sig00000158),
    .I1(sig00000159),
    .I2(sig0000015c),
    .I3(sig0000015e),
    .I4(sig0000015d),
    .I5(sig0000015b),
    .O(sig000000f9)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk00000184 (
    .I0(sig00000158),
    .I1(sig00000159),
    .I2(sig0000015d),
    .I3(sig0000015f),
    .I4(sig0000015e),
    .I5(sig0000015c),
    .O(sig000000fa)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk00000185 (
    .I0(sig00000158),
    .I1(sig00000159),
    .I2(sig0000015b),
    .I3(sig0000015d),
    .I4(sig0000015c),
    .I5(sig0000015a),
    .O(sig000000f8)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk00000186 (
    .I0(sig00000158),
    .I1(sig00000159),
    .I2(sig00000176),
    .I3(sig00000178),
    .I4(sig00000177),
    .I5(sig00000175),
    .O(sig00000113)
  );
  LUT5 #(
    .INIT ( 32'h73625140 ))
  blk00000187 (
    .I0(sig00000159),
    .I1(sig00000158),
    .I2(sig00000178),
    .I3(sig00000177),
    .I4(sig00000179),
    .O(sig00000115)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk00000188 (
    .I0(sig00000158),
    .I1(sig00000159),
    .I2(sig00000175),
    .I3(sig00000177),
    .I4(sig00000176),
    .I5(sig00000174),
    .O(sig00000112)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk00000189 (
    .I0(sig00000158),
    .I1(sig00000159),
    .I2(sig00000174),
    .I3(sig00000176),
    .I4(sig00000175),
    .I5(sig00000173),
    .O(sig00000111)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk0000018a (
    .I0(sig00000158),
    .I1(sig00000159),
    .I2(sig00000173),
    .I3(sig00000175),
    .I4(sig00000174),
    .I5(sig00000172),
    .O(sig00000110)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk0000018b (
    .I0(sig00000158),
    .I1(sig00000159),
    .I2(sig00000172),
    .I3(sig00000174),
    .I4(sig00000173),
    .I5(sig00000171),
    .O(sig0000010f)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk0000018c (
    .I0(sig00000158),
    .I1(sig00000159),
    .I2(sig00000171),
    .I3(sig00000173),
    .I4(sig00000172),
    .I5(sig00000170),
    .O(sig0000010e)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk0000018d (
    .I0(sig00000158),
    .I1(sig00000159),
    .I2(sig00000170),
    .I3(sig00000172),
    .I4(sig00000171),
    .I5(sig0000016f),
    .O(sig0000010d)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk0000018e (
    .I0(sig00000158),
    .I1(sig00000159),
    .I2(sig0000015f),
    .I3(sig00000161),
    .I4(sig00000160),
    .I5(sig0000015e),
    .O(sig000000fc)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk0000018f (
    .I0(sig0000017a),
    .I1(sig0000017b),
    .I2(sig00000191),
    .I3(sig00000199),
    .I4(sig00000195),
    .I5(sig0000018d),
    .O(sig00000129)
  );
  LUT4 #(
    .INIT ( 16'h5410 ))
  blk00000190 (
    .I0(sig0000017b),
    .I1(sig0000017a),
    .I2(sig00000195),
    .I3(sig00000199),
    .O(sig00000131)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk00000191 (
    .I0(sig0000017a),
    .I1(sig0000017b),
    .I2(sig00000190),
    .I3(sig00000198),
    .I4(sig00000194),
    .I5(sig0000018c),
    .O(sig00000128)
  );
  LUT4 #(
    .INIT ( 16'h5410 ))
  blk00000192 (
    .I0(sig0000017b),
    .I1(sig0000017a),
    .I2(sig00000194),
    .I3(sig00000198),
    .O(sig00000130)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk00000193 (
    .I0(sig0000017a),
    .I1(sig0000017b),
    .I2(sig0000018f),
    .I3(sig00000197),
    .I4(sig00000193),
    .I5(sig0000018b),
    .O(sig00000127)
  );
  LUT5 #(
    .INIT ( 32'h73625140 ))
  blk00000194 (
    .I0(sig0000017b),
    .I1(sig0000017a),
    .I2(sig00000197),
    .I3(sig00000193),
    .I4(sig0000019b),
    .O(sig0000012f)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk00000195 (
    .I0(sig0000017a),
    .I1(sig0000017b),
    .I2(sig0000018e),
    .I3(sig00000196),
    .I4(sig00000192),
    .I5(sig0000018a),
    .O(sig00000126)
  );
  LUT5 #(
    .INIT ( 32'h73625140 ))
  blk00000196 (
    .I0(sig0000017b),
    .I1(sig0000017a),
    .I2(sig00000196),
    .I3(sig00000192),
    .I4(sig0000019a),
    .O(sig0000012e)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk00000197 (
    .I0(sig0000017a),
    .I1(sig0000017b),
    .I2(sig0000018d),
    .I3(sig00000195),
    .I4(sig00000191),
    .I5(sig00000189),
    .O(sig00000125)
  );
  LUT5 #(
    .INIT ( 32'h73625140 ))
  blk00000198 (
    .I0(sig0000017b),
    .I1(sig0000017a),
    .I2(sig00000195),
    .I3(sig00000191),
    .I4(sig00000199),
    .O(sig0000012d)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk00000199 (
    .I0(sig0000017a),
    .I1(sig0000017b),
    .I2(sig0000018c),
    .I3(sig00000194),
    .I4(sig00000190),
    .I5(sig00000188),
    .O(sig00000124)
  );
  LUT5 #(
    .INIT ( 32'h73625140 ))
  blk0000019a (
    .I0(sig0000017b),
    .I1(sig0000017a),
    .I2(sig00000194),
    .I3(sig00000190),
    .I4(sig00000198),
    .O(sig0000012c)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk0000019b (
    .I0(sig0000017a),
    .I1(sig0000017b),
    .I2(sig0000018b),
    .I3(sig00000193),
    .I4(sig0000018f),
    .I5(sig00000187),
    .O(sig00000123)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk0000019c (
    .I0(sig0000017a),
    .I1(sig0000017b),
    .I2(sig00000193),
    .I3(sig0000019b),
    .I4(sig00000197),
    .I5(sig0000018f),
    .O(sig0000012b)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk0000019d (
    .I0(sig0000017a),
    .I1(sig0000017b),
    .I2(sig00000189),
    .I3(sig00000191),
    .I4(sig0000018d),
    .I5(sig00000185),
    .O(sig00000121)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk0000019e (
    .I0(sig0000017a),
    .I1(sig0000017b),
    .I2(sig00000188),
    .I3(sig00000190),
    .I4(sig0000018c),
    .I5(sig00000184),
    .O(sig00000120)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk0000019f (
    .I0(sig0000017a),
    .I1(sig0000017b),
    .I2(sig00000187),
    .I3(sig0000018f),
    .I4(sig0000018b),
    .I5(sig00000183),
    .O(sig0000011f)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk000001a0 (
    .I0(sig0000017a),
    .I1(sig0000017b),
    .I2(sig00000180),
    .I3(sig00000188),
    .I4(sig00000184),
    .I5(sig0000017c),
    .O(sig00000118)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk000001a1 (
    .I0(sig0000017a),
    .I1(sig0000017b),
    .I2(sig00000192),
    .I3(sig0000019a),
    .I4(sig00000196),
    .I5(sig0000018e),
    .O(sig0000012a)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk000001a2 (
    .I0(sig0000017a),
    .I1(sig0000017b),
    .I2(sig0000018a),
    .I3(sig00000192),
    .I4(sig0000018e),
    .I5(sig00000186),
    .O(sig00000122)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk000001a3 (
    .I0(sig0000017a),
    .I1(sig0000017b),
    .I2(sig00000186),
    .I3(sig0000018e),
    .I4(sig0000018a),
    .I5(sig00000182),
    .O(sig0000011e)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk000001a4 (
    .I0(sig0000017a),
    .I1(sig0000017b),
    .I2(sig00000185),
    .I3(sig0000018d),
    .I4(sig00000189),
    .I5(sig00000181),
    .O(sig0000011d)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk000001a5 (
    .I0(sig0000017a),
    .I1(sig0000017b),
    .I2(sig00000184),
    .I3(sig0000018c),
    .I4(sig00000188),
    .I5(sig00000180),
    .O(sig0000011c)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk000001a6 (
    .I0(sig0000017a),
    .I1(sig0000017b),
    .I2(sig00000183),
    .I3(sig0000018b),
    .I4(sig00000187),
    .I5(sig0000017f),
    .O(sig0000011b)
  );
  LUT4 #(
    .INIT ( 16'h5410 ))
  blk000001a7 (
    .I0(sig0000017b),
    .I1(sig0000017a),
    .I2(sig00000197),
    .I3(sig0000019b),
    .O(sig00000133)
  );
  LUT4 #(
    .INIT ( 16'h5410 ))
  blk000001a8 (
    .I0(sig0000017b),
    .I1(sig0000017a),
    .I2(sig00000196),
    .I3(sig0000019a),
    .O(sig00000132)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk000001a9 (
    .I0(sig0000017a),
    .I1(sig0000017b),
    .I2(sig00000182),
    .I3(sig0000018a),
    .I4(sig00000186),
    .I5(sig0000017e),
    .O(sig0000011a)
  );
  LUT6 #(
    .INIT ( 64'hFD75B931EC64A820 ))
  blk000001aa (
    .I0(sig0000017a),
    .I1(sig0000017b),
    .I2(sig00000181),
    .I3(sig00000189),
    .I4(sig00000185),
    .I5(sig0000017d),
    .O(sig00000119)
  );
  LUT3 #(
    .INIT ( 8'h10 ))
  blk000001ab (
    .I0(sig00000159),
    .I1(sig00000158),
    .I2(sig00000179),
    .O(sig00000117)
  );
  LUT3 #(
    .INIT ( 8'h10 ))
  blk000001ac (
    .I0(sig0000017b),
    .I1(sig0000017a),
    .I2(sig00000198),
    .O(sig00000134)
  );
  LUT3 #(
    .INIT ( 8'h10 ))
  blk000001ad (
    .I0(sig0000017b),
    .I1(sig0000017a),
    .I2(sig00000199),
    .O(sig00000135)
  );
  LUT3 #(
    .INIT ( 8'h10 ))
  blk000001ae (
    .I0(sig0000017b),
    .I1(sig0000017a),
    .I2(sig0000019a),
    .O(sig00000136)
  );
  LUT3 #(
    .INIT ( 8'h10 ))
  blk000001af (
    .I0(sig0000017b),
    .I1(sig0000017a),
    .I2(sig0000019b),
    .O(sig00000137)
  );
  LUT2 #(
    .INIT ( 4'h8 ))
  blk000001b0 (
    .I0(sig000000b1),
    .I1(sig000000be),
    .O(sig00000138)
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  blk000001b1 (
    .I0(sig000000b1),
    .I1(sig000000b8),
    .I2(sig000000c8),
    .O(sig00000142)
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  blk000001b2 (
    .I0(sig000000b1),
    .I1(sig000000b9),
    .I2(sig000000c9),
    .O(sig00000143)
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  blk000001b3 (
    .I0(sig000000b1),
    .I1(sig000000ba),
    .I2(sig000000ca),
    .O(sig00000144)
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  blk000001b4 (
    .I0(sig000000b1),
    .I1(sig000000bb),
    .I2(sig000000cb),
    .O(sig00000145)
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  blk000001b5 (
    .I0(sig000000b1),
    .I1(sig000000bc),
    .I2(sig000000cc),
    .O(sig00000146)
  );
  LUT2 #(
    .INIT ( 4'hE ))
  blk000001b6 (
    .I0(sig000000b1),
    .I1(sig000000bd),
    .O(sig00000147)
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  blk000001b7 (
    .I0(sig000000be),
    .I1(sig000000b1),
    .O(sig00000148)
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  blk000001b8 (
    .I0(sig000000bf),
    .I1(sig000000b1),
    .O(sig00000149)
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  blk000001b9 (
    .I0(sig000000c0),
    .I1(sig000000b1),
    .O(sig0000014a)
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  blk000001ba (
    .I0(sig000000c1),
    .I1(sig000000b1),
    .O(sig0000014b)
  );
  LUT2 #(
    .INIT ( 4'h8 ))
  blk000001bb (
    .I0(sig000000b1),
    .I1(sig000000bf),
    .O(sig00000139)
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  blk000001bc (
    .I0(sig000000c2),
    .I1(sig000000b1),
    .O(sig0000014c)
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  blk000001bd (
    .I0(sig000000c3),
    .I1(sig000000b1),
    .O(sig0000014d)
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  blk000001be (
    .I0(sig000000c4),
    .I1(sig000000b1),
    .O(sig0000014e)
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  blk000001bf (
    .I0(sig000000c5),
    .I1(sig000000b1),
    .O(sig0000014f)
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  blk000001c0 (
    .I0(sig000000c6),
    .I1(sig000000b1),
    .O(sig00000150)
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  blk000001c1 (
    .I0(sig000000c7),
    .I1(sig000000b1),
    .O(sig00000151)
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  blk000001c2 (
    .I0(sig000000c8),
    .I1(sig000000b1),
    .O(sig00000152)
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  blk000001c3 (
    .I0(sig000000c9),
    .I1(sig000000b1),
    .O(sig00000153)
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  blk000001c4 (
    .I0(sig000000ca),
    .I1(sig000000b1),
    .O(sig00000154)
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  blk000001c5 (
    .I0(sig000000cb),
    .I1(sig000000b1),
    .O(sig00000155)
  );
  LUT2 #(
    .INIT ( 4'h8 ))
  blk000001c6 (
    .I0(sig000000b1),
    .I1(sig000000c0),
    .O(sig0000013a)
  );
  LUT2 #(
    .INIT ( 4'h2 ))
  blk000001c7 (
    .I0(sig000000cc),
    .I1(sig000000b1),
    .O(sig00000156)
  );
  LUT2 #(
    .INIT ( 4'h8 ))
  blk000001c8 (
    .I0(sig000000b1),
    .I1(sig000000c1),
    .O(sig0000013b)
  );
  LUT2 #(
    .INIT ( 4'h8 ))
  blk000001c9 (
    .I0(sig000000b1),
    .I1(sig000000c2),
    .O(sig0000013c)
  );
  LUT2 #(
    .INIT ( 4'h8 ))
  blk000001ca (
    .I0(sig000000b1),
    .I1(sig000000c3),
    .O(sig0000013d)
  );
  LUT2 #(
    .INIT ( 4'h8 ))
  blk000001cb (
    .I0(sig000000b1),
    .I1(sig000000c4),
    .O(sig0000013e)
  );
  LUT2 #(
    .INIT ( 4'h8 ))
  blk000001cc (
    .I0(sig000000b1),
    .I1(sig000000c5),
    .O(sig0000013f)
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  blk000001cd (
    .I0(sig000000b1),
    .I1(sig000000b6),
    .I2(sig000000c6),
    .O(sig00000140)
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  blk000001ce (
    .I0(sig000000b1),
    .I1(sig000000b7),
    .I2(sig000000c7),
    .O(sig00000141)
  );
  LUT6 #(
    .INIT ( 64'h0000000000000001 ))
  blk000001cf (
    .I0(a[8]),
    .I1(a[9]),
    .I2(a[7]),
    .I3(a[6]),
    .I4(a[5]),
    .I5(a[4]),
    .O(sig000001dd)
  );
  LUT6 #(
    .INIT ( 64'h0000000000000001 ))
  blk000001d0 (
    .I0(a[2]),
    .I1(a[3]),
    .I2(a[22]),
    .I3(a[21]),
    .I4(a[20]),
    .I5(a[1]),
    .O(sig000001de)
  );
  LUT3 #(
    .INIT ( 8'h01 ))
  blk000001d1 (
    .I0(a[10]),
    .I1(a[11]),
    .I2(a[0]),
    .O(sig000001df)
  );
  LUT5 #(
    .INIT ( 32'h80000000 ))
  blk000001d2 (
    .I0(sig0000000e),
    .I1(sig0000000d),
    .I2(sig000001de),
    .I3(sig000001df),
    .I4(sig000001dd),
    .O(sig0000001d)
  );
  LUT3 #(
    .INIT ( 8'hFE ))
  blk000001d3 (
    .I0(sig000000b4),
    .I1(sig000000b3),
    .I2(sig000000b2),
    .O(sig000001e0)
  );
  LUT6 #(
    .INIT ( 64'hFEFFFEEEF2FFF2A2 ))
  blk000001d4 (
    .I0(sig000000ce),
    .I1(sig000000aa),
    .I2(sig000000cd),
    .I3(sig000000b5),
    .I4(sig000001e0),
    .I5(sig00000014),
    .O(sig0000001b)
  );
  LUT2 #(
    .INIT ( 4'h8 ))
  blk000001d5 (
    .I0(sig000000aa),
    .I1(sig00000014),
    .O(sig000001e1)
  );
  LUT6 #(
    .INIT ( 64'h5555555500000004 ))
  blk000001d6 (
    .I0(sig000001e1),
    .I1(sig000000ce),
    .I2(sig000000b4),
    .I3(sig000000b3),
    .I4(sig000000b2),
    .I5(sig000000b5),
    .O(sig0000001c)
  );
  LUT5 #(
    .INIT ( 32'h0FFF7777 ))
  blk000001d7 (
    .I0(sig000000e5),
    .I1(sig000000ec),
    .I2(sig000000ee),
    .I3(sig000000e7),
    .I4(sig0000017a),
    .O(sig000001e2)
  );
  LUT5 #(
    .INIT ( 32'h8880BBB3 ))
  blk000001d8 (
    .I0(sig000000e6),
    .I1(sig000000e4),
    .I2(sig0000017a),
    .I3(sig000000ed),
    .I4(sig000001e2),
    .O(sig000000d9)
  );
  LUT5 #(
    .INIT ( 32'hEA404040 ))
  blk000001d9 (
    .I0(sig000000e4),
    .I1(sig000000eb),
    .I2(sig000000f1),
    .I3(sig000000e9),
    .I4(sig000000ef),
    .O(sig000001e3)
  );
  LUT6 #(
    .INIT ( 64'hFBBBEAAA51114000 ))
  blk000001da (
    .I0(sig0000017a),
    .I1(sig000000e4),
    .I2(sig000000ea),
    .I3(sig000000f0),
    .I4(sig000000e8),
    .I5(sig000001e3),
    .O(sig000000da)
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  blk000001db (
    .I0(sig00000086),
    .O(sig000001e4)
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  blk000001dc (
    .I0(sig000000e6),
    .O(sig000001e5)
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  blk000001dd (
    .I0(sig000000e6),
    .O(sig000001e6)
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  blk000001de (
    .I0(sig000000e3),
    .O(sig000001e7)
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  blk000001df (
    .I0(sig000000e2),
    .O(sig000001e8)
  );
  LUT6 #(
    .INIT ( 64'h5C4C5F5F5C4C5C4C ))
  blk000001e0 (
    .I0(sig000000a8),
    .I1(sig00000078),
    .I2(ce),
    .I3(sig000000a9),
    .I4(sig00000065),
    .I5(sig00000085),
    .O(sig00000039)
  );
  LUT6 #(
    .INIT ( 64'h5C4C5F5F5C4C5C4C ))
  blk000001e1 (
    .I0(sig000000a8),
    .I1(sig00000077),
    .I2(ce),
    .I3(sig000000a9),
    .I4(sig00000065),
    .I5(sig00000085),
    .O(sig00000038)
  );
  LUT6 #(
    .INIT ( 64'h5C4C5F5F5C4C5C4C ))
  blk000001e2 (
    .I0(sig000000a8),
    .I1(sig00000076),
    .I2(ce),
    .I3(sig000000a9),
    .I4(sig00000065),
    .I5(sig00000085),
    .O(sig00000037)
  );
  LUT6 #(
    .INIT ( 64'h5C4C5F5F5C4C5C4C ))
  blk000001e3 (
    .I0(sig000000a8),
    .I1(sig00000075),
    .I2(ce),
    .I3(sig000000a9),
    .I4(sig00000065),
    .I5(sig00000085),
    .O(sig00000036)
  );
  LUT6 #(
    .INIT ( 64'h5C4C5F5F5C4C5C4C ))
  blk000001e4 (
    .I0(sig000000a8),
    .I1(sig00000074),
    .I2(ce),
    .I3(sig000000a9),
    .I4(sig00000065),
    .I5(sig00000085),
    .O(sig00000035)
  );
  LUT6 #(
    .INIT ( 64'h5C4C5F5F5C4C5C4C ))
  blk000001e5 (
    .I0(sig000000a8),
    .I1(sig00000073),
    .I2(ce),
    .I3(sig000000a9),
    .I4(sig00000065),
    .I5(sig00000085),
    .O(sig00000034)
  );
  LUT6 #(
    .INIT ( 64'h5C4C5F5F5C4C5C4C ))
  blk000001e6 (
    .I0(sig000000a8),
    .I1(sig00000066),
    .I2(ce),
    .I3(sig000000a9),
    .I4(sig00000065),
    .I5(sig00000085),
    .O(sig00000027)
  );
  LUT6 #(
    .INIT ( 64'h5C4C5F5F5C4C5C4C ))
  blk000001e7 (
    .I0(sig000000a8),
    .I1(sig0000006f),
    .I2(ce),
    .I3(sig000000a9),
    .I4(sig00000065),
    .I5(sig00000085),
    .O(sig00000030)
  );
  LUT6 #(
    .INIT ( 64'h5C4C5F5F5C4C5C4C ))
  blk000001e8 (
    .I0(sig000000a8),
    .I1(sig00000072),
    .I2(ce),
    .I3(sig000000a9),
    .I4(sig00000065),
    .I5(sig00000085),
    .O(sig00000033)
  );
  LUT6 #(
    .INIT ( 64'h5C4C5F5F5C4C5C4C ))
  blk000001e9 (
    .I0(sig000000a8),
    .I1(sig0000006e),
    .I2(ce),
    .I3(sig000000a9),
    .I4(sig00000065),
    .I5(sig00000085),
    .O(sig0000002f)
  );
  LUT6 #(
    .INIT ( 64'h5C4C5F5F5C4C5C4C ))
  blk000001ea (
    .I0(sig000000a8),
    .I1(sig0000006d),
    .I2(ce),
    .I3(sig000000a9),
    .I4(sig00000065),
    .I5(sig00000085),
    .O(sig0000002e)
  );
  LUT6 #(
    .INIT ( 64'h5C4C5F5F5C4C5C4C ))
  blk000001eb (
    .I0(sig000000a8),
    .I1(sig0000006c),
    .I2(ce),
    .I3(sig000000a9),
    .I4(sig00000065),
    .I5(sig00000085),
    .O(sig0000002d)
  );
  LUT6 #(
    .INIT ( 64'h5C4C5F5F5C4C5C4C ))
  blk000001ec (
    .I0(sig000000a8),
    .I1(sig0000006b),
    .I2(ce),
    .I3(sig000000a9),
    .I4(sig00000065),
    .I5(sig00000085),
    .O(sig0000002c)
  );
  LUT6 #(
    .INIT ( 64'h5C4C5F5F5C4C5C4C ))
  blk000001ed (
    .I0(sig000000a8),
    .I1(sig0000006a),
    .I2(ce),
    .I3(sig000000a9),
    .I4(sig00000065),
    .I5(sig00000085),
    .O(sig0000002b)
  );
  LUT6 #(
    .INIT ( 64'h5C4C5F5F5C4C5C4C ))
  blk000001ee (
    .I0(sig000000a8),
    .I1(sig00000069),
    .I2(ce),
    .I3(sig000000a9),
    .I4(sig00000065),
    .I5(sig00000085),
    .O(sig0000002a)
  );
  LUT6 #(
    .INIT ( 64'h5C4C5F5F5C4C5C4C ))
  blk000001ef (
    .I0(sig000000a8),
    .I1(sig00000084),
    .I2(ce),
    .I3(sig000000a9),
    .I4(sig00000065),
    .I5(sig00000085),
    .O(sig00000045)
  );
  LUT6 #(
    .INIT ( 64'h5C4C5F5F5C4C5C4C ))
  blk000001f0 (
    .I0(sig000000a8),
    .I1(sig00000068),
    .I2(ce),
    .I3(sig000000a9),
    .I4(sig00000065),
    .I5(sig00000085),
    .O(sig00000029)
  );
  LUT6 #(
    .INIT ( 64'h5C4C5F5F5C4C5C4C ))
  blk000001f1 (
    .I0(sig000000a8),
    .I1(sig00000083),
    .I2(ce),
    .I3(sig000000a9),
    .I4(sig00000065),
    .I5(sig00000085),
    .O(sig00000044)
  );
  LUT6 #(
    .INIT ( 64'h5C4C5F5F5C4C5C4C ))
  blk000001f2 (
    .I0(sig000000a8),
    .I1(sig00000082),
    .I2(ce),
    .I3(sig000000a9),
    .I4(sig00000065),
    .I5(sig00000085),
    .O(sig00000043)
  );
  LUT6 #(
    .INIT ( 64'h5C4C5F5F5C4C5C4C ))
  blk000001f3 (
    .I0(sig000000a8),
    .I1(sig00000071),
    .I2(ce),
    .I3(sig000000a9),
    .I4(sig00000065),
    .I5(sig00000085),
    .O(sig00000032)
  );
  LUT6 #(
    .INIT ( 64'h5C4C5F5F5C4C5C4C ))
  blk000001f4 (
    .I0(sig000000a8),
    .I1(sig00000081),
    .I2(ce),
    .I3(sig000000a9),
    .I4(sig00000065),
    .I5(sig00000085),
    .O(sig00000042)
  );
  LUT6 #(
    .INIT ( 64'h5C4C5F5F5C4C5C4C ))
  blk000001f5 (
    .I0(sig000000a8),
    .I1(sig00000080),
    .I2(ce),
    .I3(sig000000a9),
    .I4(sig00000065),
    .I5(sig00000085),
    .O(sig00000041)
  );
  LUT6 #(
    .INIT ( 64'h5C4C5F5F5C4C5C4C ))
  blk000001f6 (
    .I0(sig000000a8),
    .I1(sig0000007f),
    .I2(ce),
    .I3(sig000000a9),
    .I4(sig00000065),
    .I5(sig00000085),
    .O(sig00000040)
  );
  LUT6 #(
    .INIT ( 64'h5C4C5F5F5C4C5C4C ))
  blk000001f7 (
    .I0(sig000000a8),
    .I1(sig0000007e),
    .I2(ce),
    .I3(sig000000a9),
    .I4(sig00000065),
    .I5(sig00000085),
    .O(sig0000003f)
  );
  LUT6 #(
    .INIT ( 64'h5C4C5F5F5C4C5C4C ))
  blk000001f8 (
    .I0(sig000000a8),
    .I1(sig0000007d),
    .I2(ce),
    .I3(sig000000a9),
    .I4(sig00000065),
    .I5(sig00000085),
    .O(sig0000003e)
  );
  LUT6 #(
    .INIT ( 64'h5C4C5F5F5C4C5C4C ))
  blk000001f9 (
    .I0(sig000000a8),
    .I1(sig0000007c),
    .I2(ce),
    .I3(sig000000a9),
    .I4(sig00000065),
    .I5(sig00000085),
    .O(sig0000003d)
  );
  LUT6 #(
    .INIT ( 64'h5C4C5F5F5C4C5C4C ))
  blk000001fa (
    .I0(sig000000a8),
    .I1(sig0000007b),
    .I2(ce),
    .I3(sig000000a9),
    .I4(sig00000065),
    .I5(sig00000085),
    .O(sig0000003c)
  );
  LUT6 #(
    .INIT ( 64'h5C4C5F5F5C4C5C4C ))
  blk000001fb (
    .I0(sig000000a8),
    .I1(sig0000007a),
    .I2(ce),
    .I3(sig000000a9),
    .I4(sig00000065),
    .I5(sig00000085),
    .O(sig0000003b)
  );
  LUT6 #(
    .INIT ( 64'h5C4C5F5F5C4C5C4C ))
  blk000001fc (
    .I0(sig000000a8),
    .I1(sig00000067),
    .I2(ce),
    .I3(sig000000a9),
    .I4(sig00000065),
    .I5(sig00000085),
    .O(sig00000028)
  );
  LUT6 #(
    .INIT ( 64'h5C4C5F5F5C4C5C4C ))
  blk000001fd (
    .I0(sig000000a8),
    .I1(sig00000079),
    .I2(ce),
    .I3(sig000000a9),
    .I4(sig00000065),
    .I5(sig00000085),
    .O(sig0000003a)
  );
  LUT6 #(
    .INIT ( 64'h5C4C5F5F5C4C5C4C ))
  blk000001fe (
    .I0(sig000000a8),
    .I1(sig00000070),
    .I2(ce),
    .I3(sig000000a9),
    .I4(sig00000065),
    .I5(sig00000085),
    .O(sig00000031)
  );
  LUT5 #(
    .INIT ( 32'h6AAAAAAA ))
  blk000001ff (
    .I0(a[28]),
    .I1(a[24]),
    .I2(a[25]),
    .I3(a[26]),
    .I4(a[27]),
    .O(sig00000023)
  );
  LUT6 #(
    .INIT ( 64'h3666666666666666 ))
  blk00000200 (
    .I0(a[28]),
    .I1(a[29]),
    .I2(a[27]),
    .I3(a[24]),
    .I4(a[25]),
    .I5(a[26]),
    .O(sig00000024)
  );
  LUT4 #(
    .INIT ( 16'h9555 ))
  blk00000201 (
    .I0(a[27]),
    .I1(a[24]),
    .I2(a[25]),
    .I3(a[26]),
    .O(sig00000022)
  );
  LUT4 #(
    .INIT ( 16'h8000 ))
  blk00000202 (
    .I0(a[23]),
    .I1(a[24]),
    .I2(a[25]),
    .I3(a[26]),
    .O(sig00000010)
  );
  LUT3 #(
    .INIT ( 8'h6A ))
  blk00000203 (
    .I0(a[26]),
    .I1(a[25]),
    .I2(a[24]),
    .O(sig0000001e)
  );
  INV   blk00000204 (
    .I(a[23]),
    .O(sig0000000f)
  );
  INV   blk00000205 (
    .I(sig000000b1),
    .O(sig00000157)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000206 (
    .A0(sig00000001),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(ce),
    .CLK(clk),
    .D(sig000000cf),
    .Q(sig000001e9),
    .Q15(NLW_blk00000206_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000207 (
    .C(clk),
    .CE(ce),
    .D(sig000001e9),
    .Q(sig000000a8)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000208 (
    .A0(sig00000001),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(ce),
    .CLK(clk),
    .D(sig000000cd),
    .Q(sig000001ea),
    .Q15(NLW_blk00000208_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000209 (
    .C(clk),
    .CE(ce),
    .D(sig000001ea),
    .Q(sig00000086)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk0000020a (
    .A0(sig00000001),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(ce),
    .CLK(clk),
    .D(sig000000d0),
    .Q(sig000001eb),
    .Q15(NLW_blk0000020a_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000020b (
    .C(clk),
    .CE(ce),
    .D(sig000001eb),
    .Q(sig000000a9)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk0000020c (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(ce),
    .CLK(clk),
    .D(sig000000ae),
    .Q(sig000001ec),
    .Q15(NLW_blk0000020c_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000020d (
    .C(clk),
    .CE(ce),
    .D(sig000001ec),
    .Q(sig00000159)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk0000020e (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(ce),
    .CLK(clk),
    .D(sig000000ac),
    .Q(sig000001ed),
    .Q15(NLW_blk0000020e_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000020f (
    .C(clk),
    .CE(ce),
    .D(sig000001ed),
    .Q(sig000000e1)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000210 (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(ce),
    .CLK(clk),
    .D(sig000000ad),
    .Q(sig000001ee),
    .Q15(NLW_blk00000210_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000211 (
    .C(clk),
    .CE(ce),
    .D(sig000001ee),
    .Q(sig00000158)
  );
endmodule