module amiq_eth_ve_top;
	initial begin
		run_test();
	end
endmodule