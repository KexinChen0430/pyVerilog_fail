module delay (in, out);
  input  in;
  output out;
  assign out = in;
  specify
    (in => out) = (600,600);
  endspecify
endmodule