module  rtfc71e(
   sys_clk,
   rst_n,
   pse18cc,
   ls35987,
   jrc662,
   zk63316,
   lf198b2,
   yxcc596,
   os62cb4,
   fp165a1,
   xyb2d0e,
   ba96872,
   wlb4393,
   uxa1c9c,
   vke4e4,
   ay5cd66,
   `ifdef EN_VC0
      hq93919,
      ri9c8cb,
      tue465a,
   `endif
   `ifdef EN_VC1
      sj232d3,
      hd1969c,
      uicb4e7,
   `endif
   `ifdef EN_VC2
      pf5a739,
      end39ce,
      tw9ce75,
   `endif
   `ifdef EN_VC3
      kde73aa,
      ux39d54,
      kqceaa5,
   `endif
   `ifdef EN_VC4
      ip75528,
      ntaa944,
      al54a27,
   `endif
   `ifdef EN_VC5
      lfa513c,
      hd289e7,
      al44f3e,
   `endif
   `ifdef EN_VC6
      hd279f5,
      an3cfaf,
      ipe7d7d,
   `endif
   `ifdef EN_VC7
      gq3ebed,
      ykf5f68,
      phafb41,
   `endif
   os7da0f,
   tx_pmtype,
   ww683cd,
   tx_vsd_data,
   yx4e2a2,
   al7fcee,
   xw69c54,
   jce1a71,
   zx74783,
   qia3c1e,
   tw1e0f1,
   icf078a,
   ls83c50,
   ls1e282,
   yzae707,
   fa7383c,
   ng9c1e2,
   qge0f13,
   qv7898,
   ba250d2,
   wwf5804,
   vk30204,
   wyac021,
   uv60109,
   ym84d,
   pu4269,
   qi2134a,
   bn169d7,
   jpd27c8,
   do93e46,
   mt9f233,
   rib82be,
   icc15f2,
   do993fe,
   qtc9ff3,
   xjc264f,
   jr1327f,
   cm46737
   );
`ifdef LW1
parameter LANE_WIDTH = 1 ;
`else
`ifdef LW2
parameter LANE_WIDTH = 2 ;
`else
`ifdef LW4
parameter LANE_WIDTH = 4 ;
`else
parameter LANE_WIDTH = 1 ;
`endif
`endif
`endif
parameter D_WIDTH = 16 ;
parameter K27_7 = 8'hFB ;
parameter K28_0 = 8'h1C ;
parameter K28_2 = 8'h5C ;
parameter K28_3 = 8'h7C ;
parameter K28_5 = 8'hBC ;
parameter K29_7 = 8'hFD ;
parameter K30_7 = 8'hFE ;
parameter K23_7 = 8'hF7 ;
parameter K28_1 = 8'h3C ;
parameter D5_2  = 8'h45 ;
parameter D10_2 = 8'h4A ;
parameter D21_5 = 8'hB5 ;
parameter D26_5 = 8'hBA ;
parameter COM = K28_5 ;
parameter STP = K27_7 ;
parameter SDP = K28_2 ;
parameter END = K29_7 ;
parameter EDB = K30_7 ;
parameter SKP = K28_0 ;
parameter IDL = K28_3 ;
parameter PAD = K23_7 ;
parameter FTS = K28_1 ;
parameter OS_WIDTH      = 4 ;
parameter OS_T1_LIP_LAP = 4'd0 ;
parameter OS_T2_LIP_LAP = 4'd1 ;
parameter OS_COMPLI     = 4'd2 ;
parameter OS_T1         = 4'd3 ;
parameter OS_T2         = 4'd4 ;
parameter OS_IDLE       = 4'd5 ;
parameter OS_EIDLE      = 4'd6 ;
parameter OS_NFTS       = 4'd7 ;
parameter OS_BEACON     = 4'd8 ;
parameter DSM_WIDTH    = 2 ;
parameter PSM_WIDTH    = 2 ;
parameter RSM_WIDTH    = 2 ;
parameter L0SM_WIDTH   = 2 ;
parameter L0sTSM_WIDTH = 2 ;
parameter L0sRSM_WIDTH = 2 ;
parameter L1SM_WIDTH   = 1 ;
parameter L2SM_WIDTH   = 1 ;
parameter DISM_WIDTH   = 2 ;
parameter LBSM_WIDTH   = 2 ;
parameter HRSM_WIDTH   = 1 ;
parameter CFGSM_WIDTH  = 2 ;
parameter MSM_WIDTH    = 3 ;
parameter DETECT    = 4'd0 ;
parameter POLLING   = 4'd1 ;
parameter CONFIG    = 4'd2 ;
parameter L0        = 4'd3 ;
parameter L0s       = 4'd4 ;
parameter L1        = 4'd5 ;
parameter L2        = 4'd6 ;
parameter RECOVERY  = 4'd7 ;
parameter LOOPBACK  = 4'd8 ;
parameter HOTRST    = 4'd9 ;
parameter DISABLED  = 4'd10 ;
`ifdef VC1
parameter FADDR = 3 ;
`else
`ifdef VC2
parameter FADDR = 3 ;
`else
`ifdef VC3
parameter FADDR = 5 ;
`else
`ifdef VC4
parameter FADDR = 5 ;
`else
parameter FADDR = 6 ;
`endif
`endif
`endif
`endif
input                     sys_clk;
input                     rst_n;
input  [13:0]             pse18cc;
input                     ls35987;
input                     jrc662;
input                     zk63316;
input                     lf198b2;
input  [2:0]              yxcc596;
input  [1:0]              os62cb4;
input                     fp165a1;
input  [2:0]              xyb2d0e;
input  [1:0]              ba96872;
input  [`NUM_VC -1:0]     wlb4393;
input  [`NUM_VC -1:0]     uxa1c9c;
input  [`NUM_VC -1:0]     vke4e4;
input [(`NUM_VC*3)-1:0]   ay5cd66;
`ifdef EN_VC0
input  [23:0]             hq93919;
input  [23:0]             ri9c8cb;
input  [23:0]             tue465a;
`endif
`ifdef EN_VC1
input  [23:0]             sj232d3;
input  [23:0]             hd1969c;
input  [23:0]             uicb4e7;
`endif
`ifdef EN_VC2
input  [23:0]             pf5a739;
input  [23:0]             end39ce;
input  [23:0]             tw9ce75;
`endif
`ifdef EN_VC3
input  [23:0]             kde73aa;
input  [23:0]             ux39d54;
input  [23:0]             kqceaa5;
`endif
`ifdef EN_VC4
input  [23:0]             ip75528;
input  [23:0]             ntaa944;
input  [23:0]             al54a27;
`endif
`ifdef EN_VC5
input  [23:0]             lfa513c;
input  [23:0]             hd289e7;
input  [23:0]             al44f3e;
`endif
`ifdef EN_VC6
input  [23:0]             hd279f5;
input  [23:0]             an3cfaf;
input  [23:0]             ipe7d7d;
`endif
`ifdef EN_VC7
input  [23:0]             gq3ebed;
input  [23:0]             ykf5f68;
input  [23:0]             phafb41;
`endif
input                     os7da0f;
input  [2:0]              tx_pmtype;
input                     ww683cd;
input  [23:0]             tx_vsd_data;
input                     yx4e2a2;
input                     al7fcee;
input                     xw69c54;
input  [11:0]             jce1a71;
input                     zx74783;
input                     qia3c1e;
input  [2:0]              tw1e0f1;
input                     icf078a;
input  [1:0]              ls83c50;
input  [`NUM_VC -1:0]     ls1e282;
input  [15:0]             yzae707;
input                     fa7383c;
input                     ng9c1e2;
input                     qge0f13;
input                     qv7898;
output [FADDR:0]          ba250d2;
output [15:0]             wwf5804;
output                    vk30204;
output                    wyac021;
output                    uv60109;
output                    ym84d;
output                    pu4269;
output                    qi2134a;
output                    bn169d7;
output [`NUM_VC -1:0]     jpd27c8;
output [`NUM_VC -1:0]     do93e46;
output [`NUM_VC -1:0]     mt9f233;
output                    rib82be;
output                    icc15f2;
output                    do993fe;
output                    qtc9ff3;
output                    xjc264f;
output                    jr1327f;
output                    cm46737;
wire                      an3c4c4;
wire                      ene2624;
wire   [3:0]              mec4930;
wire                      wy24981;
wire                      zz13124;
wire                      aa98926;
wire   [15:0]             ks24c08;
wire   [`NUM_VC -1:0]     jpd27c8;
wire   [`NUM_VC -1:0]     do93e46;
wire   [`NUM_VC -1:0]     mt9f233;
wire                      xjc264f;
wire                      jr1327f;
wire                      cm46737;
wire                      rib82be;
wire                      icc15f2;
wire                      do993fe;
wire                      qtc9ff3;
reg                       lqe4a1a;
reg                       byd5d12;
reg                       sjae892;
reg                       pf74495;
reg   [11:0]              pua24ae;
reg                       ir12572;
reg   [2:0]               uk92b94;
reg                       sj95ca1;
reg    [23:0]             yzae50c;
reg                       ea72864;
reg                       hd94320;
wire                      sj23425;
wire                      ec1a12c;
wire   [31:0]             tud0960;
wire   [31:0]             hd84b02;
wire                      gqb98bf;
wire                      sj3cfd4;
wire                      wje7ea5;
wire                      wlb4ebf;
wire                      xya75fd;
`ifdef EN_VC0
`endif
`ifdef EN_VC1
`endif
`ifdef EN_VC2
`endif
`ifdef EN_VC3
`endif
`ifdef EN_VC4
`endif
`ifdef EN_VC5
`endif
`ifdef EN_VC6
`endif
`ifdef EN_VC7
`endif
reg [13 : 0] ldd748a;
reg bl64b01;
reg vxba456;
reg vvd22b7;
reg xl915be;
reg [2 : 0] qv8adf7;
reg [1 : 0] cm56fbc;
reg dob7de1;
reg [2 : 0] yzbef0a;
reg [1 : 0] off7854;
reg [`NUM_VC - 1 : 0] gqbc2a4;
reg [`NUM_VC - 1 : 0] zke1520;
reg [`NUM_VC - 1 : 0] mga903;
reg [(`NUM_VC * 3) - 1 : 0] cz75325;
reg uxa40c4;
reg [2 : 0] ip7f3bf;
reg ph312b;
reg [23 : 0] wl1895f;
reg ldd88f4;
reg wwc47a6;
reg co2bf0b;
reg [11 : 0] rt5f859;
reg zxfc2cf;
reg vie167e;
reg [2 : 0] hqb3f3;
reg me59f9b;
reg [1 : 0] facfcd8;
reg [`NUM_VC - 1 : 0] vv7e6c2;
reg [15 : 0] wyb31e1;
reg wy98f09;
reg jpc7848;
reg wl3c246;
reg xwe1234;
reg zz91a3;
reg xw48d1e;
reg [3 : 0] oua3cc0;
reg do1e601;
reg kq468f3;
reg co34798;
reg [15 : 0] nrf300a;
reg vvd85fe;
reg ngade42;
reg wj6f212;
reg ps79094;
reg [11 : 0] vvc84a2;
reg rg42516;
reg [2 : 0] mt128b3;
reg hd9459d;
reg [23 : 0] ria2cef;
reg db1677b;
reg gqb3bde;
reg do9918e;
reg rtc8c73;
reg [31 : 0] os4639f;
reg [31 : 0] mg31cf9;
reg uif0030;
reg ep80180;
reg gqc04;
reg vvf3617;
reg rv9b0bf;
reg [2047:0] necf6c2;
wire [59:0] ld7b613;
`ifdef LW1
`else
`ifdef LW2
`else
`ifdef LW4
`else
`endif
`endif
`endif
`ifdef VC1
`else
`ifdef VC2
`else
`ifdef VC3
`else
`ifdef VC4
`else
`endif
`endif
`endif
`endif
`ifdef EN_VC0
`endif
`ifdef EN_VC1
`endif
`ifdef EN_VC2
`endif
`ifdef EN_VC3
`endif
`ifdef EN_VC4
`endif
`ifdef EN_VC5
`endif
`ifdef EN_VC6
`endif
`ifdef EN_VC7
`endif
`ifdef EN_VC0
`endif
`ifdef EN_VC1
`endif
`ifdef EN_VC2
`endif
`ifdef EN_VC3
`endif
`ifdef EN_VC4
`endif
`ifdef EN_VC5
`endif
`ifdef EN_VC6
`endif
`ifdef EN_VC7
`endif
localparam qgdb09f = 60,nrd84f8 = 32'hfdffd42b;
localparam [31:0] thc27c7 = nrd84f8;
localparam mt9f1ff = nrd84f8 & 4'hf;
localparam [11:0] fnc7fe5 = 'h7ff;
wire  [(1 << mt9f1ff)  -1:0] suff972;
reg    [qgdb09f-1:0] cme5c87;
reg [mt9f1ff-1:0] qg721c0 [0:1];
reg [mt9f1ff-1:0] ym8700c;
reg rv38061;
integer jcc030e;
integer vk1872;
`ifdef LW1
`else
`ifdef LW2
`else
`ifdef LW4
`else
`endif
`endif
`endif
`ifdef VC1
`else
`ifdef VC2
`else
`ifdef VC3
`else
`ifdef VC4
`else
`endif
`endif
`endif
`endif
`ifdef EN_VC0
`endif
`ifdef EN_VC1
`endif
`ifdef EN_VC2
`endif
`ifdef EN_VC3
`endif
`ifdef EN_VC4
`endif
`ifdef EN_VC5
`endif
`ifdef EN_VC6
`endif
`ifdef EN_VC7
`endif
`ifdef EN_VC0
`endif
`ifdef EN_VC1
`endif
`ifdef EN_VC2
`endif
`ifdef EN_VC3
`endif
`ifdef EN_VC4
`endif
`ifdef EN_VC5
`endif
`ifdef EN_VC6
`endif
`ifdef EN_VC7
`endif
`ifdef LW1
`else
`ifdef LW2
`else
`ifdef LW4
`else
`endif
`endif
`endif
`ifdef VC1
`else
`ifdef VC2
`else
`ifdef VC3
`else
`ifdef VC4
`else
`endif
`endif
`endif
`endif
`ifdef EN_VC0
`endif
`ifdef EN_VC1
`endif
`ifdef EN_VC2
`endif
`ifdef EN_VC3
`endif
`ifdef EN_VC4
`endif
`ifdef EN_VC5
`endif
`ifdef EN_VC6
`endif
`ifdef EN_VC7
`endif
assign rib82be = ldd88f4 | wwc47a6 | uif0030;
assign icc15f2 = co2bf0b | uxa40c4 | ph312b;
always @(posedge sys_clk or negedge rst_n) begin   if (rst_n == 1'b0) begin      lqe4a1a    <= 1'b0;      byd5d12       <= 1'b0;      sjae892   <= 1'b0;      pf74495       <= 1'b0;      pua24ae       <= 12'd0;      ir12572          <= 1'b0;      uk92b94      <= 3'b000;      sj95ca1      <= 1'b0;      yzae50c     <= 24'd0;   end   else begin      lqe4a1a    <= uif0030;      byd5d12       <= ldd88f4;      sjae892   <= wwc47a6;      pf74495       <= co2bf0b;      pua24ae       <= rt5f859;      ir12572          <= uxa40c4;      uk92b94      <= ip7f3bf;      sj95ca1      <= ph312b;      yzae50c     <= wl1895f;   end
end
assign do993fe    = !(db1677b || xl915be);
assign qtc9ff3    = !(gqb3bde || dob7de1);
assign sj3cfd4  = zxfc2cf && do993fe;
assign wje7ea5 = vie167e && qtc9ff3;
always @(posedge sys_clk or negedge rst_n) begin   if (rst_n == 1'b0) begin     ea72864    <= 1'b0;     hd94320   <= 1'b0;   end   else begin     ea72864       <= ldd88f4 | wwc47a6 | uif0030;     hd94320      <= co2bf0b | uxa40c4 | ph312b;   end
end
ng8cf0c  hd3ae9(      .sys_clk                  (sys_clk),   .rst_n                    (rst_n),   .pse18cc          (ldd748a),      .jrc662             (vxba456),      .zk63316           (vvd22b7),      .lf198b2               (xl915be),   .yxcc596                 (qv8adf7),   .os62cb4                 (cm56fbc),   .fp165a1               (dob7de1),   .xyb2d0e                 (yzbef0a),   .ba96872                 (off7854),
   .wlb4393            (gqbc2a4),   .uxa1c9c           (zke1520),   .vke4e4          (mga903),   .ay5cd66                 (cz75325),
`ifdef EN_VC0
      .hq93919                   (hq93919),      .ri9c8cb                  (ri9c8cb),      .tue465a                 (tue465a),
`endif
`ifdef EN_VC1
      .sj232d3                   (sj232d3),      .hd1969c                  (hd1969c),      .uicb4e7                 (uicb4e7),
`endif
`ifdef EN_VC2
      .pf5a739                   (pf5a739),      .end39ce                  (end39ce),      .tw9ce75                 (tw9ce75),
`endif
`ifdef EN_VC3
      .kde73aa                   (kde73aa),      .ux39d54                  (ux39d54),      .kqceaa5                 (kqceaa5),
`endif
`ifdef EN_VC4
      .ip75528                   (ip75528),      .ntaa944                  (ntaa944),      .al54a27                 (al54a27),
`endif
`ifdef EN_VC5
      .lfa513c                   (lfa513c),      .hd289e7                  (hd289e7),      .al44f3e                 (al44f3e),
`endif
`ifdef EN_VC6
      .hd279f5                   (hd279f5),      .an3cfaf                  (an3cfaf),      .ipe7d7d                 (ipe7d7d),
`endif
`ifdef EN_VC7
      .gq3ebed                   (gq3ebed),      .ykf5f68                  (ykf5f68),      .phafb41                 (phafb41),
`endif
      .os7da0f                    (rg42516),   .qted079              (mt128b3),   .ww683cd                (hd9459d),   .tx_vsd_data              (ria2cef),      .yx4e2a2                 (ngade42),   .al7fcee             (wj6f212),   .xw69c54                 (ps79094),   .jce1a71                 (vvc84a2),      .ls1e282               (vv7e6c2),   .zx74783               (ep80180),   .qia3c1e              (gqc04),   .tw1e0f1              (hqb3f3),   .icf078a              (me59f9b),   .ls83c50              (facfcd8),      .wlb4ebf               (vvf3617),   .xya75fd               (rv9b0bf),   .lqe4a1a            (vvd85fe),         .ba250d2            (ba250d2),      .an3c4c4                (an3c4c4),   .ene2624                (ene2624),   .mec4930            (mec4930),      .jpd27c8              (jpd27c8),   .do93e46             (do93e46),   .mt9f233            (mt9f233),      .xjc264f                 (xjc264f),   .jr1327f                (jr1327f),      .cm46737             (cm46737),      .sj23425                (sj23425),   .ec1a12c               (ec1a12c),   .tud0960                 (tud0960),   .hd84b02              (hd84b02),   .gqb98bf              (gqb98bf)   );
aaa91a  sjab4b9(      .sys_clk                  (sys_clk),   .rst_n                    (rst_n),      .sj23425                (do9918e),   .ec1a12c               (rtc8c73),   .tud0960                 (os4639f),   .hd84b02              (mg31cf9),         .wy24981                 (wy24981),   .zz13124             (zz13124),   .aa98926            (aa98926),   .kf2ead                     (ks24c08)   );
rg66dae  ipc940f (      .sys_clk                  (sys_clk),   .rst_n                    (rst_n),      .ls35987              (bl64b01),      .yzae707               (wyb31e1),   .fa7383c           (wy98f09),   .ng9c1e2                  (jpc7848),   .qge0f13                 (wl3c246),   .qv7898                 (xwe1234),      .an3c4c4                (zz91a3),   .ene2624                (xw48d1e),   .zz13124             (kq468f3),   .aa98926            (co34798),   .mec4930            (oua3cc0),   .wy24981                 (do1e601),   .ks24c08                (nrf300a),         .wwf5804               (wwf5804),   .vk30204                (vk30204),   .wyac021                 (wyac021),   .uv60109                (uv60109),   .ym84d                (ym84d),   .pu4269            (pu4269),   .qi2134a           (qi2134a),   .bn169d7               (bn169d7),      .wlb4ebf               (wlb4ebf),   .xya75fd               (xya75fd)   );
always@* begin ldd748a<={pse18cc>>1,ld7b613[0]};bl64b01<=ld7b613[1];vxba456<=ld7b613[2];vvd22b7<=ld7b613[3];xl915be<=ld7b613[4];qv8adf7<={yxcc596>>1,ld7b613[5]};cm56fbc<={os62cb4>>1,ld7b613[6]};dob7de1<=ld7b613[7];yzbef0a<={xyb2d0e>>1,ld7b613[8]};off7854<={ba96872>>1,ld7b613[9]};gqbc2a4<={wlb4393>>1,ld7b613[10]};zke1520<={uxa1c9c>>1,ld7b613[11]};mga903<={vke4e4>>1,ld7b613[12]};cz75325<={ay5cd66>>1,ld7b613[13]};uxa40c4<=ld7b613[14];ip7f3bf<={tx_pmtype>>1,ld7b613[15]};ph312b<=ld7b613[16];wl1895f<={tx_vsd_data>>1,ld7b613[17]};ldd88f4<=ld7b613[18];wwc47a6<=ld7b613[19];co2bf0b<=ld7b613[20];rt5f859<={jce1a71>>1,ld7b613[21]};zxfc2cf<=ld7b613[22];vie167e<=ld7b613[23];hqb3f3<={tw1e0f1>>1,ld7b613[24]};me59f9b<=ld7b613[25];facfcd8<={ls83c50>>1,ld7b613[26]};vv7e6c2<={ls1e282>>1,ld7b613[27]};wyb31e1<={yzae707>>1,ld7b613[28]};wy98f09<=ld7b613[29];jpc7848<=ld7b613[30];wl3c246<=ld7b613[31];xwe1234<=ld7b613[32];zz91a3<=ld7b613[33];xw48d1e<=ld7b613[34];oua3cc0<={mec4930>>1,ld7b613[35]};do1e601<=ld7b613[36];kq468f3<=ld7b613[37];co34798<=ld7b613[38];nrf300a<={ks24c08>>1,ld7b613[39]};vvd85fe<=ld7b613[40];ngade42<=ld7b613[41];wj6f212<=ld7b613[42];ps79094<=ld7b613[43];vvc84a2<={pua24ae>>1,ld7b613[44]};rg42516<=ld7b613[45];mt128b3<={uk92b94>>1,ld7b613[46]};hd9459d<=ld7b613[47];ria2cef<={yzae50c>>1,ld7b613[48]};db1677b<=ld7b613[49];gqb3bde<=ld7b613[50];do9918e<=ld7b613[51];rtc8c73<=ld7b613[52];os4639f<={tud0960>>1,ld7b613[53]};mg31cf9<={hd84b02>>1,ld7b613[54]};uif0030<=ld7b613[55];ep80180<=ld7b613[56];gqc04<=ld7b613[57];vvf3617<=ld7b613[58];rv9b0bf<=ld7b613[59];end
always@* begin necf6c2[2047]<=ls35987;necf6c2[2046]<=jrc662;necf6c2[2044]<=zk63316;necf6c2[2041]<=lf198b2;necf6c2[2035]<=yxcc596[0];necf6c2[2029]<=wje7ea5;necf6c2[2022]<=os62cb4[0];necf6c2[2011]<=wlb4ebf;necf6c2[1996]<=fp165a1;necf6c2[1974]<=xya75fd;necf6c2[1945]<=xyb2d0e[0];necf6c2[1943]<=ea72864;necf6c2[1922]<=icf078a;necf6c2[1842]<=ba96872[0];necf6c2[1839]<=hd94320;necf6c2[1797]<=ls83c50[0];necf6c2[1778]<=uk92b94[0];necf6c2[1776]<=zx74783;necf6c2[1637]<=wlb4393[0];necf6c2[1631]<=sj23425;necf6c2[1622]<=os7da0f;necf6c2[1546]<=ls1e282[0];necf6c2[1531]<=gqb98bf;necf6c2[1509]<=sj95ca1;necf6c2[1504]<=qia3c1e;necf6c2[1468]<=xw69c54;necf6c2[1391]<=yx4e2a2;necf6c2[1312]<=ene2624;necf6c2[1226]<=uxa1c9c[0];necf6c2[1215]<=ec1a12c;necf6c2[1197]<=tx_pmtype[0];necf6c2[1153]<=wy24981;necf6c2[1044]<=yzae707[0];necf6c2[1037]<=ks24c08[0];necf6c2[1023]<=pse18cc[0];necf6c2[1014]<=sj3cfd4;necf6c2[971]<=yzae50c[0];necf6c2[961]<=tw1e0f1[0];necf6c2[889]<=ir12572;necf6c2[888]<=jce1a71[0];necf6c2[811]<=ay5cd66[0];necf6c2[765]<=hd84b02[0];necf6c2[734]<=al7fcee;necf6c2[695]<=tx_vsd_data[0];necf6c2[656]<=an3c4c4;necf6c2[576]<=mec4930[0];necf6c2[518]<=aa98926;necf6c2[444]<=pua24ae[0];necf6c2[405]<=vke4e4[0];necf6c2[382]<=tud0960[0];necf6c2[347]<=ww683cd;necf6c2[328]<=qv7898;necf6c2[259]<=zz13124;necf6c2[222]<=pf74495;necf6c2[164]<=qge0f13;necf6c2[111]<=sjae892;necf6c2[82]<=ng9c1e2;necf6c2[55]<=byd5d12;necf6c2[41]<=fa7383c;necf6c2[27]<=lqe4a1a;end         assign suff972 = necf6c2,ld7b613 = cme5c87;   initial begin   jcc030e = $fopen(".fred");   $fdisplay( jcc030e, "%3h\n%3h", (thc27c7 >> 4) & fnc7fe5, (thc27c7 >> (mt9f1ff+4)) & fnc7fe5 );   $fclose(jcc030e);   $readmemh(".fred", qg721c0);   end   always @ (suff972) begin   ym8700c = qg721c0[1];       for (vk1872=0; vk1872<qgdb09f; vk1872=vk1872+1) begin           cme5c87[vk1872] = suff972[ym8700c];       rv38061  = ^(ym8700c & qg721c0[0]);       ym8700c =  {ym8700c, rv38061};       end   end
endmodule