module %m @ time %0d:\n", $time);
        $stop(1);
      end
    end
  endtask
endmodule