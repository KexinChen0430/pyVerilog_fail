module shifterZ0 (
  input_reg,
  shift_amount_1,
  un14_pos_output,
  ret_val,
  un11_output_6_d_0,
  out_shift_amount,
  un7_output_2_0_0,
  un7_output_2_1,
  output_d,
  shift_amount_1_i,
  un11_output_1,
  un11_output_2,
  un20_output_2,
  pre_output,
  done_inv_sqrt,
  un4_overflow_0,
  output_reg_pipe_12_RNIPJ901_O6,
  un9_0_axb_8,
  un9_0_s_6,
  un9_0_s_7,
  N_414,
  N_33,
  clk,
  N_420,
  un3_shift_right,
  N_410,
  un9_0_s_5,
  un9_0_s_8,
  N_79,
  N_50,
  un9_0_s_4,
  un9_0_s_3,
  N_13_0,
  N_100_i,
  N_31,
  N_18_0,
  N_378,
  N_33_0,
  N_80,
  N_51,
  un9_0_s_0,
  un9_0_s_1,
  m9_0_0,
  N_417,
  N_62,
  N_454,
  SUM1_0_i_1_1,
  N_56,
  N_434_i,
  N_431_i,
  N_428_i,
  N_425_i,
  un9_0_s_2,
  N_419,
  N_49,
  N_413,
  un20_output_0_0_a2_0_0_lut6_2_O5,
  un1_apply_nrlt8_1,
  un1_apply_nrlt7
)
;
input [11:10] input_reg ;
input [1:1] shift_amount_1 ;
input [6:3] un14_pos_output ;
input [3:1] ret_val ;
output [9:9] un11_output_6_d_0 ;
input [1:1] out_shift_amount ;
output [6:6] un7_output_2_0_0 ;
output [6:5] un7_output_2_1 ;
output [4:4] output_d ;
input [2:2] shift_amount_1_i ;
output un11_output_1 ;
output un11_output_2 ;
input [14:14] un20_output_2 ;
output [11:1] pre_output ;
input done_inv_sqrt ;
input un4_overflow_0 ;
output output_reg_pipe_12_RNIPJ901_O6 ;
input un9_0_axb_8 ;
input un9_0_s_6 ;
input un9_0_s_7 ;
output N_414 ;
output N_33 ;
input clk ;
output N_420 ;
input un3_shift_right ;
output N_410 ;
input un9_0_s_5 ;
input un9_0_s_8 ;
output N_79 ;
output N_50 ;
input un9_0_s_4 ;
input un9_0_s_3 ;
output N_13_0 ;
input N_100_i ;
output N_31 ;
output N_18_0 ;
input N_378 ;
output N_33_0 ;
output N_80 ;
output N_51 ;
input un9_0_s_0 ;
input un9_0_s_1 ;
output m9_0_0 ;
output N_417 ;
output N_62 ;
input N_454 ;
input SUM1_0_i_1_1 ;
output N_56 ;
output N_434_i ;
output N_431_i ;
output N_428_i ;
output N_425_i ;
input un9_0_s_2 ;
input N_419 ;
output N_49 ;
output N_413 ;
input un20_output_0_0_a2_0_0_lut6_2_O5 ;
input un1_apply_nrlt8_1 ;
input un1_apply_nrlt7 ;
wire un11_output_1 ;
wire un11_output_2 ;
wire done_inv_sqrt ;
wire un4_overflow_0 ;
wire output_reg_pipe_12_RNIPJ901_O6 ;
wire un9_0_axb_8 ;
wire un9_0_s_6 ;
wire un9_0_s_7 ;
wire N_414 ;
wire N_33 ;
wire clk ;
wire N_420 ;
wire un3_shift_right ;
wire N_410 ;
wire un9_0_s_5 ;
wire un9_0_s_8 ;
wire N_79 ;
wire N_50 ;
wire un9_0_s_4 ;
wire un9_0_s_3 ;
wire N_13_0 ;
wire N_100_i ;
wire N_31 ;
wire N_18_0 ;
wire N_378 ;
wire N_33_0 ;
wire N_80 ;
wire N_51 ;
wire un9_0_s_0 ;
wire un9_0_s_1 ;
wire m9_0_0 ;
wire N_417 ;
wire N_62 ;
wire N_454 ;
wire SUM1_0_i_1_1 ;
wire N_56 ;
wire N_434_i ;
wire N_431_i ;
wire N_428_i ;
wire N_425_i ;
wire un9_0_s_2 ;
wire N_419 ;
wire N_49 ;
wire N_413 ;
wire un20_output_0_0_a2_0_0_lut6_2_O5 ;
wire un1_apply_nrlt8_1 ;
wire un1_apply_nrlt7 ;
wire [6:3] un14_pos_outputf;
wire [6:3] pre_outputf;
wire [4:4] un11_output;
wire [6:4] un11_output_1_Z;
wire un4_overflow_if ;
wire VCC ;
wire un4_overflow_i_0 ;
wire output_reg_pipe_13 ;
wire m41 ;
wire output_reg_pipe ;
wire m44 ;
wire output_reg_pipe_5 ;
wire N_427 ;
wire output_reg_pipe_10 ;
wire N_430 ;
wire output_reg_pipe_15 ;
wire N_433 ;
wire m25_0_1 ;
wire m25_0_0 ;
wire m17_0_2 ;
wire GND ;
  FD output_reg_pipe_13_Z (
	.Q(output_reg_pipe_13),
	.D(m41),
	.C(clk)
);
  FD output_reg_pipe_12_Z (
	.Q(un4_overflow_if),
	.D(un4_overflow_i_0),
	.C(clk)
);
  FD output_reg_pipe_Z (
	.Q(output_reg_pipe),
	.D(m44),
	.C(clk)
);
// @27:84
  LUT5 output_reg_pipe_RNO (
	.I0(un4_overflow_0),
	.I1(pre_output[3]),
	.I2(N_420),
	.I3(output_reg_pipe),
	.I4(done_inv_sqrt),
	.O(m44)
);
defparam output_reg_pipe_RNO.INIT=32'h0101FF00;
// @27:84
  LUT6 output_reg_pipe_13_RNO (
	.I0(input_reg[10]),
	.I1(input_reg[11]),
	.I2(un4_overflow_0),
	.I3(N_420),
	.I4(output_reg_pipe_13),
	.I5(done_inv_sqrt),
	.O(m41)
);
defparam output_reg_pipe_13_RNO.INIT=64'hEF00EF00FFFF0000;
  FDE output_reg_pipe_1_Z (
	.Q(un14_pos_outputf[3]),
	.D(un14_pos_output[3]),
	.C(clk),
	.CE(done_inv_sqrt)
);
  FDE output_reg_pipe_4_Z (
	.Q(pre_outputf[3]),
	.D(pre_output[3]),
	.C(clk),
	.CE(done_inv_sqrt)
);
  FDE output_reg_pipe_5_Z (
	.Q(output_reg_pipe_5),
	.D(N_427),
	.C(clk),
	.CE(done_inv_sqrt)
);
  FDE output_reg_pipe_6_Z (
	.Q(un14_pos_outputf[4]),
	.D(un14_pos_output[4]),
	.C(clk),
	.CE(done_inv_sqrt)
);
  FDE output_reg_pipe_9_Z (
	.Q(pre_outputf[4]),
	.D(pre_output[4]),
	.C(clk),
	.CE(done_inv_sqrt)
);
  FDE output_reg_pipe_10_Z (
	.Q(output_reg_pipe_10),
	.D(N_430),
	.C(clk),
	.CE(done_inv_sqrt)
);
  FDE output_reg_pipe_11_Z (
	.Q(un14_pos_outputf[5]),
	.D(un14_pos_output[5]),
	.C(clk),
	.CE(done_inv_sqrt)
);
  FDE output_reg_pipe_14_Z (
	.Q(pre_outputf[5]),
	.D(pre_output[5]),
	.C(clk),
	.CE(done_inv_sqrt)
);
  FDE output_reg_pipe_15_Z (
	.Q(output_reg_pipe_15),
	.D(N_433),
	.C(clk),
	.CE(done_inv_sqrt)
);
  FDE output_reg_pipe_16_Z (
	.Q(un14_pos_outputf[6]),
	.D(un14_pos_output[6]),
	.C(clk),
	.CE(done_inv_sqrt)
);
  FDE output_reg_pipe_19_Z (
	.Q(pre_outputf[6]),
	.D(pre_output[6]),
	.C(clk),
	.CE(done_inv_sqrt)
);
  LUT3 \un11_output_RNIM9LT[5]  (
	.I0(un3_shift_right),
	.I1(un7_output_2_1[5]),
	.I2(un11_output_1),
	.O(pre_output[5])
);
defparam \un11_output_RNIM9LT[5] .INIT=8'hD8;
// @27:84
  LUT4 m26 (
	.I0(ret_val[3]),
	.I1(N_410),
	.I2(m25_0_1),
	.I3(m25_0_0),
	.O(pre_output[8])
);
defparam m26.INIT=16'hFFD8;
// @8:60
  LUT5 \un11_output_6_d_0_cZ[9]  (
	.I0(ret_val[3]),
	.I1(ret_val[1]),
	.I2(shift_amount_1[1]),
	.I3(un9_0_s_5),
	.I4(un9_0_s_8),
	.O(un11_output_6_d_0[9])
);
defparam \un11_output_6_d_0_cZ[9] .INIT=32'hF8F00800;
  LUT5 \un11_output_3_RNITKM12[2]  (
	.I0(ret_val[3]),
	.I1(ret_val[1]),
	.I2(un3_shift_right),
	.I3(N_79),
	.I4(N_50),
	.O(pre_output[2])
);
defparam \un11_output_3_RNITKM12[2] .INIT=32'hFFF00700;
// @27:84
  LUT4 m19 (
	.I0(ret_val[2]),
	.I1(un9_0_axb_8),
	.I2(shift_amount_1[1]),
	.I3(un9_0_s_4),
	.O(N_410)
);
defparam m19.INIT=16'h0600;
// @27:84
  LUT4 m12 (
	.I0(ret_val[2]),
	.I1(un9_0_axb_8),
	.I2(shift_amount_1[1]),
	.I3(un9_0_s_3),
	.O(N_13_0)
);
defparam m12.INIT=16'h0600;
  LUT3 m31 (
	.I0(N_100_i),
	.I1(un9_0_s_6),
	.I2(N_31),
	.O(pre_output[10])
);
defparam m31.INIT=8'hE4;
  LUT3 m18 (
	.I0(N_100_i),
	.I1(un9_0_s_3),
	.I2(N_18_0),
	.O(pre_output[7])
);
defparam m18.INIT=8'hE4;
  LUT5 \un11_output_RNIL9QU3[4]  (
	.I0(N_378),
	.I1(un3_shift_right),
	.I2(un9_0_s_6),
	.I3(N_33_0),
	.I4(un11_output[4]),
	.O(pre_output[4])
);
defparam \un11_output_RNIL9QU3[4] .INIT=32'hF733CC80;
// @8:59
  LUT5 \un7_output_2_0[6]  (
	.I0(ret_val[3]),
	.I1(ret_val[1]),
	.I2(un9_0_axb_8),
	.I3(out_shift_amount[1]),
	.I4(un9_0_s_8),
	.O(un7_output_2_0_0[6])
);
defparam \un7_output_2_0[6] .INIT=32'h437F007F;
  LUT6 \un11_output_3_RNI53BN3[3]  (
	.I0(ret_val[3]),
	.I1(ret_val[1]),
	.I2(un9_0_axb_8),
	.I3(un3_shift_right),
	.I4(N_80),
	.I5(N_51),
	.O(pre_output[3])
);
defparam \un11_output_3_RNI53BN3[3] .INIT=64'hFF7FFF00007F0000;
// @27:84
  LUT6 m25_0_1_cZ (
	.I0(ret_val[1]),
	.I1(un9_0_axb_8),
	.I2(out_shift_amount[1]),
	.I3(un3_shift_right),
	.I4(un9_0_s_8),
	.I5(un9_0_s_7),
	.O(m25_0_1)
);
defparam m25_0_1_cZ.INIT=64'h090F000609090000;
// @27:84
  LUT6 m30 (
	.I0(ret_val[1]),
	.I1(un9_0_axb_8),
	.I2(out_shift_amount[1]),
	.I3(un3_shift_right),
	.I4(un9_0_s_8),
	.I5(un9_0_s_7),
	.O(N_31)
);
defparam m30.INIT=64'h00F0006000900000;
// @8:59
  LUT5 \un7_output_2_1_cZ[5]  (
	.I0(ret_val[1]),
	.I1(un9_0_axb_8),
	.I2(out_shift_amount[1]),
	.I3(un9_0_s_6),
	.I4(un9_0_s_7),
	.O(un7_output_2_1[5])
);
defparam \un7_output_2_1_cZ[5] .INIT=32'hFF990F09;
// @8:59
  LUT5 \un7_output_2_1_cZ[6]  (
	.I0(ret_val[1]),
	.I1(un9_0_axb_8),
	.I2(out_shift_amount[1]),
	.I3(un9_0_s_6),
	.I4(un9_0_s_7),
	.O(un7_output_2_1[6])
);
defparam \un7_output_2_1_cZ[6] .INIT=32'hFFF69990;
// @27:84
  LUT6 m25_0_0_cZ (
	.I0(ret_val[1]),
	.I1(un9_0_axb_8),
	.I2(out_shift_amount[1]),
	.I3(un3_shift_right),
	.I4(un9_0_s_5),
	.I5(un9_0_s_6),
	.O(m25_0_0)
);
defparam m25_0_0_cZ.INIT=64'h00F0009000600000;
// @8:59
  LUT5 \output_d_cZ[4]  (
	.I0(ret_val[1]),
	.I1(un9_0_axb_8),
	.I2(un3_shift_right),
	.I3(un9_0_s_6),
	.I4(un11_output[4]),
	.O(output_d[4])
);
defparam \output_d_cZ[4] .INIT=32'h9F0F9000;
// @27:84
  LUT6 m9_0_0_c (
	.I0(ret_val[1]),
	.I1(un9_0_axb_8),
	.I2(out_shift_amount[1]),
	.I3(un3_shift_right),
	.I4(un9_0_s_0),
	.I5(un9_0_s_1),
	.O(m9_0_0)
);
defparam m9_0_0_c.INIT=64'h0F09060009090000;
// @27:84
  LUT4 m33 (
	.I0(ret_val[2]),
	.I1(shift_amount_1[1]),
	.I2(un3_shift_right),
	.I3(un9_0_s_8),
	.O(N_417)
);
defparam m33.INIT=16'h0400;
// @8:60
  LUT4 \un11_output_1[7]  (
	.I0(ret_val[1]),
	.I1(un9_0_axb_8),
	.I2(un9_0_s_6),
	.I3(un9_0_s_7),
	.O(N_62)
);
defparam \un11_output_1[7] .INIT=16'hF960;
// @8:60
  LUT6 \un11_output_1[1]  (
	.I0(N_454),
	.I1(SUM1_0_i_1_1),
	.I2(ret_val[1]),
	.I3(un9_0_axb_8),
	.I4(un9_0_s_0),
	.I5(un9_0_s_1),
	.O(N_56)
);
defparam \un11_output_1[1] .INIT=64'hFFFF3013CFEC0000;
// @8:59
  LUT4 \un7_output_0[4]  (
	.I0(ret_val[1]),
	.I1(un9_0_axb_8),
	.I2(un9_0_s_4),
	.I3(un9_0_s_5),
	.O(N_33_0)
);
defparam \un7_output_0[4] .INIT=16'hF690;
// @13:37
  LUT5 output_reg_pipe_15_RNIJLNH1 (
	.I0(un14_pos_outputf[6]),
	.I1(output_reg_pipe_15),
	.I2(pre_outputf[6]),
	.I3(un4_overflow_if),
	.I4(output_reg_pipe_13),
	.O(N_434_i)
);
defparam output_reg_pipe_15_RNIJLNH1.INIT=32'h22277277;
// @13:37
  LUT5 output_reg_pipe_10_RNI4LNH1 (
	.I0(un14_pos_outputf[5]),
	.I1(output_reg_pipe_10),
	.I2(pre_outputf[5]),
	.I3(un4_overflow_if),
	.I4(output_reg_pipe_13),
	.O(N_431_i)
);
defparam output_reg_pipe_10_RNI4LNH1.INIT=32'h22277277;
// @13:37
  LUT5 output_reg_pipe_5_RNI0B2S (
	.I0(un14_pos_outputf[4]),
	.I1(output_reg_pipe_5),
	.I2(pre_outputf[4]),
	.I3(un4_overflow_if),
	.I4(output_reg_pipe_13),
	.O(N_428_i)
);
defparam output_reg_pipe_5_RNI0B2S.INIT=32'h22277277;
// @13:37
  LUT5 output_reg_pipe_1_RNI23E61 (
	.I0(un14_pos_outputf[3]),
	.I1(output_reg_pipe),
	.I2(pre_outputf[3]),
	.I3(un4_overflow_if),
	.I4(output_reg_pipe_13),
	.O(N_425_i)
);
defparam output_reg_pipe_1_RNI23E61.INIT=32'h22277277;
// @8:60
  LUT5 \un11_output_3[2]  (
	.I0(shift_amount_1_i[2]),
	.I1(shift_amount_1[1]),
	.I2(un9_0_s_0),
	.I3(un9_0_s_1),
	.I4(un9_0_s_2),
	.O(N_79)
);
defparam \un11_output_3[2] .INIT=32'hBA329810;
// @8:60
  LUT5 \un11_output_3[3]  (
	.I0(shift_amount_1_i[2]),
	.I1(shift_amount_1[1]),
	.I2(un9_0_s_2),
	.I3(N_56),
	.I4(un9_0_s_3),
	.O(N_80)
);
defparam \un11_output_3[3] .INIT=32'hF7A2D580;
// @8:60
  LUT6_L \un11_output_1[5]  (
	.I0(shift_amount_1_i[2]),
	.I1(N_100_i),
	.I2(shift_amount_1[1]),
	.I3(un9_0_s_1),
	.I4(un9_0_s_2),
	.I5(un9_0_s_3),
	.LO(un11_output_1_Z[5])
);
defparam \un11_output_1[5] .INIT=64'h4644060442400200;
// @8:60
  LUT6_L \un11_output_1[4]  (
	.I0(shift_amount_1_i[2]),
	.I1(N_100_i),
	.I2(shift_amount_1[1]),
	.I3(un9_0_s_0),
	.I4(un9_0_s_1),
	.I5(un9_0_s_2),
	.LO(un11_output_1_Z[4])
);
defparam \un11_output_1[4] .INIT=64'h4644060442400200;
// @8:59
  LUT6 \un7_output[1]  (
	.I0(N_419),
	.I1(N_378),
	.I2(N_100_i),
	.I3(un9_0_s_1),
	.I4(un9_0_s_2),
	.I5(un9_0_s_3),
	.O(N_49)
);
defparam \un7_output[1] .INIT=64'hEA62C840AA228800;
// @8:59
  LUT6 \un7_output[2]  (
	.I0(N_419),
	.I1(N_378),
	.I2(N_100_i),
	.I3(un9_0_s_2),
	.I4(un9_0_s_3),
	.I5(un9_0_s_4),
	.O(N_50)
);
defparam \un7_output[2] .INIT=64'hEA62C840AA228800;
// @8:60
  LUT6_L \un11_output_1[6]  (
	.I0(N_378),
	.I1(N_100_i),
	.I2(out_shift_amount[1]),
	.I3(un9_0_s_2),
	.I4(un9_0_s_3),
	.I5(un9_0_s_4),
	.LO(un11_output_1_Z[6])
);
defparam \un11_output_1[6] .INIT=64'hC2C0828042400200;
// @27:84
  LUT6_L m17_0_2_cZ (
	.I0(N_378),
	.I1(out_shift_amount[1]),
	.I2(un3_shift_right),
	.I3(un9_0_s_4),
	.I4(un9_0_s_5),
	.I5(un9_0_s_8),
	.LO(m17_0_2)
);
defparam m17_0_2_cZ.INIT=64'h1C1814100C080400;
// @27:84
  LUT6 m25_0 (
	.I0(N_378),
	.I1(out_shift_amount[1]),
	.I2(un3_shift_right),
	.I3(un9_0_s_8),
	.I4(un9_0_s_7),
	.I5(m25_0_0),
	.O(N_413)
);
defparam m25_0.INIT=64'hFFFFFFFF23012200;
// @8:60
  LUT6 \un11_output[5]  (
	.I0(shift_amount_1_i[2]),
	.I1(N_378),
	.I2(N_100_i),
	.I3(un9_0_s_4),
	.I4(un9_0_s_5),
	.I5(un11_output_1_Z[5]),
	.O(un11_output_1)
);
defparam \un11_output[5] .INIT=64'hFFFFFFFFA0802000;
// @8:60
  LUT6 \un11_output_cZ[4]  (
	.I0(shift_amount_1_i[2]),
	.I1(N_378),
	.I2(N_100_i),
	.I3(un9_0_s_3),
	.I4(un9_0_s_4),
	.I5(un11_output_1_Z[4]),
	.O(un11_output[4])
);
defparam \un11_output_cZ[4] .INIT=64'hFFFFFFFFA0802000;
// @8:59
  LUT6 \output_0[9]  (
	.I0(un20_output_0_0_a2_0_0_lut6_2_O5),
	.I1(N_378),
	.I2(un3_shift_right),
	.I3(un9_0_s_6),
	.I4(un9_0_s_7),
	.I5(un11_output_6_d_0[9]),
	.O(pre_output[9])
);
defparam \output_0[9] .INIT=64'h0F0D07050A080200;
// @27:84
  LUT6 m34 (
	.I0(N_100_i),
	.I1(out_shift_amount[1]),
	.I2(shift_amount_1[1]),
	.I3(un3_shift_right),
	.I4(un9_0_s_8),
	.I5(un9_0_s_7),
	.O(pre_output[11])
);
defparam m34.INIT=64'h0081000100800000;
// @8:59
  LUT6 \un7_output_2[3]  (
	.I0(N_378),
	.I1(N_100_i),
	.I2(out_shift_amount[1]),
	.I3(un9_0_s_3),
	.I4(un9_0_s_4),
	.I5(un9_0_s_5),
	.O(N_51)
);
defparam \un7_output_2[3] .INIT=64'h8C8488800C040800;
// @27:84
  LUT6 m17_0 (
	.I0(N_378),
	.I1(out_shift_amount[1]),
	.I2(un3_shift_right),
	.I3(un9_0_s_6),
	.I4(un9_0_s_7),
	.I5(m17_0_2),
	.O(N_18_0)
);
defparam m17_0.INIT=64'hFFFFFFFF23220100;
// @8:60
  LUT6 \un11_output[6]  (
	.I0(N_378),
	.I1(N_100_i),
	.I2(out_shift_amount[1]),
	.I3(un9_0_s_5),
	.I4(un9_0_s_6),
	.I5(un11_output_1_Z[6]),
	.O(un11_output_2)
);
defparam \un11_output[6] .INIT=64'hFFFFFFFF0C080400;
// @27:84
  LUT6 \output_0_RNIMQFRP[9]  (
	.I0(pre_output[11]),
	.I1(pre_output[10]),
	.I2(pre_output[9]),
	.I3(pre_output[8]),
	.I4(un1_apply_nrlt8_1),
	.I5(un1_apply_nrlt7),
	.O(N_420)
);
defparam \output_0_RNIMQFRP[9] .INIT=64'h0101011101110111;
// @27:84
  LUT5_L output_reg_pipe_5_RNO (
	.I0(input_reg[10]),
	.I1(input_reg[11]),
	.I2(un4_overflow_0),
	.I3(pre_output[4]),
	.I4(N_420),
	.LO(N_427)
);
defparam output_reg_pipe_5_RNO.INIT=32'h000000EF;
// @27:84
  LUT5_L output_reg_pipe_10_RNO (
	.I0(input_reg[10]),
	.I1(input_reg[11]),
	.I2(un4_overflow_0),
	.I3(pre_output[5]),
	.I4(N_420),
	.LO(N_430)
);
defparam output_reg_pipe_10_RNO.INIT=32'h000000EF;
// @27:84
  LUT5_L output_reg_pipe_15_RNO (
	.I0(input_reg[10]),
	.I1(input_reg[11]),
	.I2(un4_overflow_0),
	.I3(pre_output[6]),
	.I4(N_420),
	.LO(N_433)
);
defparam output_reg_pipe_15_RNO.INIT=32'h000000EF;
  LUT4 \un7_output_RNIN1BC1[1]  (
	.I0(un20_output_2[14]),
	.I1(un3_shift_right),
	.I2(N_56),
	.I3(N_49),
	.O(pre_output[1])
);
defparam \un7_output_RNIN1BC1[1] .INIT=16'hEC20;
  LUT4 \un7_output_2_0_RNI7K981[6]  (
	.I0(un3_shift_right),
	.I1(un7_output_2_0_0[6]),
	.I2(un7_output_2_1[6]),
	.I3(un11_output_2),
	.O(pre_output[6])
);
defparam \un7_output_2_0_RNI7K981[6] .INIT=16'hD580;
  VCC VCC_cZ (
	.P(VCC)
);
  GND GND_cZ (
	.G(GND)
);
// @27:84
  LUT4 m27_lut6_2_o6 (
	.I0(ret_val[2]),
	.I1(un9_0_axb_8),
	.I2(shift_amount_1[1]),
	.I3(un9_0_s_6),
	.O(N_414)
);
defparam m27_lut6_2_o6.INIT=16'h0600;
// @27:84
  LUT4 m27_lut6_2_o5 (
	.I0(ret_val[2]),
	.I1(un9_0_axb_8),
	.I2(shift_amount_1[1]),
	.I3(un9_0_s_7),
	.O(N_33)
);
defparam m27_lut6_2_o5.INIT=16'h0600;
  LUT4 output_reg_pipe_12_RNIPJ901_o6 (
	.I0(input_reg[10]),
	.I1(input_reg[11]),
	.I2(done_inv_sqrt),
	.I3(un4_overflow_0),
	.O(output_reg_pipe_12_RNIPJ901_O6)
);
defparam output_reg_pipe_12_RNIPJ901_o6.INIT=16'h1000;
  LUT5 output_reg_pipe_12_RNIPJ901_o5 (
	.I0(un4_overflow_if),
	.I1(input_reg[10]),
	.I2(input_reg[11]),
	.I3(done_inv_sqrt),
	.I4(un4_overflow_0),
	.O(un4_overflow_i_0)
);
defparam output_reg_pipe_12_RNIPJ901_o5.INIT=32'hFCAAFFAA;
endmodule