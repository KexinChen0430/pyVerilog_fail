module QL_DSP1 (
    input  [19:0] a,
    input  [17:0] b,
    input  clk0,
    (* clkbuf_sink *)
    input  clk1,
    (* clkbuf_sink *)
    input  [ 1:0] feedback0,
    input  [ 1:0] feedback1,
    input  load_acc0,
    input  load_acc1,
    input  reset0,
    input  reset1,
    output reg [37:0] z
);
    parameter MODE_BITS = 27'b00000000000000000000000000;
endmodule