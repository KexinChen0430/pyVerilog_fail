module top ;
          wire  Net_3491;
          wire  Net_3490;
          wire  Net_3489;
          wire  Net_3488;
          wire  Net_3487;
          wire  Net_3486;
          wire  Net_3485;
          wire  Net_3484;
          wire  Net_3483;
          wire  Net_3482;
          wire  Net_3481;
          wire  Net_3480;
          wire  Net_3479;
          wire  Net_3478;
          wire  Net_3477;
          wire  Net_3476;
          wire  Net_3475;
          wire  Net_3474;
          wire  Net_3473;
          wire  Net_3450;
	wire [0:0] tmpOE__LED_G_net;
	wire [0:0] tmpFB_0__LED_G_net;
	wire [0:0] tmpIO_0__LED_G_net;
	wire [0:0] tmpINTERRUPT_0__LED_G_net;
	electrical [0:0] tmpSIOVREF__LED_G_net;
	cy_psoc3_pins_v1_10
		#(.id("e851a3b9-efb8-48be-bbb8-b303b216c393"),
		  .drive_mode(3'b110),
		  .ibuf_enabled(1'b1),
		  .init_dr_st(1'b1),
		  .input_clk_en(0),
		  .input_sync(1'b1),
		  .input_sync_mode(1'b0),
		  .intr_mode(2'b00),
		  .invert_in_clock(0),
		  .invert_in_clock_en(0),
		  .invert_in_reset(0),
		  .invert_out_clock(0),
		  .invert_out_clock_en(0),
		  .invert_out_reset(0),
		  .io_voltage(""),
		  .layout_mode("CONTIGUOUS"),
		  .oe_conn(1'b0),
		  .oe_reset(0),
		  .oe_sync(1'b0),
		  .output_clk_en(0),
		  .output_clock_mode(1'b0),
		  .output_conn(1'b0),
		  .output_mode(1'b0),
		  .output_reset(0),
		  .output_sync(1'b0),
		  .pa_in_clock(-1),
		  .pa_in_clock_en(-1),
		  .pa_in_reset(-1),
		  .pa_out_clock(-1),
		  .pa_out_clock_en(-1),
		  .pa_out_reset(-1),
		  .pin_aliases(""),
		  .pin_mode("O"),
		  .por_state(4),
		  .sio_group_cnt(0),
		  .sio_hyst(1'b1),
		  .sio_ibuf(""),
		  .sio_info(2'b00),
		  .sio_obuf(""),
		  .sio_refsel(""),
		  .sio_vtrip(""),
		  .sio_hifreq(""),
		  .sio_vohsel(""),
		  .slew_rate(1'b0),
		  .spanning(0),
		  .use_annotation(1'b0),
		  .vtrip(2'b10),
		  .width(1),
		  .ovt_hyst_trim(1'b0),
		  .ovt_needed(1'b0),
		  .ovt_slew_control(2'b00),
		  .input_buffer_sel(2'b00))
		LED_G
		 (.oe(tmpOE__LED_G_net),
		  .y({1'b0}),
		  .fb({tmpFB_0__LED_G_net[0:0]}),
		  .io({tmpIO_0__LED_G_net[0:0]}),
		  .siovref(tmpSIOVREF__LED_G_net),
		  .interrupt({tmpINTERRUPT_0__LED_G_net[0:0]}),
		  .in_clock({1'b0}),
		  .in_clock_en({1'b1}),
		  .in_reset({1'b0}),
		  .out_clock({1'b0}),
		  .out_clock_en({1'b1}),
		  .out_reset({1'b0}));
	assign tmpOE__LED_G_net = (`CYDEV_CHIP_MEMBER_USED == `CYDEV_CHIP_MEMBER_3A && `CYDEV_CHIP_REVISION_USED < `CYDEV_CHIP_REVISION_3A_ES3) ? ~{1'b1} : {1'b1};
	wire [0:0] tmpOE__LED_R_net;
	wire [0:0] tmpFB_0__LED_R_net;
	wire [0:0] tmpIO_0__LED_R_net;
	wire [0:0] tmpINTERRUPT_0__LED_R_net;
	electrical [0:0] tmpSIOVREF__LED_R_net;
	cy_psoc3_pins_v1_10
		#(.id("46bcb939-fabe-42b9-90af-3e1c6577dc70"),
		  .drive_mode(3'b110),
		  .ibuf_enabled(1'b1),
		  .init_dr_st(1'b1),
		  .input_clk_en(0),
		  .input_sync(1'b1),
		  .input_sync_mode(1'b0),
		  .intr_mode(2'b00),
		  .invert_in_clock(0),
		  .invert_in_clock_en(0),
		  .invert_in_reset(0),
		  .invert_out_clock(0),
		  .invert_out_clock_en(0),
		  .invert_out_reset(0),
		  .io_voltage(""),
		  .layout_mode("CONTIGUOUS"),
		  .oe_conn(1'b0),
		  .oe_reset(0),
		  .oe_sync(1'b0),
		  .output_clk_en(0),
		  .output_clock_mode(1'b0),
		  .output_conn(1'b0),
		  .output_mode(1'b0),
		  .output_reset(0),
		  .output_sync(1'b0),
		  .pa_in_clock(-1),
		  .pa_in_clock_en(-1),
		  .pa_in_reset(-1),
		  .pa_out_clock(-1),
		  .pa_out_clock_en(-1),
		  .pa_out_reset(-1),
		  .pin_aliases(""),
		  .pin_mode("O"),
		  .por_state(4),
		  .sio_group_cnt(0),
		  .sio_hyst(1'b1),
		  .sio_ibuf(""),
		  .sio_info(2'b00),
		  .sio_obuf(""),
		  .sio_refsel(""),
		  .sio_vtrip(""),
		  .sio_hifreq(""),
		  .sio_vohsel(""),
		  .slew_rate(1'b0),
		  .spanning(0),
		  .use_annotation(1'b0),
		  .vtrip(2'b10),
		  .width(1),
		  .ovt_hyst_trim(1'b0),
		  .ovt_needed(1'b0),
		  .ovt_slew_control(2'b00),
		  .input_buffer_sel(2'b00))
		LED_R
		 (.oe(tmpOE__LED_R_net),
		  .y({1'b0}),
		  .fb({tmpFB_0__LED_R_net[0:0]}),
		  .io({tmpIO_0__LED_R_net[0:0]}),
		  .siovref(tmpSIOVREF__LED_R_net),
		  .interrupt({tmpINTERRUPT_0__LED_R_net[0:0]}),
		  .in_clock({1'b0}),
		  .in_clock_en({1'b1}),
		  .in_reset({1'b0}),
		  .out_clock({1'b0}),
		  .out_clock_en({1'b1}),
		  .out_reset({1'b0}));
	assign tmpOE__LED_R_net = (`CYDEV_CHIP_MEMBER_USED == `CYDEV_CHIP_MEMBER_3A && `CYDEV_CHIP_REVISION_USED < `CYDEV_CHIP_REVISION_3A_ES3) ? ~{1'b1} : {1'b1};
	cy_isr_v1_0
		#(.int_type(2'b10))
		WDT_isr
		 (.int_signal(Net_3450));
	cy_gsref_v1_0
		#(.guid("1563FAA8-0748-4a1c-9785-CED309984BE3"))
		WDT
		 (.sig_out(Net_3450));
    SCB_P4_v3_20_0 UART (
        .cts_in(1'b0),
        .tx_out(Net_3474),
        .rts_out(Net_3475),
        .interrupt(Net_3476),
        .clock(1'b0),
        .rx_tr_out(Net_3478),
        .tx_tr_out(Net_3479),
        .s_mosi(1'b0),
        .s_sclk(1'b0),
        .s_ss(1'b0),
        .m_miso(1'b0),
        .m_mosi(Net_3484),
        .m_sclk(Net_3485),
        .m_ss0(Net_3486),
        .m_ss1(Net_3487),
        .m_ss2(Net_3488),
        .m_ss3(Net_3489),
        .s_miso(Net_3490),
        .rx_in(1'b0));
	wire [0:0] tmpOE__LED_B_net;
	wire [0:0] tmpFB_0__LED_B_net;
	wire [0:0] tmpIO_0__LED_B_net;
	wire [0:0] tmpINTERRUPT_0__LED_B_net;
	electrical [0:0] tmpSIOVREF__LED_B_net;
	cy_psoc3_pins_v1_10
		#(.id("3b8d3c3c-27ec-4327-b3ef-9251ee2d52b4"),
		  .drive_mode(3'b110),
		  .ibuf_enabled(1'b1),
		  .init_dr_st(1'b1),
		  .input_clk_en(0),
		  .input_sync(1'b1),
		  .input_sync_mode(1'b0),
		  .intr_mode(2'b00),
		  .invert_in_clock(0),
		  .invert_in_clock_en(0),
		  .invert_in_reset(0),
		  .invert_out_clock(0),
		  .invert_out_clock_en(0),
		  .invert_out_reset(0),
		  .io_voltage(""),
		  .layout_mode("CONTIGUOUS"),
		  .oe_conn(1'b0),
		  .oe_reset(0),
		  .oe_sync(1'b0),
		  .output_clk_en(0),
		  .output_clock_mode(1'b0),
		  .output_conn(1'b0),
		  .output_mode(1'b0),
		  .output_reset(0),
		  .output_sync(1'b0),
		  .pa_in_clock(-1),
		  .pa_in_clock_en(-1),
		  .pa_in_reset(-1),
		  .pa_out_clock(-1),
		  .pa_out_clock_en(-1),
		  .pa_out_reset(-1),
		  .pin_aliases(""),
		  .pin_mode("O"),
		  .por_state(4),
		  .sio_group_cnt(0),
		  .sio_hyst(1'b1),
		  .sio_ibuf(""),
		  .sio_info(2'b00),
		  .sio_obuf(""),
		  .sio_refsel(""),
		  .sio_vtrip(""),
		  .sio_hifreq(""),
		  .sio_vohsel(""),
		  .slew_rate(1'b0),
		  .spanning(0),
		  .use_annotation(1'b0),
		  .vtrip(2'b10),
		  .width(1),
		  .ovt_hyst_trim(1'b0),
		  .ovt_needed(1'b0),
		  .ovt_slew_control(2'b00),
		  .input_buffer_sel(2'b00))
		LED_B
		 (.oe(tmpOE__LED_B_net),
		  .y({1'b0}),
		  .fb({tmpFB_0__LED_B_net[0:0]}),
		  .io({tmpIO_0__LED_B_net[0:0]}),
		  .siovref(tmpSIOVREF__LED_B_net),
		  .interrupt({tmpINTERRUPT_0__LED_B_net[0:0]}),
		  .in_clock({1'b0}),
		  .in_clock_en({1'b1}),
		  .in_reset({1'b0}),
		  .out_clock({1'b0}),
		  .out_clock_en({1'b1}),
		  .out_reset({1'b0}));
	assign tmpOE__LED_B_net = (`CYDEV_CHIP_MEMBER_USED == `CYDEV_CHIP_MEMBER_3A && `CYDEV_CHIP_REVISION_USED < `CYDEV_CHIP_REVISION_3A_ES3) ? ~{1'b1} : {1'b1};
	cy_isr_v1_0
		#(.int_type(2'b10))
		UART_isr
		 (.int_signal(Net_3476));
endmodule