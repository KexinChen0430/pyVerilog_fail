module SCB_P4_v3_0_0 (
    interrupt,
    clock,
    rx_tr_out,
    tx_tr_out);
    output      interrupt;
    input       clock;
    output      rx_tr_out;
    output      tx_tr_out;
          wire  uncfg_rx_irq;
          wire  Net_1191;
          wire  Net_1258;
          wire  Net_1099;
          wire  rx_irq;
          wire [3:0] ss;
          wire  Net_1257;
          wire  Net_1197;
          wire  Net_1196;
          wire  Net_1195;
          wire  Net_1194;
          wire  Net_1193;
          wire  Net_1263;
          wire  Net_663;
          wire  Net_547;
          wire  Net_467;
          wire  Net_1090;
          wire  Net_1091;
          wire  Net_1172;
          wire  Net_1089;
          wire  Net_1088;
          wire  Net_387;
          wire  Net_252;
          wire  Net_1087;
          wire  Net_1086;
          wire  Net_1000;
          wire  Net_915;
          wire  Net_916;
          wire  Net_1175;
          wire  Net_654;
          wire  Net_990;
          wire  Net_652;
          wire  Net_459;
          wire  Net_580;
          wire  Net_581;
          wire  Net_452;
          wire  Net_909;
          wire  Net_1001;
          wire  Net_899;
          wire  Net_747;
          wire  Net_891;
          wire  Net_1028;
          wire  Net_1170;
          wire  Net_1061;
          wire  Net_1053;
          wire  Net_1055;
          wire  Net_1062;
          wire  Net_1059;
          wire  Net_847;
	cy_clock_v1_0
		#(.id("43ec2fa1-bf22-4b71-9477-b6ca7b97f0b0/2dc2d7a8-ce2b-43c7-af4a-821c8cd73ccf"),
		  .source_clock_id(""),
		  .divisor(0),
		  .period("667735042.735043"),
		  .is_direct(0),
		  .is_digital(0))
		SCBCLK
		 (.clock_out(Net_847));
    ZeroTerminal ZeroTerminal_5 (
        .z(Net_459));
	// select_s_VM (cy_virtualmux_v1_0)
	assign Net_652 = Net_459;
    ZeroTerminal ZeroTerminal_4 (
        .z(Net_452));
    ZeroTerminal ZeroTerminal_3 (
        .z(Net_1194));
    ZeroTerminal ZeroTerminal_2 (
        .z(Net_1195));
    ZeroTerminal ZeroTerminal_1 (
        .z(Net_1196));
	// rx_VM (cy_virtualmux_v1_0)
	assign Net_654 = Net_1197;
	// rx_wake_VM (cy_virtualmux_v1_0)
	assign Net_1257 = uncfg_rx_irq;
	// clock_VM (cy_virtualmux_v1_0)
	assign Net_1170 = Net_847;
	// sclk_s_VM (cy_virtualmux_v1_0)
	assign Net_990 = Net_1196;
	// mosi_s_VM (cy_virtualmux_v1_0)
	assign Net_909 = Net_1194;
	// miso_m_VM (cy_virtualmux_v1_0)
	assign Net_663 = Net_1195;
	wire [0:0] tmpOE__tx_net;
	wire [0:0] tmpFB_0__tx_net;
	wire [0:0] tmpIO_0__tx_net;
	wire [0:0] tmpINTERRUPT_0__tx_net;
	electrical [0:0] tmpSIOVREF__tx_net;
	cy_psoc3_pins_v1_10
		#(.id("43ec2fa1-bf22-4b71-9477-b6ca7b97f0b0/23b8206d-1c77-4e61-be4a-b4037d5de5fc"),
		  .drive_mode(3'b110),
		  .ibuf_enabled(1'b0),
		  .init_dr_st(1'b1),
		  .input_clk_en(0),
		  .input_sync(1'b0),
		  .input_sync_mode(1'b0),
		  .intr_mode(2'b00),
		  .invert_in_clock(0),
		  .invert_in_clock_en(0),
		  .invert_in_reset(0),
		  .invert_out_clock(0),
		  .invert_out_clock_en(0),
		  .invert_out_reset(0),
		  .io_voltage(""),
		  .layout_mode("CONTIGUOUS"),
		  .oe_conn(1'b0),
		  .oe_reset(0),
		  .oe_sync(1'b0),
		  .output_clk_en(0),
		  .output_clock_mode(1'b0),
		  .output_conn(1'b1),
		  .output_mode(1'b0),
		  .output_reset(0),
		  .output_sync(1'b0),
		  .pa_in_clock(-1),
		  .pa_in_clock_en(-1),
		  .pa_in_reset(-1),
		  .pa_out_clock(-1),
		  .pa_out_clock_en(-1),
		  .pa_out_reset(-1),
		  .pin_aliases(""),
		  .pin_mode("B"),
		  .por_state(4),
		  .sio_group_cnt(0),
		  .sio_hyst(1'b1),
		  .sio_ibuf(""),
		  .sio_info(2'b00),
		  .sio_obuf(""),
		  .sio_refsel(""),
		  .sio_vtrip(""),
		  .slew_rate(1'b0),
		  .spanning(0),
		  .use_annotation(1'b0),
		  .vtrip(2'b00),
		  .width(1),
		  .ovt_hyst_trim(1'b0),
		  .ovt_needed(1'b0),
		  .ovt_slew_control(2'b00),
		  .input_buffer_sel(2'b00))
		tx
		 (.oe(tmpOE__tx_net),
		  .y({Net_1062}),
		  .fb({tmpFB_0__tx_net[0:0]}),
		  .io({tmpIO_0__tx_net[0:0]}),
		  .siovref(tmpSIOVREF__tx_net),
		  .interrupt({tmpINTERRUPT_0__tx_net[0:0]}),
		  .in_clock({1'b0}),
		  .in_clock_en({1'b1}),
		  .in_reset({1'b0}),
		  .out_clock({1'b0}),
		  .out_clock_en({1'b1}),
		  .out_reset({1'b0}));
	assign tmpOE__tx_net = (`CYDEV_CHIP_MEMBER_USED == `CYDEV_CHIP_MEMBER_3A && `CYDEV_CHIP_REVISION_USED < `CYDEV_CHIP_REVISION_3A_ES3) ? ~{1'b1} : {1'b1};
    ZeroTerminal ZeroTerminal_7 (
        .z(Net_1099));
    assign Net_1258 = Net_847 | Net_1099;
	wire [0:0] tmpOE__rx_net;
	wire [0:0] tmpIO_0__rx_net;
	wire [0:0] tmpINTERRUPT_0__rx_net;
	electrical [0:0] tmpSIOVREF__rx_net;
	cy_psoc3_pins_v1_10
		#(.id("43ec2fa1-bf22-4b71-9477-b6ca7b97f0b0/78e33e5d-45ea-4b75-88d5-73274e8a7ce4"),
		  .drive_mode(3'b001),
		  .ibuf_enabled(1'b1),
		  .init_dr_st(1'b0),
		  .input_clk_en(0),
		  .input_sync(1'b0),
		  .input_sync_mode(1'b0),
		  .intr_mode(2'b00),
		  .invert_in_clock(0),
		  .invert_in_clock_en(0),
		  .invert_in_reset(0),
		  .invert_out_clock(0),
		  .invert_out_clock_en(0),
		  .invert_out_reset(0),
		  .io_voltage(""),
		  .layout_mode("CONTIGUOUS"),
		  .oe_conn(1'b0),
		  .oe_reset(0),
		  .oe_sync(1'b0),
		  .output_clk_en(0),
		  .output_clock_mode(1'b0),
		  .output_conn(1'b0),
		  .output_mode(1'b0),
		  .output_reset(0),
		  .output_sync(1'b0),
		  .pa_in_clock(-1),
		  .pa_in_clock_en(-1),
		  .pa_in_reset(-1),
		  .pa_out_clock(-1),
		  .pa_out_clock_en(-1),
		  .pa_out_reset(-1),
		  .pin_aliases(""),
		  .pin_mode("I"),
		  .por_state(4),
		  .sio_group_cnt(0),
		  .sio_hyst(1'b1),
		  .sio_ibuf(""),
		  .sio_info(2'b00),
		  .sio_obuf(""),
		  .sio_refsel(""),
		  .sio_vtrip(""),
		  .slew_rate(1'b0),
		  .spanning(0),
		  .use_annotation(1'b0),
		  .vtrip(2'b00),
		  .width(1),
		  .ovt_hyst_trim(1'b0),
		  .ovt_needed(1'b0),
		  .ovt_slew_control(2'b00),
		  .input_buffer_sel(2'b00))
		rx
		 (.oe(tmpOE__rx_net),
		  .y({1'b0}),
		  .fb({Net_1197}),
		  .io({tmpIO_0__rx_net[0:0]}),
		  .siovref(tmpSIOVREF__rx_net),
		  .interrupt({tmpINTERRUPT_0__rx_net[0:0]}),
		  .in_clock({1'b0}),
		  .in_clock_en({1'b1}),
		  .in_reset({1'b0}),
		  .out_clock({1'b0}),
		  .out_clock_en({1'b1}),
		  .out_reset({1'b0}));
	assign tmpOE__rx_net = (`CYDEV_CHIP_MEMBER_USED == `CYDEV_CHIP_MEMBER_3A && `CYDEV_CHIP_REVISION_USED < `CYDEV_CHIP_REVISION_3A_ES3) ? ~{1'b1} : {1'b1};
	// cts_VM (cy_virtualmux_v1_0)
	assign Net_1175 = Net_747;
    cy_m0s8_scb_v2_0 SCB (
        .rx(Net_654),
        .miso_m(Net_663),
        .select_m(ss[3:0]),
        .sclk_m(Net_1059),
        .mosi_s(Net_909),
        .select_s(Net_652),
        .sclk_s(Net_990),
        .mosi_m(Net_1061),
        .scl(Net_580),
        .sda(Net_581),
        .tx(Net_1062),
        .miso_s(Net_1055),
        .interrupt(interrupt),
        .cts(Net_1175),
        .rts(Net_1053),
        .tx_req(tx_tr_out),
        .rx_req(rx_tr_out),
        .clock(Net_1170));
    defparam SCB.scb_mode = 2;
    ZeroTerminal ZeroTerminal_6 (
        .z(Net_747));
	// Device_VM1 (cy_virtualmux_v1_0)
	assign Net_547 = Net_1090;
	// Device_VM5 (cy_virtualmux_v1_0)
	assign Net_891 = Net_1089;
	// Device_VM2 (cy_virtualmux_v1_0)
	assign Net_1001 = Net_1086;
	// Device_VM3 (cy_virtualmux_v1_0)
	assign Net_899 = Net_916;
	// Device_VM4 (cy_virtualmux_v1_0)
	assign uncfg_rx_irq = Net_1000;
endmodule