module v95;
  integer signed; initial signed = 1;
endmodule