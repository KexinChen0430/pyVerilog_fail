module add_float32_float32_float32 (
                                      CLK, ce, inp, out
);
            parameter INSTANCE_NAME="INST";
  input wire CLK;
  input wire ce;
  input [63 : 0] inp;
  output [31 : 0] out;
   wire           clk;
   assign clk=CLK;
   wire [31:0]    a;
   wire [31:0]    b;
   wire [31:0]    result;
   assign a = inp[31:0];
   assign b = inp[63:32];
   assign out = result;
  wire \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.DSP.OP/OP/sign_op ;
  wire sig00000001;
  wire sig00000002;
  wire sig00000003;
  wire sig00000004;
  wire sig00000005;
  wire sig00000006;
  wire sig00000007;
  wire sig00000008;
  wire sig00000009;
  wire sig0000000a;
  wire sig0000000b;
  wire sig0000000c;
  wire sig0000000d;
  wire sig0000000e;
  wire sig0000000f;
  wire sig00000010;
  wire sig00000011;
  wire sig00000012;
  wire sig00000013;
  wire sig00000014;
  wire sig00000015;
  wire sig00000016;
  wire sig00000017;
  wire sig00000018;
  wire sig00000019;
  wire sig0000001a;
  wire sig0000001b;
  wire sig0000001c;
  wire sig0000001d;
  wire sig0000001e;
  wire sig0000001f;
  wire sig00000020;
  wire sig00000021;
  wire sig00000022;
  wire sig00000023;
  wire sig00000024;
  wire sig00000025;
  wire sig00000026;
  wire sig00000027;
  wire sig00000028;
  wire sig00000029;
  wire sig0000002a;
  wire sig0000002b;
  wire sig0000002c;
  wire sig0000002d;
  wire sig0000002e;
  wire sig0000002f;
  wire sig00000030;
  wire sig00000031;
  wire sig00000032;
  wire sig00000033;
  wire sig00000034;
  wire sig00000035;
  wire sig00000036;
  wire sig00000037;
  wire sig00000038;
  wire sig00000039;
  wire sig0000003a;
  wire sig0000003b;
  wire sig0000003c;
  wire sig0000003d;
  wire sig0000003e;
  wire sig0000003f;
  wire sig00000040;
  wire sig00000041;
  wire sig00000042;
  wire sig00000043;
  wire sig00000044;
  wire sig00000045;
  wire sig00000046;
  wire sig00000047;
  wire sig00000048;
  wire sig00000049;
  wire sig0000004a;
  wire sig0000004b;
  wire sig0000004c;
  wire sig0000004d;
  wire sig0000004e;
  wire sig0000004f;
  wire sig00000050;
  wire sig00000051;
  wire sig00000052;
  wire sig00000053;
  wire sig00000054;
  wire sig00000055;
  wire sig00000056;
  wire sig00000057;
  wire sig00000058;
  wire sig00000059;
  wire sig0000005a;
  wire sig0000005b;
  wire sig0000005c;
  wire sig0000005d;
  wire sig0000005e;
  wire sig0000005f;
  wire sig00000060;
  wire sig00000061;
  wire sig00000062;
  wire sig00000063;
  wire sig00000064;
  wire sig00000065;
  wire sig00000066;
  wire sig00000067;
  wire sig00000068;
  wire sig00000069;
  wire sig0000006a;
  wire sig0000006b;
  wire sig0000006c;
  wire sig0000006d;
  wire sig0000006e;
  wire sig0000006f;
  wire sig00000070;
  wire sig00000071;
  wire sig00000072;
  wire sig00000073;
  wire sig00000074;
  wire sig00000075;
  wire sig00000076;
  wire sig00000077;
  wire sig00000078;
  wire sig00000079;
  wire sig0000007a;
  wire sig0000007b;
  wire sig0000007c;
  wire sig0000007d;
  wire sig0000007e;
  wire sig0000007f;
  wire sig00000080;
  wire sig00000081;
  wire sig00000082;
  wire sig00000083;
  wire sig00000084;
  wire sig00000085;
  wire sig00000086;
  wire sig00000087;
  wire sig00000088;
  wire sig00000089;
  wire sig0000008a;
  wire sig0000008b;
  wire sig0000008c;
  wire sig0000008d;
  wire sig0000008e;
  wire sig0000008f;
  wire sig00000090;
  wire sig00000091;
  wire sig00000092;
  wire sig00000093;
  wire sig00000094;
  wire sig00000095;
  wire sig00000096;
  wire sig00000097;
  wire sig00000098;
  wire sig00000099;
  wire sig0000009a;
  wire sig0000009b;
  wire sig0000009c;
  wire sig0000009d;
  wire sig0000009e;
  wire sig0000009f;
  wire sig000000a0;
  wire sig000000a1;
  wire sig000000a2;
  wire sig000000a3;
  wire sig000000a4;
  wire sig000000a5;
  wire sig000000a6;
  wire sig000000a7;
  wire sig000000a8;
  wire sig000000a9;
  wire sig000000aa;
  wire sig000000ab;
  wire sig000000ac;
  wire sig000000ad;
  wire sig000000ae;
  wire sig000000af;
  wire sig000000b0;
  wire sig000000b1;
  wire sig000000b2;
  wire sig000000b3;
  wire sig000000b4;
  wire sig000000b5;
  wire sig000000b6;
  wire sig000000b7;
  wire sig000000b8;
  wire sig000000b9;
  wire sig000000ba;
  wire sig000000bb;
  wire sig000000bc;
  wire sig000000bd;
  wire sig000000be;
  wire sig000000bf;
  wire sig000000c0;
  wire sig000000c1;
  wire sig000000c2;
  wire sig000000c3;
  wire sig000000c4;
  wire sig000000c5;
  wire sig000000c6;
  wire sig000000c7;
  wire sig000000c8;
  wire sig000000c9;
  wire sig000000ca;
  wire sig000000cb;
  wire sig000000cc;
  wire sig000000cd;
  wire sig000000ce;
  wire sig000000cf;
  wire sig000000d0;
  wire sig000000d1;
  wire sig000000d2;
  wire sig000000d3;
  wire sig000000d4;
  wire sig000000d5;
  wire sig000000d6;
  wire sig000000d7;
  wire sig000000d8;
  wire sig000000d9;
  wire sig000000da;
  wire sig000000db;
  wire sig000000dc;
  wire sig000000dd;
  wire sig000000de;
  wire sig000000df;
  wire sig000000e0;
  wire sig000000e1;
  wire sig000000e2;
  wire sig000000e3;
  wire sig000000e4;
  wire sig000000e5;
  wire sig000000e6;
  wire sig000000e7;
  wire sig000000e8;
  wire sig000000e9;
  wire sig000000ea;
  wire sig000000eb;
  wire sig000000ec;
  wire sig000000ed;
  wire sig000000ee;
  wire sig000000ef;
  wire sig000000f0;
  wire sig000000f1;
  wire sig000000f2;
  wire sig000000f3;
  wire sig000000f4;
  wire sig000000f5;
  wire sig000000f6;
  wire sig000000f7;
  wire sig000000f8;
  wire sig000000f9;
  wire sig000000fa;
  wire sig000000fb;
  wire sig000000fc;
  wire sig000000fd;
  wire sig000000fe;
  wire sig000000ff;
  wire sig00000100;
  wire sig00000101;
  wire sig00000102;
  wire sig00000103;
  wire sig00000104;
  wire sig00000105;
  wire sig00000106;
  wire sig00000107;
  wire sig00000108;
  wire sig00000109;
  wire sig0000010a;
  wire sig0000010b;
  wire sig0000010c;
  wire sig0000010d;
  wire sig0000010e;
  wire sig0000010f;
  wire sig00000110;
  wire sig00000111;
  wire sig00000112;
  wire sig00000113;
  wire sig00000114;
  wire sig00000115;
  wire sig00000116;
  wire sig00000117;
  wire sig00000118;
  wire sig00000119;
  wire sig0000011a;
  wire sig0000011b;
  wire sig0000011c;
  wire sig0000011d;
  wire sig0000011e;
  wire sig0000011f;
  wire sig00000120;
  wire sig00000121;
  wire sig00000122;
  wire sig00000123;
  wire sig00000124;
  wire sig00000125;
  wire sig00000126;
  wire sig00000127;
  wire sig00000128;
  wire sig00000129;
  wire sig0000012a;
  wire sig0000012b;
  wire sig0000012c;
  wire sig0000012d;
  wire sig0000012e;
  wire sig0000012f;
  wire sig00000130;
  wire sig00000131;
  wire sig00000132;
  wire sig00000133;
  wire sig00000134;
  wire sig00000135;
  wire sig00000136;
  wire sig00000137;
  wire sig00000138;
  wire sig00000139;
  wire sig0000013a;
  wire sig0000013b;
  wire sig0000013c;
  wire sig0000013d;
  wire sig0000013e;
  wire sig0000013f;
  wire sig00000140;
  wire sig00000141;
  wire sig00000142;
  wire sig00000143;
  wire sig00000144;
  wire sig00000145;
  wire sig00000146;
  wire sig00000147;
  wire sig00000148;
  wire sig00000149;
  wire sig0000014a;
  wire sig0000014b;
  wire sig0000014c;
  wire sig0000014d;
  wire sig0000014e;
  wire sig0000014f;
  wire sig00000150;
  wire sig00000151;
  wire sig00000152;
  wire sig00000153;
  wire sig00000154;
  wire sig00000155;
  wire sig00000156;
  wire sig00000157;
  wire sig00000158;
  wire sig00000159;
  wire sig0000015a;
  wire sig0000015b;
  wire sig0000015c;
  wire sig0000015d;
  wire sig0000015e;
  wire sig0000015f;
  wire sig00000160;
  wire sig00000161;
  wire sig00000162;
  wire sig00000163;
  wire sig00000164;
  wire sig00000165;
  wire sig00000166;
  wire sig00000167;
  wire sig00000168;
  wire sig00000169;
  wire sig0000016a;
  wire sig0000016b;
  wire sig0000016c;
  wire sig0000016d;
  wire sig0000016e;
  wire sig0000016f;
  wire sig00000170;
  wire sig00000171;
  wire sig00000172;
  wire sig00000173;
  wire sig00000174;
  wire sig00000175;
  wire sig00000176;
  wire sig00000177;
  wire sig00000178;
  wire sig00000179;
  wire sig0000017a;
  wire sig0000017b;
  wire sig0000017c;
  wire sig0000017d;
  wire sig0000017e;
  wire sig0000017f;
  wire sig00000180;
  wire sig00000181;
  wire sig00000182;
  wire sig00000183;
  wire sig00000184;
  wire sig00000185;
  wire sig00000186;
  wire sig00000187;
  wire sig00000188;
  wire sig00000189;
  wire sig0000018a;
  wire sig0000018b;
  wire sig0000018c;
  wire sig0000018d;
  wire sig0000018e;
  wire sig0000018f;
  wire sig00000190;
  wire sig00000191;
  wire sig00000192;
  wire sig00000193;
  wire sig00000194;
  wire sig00000195;
  wire sig00000196;
  wire sig00000197;
  wire sig00000198;
  wire sig00000199;
  wire sig0000019a;
  wire sig0000019b;
  wire sig0000019c;
  wire sig0000019d;
  wire sig0000019e;
  wire sig0000019f;
  wire sig000001a0;
  wire sig000001a1;
  wire sig000001a2;
  wire sig000001a3;
  wire sig000001a4;
  wire sig000001a5;
  wire sig000001a6;
  wire sig000001a7;
  wire sig000001a8;
  wire sig000001a9;
  wire sig000001aa;
  wire sig000001ab;
  wire sig000001ac;
  wire sig000001ad;
  wire sig000001ae;
  wire sig000001af;
  wire sig000001b0;
  wire sig000001b1;
  wire sig000001b2;
  wire sig000001b3;
  wire sig000001b4;
  wire sig000001b5;
  wire sig000001b6;
  wire sig000001b7;
  wire sig000001b8;
  wire sig000001b9;
  wire sig000001ba;
  wire sig000001bb;
  wire sig000001bc;
  wire sig000001bd;
  wire sig000001be;
  wire sig000001bf;
  wire sig000001c0;
  wire sig000001c1;
  wire sig000001c2;
  wire sig000001c3;
  wire sig000001c4;
  wire sig000001c5;
  wire sig000001c6;
  wire sig000001c7;
  wire sig000001c8;
  wire sig000001c9;
  wire sig000001ca;
  wire sig000001cb;
  wire sig000001cc;
  wire sig000001cd;
  wire sig000001ce;
  wire sig000001cf;
  wire sig000001d0;
  wire sig000001d1;
  wire sig000001d2;
  wire sig000001d3;
  wire sig000001d4;
  wire sig000001d5;
  wire sig000001d6;
  wire sig000001d7;
  wire sig000001d8;
  wire sig000001d9;
  wire sig000001da;
  wire sig000001db;
  wire sig000001dc;
  wire sig000001dd;
  wire sig000001de;
  wire sig000001df;
  wire sig000001e0;
  wire sig000001e1;
  wire sig000001e2;
  wire sig000001e3;
  wire sig000001e4;
  wire sig000001e5;
  wire sig000001e6;
  wire sig000001e7;
  wire sig000001e8;
  wire sig000001e9;
  wire sig000001ea;
  wire sig000001eb;
  wire sig000001ec;
  wire sig000001ed;
  wire sig000001ee;
  wire sig000001ef;
  wire sig000001f0;
  wire sig000001f1;
  wire sig000001f2;
  wire sig000001f3;
  wire sig000001f4;
  wire sig000001f5;
  wire sig000001f6;
  wire sig000001f7;
  wire sig000001f8;
  wire sig000001f9;
  wire sig000001fa;
  wire sig000001fb;
  wire sig000001fc;
  wire sig000001fd;
  wire sig000001fe;
  wire sig000001ff;
  wire sig00000200;
  wire sig00000201;
  wire sig00000202;
  wire sig00000203;
  wire sig00000204;
  wire sig00000205;
  wire sig00000206;
  wire sig00000207;
  wire sig00000208;
  wire sig00000209;
  wire sig0000020a;
  wire sig0000020b;
  wire sig0000020c;
  wire sig0000020d;
  wire sig0000020e;
  wire sig0000020f;
  wire sig00000210;
  wire sig00000211;
  wire sig00000212;
  wire sig00000213;
  wire sig00000214;
  wire sig00000215;
  wire sig00000216;
  wire sig00000217;
  wire sig00000218;
  wire sig00000219;
  wire sig0000021a;
  wire sig0000021b;
  wire sig0000021c;
  wire sig0000021d;
  wire sig0000021e;
  wire sig0000021f;
  wire sig00000220;
  wire sig00000221;
  wire sig00000222;
  wire sig00000223;
  wire sig00000224;
  wire sig00000225;
  wire sig00000226;
  wire sig00000227;
  wire sig00000228;
  wire sig00000229;
  wire sig0000022a;
  wire sig0000022b;
  wire sig0000022c;
  wire sig0000022d;
  wire sig0000022e;
  wire sig0000022f;
  wire sig00000230;
  wire sig00000231;
  wire sig00000232;
  wire sig00000233;
  wire sig00000234;
  wire sig00000235;
  wire sig00000236;
  wire sig00000237;
  wire sig00000238;
  wire sig00000239;
  wire sig0000023a;
  wire sig0000023b;
  wire sig0000023c;
  wire sig0000023d;
  wire sig0000023e;
  wire sig0000023f;
  wire sig00000240;
  wire sig00000241;
  wire sig00000242;
  wire sig00000243;
  wire sig00000244;
  wire sig00000245;
  wire sig00000246;
  wire sig00000247;
  wire sig00000248;
  wire sig00000249;
  wire sig0000024a;
  wire sig0000024b;
  wire sig0000024c;
  wire sig0000024d;
  wire sig0000024e;
  wire sig0000024f;
  wire sig00000250;
  wire sig00000251;
  wire sig00000252;
  wire sig00000253;
  wire sig00000254;
  wire sig00000255;
  wire sig00000256;
  wire sig00000257;
  wire sig00000258;
  wire sig00000259;
  wire sig0000025a;
  wire sig0000025b;
  wire sig0000025c;
  wire sig0000025d;
  wire sig0000025e;
  wire sig0000025f;
  wire sig00000260;
  wire sig00000261;
  wire sig00000262;
  wire sig00000263;
  wire sig00000264;
  wire sig00000265;
  wire sig00000266;
  wire sig00000267;
  wire sig00000268;
  wire sig00000269;
  wire sig0000026a;
  wire sig0000026b;
  wire sig0000026c;
  wire sig0000026d;
  wire sig0000026e;
  wire sig0000026f;
  wire sig00000270;
  wire sig00000271;
  wire sig00000272;
  wire sig00000273;
  wire sig00000274;
  wire sig00000275;
  wire sig00000276;
  wire sig00000277;
  wire sig00000278;
  wire sig00000279;
  wire sig0000027a;
  wire sig0000027b;
  wire sig0000027c;
  wire sig0000027d;
  wire sig0000027e;
  wire sig0000027f;
  wire sig00000280;
  wire sig00000281;
  wire sig00000282;
  wire sig00000283;
  wire sig00000284;
  wire sig00000285;
  wire sig00000286;
  wire sig00000287;
  wire sig00000288;
  wire sig00000289;
  wire sig0000028a;
  wire sig0000028b;
  wire sig0000028c;
  wire sig0000028d;
  wire sig0000028e;
  wire sig0000028f;
  wire sig00000290;
  wire sig00000291;
  wire sig00000292;
  wire sig00000293;
  wire sig00000294;
  wire sig00000295;
  wire sig00000296;
  wire sig00000297;
  wire sig00000298;
  wire sig00000299;
  wire sig0000029a;
  wire sig0000029b;
  wire sig0000029c;
  wire sig0000029d;
  wire sig0000029e;
  wire sig0000029f;
  wire sig000002a0;
  wire sig000002a1;
  wire sig000002a2;
  wire sig000002a3;
  wire sig000002a4;
  wire sig000002a5;
  wire sig000002a6;
  wire sig000002a7;
  wire sig000002a8;
  wire sig000002a9;
  wire sig000002aa;
  wire sig000002ab;
  wire sig000002ac;
  wire sig000002ad;
  wire sig000002ae;
  wire sig000002af;
  wire sig000002b0;
  wire sig000002b1;
  wire sig000002b2;
  wire sig000002b3;
  wire sig000002b4;
  wire sig000002b5;
  wire sig000002b6;
  wire sig000002b7;
  wire sig000002b8;
  wire sig000002b9;
  wire sig000002ba;
  wire sig000002bb;
  wire sig000002bc;
  wire sig000002bd;
  wire sig000002be;
  wire sig000002bf;
  wire sig000002c0;
  wire sig000002c1;
  wire sig000002c2;
  wire sig000002c3;
  wire sig000002c4;
  wire sig000002c5;
  wire sig000002c6;
  wire sig000002c7;
  wire sig000002c8;
  wire sig000002c9;
  wire sig000002ca;
  wire sig000002cb;
  wire sig000002cc;
  wire sig000002cd;
  wire sig000002ce;
  wire sig000002cf;
  wire sig000002d0;
  wire sig000002d1;
  wire sig000002d2;
  wire sig000002d3;
  wire sig000002d4;
  wire sig000002d5;
  wire sig000002d6;
  wire sig000002d7;
  wire sig000002d8;
  wire sig000002d9;
  wire sig000002da;
  wire sig000002db;
  wire sig000002dc;
  wire sig000002dd;
  wire sig000002de;
  wire sig000002df;
  wire sig000002e0;
  wire sig000002e1;
  wire sig000002e2;
  wire sig000002e3;
  wire sig000002e4;
  wire NLW_blk00000082_O_UNCONNECTED;
  wire NLW_blk000000cb_O_UNCONNECTED;
  wire NLW_blk000002a3_Q15_UNCONNECTED;
  wire NLW_blk000002a5_Q15_UNCONNECTED;
  wire NLW_blk000002a7_Q15_UNCONNECTED;
  wire NLW_blk000002a9_Q15_UNCONNECTED;
  wire NLW_blk000002ab_Q15_UNCONNECTED;
  wire NLW_blk000002ad_Q15_UNCONNECTED;
  wire NLW_blk000002af_Q15_UNCONNECTED;
  wire NLW_blk000002b1_Q15_UNCONNECTED;
  wire NLW_blk000002b3_Q15_UNCONNECTED;
  wire NLW_blk000002b5_Q15_UNCONNECTED;
  wire NLW_blk000002b7_Q15_UNCONNECTED;
  wire NLW_blk000002b9_Q15_UNCONNECTED;
  wire NLW_blk000002bb_Q15_UNCONNECTED;
  wire NLW_blk000002bd_Q15_UNCONNECTED;
  wire NLW_blk000002bf_PATTERNBDETECT_UNCONNECTED;
  wire NLW_blk000002bf_MULTSIGNOUT_UNCONNECTED;
  wire NLW_blk000002bf_CARRYCASCOUT_UNCONNECTED;
  wire NLW_blk000002bf_UNDERFLOW_UNCONNECTED;
  wire NLW_blk000002bf_OVERFLOW_UNCONNECTED;
  wire \NLW_blk000002bf_ACOUT<29>_UNCONNECTED ;
  wire \NLW_blk000002bf_ACOUT<28>_UNCONNECTED ;
  wire \NLW_blk000002bf_ACOUT<27>_UNCONNECTED ;
  wire \NLW_blk000002bf_ACOUT<26>_UNCONNECTED ;
  wire \NLW_blk000002bf_ACOUT<25>_UNCONNECTED ;
  wire \NLW_blk000002bf_ACOUT<24>_UNCONNECTED ;
  wire \NLW_blk000002bf_ACOUT<23>_UNCONNECTED ;
  wire \NLW_blk000002bf_ACOUT<22>_UNCONNECTED ;
  wire \NLW_blk000002bf_ACOUT<21>_UNCONNECTED ;
  wire \NLW_blk000002bf_ACOUT<20>_UNCONNECTED ;
  wire \NLW_blk000002bf_ACOUT<19>_UNCONNECTED ;
  wire \NLW_blk000002bf_ACOUT<18>_UNCONNECTED ;
  wire \NLW_blk000002bf_ACOUT<17>_UNCONNECTED ;
  wire \NLW_blk000002bf_ACOUT<16>_UNCONNECTED ;
  wire \NLW_blk000002bf_ACOUT<15>_UNCONNECTED ;
  wire \NLW_blk000002bf_ACOUT<14>_UNCONNECTED ;
  wire \NLW_blk000002bf_ACOUT<13>_UNCONNECTED ;
  wire \NLW_blk000002bf_ACOUT<12>_UNCONNECTED ;
  wire \NLW_blk000002bf_ACOUT<11>_UNCONNECTED ;
  wire \NLW_blk000002bf_ACOUT<10>_UNCONNECTED ;
  wire \NLW_blk000002bf_ACOUT<9>_UNCONNECTED ;
  wire \NLW_blk000002bf_ACOUT<8>_UNCONNECTED ;
  wire \NLW_blk000002bf_ACOUT<7>_UNCONNECTED ;
  wire \NLW_blk000002bf_ACOUT<6>_UNCONNECTED ;
  wire \NLW_blk000002bf_ACOUT<5>_UNCONNECTED ;
  wire \NLW_blk000002bf_ACOUT<4>_UNCONNECTED ;
  wire \NLW_blk000002bf_ACOUT<3>_UNCONNECTED ;
  wire \NLW_blk000002bf_ACOUT<2>_UNCONNECTED ;
  wire \NLW_blk000002bf_ACOUT<1>_UNCONNECTED ;
  wire \NLW_blk000002bf_ACOUT<0>_UNCONNECTED ;
  wire \NLW_blk000002bf_CARRYOUT<3>_UNCONNECTED ;
  wire \NLW_blk000002bf_CARRYOUT<2>_UNCONNECTED ;
  wire \NLW_blk000002bf_CARRYOUT<1>_UNCONNECTED ;
  wire \NLW_blk000002bf_CARRYOUT<0>_UNCONNECTED ;
  wire \NLW_blk000002bf_BCOUT<17>_UNCONNECTED ;
  wire \NLW_blk000002bf_BCOUT<16>_UNCONNECTED ;
  wire \NLW_blk000002bf_BCOUT<15>_UNCONNECTED ;
  wire \NLW_blk000002bf_BCOUT<14>_UNCONNECTED ;
  wire \NLW_blk000002bf_BCOUT<13>_UNCONNECTED ;
  wire \NLW_blk000002bf_BCOUT<12>_UNCONNECTED ;
  wire \NLW_blk000002bf_BCOUT<11>_UNCONNECTED ;
  wire \NLW_blk000002bf_BCOUT<10>_UNCONNECTED ;
  wire \NLW_blk000002bf_BCOUT<9>_UNCONNECTED ;
  wire \NLW_blk000002bf_BCOUT<8>_UNCONNECTED ;
  wire \NLW_blk000002bf_BCOUT<7>_UNCONNECTED ;
  wire \NLW_blk000002bf_BCOUT<6>_UNCONNECTED ;
  wire \NLW_blk000002bf_BCOUT<5>_UNCONNECTED ;
  wire \NLW_blk000002bf_BCOUT<4>_UNCONNECTED ;
  wire \NLW_blk000002bf_BCOUT<3>_UNCONNECTED ;
  wire \NLW_blk000002bf_BCOUT<2>_UNCONNECTED ;
  wire \NLW_blk000002bf_BCOUT<1>_UNCONNECTED ;
  wire \NLW_blk000002bf_BCOUT<0>_UNCONNECTED ;
  wire \NLW_blk000002bf_P<47>_UNCONNECTED ;
  wire \NLW_blk000002bf_P<46>_UNCONNECTED ;
  wire \NLW_blk000002bf_P<45>_UNCONNECTED ;
  wire \NLW_blk000002bf_P<44>_UNCONNECTED ;
  wire \NLW_blk000002bf_P<43>_UNCONNECTED ;
  wire \NLW_blk000002bf_P<42>_UNCONNECTED ;
  wire \NLW_blk000002bf_P<41>_UNCONNECTED ;
  wire \NLW_blk000002bf_P<40>_UNCONNECTED ;
  wire \NLW_blk000002bf_PCOUT<47>_UNCONNECTED ;
  wire \NLW_blk000002bf_PCOUT<46>_UNCONNECTED ;
  wire \NLW_blk000002bf_PCOUT<45>_UNCONNECTED ;
  wire \NLW_blk000002bf_PCOUT<44>_UNCONNECTED ;
  wire \NLW_blk000002bf_PCOUT<43>_UNCONNECTED ;
  wire \NLW_blk000002bf_PCOUT<42>_UNCONNECTED ;
  wire \NLW_blk000002bf_PCOUT<41>_UNCONNECTED ;
  wire \NLW_blk000002bf_PCOUT<40>_UNCONNECTED ;
  wire \NLW_blk000002bf_PCOUT<39>_UNCONNECTED ;
  wire \NLW_blk000002bf_PCOUT<38>_UNCONNECTED ;
  wire \NLW_blk000002bf_PCOUT<37>_UNCONNECTED ;
  wire \NLW_blk000002bf_PCOUT<36>_UNCONNECTED ;
  wire \NLW_blk000002bf_PCOUT<35>_UNCONNECTED ;
  wire \NLW_blk000002bf_PCOUT<34>_UNCONNECTED ;
  wire \NLW_blk000002bf_PCOUT<33>_UNCONNECTED ;
  wire \NLW_blk000002bf_PCOUT<32>_UNCONNECTED ;
  wire \NLW_blk000002bf_PCOUT<31>_UNCONNECTED ;
  wire \NLW_blk000002bf_PCOUT<30>_UNCONNECTED ;
  wire \NLW_blk000002bf_PCOUT<29>_UNCONNECTED ;
  wire \NLW_blk000002bf_PCOUT<28>_UNCONNECTED ;
  wire \NLW_blk000002bf_PCOUT<27>_UNCONNECTED ;
  wire \NLW_blk000002bf_PCOUT<26>_UNCONNECTED ;
  wire \NLW_blk000002bf_PCOUT<25>_UNCONNECTED ;
  wire \NLW_blk000002bf_PCOUT<24>_UNCONNECTED ;
  wire \NLW_blk000002bf_PCOUT<23>_UNCONNECTED ;
  wire \NLW_blk000002bf_PCOUT<22>_UNCONNECTED ;
  wire \NLW_blk000002bf_PCOUT<21>_UNCONNECTED ;
  wire \NLW_blk000002bf_PCOUT<20>_UNCONNECTED ;
  wire \NLW_blk000002bf_PCOUT<19>_UNCONNECTED ;
  wire \NLW_blk000002bf_PCOUT<18>_UNCONNECTED ;
  wire \NLW_blk000002bf_PCOUT<17>_UNCONNECTED ;
  wire \NLW_blk000002bf_PCOUT<16>_UNCONNECTED ;
  wire \NLW_blk000002bf_PCOUT<15>_UNCONNECTED ;
  wire \NLW_blk000002bf_PCOUT<14>_UNCONNECTED ;
  wire \NLW_blk000002bf_PCOUT<13>_UNCONNECTED ;
  wire \NLW_blk000002bf_PCOUT<12>_UNCONNECTED ;
  wire \NLW_blk000002bf_PCOUT<11>_UNCONNECTED ;
  wire \NLW_blk000002bf_PCOUT<10>_UNCONNECTED ;
  wire \NLW_blk000002bf_PCOUT<9>_UNCONNECTED ;
  wire \NLW_blk000002bf_PCOUT<8>_UNCONNECTED ;
  wire \NLW_blk000002bf_PCOUT<7>_UNCONNECTED ;
  wire \NLW_blk000002bf_PCOUT<6>_UNCONNECTED ;
  wire \NLW_blk000002bf_PCOUT<5>_UNCONNECTED ;
  wire \NLW_blk000002bf_PCOUT<4>_UNCONNECTED ;
  wire \NLW_blk000002bf_PCOUT<3>_UNCONNECTED ;
  wire \NLW_blk000002bf_PCOUT<2>_UNCONNECTED ;
  wire \NLW_blk000002bf_PCOUT<1>_UNCONNECTED ;
  wire \NLW_blk000002bf_PCOUT<0>_UNCONNECTED ;
  wire \NLW_blk000002c0_P<26>_UNCONNECTED ;
  wire NLW_blk000002c0_PATTERNBDETECT_UNCONNECTED;
  wire NLW_blk000002c0_MULTSIGNOUT_UNCONNECTED;
  wire NLW_blk000002c0_CARRYCASCOUT_UNCONNECTED;
  wire NLW_blk000002c0_UNDERFLOW_UNCONNECTED;
  wire NLW_blk000002c0_PATTERNDETECT_UNCONNECTED;
  wire NLW_blk000002c0_OVERFLOW_UNCONNECTED;
  wire \NLW_blk000002c0_ACOUT<29>_UNCONNECTED ;
  wire \NLW_blk000002c0_ACOUT<28>_UNCONNECTED ;
  wire \NLW_blk000002c0_ACOUT<27>_UNCONNECTED ;
  wire \NLW_blk000002c0_ACOUT<26>_UNCONNECTED ;
  wire \NLW_blk000002c0_ACOUT<25>_UNCONNECTED ;
  wire \NLW_blk000002c0_ACOUT<24>_UNCONNECTED ;
  wire \NLW_blk000002c0_ACOUT<23>_UNCONNECTED ;
  wire \NLW_blk000002c0_ACOUT<22>_UNCONNECTED ;
  wire \NLW_blk000002c0_ACOUT<21>_UNCONNECTED ;
  wire \NLW_blk000002c0_ACOUT<20>_UNCONNECTED ;
  wire \NLW_blk000002c0_ACOUT<19>_UNCONNECTED ;
  wire \NLW_blk000002c0_ACOUT<18>_UNCONNECTED ;
  wire \NLW_blk000002c0_ACOUT<17>_UNCONNECTED ;
  wire \NLW_blk000002c0_ACOUT<16>_UNCONNECTED ;
  wire \NLW_blk000002c0_ACOUT<15>_UNCONNECTED ;
  wire \NLW_blk000002c0_ACOUT<14>_UNCONNECTED ;
  wire \NLW_blk000002c0_ACOUT<13>_UNCONNECTED ;
  wire \NLW_blk000002c0_ACOUT<12>_UNCONNECTED ;
  wire \NLW_blk000002c0_ACOUT<11>_UNCONNECTED ;
  wire \NLW_blk000002c0_ACOUT<10>_UNCONNECTED ;
  wire \NLW_blk000002c0_ACOUT<9>_UNCONNECTED ;
  wire \NLW_blk000002c0_ACOUT<8>_UNCONNECTED ;
  wire \NLW_blk000002c0_ACOUT<7>_UNCONNECTED ;
  wire \NLW_blk000002c0_ACOUT<6>_UNCONNECTED ;
  wire \NLW_blk000002c0_ACOUT<5>_UNCONNECTED ;
  wire \NLW_blk000002c0_ACOUT<4>_UNCONNECTED ;
  wire \NLW_blk000002c0_ACOUT<3>_UNCONNECTED ;
  wire \NLW_blk000002c0_ACOUT<2>_UNCONNECTED ;
  wire \NLW_blk000002c0_ACOUT<1>_UNCONNECTED ;
  wire \NLW_blk000002c0_ACOUT<0>_UNCONNECTED ;
  wire \NLW_blk000002c0_CARRYOUT<3>_UNCONNECTED ;
  wire \NLW_blk000002c0_CARRYOUT<2>_UNCONNECTED ;
  wire \NLW_blk000002c0_CARRYOUT<1>_UNCONNECTED ;
  wire \NLW_blk000002c0_CARRYOUT<0>_UNCONNECTED ;
  wire \NLW_blk000002c0_BCOUT<17>_UNCONNECTED ;
  wire \NLW_blk000002c0_BCOUT<16>_UNCONNECTED ;
  wire \NLW_blk000002c0_BCOUT<15>_UNCONNECTED ;
  wire \NLW_blk000002c0_BCOUT<14>_UNCONNECTED ;
  wire \NLW_blk000002c0_BCOUT<13>_UNCONNECTED ;
  wire \NLW_blk000002c0_BCOUT<12>_UNCONNECTED ;
  wire \NLW_blk000002c0_BCOUT<11>_UNCONNECTED ;
  wire \NLW_blk000002c0_BCOUT<10>_UNCONNECTED ;
  wire \NLW_blk000002c0_BCOUT<9>_UNCONNECTED ;
  wire \NLW_blk000002c0_BCOUT<8>_UNCONNECTED ;
  wire \NLW_blk000002c0_BCOUT<7>_UNCONNECTED ;
  wire \NLW_blk000002c0_BCOUT<6>_UNCONNECTED ;
  wire \NLW_blk000002c0_BCOUT<5>_UNCONNECTED ;
  wire \NLW_blk000002c0_BCOUT<4>_UNCONNECTED ;
  wire \NLW_blk000002c0_BCOUT<3>_UNCONNECTED ;
  wire \NLW_blk000002c0_BCOUT<2>_UNCONNECTED ;
  wire \NLW_blk000002c0_BCOUT<1>_UNCONNECTED ;
  wire \NLW_blk000002c0_BCOUT<0>_UNCONNECTED ;
  wire \NLW_blk000002c0_P<47>_UNCONNECTED ;
  wire \NLW_blk000002c0_P<46>_UNCONNECTED ;
  wire \NLW_blk000002c0_P<45>_UNCONNECTED ;
  wire \NLW_blk000002c0_P<44>_UNCONNECTED ;
  wire \NLW_blk000002c0_P<43>_UNCONNECTED ;
  wire \NLW_blk000002c0_P<42>_UNCONNECTED ;
  wire \NLW_blk000002c0_P<41>_UNCONNECTED ;
  wire \NLW_blk000002c0_P<40>_UNCONNECTED ;
  wire \NLW_blk000002c0_P<39>_UNCONNECTED ;
  wire \NLW_blk000002c0_P<38>_UNCONNECTED ;
  wire \NLW_blk000002c0_P<37>_UNCONNECTED ;
  wire \NLW_blk000002c0_P<36>_UNCONNECTED ;
  wire \NLW_blk000002c0_P<35>_UNCONNECTED ;
  wire \NLW_blk000002c0_P<25>_UNCONNECTED ;
  wire \NLW_blk000002c0_P<1>_UNCONNECTED ;
  wire \NLW_blk000002c0_P<0>_UNCONNECTED ;
  wire \NLW_blk000002c0_PCOUT<47>_UNCONNECTED ;
  wire \NLW_blk000002c0_PCOUT<46>_UNCONNECTED ;
  wire \NLW_blk000002c0_PCOUT<45>_UNCONNECTED ;
  wire \NLW_blk000002c0_PCOUT<44>_UNCONNECTED ;
  wire \NLW_blk000002c0_PCOUT<43>_UNCONNECTED ;
  wire \NLW_blk000002c0_PCOUT<42>_UNCONNECTED ;
  wire \NLW_blk000002c0_PCOUT<41>_UNCONNECTED ;
  wire \NLW_blk000002c0_PCOUT<40>_UNCONNECTED ;
  wire \NLW_blk000002c0_PCOUT<39>_UNCONNECTED ;
  wire \NLW_blk000002c0_PCOUT<38>_UNCONNECTED ;
  wire \NLW_blk000002c0_PCOUT<37>_UNCONNECTED ;
  wire \NLW_blk000002c0_PCOUT<36>_UNCONNECTED ;
  wire \NLW_blk000002c0_PCOUT<35>_UNCONNECTED ;
  wire \NLW_blk000002c0_PCOUT<34>_UNCONNECTED ;
  wire \NLW_blk000002c0_PCOUT<33>_UNCONNECTED ;
  wire \NLW_blk000002c0_PCOUT<32>_UNCONNECTED ;
  wire \NLW_blk000002c0_PCOUT<31>_UNCONNECTED ;
  wire \NLW_blk000002c0_PCOUT<30>_UNCONNECTED ;
  wire \NLW_blk000002c0_PCOUT<29>_UNCONNECTED ;
  wire \NLW_blk000002c0_PCOUT<28>_UNCONNECTED ;
  wire \NLW_blk000002c0_PCOUT<27>_UNCONNECTED ;
  wire \NLW_blk000002c0_PCOUT<26>_UNCONNECTED ;
  wire \NLW_blk000002c0_PCOUT<25>_UNCONNECTED ;
  wire \NLW_blk000002c0_PCOUT<24>_UNCONNECTED ;
  wire \NLW_blk000002c0_PCOUT<23>_UNCONNECTED ;
  wire \NLW_blk000002c0_PCOUT<22>_UNCONNECTED ;
  wire \NLW_blk000002c0_PCOUT<21>_UNCONNECTED ;
  wire \NLW_blk000002c0_PCOUT<20>_UNCONNECTED ;
  wire \NLW_blk000002c0_PCOUT<19>_UNCONNECTED ;
  wire \NLW_blk000002c0_PCOUT<18>_UNCONNECTED ;
  wire \NLW_blk000002c0_PCOUT<17>_UNCONNECTED ;
  wire \NLW_blk000002c0_PCOUT<16>_UNCONNECTED ;
  wire \NLW_blk000002c0_PCOUT<15>_UNCONNECTED ;
  wire \NLW_blk000002c0_PCOUT<14>_UNCONNECTED ;
  wire \NLW_blk000002c0_PCOUT<13>_UNCONNECTED ;
  wire \NLW_blk000002c0_PCOUT<12>_UNCONNECTED ;
  wire \NLW_blk000002c0_PCOUT<11>_UNCONNECTED ;
  wire \NLW_blk000002c0_PCOUT<10>_UNCONNECTED ;
  wire \NLW_blk000002c0_PCOUT<9>_UNCONNECTED ;
  wire \NLW_blk000002c0_PCOUT<8>_UNCONNECTED ;
  wire \NLW_blk000002c0_PCOUT<7>_UNCONNECTED ;
  wire \NLW_blk000002c0_PCOUT<6>_UNCONNECTED ;
  wire \NLW_blk000002c0_PCOUT<5>_UNCONNECTED ;
  wire \NLW_blk000002c0_PCOUT<4>_UNCONNECTED ;
  wire \NLW_blk000002c0_PCOUT<3>_UNCONNECTED ;
  wire \NLW_blk000002c0_PCOUT<2>_UNCONNECTED ;
  wire \NLW_blk000002c0_PCOUT<1>_UNCONNECTED ;
  wire \NLW_blk000002c0_PCOUT<0>_UNCONNECTED ;
  wire [7 : 0] \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.DSP.OP/OP/exp_op ;
  wire [22 : 0] \NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.DSP.OP/OP/mant_op ;
  assign
    result[31] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.DSP.OP/OP/sign_op ,
    result[30] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.DSP.OP/OP/exp_op [7],
    result[29] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.DSP.OP/OP/exp_op [6],
    result[28] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.DSP.OP/OP/exp_op [5],
    result[27] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.DSP.OP/OP/exp_op [4],
    result[26] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.DSP.OP/OP/exp_op [3],
    result[25] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.DSP.OP/OP/exp_op [2],
    result[24] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.DSP.OP/OP/exp_op [1],
    result[23] = \U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.DSP.OP/OP/exp_op [0],
    result[22] = \NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.DSP.OP/OP/mant_op [22],
    result[21] = \NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.DSP.OP/OP/mant_op [21],
    result[20] = \NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.DSP.OP/OP/mant_op [20],
    result[19] = \NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.DSP.OP/OP/mant_op [19],
    result[18] = \NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.DSP.OP/OP/mant_op [18],
    result[17] = \NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.DSP.OP/OP/mant_op [17],
    result[16] = \NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.DSP.OP/OP/mant_op [16],
    result[15] = \NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.DSP.OP/OP/mant_op [15],
    result[14] = \NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.DSP.OP/OP/mant_op [14],
    result[13] = \NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.DSP.OP/OP/mant_op [13],
    result[12] = \NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.DSP.OP/OP/mant_op [12],
    result[11] = \NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.DSP.OP/OP/mant_op [11],
    result[10] = \NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.DSP.OP/OP/mant_op [10],
    result[9] = \NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.DSP.OP/OP/mant_op [9],
    result[8] = \NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.DSP.OP/OP/mant_op [8],
    result[7] = \NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.DSP.OP/OP/mant_op [7],
    result[6] = \NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.DSP.OP/OP/mant_op [6],
    result[5] = \NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.DSP.OP/OP/mant_op [5],
    result[4] = \NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.DSP.OP/OP/mant_op [4],
    result[3] = \NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.DSP.OP/OP/mant_op [3],
    result[2] = \NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.DSP.OP/OP/mant_op [2],
    result[1] = \NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.DSP.OP/OP/mant_op [1],
    result[0] = \NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.DSP.OP/OP/mant_op [0];
  VCC   blk00000001 (
    .P(sig00000001)
  );
  GND   blk00000002 (
    .G(sig00000002)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000003 (
    .C(clk),
    .CE(ce),
    .D(sig000000af),
    .Q(sig0000000f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000004 (
    .C(clk),
    .CE(ce),
    .D(sig000000ae),
    .Q(sig0000000e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000005 (
    .C(clk),
    .CE(ce),
    .D(sig000000ad),
    .Q(sig0000000c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000006 (
    .C(clk),
    .CE(ce),
    .D(sig000000dd),
    .Q(sig00000010)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000007 (
    .C(clk),
    .CE(ce),
    .D(sig000000de),
    .Q(sig0000000d)
  );
  XORCY   blk00000008 (
    .CI(sig0000008c),
    .LI(sig00000001),
    .O(sig000000dc)
  );
  MUXCY   blk00000009 (
    .CI(sig0000008d),
    .DI(sig00000002),
    .S(sig00000001),
    .O(sig0000008c)
  );
  XORCY   blk0000000a (
    .CI(sig0000008f),
    .LI(sig0000008e),
    .O(sig000000db)
  );
  MUXCY   blk0000000b (
    .CI(sig0000008f),
    .DI(sig000000ea),
    .S(sig0000008e),
    .O(sig0000008d)
  );
  XORCY   blk0000000c (
    .CI(sig00000091),
    .LI(sig00000090),
    .O(sig000000da)
  );
  MUXCY   blk0000000d (
    .CI(sig00000091),
    .DI(sig000000e9),
    .S(sig00000090),
    .O(sig0000008f)
  );
  XORCY   blk0000000e (
    .CI(sig00000093),
    .LI(sig00000092),
    .O(sig000000d9)
  );
  MUXCY   blk0000000f (
    .CI(sig00000093),
    .DI(sig000000e8),
    .S(sig00000092),
    .O(sig00000091)
  );
  XORCY   blk00000010 (
    .CI(sig00000095),
    .LI(sig00000094),
    .O(sig000000d8)
  );
  MUXCY   blk00000011 (
    .CI(sig00000095),
    .DI(sig000000e7),
    .S(sig00000094),
    .O(sig00000093)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000012 (
    .I0(sig000000e7),
    .I1(sig00000067),
    .O(sig00000094)
  );
  XORCY   blk00000013 (
    .CI(sig00000097),
    .LI(sig00000096),
    .O(sig000000d7)
  );
  MUXCY   blk00000014 (
    .CI(sig00000097),
    .DI(sig000000e6),
    .S(sig00000096),
    .O(sig00000095)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000015 (
    .I0(sig000000e6),
    .I1(sig00000068),
    .O(sig00000096)
  );
  XORCY   blk00000016 (
    .CI(sig00000099),
    .LI(sig00000098),
    .O(sig000000d6)
  );
  MUXCY   blk00000017 (
    .CI(sig00000099),
    .DI(sig000000e5),
    .S(sig00000098),
    .O(sig00000097)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000018 (
    .I0(sig000000e5),
    .I1(sig00000069),
    .O(sig00000098)
  );
  XORCY   blk00000019 (
    .CI(sig0000009b),
    .LI(sig0000009a),
    .O(sig000000d5)
  );
  MUXCY   blk0000001a (
    .CI(sig0000009b),
    .DI(sig000000e4),
    .S(sig0000009a),
    .O(sig00000099)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk0000001b (
    .I0(sig000000e4),
    .I1(sig0000006a),
    .O(sig0000009a)
  );
  XORCY   blk0000001c (
    .CI(sig00000001),
    .LI(sig0000009c),
    .O(sig000000d4)
  );
  MUXCY   blk0000001d (
    .CI(sig00000001),
    .DI(sig000000e3),
    .S(sig0000009c),
    .O(sig0000009b)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk0000001e (
    .I0(sig000000e3),
    .I1(sig0000006b),
    .O(sig0000009c)
  );
  XORCY   blk0000001f (
    .CI(sig0000009d),
    .LI(sig00000001),
    .O(sig000000cc)
  );
  XORCY   blk00000020 (
    .CI(sig0000009f),
    .LI(sig0000009e),
    .O(sig000000cb)
  );
  MUXCY   blk00000021 (
    .CI(sig0000009f),
    .DI(b[30]),
    .S(sig0000009e),
    .O(sig0000009d)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000022 (
    .I0(b[30]),
    .I1(a[30]),
    .O(sig0000009e)
  );
  XORCY   blk00000023 (
    .CI(sig000000a1),
    .LI(sig000000a0),
    .O(sig000000ca)
  );
  MUXCY   blk00000024 (
    .CI(sig000000a1),
    .DI(b[29]),
    .S(sig000000a0),
    .O(sig0000009f)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000025 (
    .I0(b[29]),
    .I1(a[29]),
    .O(sig000000a0)
  );
  XORCY   blk00000026 (
    .CI(sig000000a3),
    .LI(sig000000a2),
    .O(sig000000c9)
  );
  MUXCY   blk00000027 (
    .CI(sig000000a3),
    .DI(b[28]),
    .S(sig000000a2),
    .O(sig000000a1)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000028 (
    .I0(b[28]),
    .I1(a[28]),
    .O(sig000000a2)
  );
  XORCY   blk00000029 (
    .CI(sig000000a5),
    .LI(sig000000a4),
    .O(sig000000c8)
  );
  MUXCY   blk0000002a (
    .CI(sig000000a5),
    .DI(b[27]),
    .S(sig000000a4),
    .O(sig000000a3)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk0000002b (
    .I0(b[27]),
    .I1(a[27]),
    .O(sig000000a4)
  );
  XORCY   blk0000002c (
    .CI(sig000000a7),
    .LI(sig000000a6),
    .O(sig000000c7)
  );
  MUXCY   blk0000002d (
    .CI(sig000000a7),
    .DI(b[26]),
    .S(sig000000a6),
    .O(sig000000a5)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk0000002e (
    .I0(b[26]),
    .I1(a[26]),
    .O(sig000000a6)
  );
  XORCY   blk0000002f (
    .CI(sig000000a9),
    .LI(sig000000a8),
    .O(sig000000c6)
  );
  MUXCY   blk00000030 (
    .CI(sig000000a9),
    .DI(b[25]),
    .S(sig000000a8),
    .O(sig000000a7)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000031 (
    .I0(b[25]),
    .I1(a[25]),
    .O(sig000000a8)
  );
  XORCY   blk00000032 (
    .CI(sig000000ab),
    .LI(sig000000aa),
    .O(sig000000c5)
  );
  MUXCY   blk00000033 (
    .CI(sig000000ab),
    .DI(b[24]),
    .S(sig000000aa),
    .O(sig000000a9)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000034 (
    .I0(b[24]),
    .I1(a[24]),
    .O(sig000000aa)
  );
  XORCY   blk00000035 (
    .CI(sig00000001),
    .LI(sig000000ac),
    .O(sig000000c4)
  );
  MUXCY   blk00000036 (
    .CI(sig00000001),
    .DI(b[23]),
    .S(sig000000ac),
    .O(sig000000ab)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000037 (
    .I0(b[23]),
    .I1(a[23]),
    .O(sig000000ac)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000038 (
    .C(clk),
    .CE(ce),
    .D(sig000000bf),
    .Q(sig000000df)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000039 (
    .C(clk),
    .CE(ce),
    .D(sig000000e2),
    .Q(sig000000e1)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000003a (
    .C(clk),
    .CE(ce),
    .D(sig000000be),
    .Q(sig000000e0)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000003b (
    .C(clk),
    .CE(ce),
    .D(sig000000ce),
    .Q(sig000000b0)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000003c (
    .C(clk),
    .CE(ce),
    .D(a[31]),
    .Q(sig000000fe)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000003d (
    .C(clk),
    .CE(ce),
    .D(b[31]),
    .Q(sig000000fd)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000003e (
    .C(clk),
    .CE(ce),
    .D(sig0000008b),
    .Q(sig000000b1)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000003f (
    .C(clk),
    .CE(ce),
    .D(sig0000001a),
    .Q(sig000000fc)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000040 (
    .C(clk),
    .CE(ce),
    .D(sig000000c1),
    .Q(sig000000fb)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000041 (
    .C(clk),
    .CE(ce),
    .D(sig000000c3),
    .Q(sig000000fa)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000042 (
    .C(clk),
    .CE(ce),
    .D(sig000000c2),
    .Q(sig000000f8)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000043 (
    .C(clk),
    .CE(ce),
    .D(sig000000c0),
    .Q(sig000001a3)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000044 (
    .C(clk),
    .CE(ce),
    .D(sig000000d1),
    .Q(sig000000f7)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000045 (
    .C(clk),
    .CE(ce),
    .D(sig000000d2),
    .Q(sig000000f9)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000046 (
    .C(clk),
    .CE(ce),
    .D(sig000000d3),
    .Q(sig000000f6)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000047 (
    .C(clk),
    .CE(ce),
    .D(sig000000cd),
    .Q(sig0000001b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000048 (
    .C(clk),
    .CE(ce),
    .D(sig000000b5),
    .Q(sig00000110)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000049 (
    .C(clk),
    .CE(ce),
    .D(sig000000b4),
    .Q(sig00000111)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000004a (
    .C(clk),
    .CE(ce),
    .D(sig000000b3),
    .Q(sig00000113)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000004b (
    .C(clk),
    .CE(ce),
    .D(sig000000b2),
    .Q(sig00000114)
  );
  MUXCY   blk0000004c (
    .CI(sig00000001),
    .DI(sig00000002),
    .S(sig0000011c),
    .O(sig00000116)
  );
  MUXCY   blk0000004d (
    .CI(sig00000116),
    .DI(sig00000002),
    .S(sig0000011b),
    .O(sig00000117)
  );
  MUXCY   blk0000004e (
    .CI(sig00000117),
    .DI(sig00000002),
    .S(sig0000011a),
    .O(sig00000118)
  );
  MUXCY   blk0000004f (
    .CI(sig00000118),
    .DI(sig00000002),
    .S(sig0000011d),
    .O(sig00000119)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000050 (
    .C(clk),
    .CE(ce),
    .D(sig00000119),
    .Q(sig00000115)
  );
  MUXCY   blk00000051 (
    .CI(sig00000001),
    .DI(sig00000002),
    .S(sig00000124),
    .O(sig0000011e)
  );
  MUXCY   blk00000052 (
    .CI(sig0000011e),
    .DI(sig00000002),
    .S(sig00000123),
    .O(sig0000011f)
  );
  MUXCY   blk00000053 (
    .CI(sig0000011f),
    .DI(sig00000002),
    .S(sig00000122),
    .O(sig00000120)
  );
  MUXCY   blk00000054 (
    .CI(sig00000120),
    .DI(sig00000002),
    .S(sig00000125),
    .O(sig00000121)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000055 (
    .C(clk),
    .CE(ce),
    .D(sig00000121),
    .Q(sig00000112)
  );
  MUXCY   blk00000056 (
    .CI(sig00000147),
    .DI(sig00000126),
    .S(sig00000127),
    .O(sig00000146)
  );
  MUXCY   blk00000057 (
    .CI(sig00000148),
    .DI(sig00000128),
    .S(sig00000129),
    .O(sig00000147)
  );
  MUXCY   blk00000058 (
    .CI(sig00000149),
    .DI(sig0000012a),
    .S(sig0000012b),
    .O(sig00000148)
  );
  MUXCY   blk00000059 (
    .CI(sig0000014a),
    .DI(sig0000012c),
    .S(sig0000012d),
    .O(sig00000149)
  );
  MUXCY   blk0000005a (
    .CI(sig0000014b),
    .DI(sig0000012e),
    .S(sig0000012f),
    .O(sig0000014a)
  );
  MUXCY   blk0000005b (
    .CI(sig0000014c),
    .DI(sig00000130),
    .S(sig00000131),
    .O(sig0000014b)
  );
  MUXCY   blk0000005c (
    .CI(sig0000014d),
    .DI(sig00000132),
    .S(sig00000133),
    .O(sig0000014c)
  );
  MUXCY   blk0000005d (
    .CI(sig0000014e),
    .DI(sig00000134),
    .S(sig00000135),
    .O(sig0000014d)
  );
  MUXCY   blk0000005e (
    .CI(sig0000014f),
    .DI(sig00000136),
    .S(sig00000137),
    .O(sig0000014e)
  );
  MUXCY   blk0000005f (
    .CI(sig00000150),
    .DI(sig00000138),
    .S(sig00000139),
    .O(sig0000014f)
  );
  MUXCY   blk00000060 (
    .CI(sig00000151),
    .DI(sig0000013a),
    .S(sig0000013b),
    .O(sig00000150)
  );
  MUXCY   blk00000061 (
    .CI(sig00000152),
    .DI(sig0000013c),
    .S(sig0000013d),
    .O(sig00000151)
  );
  MUXCY   blk00000062 (
    .CI(sig00000153),
    .DI(sig0000013e),
    .S(sig0000013f),
    .O(sig00000152)
  );
  MUXCY   blk00000063 (
    .CI(sig00000154),
    .DI(sig00000140),
    .S(sig00000141),
    .O(sig00000153)
  );
  MUXCY   blk00000064 (
    .CI(sig00000155),
    .DI(sig00000142),
    .S(sig00000143),
    .O(sig00000154)
  );
  MUXCY   blk00000065 (
    .CI(sig00000002),
    .DI(sig00000144),
    .S(sig00000145),
    .O(sig00000155)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000066 (
    .C(clk),
    .CE(ce),
    .D(sig00000146),
    .Q(sig00000019)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000067 (
    .C(clk),
    .CE(ce),
    .D(b[30]),
    .Q(sig00000106)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000068 (
    .C(clk),
    .CE(ce),
    .D(b[29]),
    .Q(sig00000105)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000069 (
    .C(clk),
    .CE(ce),
    .D(b[28]),
    .Q(sig00000104)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000006a (
    .C(clk),
    .CE(ce),
    .D(b[27]),
    .Q(sig00000103)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000006b (
    .C(clk),
    .CE(ce),
    .D(b[26]),
    .Q(sig00000102)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000006c (
    .C(clk),
    .CE(ce),
    .D(b[25]),
    .Q(sig00000101)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000006d (
    .C(clk),
    .CE(ce),
    .D(b[24]),
    .Q(sig00000100)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000006e (
    .C(clk),
    .CE(ce),
    .D(b[23]),
    .Q(sig000000ff)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000006f (
    .C(clk),
    .CE(ce),
    .D(a[30]),
    .Q(sig0000010e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000070 (
    .C(clk),
    .CE(ce),
    .D(a[29]),
    .Q(sig0000010d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000071 (
    .C(clk),
    .CE(ce),
    .D(a[28]),
    .Q(sig0000010c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000072 (
    .C(clk),
    .CE(ce),
    .D(a[27]),
    .Q(sig0000010b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000073 (
    .C(clk),
    .CE(ce),
    .D(a[26]),
    .Q(sig0000010a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000074 (
    .C(clk),
    .CE(ce),
    .D(a[25]),
    .Q(sig00000109)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000075 (
    .C(clk),
    .CE(ce),
    .D(a[24]),
    .Q(sig00000108)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000076 (
    .C(clk),
    .CE(ce),
    .D(a[23]),
    .Q(sig00000107)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000077 (
    .C(clk),
    .CE(ce),
    .D(sig000000cc),
    .Q(sig00000003)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000078 (
    .C(clk),
    .CE(ce),
    .D(sig000000cb),
    .Q(sig00000004)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000079 (
    .C(clk),
    .CE(ce),
    .D(sig000000ca),
    .Q(sig00000005)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000007a (
    .C(clk),
    .CE(ce),
    .D(sig000000c9),
    .Q(sig00000006)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000007b (
    .C(clk),
    .CE(ce),
    .D(sig000000c8),
    .Q(sig00000007)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000007c (
    .C(clk),
    .CE(ce),
    .D(sig000000c7),
    .Q(sig00000008)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000007d (
    .C(clk),
    .CE(ce),
    .D(sig000000c6),
    .Q(sig00000009)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000007e (
    .C(clk),
    .CE(ce),
    .D(sig000000c5),
    .Q(sig0000000a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000007f (
    .C(clk),
    .CE(ce),
    .D(sig000000c4),
    .Q(sig0000000b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000080 (
    .C(clk),
    .CE(ce),
    .D(sig000000d0),
    .Q(sig00000157)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000081 (
    .C(clk),
    .CE(ce),
    .D(sig000000cf),
    .Q(sig00000156)
  );
  XORCY   blk00000082 (
    .CI(sig00000158),
    .LI(sig00000002),
    .O(NLW_blk00000082_O_UNCONNECTED)
  );
  XORCY   blk00000083 (
    .CI(sig00000159),
    .LI(sig000000bd),
    .O(sig000000f2)
  );
  MUXCY   blk00000084 (
    .CI(sig00000159),
    .DI(sig00000002),
    .S(sig000000bd),
    .O(sig00000158)
  );
  XORCY   blk00000085 (
    .CI(sig0000015a),
    .LI(sig000000bc),
    .O(sig000000f1)
  );
  MUXCY   blk00000086 (
    .CI(sig0000015a),
    .DI(sig00000002),
    .S(sig000000bc),
    .O(sig00000159)
  );
  XORCY   blk00000087 (
    .CI(sig0000015b),
    .LI(sig000000bb),
    .O(sig000000f0)
  );
  MUXCY   blk00000088 (
    .CI(sig0000015b),
    .DI(sig00000002),
    .S(sig000000bb),
    .O(sig0000015a)
  );
  XORCY   blk00000089 (
    .CI(sig0000015c),
    .LI(sig000000ba),
    .O(sig000000ef)
  );
  MUXCY   blk0000008a (
    .CI(sig0000015c),
    .DI(sig00000002),
    .S(sig000000ba),
    .O(sig0000015b)
  );
  XORCY   blk0000008b (
    .CI(sig0000015d),
    .LI(sig000000b9),
    .O(sig000000ee)
  );
  MUXCY   blk0000008c (
    .CI(sig0000015d),
    .DI(sig00000002),
    .S(sig000000b9),
    .O(sig0000015c)
  );
  XORCY   blk0000008d (
    .CI(sig0000015e),
    .LI(sig000000b8),
    .O(sig000000ed)
  );
  MUXCY   blk0000008e (
    .CI(sig0000015e),
    .DI(sig00000002),
    .S(sig000000b8),
    .O(sig0000015d)
  );
  XORCY   blk0000008f (
    .CI(sig0000015f),
    .LI(sig000000b7),
    .O(sig000000ec)
  );
  MUXCY   blk00000090 (
    .CI(sig0000015f),
    .DI(sig00000002),
    .S(sig000000b7),
    .O(sig0000015e)
  );
  XORCY   blk00000091 (
    .CI(sig00000002),
    .LI(sig000000b6),
    .O(sig000000eb)
  );
  MUXCY   blk00000092 (
    .CI(sig00000002),
    .DI(sig00000001),
    .S(sig000000b6),
    .O(sig0000015f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000093 (
    .C(clk),
    .CE(ce),
    .D(sig000000dc),
    .Q(sig000000e2)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000094 (
    .C(clk),
    .CE(ce),
    .D(sig000000db),
    .Q(sig00000011)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000095 (
    .C(clk),
    .CE(ce),
    .D(sig000000da),
    .Q(sig00000012)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000096 (
    .C(clk),
    .CE(ce),
    .D(sig000000d9),
    .Q(sig00000013)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000097 (
    .C(clk),
    .CE(ce),
    .D(sig000000d8),
    .Q(sig00000014)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000098 (
    .C(clk),
    .CE(ce),
    .D(sig000000d7),
    .Q(sig00000015)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000099 (
    .C(clk),
    .CE(ce),
    .D(sig000000d6),
    .Q(sig00000016)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000009a (
    .C(clk),
    .CE(ce),
    .D(sig000000d5),
    .Q(sig00000017)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000009b (
    .C(clk),
    .CE(ce),
    .D(sig000000d4),
    .Q(sig00000018)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000009c (
    .C(clk),
    .CE(ce),
    .D(a[22]),
    .Q(sig0000001c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000009d (
    .C(clk),
    .CE(ce),
    .D(a[21]),
    .Q(sig0000001d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000009e (
    .C(clk),
    .CE(ce),
    .D(a[20]),
    .Q(sig0000001e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000009f (
    .C(clk),
    .CE(ce),
    .D(a[19]),
    .Q(sig0000001f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000a0 (
    .C(clk),
    .CE(ce),
    .D(a[18]),
    .Q(sig00000020)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000a1 (
    .C(clk),
    .CE(ce),
    .D(a[17]),
    .Q(sig00000021)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000a2 (
    .C(clk),
    .CE(ce),
    .D(a[16]),
    .Q(sig00000022)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000a3 (
    .C(clk),
    .CE(ce),
    .D(a[15]),
    .Q(sig00000023)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000a4 (
    .C(clk),
    .CE(ce),
    .D(a[14]),
    .Q(sig00000024)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000a5 (
    .C(clk),
    .CE(ce),
    .D(a[13]),
    .Q(sig00000025)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000a6 (
    .C(clk),
    .CE(ce),
    .D(a[12]),
    .Q(sig00000026)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000a7 (
    .C(clk),
    .CE(ce),
    .D(a[11]),
    .Q(sig00000027)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000a8 (
    .C(clk),
    .CE(ce),
    .D(a[10]),
    .Q(sig00000028)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000a9 (
    .C(clk),
    .CE(ce),
    .D(a[9]),
    .Q(sig00000029)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000aa (
    .C(clk),
    .CE(ce),
    .D(a[8]),
    .Q(sig0000002a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000ab (
    .C(clk),
    .CE(ce),
    .D(a[7]),
    .Q(sig0000002b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000ac (
    .C(clk),
    .CE(ce),
    .D(a[6]),
    .Q(sig0000002c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000ad (
    .C(clk),
    .CE(ce),
    .D(a[5]),
    .Q(sig0000002d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000ae (
    .C(clk),
    .CE(ce),
    .D(a[4]),
    .Q(sig0000002e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000af (
    .C(clk),
    .CE(ce),
    .D(a[3]),
    .Q(sig0000002f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000b0 (
    .C(clk),
    .CE(ce),
    .D(a[2]),
    .Q(sig00000030)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000b1 (
    .C(clk),
    .CE(ce),
    .D(a[1]),
    .Q(sig00000031)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000b2 (
    .C(clk),
    .CE(ce),
    .D(a[0]),
    .Q(sig00000032)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000b3 (
    .C(clk),
    .CE(ce),
    .D(b[22]),
    .Q(sig00000033)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000b4 (
    .C(clk),
    .CE(ce),
    .D(b[21]),
    .Q(sig00000034)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000b5 (
    .C(clk),
    .CE(ce),
    .D(b[20]),
    .Q(sig00000035)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000b6 (
    .C(clk),
    .CE(ce),
    .D(b[19]),
    .Q(sig00000036)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000b7 (
    .C(clk),
    .CE(ce),
    .D(b[18]),
    .Q(sig00000037)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000b8 (
    .C(clk),
    .CE(ce),
    .D(b[17]),
    .Q(sig00000038)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000b9 (
    .C(clk),
    .CE(ce),
    .D(b[16]),
    .Q(sig00000039)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000ba (
    .C(clk),
    .CE(ce),
    .D(b[15]),
    .Q(sig0000003a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000bb (
    .C(clk),
    .CE(ce),
    .D(b[14]),
    .Q(sig0000003b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000bc (
    .C(clk),
    .CE(ce),
    .D(b[13]),
    .Q(sig0000003c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000bd (
    .C(clk),
    .CE(ce),
    .D(b[12]),
    .Q(sig0000003d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000be (
    .C(clk),
    .CE(ce),
    .D(b[11]),
    .Q(sig0000003e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000bf (
    .C(clk),
    .CE(ce),
    .D(b[10]),
    .Q(sig0000003f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000c0 (
    .C(clk),
    .CE(ce),
    .D(b[9]),
    .Q(sig00000040)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000c1 (
    .C(clk),
    .CE(ce),
    .D(b[8]),
    .Q(sig00000041)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000c2 (
    .C(clk),
    .CE(ce),
    .D(b[7]),
    .Q(sig00000042)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000c3 (
    .C(clk),
    .CE(ce),
    .D(b[6]),
    .Q(sig00000043)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000c4 (
    .C(clk),
    .CE(ce),
    .D(b[5]),
    .Q(sig00000044)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000c5 (
    .C(clk),
    .CE(ce),
    .D(b[4]),
    .Q(sig00000045)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000c6 (
    .C(clk),
    .CE(ce),
    .D(b[3]),
    .Q(sig00000046)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000c7 (
    .C(clk),
    .CE(ce),
    .D(b[2]),
    .Q(sig00000047)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000c8 (
    .C(clk),
    .CE(ce),
    .D(b[1]),
    .Q(sig00000048)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000c9 (
    .C(clk),
    .CE(ce),
    .D(b[0]),
    .Q(sig00000049)
  );
  MUXCY   blk000000ca (
    .CI(sig000001fa),
    .DI(sig00000001),
    .S(sig000002d6),
    .O(sig000001a2)
  );
  XORCY   blk000000cb (
    .CI(sig000001fa),
    .LI(sig000002d6),
    .O(NLW_blk000000cb_O_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000cc (
    .C(clk),
    .CE(ce),
    .D(sig000001a2),
    .Q(sig000001f9)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000cd (
    .C(clk),
    .CE(ce),
    .D(sig000001a3),
    .Q(sig000001fb)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000ce (
    .C(clk),
    .CE(ce),
    .D(sig000001c0),
    .Q(sig000001a4)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000cf (
    .C(clk),
    .CE(ce),
    .D(sig000001a4),
    .Q(sig000001a1)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000d0 (
    .C(clk),
    .CE(ce),
    .D(sig000001fc),
    .Q(sig000001a5)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000d1 (
    .C(clk),
    .CE(ce),
    .D(sig000001a5),
    .Q(sig000001a0)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000d2 (
    .C(clk),
    .CE(ce),
    .D(sig000001bf),
    .Q(sig000001f8)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000d3 (
    .C(clk),
    .CE(ce),
    .D(sig000001be),
    .Q(sig00000065)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000d4 (
    .C(clk),
    .CE(ce),
    .D(sig00000214),
    .Q(sig00000188)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000d5 (
    .C(clk),
    .CE(ce),
    .D(sig00000213),
    .Q(sig00000189)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000d6 (
    .C(clk),
    .CE(ce),
    .D(sig00000212),
    .Q(sig0000018a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000d7 (
    .C(clk),
    .CE(ce),
    .D(sig00000211),
    .Q(sig0000018b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000d8 (
    .C(clk),
    .CE(ce),
    .D(sig00000210),
    .Q(sig0000018c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000d9 (
    .C(clk),
    .CE(ce),
    .D(sig0000020f),
    .Q(sig0000018d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000da (
    .C(clk),
    .CE(ce),
    .D(sig0000020e),
    .Q(sig0000018e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000db (
    .C(clk),
    .CE(ce),
    .D(sig0000020d),
    .Q(sig0000018f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000dc (
    .C(clk),
    .CE(ce),
    .D(sig0000020c),
    .Q(sig00000190)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000dd (
    .C(clk),
    .CE(ce),
    .D(sig0000020b),
    .Q(sig00000191)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000de (
    .C(clk),
    .CE(ce),
    .D(sig0000020a),
    .Q(sig00000192)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000df (
    .C(clk),
    .CE(ce),
    .D(sig00000209),
    .Q(sig00000193)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000e0 (
    .C(clk),
    .CE(ce),
    .D(sig00000208),
    .Q(sig00000194)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000e1 (
    .C(clk),
    .CE(ce),
    .D(sig00000207),
    .Q(sig00000195)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000e2 (
    .C(clk),
    .CE(ce),
    .D(sig00000206),
    .Q(sig00000196)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000e3 (
    .C(clk),
    .CE(ce),
    .D(sig00000205),
    .Q(sig00000197)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000e4 (
    .C(clk),
    .CE(ce),
    .D(sig00000204),
    .Q(sig00000198)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000e5 (
    .C(clk),
    .CE(ce),
    .D(sig00000203),
    .Q(sig00000199)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000e6 (
    .C(clk),
    .CE(ce),
    .D(sig00000202),
    .Q(sig0000019a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000e7 (
    .C(clk),
    .CE(ce),
    .D(sig00000201),
    .Q(sig0000019b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000e8 (
    .C(clk),
    .CE(ce),
    .D(sig00000200),
    .Q(sig0000019c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000e9 (
    .C(clk),
    .CE(ce),
    .D(sig000001ff),
    .Q(sig0000019d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000ea (
    .C(clk),
    .CE(ce),
    .D(sig000001fe),
    .Q(sig0000019e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000eb (
    .C(clk),
    .CE(ce),
    .D(sig000001fd),
    .Q(sig0000019f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000ec (
    .C(clk),
    .CE(ce),
    .D(sig00000001),
    .Q(sig00000214)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000ed (
    .C(clk),
    .CE(ce),
    .D(sig000001e9),
    .Q(sig00000213)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000ee (
    .C(clk),
    .CE(ce),
    .D(sig000001e8),
    .Q(sig00000212)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000ef (
    .C(clk),
    .CE(ce),
    .D(sig000001e7),
    .Q(sig00000211)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000f0 (
    .C(clk),
    .CE(ce),
    .D(sig000001e6),
    .Q(sig00000210)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000f1 (
    .C(clk),
    .CE(ce),
    .D(sig000001e5),
    .Q(sig0000020f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000f2 (
    .C(clk),
    .CE(ce),
    .D(sig000001e4),
    .Q(sig0000020e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000f3 (
    .C(clk),
    .CE(ce),
    .D(sig000001e3),
    .Q(sig0000020d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000f4 (
    .C(clk),
    .CE(ce),
    .D(sig000001e2),
    .Q(sig0000020c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000f5 (
    .C(clk),
    .CE(ce),
    .D(sig000001e1),
    .Q(sig0000020b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000f6 (
    .C(clk),
    .CE(ce),
    .D(sig000001e0),
    .Q(sig0000020a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000f7 (
    .C(clk),
    .CE(ce),
    .D(sig000001df),
    .Q(sig00000209)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000f8 (
    .C(clk),
    .CE(ce),
    .D(sig000001de),
    .Q(sig00000208)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000f9 (
    .C(clk),
    .CE(ce),
    .D(sig000001dd),
    .Q(sig00000207)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000fa (
    .C(clk),
    .CE(ce),
    .D(sig000001dc),
    .Q(sig00000206)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000fb (
    .C(clk),
    .CE(ce),
    .D(sig000001db),
    .Q(sig00000205)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000fc (
    .C(clk),
    .CE(ce),
    .D(sig000001da),
    .Q(sig00000204)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000fd (
    .C(clk),
    .CE(ce),
    .D(sig000001d9),
    .Q(sig00000203)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000fe (
    .C(clk),
    .CE(ce),
    .D(sig000001d8),
    .Q(sig00000202)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000000ff (
    .C(clk),
    .CE(ce),
    .D(sig000001d7),
    .Q(sig00000201)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000100 (
    .C(clk),
    .CE(ce),
    .D(sig000001d6),
    .Q(sig00000200)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000101 (
    .C(clk),
    .CE(ce),
    .D(sig000001d5),
    .Q(sig000001ff)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000102 (
    .C(clk),
    .CE(ce),
    .D(sig000001d4),
    .Q(sig000001fe)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000103 (
    .C(clk),
    .CE(ce),
    .D(sig000001d3),
    .Q(sig000001fd)
  );
  MUXCY   blk00000104 (
    .CI(sig00000001),
    .DI(sig00000002),
    .S(sig00000221),
    .O(sig00000215)
  );
  MUXCY   blk00000105 (
    .CI(sig00000215),
    .DI(sig00000002),
    .S(sig00000220),
    .O(sig00000216)
  );
  MUXCY   blk00000106 (
    .CI(sig00000216),
    .DI(sig00000002),
    .S(sig0000021f),
    .O(sig00000217)
  );
  MUXCY   blk00000107 (
    .CI(sig00000217),
    .DI(sig00000002),
    .S(sig0000021e),
    .O(sig00000218)
  );
  MUXCY   blk00000108 (
    .CI(sig00000218),
    .DI(sig00000002),
    .S(sig0000021d),
    .O(sig00000219)
  );
  MUXCY   blk00000109 (
    .CI(sig00000219),
    .DI(sig00000002),
    .S(sig0000021c),
    .O(sig0000021a)
  );
  MUXCY   blk0000010a (
    .CI(sig0000021a),
    .DI(sig00000002),
    .S(sig0000021b),
    .O(sig000001fa)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000010b (
    .C(clk),
    .CE(ce),
    .D(sig000001d0),
    .Q(sig00000178)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000010c (
    .C(clk),
    .CE(ce),
    .D(sig000001cf),
    .Q(sig00000179)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000010d (
    .C(clk),
    .CE(ce),
    .D(sig000001ce),
    .Q(sig0000017a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000010e (
    .C(clk),
    .CE(ce),
    .D(sig000001cd),
    .Q(sig0000017b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000010f (
    .C(clk),
    .CE(ce),
    .D(sig000001cc),
    .Q(sig0000017c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000110 (
    .C(clk),
    .CE(ce),
    .D(sig000001cb),
    .Q(sig0000017d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000111 (
    .C(clk),
    .CE(ce),
    .D(sig000001ca),
    .Q(sig0000017e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000112 (
    .C(clk),
    .CE(ce),
    .D(sig000001c9),
    .Q(sig0000017f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000113 (
    .C(clk),
    .CE(ce),
    .D(sig000001c8),
    .Q(sig00000180)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000114 (
    .C(clk),
    .CE(ce),
    .D(sig000001c7),
    .Q(sig00000181)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000115 (
    .C(clk),
    .CE(ce),
    .D(sig000001c6),
    .Q(sig00000182)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000116 (
    .C(clk),
    .CE(ce),
    .D(sig000001c5),
    .Q(sig00000183)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000117 (
    .C(clk),
    .CE(ce),
    .D(sig000001c4),
    .Q(sig00000184)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000118 (
    .C(clk),
    .CE(ce),
    .D(sig000001c3),
    .Q(sig00000185)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000119 (
    .C(clk),
    .CE(ce),
    .D(sig000001c2),
    .Q(sig00000186)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000011a (
    .C(clk),
    .CE(ce),
    .D(sig000001c1),
    .Q(sig00000187)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000011b (
    .C(clk),
    .CE(ce),
    .D(sig000001bd),
    .Q(sig00000160)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000011c (
    .C(clk),
    .CE(ce),
    .D(sig000001bc),
    .Q(sig00000161)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000011d (
    .C(clk),
    .CE(ce),
    .D(sig000001bb),
    .Q(sig00000162)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000011e (
    .C(clk),
    .CE(ce),
    .D(sig000001ba),
    .Q(sig00000163)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000011f (
    .C(clk),
    .CE(ce),
    .D(sig000001b9),
    .Q(sig00000164)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000120 (
    .C(clk),
    .CE(ce),
    .D(sig000001b8),
    .Q(sig00000165)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000121 (
    .C(clk),
    .CE(ce),
    .D(sig000001b7),
    .Q(sig00000166)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000122 (
    .C(clk),
    .CE(ce),
    .D(sig000001b6),
    .Q(sig00000167)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000123 (
    .C(clk),
    .CE(ce),
    .D(sig000001b5),
    .Q(sig00000168)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000124 (
    .C(clk),
    .CE(ce),
    .D(sig000001b4),
    .Q(sig00000169)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000125 (
    .C(clk),
    .CE(ce),
    .D(sig000001b3),
    .Q(sig0000016a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000126 (
    .C(clk),
    .CE(ce),
    .D(sig000001b2),
    .Q(sig0000016b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000127 (
    .C(clk),
    .CE(ce),
    .D(sig000001b1),
    .Q(sig0000016c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000128 (
    .C(clk),
    .CE(ce),
    .D(sig000001b0),
    .Q(sig0000016d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000129 (
    .C(clk),
    .CE(ce),
    .D(sig000001af),
    .Q(sig0000016e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000012a (
    .C(clk),
    .CE(ce),
    .D(sig000001ae),
    .Q(sig0000016f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000012b (
    .C(clk),
    .CE(ce),
    .D(sig000001ad),
    .Q(sig00000170)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000012c (
    .C(clk),
    .CE(ce),
    .D(sig000001ac),
    .Q(sig00000171)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000012d (
    .C(clk),
    .CE(ce),
    .D(sig000001ab),
    .Q(sig00000172)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000012e (
    .C(clk),
    .CE(ce),
    .D(sig000001aa),
    .Q(sig00000173)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000012f (
    .C(clk),
    .CE(ce),
    .D(sig000001a9),
    .Q(sig00000174)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000130 (
    .C(clk),
    .CE(ce),
    .D(sig000001a8),
    .Q(sig00000175)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000131 (
    .C(clk),
    .CE(ce),
    .D(sig000001a7),
    .Q(sig00000176)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000132 (
    .C(clk),
    .CE(ce),
    .D(sig000001a6),
    .Q(sig00000177)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000133 (
    .C(clk),
    .CE(ce),
    .D(sig00000229),
    .Q(sig00000222)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000134 (
    .C(clk),
    .CE(ce),
    .D(sig00000222),
    .Q(sig0000022a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000135 (
    .C(clk),
    .CE(ce),
    .D(sig00000228),
    .Q(sig00000223)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000136 (
    .C(clk),
    .CE(ce),
    .D(sig00000223),
    .Q(sig0000022e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000137 (
    .C(clk),
    .CE(ce),
    .D(sig00000227),
    .Q(sig00000224)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000138 (
    .C(clk),
    .CE(ce),
    .D(sig00000224),
    .Q(sig0000022d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000139 (
    .C(clk),
    .CE(ce),
    .D(sig00000226),
    .Q(sig00000230)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000013a (
    .C(clk),
    .CE(ce),
    .D(sig00000231),
    .Q(sig0000022f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000013b (
    .C(clk),
    .CE(ce),
    .D(sig00000225),
    .Q(sig0000022c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000013c (
    .C(clk),
    .CE(ce),
    .D(sig00000285),
    .Q(sig0000024c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000013d (
    .C(clk),
    .CE(ce),
    .D(sig00000282),
    .Q(sig0000024d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000013e (
    .C(clk),
    .CE(ce),
    .D(sig00000281),
    .Q(sig0000024e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000013f (
    .C(clk),
    .CE(ce),
    .D(sig00000280),
    .Q(sig0000024f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000140 (
    .C(clk),
    .CE(ce),
    .D(sig0000027f),
    .Q(sig00000250)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000141 (
    .C(clk),
    .CE(ce),
    .D(sig0000027c),
    .Q(sig00000251)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000142 (
    .C(clk),
    .CE(ce),
    .D(sig0000027b),
    .Q(sig00000252)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000143 (
    .C(clk),
    .CE(ce),
    .D(sig0000027a),
    .Q(sig00000253)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000144 (
    .C(clk),
    .CE(ce),
    .D(sig00000279),
    .Q(sig00000254)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000145 (
    .C(clk),
    .CE(ce),
    .D(sig00000276),
    .Q(sig00000255)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000146 (
    .C(clk),
    .CE(ce),
    .D(sig00000275),
    .Q(sig00000256)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000147 (
    .C(clk),
    .CE(ce),
    .D(sig00000274),
    .Q(sig00000257)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000148 (
    .C(clk),
    .CE(ce),
    .D(sig00000273),
    .Q(sig00000258)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000149 (
    .C(clk),
    .CE(ce),
    .D(sig00000270),
    .Q(sig00000259)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000014a (
    .C(clk),
    .CE(ce),
    .D(sig0000026f),
    .Q(sig0000025a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000014b (
    .C(clk),
    .CE(ce),
    .D(sig0000026e),
    .Q(sig0000025b)
  );
  MUXCY   blk0000014c (
    .CI(sig0000025d),
    .DI(sig00000002),
    .S(sig00000264),
    .O(sig0000025c)
  );
  MUXCY   blk0000014d (
    .CI(sig0000025e),
    .DI(sig00000002),
    .S(sig00000265),
    .O(sig0000025d)
  );
  MUXCY   blk0000014e (
    .CI(sig0000025f),
    .DI(sig00000002),
    .S(sig00000266),
    .O(sig0000025e)
  );
  MUXCY   blk0000014f (
    .CI(sig00000260),
    .DI(sig00000002),
    .S(sig00000267),
    .O(sig0000025f)
  );
  MUXCY   blk00000150 (
    .CI(sig00000261),
    .DI(sig00000002),
    .S(sig00000268),
    .O(sig00000260)
  );
  MUXCY   blk00000151 (
    .CI(sig00000262),
    .DI(sig00000002),
    .S(sig00000269),
    .O(sig00000261)
  );
  MUXCY   blk00000152 (
    .CI(sig00000263),
    .DI(sig00000002),
    .S(sig0000026a),
    .O(sig00000262)
  );
  MUXCY   blk00000153 (
    .CI(sig00000001),
    .DI(sig00000002),
    .S(sig0000026b),
    .O(sig00000263)
  );
  LUT5 #(
    .INIT ( 32'h000000FC ))
  blk00000154 (
    .I0(sig00000002),
    .I1(sig0000023c),
    .I2(sig0000023d),
    .I3(sig0000023e),
    .I4(sig0000023f),
    .O(sig00000271)
  );
  LUT5 #(
    .INIT ( 32'h0000FF0C ))
  blk00000155 (
    .I0(sig00000002),
    .I1(sig0000023c),
    .I2(sig0000023d),
    .I3(sig0000023e),
    .I4(sig0000023f),
    .O(sig00000272)
  );
  LUT5 #(
    .INIT ( 32'h000000FC ))
  blk00000156 (
    .I0(sig00000002),
    .I1(sig00000240),
    .I2(sig00000241),
    .I3(sig00000242),
    .I4(sig00000243),
    .O(sig00000277)
  );
  LUT5 #(
    .INIT ( 32'h0000FF0C ))
  blk00000157 (
    .I0(sig00000002),
    .I1(sig00000240),
    .I2(sig00000241),
    .I3(sig00000242),
    .I4(sig00000243),
    .O(sig00000278)
  );
  LUT5 #(
    .INIT ( 32'h000000FC ))
  blk00000158 (
    .I0(sig00000002),
    .I1(sig00000244),
    .I2(sig00000245),
    .I3(sig00000246),
    .I4(sig00000247),
    .O(sig0000027d)
  );
  LUT5 #(
    .INIT ( 32'h0000FF0C ))
  blk00000159 (
    .I0(sig00000002),
    .I1(sig00000244),
    .I2(sig00000245),
    .I3(sig00000246),
    .I4(sig00000247),
    .O(sig0000027e)
  );
  LUT5 #(
    .INIT ( 32'h000000FC ))
  blk0000015a (
    .I0(sig00000002),
    .I1(sig00000248),
    .I2(sig00000249),
    .I3(sig0000024b),
    .I4(sig0000024a),
    .O(sig00000283)
  );
  LUT5 #(
    .INIT ( 32'h0000FF0C ))
  blk0000015b (
    .I0(sig00000002),
    .I1(sig00000248),
    .I2(sig00000249),
    .I3(sig0000024b),
    .I4(sig0000024a),
    .O(sig00000284)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000015c (
    .C(clk),
    .CE(ce),
    .D(sig0000026d),
    .Q(sig0000006b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000015d (
    .C(clk),
    .CE(ce),
    .D(sig0000026c),
    .Q(sig0000006a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000015e (
    .C(clk),
    .CE(ce),
    .D(sig00000286),
    .Q(sig00000069)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000015f (
    .C(clk),
    .CE(ce),
    .D(sig0000028b),
    .Q(sig00000068)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000160 (
    .C(clk),
    .CE(ce),
    .D(sig0000028f),
    .Q(sig00000067)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000161 (
    .C(clk),
    .CE(ce),
    .D(sig00000066),
    .Q(sig0000028f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000162 (
    .C(clk),
    .CE(ce),
    .D(sig0000025c),
    .Q(sig00000287)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000163 (
    .C(clk),
    .CE(ce),
    .D(sig0000025d),
    .Q(sig00000288)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000164 (
    .C(clk),
    .CE(ce),
    .D(sig0000025e),
    .Q(sig00000289)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000165 (
    .C(clk),
    .CE(ce),
    .D(sig0000025f),
    .Q(sig0000028a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000166 (
    .C(clk),
    .CE(ce),
    .D(sig00000260),
    .Q(sig0000028b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000167 (
    .C(clk),
    .CE(ce),
    .D(sig00000261),
    .Q(sig0000028c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000168 (
    .C(clk),
    .CE(ce),
    .D(sig00000262),
    .Q(sig0000028d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000169 (
    .C(clk),
    .CE(ce),
    .D(sig00000263),
    .Q(sig0000028e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000016a (
    .C(clk),
    .CE(ce),
    .D(sig000002a9),
    .Q(sig0000024a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000016b (
    .C(clk),
    .CE(ce),
    .D(sig000002a8),
    .Q(sig0000024b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000016c (
    .C(clk),
    .CE(ce),
    .D(sig000002a7),
    .Q(sig00000249)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000016d (
    .C(clk),
    .CE(ce),
    .D(sig000002a6),
    .Q(sig00000248)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000016e (
    .C(clk),
    .CE(ce),
    .D(sig000002a5),
    .Q(sig00000247)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000016f (
    .C(clk),
    .CE(ce),
    .D(sig000002a4),
    .Q(sig00000246)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000170 (
    .C(clk),
    .CE(ce),
    .D(sig000002a3),
    .Q(sig00000245)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000171 (
    .C(clk),
    .CE(ce),
    .D(sig000002a2),
    .Q(sig00000244)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000172 (
    .C(clk),
    .CE(ce),
    .D(sig000002a1),
    .Q(sig00000243)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000173 (
    .C(clk),
    .CE(ce),
    .D(sig000002a0),
    .Q(sig00000242)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000174 (
    .C(clk),
    .CE(ce),
    .D(sig0000029f),
    .Q(sig00000241)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000175 (
    .C(clk),
    .CE(ce),
    .D(sig0000029e),
    .Q(sig00000240)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000176 (
    .C(clk),
    .CE(ce),
    .D(sig0000029d),
    .Q(sig0000023f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000177 (
    .C(clk),
    .CE(ce),
    .D(sig0000029c),
    .Q(sig0000023e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000178 (
    .C(clk),
    .CE(ce),
    .D(sig0000029b),
    .Q(sig0000023d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000179 (
    .C(clk),
    .CE(ce),
    .D(sig0000029a),
    .Q(sig0000023c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000017a (
    .C(clk),
    .CE(ce),
    .D(sig00000299),
    .Q(sig0000023b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000017b (
    .C(clk),
    .CE(ce),
    .D(sig00000298),
    .Q(sig0000023a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000017c (
    .C(clk),
    .CE(ce),
    .D(sig00000297),
    .Q(sig00000239)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000017d (
    .C(clk),
    .CE(ce),
    .D(sig00000296),
    .Q(sig00000238)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000017e (
    .C(clk),
    .CE(ce),
    .D(sig00000295),
    .Q(sig00000237)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000017f (
    .C(clk),
    .CE(ce),
    .D(sig00000294),
    .Q(sig00000236)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000180 (
    .C(clk),
    .CE(ce),
    .D(sig00000293),
    .Q(sig00000235)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000181 (
    .C(clk),
    .CE(ce),
    .D(sig00000292),
    .Q(sig00000234)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000182 (
    .C(clk),
    .CE(ce),
    .D(sig00000291),
    .Q(sig00000233)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000183 (
    .C(clk),
    .CE(ce),
    .D(sig00000290),
    .Q(sig00000232)
  );
  FD   blk00000184 (
    .C(clk),
    .D(sig000002c0),
    .Q(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.DSP.OP/OP/mant_op [22])
  );
  FD   blk00000185 (
    .C(clk),
    .D(sig000002bf),
    .Q(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.DSP.OP/OP/mant_op [21])
  );
  FD   blk00000186 (
    .C(clk),
    .D(sig000002be),
    .Q(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.DSP.OP/OP/mant_op [20])
  );
  FD   blk00000187 (
    .C(clk),
    .D(sig000002bd),
    .Q(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.DSP.OP/OP/mant_op [19])
  );
  FD   blk00000188 (
    .C(clk),
    .D(sig000002bc),
    .Q(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.DSP.OP/OP/mant_op [18])
  );
  FD   blk00000189 (
    .C(clk),
    .D(sig000002bb),
    .Q(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.DSP.OP/OP/mant_op [17])
  );
  FD   blk0000018a (
    .C(clk),
    .D(sig000002ba),
    .Q(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.DSP.OP/OP/mant_op [16])
  );
  FD   blk0000018b (
    .C(clk),
    .D(sig000002b9),
    .Q(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.DSP.OP/OP/mant_op [15])
  );
  FD   blk0000018c (
    .C(clk),
    .D(sig000002b8),
    .Q(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.DSP.OP/OP/mant_op [14])
  );
  FD   blk0000018d (
    .C(clk),
    .D(sig000002b7),
    .Q(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.DSP.OP/OP/mant_op [13])
  );
  FD   blk0000018e (
    .C(clk),
    .D(sig000002b6),
    .Q(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.DSP.OP/OP/mant_op [12])
  );
  FD   blk0000018f (
    .C(clk),
    .D(sig000002b5),
    .Q(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.DSP.OP/OP/mant_op [11])
  );
  FD   blk00000190 (
    .C(clk),
    .D(sig000002b4),
    .Q(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.DSP.OP/OP/mant_op [10])
  );
  FD   blk00000191 (
    .C(clk),
    .D(sig000002b3),
    .Q(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.DSP.OP/OP/mant_op [9])
  );
  FD   blk00000192 (
    .C(clk),
    .D(sig000002b2),
    .Q(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.DSP.OP/OP/mant_op [8])
  );
  FD   blk00000193 (
    .C(clk),
    .D(sig000002b1),
    .Q(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.DSP.OP/OP/mant_op [7])
  );
  FD   blk00000194 (
    .C(clk),
    .D(sig000002b0),
    .Q(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.DSP.OP/OP/mant_op [6])
  );
  FD   blk00000195 (
    .C(clk),
    .D(sig000002af),
    .Q(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.DSP.OP/OP/mant_op [5])
  );
  FD   blk00000196 (
    .C(clk),
    .D(sig000002ae),
    .Q(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.DSP.OP/OP/mant_op [4])
  );
  FD   blk00000197 (
    .C(clk),
    .D(sig000002ad),
    .Q(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.DSP.OP/OP/mant_op [3])
  );
  FD   blk00000198 (
    .C(clk),
    .D(sig000002ac),
    .Q(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.DSP.OP/OP/mant_op [2])
  );
  FD   blk00000199 (
    .C(clk),
    .D(sig000002ab),
    .Q(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.DSP.OP/OP/mant_op [1])
  );
  FD   blk0000019a (
    .C(clk),
    .D(sig000002aa),
    .Q(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.DSP.OP/OP/mant_op [0])
  );
  LUT4 #(
    .INIT ( 16'hAA8A ))
  blk0000019b (
    .I0(sig000000f3),
    .I1(sig000000f5),
    .I2(sig0000010f),
    .I3(sig000000f4),
    .O(sig000000cd)
  );
  LUT4 #(
    .INIT ( 16'hEA2A ))
  blk0000019c (
    .I0(sig000000fd),
    .I1(sig00000114),
    .I2(sig00000115),
    .I3(sig000000fe),
    .O(sig000000d1)
  );
  LUT4 #(
    .INIT ( 16'hF888 ))
  blk0000019d (
    .I0(sig00000111),
    .I1(sig00000112),
    .I2(sig00000114),
    .I3(sig00000115),
    .O(sig000000c2)
  );
  LUT4 #(
    .INIT ( 16'h8000 ))
  blk0000019e (
    .I0(sig00000111),
    .I1(sig00000112),
    .I2(sig00000114),
    .I3(sig00000115),
    .O(sig000000c3)
  );
  LUT6 #(
    .INIT ( 64'hFFFFFFFFFFFFFFFE ))
  blk0000019f (
    .I0(sig0000010f),
    .I1(sig000000df),
    .I2(sig000000e1),
    .I3(sig000000e0),
    .I4(sig000000f4),
    .I5(sig000000f5),
    .O(sig000000ad)
  );
  LUT5 #(
    .INIT ( 32'h55555554 ))
  blk000001a0 (
    .I0(sig000000f4),
    .I1(sig0000010f),
    .I2(sig000000f5),
    .I3(sig000000e1),
    .I4(sig000000e0),
    .O(sig000000af)
  );
  LUT5 #(
    .INIT ( 32'hFFFF1504 ))
  blk000001a1 (
    .I0(sig000000fb),
    .I1(sig000000fa),
    .I2(sig000001a3),
    .I3(sig000000f8),
    .I4(sig000000fc),
    .O(sig000000d0)
  );
  LUT4 #(
    .INIT ( 16'h5554 ))
  blk000001a2 (
    .I0(sig000000fc),
    .I1(sig000000fa),
    .I2(sig000000f8),
    .I3(sig000000fb),
    .O(sig000000cf)
  );
  LUT6 #(
    .INIT ( 64'hFFFFFFFF55555554 ))
  blk000001a3 (
    .I0(sig000000f4),
    .I1(sig0000010f),
    .I2(sig000000df),
    .I3(sig000000e1),
    .I4(sig000000e0),
    .I5(sig000000f5),
    .O(sig000000de)
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  blk000001a4 (
    .I0(sig000000f5),
    .I1(sig000000f4),
    .O(sig000000ae)
  );
  LUT6 #(
    .INIT ( 64'hAAAAAAAAAAAAABAA ))
  blk000001a5 (
    .I0(sig000000f4),
    .I1(sig0000010f),
    .I2(sig000000f5),
    .I3(sig000000df),
    .I4(sig000000e1),
    .I5(sig000000e0),
    .O(sig000000dd)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk000001a6 (
    .I0(sig00000003),
    .I1(sig00000108),
    .I2(sig00000100),
    .O(sig000000b7)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk000001a7 (
    .I0(sig00000003),
    .I1(sig00000109),
    .I2(sig00000101),
    .O(sig000000b8)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk000001a8 (
    .I0(sig00000003),
    .I1(sig0000010a),
    .I2(sig00000102),
    .O(sig000000b9)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk000001a9 (
    .I0(sig00000003),
    .I1(sig0000010b),
    .I2(sig00000103),
    .O(sig000000ba)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk000001aa (
    .I0(sig00000003),
    .I1(sig0000010c),
    .I2(sig00000104),
    .O(sig000000bb)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk000001ab (
    .I0(sig00000003),
    .I1(sig0000010d),
    .I2(sig00000105),
    .O(sig000000bc)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk000001ac (
    .I0(sig00000003),
    .I1(sig0000010e),
    .I2(sig00000106),
    .O(sig000000bd)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk000001ad (
    .I0(sig00000019),
    .I1(sig000000fd),
    .I2(sig000000fe),
    .O(sig000000d3)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk000001ae (
    .I0(sig000000fe),
    .I1(sig000000fd),
    .O(sig000000c0)
  );
  LUT3 #(
    .INIT ( 8'h1B ))
  blk000001af (
    .I0(sig00000003),
    .I1(sig000000ff),
    .I2(sig00000107),
    .O(sig000000b6)
  );
  LUT4 #(
    .INIT ( 16'h22F2 ))
  blk000001b0 (
    .I0(sig00000114),
    .I1(sig00000115),
    .I2(sig00000111),
    .I3(sig00000112),
    .O(sig000000c1)
  );
  LUT2 #(
    .INIT ( 4'h8 ))
  blk000001b1 (
    .I0(sig000000fe),
    .I1(sig000000fd),
    .O(sig000000d2)
  );
  LUT2 #(
    .INIT ( 4'h8 ))
  blk000001b2 (
    .I0(sig00000110),
    .I1(sig00000113),
    .O(sig0000001a)
  );
  LUT6 #(
    .INIT ( 64'h0000000000000001 ))
  blk000001b3 (
    .I0(a[12]),
    .I1(a[13]),
    .I2(a[14]),
    .I3(a[15]),
    .I4(a[16]),
    .I5(a[17]),
    .O(sig0000011a)
  );
  LUT6 #(
    .INIT ( 64'h0000000000000001 ))
  blk000001b4 (
    .I0(a[6]),
    .I1(a[7]),
    .I2(a[8]),
    .I3(a[9]),
    .I4(a[10]),
    .I5(a[11]),
    .O(sig0000011b)
  );
  LUT6 #(
    .INIT ( 64'h0000000000000001 ))
  blk000001b5 (
    .I0(a[0]),
    .I1(a[1]),
    .I2(a[2]),
    .I3(a[3]),
    .I4(a[4]),
    .I5(a[5]),
    .O(sig0000011c)
  );
  LUT5 #(
    .INIT ( 32'h00000001 ))
  blk000001b6 (
    .I0(a[18]),
    .I1(a[19]),
    .I2(a[20]),
    .I3(a[21]),
    .I4(a[22]),
    .O(sig0000011d)
  );
  LUT6 #(
    .INIT ( 64'h0000000000000001 ))
  blk000001b7 (
    .I0(b[12]),
    .I1(b[13]),
    .I2(b[14]),
    .I3(b[15]),
    .I4(b[16]),
    .I5(b[17]),
    .O(sig00000122)
  );
  LUT6 #(
    .INIT ( 64'h0000000000000001 ))
  blk000001b8 (
    .I0(b[6]),
    .I1(b[7]),
    .I2(b[8]),
    .I3(b[9]),
    .I4(b[10]),
    .I5(b[11]),
    .O(sig00000123)
  );
  LUT6 #(
    .INIT ( 64'h0000000000000001 ))
  blk000001b9 (
    .I0(b[0]),
    .I1(b[1]),
    .I2(b[2]),
    .I3(b[3]),
    .I4(b[4]),
    .I5(b[5]),
    .O(sig00000124)
  );
  LUT5 #(
    .INIT ( 32'h00000001 ))
  blk000001ba (
    .I0(b[18]),
    .I1(b[19]),
    .I2(b[20]),
    .I3(b[21]),
    .I4(b[22]),
    .O(sig00000125)
  );
  LUT4 #(
    .INIT ( 16'h9009 ))
  blk000001bb (
    .I0(b[19]),
    .I1(a[19]),
    .I2(b[18]),
    .I3(a[18]),
    .O(sig00000133)
  );
  LUT4 #(
    .INIT ( 16'h9009 ))
  blk000001bc (
    .I0(b[17]),
    .I1(a[17]),
    .I2(b[16]),
    .I3(a[16]),
    .O(sig00000135)
  );
  LUT4 #(
    .INIT ( 16'h9009 ))
  blk000001bd (
    .I0(b[15]),
    .I1(a[15]),
    .I2(b[14]),
    .I3(a[14]),
    .O(sig00000137)
  );
  LUT4 #(
    .INIT ( 16'h9009 ))
  blk000001be (
    .I0(b[13]),
    .I1(a[13]),
    .I2(b[12]),
    .I3(a[12]),
    .O(sig00000139)
  );
  LUT4 #(
    .INIT ( 16'h9009 ))
  blk000001bf (
    .I0(b[11]),
    .I1(a[11]),
    .I2(b[10]),
    .I3(a[10]),
    .O(sig0000013b)
  );
  LUT4 #(
    .INIT ( 16'h9009 ))
  blk000001c0 (
    .I0(b[9]),
    .I1(a[9]),
    .I2(b[8]),
    .I3(a[8]),
    .O(sig0000013d)
  );
  LUT4 #(
    .INIT ( 16'h9009 ))
  blk000001c1 (
    .I0(b[7]),
    .I1(a[7]),
    .I2(b[6]),
    .I3(a[6]),
    .O(sig0000013f)
  );
  LUT4 #(
    .INIT ( 16'h9009 ))
  blk000001c2 (
    .I0(b[5]),
    .I1(a[5]),
    .I2(b[4]),
    .I3(a[4]),
    .O(sig00000141)
  );
  LUT4 #(
    .INIT ( 16'h9009 ))
  blk000001c3 (
    .I0(b[3]),
    .I1(a[3]),
    .I2(b[2]),
    .I3(a[2]),
    .O(sig00000143)
  );
  LUT4 #(
    .INIT ( 16'h9009 ))
  blk000001c4 (
    .I0(b[29]),
    .I1(a[29]),
    .I2(b[28]),
    .I3(a[28]),
    .O(sig00000129)
  );
  LUT4 #(
    .INIT ( 16'h9009 ))
  blk000001c5 (
    .I0(b[27]),
    .I1(a[27]),
    .I2(b[26]),
    .I3(a[26]),
    .O(sig0000012b)
  );
  LUT4 #(
    .INIT ( 16'h9009 ))
  blk000001c6 (
    .I0(b[25]),
    .I1(a[25]),
    .I2(b[24]),
    .I3(a[24]),
    .O(sig0000012d)
  );
  LUT4 #(
    .INIT ( 16'h9009 ))
  blk000001c7 (
    .I0(b[23]),
    .I1(a[23]),
    .I2(b[22]),
    .I3(a[22]),
    .O(sig0000012f)
  );
  LUT4 #(
    .INIT ( 16'h9009 ))
  blk000001c8 (
    .I0(b[21]),
    .I1(a[21]),
    .I2(b[20]),
    .I3(a[20]),
    .O(sig00000131)
  );
  LUT4 #(
    .INIT ( 16'h9009 ))
  blk000001c9 (
    .I0(b[1]),
    .I1(a[1]),
    .I2(b[0]),
    .I3(a[0]),
    .O(sig00000145)
  );
  LUT4 #(
    .INIT ( 16'h22B2 ))
  blk000001ca (
    .I0(b[29]),
    .I1(a[29]),
    .I2(b[28]),
    .I3(a[28]),
    .O(sig00000128)
  );
  LUT4 #(
    .INIT ( 16'h22B2 ))
  blk000001cb (
    .I0(b[27]),
    .I1(a[27]),
    .I2(b[26]),
    .I3(a[26]),
    .O(sig0000012a)
  );
  LUT4 #(
    .INIT ( 16'h22B2 ))
  blk000001cc (
    .I0(b[25]),
    .I1(a[25]),
    .I2(b[24]),
    .I3(a[24]),
    .O(sig0000012c)
  );
  LUT4 #(
    .INIT ( 16'h22B2 ))
  blk000001cd (
    .I0(b[23]),
    .I1(a[23]),
    .I2(b[22]),
    .I3(a[22]),
    .O(sig0000012e)
  );
  LUT4 #(
    .INIT ( 16'h22B2 ))
  blk000001ce (
    .I0(b[21]),
    .I1(a[21]),
    .I2(b[20]),
    .I3(a[20]),
    .O(sig00000130)
  );
  LUT4 #(
    .INIT ( 16'h22B2 ))
  blk000001cf (
    .I0(b[19]),
    .I1(a[19]),
    .I2(b[18]),
    .I3(a[18]),
    .O(sig00000132)
  );
  LUT4 #(
    .INIT ( 16'h22B2 ))
  blk000001d0 (
    .I0(b[17]),
    .I1(a[17]),
    .I2(b[16]),
    .I3(a[16]),
    .O(sig00000134)
  );
  LUT4 #(
    .INIT ( 16'h22B2 ))
  blk000001d1 (
    .I0(b[15]),
    .I1(a[15]),
    .I2(b[14]),
    .I3(a[14]),
    .O(sig00000136)
  );
  LUT4 #(
    .INIT ( 16'h22B2 ))
  blk000001d2 (
    .I0(b[13]),
    .I1(a[13]),
    .I2(b[12]),
    .I3(a[12]),
    .O(sig00000138)
  );
  LUT4 #(
    .INIT ( 16'h22B2 ))
  blk000001d3 (
    .I0(b[11]),
    .I1(a[11]),
    .I2(b[10]),
    .I3(a[10]),
    .O(sig0000013a)
  );
  LUT4 #(
    .INIT ( 16'h22B2 ))
  blk000001d4 (
    .I0(b[9]),
    .I1(a[9]),
    .I2(b[8]),
    .I3(a[8]),
    .O(sig0000013c)
  );
  LUT4 #(
    .INIT ( 16'h22B2 ))
  blk000001d5 (
    .I0(b[7]),
    .I1(a[7]),
    .I2(b[6]),
    .I3(a[6]),
    .O(sig0000013e)
  );
  LUT4 #(
    .INIT ( 16'h22B2 ))
  blk000001d6 (
    .I0(b[5]),
    .I1(a[5]),
    .I2(b[4]),
    .I3(a[4]),
    .O(sig00000140)
  );
  LUT4 #(
    .INIT ( 16'h22B2 ))
  blk000001d7 (
    .I0(b[3]),
    .I1(a[3]),
    .I2(b[2]),
    .I3(a[2]),
    .O(sig00000142)
  );
  LUT4 #(
    .INIT ( 16'h22B2 ))
  blk000001d8 (
    .I0(b[1]),
    .I1(a[1]),
    .I2(b[0]),
    .I3(a[0]),
    .O(sig00000144)
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  blk000001d9 (
    .I0(a[30]),
    .I1(b[30]),
    .O(sig00000126)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk000001da (
    .I0(a[30]),
    .I1(b[30]),
    .O(sig00000127)
  );
  LUT4 #(
    .INIT ( 16'h00AC ))
  blk000001db (
    .I0(sig0000001c),
    .I1(sig00000033),
    .I2(sig00000019),
    .I3(sig000001d2),
    .O(sig000001bc)
  );
  LUT4 #(
    .INIT ( 16'h00AC ))
  blk000001dc (
    .I0(sig0000001d),
    .I1(sig00000034),
    .I2(sig00000019),
    .I3(sig000001d2),
    .O(sig000001bb)
  );
  LUT4 #(
    .INIT ( 16'h00AC ))
  blk000001dd (
    .I0(sig0000001e),
    .I1(sig00000035),
    .I2(sig00000019),
    .I3(sig000001d2),
    .O(sig000001ba)
  );
  LUT4 #(
    .INIT ( 16'h00AC ))
  blk000001de (
    .I0(sig0000001f),
    .I1(sig00000036),
    .I2(sig00000019),
    .I3(sig000001d2),
    .O(sig000001b9)
  );
  LUT4 #(
    .INIT ( 16'h00AC ))
  blk000001df (
    .I0(sig00000020),
    .I1(sig00000037),
    .I2(sig00000019),
    .I3(sig000001d2),
    .O(sig000001b8)
  );
  LUT4 #(
    .INIT ( 16'h00AC ))
  blk000001e0 (
    .I0(sig00000021),
    .I1(sig00000038),
    .I2(sig00000019),
    .I3(sig000001d2),
    .O(sig000001b7)
  );
  LUT4 #(
    .INIT ( 16'h00AC ))
  blk000001e1 (
    .I0(sig00000022),
    .I1(sig00000039),
    .I2(sig00000019),
    .I3(sig000001d2),
    .O(sig000001b6)
  );
  LUT4 #(
    .INIT ( 16'h00AC ))
  blk000001e2 (
    .I0(sig00000023),
    .I1(sig0000003a),
    .I2(sig00000019),
    .I3(sig000001d2),
    .O(sig000001b5)
  );
  LUT4 #(
    .INIT ( 16'h00AC ))
  blk000001e3 (
    .I0(sig00000024),
    .I1(sig0000003b),
    .I2(sig00000019),
    .I3(sig000001d2),
    .O(sig000001b4)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk000001e4 (
    .I0(sig00000019),
    .I1(sig00000049),
    .I2(sig00000032),
    .O(sig000001d3)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk000001e5 (
    .I0(sig00000019),
    .I1(sig0000003f),
    .I2(sig00000028),
    .O(sig000001dd)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk000001e6 (
    .I0(sig00000019),
    .I1(sig0000003e),
    .I2(sig00000027),
    .O(sig000001de)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk000001e7 (
    .I0(sig00000019),
    .I1(sig0000003d),
    .I2(sig00000026),
    .O(sig000001df)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk000001e8 (
    .I0(sig00000019),
    .I1(sig0000003c),
    .I2(sig00000025),
    .O(sig000001e0)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk000001e9 (
    .I0(sig00000019),
    .I1(sig0000003b),
    .I2(sig00000024),
    .O(sig000001e1)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk000001ea (
    .I0(sig00000019),
    .I1(sig0000003a),
    .I2(sig00000023),
    .O(sig000001e2)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk000001eb (
    .I0(sig00000019),
    .I1(sig00000039),
    .I2(sig00000022),
    .O(sig000001e3)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk000001ec (
    .I0(sig00000019),
    .I1(sig00000038),
    .I2(sig00000021),
    .O(sig000001e4)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk000001ed (
    .I0(sig00000019),
    .I1(sig00000037),
    .I2(sig00000020),
    .O(sig000001e5)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk000001ee (
    .I0(sig00000019),
    .I1(sig00000036),
    .I2(sig0000001f),
    .O(sig000001e6)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk000001ef (
    .I0(sig00000019),
    .I1(sig00000048),
    .I2(sig00000031),
    .O(sig000001d4)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk000001f0 (
    .I0(sig00000019),
    .I1(sig00000035),
    .I2(sig0000001e),
    .O(sig000001e7)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk000001f1 (
    .I0(sig00000019),
    .I1(sig00000034),
    .I2(sig0000001d),
    .O(sig000001e8)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk000001f2 (
    .I0(sig00000019),
    .I1(sig00000033),
    .I2(sig0000001c),
    .O(sig000001e9)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk000001f3 (
    .I0(sig00000019),
    .I1(sig00000047),
    .I2(sig00000030),
    .O(sig000001d5)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk000001f4 (
    .I0(sig00000019),
    .I1(sig00000046),
    .I2(sig0000002f),
    .O(sig000001d6)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk000001f5 (
    .I0(sig00000019),
    .I1(sig00000045),
    .I2(sig0000002e),
    .O(sig000001d7)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk000001f6 (
    .I0(sig00000019),
    .I1(sig00000044),
    .I2(sig0000002d),
    .O(sig000001d8)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk000001f7 (
    .I0(sig00000019),
    .I1(sig00000043),
    .I2(sig0000002c),
    .O(sig000001d9)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk000001f8 (
    .I0(sig00000019),
    .I1(sig00000042),
    .I2(sig0000002b),
    .O(sig000001da)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk000001f9 (
    .I0(sig00000019),
    .I1(sig00000041),
    .I2(sig0000002a),
    .O(sig000001db)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk000001fa (
    .I0(sig00000019),
    .I1(sig00000040),
    .I2(sig00000029),
    .O(sig000001dc)
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  blk000001fb (
    .I0(sig000001f9),
    .I1(sig000001a3),
    .O(sig000001bf)
  );
  LUT4 #(
    .INIT ( 16'h1537 ))
  blk000001fc (
    .I0(sig0000004a),
    .I1(sig00000064),
    .I2(sig0000004b),
    .I3(sig00000063),
    .O(sig00000226)
  );
  LUT3 #(
    .INIT ( 8'hA2 ))
  blk000001fd (
    .I0(sig0000022e),
    .I1(sig0000022f),
    .I2(sig0000022d),
    .O(sig00000225)
  );
  LUT6 #(
    .INIT ( 64'hFBEAEAEA51404040 ))
  blk000001fe (
    .I0(sig0000004a),
    .I1(sig0000004b),
    .I2(sig00000062),
    .I3(sig00000063),
    .I4(sig0000004c),
    .I5(sig00000061),
    .O(sig00000227)
  );
  LUT6 #(
    .INIT ( 64'hFBEAEAEA51404040 ))
  blk000001ff (
    .I0(sig0000004a),
    .I1(sig0000004b),
    .I2(sig00000063),
    .I3(sig00000064),
    .I4(sig0000004c),
    .I5(sig00000062),
    .O(sig00000228)
  );
  LUT2 #(
    .INIT ( 4'h8 ))
  blk00000200 (
    .I0(sig0000024b),
    .I1(sig0000024a),
    .O(sig00000229)
  );
  LUT2 #(
    .INIT ( 4'h8 ))
  blk00000201 (
    .I0(sig00000230),
    .I1(sig00000065),
    .O(sig00000231)
  );
  LUT3 #(
    .INIT ( 8'hF1 ))
  blk00000202 (
    .I0(sig00000059),
    .I1(sig00000058),
    .I2(sig00000066),
    .O(sig00000264)
  );
  LUT3 #(
    .INIT ( 8'hF1 ))
  blk00000203 (
    .I0(sig00000057),
    .I1(sig00000056),
    .I2(sig00000066),
    .O(sig00000265)
  );
  LUT4 #(
    .INIT ( 16'h0F11 ))
  blk00000204 (
    .I0(sig00000055),
    .I1(sig00000054),
    .I2(sig00000064),
    .I3(sig00000066),
    .O(sig00000266)
  );
  LUT5 #(
    .INIT ( 32'h000F1111 ))
  blk00000205 (
    .I0(sig00000053),
    .I1(sig00000052),
    .I2(sig00000062),
    .I3(sig00000063),
    .I4(sig00000066),
    .O(sig00000267)
  );
  LUT5 #(
    .INIT ( 32'h000F1111 ))
  blk00000206 (
    .I0(sig0000004f),
    .I1(sig0000004e),
    .I2(sig0000005f),
    .I3(sig0000005e),
    .I4(sig00000066),
    .O(sig00000269)
  );
  LUT5 #(
    .INIT ( 32'h03030055 ))
  blk00000207 (
    .I0(sig0000004d),
    .I1(sig0000005d),
    .I2(sig0000005c),
    .I3(sig0000004c),
    .I4(sig00000066),
    .O(sig0000026a)
  );
  LUT5 #(
    .INIT ( 32'h000F1111 ))
  blk00000208 (
    .I0(sig00000051),
    .I1(sig00000050),
    .I2(sig00000060),
    .I3(sig00000061),
    .I4(sig00000066),
    .O(sig00000268)
  );
  LUT5 #(
    .INIT ( 32'h1111000F ))
  blk00000209 (
    .I0(sig0000005b),
    .I1(sig0000005a),
    .I2(sig0000004b),
    .I3(sig0000004a),
    .I4(sig00000066),
    .O(sig0000026b)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk0000020a (
    .I0(sig0000028b),
    .I1(sig00000289),
    .I2(sig0000028d),
    .O(sig00000286)
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  blk0000020b (
    .I0(sig00000066),
    .I1(sig0000005a),
    .O(sig00000299)
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  blk0000020c (
    .I0(sig00000066),
    .I1(sig00000059),
    .O(sig0000029a)
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  blk0000020d (
    .I0(sig00000066),
    .I1(sig00000058),
    .O(sig0000029b)
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  blk0000020e (
    .I0(sig00000066),
    .I1(sig00000057),
    .O(sig0000029c)
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  blk0000020f (
    .I0(sig00000066),
    .I1(sig00000056),
    .O(sig0000029d)
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  blk00000210 (
    .I0(sig00000066),
    .I1(sig00000055),
    .O(sig0000029e)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk00000211 (
    .I0(sig00000066),
    .I1(sig00000064),
    .I2(sig00000054),
    .O(sig0000029f)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk00000212 (
    .I0(sig00000066),
    .I1(sig00000063),
    .I2(sig00000053),
    .O(sig000002a0)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk00000213 (
    .I0(sig00000066),
    .I1(sig00000062),
    .I2(sig00000052),
    .O(sig000002a1)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk00000214 (
    .I0(sig00000066),
    .I1(sig00000061),
    .I2(sig00000051),
    .O(sig000002a2)
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  blk00000215 (
    .I0(sig00000066),
    .I1(sig00000063),
    .O(sig00000290)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk00000216 (
    .I0(sig00000066),
    .I1(sig00000060),
    .I2(sig00000050),
    .O(sig000002a3)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk00000217 (
    .I0(sig00000066),
    .I1(sig0000005f),
    .I2(sig0000004f),
    .O(sig000002a4)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk00000218 (
    .I0(sig00000066),
    .I1(sig0000005e),
    .I2(sig0000004e),
    .O(sig000002a5)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk00000219 (
    .I0(sig00000066),
    .I1(sig0000005d),
    .I2(sig0000004d),
    .O(sig000002a6)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk0000021a (
    .I0(sig00000066),
    .I1(sig0000005c),
    .I2(sig0000004c),
    .O(sig000002a7)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk0000021b (
    .I0(sig00000066),
    .I1(sig0000005b),
    .I2(sig0000004b),
    .O(sig000002a8)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk0000021c (
    .I0(sig00000066),
    .I1(sig0000005a),
    .I2(sig0000004a),
    .O(sig000002a9)
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  blk0000021d (
    .I0(sig00000066),
    .I1(sig00000062),
    .O(sig00000291)
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  blk0000021e (
    .I0(sig00000066),
    .I1(sig00000061),
    .O(sig00000292)
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  blk0000021f (
    .I0(sig00000066),
    .I1(sig00000060),
    .O(sig00000293)
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  blk00000220 (
    .I0(sig00000066),
    .I1(sig0000005f),
    .O(sig00000294)
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  blk00000221 (
    .I0(sig00000066),
    .I1(sig0000005e),
    .O(sig00000295)
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  blk00000222 (
    .I0(sig00000066),
    .I1(sig0000005d),
    .O(sig00000296)
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  blk00000223 (
    .I0(sig00000066),
    .I1(sig0000005c),
    .O(sig00000297)
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  blk00000224 (
    .I0(sig00000066),
    .I1(sig0000005b),
    .O(sig00000298)
  );
  LUT4 #(
    .INIT ( 16'h0020 ))
  blk00000225 (
    .I0(sig0000023c),
    .I1(sig0000023d),
    .I2(sig00000288),
    .I3(sig00000287),
    .O(sig0000026e)
  );
  LUT3 #(
    .INIT ( 8'h08 ))
  blk00000226 (
    .I0(sig0000023d),
    .I1(sig00000288),
    .I2(sig00000287),
    .O(sig0000026f)
  );
  LUT4 #(
    .INIT ( 16'h0020 ))
  blk00000227 (
    .I0(sig0000023e),
    .I1(sig0000023f),
    .I2(sig00000289),
    .I3(sig00000288),
    .O(sig00000270)
  );
  LUT3 #(
    .INIT ( 8'h08 ))
  blk00000228 (
    .I0(sig0000023f),
    .I1(sig00000289),
    .I2(sig00000288),
    .O(sig00000273)
  );
  LUT4 #(
    .INIT ( 16'h0020 ))
  blk00000229 (
    .I0(sig00000240),
    .I1(sig00000241),
    .I2(sig0000028a),
    .I3(sig00000289),
    .O(sig00000274)
  );
  LUT3 #(
    .INIT ( 8'h08 ))
  blk0000022a (
    .I0(sig00000241),
    .I1(sig0000028a),
    .I2(sig00000289),
    .O(sig00000275)
  );
  LUT4 #(
    .INIT ( 16'h0020 ))
  blk0000022b (
    .I0(sig00000242),
    .I1(sig00000243),
    .I2(sig0000028b),
    .I3(sig0000028a),
    .O(sig00000276)
  );
  LUT3 #(
    .INIT ( 8'h08 ))
  blk0000022c (
    .I0(sig00000243),
    .I1(sig0000028b),
    .I2(sig0000028a),
    .O(sig00000279)
  );
  LUT4 #(
    .INIT ( 16'h0020 ))
  blk0000022d (
    .I0(sig00000244),
    .I1(sig00000245),
    .I2(sig0000028c),
    .I3(sig0000028b),
    .O(sig0000027a)
  );
  LUT3 #(
    .INIT ( 8'h08 ))
  blk0000022e (
    .I0(sig00000245),
    .I1(sig0000028c),
    .I2(sig0000028b),
    .O(sig0000027b)
  );
  LUT4 #(
    .INIT ( 16'h0020 ))
  blk0000022f (
    .I0(sig00000246),
    .I1(sig00000247),
    .I2(sig0000028d),
    .I3(sig0000028c),
    .O(sig0000027c)
  );
  LUT3 #(
    .INIT ( 8'h08 ))
  blk00000230 (
    .I0(sig00000247),
    .I1(sig0000028d),
    .I2(sig0000028c),
    .O(sig0000027f)
  );
  LUT4 #(
    .INIT ( 16'h0020 ))
  blk00000231 (
    .I0(sig00000248),
    .I1(sig00000249),
    .I2(sig0000028e),
    .I3(sig0000028d),
    .O(sig00000280)
  );
  LUT3 #(
    .INIT ( 8'h08 ))
  blk00000232 (
    .I0(sig00000249),
    .I1(sig0000028e),
    .I2(sig0000028d),
    .O(sig00000281)
  );
  LUT3 #(
    .INIT ( 8'h02 ))
  blk00000233 (
    .I0(sig0000024b),
    .I1(sig0000024a),
    .I2(sig0000028e),
    .O(sig00000282)
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  blk00000234 (
    .I0(sig0000028e),
    .I1(sig0000024a),
    .O(sig00000285)
  );
  LUT2 #(
    .INIT ( 4'h8 ))
  blk00000235 (
    .I0(sig0000028f),
    .I1(sig00000287),
    .O(sig0000008b)
  );
  LUT4 #(
    .INIT ( 16'h7520 ))
  blk00000236 (
    .I0(ce),
    .I1(sig0000000c),
    .I2(sig00000082),
    .I3(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.DSP.OP/OP/mant_op [0]),
    .O(sig000002aa)
  );
  LUT4 #(
    .INIT ( 16'h7520 ))
  blk00000237 (
    .I0(ce),
    .I1(sig0000000c),
    .I2(sig00000081),
    .I3(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.DSP.OP/OP/mant_op [1]),
    .O(sig000002ab)
  );
  LUT4 #(
    .INIT ( 16'h7520 ))
  blk00000238 (
    .I0(ce),
    .I1(sig0000000c),
    .I2(sig0000007f),
    .I3(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.DSP.OP/OP/mant_op [3]),
    .O(sig000002ad)
  );
  LUT4 #(
    .INIT ( 16'h7520 ))
  blk00000239 (
    .I0(ce),
    .I1(sig0000000c),
    .I2(sig0000007e),
    .I3(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.DSP.OP/OP/mant_op [4]),
    .O(sig000002ae)
  );
  LUT4 #(
    .INIT ( 16'h7520 ))
  blk0000023a (
    .I0(ce),
    .I1(sig0000000c),
    .I2(sig00000080),
    .I3(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.DSP.OP/OP/mant_op [2]),
    .O(sig000002ac)
  );
  LUT4 #(
    .INIT ( 16'h7520 ))
  blk0000023b (
    .I0(ce),
    .I1(sig0000000c),
    .I2(sig0000007d),
    .I3(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.DSP.OP/OP/mant_op [5]),
    .O(sig000002af)
  );
  LUT4 #(
    .INIT ( 16'h7520 ))
  blk0000023c (
    .I0(ce),
    .I1(sig0000000c),
    .I2(sig0000007c),
    .I3(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.DSP.OP/OP/mant_op [6]),
    .O(sig000002b0)
  );
  LUT4 #(
    .INIT ( 16'h7520 ))
  blk0000023d (
    .I0(ce),
    .I1(sig0000000c),
    .I2(sig0000007b),
    .I3(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.DSP.OP/OP/mant_op [7]),
    .O(sig000002b1)
  );
  LUT4 #(
    .INIT ( 16'h7520 ))
  blk0000023e (
    .I0(ce),
    .I1(sig0000000c),
    .I2(sig0000007a),
    .I3(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.DSP.OP/OP/mant_op [8]),
    .O(sig000002b2)
  );
  LUT4 #(
    .INIT ( 16'h7520 ))
  blk0000023f (
    .I0(ce),
    .I1(sig0000000c),
    .I2(sig00000079),
    .I3(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.DSP.OP/OP/mant_op [9]),
    .O(sig000002b3)
  );
  LUT4 #(
    .INIT ( 16'h7520 ))
  blk00000240 (
    .I0(ce),
    .I1(sig0000000c),
    .I2(sig00000078),
    .I3(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.DSP.OP/OP/mant_op [10]),
    .O(sig000002b4)
  );
  LUT4 #(
    .INIT ( 16'h7520 ))
  blk00000241 (
    .I0(ce),
    .I1(sig0000000c),
    .I2(sig00000076),
    .I3(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.DSP.OP/OP/mant_op [12]),
    .O(sig000002b6)
  );
  LUT4 #(
    .INIT ( 16'h7520 ))
  blk00000242 (
    .I0(ce),
    .I1(sig0000000c),
    .I2(sig00000075),
    .I3(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.DSP.OP/OP/mant_op [13]),
    .O(sig000002b7)
  );
  LUT4 #(
    .INIT ( 16'h7520 ))
  blk00000243 (
    .I0(ce),
    .I1(sig0000000c),
    .I2(sig00000077),
    .I3(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.DSP.OP/OP/mant_op [11]),
    .O(sig000002b5)
  );
  LUT4 #(
    .INIT ( 16'h7520 ))
  blk00000244 (
    .I0(ce),
    .I1(sig0000000c),
    .I2(sig00000074),
    .I3(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.DSP.OP/OP/mant_op [14]),
    .O(sig000002b8)
  );
  LUT4 #(
    .INIT ( 16'h7520 ))
  blk00000245 (
    .I0(ce),
    .I1(sig0000000c),
    .I2(sig00000073),
    .I3(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.DSP.OP/OP/mant_op [15]),
    .O(sig000002b9)
  );
  LUT4 #(
    .INIT ( 16'h7520 ))
  blk00000246 (
    .I0(ce),
    .I1(sig0000000c),
    .I2(sig00000072),
    .I3(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.DSP.OP/OP/mant_op [16]),
    .O(sig000002ba)
  );
  LUT4 #(
    .INIT ( 16'h7520 ))
  blk00000247 (
    .I0(ce),
    .I1(sig0000000c),
    .I2(sig00000071),
    .I3(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.DSP.OP/OP/mant_op [17]),
    .O(sig000002bb)
  );
  LUT4 #(
    .INIT ( 16'h7520 ))
  blk00000248 (
    .I0(ce),
    .I1(sig0000000c),
    .I2(sig00000070),
    .I3(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.DSP.OP/OP/mant_op [18]),
    .O(sig000002bc)
  );
  LUT4 #(
    .INIT ( 16'h7520 ))
  blk00000249 (
    .I0(ce),
    .I1(sig0000000c),
    .I2(sig0000006f),
    .I3(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.DSP.OP/OP/mant_op [19]),
    .O(sig000002bd)
  );
  LUT4 #(
    .INIT ( 16'h7520 ))
  blk0000024a (
    .I0(ce),
    .I1(sig0000000c),
    .I2(sig0000006d),
    .I3(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.DSP.OP/OP/mant_op [21]),
    .O(sig000002bf)
  );
  LUT4 #(
    .INIT ( 16'h7520 ))
  blk0000024b (
    .I0(ce),
    .I1(sig0000000c),
    .I2(sig0000006e),
    .I3(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.DSP.OP/OP/mant_op [20]),
    .O(sig000002be)
  );
  LUT5 #(
    .INIT ( 32'h77752220 ))
  blk0000024c (
    .I0(ce),
    .I1(sig0000000d),
    .I2(sig0000000e),
    .I3(sig0000006c),
    .I4(\NlwRenamedSig_OI_U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.DSP.OP/OP/mant_op [22]),
    .O(sig000002c0)
  );
  LUT2 #(
    .INIT ( 4'h8 ))
  blk0000024d (
    .I0(sig0000000f),
    .I1(ce),
    .O(sig000002c1)
  );
  LUT4 #(
    .INIT ( 16'hF7FF ))
  blk0000024e (
    .I0(sig00000013),
    .I1(sig00000015),
    .I2(sig000000e2),
    .I3(sig00000014),
    .O(sig000002c2)
  );
  LUT6 #(
    .INIT ( 64'h0000000080000000 ))
  blk0000024f (
    .I0(sig00000017),
    .I1(sig00000018),
    .I2(sig00000016),
    .I3(sig00000011),
    .I4(sig00000012),
    .I5(sig000002c2),
    .O(sig000000bf)
  );
  LUT3 #(
    .INIT ( 8'hD8 ))
  blk00000250 (
    .I0(sig000000f8),
    .I1(sig000000f7),
    .I2(sig000000f6),
    .O(sig000002c3)
  );
  LUT5 #(
    .INIT ( 32'hAA0BAA08 ))
  blk00000251 (
    .I0(sig000000f9),
    .I1(sig000000fa),
    .I2(sig000000fb),
    .I3(sig000000fc),
    .I4(sig000002c3),
    .O(sig000000ce)
  );
  LUT3 #(
    .INIT ( 8'h80 ))
  blk00000252 (
    .I0(a[25]),
    .I1(a[24]),
    .I2(a[23]),
    .O(sig000002c4)
  );
  LUT6 #(
    .INIT ( 64'h8000000000000000 ))
  blk00000253 (
    .I0(a[30]),
    .I1(a[29]),
    .I2(a[28]),
    .I3(a[27]),
    .I4(a[26]),
    .I5(sig000002c4),
    .O(sig000000b2)
  );
  LUT3 #(
    .INIT ( 8'hFE ))
  blk00000254 (
    .I0(a[25]),
    .I1(a[24]),
    .I2(a[23]),
    .O(sig000002c5)
  );
  LUT6 #(
    .INIT ( 64'h0000000000000001 ))
  blk00000255 (
    .I0(a[30]),
    .I1(a[29]),
    .I2(a[28]),
    .I3(a[27]),
    .I4(a[26]),
    .I5(sig000002c5),
    .O(sig000000b3)
  );
  LUT3 #(
    .INIT ( 8'h80 ))
  blk00000256 (
    .I0(b[25]),
    .I1(b[24]),
    .I2(b[23]),
    .O(sig000002c6)
  );
  LUT6 #(
    .INIT ( 64'h8000000000000000 ))
  blk00000257 (
    .I0(b[30]),
    .I1(b[29]),
    .I2(b[28]),
    .I3(b[27]),
    .I4(b[26]),
    .I5(sig000002c6),
    .O(sig000000b4)
  );
  LUT3 #(
    .INIT ( 8'hFE ))
  blk00000258 (
    .I0(b[25]),
    .I1(b[24]),
    .I2(b[23]),
    .O(sig000002c7)
  );
  LUT6 #(
    .INIT ( 64'h0000000000000001 ))
  blk00000259 (
    .I0(b[30]),
    .I1(b[29]),
    .I2(b[28]),
    .I3(b[27]),
    .I4(b[26]),
    .I5(sig000002c7),
    .O(sig000000b5)
  );
  LUT4 #(
    .INIT ( 16'hFFFE ))
  blk0000025a (
    .I0(sig00000013),
    .I1(sig00000015),
    .I2(sig00000014),
    .I3(sig000000e2),
    .O(sig000002c8)
  );
  LUT6 #(
    .INIT ( 64'h0000000000000001 ))
  blk0000025b (
    .I0(sig00000017),
    .I1(sig00000018),
    .I2(sig00000016),
    .I3(sig00000011),
    .I4(sig00000012),
    .I5(sig000002c8),
    .O(sig000000be)
  );
  LUT2 #(
    .INIT ( 4'hE ))
  blk0000025c (
    .I0(sig00000110),
    .I1(sig00000113),
    .O(sig000002c9)
  );
  LUT6 #(
    .INIT ( 64'h0000000000008001 ))
  blk0000025d (
    .I0(sig00000005),
    .I1(sig00000004),
    .I2(sig00000003),
    .I3(sig00000006),
    .I4(sig000002c9),
    .I5(sig000001d1),
    .O(sig000001c0)
  );
  LUT6 #(
    .INIT ( 64'h0000000000010000 ))
  blk0000025e (
    .I0(sig000001ed),
    .I1(sig000001ee),
    .I2(sig000001ef),
    .I3(sig000001f0),
    .I4(sig000001f7),
    .I5(sig000001f1),
    .O(sig000002ca)
  );
  LUT6 #(
    .INIT ( 64'h0000000000000001 ))
  blk0000025f (
    .I0(sig000001f3),
    .I1(sig000001f2),
    .I2(sig000001f4),
    .I3(sig000001f5),
    .I4(sig000001ea),
    .I5(sig000001eb),
    .O(sig000002cb)
  );
  LUT4 #(
    .INIT ( 16'h0020 ))
  blk00000260 (
    .I0(sig000002cb),
    .I1(sig000001f6),
    .I2(sig000002ca),
    .I3(sig000001ec),
    .O(sig000001be)
  );
  LUT3 #(
    .INIT ( 8'h1B ))
  blk00000261 (
    .I0(sig0000028d),
    .I1(sig00000283),
    .I2(sig0000027d),
    .O(sig000002cc)
  );
  LUT5 #(
    .INIT ( 32'h8A80DFD5 ))
  blk00000262 (
    .I0(sig0000028b),
    .I1(sig00000271),
    .I2(sig00000289),
    .I3(sig00000277),
    .I4(sig000002cc),
    .O(sig0000026c)
  );
  LUT3 #(
    .INIT ( 8'h1B ))
  blk00000263 (
    .I0(sig0000028d),
    .I1(sig00000284),
    .I2(sig0000027e),
    .O(sig000002cd)
  );
  LUT5 #(
    .INIT ( 32'h8A80DFD5 ))
  blk00000264 (
    .I0(sig0000028b),
    .I1(sig00000272),
    .I2(sig00000289),
    .I3(sig00000278),
    .I4(sig000002cd),
    .O(sig0000026d)
  );
  FDRE   blk00000265 (
    .C(clk),
    .CE(ce),
    .D(sig000002ce),
    .R(sig000002c1),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.DSP.OP/OP/exp_op [7])
  );
  LUT2 #(
    .INIT ( 4'hE ))
  blk00000266 (
    .I0(sig00000083),
    .I1(sig00000010),
    .O(sig000002ce)
  );
  FDRE   blk00000267 (
    .C(clk),
    .CE(ce),
    .D(sig000002cf),
    .R(sig000002c1),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.DSP.OP/OP/exp_op [6])
  );
  LUT2 #(
    .INIT ( 4'hE ))
  blk00000268 (
    .I0(sig00000084),
    .I1(sig00000010),
    .O(sig000002cf)
  );
  FDRE   blk00000269 (
    .C(clk),
    .CE(ce),
    .D(sig000002d0),
    .R(sig000002c1),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.DSP.OP/OP/exp_op [5])
  );
  LUT2 #(
    .INIT ( 4'hE ))
  blk0000026a (
    .I0(sig00000085),
    .I1(sig00000010),
    .O(sig000002d0)
  );
  FDRE   blk0000026b (
    .C(clk),
    .CE(ce),
    .D(sig000002d1),
    .R(sig000002c1),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.DSP.OP/OP/exp_op [4])
  );
  LUT2 #(
    .INIT ( 4'hE ))
  blk0000026c (
    .I0(sig00000086),
    .I1(sig00000010),
    .O(sig000002d1)
  );
  FDRE   blk0000026d (
    .C(clk),
    .CE(ce),
    .D(sig000002d2),
    .R(sig000002c1),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.DSP.OP/OP/exp_op [3])
  );
  LUT2 #(
    .INIT ( 4'hE ))
  blk0000026e (
    .I0(sig00000087),
    .I1(sig00000010),
    .O(sig000002d2)
  );
  FDRE   blk0000026f (
    .C(clk),
    .CE(ce),
    .D(sig000002d3),
    .R(sig000002c1),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.DSP.OP/OP/exp_op [2])
  );
  LUT2 #(
    .INIT ( 4'hE ))
  blk00000270 (
    .I0(sig00000088),
    .I1(sig00000010),
    .O(sig000002d3)
  );
  FDRE   blk00000271 (
    .C(clk),
    .CE(ce),
    .D(sig000002d4),
    .R(sig000002c1),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.DSP.OP/OP/exp_op [1])
  );
  LUT2 #(
    .INIT ( 4'hE ))
  blk00000272 (
    .I0(sig00000089),
    .I1(sig00000010),
    .O(sig000002d4)
  );
  FDRE   blk00000273 (
    .C(clk),
    .CE(ce),
    .D(sig000002d5),
    .R(sig000002c1),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.DSP.OP/OP/exp_op [0])
  );
  LUT2 #(
    .INIT ( 4'hE ))
  blk00000274 (
    .I0(sig0000008a),
    .I1(sig00000010),
    .O(sig000002d5)
  );
  FDE   blk00000275 (
    .C(clk),
    .CE(ce),
    .D(sig0000001b),
    .Q(\U0/op_inst/FLT_PT_OP/ADDSUB_OP.SPEED_OP.DSP.OP/OP/sign_op )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  blk00000276 (
    .I0(sig000001d2),
    .O(sig000002d6)
  );
  LUT5 #(
    .INIT ( 32'h02020257 ))
  blk00000277 (
    .I0(sig00000019),
    .I1(sig00000031),
    .I2(sig00000032),
    .I3(sig00000048),
    .I4(sig00000049),
    .O(sig00000221)
  );
  LUT5 #(
    .INIT ( 32'h02020257 ))
  blk00000278 (
    .I0(sig00000019),
    .I1(sig0000002f),
    .I2(sig00000030),
    .I3(sig00000046),
    .I4(sig00000047),
    .O(sig00000220)
  );
  LUT6 #(
    .INIT ( 64'hF0F0FF00CCCCAAAA ))
  blk00000279 (
    .I0(sig00000046),
    .I1(sig0000002f),
    .I2(sig00000021),
    .I3(sig00000038),
    .I4(sig00000019),
    .I5(sig000001d2),
    .O(sig000001a9)
  );
  LUT6 #(
    .INIT ( 64'hF0F0FF00CCCCAAAA ))
  blk0000027a (
    .I0(sig00000047),
    .I1(sig00000030),
    .I2(sig00000022),
    .I3(sig00000039),
    .I4(sig00000019),
    .I5(sig000001d2),
    .O(sig000001a8)
  );
  LUT6 #(
    .INIT ( 64'hF0F0FF00CCCCAAAA ))
  blk0000027b (
    .I0(sig00000048),
    .I1(sig00000031),
    .I2(sig00000023),
    .I3(sig0000003a),
    .I4(sig00000019),
    .I5(sig000001d2),
    .O(sig000001a7)
  );
  LUT6 #(
    .INIT ( 64'hF0F0FF00CCCCAAAA ))
  blk0000027c (
    .I0(sig00000049),
    .I1(sig00000032),
    .I2(sig00000024),
    .I3(sig0000003b),
    .I4(sig00000019),
    .I5(sig000001d2),
    .O(sig000001a6)
  );
  LUT5 #(
    .INIT ( 32'h02020257 ))
  blk0000027d (
    .I0(sig00000019),
    .I1(sig0000002e),
    .I2(sig0000002d),
    .I3(sig00000045),
    .I4(sig00000044),
    .O(sig0000021f)
  );
  LUT5 #(
    .INIT ( 32'h02020257 ))
  blk0000027e (
    .I0(sig00000019),
    .I1(sig0000002c),
    .I2(sig0000002b),
    .I3(sig00000043),
    .I4(sig00000042),
    .O(sig0000021e)
  );
  LUT5 #(
    .INIT ( 32'h02020257 ))
  blk0000027f (
    .I0(sig00000019),
    .I1(sig0000002a),
    .I2(sig00000029),
    .I3(sig00000041),
    .I4(sig00000040),
    .O(sig0000021d)
  );
  LUT5 #(
    .INIT ( 32'h02020257 ))
  blk00000280 (
    .I0(sig00000019),
    .I1(sig00000028),
    .I2(sig00000027),
    .I3(sig0000003f),
    .I4(sig0000003e),
    .O(sig0000021c)
  );
  LUT5 #(
    .INIT ( 32'h02020257 ))
  blk00000281 (
    .I0(sig00000019),
    .I1(sig00000026),
    .I2(sig00000025),
    .I3(sig0000003d),
    .I4(sig0000003c),
    .O(sig0000021b)
  );
  LUT2 #(
    .INIT ( 4'h7 ))
  blk00000282 (
    .I0(sig00000110),
    .I1(sig00000113),
    .O(sig000001fc)
  );
  LUT6 #(
    .INIT ( 64'hF0F0FF00CCCCAAAA ))
  blk00000283 (
    .I0(sig00000041),
    .I1(sig0000002a),
    .I2(sig0000001c),
    .I3(sig00000033),
    .I4(sig00000019),
    .I5(sig000001d2),
    .O(sig000001ae)
  );
  LUT6 #(
    .INIT ( 64'hF0F0FF00CCCCAAAA ))
  blk00000284 (
    .I0(sig00000042),
    .I1(sig0000002b),
    .I2(sig0000001d),
    .I3(sig00000034),
    .I4(sig00000019),
    .I5(sig000001d2),
    .O(sig000001ad)
  );
  LUT6 #(
    .INIT ( 64'hF0F0FF00CCCCAAAA ))
  blk00000285 (
    .I0(sig00000043),
    .I1(sig0000002c),
    .I2(sig0000001e),
    .I3(sig00000035),
    .I4(sig00000019),
    .I5(sig000001d2),
    .O(sig000001ac)
  );
  LUT6 #(
    .INIT ( 64'hF0F0FF00CCCCAAAA ))
  blk00000286 (
    .I0(sig00000044),
    .I1(sig0000002d),
    .I2(sig0000001f),
    .I3(sig00000036),
    .I4(sig00000019),
    .I5(sig000001d2),
    .O(sig000001ab)
  );
  LUT6 #(
    .INIT ( 64'hF0F0FF00CCCCAAAA ))
  blk00000287 (
    .I0(sig00000045),
    .I1(sig0000002e),
    .I2(sig00000020),
    .I3(sig00000037),
    .I4(sig00000019),
    .I5(sig000001d2),
    .O(sig000001aa)
  );
  LUT4 #(
    .INIT ( 16'h00AC ))
  blk00000288 (
    .I0(sig00000028),
    .I1(sig0000003f),
    .I2(sig00000019),
    .I3(sig000001d2),
    .O(sig000001b0)
  );
  LUT4 #(
    .INIT ( 16'h00AC ))
  blk00000289 (
    .I0(sig00000027),
    .I1(sig0000003e),
    .I2(sig00000019),
    .I3(sig000001d2),
    .O(sig000001b1)
  );
  LUT4 #(
    .INIT ( 16'h00AC ))
  blk0000028a (
    .I0(sig00000026),
    .I1(sig0000003d),
    .I2(sig00000019),
    .I3(sig000001d2),
    .O(sig000001b2)
  );
  LUT4 #(
    .INIT ( 16'h00AC ))
  blk0000028b (
    .I0(sig00000025),
    .I1(sig0000003c),
    .I2(sig00000019),
    .I3(sig000001d2),
    .O(sig000001b3)
  );
  LUT4 #(
    .INIT ( 16'hFFD8 ))
  blk0000028c (
    .I0(sig00000019),
    .I1(sig00000029),
    .I2(sig00000040),
    .I3(sig000001d2),
    .O(sig000001af)
  );
  INV   blk0000028d (
    .I(sig000001d2),
    .O(sig000001bd)
  );
  INV   blk0000028e (
    .I(sig000000e8),
    .O(sig00000092)
  );
  INV   blk0000028f (
    .I(sig000000e9),
    .O(sig00000090)
  );
  INV   blk00000290 (
    .I(sig000000ea),
    .O(sig0000008e)
  );
  LUT6 #(
    .INIT ( 64'h0818181018181810 ))
  blk00000291 (
    .I0(sig00000008),
    .I1(sig00000007),
    .I2(sig00000006),
    .I3(sig0000000a),
    .I4(sig00000009),
    .I5(sig0000000b),
    .O(sig000001d1)
  );
  LUT6 #(
    .INIT ( 64'h666666666666666A ))
  blk00000292 (
    .I0(sig00000007),
    .I1(sig00000006),
    .I2(sig00000008),
    .I3(sig00000009),
    .I4(sig0000000a),
    .I5(sig0000000b),
    .O(sig000001d2)
  );
  LUT5 #(
    .INIT ( 32'h00000001 ))
  blk00000293 (
    .I0(sig0000000b),
    .I1(sig0000000a),
    .I2(sig00000009),
    .I3(sig00000008),
    .I4(sig00000007),
    .O(sig000001d0)
  );
  LUT6 #(
    .INIT ( 64'h8000000000000002 ))
  blk00000294 (
    .I0(sig0000000b),
    .I1(sig0000000a),
    .I2(sig00000009),
    .I3(sig00000008),
    .I4(sig00000007),
    .I5(sig00000006),
    .O(sig000001cf)
  );
  LUT6 #(
    .INIT ( 64'h4001000000010004 ))
  blk00000295 (
    .I0(sig0000000b),
    .I1(sig0000000a),
    .I2(sig00000009),
    .I3(sig00000008),
    .I4(sig00000007),
    .I5(sig00000006),
    .O(sig000001ce)
  );
  LUT6 #(
    .INIT ( 64'h2800000000000028 ))
  blk00000296 (
    .I0(sig0000000b),
    .I1(sig0000000a),
    .I2(sig00000007),
    .I3(sig00000009),
    .I4(sig00000008),
    .I5(sig00000006),
    .O(sig000001cd)
  );
  LUT6 #(
    .INIT ( 64'h0400400000100004 ))
  blk00000297 (
    .I0(sig0000000b),
    .I1(sig00000009),
    .I2(sig0000000a),
    .I3(sig00000008),
    .I4(sig00000007),
    .I5(sig00000006),
    .O(sig000001cc)
  );
  LUT6 #(
    .INIT ( 64'h0820000000000820 ))
  blk00000298 (
    .I0(sig0000000b),
    .I1(sig0000000a),
    .I2(sig00000009),
    .I3(sig00000007),
    .I4(sig00000008),
    .I5(sig00000006),
    .O(sig000001cb)
  );
  LUT6 #(
    .INIT ( 64'h1000040000040040 ))
  blk00000299 (
    .I0(sig0000000b),
    .I1(sig00000009),
    .I2(sig0000000a),
    .I3(sig00000008),
    .I4(sig00000007),
    .I5(sig00000006),
    .O(sig000001ca)
  );
  LUT6 #(
    .INIT ( 64'h0000002828000000 ))
  blk0000029a (
    .I0(sig0000000b),
    .I1(sig00000007),
    .I2(sig0000000a),
    .I3(sig00000006),
    .I4(sig00000008),
    .I5(sig00000009),
    .O(sig000001c9)
  );
  LUT6 #(
    .INIT ( 64'h0010100004000010 ))
  blk0000029b (
    .I0(sig0000000b),
    .I1(sig00000009),
    .I2(sig00000008),
    .I3(sig0000000a),
    .I4(sig00000007),
    .I5(sig00000006),
    .O(sig000001c8)
  );
  LUT5 #(
    .INIT ( 32'h00800200 ))
  blk0000029c (
    .I0(sig0000000b),
    .I1(sig0000000a),
    .I2(sig00000009),
    .I3(sig00000008),
    .I4(sig00000007),
    .O(sig000001c7)
  );
  LUT6 #(
    .INIT ( 64'h0400001000101000 ))
  blk0000029d (
    .I0(sig0000000b),
    .I1(sig00000009),
    .I2(sig00000008),
    .I3(sig0000000a),
    .I4(sig00000007),
    .I5(sig00000006),
    .O(sig000001c6)
  );
  LUT6 #(
    .INIT ( 64'h0000002828000000 ))
  blk0000029e (
    .I0(sig0000000b),
    .I1(sig00000007),
    .I2(sig0000000a),
    .I3(sig00000006),
    .I4(sig00000009),
    .I5(sig00000008),
    .O(sig000001c5)
  );
  LUT6 #(
    .INIT ( 64'h0010000404004000 ))
  blk0000029f (
    .I0(sig0000000b),
    .I1(sig00000009),
    .I2(sig0000000a),
    .I3(sig00000006),
    .I4(sig00000007),
    .I5(sig00000008),
    .O(sig000001c4)
  );
  LUT6 #(
    .INIT ( 64'h0000002828000000 ))
  blk000002a0 (
    .I0(sig0000000b),
    .I1(sig00000006),
    .I2(sig00000008),
    .I3(sig00000007),
    .I4(sig0000000a),
    .I5(sig00000009),
    .O(sig000001c3)
  );
  LUT6 #(
    .INIT ( 64'h0010000404004000 ))
  blk000002a1 (
    .I0(sig0000000b),
    .I1(sig00000009),
    .I2(sig0000000a),
    .I3(sig00000008),
    .I4(sig00000007),
    .I5(sig00000006),
    .O(sig000001c2)
  );
  LUT6 #(
    .INIT ( 64'h0000002828000000 ))
  blk000002a2 (
    .I0(sig0000000b),
    .I1(sig00000007),
    .I2(sig0000000a),
    .I3(sig00000008),
    .I4(sig00000009),
    .I5(sig00000006),
    .O(sig000001c1)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000002a3 (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000001),
    .A3(sig00000002),
    .CE(ce),
    .CLK(clk),
    .D(sig000000b0),
    .Q(sig000002d7),
    .Q15(NLW_blk000002a3_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002a4 (
    .C(clk),
    .CE(ce),
    .D(sig000002d7),
    .Q(sig000000f3)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000002a5 (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(ce),
    .CLK(clk),
    .D(sig000000b1),
    .Q(sig000002d8),
    .Q15(NLW_blk000002a5_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002a6 (
    .C(clk),
    .CE(ce),
    .D(sig000002d8),
    .Q(sig0000010f)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000002a7 (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000001),
    .A3(sig00000002),
    .CE(ce),
    .CLK(clk),
    .D(sig00000157),
    .Q(sig000002d9),
    .Q15(NLW_blk000002a7_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002a8 (
    .C(clk),
    .CE(ce),
    .D(sig000002d9),
    .Q(sig000000f5)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000002a9 (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000001),
    .A3(sig00000002),
    .CE(ce),
    .CLK(clk),
    .D(sig00000156),
    .Q(sig000002da),
    .Q15(NLW_blk000002a9_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002aa (
    .C(clk),
    .CE(ce),
    .D(sig000002da),
    .Q(sig000000f4)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000002ab (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000001),
    .A3(sig00000002),
    .CE(ce),
    .CLK(clk),
    .D(sig000000f0),
    .Q(sig000002db),
    .Q15(NLW_blk000002ab_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002ac (
    .C(clk),
    .CE(ce),
    .D(sig000002db),
    .Q(sig000000e8)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000002ad (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000001),
    .A3(sig00000002),
    .CE(ce),
    .CLK(clk),
    .D(sig000000f2),
    .Q(sig000002dc),
    .Q15(NLW_blk000002ad_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002ae (
    .C(clk),
    .CE(ce),
    .D(sig000002dc),
    .Q(sig000000ea)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000002af (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000001),
    .A3(sig00000002),
    .CE(ce),
    .CLK(clk),
    .D(sig000000f1),
    .Q(sig000002dd),
    .Q15(NLW_blk000002af_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002b0 (
    .C(clk),
    .CE(ce),
    .D(sig000002dd),
    .Q(sig000000e9)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000002b1 (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000001),
    .A3(sig00000002),
    .CE(ce),
    .CLK(clk),
    .D(sig000000ef),
    .Q(sig000002de),
    .Q15(NLW_blk000002b1_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002b2 (
    .C(clk),
    .CE(ce),
    .D(sig000002de),
    .Q(sig000000e7)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000002b3 (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000001),
    .A3(sig00000002),
    .CE(ce),
    .CLK(clk),
    .D(sig000000ee),
    .Q(sig000002df),
    .Q15(NLW_blk000002b3_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002b4 (
    .C(clk),
    .CE(ce),
    .D(sig000002df),
    .Q(sig000000e6)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000002b5 (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000001),
    .A3(sig00000002),
    .CE(ce),
    .CLK(clk),
    .D(sig000000ed),
    .Q(sig000002e0),
    .Q15(NLW_blk000002b5_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002b6 (
    .C(clk),
    .CE(ce),
    .D(sig000002e0),
    .Q(sig000000e5)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000002b7 (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000001),
    .A3(sig00000002),
    .CE(ce),
    .CLK(clk),
    .D(sig000000ec),
    .Q(sig000002e1),
    .Q15(NLW_blk000002b7_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002b8 (
    .C(clk),
    .CE(ce),
    .D(sig000002e1),
    .Q(sig000000e4)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000002b9 (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(ce),
    .CLK(clk),
    .D(sig0000024b),
    .Q(sig000002e2),
    .Q15(NLW_blk000002b9_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002ba (
    .C(clk),
    .CE(ce),
    .D(sig000002e2),
    .Q(sig0000022b)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000002bb (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000001),
    .A3(sig00000002),
    .CE(ce),
    .CLK(clk),
    .D(sig000000eb),
    .Q(sig000002e3),
    .Q15(NLW_blk000002bb_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002bc (
    .C(clk),
    .CE(ce),
    .D(sig000002e3),
    .Q(sig000000e3)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk000002bd (
    .A0(sig00000001),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(ce),
    .CLK(clk),
    .D(sig000001f9),
    .Q(sig000002e4),
    .Q15(NLW_blk000002bd_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000002be (
    .C(clk),
    .CE(ce),
    .D(sig000002e4),
    .Q(sig000001f7)
  );
  DSP48E #(
    .ACASCREG ( 1 ),
    .ALUMODEREG ( 1 ),
    .AREG ( 1 ),
    .AUTORESET_PATTERN_DETECT ( 0 ),
    .AUTORESET_PATTERN_DETECT_OPTINV ( "MATCH" ),
    .A_INPUT ( "DIRECT" ),
    .BCASCREG ( 1 ),
    .BREG ( 1 ),
    .B_INPUT ( "DIRECT" ),
    .CARRYINREG ( 1 ),
    .CARRYINSELREG ( 1 ),
    .CREG ( 1 ),
    .MASK ( 48'hFF0000FFFFFF ),
    .MREG ( 1 ),
    .MULTCARRYINREG ( 0 ),
    .OPMODEREG ( 1 ),
    .PATTERN ( 48'h000000000000 ),
    .PREG ( 1 ),
    .SEL_MASK ( "MASK" ),
    .SEL_PATTERN ( "PATTERN" ),
    .SEL_ROUNDING_MASK ( "SEL_MASK" ),
    .SIM_MODE ( "SAFE" ),
    .USE_MULT ( "MULT_S" ),
    .USE_PATTERN_DETECT ( "PATDET" ),
    .USE_SIMD ( "ONE48" ))
  blk000002bf (
    .CEM(ce),
    .PATTERNDETECT(sig00000066),
    .CLK(clk),
    .CARRYIN(sig000001f8),
    .PATTERNBDETECT(NLW_blk000002bf_PATTERNBDETECT_UNCONNECTED),
    .RSTC(sig00000002),
    .CEB1(sig00000002),
    .MULTSIGNOUT(NLW_blk000002bf_MULTSIGNOUT_UNCONNECTED),
    .CEC(ce),
    .RSTM(sig00000002),
    .MULTSIGNIN(sig00000002),
    .CEB2(ce),
    .RSTCTRL(sig00000002),
    .CEP(ce),
    .CARRYCASCOUT(NLW_blk000002bf_CARRYCASCOUT_UNCONNECTED),
    .RSTA(sig00000002),
    .CECARRYIN(ce),
    .UNDERFLOW(NLW_blk000002bf_UNDERFLOW_UNCONNECTED),
    .RSTALUMODE(sig00000002),
    .RSTALLCARRYIN(sig00000002),
    .CEALUMODE(ce),
    .CEA2(ce),
    .CEA1(sig00000002),
    .RSTB(sig00000002),
    .CEMULTCARRYIN(sig00000002),
    .OVERFLOW(NLW_blk000002bf_OVERFLOW_UNCONNECTED),
    .CECTRL(ce),
    .CARRYCASCIN(sig00000002),
    .RSTP(sig00000002),
    .CARRYINSEL({sig00000002, sig00000002, sig00000002}),
    .OPMODE({sig00000002, sig000001a0, sig000001a0, sig00000002, sig000001a1, sig00000002, sig000001a1}),
    .ALUMODE({sig00000002, sig00000002, sig000001fb, sig000001fb}),
    .C({sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000188, sig00000189
, sig0000018a, sig0000018b, sig0000018c, sig0000018d, sig0000018e, sig0000018f, sig00000190, sig00000191, sig00000192, sig00000193, sig00000194,
sig00000195, sig00000196, sig00000197, sig00000198, sig00000199, sig0000019a, sig0000019b, sig0000019c, sig0000019d, sig0000019e, sig0000019f,
sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002,
sig00000002, sig00000002, sig00000002, sig00000002}),
    .B({sig00000002, sig00000002, sig00000178, sig00000179, sig0000017a, sig0000017b, sig0000017c, sig0000017d, sig0000017e, sig0000017f, sig00000180
, sig00000181, sig00000182, sig00000183, sig00000184, sig00000185, sig00000186, sig00000187}),
    .P({\NLW_blk000002bf_P<47>_UNCONNECTED , \NLW_blk000002bf_P<46>_UNCONNECTED , \NLW_blk000002bf_P<45>_UNCONNECTED ,
\NLW_blk000002bf_P<44>_UNCONNECTED , \NLW_blk000002bf_P<43>_UNCONNECTED , \NLW_blk000002bf_P<42>_UNCONNECTED , \NLW_blk000002bf_P<41>_UNCONNECTED ,
\NLW_blk000002bf_P<40>_UNCONNECTED , sig0000004a, sig0000004b, sig0000004c, sig0000004d, sig0000004e, sig0000004f, sig00000050, sig00000051,
sig00000052, sig00000053, sig00000054, sig00000055, sig00000056, sig00000057, sig00000058, sig00000059, sig0000005a, sig0000005b, sig0000005c,
sig0000005d, sig0000005e, sig0000005f, sig00000060, sig00000061, sig00000062, sig00000063, sig00000064, sig000001ea, sig000001eb, sig000001ec,
sig000001ed, sig000001ee, sig000001ef, sig000001f0, sig000001f1, sig000001f2, sig000001f3, sig000001f4, sig000001f5, sig000001f6}),
    .A({sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000160, sig00000161, sig00000162, sig00000163, sig00000164
, sig00000165, sig00000166, sig00000167, sig00000168, sig00000169, sig0000016a, sig0000016b, sig0000016c, sig0000016d, sig0000016e, sig0000016f,
sig00000170, sig00000171, sig00000172, sig00000173, sig00000174, sig00000175, sig00000176, sig00000177}),
    .ACOUT({\NLW_blk000002bf_ACOUT<29>_UNCONNECTED , \NLW_blk000002bf_ACOUT<28>_UNCONNECTED , \NLW_blk000002bf_ACOUT<27>_UNCONNECTED ,
\NLW_blk000002bf_ACOUT<26>_UNCONNECTED , \NLW_blk000002bf_ACOUT<25>_UNCONNECTED , \NLW_blk000002bf_ACOUT<24>_UNCONNECTED ,
\NLW_blk000002bf_ACOUT<23>_UNCONNECTED , \NLW_blk000002bf_ACOUT<22>_UNCONNECTED , \NLW_blk000002bf_ACOUT<21>_UNCONNECTED ,
\NLW_blk000002bf_ACOUT<20>_UNCONNECTED , \NLW_blk000002bf_ACOUT<19>_UNCONNECTED , \NLW_blk000002bf_ACOUT<18>_UNCONNECTED ,
\NLW_blk000002bf_ACOUT<17>_UNCONNECTED , \NLW_blk000002bf_ACOUT<16>_UNCONNECTED , \NLW_blk000002bf_ACOUT<15>_UNCONNECTED ,
\NLW_blk000002bf_ACOUT<14>_UNCONNECTED , \NLW_blk000002bf_ACOUT<13>_UNCONNECTED , \NLW_blk000002bf_ACOUT<12>_UNCONNECTED ,
\NLW_blk000002bf_ACOUT<11>_UNCONNECTED , \NLW_blk000002bf_ACOUT<10>_UNCONNECTED , \NLW_blk000002bf_ACOUT<9>_UNCONNECTED ,
\NLW_blk000002bf_ACOUT<8>_UNCONNECTED , \NLW_blk000002bf_ACOUT<7>_UNCONNECTED , \NLW_blk000002bf_ACOUT<6>_UNCONNECTED ,
\NLW_blk000002bf_ACOUT<5>_UNCONNECTED , \NLW_blk000002bf_ACOUT<4>_UNCONNECTED , \NLW_blk000002bf_ACOUT<3>_UNCONNECTED ,
\NLW_blk000002bf_ACOUT<2>_UNCONNECTED , \NLW_blk000002bf_ACOUT<1>_UNCONNECTED , \NLW_blk000002bf_ACOUT<0>_UNCONNECTED }),
    .PCIN({sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002,
sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002,
sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002,
sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002,
sig00000002, sig00000002, sig00000002, sig00000002, sig00000002}),
    .CARRYOUT({\NLW_blk000002bf_CARRYOUT<3>_UNCONNECTED , \NLW_blk000002bf_CARRYOUT<2>_UNCONNECTED , \NLW_blk000002bf_CARRYOUT<1>_UNCONNECTED ,
\NLW_blk000002bf_CARRYOUT<0>_UNCONNECTED }),
    .BCIN({sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002,
sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002}),
    .BCOUT({\NLW_blk000002bf_BCOUT<17>_UNCONNECTED , \NLW_blk000002bf_BCOUT<16>_UNCONNECTED , \NLW_blk000002bf_BCOUT<15>_UNCONNECTED ,
\NLW_blk000002bf_BCOUT<14>_UNCONNECTED , \NLW_blk000002bf_BCOUT<13>_UNCONNECTED , \NLW_blk000002bf_BCOUT<12>_UNCONNECTED ,
\NLW_blk000002bf_BCOUT<11>_UNCONNECTED , \NLW_blk000002bf_BCOUT<10>_UNCONNECTED , \NLW_blk000002bf_BCOUT<9>_UNCONNECTED ,
\NLW_blk000002bf_BCOUT<8>_UNCONNECTED , \NLW_blk000002bf_BCOUT<7>_UNCONNECTED , \NLW_blk000002bf_BCOUT<6>_UNCONNECTED ,
\NLW_blk000002bf_BCOUT<5>_UNCONNECTED , \NLW_blk000002bf_BCOUT<4>_UNCONNECTED , \NLW_blk000002bf_BCOUT<3>_UNCONNECTED ,
\NLW_blk000002bf_BCOUT<2>_UNCONNECTED , \NLW_blk000002bf_BCOUT<1>_UNCONNECTED , \NLW_blk000002bf_BCOUT<0>_UNCONNECTED }),
    .PCOUT({\NLW_blk000002bf_PCOUT<47>_UNCONNECTED , \NLW_blk000002bf_PCOUT<46>_UNCONNECTED , \NLW_blk000002bf_PCOUT<45>_UNCONNECTED ,
\NLW_blk000002bf_PCOUT<44>_UNCONNECTED , \NLW_blk000002bf_PCOUT<43>_UNCONNECTED , \NLW_blk000002bf_PCOUT<42>_UNCONNECTED ,
\NLW_blk000002bf_PCOUT<41>_UNCONNECTED , \NLW_blk000002bf_PCOUT<40>_UNCONNECTED , \NLW_blk000002bf_PCOUT<39>_UNCONNECTED ,
\NLW_blk000002bf_PCOUT<38>_UNCONNECTED , \NLW_blk000002bf_PCOUT<37>_UNCONNECTED , \NLW_blk000002bf_PCOUT<36>_UNCONNECTED ,
\NLW_blk000002bf_PCOUT<35>_UNCONNECTED , \NLW_blk000002bf_PCOUT<34>_UNCONNECTED , \NLW_blk000002bf_PCOUT<33>_UNCONNECTED ,
\NLW_blk000002bf_PCOUT<32>_UNCONNECTED , \NLW_blk000002bf_PCOUT<31>_UNCONNECTED , \NLW_blk000002bf_PCOUT<30>_UNCONNECTED ,
\NLW_blk000002bf_PCOUT<29>_UNCONNECTED , \NLW_blk000002bf_PCOUT<28>_UNCONNECTED , \NLW_blk000002bf_PCOUT<27>_UNCONNECTED ,
\NLW_blk000002bf_PCOUT<26>_UNCONNECTED , \NLW_blk000002bf_PCOUT<25>_UNCONNECTED , \NLW_blk000002bf_PCOUT<24>_UNCONNECTED ,
\NLW_blk000002bf_PCOUT<23>_UNCONNECTED , \NLW_blk000002bf_PCOUT<22>_UNCONNECTED , \NLW_blk000002bf_PCOUT<21>_UNCONNECTED ,
\NLW_blk000002bf_PCOUT<20>_UNCONNECTED , \NLW_blk000002bf_PCOUT<19>_UNCONNECTED , \NLW_blk000002bf_PCOUT<18>_UNCONNECTED ,
\NLW_blk000002bf_PCOUT<17>_UNCONNECTED , \NLW_blk000002bf_PCOUT<16>_UNCONNECTED , \NLW_blk000002bf_PCOUT<15>_UNCONNECTED ,
\NLW_blk000002bf_PCOUT<14>_UNCONNECTED , \NLW_blk000002bf_PCOUT<13>_UNCONNECTED , \NLW_blk000002bf_PCOUT<12>_UNCONNECTED ,
\NLW_blk000002bf_PCOUT<11>_UNCONNECTED , \NLW_blk000002bf_PCOUT<10>_UNCONNECTED , \NLW_blk000002bf_PCOUT<9>_UNCONNECTED ,
\NLW_blk000002bf_PCOUT<8>_UNCONNECTED , \NLW_blk000002bf_PCOUT<7>_UNCONNECTED , \NLW_blk000002bf_PCOUT<6>_UNCONNECTED ,
\NLW_blk000002bf_PCOUT<5>_UNCONNECTED , \NLW_blk000002bf_PCOUT<4>_UNCONNECTED , \NLW_blk000002bf_PCOUT<3>_UNCONNECTED ,
\NLW_blk000002bf_PCOUT<2>_UNCONNECTED , \NLW_blk000002bf_PCOUT<1>_UNCONNECTED , \NLW_blk000002bf_PCOUT<0>_UNCONNECTED }),
    .ACIN({sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002,
sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002,
sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002})
  );
  DSP48E #(
    .ACASCREG ( 2 ),
    .ALUMODEREG ( 1 ),
    .AREG ( 2 ),
    .AUTORESET_PATTERN_DETECT ( 0 ),
    .AUTORESET_PATTERN_DETECT_OPTINV ( "MATCH" ),
    .A_INPUT ( "DIRECT" ),
    .BCASCREG ( 1 ),
    .BREG ( 1 ),
    .B_INPUT ( "DIRECT" ),
    .CARRYINREG ( 1 ),
    .CARRYINSELREG ( 1 ),
    .CREG ( 1 ),
    .MASK ( 48'h3FFFFFFFFFFF ),
    .MREG ( 1 ),
    .MULTCARRYINREG ( 0 ),
    .OPMODEREG ( 1 ),
    .PATTERN ( 48'h000000000000 ),
    .PREG ( 1 ),
    .SEL_MASK ( "MASK" ),
    .SEL_PATTERN ( "PATTERN" ),
    .SEL_ROUNDING_MASK ( "SEL_MASK" ),
    .SIM_MODE ( "SAFE" ),
    .USE_MULT ( "MULT_S" ),
    .USE_PATTERN_DETECT ( "NO_PATDET" ),
    .USE_SIMD ( "ONE48" ))
  blk000002c0 (
    .CEM(ce),
    .CLK(clk),
    .PATTERNBDETECT(NLW_blk000002c0_PATTERNBDETECT_UNCONNECTED),
    .RSTC(sig00000002),
    .CEB1(sig00000002),
    .MULTSIGNOUT(NLW_blk000002c0_MULTSIGNOUT_UNCONNECTED),
    .CEC(ce),
    .RSTM(sig00000002),
    .MULTSIGNIN(sig00000002),
    .CEB2(ce),
    .RSTCTRL(sig00000002),
    .CEP(ce),
    .CARRYCASCOUT(NLW_blk000002c0_CARRYCASCOUT_UNCONNECTED),
    .RSTA(sig00000002),
    .CECARRYIN(ce),
    .UNDERFLOW(NLW_blk000002c0_UNDERFLOW_UNCONNECTED),
    .PATTERNDETECT(NLW_blk000002c0_PATTERNDETECT_UNCONNECTED),
    .RSTALUMODE(sig00000002),
    .RSTALLCARRYIN(sig00000002),
    .CEALUMODE(ce),
    .CEA2(ce),
    .CEA1(ce),
    .RSTB(sig00000002),
    .CEMULTCARRYIN(sig00000002),
    .OVERFLOW(NLW_blk000002c0_OVERFLOW_UNCONNECTED),
    .CECTRL(ce),
    .CARRYIN(sig00000002),
    .CARRYCASCIN(sig00000002),
    .RSTP(sig00000002),
    .CARRYINSEL({sig00000002, sig00000002, sig00000002}),
    .C({sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002
, sig00000002, sig00000002, sig00000011, sig00000012, sig00000013, sig00000014, sig00000015, sig00000016, sig00000017, sig00000018, sig00000001,
sig0000022b, sig0000022a, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002,
sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002,
sig00000002, sig0000022c, sig00000002, sig00000002}),
    .B({sig00000002, sig00000002, sig0000025b, sig0000025a, sig00000259, sig00000258, sig00000257, sig00000256, sig00000255, sig00000254, sig00000253
, sig00000252, sig00000251, sig00000250, sig0000024f, sig0000024e, sig0000024d, sig0000024c}),
    .P({\NLW_blk000002c0_P<47>_UNCONNECTED , \NLW_blk000002c0_P<46>_UNCONNECTED , \NLW_blk000002c0_P<45>_UNCONNECTED ,
\NLW_blk000002c0_P<44>_UNCONNECTED , \NLW_blk000002c0_P<43>_UNCONNECTED , \NLW_blk000002c0_P<42>_UNCONNECTED , \NLW_blk000002c0_P<41>_UNCONNECTED ,
\NLW_blk000002c0_P<40>_UNCONNECTED , \NLW_blk000002c0_P<39>_UNCONNECTED , \NLW_blk000002c0_P<38>_UNCONNECTED , \NLW_blk000002c0_P<37>_UNCONNECTED ,
\NLW_blk000002c0_P<36>_UNCONNECTED , \NLW_blk000002c0_P<35>_UNCONNECTED , sig00000083, sig00000084, sig00000085, sig00000086, sig00000087, sig00000088
, sig00000089, sig0000008a, \NLW_blk000002c0_P<26>_UNCONNECTED , \NLW_blk000002c0_P<25>_UNCONNECTED , sig0000006c, sig0000006d, sig0000006e,
sig0000006f, sig00000070, sig00000071, sig00000072, sig00000073, sig00000074, sig00000075, sig00000076, sig00000077, sig00000078, sig00000079,
sig0000007a, sig0000007b, sig0000007c, sig0000007d, sig0000007e, sig0000007f, sig00000080, sig00000081, sig00000082,
\NLW_blk000002c0_P<1>_UNCONNECTED , \NLW_blk000002c0_P<0>_UNCONNECTED }),
    .A({sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000249, sig00000248, sig00000247, sig00000246, sig00000245
, sig00000244, sig00000243, sig00000242, sig00000241, sig00000240, sig0000023f, sig0000023e, sig0000023d, sig0000023c, sig0000023b, sig0000023a,
sig00000239, sig00000238, sig00000237, sig00000236, sig00000235, sig00000234, sig00000233, sig00000232}),
    .ACOUT({\NLW_blk000002c0_ACOUT<29>_UNCONNECTED , \NLW_blk000002c0_ACOUT<28>_UNCONNECTED , \NLW_blk000002c0_ACOUT<27>_UNCONNECTED ,
\NLW_blk000002c0_ACOUT<26>_UNCONNECTED , \NLW_blk000002c0_ACOUT<25>_UNCONNECTED , \NLW_blk000002c0_ACOUT<24>_UNCONNECTED ,
\NLW_blk000002c0_ACOUT<23>_UNCONNECTED , \NLW_blk000002c0_ACOUT<22>_UNCONNECTED , \NLW_blk000002c0_ACOUT<21>_UNCONNECTED ,
\NLW_blk000002c0_ACOUT<20>_UNCONNECTED , \NLW_blk000002c0_ACOUT<19>_UNCONNECTED , \NLW_blk000002c0_ACOUT<18>_UNCONNECTED ,
\NLW_blk000002c0_ACOUT<17>_UNCONNECTED , \NLW_blk000002c0_ACOUT<16>_UNCONNECTED , \NLW_blk000002c0_ACOUT<15>_UNCONNECTED ,
\NLW_blk000002c0_ACOUT<14>_UNCONNECTED , \NLW_blk000002c0_ACOUT<13>_UNCONNECTED , \NLW_blk000002c0_ACOUT<12>_UNCONNECTED ,
\NLW_blk000002c0_ACOUT<11>_UNCONNECTED , \NLW_blk000002c0_ACOUT<10>_UNCONNECTED , \NLW_blk000002c0_ACOUT<9>_UNCONNECTED ,
\NLW_blk000002c0_ACOUT<8>_UNCONNECTED , \NLW_blk000002c0_ACOUT<7>_UNCONNECTED , \NLW_blk000002c0_ACOUT<6>_UNCONNECTED ,
\NLW_blk000002c0_ACOUT<5>_UNCONNECTED , \NLW_blk000002c0_ACOUT<4>_UNCONNECTED , \NLW_blk000002c0_ACOUT<3>_UNCONNECTED ,
\NLW_blk000002c0_ACOUT<2>_UNCONNECTED , \NLW_blk000002c0_ACOUT<1>_UNCONNECTED , \NLW_blk000002c0_ACOUT<0>_UNCONNECTED }),
    .OPMODE({sig00000002, sig00000001, sig00000001, sig00000002, sig00000001, sig00000002, sig00000001}),
    .PCIN({sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002,
sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002,
sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002,
sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002,
sig00000002, sig00000002, sig00000002, sig00000002, sig00000002}),
    .ALUMODE({sig00000002, sig00000002, sig00000002, sig00000002}),
    .CARRYOUT({\NLW_blk000002c0_CARRYOUT<3>_UNCONNECTED , \NLW_blk000002c0_CARRYOUT<2>_UNCONNECTED , \NLW_blk000002c0_CARRYOUT<1>_UNCONNECTED ,
\NLW_blk000002c0_CARRYOUT<0>_UNCONNECTED }),
    .BCIN({sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002,
sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002}),
    .BCOUT({\NLW_blk000002c0_BCOUT<17>_UNCONNECTED , \NLW_blk000002c0_BCOUT<16>_UNCONNECTED , \NLW_blk000002c0_BCOUT<15>_UNCONNECTED ,
\NLW_blk000002c0_BCOUT<14>_UNCONNECTED , \NLW_blk000002c0_BCOUT<13>_UNCONNECTED , \NLW_blk000002c0_BCOUT<12>_UNCONNECTED ,
\NLW_blk000002c0_BCOUT<11>_UNCONNECTED , \NLW_blk000002c0_BCOUT<10>_UNCONNECTED , \NLW_blk000002c0_BCOUT<9>_UNCONNECTED ,
\NLW_blk000002c0_BCOUT<8>_UNCONNECTED , \NLW_blk000002c0_BCOUT<7>_UNCONNECTED , \NLW_blk000002c0_BCOUT<6>_UNCONNECTED ,
\NLW_blk000002c0_BCOUT<5>_UNCONNECTED , \NLW_blk000002c0_BCOUT<4>_UNCONNECTED , \NLW_blk000002c0_BCOUT<3>_UNCONNECTED ,
\NLW_blk000002c0_BCOUT<2>_UNCONNECTED , \NLW_blk000002c0_BCOUT<1>_UNCONNECTED , \NLW_blk000002c0_BCOUT<0>_UNCONNECTED }),
    .PCOUT({\NLW_blk000002c0_PCOUT<47>_UNCONNECTED , \NLW_blk000002c0_PCOUT<46>_UNCONNECTED , \NLW_blk000002c0_PCOUT<45>_UNCONNECTED ,
\NLW_blk000002c0_PCOUT<44>_UNCONNECTED , \NLW_blk000002c0_PCOUT<43>_UNCONNECTED , \NLW_blk000002c0_PCOUT<42>_UNCONNECTED ,
\NLW_blk000002c0_PCOUT<41>_UNCONNECTED , \NLW_blk000002c0_PCOUT<40>_UNCONNECTED , \NLW_blk000002c0_PCOUT<39>_UNCONNECTED ,
\NLW_blk000002c0_PCOUT<38>_UNCONNECTED , \NLW_blk000002c0_PCOUT<37>_UNCONNECTED , \NLW_blk000002c0_PCOUT<36>_UNCONNECTED ,
\NLW_blk000002c0_PCOUT<35>_UNCONNECTED , \NLW_blk000002c0_PCOUT<34>_UNCONNECTED , \NLW_blk000002c0_PCOUT<33>_UNCONNECTED ,
\NLW_blk000002c0_PCOUT<32>_UNCONNECTED , \NLW_blk000002c0_PCOUT<31>_UNCONNECTED , \NLW_blk000002c0_PCOUT<30>_UNCONNECTED ,
\NLW_blk000002c0_PCOUT<29>_UNCONNECTED , \NLW_blk000002c0_PCOUT<28>_UNCONNECTED , \NLW_blk000002c0_PCOUT<27>_UNCONNECTED ,
\NLW_blk000002c0_PCOUT<26>_UNCONNECTED , \NLW_blk000002c0_PCOUT<25>_UNCONNECTED , \NLW_blk000002c0_PCOUT<24>_UNCONNECTED ,
\NLW_blk000002c0_PCOUT<23>_UNCONNECTED , \NLW_blk000002c0_PCOUT<22>_UNCONNECTED , \NLW_blk000002c0_PCOUT<21>_UNCONNECTED ,
\NLW_blk000002c0_PCOUT<20>_UNCONNECTED , \NLW_blk000002c0_PCOUT<19>_UNCONNECTED , \NLW_blk000002c0_PCOUT<18>_UNCONNECTED ,
\NLW_blk000002c0_PCOUT<17>_UNCONNECTED , \NLW_blk000002c0_PCOUT<16>_UNCONNECTED , \NLW_blk000002c0_PCOUT<15>_UNCONNECTED ,
\NLW_blk000002c0_PCOUT<14>_UNCONNECTED , \NLW_blk000002c0_PCOUT<13>_UNCONNECTED , \NLW_blk000002c0_PCOUT<12>_UNCONNECTED ,
\NLW_blk000002c0_PCOUT<11>_UNCONNECTED , \NLW_blk000002c0_PCOUT<10>_UNCONNECTED , \NLW_blk000002c0_PCOUT<9>_UNCONNECTED ,
\NLW_blk000002c0_PCOUT<8>_UNCONNECTED , \NLW_blk000002c0_PCOUT<7>_UNCONNECTED , \NLW_blk000002c0_PCOUT<6>_UNCONNECTED ,
\NLW_blk000002c0_PCOUT<5>_UNCONNECTED , \NLW_blk000002c0_PCOUT<4>_UNCONNECTED , \NLW_blk000002c0_PCOUT<3>_UNCONNECTED ,
\NLW_blk000002c0_PCOUT<2>_UNCONNECTED , \NLW_blk000002c0_PCOUT<1>_UNCONNECTED , \NLW_blk000002c0_PCOUT<0>_UNCONNECTED }),
    .ACIN({sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002,
sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002,
sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002})
  );
endmodule