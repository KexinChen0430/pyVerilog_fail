module div (
  aclk, s_axis_divisor_tvalid, s_axis_dividend_tvalid, s_axis_divisor_tready, s_axis_dividend_tready, m_axis_dout_tvalid, s_axis_divisor_tdata,
s_axis_dividend_tdata, m_axis_dout_tdata
)/* synthesis syn_black_box syn_noprune=1 */;
  input aclk;
  input s_axis_divisor_tvalid;
  input s_axis_dividend_tvalid;
  output s_axis_divisor_tready;
  output s_axis_dividend_tready;
  output m_axis_dout_tvalid;
  input [15 : 0] s_axis_divisor_tdata;
  input [15 : 0] s_axis_dividend_tdata;
  output [31 : 0] m_axis_dout_tdata;
  // synthesis translate_off
  wire NlwRenamedSignal_s_axis_dividend_tready;
  wire \blk00000001/sig000005f5 ;
  wire \blk00000001/sig000005f4 ;
  wire \blk00000001/sig000005f3 ;
  wire \blk00000001/sig000005f2 ;
  wire \blk00000001/sig000005f1 ;
  wire \blk00000001/sig000005f0 ;
  wire \blk00000001/sig000005ef ;
  wire \blk00000001/sig000005ee ;
  wire \blk00000001/sig000005ed ;
  wire \blk00000001/sig000005ec ;
  wire \blk00000001/sig000005eb ;
  wire \blk00000001/sig000005ea ;
  wire \blk00000001/sig000005e9 ;
  wire \blk00000001/sig000005e8 ;
  wire \blk00000001/sig000005e7 ;
  wire \blk00000001/sig000005e6 ;
  wire \blk00000001/sig000005e5 ;
  wire \blk00000001/sig000005e4 ;
  wire \blk00000001/sig000005e3 ;
  wire \blk00000001/sig000005e2 ;
  wire \blk00000001/sig000005e1 ;
  wire \blk00000001/sig000005e0 ;
  wire \blk00000001/sig000005df ;
  wire \blk00000001/sig000005de ;
  wire \blk00000001/sig000005dd ;
  wire \blk00000001/sig000005dc ;
  wire \blk00000001/sig000005db ;
  wire \blk00000001/sig000005da ;
  wire \blk00000001/sig000005d9 ;
  wire \blk00000001/sig000005d8 ;
  wire \blk00000001/sig000005d7 ;
  wire \blk00000001/sig000005d6 ;
  wire \blk00000001/sig000005d5 ;
  wire \blk00000001/sig000005d4 ;
  wire \blk00000001/sig000005d3 ;
  wire \blk00000001/sig000005d2 ;
  wire \blk00000001/sig000005d1 ;
  wire \blk00000001/sig000005d0 ;
  wire \blk00000001/sig000005cf ;
  wire \blk00000001/sig000005ce ;
  wire \blk00000001/sig000005cd ;
  wire \blk00000001/sig000005cc ;
  wire \blk00000001/sig000005cb ;
  wire \blk00000001/sig000005ca ;
  wire \blk00000001/sig000005c9 ;
  wire \blk00000001/sig000005c8 ;
  wire \blk00000001/sig000005c7 ;
  wire \blk00000001/sig000005c6 ;
  wire \blk00000001/sig000005c5 ;
  wire \blk00000001/sig000005c4 ;
  wire \blk00000001/sig000005c3 ;
  wire \blk00000001/sig000005c2 ;
  wire \blk00000001/sig000005c1 ;
  wire \blk00000001/sig000005c0 ;
  wire \blk00000001/sig000005bf ;
  wire \blk00000001/sig000005be ;
  wire \blk00000001/sig000005bd ;
  wire \blk00000001/sig000005bc ;
  wire \blk00000001/sig000005bb ;
  wire \blk00000001/sig000005ba ;
  wire \blk00000001/sig000005b9 ;
  wire \blk00000001/sig000005b8 ;
  wire \blk00000001/sig000005b7 ;
  wire \blk00000001/sig000005b6 ;
  wire \blk00000001/sig000005b5 ;
  wire \blk00000001/sig000005b4 ;
  wire \blk00000001/sig000005b3 ;
  wire \blk00000001/sig000005b2 ;
  wire \blk00000001/sig000005b1 ;
  wire \blk00000001/sig000005b0 ;
  wire \blk00000001/sig000005af ;
  wire \blk00000001/sig000005ae ;
  wire \blk00000001/sig000005ad ;
  wire \blk00000001/sig000005ac ;
  wire \blk00000001/sig000005ab ;
  wire \blk00000001/sig000005aa ;
  wire \blk00000001/sig000005a9 ;
  wire \blk00000001/sig000005a8 ;
  wire \blk00000001/sig000005a7 ;
  wire \blk00000001/sig000005a6 ;
  wire \blk00000001/sig000005a5 ;
  wire \blk00000001/sig000005a4 ;
  wire \blk00000001/sig000005a3 ;
  wire \blk00000001/sig000005a2 ;
  wire \blk00000001/sig000005a1 ;
  wire \blk00000001/sig000005a0 ;
  wire \blk00000001/sig0000059f ;
  wire \blk00000001/sig0000059e ;
  wire \blk00000001/sig0000059d ;
  wire \blk00000001/sig0000059c ;
  wire \blk00000001/sig0000059b ;
  wire \blk00000001/sig0000059a ;
  wire \blk00000001/sig00000599 ;
  wire \blk00000001/sig00000598 ;
  wire \blk00000001/sig00000597 ;
  wire \blk00000001/sig00000596 ;
  wire \blk00000001/sig00000595 ;
  wire \blk00000001/sig00000594 ;
  wire \blk00000001/sig00000593 ;
  wire \blk00000001/sig00000592 ;
  wire \blk00000001/sig00000591 ;
  wire \blk00000001/sig00000590 ;
  wire \blk00000001/sig0000058f ;
  wire \blk00000001/sig0000058e ;
  wire \blk00000001/sig0000058d ;
  wire \blk00000001/sig0000058c ;
  wire \blk00000001/sig0000058b ;
  wire \blk00000001/sig0000058a ;
  wire \blk00000001/sig00000589 ;
  wire \blk00000001/sig00000588 ;
  wire \blk00000001/sig00000587 ;
  wire \blk00000001/sig00000586 ;
  wire \blk00000001/sig00000585 ;
  wire \blk00000001/sig00000584 ;
  wire \blk00000001/sig00000583 ;
  wire \blk00000001/sig00000582 ;
  wire \blk00000001/sig00000581 ;
  wire \blk00000001/sig00000580 ;
  wire \blk00000001/sig0000057f ;
  wire \blk00000001/sig0000057e ;
  wire \blk00000001/sig0000057d ;
  wire \blk00000001/sig0000057c ;
  wire \blk00000001/sig0000057b ;
  wire \blk00000001/sig0000057a ;
  wire \blk00000001/sig00000579 ;
  wire \blk00000001/sig00000578 ;
  wire \blk00000001/sig00000577 ;
  wire \blk00000001/sig00000576 ;
  wire \blk00000001/sig00000575 ;
  wire \blk00000001/sig00000574 ;
  wire \blk00000001/sig00000573 ;
  wire \blk00000001/sig00000572 ;
  wire \blk00000001/sig00000571 ;
  wire \blk00000001/sig00000570 ;
  wire \blk00000001/sig0000056f ;
  wire \blk00000001/sig0000056e ;
  wire \blk00000001/sig0000056d ;
  wire \blk00000001/sig0000056c ;
  wire \blk00000001/sig0000056b ;
  wire \blk00000001/sig0000056a ;
  wire \blk00000001/sig00000569 ;
  wire \blk00000001/sig00000568 ;
  wire \blk00000001/sig00000567 ;
  wire \blk00000001/sig00000566 ;
  wire \blk00000001/sig00000565 ;
  wire \blk00000001/sig00000564 ;
  wire \blk00000001/sig00000563 ;
  wire \blk00000001/sig00000562 ;
  wire \blk00000001/sig00000561 ;
  wire \blk00000001/sig00000560 ;
  wire \blk00000001/sig0000055f ;
  wire \blk00000001/sig0000055e ;
  wire \blk00000001/sig0000055d ;
  wire \blk00000001/sig0000055c ;
  wire \blk00000001/sig0000055b ;
  wire \blk00000001/sig0000055a ;
  wire \blk00000001/sig00000559 ;
  wire \blk00000001/sig00000558 ;
  wire \blk00000001/sig00000557 ;
  wire \blk00000001/sig00000556 ;
  wire \blk00000001/sig00000555 ;
  wire \blk00000001/sig00000554 ;
  wire \blk00000001/sig00000553 ;
  wire \blk00000001/sig00000552 ;
  wire \blk00000001/sig00000551 ;
  wire \blk00000001/sig00000550 ;
  wire \blk00000001/sig0000054f ;
  wire \blk00000001/sig0000054e ;
  wire \blk00000001/sig0000054d ;
  wire \blk00000001/sig0000054c ;
  wire \blk00000001/sig0000054b ;
  wire \blk00000001/sig0000054a ;
  wire \blk00000001/sig00000549 ;
  wire \blk00000001/sig00000548 ;
  wire \blk00000001/sig00000547 ;
  wire \blk00000001/sig00000546 ;
  wire \blk00000001/sig00000545 ;
  wire \blk00000001/sig00000544 ;
  wire \blk00000001/sig00000543 ;
  wire \blk00000001/sig00000542 ;
  wire \blk00000001/sig00000541 ;
  wire \blk00000001/sig00000540 ;
  wire \blk00000001/sig0000053f ;
  wire \blk00000001/sig0000053e ;
  wire \blk00000001/sig0000053d ;
  wire \blk00000001/sig0000053c ;
  wire \blk00000001/sig0000053b ;
  wire \blk00000001/sig0000053a ;
  wire \blk00000001/sig00000539 ;
  wire \blk00000001/sig00000538 ;
  wire \blk00000001/sig00000537 ;
  wire \blk00000001/sig00000536 ;
  wire \blk00000001/sig00000535 ;
  wire \blk00000001/sig00000534 ;
  wire \blk00000001/sig00000533 ;
  wire \blk00000001/sig00000532 ;
  wire \blk00000001/sig00000531 ;
  wire \blk00000001/sig00000530 ;
  wire \blk00000001/sig0000052f ;
  wire \blk00000001/sig0000052e ;
  wire \blk00000001/sig0000052d ;
  wire \blk00000001/sig0000052c ;
  wire \blk00000001/sig0000052b ;
  wire \blk00000001/sig0000052a ;
  wire \blk00000001/sig00000529 ;
  wire \blk00000001/sig00000528 ;
  wire \blk00000001/sig00000527 ;
  wire \blk00000001/sig00000526 ;
  wire \blk00000001/sig00000525 ;
  wire \blk00000001/sig00000524 ;
  wire \blk00000001/sig00000523 ;
  wire \blk00000001/sig00000522 ;
  wire \blk00000001/sig00000521 ;
  wire \blk00000001/sig00000520 ;
  wire \blk00000001/sig0000051f ;
  wire \blk00000001/sig0000051e ;
  wire \blk00000001/sig0000051d ;
  wire \blk00000001/sig0000051c ;
  wire \blk00000001/sig0000051b ;
  wire \blk00000001/sig0000051a ;
  wire \blk00000001/sig00000519 ;
  wire \blk00000001/sig00000518 ;
  wire \blk00000001/sig00000517 ;
  wire \blk00000001/sig00000516 ;
  wire \blk00000001/sig00000515 ;
  wire \blk00000001/sig00000514 ;
  wire \blk00000001/sig00000513 ;
  wire \blk00000001/sig00000512 ;
  wire \blk00000001/sig00000511 ;
  wire \blk00000001/sig00000510 ;
  wire \blk00000001/sig0000050f ;
  wire \blk00000001/sig0000050e ;
  wire \blk00000001/sig0000050d ;
  wire \blk00000001/sig0000050c ;
  wire \blk00000001/sig0000050b ;
  wire \blk00000001/sig0000050a ;
  wire \blk00000001/sig00000509 ;
  wire \blk00000001/sig00000508 ;
  wire \blk00000001/sig00000507 ;
  wire \blk00000001/sig00000506 ;
  wire \blk00000001/sig00000505 ;
  wire \blk00000001/sig00000504 ;
  wire \blk00000001/sig00000503 ;
  wire \blk00000001/sig00000502 ;
  wire \blk00000001/sig00000501 ;
  wire \blk00000001/sig00000500 ;
  wire \blk00000001/sig000004ff ;
  wire \blk00000001/sig000004fe ;
  wire \blk00000001/sig000004fd ;
  wire \blk00000001/sig000004fc ;
  wire \blk00000001/sig000004fb ;
  wire \blk00000001/sig000004fa ;
  wire \blk00000001/sig000004f9 ;
  wire \blk00000001/sig000004f8 ;
  wire \blk00000001/sig000004f7 ;
  wire \blk00000001/sig000004f6 ;
  wire \blk00000001/sig000004f5 ;
  wire \blk00000001/sig000004f4 ;
  wire \blk00000001/sig000004f3 ;
  wire \blk00000001/sig000004f2 ;
  wire \blk00000001/sig000004f1 ;
  wire \blk00000001/sig000004f0 ;
  wire \blk00000001/sig000004ef ;
  wire \blk00000001/sig000004ee ;
  wire \blk00000001/sig000004ed ;
  wire \blk00000001/sig000004ec ;
  wire \blk00000001/sig000004eb ;
  wire \blk00000001/sig000004ea ;
  wire \blk00000001/sig000004e9 ;
  wire \blk00000001/sig000004e8 ;
  wire \blk00000001/sig000004e7 ;
  wire \blk00000001/sig000004e6 ;
  wire \blk00000001/sig000004e5 ;
  wire \blk00000001/sig000004e4 ;
  wire \blk00000001/sig000004e3 ;
  wire \blk00000001/sig000004e2 ;
  wire \blk00000001/sig000004e1 ;
  wire \blk00000001/sig000004e0 ;
  wire \blk00000001/sig000004df ;
  wire \blk00000001/sig000004de ;
  wire \blk00000001/sig000004dd ;
  wire \blk00000001/sig000004dc ;
  wire \blk00000001/sig000004db ;
  wire \blk00000001/sig000004da ;
  wire \blk00000001/sig000004d9 ;
  wire \blk00000001/sig000004d8 ;
  wire \blk00000001/sig000004d7 ;
  wire \blk00000001/sig000004d6 ;
  wire \blk00000001/sig000004d5 ;
  wire \blk00000001/sig000004d4 ;
  wire \blk00000001/sig000004d3 ;
  wire \blk00000001/sig000004d2 ;
  wire \blk00000001/sig000004d1 ;
  wire \blk00000001/sig000004d0 ;
  wire \blk00000001/sig000004cf ;
  wire \blk00000001/sig000004ce ;
  wire \blk00000001/sig000004cd ;
  wire \blk00000001/sig000004cc ;
  wire \blk00000001/sig000004cb ;
  wire \blk00000001/sig000004ca ;
  wire \blk00000001/sig000004c9 ;
  wire \blk00000001/sig000004c8 ;
  wire \blk00000001/sig000004c7 ;
  wire \blk00000001/sig000004c6 ;
  wire \blk00000001/sig000004c5 ;
  wire \blk00000001/sig000004c4 ;
  wire \blk00000001/sig000004c3 ;
  wire \blk00000001/sig000004c2 ;
  wire \blk00000001/sig000004c1 ;
  wire \blk00000001/sig000004c0 ;
  wire \blk00000001/sig000004bf ;
  wire \blk00000001/sig000004be ;
  wire \blk00000001/sig000004bd ;
  wire \blk00000001/sig000004bc ;
  wire \blk00000001/sig000004bb ;
  wire \blk00000001/sig000004ba ;
  wire \blk00000001/sig000004b9 ;
  wire \blk00000001/sig000004b8 ;
  wire \blk00000001/sig000004b7 ;
  wire \blk00000001/sig000004b6 ;
  wire \blk00000001/sig000004b5 ;
  wire \blk00000001/sig000004b4 ;
  wire \blk00000001/sig000004b3 ;
  wire \blk00000001/sig000004b2 ;
  wire \blk00000001/sig000004b1 ;
  wire \blk00000001/sig000004b0 ;
  wire \blk00000001/sig000004af ;
  wire \blk00000001/sig000004ae ;
  wire \blk00000001/sig000004ad ;
  wire \blk00000001/sig000004ac ;
  wire \blk00000001/sig000004ab ;
  wire \blk00000001/sig000004aa ;
  wire \blk00000001/sig000004a9 ;
  wire \blk00000001/sig000004a8 ;
  wire \blk00000001/sig000004a7 ;
  wire \blk00000001/sig000004a6 ;
  wire \blk00000001/sig000004a5 ;
  wire \blk00000001/sig000004a4 ;
  wire \blk00000001/sig000004a3 ;
  wire \blk00000001/sig000004a2 ;
  wire \blk00000001/sig000004a1 ;
  wire \blk00000001/sig000004a0 ;
  wire \blk00000001/sig0000049f ;
  wire \blk00000001/sig0000049e ;
  wire \blk00000001/sig0000049d ;
  wire \blk00000001/sig0000049c ;
  wire \blk00000001/sig0000049b ;
  wire \blk00000001/sig0000049a ;
  wire \blk00000001/sig00000499 ;
  wire \blk00000001/sig00000498 ;
  wire \blk00000001/sig00000497 ;
  wire \blk00000001/sig00000496 ;
  wire \blk00000001/sig00000495 ;
  wire \blk00000001/sig00000494 ;
  wire \blk00000001/sig00000493 ;
  wire \blk00000001/sig00000492 ;
  wire \blk00000001/sig00000491 ;
  wire \blk00000001/sig00000490 ;
  wire \blk00000001/sig0000048f ;
  wire \blk00000001/sig0000048e ;
  wire \blk00000001/sig0000048d ;
  wire \blk00000001/sig0000048c ;
  wire \blk00000001/sig0000048b ;
  wire \blk00000001/sig0000048a ;
  wire \blk00000001/sig00000489 ;
  wire \blk00000001/sig00000488 ;
  wire \blk00000001/sig00000487 ;
  wire \blk00000001/sig00000486 ;
  wire \blk00000001/sig00000485 ;
  wire \blk00000001/sig00000484 ;
  wire \blk00000001/sig00000483 ;
  wire \blk00000001/sig00000482 ;
  wire \blk00000001/sig00000481 ;
  wire \blk00000001/sig00000480 ;
  wire \blk00000001/sig0000047f ;
  wire \blk00000001/sig0000047e ;
  wire \blk00000001/sig0000047d ;
  wire \blk00000001/sig0000047c ;
  wire \blk00000001/sig0000047b ;
  wire \blk00000001/sig0000047a ;
  wire \blk00000001/sig00000479 ;
  wire \blk00000001/sig00000478 ;
  wire \blk00000001/sig00000477 ;
  wire \blk00000001/sig00000476 ;
  wire \blk00000001/sig00000475 ;
  wire \blk00000001/sig00000474 ;
  wire \blk00000001/sig00000473 ;
  wire \blk00000001/sig00000472 ;
  wire \blk00000001/sig00000471 ;
  wire \blk00000001/sig00000470 ;
  wire \blk00000001/sig0000046f ;
  wire \blk00000001/sig0000046e ;
  wire \blk00000001/sig0000046d ;
  wire \blk00000001/sig0000046c ;
  wire \blk00000001/sig0000046b ;
  wire \blk00000001/sig0000046a ;
  wire \blk00000001/sig00000469 ;
  wire \blk00000001/sig00000468 ;
  wire \blk00000001/sig00000467 ;
  wire \blk00000001/sig00000466 ;
  wire \blk00000001/sig00000465 ;
  wire \blk00000001/sig00000464 ;
  wire \blk00000001/sig00000463 ;
  wire \blk00000001/sig00000462 ;
  wire \blk00000001/sig00000461 ;
  wire \blk00000001/sig00000460 ;
  wire \blk00000001/sig0000045f ;
  wire \blk00000001/sig0000045e ;
  wire \blk00000001/sig0000045d ;
  wire \blk00000001/sig0000045c ;
  wire \blk00000001/sig0000045b ;
  wire \blk00000001/sig0000045a ;
  wire \blk00000001/sig00000459 ;
  wire \blk00000001/sig00000458 ;
  wire \blk00000001/sig00000457 ;
  wire \blk00000001/sig00000456 ;
  wire \blk00000001/sig00000455 ;
  wire \blk00000001/sig00000454 ;
  wire \blk00000001/sig00000453 ;
  wire \blk00000001/sig00000452 ;
  wire \blk00000001/sig00000451 ;
  wire \blk00000001/sig00000450 ;
  wire \blk00000001/sig0000044f ;
  wire \blk00000001/sig0000044e ;
  wire \blk00000001/sig0000044d ;
  wire \blk00000001/sig0000044c ;
  wire \blk00000001/sig0000044b ;
  wire \blk00000001/sig0000044a ;
  wire \blk00000001/sig00000449 ;
  wire \blk00000001/sig00000448 ;
  wire \blk00000001/sig00000447 ;
  wire \blk00000001/sig00000446 ;
  wire \blk00000001/sig00000445 ;
  wire \blk00000001/sig00000444 ;
  wire \blk00000001/sig00000443 ;
  wire \blk00000001/sig00000442 ;
  wire \blk00000001/sig00000441 ;
  wire \blk00000001/sig00000440 ;
  wire \blk00000001/sig0000043f ;
  wire \blk00000001/sig0000043e ;
  wire \blk00000001/sig0000043d ;
  wire \blk00000001/sig0000043c ;
  wire \blk00000001/sig0000043b ;
  wire \blk00000001/sig0000043a ;
  wire \blk00000001/sig00000439 ;
  wire \blk00000001/sig00000438 ;
  wire \blk00000001/sig00000437 ;
  wire \blk00000001/sig00000436 ;
  wire \blk00000001/sig00000435 ;
  wire \blk00000001/sig00000434 ;
  wire \blk00000001/sig00000433 ;
  wire \blk00000001/sig00000432 ;
  wire \blk00000001/sig00000431 ;
  wire \blk00000001/sig00000430 ;
  wire \blk00000001/sig0000042f ;
  wire \blk00000001/sig0000042e ;
  wire \blk00000001/sig0000042d ;
  wire \blk00000001/sig0000042c ;
  wire \blk00000001/sig0000042b ;
  wire \blk00000001/sig0000042a ;
  wire \blk00000001/sig00000429 ;
  wire \blk00000001/sig00000428 ;
  wire \blk00000001/sig00000427 ;
  wire \blk00000001/sig00000426 ;
  wire \blk00000001/sig00000425 ;
  wire \blk00000001/sig00000424 ;
  wire \blk00000001/sig00000423 ;
  wire \blk00000001/sig00000422 ;
  wire \blk00000001/sig00000421 ;
  wire \blk00000001/sig00000420 ;
  wire \blk00000001/sig0000041f ;
  wire \blk00000001/sig0000041e ;
  wire \blk00000001/sig0000041d ;
  wire \blk00000001/sig0000041c ;
  wire \blk00000001/sig0000041b ;
  wire \blk00000001/sig0000041a ;
  wire \blk00000001/sig00000419 ;
  wire \blk00000001/sig00000418 ;
  wire \blk00000001/sig00000417 ;
  wire \blk00000001/sig00000416 ;
  wire \blk00000001/sig00000415 ;
  wire \blk00000001/sig00000414 ;
  wire \blk00000001/sig00000413 ;
  wire \blk00000001/sig00000412 ;
  wire \blk00000001/sig00000411 ;
  wire \blk00000001/sig00000410 ;
  wire \blk00000001/sig0000040f ;
  wire \blk00000001/sig0000040e ;
  wire \blk00000001/sig0000040d ;
  wire \blk00000001/sig0000040c ;
  wire \blk00000001/sig0000040b ;
  wire \blk00000001/sig0000040a ;
  wire \blk00000001/sig00000409 ;
  wire \blk00000001/sig00000408 ;
  wire \blk00000001/sig00000407 ;
  wire \blk00000001/sig00000406 ;
  wire \blk00000001/sig00000405 ;
  wire \blk00000001/sig00000404 ;
  wire \blk00000001/sig00000403 ;
  wire \blk00000001/sig00000402 ;
  wire \blk00000001/sig00000401 ;
  wire \blk00000001/sig00000400 ;
  wire \blk00000001/sig000003ff ;
  wire \blk00000001/sig000003fe ;
  wire \blk00000001/sig000003fd ;
  wire \blk00000001/sig000003fc ;
  wire \blk00000001/sig000003fb ;
  wire \blk00000001/sig000003fa ;
  wire \blk00000001/sig000003f9 ;
  wire \blk00000001/sig000003f8 ;
  wire \blk00000001/sig000003f7 ;
  wire \blk00000001/sig000003f6 ;
  wire \blk00000001/sig000003f5 ;
  wire \blk00000001/sig000003f4 ;
  wire \blk00000001/sig000003f3 ;
  wire \blk00000001/sig000003f2 ;
  wire \blk00000001/sig000003f1 ;
  wire \blk00000001/sig000003f0 ;
  wire \blk00000001/sig000003ef ;
  wire \blk00000001/sig000003ee ;
  wire \blk00000001/sig000003ed ;
  wire \blk00000001/sig000003ec ;
  wire \blk00000001/sig000003eb ;
  wire \blk00000001/sig000003ea ;
  wire \blk00000001/sig000003e9 ;
  wire \blk00000001/sig000003e8 ;
  wire \blk00000001/sig000003e7 ;
  wire \blk00000001/sig000003e6 ;
  wire \blk00000001/sig000003e5 ;
  wire \blk00000001/sig000003e4 ;
  wire \blk00000001/sig000003e3 ;
  wire \blk00000001/sig000003e2 ;
  wire \blk00000001/sig000003e1 ;
  wire \blk00000001/sig000003e0 ;
  wire \blk00000001/sig000003df ;
  wire \blk00000001/sig000003de ;
  wire \blk00000001/sig000003dd ;
  wire \blk00000001/sig000003dc ;
  wire \blk00000001/sig000003db ;
  wire \blk00000001/sig000003da ;
  wire \blk00000001/sig000003d9 ;
  wire \blk00000001/sig000003d8 ;
  wire \blk00000001/sig000003d7 ;
  wire \blk00000001/sig000003d6 ;
  wire \blk00000001/sig000003d5 ;
  wire \blk00000001/sig000003d4 ;
  wire \blk00000001/sig000003d3 ;
  wire \blk00000001/sig000003d2 ;
  wire \blk00000001/sig000003d1 ;
  wire \blk00000001/sig000003d0 ;
  wire \blk00000001/sig000003cf ;
  wire \blk00000001/sig000003ce ;
  wire \blk00000001/sig000003cd ;
  wire \blk00000001/sig000003cc ;
  wire \blk00000001/sig000003cb ;
  wire \blk00000001/sig000003ca ;
  wire \blk00000001/sig000003c9 ;
  wire \blk00000001/sig000003c8 ;
  wire \blk00000001/sig000003c7 ;
  wire \blk00000001/sig000003c6 ;
  wire \blk00000001/sig000003c5 ;
  wire \blk00000001/sig000003c4 ;
  wire \blk00000001/sig000003c3 ;
  wire \blk00000001/sig000003c2 ;
  wire \blk00000001/sig000003c1 ;
  wire \blk00000001/sig000003c0 ;
  wire \blk00000001/sig000003bf ;
  wire \blk00000001/sig000003be ;
  wire \blk00000001/sig000003bd ;
  wire \blk00000001/sig000003bc ;
  wire \blk00000001/sig000003bb ;
  wire \blk00000001/sig000003ba ;
  wire \blk00000001/sig000003b9 ;
  wire \blk00000001/sig000003b8 ;
  wire \blk00000001/sig000003b7 ;
  wire \blk00000001/sig000003b6 ;
  wire \blk00000001/sig000003b5 ;
  wire \blk00000001/sig000003b4 ;
  wire \blk00000001/sig000003b3 ;
  wire \blk00000001/sig000003b2 ;
  wire \blk00000001/sig000003b1 ;
  wire \blk00000001/sig000003b0 ;
  wire \blk00000001/sig000003af ;
  wire \blk00000001/sig000003ae ;
  wire \blk00000001/sig000003ad ;
  wire \blk00000001/sig000003ac ;
  wire \blk00000001/sig000003ab ;
  wire \blk00000001/sig000003aa ;
  wire \blk00000001/sig000003a9 ;
  wire \blk00000001/sig000003a8 ;
  wire \blk00000001/sig000003a7 ;
  wire \blk00000001/sig000003a6 ;
  wire \blk00000001/sig000003a5 ;
  wire \blk00000001/sig000003a4 ;
  wire \blk00000001/sig000003a3 ;
  wire \blk00000001/sig000003a2 ;
  wire \blk00000001/sig000003a1 ;
  wire \blk00000001/sig000003a0 ;
  wire \blk00000001/sig0000039f ;
  wire \blk00000001/sig0000039e ;
  wire \blk00000001/sig0000039d ;
  wire \blk00000001/sig0000039c ;
  wire \blk00000001/sig0000039b ;
  wire \blk00000001/sig0000039a ;
  wire \blk00000001/sig00000399 ;
  wire \blk00000001/sig00000398 ;
  wire \blk00000001/sig00000397 ;
  wire \blk00000001/sig00000396 ;
  wire \blk00000001/sig00000395 ;
  wire \blk00000001/sig00000394 ;
  wire \blk00000001/sig00000393 ;
  wire \blk00000001/sig00000392 ;
  wire \blk00000001/sig00000391 ;
  wire \blk00000001/sig00000390 ;
  wire \blk00000001/sig0000038f ;
  wire \blk00000001/sig0000038e ;
  wire \blk00000001/sig0000038d ;
  wire \blk00000001/sig0000038c ;
  wire \blk00000001/sig0000038b ;
  wire \blk00000001/sig0000038a ;
  wire \blk00000001/sig00000389 ;
  wire \blk00000001/sig00000388 ;
  wire \blk00000001/sig00000387 ;
  wire \blk00000001/sig00000386 ;
  wire \blk00000001/sig00000385 ;
  wire \blk00000001/sig00000384 ;
  wire \blk00000001/sig00000383 ;
  wire \blk00000001/sig00000382 ;
  wire \blk00000001/sig00000381 ;
  wire \blk00000001/sig00000380 ;
  wire \blk00000001/sig0000037f ;
  wire \blk00000001/sig0000037e ;
  wire \blk00000001/sig0000037d ;
  wire \blk00000001/sig0000037c ;
  wire \blk00000001/sig0000037b ;
  wire \blk00000001/sig0000037a ;
  wire \blk00000001/sig00000379 ;
  wire \blk00000001/sig00000378 ;
  wire \blk00000001/sig00000377 ;
  wire \blk00000001/sig00000376 ;
  wire \blk00000001/sig00000375 ;
  wire \blk00000001/sig00000374 ;
  wire \blk00000001/sig00000373 ;
  wire \blk00000001/sig00000372 ;
  wire \blk00000001/sig00000371 ;
  wire \blk00000001/sig00000370 ;
  wire \blk00000001/sig0000036f ;
  wire \blk00000001/sig0000036e ;
  wire \blk00000001/sig0000036d ;
  wire \blk00000001/sig0000036c ;
  wire \blk00000001/sig0000036b ;
  wire \blk00000001/sig0000036a ;
  wire \blk00000001/sig00000369 ;
  wire \blk00000001/sig00000368 ;
  wire \blk00000001/sig00000367 ;
  wire \blk00000001/sig00000366 ;
  wire \blk00000001/sig00000365 ;
  wire \blk00000001/sig00000364 ;
  wire \blk00000001/sig00000363 ;
  wire \blk00000001/sig00000362 ;
  wire \blk00000001/sig00000361 ;
  wire \blk00000001/sig00000360 ;
  wire \blk00000001/sig0000035f ;
  wire \blk00000001/sig0000035e ;
  wire \blk00000001/sig0000035d ;
  wire \blk00000001/sig0000035c ;
  wire \blk00000001/sig0000035b ;
  wire \blk00000001/sig0000035a ;
  wire \blk00000001/sig00000359 ;
  wire \blk00000001/sig00000358 ;
  wire \blk00000001/sig00000357 ;
  wire \blk00000001/sig00000356 ;
  wire \blk00000001/sig00000355 ;
  wire \blk00000001/sig00000354 ;
  wire \blk00000001/sig00000353 ;
  wire \blk00000001/sig00000352 ;
  wire \blk00000001/sig00000351 ;
  wire \blk00000001/sig00000350 ;
  wire \blk00000001/sig0000034f ;
  wire \blk00000001/sig0000034e ;
  wire \blk00000001/sig0000034d ;
  wire \blk00000001/sig0000034c ;
  wire \blk00000001/sig0000034b ;
  wire \blk00000001/sig0000034a ;
  wire \blk00000001/sig00000349 ;
  wire \blk00000001/sig00000348 ;
  wire \blk00000001/sig00000347 ;
  wire \blk00000001/sig00000346 ;
  wire \blk00000001/sig00000345 ;
  wire \blk00000001/sig00000344 ;
  wire \blk00000001/sig00000343 ;
  wire \blk00000001/sig00000342 ;
  wire \blk00000001/sig00000341 ;
  wire \blk00000001/sig00000340 ;
  wire \blk00000001/sig0000033f ;
  wire \blk00000001/sig0000033e ;
  wire \blk00000001/sig0000033d ;
  wire \blk00000001/sig0000033c ;
  wire \blk00000001/sig0000033b ;
  wire \blk00000001/sig0000033a ;
  wire \blk00000001/sig00000339 ;
  wire \blk00000001/sig00000338 ;
  wire \blk00000001/sig00000337 ;
  wire \blk00000001/sig00000336 ;
  wire \blk00000001/sig00000335 ;
  wire \blk00000001/sig00000334 ;
  wire \blk00000001/sig00000333 ;
  wire \blk00000001/sig00000332 ;
  wire \blk00000001/sig00000331 ;
  wire \blk00000001/sig00000330 ;
  wire \blk00000001/sig0000032f ;
  wire \blk00000001/sig0000032e ;
  wire \blk00000001/sig0000032d ;
  wire \blk00000001/sig0000032c ;
  wire \blk00000001/sig0000032b ;
  wire \blk00000001/sig0000032a ;
  wire \blk00000001/sig00000329 ;
  wire \blk00000001/sig00000328 ;
  wire \blk00000001/sig00000327 ;
  wire \blk00000001/sig00000326 ;
  wire \blk00000001/sig00000325 ;
  wire \blk00000001/sig00000324 ;
  wire \blk00000001/sig00000323 ;
  wire \blk00000001/sig00000322 ;
  wire \blk00000001/sig00000321 ;
  wire \blk00000001/sig00000320 ;
  wire \blk00000001/sig0000031f ;
  wire \blk00000001/sig0000031e ;
  wire \blk00000001/sig0000031d ;
  wire \blk00000001/sig0000031c ;
  wire \blk00000001/sig0000031b ;
  wire \blk00000001/sig0000031a ;
  wire \blk00000001/sig00000319 ;
  wire \blk00000001/sig00000318 ;
  wire \blk00000001/sig00000317 ;
  wire \blk00000001/sig00000316 ;
  wire \blk00000001/sig00000315 ;
  wire \blk00000001/sig00000314 ;
  wire \blk00000001/sig00000313 ;
  wire \blk00000001/sig00000312 ;
  wire \blk00000001/sig00000311 ;
  wire \blk00000001/sig00000310 ;
  wire \blk00000001/sig0000030f ;
  wire \blk00000001/sig0000030e ;
  wire \blk00000001/sig0000030d ;
  wire \blk00000001/sig0000030c ;
  wire \blk00000001/sig0000030b ;
  wire \blk00000001/sig0000030a ;
  wire \blk00000001/sig00000309 ;
  wire \blk00000001/sig00000308 ;
  wire \blk00000001/sig00000307 ;
  wire \blk00000001/sig00000306 ;
  wire \blk00000001/sig00000305 ;
  wire \blk00000001/sig00000304 ;
  wire \blk00000001/sig00000303 ;
  wire \blk00000001/sig00000302 ;
  wire \blk00000001/sig00000301 ;
  wire \blk00000001/sig00000300 ;
  wire \blk00000001/sig000002ff ;
  wire \blk00000001/sig000002fe ;
  wire \blk00000001/sig000002fd ;
  wire \blk00000001/sig000002fc ;
  wire \blk00000001/sig000002fb ;
  wire \blk00000001/sig000002fa ;
  wire \blk00000001/sig000002f9 ;
  wire \blk00000001/sig000002f8 ;
  wire \blk00000001/sig000002f7 ;
  wire \blk00000001/sig000002f6 ;
  wire \blk00000001/sig000002f5 ;
  wire \blk00000001/sig000002f4 ;
  wire \blk00000001/sig000002f3 ;
  wire \blk00000001/sig000002f2 ;
  wire \blk00000001/sig000002f1 ;
  wire \blk00000001/sig000002f0 ;
  wire \blk00000001/sig000002ef ;
  wire \blk00000001/sig000002ee ;
  wire \blk00000001/sig000002ed ;
  wire \blk00000001/sig000002ec ;
  wire \blk00000001/sig000002eb ;
  wire \blk00000001/sig000002ea ;
  wire \blk00000001/sig000002e9 ;
  wire \blk00000001/sig000002e8 ;
  wire \blk00000001/sig000002e7 ;
  wire \blk00000001/sig000002e6 ;
  wire \blk00000001/sig000002e5 ;
  wire \blk00000001/sig000002e4 ;
  wire \blk00000001/sig000002e3 ;
  wire \blk00000001/sig000002e2 ;
  wire \blk00000001/sig000002e1 ;
  wire \blk00000001/sig000002e0 ;
  wire \blk00000001/sig000002df ;
  wire \blk00000001/sig000002de ;
  wire \blk00000001/sig000002dd ;
  wire \blk00000001/sig000002dc ;
  wire \blk00000001/sig000002db ;
  wire \blk00000001/sig000002da ;
  wire \blk00000001/sig000002d9 ;
  wire \blk00000001/sig000002d8 ;
  wire \blk00000001/sig000002d7 ;
  wire \blk00000001/sig000002d6 ;
  wire \blk00000001/sig000002d5 ;
  wire \blk00000001/sig000002d4 ;
  wire \blk00000001/sig000002d3 ;
  wire \blk00000001/sig000002d2 ;
  wire \blk00000001/sig000002d1 ;
  wire \blk00000001/sig000002d0 ;
  wire \blk00000001/sig000002cf ;
  wire \blk00000001/sig000002ce ;
  wire \blk00000001/sig000002cd ;
  wire \blk00000001/sig000002cc ;
  wire \blk00000001/sig000002cb ;
  wire \blk00000001/sig000002ca ;
  wire \blk00000001/sig000002c9 ;
  wire \blk00000001/sig000002c8 ;
  wire \blk00000001/sig000002c7 ;
  wire \blk00000001/sig000002c6 ;
  wire \blk00000001/sig000002c5 ;
  wire \blk00000001/sig000002c4 ;
  wire \blk00000001/sig000002c3 ;
  wire \blk00000001/sig000002c2 ;
  wire \blk00000001/sig000002c1 ;
  wire \blk00000001/sig000002c0 ;
  wire \blk00000001/sig000002bf ;
  wire \blk00000001/sig000002be ;
  wire \blk00000001/sig000002bd ;
  wire \blk00000001/sig000002bc ;
  wire \blk00000001/sig000002bb ;
  wire \blk00000001/sig000002ba ;
  wire \blk00000001/sig000002b9 ;
  wire \blk00000001/sig000002b8 ;
  wire \blk00000001/sig000002b7 ;
  wire \blk00000001/sig000002b6 ;
  wire \blk00000001/sig000002b5 ;
  wire \blk00000001/sig000002b4 ;
  wire \blk00000001/sig000002b3 ;
  wire \blk00000001/sig000002b2 ;
  wire \blk00000001/sig000002b1 ;
  wire \blk00000001/sig000002b0 ;
  wire \blk00000001/sig000002af ;
  wire \blk00000001/sig000002ae ;
  wire \blk00000001/sig000002ad ;
  wire \blk00000001/sig000002ac ;
  wire \blk00000001/sig000002ab ;
  wire \blk00000001/sig000002aa ;
  wire \blk00000001/sig000002a9 ;
  wire \blk00000001/sig000002a8 ;
  wire \blk00000001/sig000002a7 ;
  wire \blk00000001/sig000002a6 ;
  wire \blk00000001/sig000002a5 ;
  wire \blk00000001/sig000002a4 ;
  wire \blk00000001/sig000002a3 ;
  wire \blk00000001/sig000002a2 ;
  wire \blk00000001/sig000002a1 ;
  wire \blk00000001/sig000002a0 ;
  wire \blk00000001/sig0000029f ;
  wire \blk00000001/sig0000029e ;
  wire \blk00000001/sig0000029d ;
  wire \blk00000001/sig0000029c ;
  wire \blk00000001/sig0000029b ;
  wire \blk00000001/sig0000029a ;
  wire \blk00000001/sig00000299 ;
  wire \blk00000001/sig00000298 ;
  wire \blk00000001/sig00000297 ;
  wire \blk00000001/sig00000296 ;
  wire \blk00000001/sig00000295 ;
  wire \blk00000001/sig00000294 ;
  wire \blk00000001/sig00000293 ;
  wire \blk00000001/sig00000292 ;
  wire \blk00000001/sig00000291 ;
  wire \blk00000001/sig00000290 ;
  wire \blk00000001/sig0000028f ;
  wire \blk00000001/sig0000028e ;
  wire \blk00000001/sig0000028d ;
  wire \blk00000001/sig0000028c ;
  wire \blk00000001/sig0000028b ;
  wire \blk00000001/sig0000028a ;
  wire \blk00000001/sig00000289 ;
  wire \blk00000001/sig00000288 ;
  wire \blk00000001/sig00000287 ;
  wire \blk00000001/sig00000286 ;
  wire \blk00000001/sig00000285 ;
  wire \blk00000001/sig00000284 ;
  wire \blk00000001/sig00000283 ;
  wire \blk00000001/sig00000282 ;
  wire \blk00000001/sig00000281 ;
  wire \blk00000001/sig00000280 ;
  wire \blk00000001/sig0000027f ;
  wire \blk00000001/sig0000027e ;
  wire \blk00000001/sig0000027d ;
  wire \blk00000001/sig0000027c ;
  wire \blk00000001/sig0000027b ;
  wire \blk00000001/sig0000027a ;
  wire \blk00000001/sig00000279 ;
  wire \blk00000001/sig00000278 ;
  wire \blk00000001/sig00000277 ;
  wire \blk00000001/sig00000276 ;
  wire \blk00000001/sig00000275 ;
  wire \blk00000001/sig00000274 ;
  wire \blk00000001/sig00000273 ;
  wire \blk00000001/sig00000272 ;
  wire \blk00000001/sig00000271 ;
  wire \blk00000001/sig00000270 ;
  wire \blk00000001/sig0000026f ;
  wire \blk00000001/sig0000026e ;
  wire \blk00000001/sig0000026d ;
  wire \blk00000001/sig0000026c ;
  wire \blk00000001/sig0000026b ;
  wire \blk00000001/sig0000026a ;
  wire \blk00000001/sig00000269 ;
  wire \blk00000001/sig00000268 ;
  wire \blk00000001/sig00000267 ;
  wire \blk00000001/sig00000266 ;
  wire \blk00000001/sig00000265 ;
  wire \blk00000001/sig00000264 ;
  wire \blk00000001/sig00000263 ;
  wire \blk00000001/sig00000262 ;
  wire \blk00000001/sig00000261 ;
  wire \blk00000001/sig00000260 ;
  wire \blk00000001/sig0000025f ;
  wire \blk00000001/sig0000025e ;
  wire \blk00000001/sig0000025d ;
  wire \blk00000001/sig0000025c ;
  wire \blk00000001/sig0000025b ;
  wire \blk00000001/sig0000025a ;
  wire \blk00000001/sig00000259 ;
  wire \blk00000001/sig00000258 ;
  wire \blk00000001/sig00000257 ;
  wire \blk00000001/sig00000256 ;
  wire \blk00000001/sig00000255 ;
  wire \blk00000001/sig00000254 ;
  wire \blk00000001/sig00000253 ;
  wire \blk00000001/sig00000252 ;
  wire \blk00000001/sig00000251 ;
  wire \blk00000001/sig00000250 ;
  wire \blk00000001/sig0000024f ;
  wire \blk00000001/sig0000024e ;
  wire \blk00000001/sig0000024d ;
  wire \blk00000001/sig0000024c ;
  wire \blk00000001/sig0000024b ;
  wire \blk00000001/sig0000024a ;
  wire \blk00000001/sig00000249 ;
  wire \blk00000001/sig00000248 ;
  wire \blk00000001/sig00000247 ;
  wire \blk00000001/sig00000246 ;
  wire \blk00000001/sig00000245 ;
  wire \blk00000001/sig00000244 ;
  wire \blk00000001/sig00000243 ;
  wire \blk00000001/sig00000242 ;
  wire \blk00000001/sig00000241 ;
  wire \blk00000001/sig00000240 ;
  wire \blk00000001/sig0000023f ;
  wire \blk00000001/sig0000023e ;
  wire \blk00000001/sig0000023d ;
  wire \blk00000001/sig0000023c ;
  wire \blk00000001/sig0000023b ;
  wire \blk00000001/sig0000023a ;
  wire \blk00000001/sig00000239 ;
  wire \blk00000001/sig00000238 ;
  wire \blk00000001/sig00000237 ;
  wire \blk00000001/sig00000236 ;
  wire \blk00000001/sig00000235 ;
  wire \blk00000001/sig00000234 ;
  wire \blk00000001/sig00000233 ;
  wire \blk00000001/sig00000232 ;
  wire \blk00000001/sig00000231 ;
  wire \blk00000001/sig00000230 ;
  wire \blk00000001/sig0000022f ;
  wire \blk00000001/sig0000022e ;
  wire \blk00000001/sig0000022d ;
  wire \blk00000001/sig0000022c ;
  wire \blk00000001/sig0000022b ;
  wire \blk00000001/sig0000022a ;
  wire \blk00000001/sig00000229 ;
  wire \blk00000001/sig00000228 ;
  wire \blk00000001/sig00000227 ;
  wire \blk00000001/sig00000226 ;
  wire \blk00000001/sig00000225 ;
  wire \blk00000001/sig00000224 ;
  wire \blk00000001/sig00000223 ;
  wire \blk00000001/sig00000222 ;
  wire \blk00000001/sig00000221 ;
  wire \blk00000001/sig00000220 ;
  wire \blk00000001/sig0000021f ;
  wire \blk00000001/sig0000021e ;
  wire \blk00000001/sig0000021d ;
  wire \blk00000001/sig0000021c ;
  wire \blk00000001/sig0000021b ;
  wire \blk00000001/sig0000021a ;
  wire \blk00000001/sig00000219 ;
  wire \blk00000001/sig00000218 ;
  wire \blk00000001/sig00000217 ;
  wire \blk00000001/sig00000216 ;
  wire \blk00000001/sig00000215 ;
  wire \blk00000001/sig00000214 ;
  wire \blk00000001/sig00000213 ;
  wire \blk00000001/sig00000212 ;
  wire \blk00000001/sig00000211 ;
  wire \blk00000001/sig00000210 ;
  wire \blk00000001/sig0000020f ;
  wire \blk00000001/sig0000020e ;
  wire \blk00000001/sig0000020d ;
  wire \blk00000001/sig0000020c ;
  wire \blk00000001/sig0000020b ;
  wire \blk00000001/sig0000020a ;
  wire \blk00000001/sig00000209 ;
  wire \blk00000001/sig00000208 ;
  wire \blk00000001/sig00000207 ;
  wire \blk00000001/sig00000206 ;
  wire \blk00000001/sig00000205 ;
  wire \blk00000001/sig00000204 ;
  wire \blk00000001/sig00000203 ;
  wire \blk00000001/sig00000202 ;
  wire \blk00000001/sig00000201 ;
  wire \blk00000001/sig00000200 ;
  wire \blk00000001/sig000001ff ;
  wire \blk00000001/sig000001fe ;
  wire \blk00000001/sig000001fd ;
  wire \blk00000001/sig000001fc ;
  wire \blk00000001/sig000001fb ;
  wire \blk00000001/sig000001fa ;
  wire \blk00000001/sig000001f9 ;
  wire \blk00000001/sig000001f8 ;
  wire \blk00000001/sig000001f7 ;
  wire \blk00000001/sig000001f6 ;
  wire \blk00000001/sig000001f5 ;
  wire \blk00000001/sig000001f4 ;
  wire \blk00000001/sig000001f3 ;
  wire \blk00000001/sig000001f2 ;
  wire \blk00000001/sig000001f1 ;
  wire \blk00000001/sig000001f0 ;
  wire \blk00000001/sig000001ef ;
  wire \blk00000001/sig000001ee ;
  wire \blk00000001/sig000001ed ;
  wire \blk00000001/sig000001ec ;
  wire \blk00000001/sig000001eb ;
  wire \blk00000001/sig000001ea ;
  wire \blk00000001/sig000001e9 ;
  wire \blk00000001/sig000001e8 ;
  wire \blk00000001/sig000001e7 ;
  wire \blk00000001/sig000001e6 ;
  wire \blk00000001/sig000001e5 ;
  wire \blk00000001/sig000001e4 ;
  wire \blk00000001/sig000001e3 ;
  wire \blk00000001/sig000001e2 ;
  wire \blk00000001/sig000001e1 ;
  wire \blk00000001/sig000001e0 ;
  wire \blk00000001/sig000001df ;
  wire \blk00000001/sig000001de ;
  wire \blk00000001/sig000001dd ;
  wire \blk00000001/sig000001dc ;
  wire \blk00000001/sig000001db ;
  wire \blk00000001/sig000001da ;
  wire \blk00000001/sig000001d9 ;
  wire \blk00000001/sig000001d8 ;
  wire \blk00000001/sig000001d7 ;
  wire \blk00000001/sig000001d6 ;
  wire \blk00000001/sig000001d5 ;
  wire \blk00000001/sig000001d4 ;
  wire \blk00000001/sig000001d3 ;
  wire \blk00000001/sig000001d2 ;
  wire \blk00000001/sig000001d1 ;
  wire \blk00000001/sig000001d0 ;
  wire \blk00000001/sig000001cf ;
  wire \blk00000001/sig000001ce ;
  wire \blk00000001/sig000001cd ;
  wire \blk00000001/sig000001cc ;
  wire \blk00000001/sig000001cb ;
  wire \blk00000001/sig000001ca ;
  wire \blk00000001/sig000001c9 ;
  wire \blk00000001/sig000001c8 ;
  wire \blk00000001/sig000001c7 ;
  wire \blk00000001/sig000001c6 ;
  wire \blk00000001/sig000001c5 ;
  wire \blk00000001/sig000001c4 ;
  wire \blk00000001/sig000001c3 ;
  wire \blk00000001/sig000001c2 ;
  wire \blk00000001/sig000001c1 ;
  wire \blk00000001/sig000001c0 ;
  wire \blk00000001/sig000001bf ;
  wire \blk00000001/sig000001be ;
  wire \blk00000001/sig000001bd ;
  wire \blk00000001/sig000001bc ;
  wire \blk00000001/sig000001bb ;
  wire \blk00000001/sig000001ba ;
  wire \blk00000001/sig000001b9 ;
  wire \blk00000001/sig000001b8 ;
  wire \blk00000001/sig000001b7 ;
  wire \blk00000001/sig000001b6 ;
  wire \blk00000001/sig000001b5 ;
  wire \blk00000001/sig000001b4 ;
  wire \blk00000001/sig000001b3 ;
  wire \blk00000001/sig000001b2 ;
  wire \blk00000001/sig000001b1 ;
  wire \blk00000001/sig000001b0 ;
  wire \blk00000001/sig000001af ;
  wire \blk00000001/sig000001ae ;
  wire \blk00000001/sig000001ad ;
  wire \blk00000001/sig000001ac ;
  wire \blk00000001/sig000001ab ;
  wire \blk00000001/sig000001aa ;
  wire \blk00000001/sig000001a9 ;
  wire \blk00000001/sig000001a8 ;
  wire \blk00000001/sig000001a7 ;
  wire \blk00000001/sig000001a6 ;
  wire \blk00000001/sig000001a5 ;
  wire \blk00000001/sig000001a4 ;
  wire \blk00000001/sig000001a3 ;
  wire \blk00000001/sig000001a2 ;
  wire \blk00000001/sig000001a1 ;
  wire \blk00000001/sig000001a0 ;
  wire \blk00000001/sig0000019f ;
  wire \blk00000001/sig0000019e ;
  wire \blk00000001/sig0000019d ;
  wire \blk00000001/sig0000019c ;
  wire \blk00000001/sig0000019b ;
  wire \blk00000001/sig0000019a ;
  wire \blk00000001/sig00000199 ;
  wire \blk00000001/sig00000198 ;
  wire \blk00000001/sig00000197 ;
  wire \blk00000001/sig00000196 ;
  wire \blk00000001/sig00000195 ;
  wire \blk00000001/sig00000194 ;
  wire \blk00000001/sig00000193 ;
  wire \blk00000001/sig00000192 ;
  wire \blk00000001/sig00000191 ;
  wire \blk00000001/sig00000190 ;
  wire \blk00000001/sig0000018f ;
  wire \blk00000001/sig0000018e ;
  wire \blk00000001/sig0000018d ;
  wire \blk00000001/sig0000018c ;
  wire \blk00000001/sig0000018b ;
  wire \blk00000001/sig0000018a ;
  wire \blk00000001/sig00000189 ;
  wire \blk00000001/sig00000188 ;
  wire \blk00000001/sig00000187 ;
  wire \blk00000001/sig00000186 ;
  wire \blk00000001/sig00000185 ;
  wire \blk00000001/sig00000184 ;
  wire \blk00000001/sig00000183 ;
  wire \blk00000001/sig00000182 ;
  wire \blk00000001/sig00000181 ;
  wire \blk00000001/sig00000180 ;
  wire \blk00000001/sig0000017f ;
  wire \blk00000001/sig0000017e ;
  wire \blk00000001/sig0000017d ;
  wire \blk00000001/sig0000017c ;
  wire \blk00000001/sig0000017b ;
  wire \blk00000001/sig0000017a ;
  wire \blk00000001/sig00000179 ;
  wire \blk00000001/sig00000178 ;
  wire \blk00000001/sig00000177 ;
  wire \blk00000001/sig00000176 ;
  wire \blk00000001/sig00000175 ;
  wire \blk00000001/sig00000174 ;
  wire \blk00000001/sig00000173 ;
  wire \blk00000001/sig00000172 ;
  wire \blk00000001/sig00000171 ;
  wire \blk00000001/sig00000170 ;
  wire \blk00000001/sig0000016f ;
  wire \blk00000001/sig0000016e ;
  wire \blk00000001/sig0000016d ;
  wire \blk00000001/sig0000016c ;
  wire \blk00000001/sig0000016b ;
  wire \blk00000001/sig0000016a ;
  wire \blk00000001/sig00000169 ;
  wire \blk00000001/sig00000168 ;
  wire \blk00000001/sig00000167 ;
  wire \blk00000001/sig00000166 ;
  wire \blk00000001/sig00000165 ;
  wire \blk00000001/sig00000164 ;
  wire \blk00000001/sig00000163 ;
  wire \blk00000001/sig00000162 ;
  wire \blk00000001/sig00000161 ;
  wire \blk00000001/sig00000160 ;
  wire \blk00000001/sig0000015f ;
  wire \blk00000001/sig0000015e ;
  wire \blk00000001/sig0000015d ;
  wire \blk00000001/sig0000015c ;
  wire \blk00000001/sig0000015b ;
  wire \blk00000001/sig0000015a ;
  wire \blk00000001/sig00000159 ;
  wire \blk00000001/sig00000158 ;
  wire \blk00000001/sig00000157 ;
  wire \blk00000001/sig00000156 ;
  wire \blk00000001/sig00000155 ;
  wire \blk00000001/sig00000154 ;
  wire \blk00000001/sig00000153 ;
  wire \blk00000001/sig00000152 ;
  wire \blk00000001/sig00000151 ;
  wire \blk00000001/sig00000150 ;
  wire \blk00000001/sig0000014f ;
  wire \blk00000001/sig0000014e ;
  wire \blk00000001/sig0000014d ;
  wire \blk00000001/sig0000014c ;
  wire \blk00000001/sig0000014b ;
  wire \blk00000001/sig0000014a ;
  wire \blk00000001/sig00000149 ;
  wire \blk00000001/sig00000148 ;
  wire \blk00000001/sig00000147 ;
  wire \blk00000001/sig00000146 ;
  wire \blk00000001/sig00000145 ;
  wire \blk00000001/sig00000144 ;
  wire \blk00000001/sig00000143 ;
  wire \blk00000001/sig00000142 ;
  wire \blk00000001/sig00000141 ;
  wire \blk00000001/sig00000140 ;
  wire \blk00000001/sig0000013f ;
  wire \blk00000001/sig0000013e ;
  wire \blk00000001/sig0000013d ;
  wire \blk00000001/sig0000013c ;
  wire \blk00000001/sig0000013b ;
  wire \blk00000001/sig0000013a ;
  wire \blk00000001/sig00000139 ;
  wire \blk00000001/sig00000138 ;
  wire \blk00000001/sig00000137 ;
  wire \blk00000001/sig00000136 ;
  wire \blk00000001/sig00000135 ;
  wire \blk00000001/sig00000134 ;
  wire \blk00000001/sig00000133 ;
  wire \blk00000001/sig00000132 ;
  wire \blk00000001/sig00000131 ;
  wire \blk00000001/sig00000130 ;
  wire \blk00000001/sig0000012f ;
  wire \blk00000001/sig0000012e ;
  wire \blk00000001/sig0000012d ;
  wire \blk00000001/sig0000012c ;
  wire \blk00000001/sig0000012b ;
  wire \blk00000001/sig0000012a ;
  wire \blk00000001/sig00000129 ;
  wire \blk00000001/sig00000128 ;
  wire \blk00000001/sig00000127 ;
  wire \blk00000001/sig00000126 ;
  wire \blk00000001/sig00000125 ;
  wire \blk00000001/sig00000124 ;
  wire \blk00000001/sig00000123 ;
  wire \blk00000001/sig00000122 ;
  wire \blk00000001/sig00000121 ;
  wire \blk00000001/sig00000120 ;
  wire \blk00000001/sig0000011f ;
  wire \blk00000001/sig0000011e ;
  wire \blk00000001/sig0000011d ;
  wire \blk00000001/sig0000011c ;
  wire \blk00000001/sig0000011b ;
  wire \blk00000001/sig0000011a ;
  wire \blk00000001/sig00000119 ;
  wire \blk00000001/sig00000118 ;
  wire \blk00000001/sig00000117 ;
  wire \blk00000001/sig00000116 ;
  wire \blk00000001/sig00000115 ;
  wire \blk00000001/sig00000114 ;
  wire \blk00000001/sig00000113 ;
  wire \blk00000001/sig00000112 ;
  wire \blk00000001/sig00000111 ;
  wire \blk00000001/sig00000110 ;
  wire \blk00000001/sig0000010f ;
  wire \blk00000001/sig0000010e ;
  wire \blk00000001/sig0000010d ;
  wire \blk00000001/sig0000010c ;
  wire \blk00000001/sig0000010b ;
  wire \blk00000001/sig0000010a ;
  wire \blk00000001/sig00000109 ;
  wire \blk00000001/sig00000108 ;
  wire \blk00000001/sig00000107 ;
  wire \blk00000001/sig00000106 ;
  wire \blk00000001/sig00000105 ;
  wire \blk00000001/sig00000104 ;
  wire \blk00000001/sig00000103 ;
  wire \blk00000001/sig00000102 ;
  wire \blk00000001/sig00000101 ;
  wire \blk00000001/sig00000100 ;
  wire \blk00000001/sig000000ff ;
  wire \blk00000001/sig000000fe ;
  wire \blk00000001/sig000000fd ;
  wire \blk00000001/sig000000fc ;
  wire \blk00000001/sig000000fb ;
  wire \blk00000001/sig000000fa ;
  wire \blk00000001/sig000000f9 ;
  wire \blk00000001/sig000000f8 ;
  wire \blk00000001/sig000000f7 ;
  wire \blk00000001/sig000000f6 ;
  wire \blk00000001/sig000000f5 ;
  wire \blk00000001/sig000000f4 ;
  wire \blk00000001/sig000000f3 ;
  wire \blk00000001/sig000000f2 ;
  wire \blk00000001/sig000000f1 ;
  wire \blk00000001/sig000000f0 ;
  wire \blk00000001/sig000000ef ;
  wire \blk00000001/sig000000ee ;
  wire \blk00000001/sig000000ed ;
  wire \blk00000001/sig000000ec ;
  wire \blk00000001/sig000000eb ;
  wire \blk00000001/sig000000ea ;
  wire \blk00000001/sig000000e9 ;
  wire \blk00000001/sig000000e8 ;
  wire \blk00000001/sig000000e7 ;
  wire \blk00000001/sig000000e6 ;
  wire \blk00000001/sig000000e5 ;
  wire \blk00000001/sig000000e4 ;
  wire \blk00000001/sig000000e3 ;
  wire \blk00000001/sig000000e2 ;
  wire \blk00000001/sig000000e1 ;
  wire \blk00000001/sig000000e0 ;
  wire \blk00000001/sig000000df ;
  wire \blk00000001/sig000000de ;
  wire \blk00000001/sig000000dd ;
  wire \blk00000001/sig000000dc ;
  wire \blk00000001/sig000000db ;
  wire \blk00000001/sig000000da ;
  wire \blk00000001/sig000000d9 ;
  wire \blk00000001/sig000000d8 ;
  wire \blk00000001/sig000000d7 ;
  wire \blk00000001/sig000000d6 ;
  wire \blk00000001/sig000000d5 ;
  wire \blk00000001/sig000000d4 ;
  wire \blk00000001/sig000000d3 ;
  wire \blk00000001/sig000000d2 ;
  wire \blk00000001/sig000000d1 ;
  wire \blk00000001/sig000000d0 ;
  wire \blk00000001/sig000000cf ;
  wire \blk00000001/sig000000ce ;
  wire \blk00000001/sig000000cd ;
  wire \blk00000001/sig000000cc ;
  wire \blk00000001/sig000000cb ;
  wire \blk00000001/sig000000ca ;
  wire \blk00000001/sig000000c9 ;
  wire \blk00000001/sig000000c8 ;
  wire \blk00000001/sig000000c7 ;
  wire \blk00000001/sig000000c6 ;
  wire \blk00000001/sig000000c5 ;
  wire \blk00000001/sig000000c4 ;
  wire \blk00000001/sig000000c3 ;
  wire \blk00000001/sig000000c2 ;
  wire \blk00000001/sig000000c1 ;
  wire \blk00000001/sig000000c0 ;
  wire \blk00000001/sig000000bf ;
  wire \blk00000001/sig000000be ;
  wire \blk00000001/sig000000bd ;
  wire \blk00000001/sig000000bc ;
  wire \blk00000001/sig000000bb ;
  wire \blk00000001/sig000000ba ;
  wire \blk00000001/sig000000b9 ;
  wire \blk00000001/sig000000b8 ;
  wire \blk00000001/sig000000b7 ;
  wire \blk00000001/sig000000b6 ;
  wire \blk00000001/sig000000b5 ;
  wire \blk00000001/sig000000b4 ;
  wire \blk00000001/sig000000b3 ;
  wire \blk00000001/sig000000b2 ;
  wire \blk00000001/sig000000b1 ;
  wire \blk00000001/sig000000b0 ;
  wire \blk00000001/sig000000af ;
  wire \blk00000001/sig000000ae ;
  wire \blk00000001/sig000000ad ;
  wire \blk00000001/sig000000ac ;
  wire \blk00000001/sig000000ab ;
  wire \blk00000001/sig000000aa ;
  wire \blk00000001/sig000000a9 ;
  wire \blk00000001/sig000000a8 ;
  wire \blk00000001/sig000000a7 ;
  wire \blk00000001/sig000000a6 ;
  wire \blk00000001/sig000000a5 ;
  wire \blk00000001/sig000000a4 ;
  wire \blk00000001/sig000000a3 ;
  wire \blk00000001/sig000000a2 ;
  wire \blk00000001/sig000000a1 ;
  wire \blk00000001/sig000000a0 ;
  wire \blk00000001/sig0000009f ;
  wire \blk00000001/sig0000009e ;
  wire \blk00000001/sig0000009d ;
  wire \blk00000001/sig0000009c ;
  wire \blk00000001/sig0000009b ;
  wire \blk00000001/sig0000009a ;
  wire \blk00000001/sig00000099 ;
  wire \blk00000001/sig00000098 ;
  wire \blk00000001/sig00000097 ;
  wire \blk00000001/sig00000096 ;
  wire \blk00000001/sig00000095 ;
  wire \blk00000001/sig00000094 ;
  wire \blk00000001/sig00000093 ;
  wire \blk00000001/sig00000092 ;
  wire \blk00000001/sig00000091 ;
  wire \blk00000001/sig00000090 ;
  wire \blk00000001/sig0000008f ;
  wire \blk00000001/sig0000008e ;
  wire \blk00000001/sig0000008d ;
  wire \blk00000001/sig0000008c ;
  wire \blk00000001/sig0000008b ;
  wire \blk00000001/sig0000008a ;
  wire \blk00000001/sig00000089 ;
  wire \blk00000001/sig00000088 ;
  wire \blk00000001/sig00000087 ;
  wire \blk00000001/sig00000086 ;
  wire \blk00000001/sig00000085 ;
  wire \blk00000001/sig00000084 ;
  wire \blk00000001/sig00000083 ;
  wire \blk00000001/sig00000082 ;
  wire \blk00000001/sig00000081 ;
  wire \blk00000001/sig00000080 ;
  wire \blk00000001/sig0000007f ;
  wire \blk00000001/sig0000007e ;
  wire \blk00000001/sig0000007d ;
  wire \blk00000001/sig0000007c ;
  wire \blk00000001/sig0000007b ;
  wire \blk00000001/sig0000007a ;
  wire \blk00000001/sig00000079 ;
  wire \blk00000001/sig00000078 ;
  wire \blk00000001/sig00000077 ;
  wire \blk00000001/sig00000076 ;
  wire \blk00000001/sig00000075 ;
  wire \blk00000001/sig00000074 ;
  wire \blk00000001/sig00000073 ;
  wire \blk00000001/sig00000072 ;
  wire \blk00000001/sig00000071 ;
  wire \blk00000001/sig00000070 ;
  wire \blk00000001/sig0000006f ;
  wire \blk00000001/sig0000006e ;
  wire \blk00000001/sig0000006d ;
  wire \blk00000001/sig0000006c ;
  wire \blk00000001/sig0000006b ;
  wire \blk00000001/sig0000006a ;
  wire \blk00000001/sig00000069 ;
  wire \blk00000001/sig00000068 ;
  wire \blk00000001/sig00000067 ;
  wire \blk00000001/sig00000066 ;
  wire \blk00000001/sig00000065 ;
  wire \blk00000001/sig00000064 ;
  wire \blk00000001/sig00000063 ;
  wire \blk00000001/sig00000062 ;
  wire \blk00000001/sig00000061 ;
  wire \blk00000001/sig00000060 ;
  wire \blk00000001/sig0000005f ;
  wire \blk00000001/sig0000005e ;
  wire \blk00000001/sig0000005d ;
  wire \blk00000001/sig0000005c ;
  wire \blk00000001/sig0000005b ;
  wire \blk00000001/sig0000005a ;
  wire \blk00000001/sig00000059 ;
  wire \blk00000001/sig00000058 ;
  wire \blk00000001/sig00000057 ;
  wire \blk00000001/sig00000056 ;
  wire \blk00000001/sig00000055 ;
  wire \blk00000001/sig00000054 ;
  wire \blk00000001/sig00000053 ;
  wire \blk00000001/sig00000052 ;
  wire \blk00000001/sig00000051 ;
  wire \blk00000001/sig00000050 ;
  wire \blk00000001/sig0000004f ;
  wire \blk00000001/sig0000004e ;
  wire \blk00000001/sig0000004d ;
  wire \blk00000001/sig0000004c ;
  wire \blk00000001/sig0000004b ;
  wire \blk00000001/sig0000004a ;
  wire \blk00000001/sig00000049 ;
  wire \blk00000001/sig00000048 ;
  wire \blk00000001/sig00000047 ;
  wire \blk00000001/sig00000046 ;
  wire \blk00000001/sig00000045 ;
  wire \blk00000001/sig00000044 ;
  wire \blk00000001/sig00000043 ;
  wire \blk00000001/sig00000042 ;
  wire \blk00000001/sig00000041 ;
  wire \blk00000001/sig00000040 ;
  wire \blk00000001/sig0000003f ;
  wire \blk00000001/sig0000003e ;
  wire \blk00000001/sig0000003d ;
  wire \blk00000001/sig0000003c ;
  wire \blk00000001/sig0000003b ;
  wire \blk00000001/sig0000003a ;
  wire \blk00000001/sig00000039 ;
  wire \blk00000001/blk000000ae/sig000006d6 ;
  wire \blk00000001/blk000000ae/sig000006d5 ;
  wire \blk00000001/blk000000ae/sig000006d4 ;
  wire \blk00000001/blk000000ae/sig000006d3 ;
  wire \blk00000001/blk000000ae/sig000006d2 ;
  wire \blk00000001/blk000000ae/sig000006d1 ;
  wire \blk00000001/blk000000ae/sig000006d0 ;
  wire \blk00000001/blk000000ae/sig000006cf ;
  wire \blk00000001/blk000000ae/sig000006ce ;
  wire \blk00000001/blk000000ae/sig000006cd ;
  wire \blk00000001/blk000000ae/sig000006cc ;
  wire \blk00000001/blk000000ae/sig000006cb ;
  wire \blk00000001/blk000000ae/sig000006ca ;
  wire \blk00000001/blk000000ae/sig000006c9 ;
  wire \blk00000001/blk000000ae/sig000006c8 ;
  wire \blk00000001/blk000000ae/sig000006c7 ;
  wire \blk00000001/blk000000ae/sig000006c6 ;
  wire \blk00000001/blk000000ae/sig000006c5 ;
  wire \blk00000001/blk000000ae/sig000006c4 ;
  wire \blk00000001/blk000000ae/sig000006c3 ;
  wire \blk00000001/blk000000ae/sig000006c2 ;
  wire \blk00000001/blk000000ae/sig000006c1 ;
  wire \blk00000001/blk000000ae/sig000006c0 ;
  wire \blk00000001/blk000000ae/sig000006bf ;
  wire \blk00000001/blk000000ae/sig000006be ;
  wire \blk00000001/blk000000ae/sig000006bd ;
  wire \blk00000001/blk000000ae/sig000006bc ;
  wire \blk00000001/blk000000ae/sig000006bb ;
  wire \blk00000001/blk000000ae/sig000006ba ;
  wire \blk00000001/blk000000ae/sig000006b9 ;
  wire \blk00000001/blk000000ae/sig000006b8 ;
  wire \blk00000001/blk000000ae/sig000006b7 ;
  wire \blk00000001/blk000000ae/sig000006b6 ;
  wire \blk00000001/blk000000ae/sig000006b5 ;
  wire \blk00000001/blk000000ae/sig000006b4 ;
  wire \blk00000001/blk000000ae/sig000006b3 ;
  wire \blk00000001/blk000000ae/sig000006b2 ;
  wire \blk00000001/blk000000ae/sig000006b1 ;
  wire \blk00000001/blk000000ae/sig000006b0 ;
  wire \blk00000001/blk000000ae/sig000006af ;
  wire \blk00000001/blk000000ae/sig000006ae ;
  wire \blk00000001/blk000000ae/sig000006ad ;
  wire \blk00000001/blk000000ae/sig000006ac ;
  wire \blk00000001/blk000000ae/sig000006ab ;
  wire \blk00000001/blk000000ae/sig000006aa ;
  wire \blk00000001/blk000000ae/sig000006a9 ;
  wire \blk00000001/blk000000ae/sig000006a8 ;
  wire \blk00000001/blk000000ae/sig000006a7 ;
  wire \blk00000001/blk000000ae/sig000006a6 ;
  wire \blk00000001/blk000000ae/sig000006a5 ;
  wire \blk00000001/blk000000ae/sig000006a4 ;
  wire \blk00000001/blk000000ae/sig000006a3 ;
  wire \blk00000001/blk000000ae/sig000006a2 ;
  wire \blk00000001/blk000000ae/sig000006a1 ;
  wire \blk00000001/blk000000ae/sig000006a0 ;
  wire \blk00000001/blk000000ae/sig0000069f ;
  wire \blk00000001/blk000000ae/sig0000069e ;
  wire \blk00000001/blk000000ae/sig0000069d ;
  wire \blk00000001/blk000000ae/sig0000069c ;
  wire \blk00000001/blk000000ae/sig0000069b ;
  wire \blk00000001/blk000000ae/sig0000069a ;
  wire \blk00000001/blk000000ae/sig00000699 ;
  wire \blk00000001/blk000000ae/sig00000698 ;
  wire \blk00000001/blk000000ae/sig00000697 ;
  wire \blk00000001/blk000000ae/sig00000696 ;
  wire \blk00000001/blk000000ae/sig00000695 ;
  wire \blk00000001/blk000000ae/sig00000694 ;
  wire \blk00000001/blk000000ae/sig00000693 ;
  wire \blk00000001/blk000000ae/sig00000692 ;
  wire \blk00000001/blk000000ae/sig00000691 ;
  wire \blk00000001/blk000000ae/sig00000690 ;
  wire \blk00000001/blk000000ae/sig0000068f ;
  wire \blk00000001/blk000000ae/sig0000068e ;
  wire \blk00000001/blk000000ae/sig0000068d ;
  wire \blk00000001/blk000000ae/sig0000068c ;
  wire \blk00000001/blk000000ae/sig0000068b ;
  wire \blk00000001/blk000000ae/sig0000068a ;
  wire \blk00000001/blk000000ae/sig00000689 ;
  wire \blk00000001/blk000000ae/sig00000688 ;
  wire \blk00000001/blk000000ae/sig00000687 ;
  wire \blk00000001/blk000000ae/sig00000686 ;
  wire \blk00000001/blk000000ae/sig00000685 ;
  wire \blk00000001/blk000000ae/sig00000684 ;
  wire \blk00000001/blk000000ae/sig00000683 ;
  wire \blk00000001/blk000000ae/sig00000682 ;
  wire \blk00000001/blk000000ae/sig00000681 ;
  wire \blk00000001/blk000000ae/sig00000680 ;
  wire \blk00000001/blk000000ae/sig0000067f ;
  wire \blk00000001/blk000000ae/sig0000067e ;
  wire \blk00000001/blk000000ae/sig0000067d ;
  wire \blk00000001/blk000000ae/sig0000067c ;
  wire \blk00000001/blk000000ae/sig0000067b ;
  wire \blk00000001/blk000000ae/sig0000067a ;
  wire \blk00000001/blk000000ae/sig00000679 ;
  wire \blk00000001/blk000000ae/sig00000678 ;
  wire \blk00000001/blk000000ae/sig00000677 ;
  wire \blk00000001/blk000000ae/sig00000676 ;
  wire \blk00000001/blk000000ae/sig00000675 ;
  wire \blk00000001/blk000000ae/sig00000674 ;
  wire \blk00000001/blk000000ae/sig00000673 ;
  wire \blk00000001/blk000000ae/sig00000672 ;
  wire \blk00000001/blk000000ae/sig00000671 ;
  wire \blk00000001/blk000000ae/sig00000670 ;
  wire \blk00000001/blk000000ae/sig0000066f ;
  wire \blk00000001/blk000000ae/sig0000066e ;
  wire \blk00000001/blk000000ae/sig0000066d ;
  wire \blk00000001/blk000000ae/sig0000066c ;
  wire \blk00000001/blk000000ae/sig0000066b ;
  wire \blk00000001/blk000000ae/sig0000066a ;
  wire \blk00000001/blk000000ae/sig00000669 ;
  wire \blk00000001/blk000000ae/sig00000668 ;
  wire \blk00000001/blk000000ae/sig00000667 ;
  wire \blk00000001/blk000000ae/sig00000666 ;
  wire \blk00000001/blk000000ae/sig00000665 ;
  wire \blk00000001/blk000000ae/sig00000664 ;
  wire \blk00000001/blk000000ae/sig00000663 ;
  wire \blk00000001/blk000000ae/sig00000662 ;
  wire \blk00000001/blk000000ae/sig00000661 ;
  wire \blk00000001/blk000000ae/sig00000660 ;
  wire \blk00000001/blk000000ae/sig0000065f ;
  wire \blk00000001/blk000000ae/sig0000065e ;
  wire \blk00000001/blk000000ae/sig0000065d ;
  wire \blk00000001/blk000000ae/sig0000065c ;
  wire \blk00000001/blk000000ae/sig0000065b ;
  wire \blk00000001/blk000000ae/sig0000065a ;
  wire \blk00000001/blk000000ae/sig00000659 ;
  wire \blk00000001/blk000000ae/sig00000658 ;
  wire \blk00000001/blk000000ae/sig00000657 ;
  wire \blk00000001/blk000000ae/sig00000656 ;
  wire \blk00000001/blk000000ae/sig00000655 ;
  wire \blk00000001/blk000000ae/sig00000654 ;
  wire \blk00000001/blk000000ae/sig00000653 ;
  wire \blk00000001/blk000000ae/sig00000652 ;
  wire \blk00000001/blk000000ae/sig00000651 ;
  wire \blk00000001/blk000000ae/sig00000650 ;
  wire \blk00000001/blk000000ae/sig0000064f ;
  wire \blk00000001/blk000000ae/sig0000064e ;
  wire \blk00000001/blk000000ae/sig0000064d ;
  wire \blk00000001/blk000000ae/sig0000064c ;
  wire \blk00000001/blk000000ae/sig0000064b ;
  wire \blk00000001/blk000000ae/sig0000064a ;
  wire \blk00000001/blk000000ae/sig00000649 ;
  wire \blk00000001/blk000000ae/sig00000648 ;
  wire \blk00000001/blk000000ae/sig00000647 ;
  wire \blk00000001/blk000000ae/sig00000646 ;
  wire \blk00000001/blk000000ae/sig00000645 ;
  wire \blk00000001/blk000000ae/sig00000644 ;
  wire \blk00000001/blk000000ae/sig00000643 ;
  wire \blk00000001/blk000000ae/sig00000642 ;
  wire \blk00000001/blk000000ae/sig00000641 ;
  wire \blk00000001/blk000000ae/sig00000640 ;
  wire \blk00000001/blk000000ae/sig0000063f ;
  wire \blk00000001/blk000000ae/sig0000063e ;
  wire \blk00000001/blk000000ae/sig0000063d ;
  wire \blk00000001/blk000000ae/sig0000063c ;
  wire \blk00000001/blk000000ae/sig0000063b ;
  wire \blk00000001/blk000000ae/sig0000063a ;
  wire \blk00000001/blk000000ae/sig00000639 ;
  wire \blk00000001/blk000000ae/sig00000638 ;
  wire \blk00000001/blk000000ae/sig00000637 ;
  wire \blk00000001/blk000000ae/sig00000636 ;
  wire \blk00000001/blk000000ae/sig00000627 ;
  wire \blk00000001/blk000000ae/sig00000626 ;
  wire \blk00000001/blk000000ae/sig00000625 ;
  wire \blk00000001/blk000000ae/sig00000624 ;
  wire \blk00000001/blk000000ae/sig00000623 ;
  wire \blk00000001/blk000000ae/sig00000622 ;
  wire \blk00000001/blk000000ae/sig00000621 ;
  wire \blk00000001/blk000000ae/sig00000620 ;
  wire \blk00000001/blk000000ae/sig0000061f ;
  wire \blk00000001/blk000000ae/sig0000061e ;
  wire \blk00000001/blk000000ae/sig0000061d ;
  wire \blk00000001/blk000000ae/sig0000061c ;
  wire \blk00000001/blk000000ae/sig0000061b ;
  wire \blk00000001/blk000000ae/sig0000061a ;
  wire \blk00000001/blk000000ae/sig00000619 ;
  wire \blk00000001/blk000000ae/sig00000618 ;
  wire \NLW_blk00000001/blk000004ac_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk000004aa_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk000004a8_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk000004a6_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk000004a4_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk000004a2_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk000004a0_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000049e_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000049c_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000049a_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk00000498_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk00000496_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk00000494_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk00000492_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk00000490_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000048e_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000048c_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000048a_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk00000488_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk00000486_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk00000484_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk00000482_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk00000480_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000047e_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000047c_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000047a_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk00000478_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk00000476_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk00000474_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk00000472_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk00000470_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000046e_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000046c_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000046a_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk00000468_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk00000466_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk00000464_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk00000462_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk00000460_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000045e_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000045c_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000045a_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk00000458_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk00000456_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk00000454_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk00000452_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk00000450_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000044e_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000044c_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000044a_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk00000448_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk00000446_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk00000444_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk00000442_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk00000440_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000043e_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000043c_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000043a_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk00000438_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk00000436_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk00000434_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk00000432_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk00000430_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000042e_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000042c_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000042a_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk00000428_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk00000426_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk00000424_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk00000422_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk00000420_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000041e_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000041c_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000041a_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk00000418_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk00000416_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk00000414_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk00000412_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk00000410_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000040e_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000040c_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000040a_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk00000408_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk00000406_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk00000404_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk00000402_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk00000400_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk000003fe_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk000003fc_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk000003fa_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk000003f8_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk000003f6_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk000003f4_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk000003f2_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk000003f0_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk000003ee_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk000003ec_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk000003ea_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk000003e8_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk000003e6_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk000003e4_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk000003e2_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk000003e0_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk000003de_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk000003dc_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk000003da_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk000003d8_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk000003d6_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk000003d4_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk000003d2_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk000003d0_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk000003ce_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk000003cc_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk000003ca_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk000003c8_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk000003c6_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk000003c4_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk000003c2_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk000003c0_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk000003be_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk000003bc_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk000003ba_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk000003b8_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk000003b6_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk000003b4_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk000003b2_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk000003b0_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk000003ae_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk000003ac_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk000003aa_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk000003a8_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk000003a6_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk000003a4_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk000003a2_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk000003a0_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000039e_Q15_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000039d_DIPA<3>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000039d_DIPA<2>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000039d_DOA<31>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000039d_DOA<30>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000039d_DOA<29>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000039d_DOA<28>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000039d_DOA<27>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000039d_DOA<26>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000039d_DOA<25>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000039d_DOA<24>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000039d_DOA<23>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000039d_DOA<22>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000039d_DOA<21>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000039d_DOA<20>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000039d_DOA<19>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000039d_DOA<18>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000039d_DOA<17>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000039d_DOA<16>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000039d_ADDRA<3>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000039d_ADDRA<2>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000039d_ADDRA<1>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000039d_ADDRA<0>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000039d_ADDRB<3>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000039d_ADDRB<2>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000039d_ADDRB<1>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000039d_ADDRB<0>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000039d_DIB<31>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000039d_DIB<30>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000039d_DIB<29>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000039d_DIB<28>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000039d_DIB<27>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000039d_DIB<26>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000039d_DIB<25>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000039d_DIB<24>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000039d_DIB<23>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000039d_DIB<22>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000039d_DIB<21>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000039d_DIB<20>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000039d_DIB<19>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000039d_DIB<18>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000039d_DIB<17>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000039d_DIB<16>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000039d_DOPA<3>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000039d_DOPA<2>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000039d_DIPB<3>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000039d_DIPB<2>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000039d_DOPB<3>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000039d_DOPB<2>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000039d_DOB<31>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000039d_DOB<30>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000039d_DOB<29>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000039d_DOB<28>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000039d_DOB<27>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000039d_DOB<26>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000039d_DOB<25>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000039d_DOB<24>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000039d_DOB<23>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000039d_DOB<22>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000039d_DOB<21>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000039d_DOB<20>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000039d_DOB<19>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000039d_DOB<18>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000039d_DOB<17>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000039d_DOB<16>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000039d_DIA<31>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000039d_DIA<30>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000039d_DIA<29>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000039d_DIA<28>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000039d_DIA<27>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000039d_DIA<26>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000039d_DIA<25>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000039d_DIA<24>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000039d_DIA<23>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000039d_DIA<22>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000039d_DIA<21>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000039d_DIA<20>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000039d_DIA<19>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000039d_DIA<18>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000039d_DIA<17>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000039d_DIA<16>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_CARRYOUTF_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_CARRYOUT_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_BCOUT<17>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_BCOUT<16>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_BCOUT<15>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_BCOUT<14>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_BCOUT<13>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_BCOUT<12>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_BCOUT<11>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_BCOUT<10>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_BCOUT<9>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_BCOUT<8>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_BCOUT<7>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_BCOUT<6>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_BCOUT<5>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_BCOUT<4>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_BCOUT<3>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_BCOUT<2>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_BCOUT<1>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_BCOUT<0>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_P<47>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_P<46>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_P<45>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_P<44>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_P<43>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_P<42>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_P<41>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_P<40>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_P<39>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_P<38>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_P<37>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_P<36>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_P<35>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_P<34>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_P<33>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_P<32>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_P<31>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_P<30>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_P<29>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_PCOUT<47>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_PCOUT<46>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_PCOUT<45>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_PCOUT<44>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_PCOUT<43>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_PCOUT<42>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_PCOUT<41>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_PCOUT<40>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_PCOUT<39>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_PCOUT<38>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_PCOUT<37>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_PCOUT<36>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_PCOUT<35>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_PCOUT<34>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_PCOUT<33>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_PCOUT<32>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_PCOUT<31>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_PCOUT<30>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_PCOUT<29>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_PCOUT<28>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_PCOUT<27>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_PCOUT<26>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_PCOUT<25>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_PCOUT<24>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_PCOUT<23>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_PCOUT<22>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_PCOUT<21>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_PCOUT<20>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_PCOUT<19>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_PCOUT<18>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_PCOUT<17>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_PCOUT<16>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_PCOUT<15>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_PCOUT<14>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_PCOUT<13>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_PCOUT<12>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_PCOUT<11>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_PCOUT<10>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_PCOUT<9>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_PCOUT<8>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_PCOUT<7>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_PCOUT<6>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_PCOUT<5>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_PCOUT<4>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_PCOUT<3>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_PCOUT<2>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_PCOUT<1>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_PCOUT<0>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_M<35>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_M<34>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_M<33>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_M<32>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_M<31>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_M<30>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_M<29>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_M<28>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_M<27>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_M<26>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_M<25>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_M<24>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_M<23>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_M<22>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_M<21>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_M<20>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_M<19>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_M<18>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_M<17>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_M<16>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_M<15>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_M<14>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_M<13>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_M<12>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_M<11>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_M<10>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_M<9>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_M<8>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_M<7>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_M<6>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_M<5>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_M<4>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_M<3>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_M<2>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_M<1>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000020e_M<0>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_CARRYOUTF_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_CARRYOUT_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_BCOUT<17>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_BCOUT<16>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_BCOUT<15>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_BCOUT<14>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_BCOUT<13>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_BCOUT<12>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_BCOUT<11>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_BCOUT<10>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_BCOUT<9>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_BCOUT<8>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_BCOUT<7>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_BCOUT<6>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_BCOUT<5>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_BCOUT<4>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_BCOUT<3>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_BCOUT<2>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_BCOUT<1>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_BCOUT<0>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_P<46>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_P<45>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_P<44>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_P<43>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_P<42>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_P<41>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_P<40>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_P<39>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_P<38>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_P<37>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_P<36>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_P<35>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_P<34>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_PCOUT<47>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_PCOUT<46>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_PCOUT<45>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_PCOUT<44>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_PCOUT<43>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_PCOUT<42>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_PCOUT<41>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_PCOUT<40>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_PCOUT<39>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_PCOUT<38>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_PCOUT<37>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_PCOUT<36>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_PCOUT<35>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_PCOUT<34>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_PCOUT<33>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_PCOUT<32>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_PCOUT<31>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_PCOUT<30>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_PCOUT<29>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_PCOUT<28>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_PCOUT<27>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_PCOUT<26>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_PCOUT<25>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_PCOUT<24>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_PCOUT<23>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_PCOUT<22>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_PCOUT<21>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_PCOUT<20>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_PCOUT<19>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_PCOUT<18>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_PCOUT<17>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_PCOUT<16>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_PCOUT<15>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_PCOUT<14>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_PCOUT<13>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_PCOUT<12>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_PCOUT<11>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_PCOUT<10>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_PCOUT<9>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_PCOUT<8>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_PCOUT<7>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_PCOUT<6>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_PCOUT<5>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_PCOUT<4>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_PCOUT<3>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_PCOUT<2>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_PCOUT<1>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_PCOUT<0>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_M<35>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_M<34>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_M<33>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_M<32>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_M<31>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_M<30>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_M<29>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_M<28>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_M<27>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_M<26>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_M<25>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_M<24>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_M<23>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_M<22>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_M<21>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_M<20>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_M<19>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_M<18>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_M<17>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_M<16>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_M<15>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_M<14>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_M<13>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_M<12>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_M<11>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_M<10>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_M<9>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_M<8>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_M<7>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_M<6>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_M<5>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_M<4>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_M<3>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_M<2>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_M<1>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001da_M<0>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_CARRYOUTF_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_CARRYOUT_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_BCOUT<17>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_BCOUT<16>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_BCOUT<15>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_BCOUT<14>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_BCOUT<13>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_BCOUT<12>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_BCOUT<11>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_BCOUT<10>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_BCOUT<9>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_BCOUT<8>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_BCOUT<7>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_BCOUT<6>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_BCOUT<5>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_BCOUT<4>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_BCOUT<3>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_BCOUT<2>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_BCOUT<1>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_BCOUT<0>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_P<47>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_P<46>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_P<45>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_P<44>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_P<43>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_P<42>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_P<41>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_P<40>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_P<39>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_P<38>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_P<37>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_P<36>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_P<35>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_P<34>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_P<33>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_P<32>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_P<31>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_P<30>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_P<29>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_P<28>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_P<27>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_P<26>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_P<25>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_P<24>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_P<23>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_P<22>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_P<21>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_P<20>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_P<19>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_PCOUT<47>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_PCOUT<46>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_PCOUT<45>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_PCOUT<44>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_PCOUT<43>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_PCOUT<42>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_PCOUT<41>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_PCOUT<40>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_PCOUT<39>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_PCOUT<38>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_PCOUT<37>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_PCOUT<36>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_PCOUT<35>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_PCOUT<34>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_PCOUT<33>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_PCOUT<32>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_PCOUT<31>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_PCOUT<30>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_PCOUT<29>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_PCOUT<28>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_PCOUT<27>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_PCOUT<26>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_PCOUT<25>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_PCOUT<24>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_PCOUT<23>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_PCOUT<22>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_PCOUT<21>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_PCOUT<20>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_PCOUT<19>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_PCOUT<18>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_PCOUT<17>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_PCOUT<16>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_PCOUT<15>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_PCOUT<14>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_PCOUT<13>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_PCOUT<12>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_PCOUT<11>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_PCOUT<10>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_PCOUT<9>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_PCOUT<8>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_PCOUT<7>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_PCOUT<6>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_PCOUT<5>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_PCOUT<4>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_PCOUT<3>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_PCOUT<2>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_PCOUT<1>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_PCOUT<0>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_M<35>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_M<34>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_M<33>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_M<32>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_M<31>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_M<30>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_M<29>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_M<28>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_M<27>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_M<26>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_M<25>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_M<24>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_M<23>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_M<22>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_M<21>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_M<20>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_M<19>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_M<18>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_M<17>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_M<16>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_M<15>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_M<14>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_M<13>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_M<12>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_M<11>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_M<10>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_M<9>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_M<8>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_M<7>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_M<6>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_M<5>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_M<4>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_M<3>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_M<2>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_M<1>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d9_M<0>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_CARRYOUTF_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_CARRYOUT_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_BCOUT<17>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_BCOUT<16>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_BCOUT<15>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_BCOUT<14>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_BCOUT<13>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_BCOUT<12>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_BCOUT<11>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_BCOUT<10>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_BCOUT<9>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_BCOUT<8>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_BCOUT<7>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_BCOUT<6>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_BCOUT<5>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_BCOUT<4>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_BCOUT<3>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_BCOUT<2>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_BCOUT<1>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_BCOUT<0>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_P<47>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_P<46>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_P<45>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_P<44>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_P<43>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_P<42>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_P<41>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_P<40>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_P<39>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_P<38>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_P<37>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_P<36>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_P<35>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_P<34>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_PCOUT<47>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_PCOUT<46>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_PCOUT<45>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_PCOUT<44>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_PCOUT<43>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_PCOUT<42>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_PCOUT<41>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_PCOUT<40>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_PCOUT<39>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_PCOUT<38>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_PCOUT<37>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_PCOUT<36>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_PCOUT<35>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_PCOUT<34>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_PCOUT<33>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_PCOUT<32>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_PCOUT<31>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_PCOUT<30>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_PCOUT<29>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_PCOUT<28>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_PCOUT<27>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_PCOUT<26>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_PCOUT<25>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_PCOUT<24>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_PCOUT<23>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_PCOUT<22>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_PCOUT<21>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_PCOUT<20>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_PCOUT<19>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_PCOUT<18>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_PCOUT<17>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_PCOUT<16>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_PCOUT<15>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_PCOUT<14>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_PCOUT<13>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_PCOUT<12>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_PCOUT<11>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_PCOUT<10>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_PCOUT<9>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_PCOUT<8>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_PCOUT<7>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_PCOUT<6>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_PCOUT<5>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_PCOUT<4>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_PCOUT<3>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_PCOUT<2>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_PCOUT<1>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_PCOUT<0>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_M<35>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_M<34>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_M<33>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_M<32>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_M<31>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_M<30>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_M<29>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_M<28>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_M<27>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_M<26>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_M<25>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_M<24>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_M<23>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_M<22>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_M<21>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_M<20>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_M<19>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_M<18>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_M<17>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_M<16>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_M<15>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_M<14>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_M<13>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_M<12>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_M<11>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_M<10>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_M<9>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_M<8>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_M<7>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_M<6>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_M<5>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_M<4>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_M<3>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_M<2>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_M<1>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d8_M<0>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_CARRYOUTF_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_CARRYOUT_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_BCOUT<17>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_BCOUT<16>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_BCOUT<15>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_BCOUT<14>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_BCOUT<13>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_BCOUT<12>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_BCOUT<11>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_BCOUT<10>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_BCOUT<9>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_BCOUT<8>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_BCOUT<7>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_BCOUT<6>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_BCOUT<5>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_BCOUT<4>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_BCOUT<3>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_BCOUT<2>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_BCOUT<1>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_BCOUT<0>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_P<47>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_P<46>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_P<45>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_P<44>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_P<43>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_P<42>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_P<41>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_P<40>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_P<39>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_P<38>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_P<37>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_P<36>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_P<35>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_P<34>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_P<33>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_P<32>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_P<31>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_P<30>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_P<29>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_P<28>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_P<27>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_P<26>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_P<25>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_P<24>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_P<23>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_P<22>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_P<21>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_P<20>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_P<19>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_P<18>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_P<17>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_P<16>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_P<15>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_P<14>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_P<13>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_P<12>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_P<11>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_P<10>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_P<9>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_P<8>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_P<7>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_P<6>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_P<5>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_P<4>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_P<3>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_P<2>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_P<1>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_P<0>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_M<35>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_M<34>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_M<33>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_M<32>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_M<31>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_M<30>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_M<29>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_M<28>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_M<27>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_M<26>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_M<25>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_M<24>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_M<23>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_M<22>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_M<21>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_M<20>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_M<19>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_M<18>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_M<17>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_M<16>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_M<15>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_M<14>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_M<13>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_M<12>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_M<11>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_M<10>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_M<9>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_M<8>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_M<7>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_M<6>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_M<5>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_M<4>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_M<3>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_M<2>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_M<1>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d7_M<0>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_CARRYOUTF_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_CARRYOUT_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_BCOUT<17>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_BCOUT<16>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_BCOUT<15>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_BCOUT<14>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_BCOUT<13>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_BCOUT<12>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_BCOUT<11>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_BCOUT<10>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_BCOUT<9>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_BCOUT<8>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_BCOUT<7>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_BCOUT<6>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_BCOUT<5>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_BCOUT<4>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_BCOUT<3>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_BCOUT<2>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_BCOUT<1>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_BCOUT<0>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_P<47>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_P<46>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_P<45>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_P<44>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_P<43>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_P<42>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_P<41>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_P<40>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_P<39>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_P<38>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_P<37>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_P<36>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_P<35>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_P<34>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_P<33>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_P<32>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_P<31>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_P<30>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_P<29>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_P<28>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_P<27>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_P<26>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_P<25>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_P<24>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_P<23>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_P<22>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_P<21>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_P<20>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_P<19>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_P<18>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_P<17>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_P<16>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_P<15>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_P<14>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_P<13>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_P<12>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_P<11>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_P<10>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_P<9>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_P<8>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_P<7>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_P<6>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_P<5>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_P<4>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_P<3>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_P<2>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_P<1>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_P<0>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_M<35>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_M<34>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_M<33>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_M<32>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_M<31>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_M<30>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_M<29>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_M<28>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_M<27>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_M<26>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_M<25>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_M<24>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_M<23>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_M<22>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_M<21>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_M<20>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_M<19>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_M<18>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_M<17>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_M<16>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_M<15>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_M<14>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_M<13>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_M<12>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_M<11>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_M<10>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_M<9>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_M<8>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_M<7>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_M<6>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_M<5>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_M<4>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_M<3>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_M<2>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_M<1>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d6_M<0>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_CARRYOUTF_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_CARRYOUT_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_BCOUT<17>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_BCOUT<16>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_BCOUT<15>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_BCOUT<14>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_BCOUT<13>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_BCOUT<12>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_BCOUT<11>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_BCOUT<10>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_BCOUT<9>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_BCOUT<8>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_BCOUT<7>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_BCOUT<6>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_BCOUT<5>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_BCOUT<4>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_BCOUT<3>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_BCOUT<2>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_BCOUT<1>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_BCOUT<0>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_P<47>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_P<46>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_P<45>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_P<44>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_P<43>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_P<42>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_P<41>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_P<40>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_P<39>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_P<38>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_P<37>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_P<36>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_P<35>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_P<34>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_P<33>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_P<32>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_P<31>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_P<30>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_P<29>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_P<28>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_P<27>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_P<26>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_P<25>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_P<24>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_P<23>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_P<22>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_P<21>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_P<20>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_P<19>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_P<18>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_P<17>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_P<16>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_P<15>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_P<14>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_P<13>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_P<12>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_P<11>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_P<10>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_P<9>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_P<8>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_P<7>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_P<6>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_P<5>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_P<4>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_P<3>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_P<2>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_P<1>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_P<0>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_M<35>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_M<34>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_M<33>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_M<32>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_M<31>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_M<30>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_M<29>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_M<28>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_M<27>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_M<26>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_M<25>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_M<24>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_M<23>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_M<22>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_M<21>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_M<20>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_M<19>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_M<18>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_M<17>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_M<16>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_M<15>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_M<14>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_M<13>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_M<12>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_M<11>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_M<10>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_M<9>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_M<8>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_M<7>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_M<6>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_M<5>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_M<4>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_M<3>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_M<2>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_M<1>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000001d5_M<0>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_CARRYOUTF_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_CARRYOUT_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_BCOUT<17>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_BCOUT<16>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_BCOUT<15>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_BCOUT<14>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_BCOUT<13>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_BCOUT<12>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_BCOUT<11>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_BCOUT<10>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_BCOUT<9>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_BCOUT<8>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_BCOUT<7>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_BCOUT<6>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_BCOUT<5>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_BCOUT<4>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_BCOUT<3>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_BCOUT<2>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_BCOUT<1>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_BCOUT<0>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_P<47>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_P<46>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_P<45>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_P<44>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_P<43>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_P<42>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_P<41>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_P<21>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_P<20>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_P<19>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_P<18>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_P<17>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_P<16>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_P<15>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_P<14>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_P<13>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_P<12>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_P<11>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_P<10>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_P<9>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_P<8>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_P<7>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_P<6>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_P<5>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_P<4>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_P<3>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_P<2>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_P<1>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_P<0>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_PCOUT<47>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_PCOUT<46>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_PCOUT<45>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_PCOUT<44>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_PCOUT<43>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_PCOUT<42>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_PCOUT<41>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_PCOUT<40>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_PCOUT<39>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_PCOUT<38>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_PCOUT<37>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_PCOUT<36>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_PCOUT<35>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_PCOUT<34>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_PCOUT<33>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_PCOUT<32>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_PCOUT<31>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_PCOUT<30>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_PCOUT<29>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_PCOUT<28>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_PCOUT<27>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_PCOUT<26>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_PCOUT<25>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_PCOUT<24>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_PCOUT<23>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_PCOUT<22>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_PCOUT<21>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_PCOUT<20>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_PCOUT<19>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_PCOUT<18>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_PCOUT<17>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_PCOUT<16>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_PCOUT<15>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_PCOUT<14>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_PCOUT<13>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_PCOUT<12>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_PCOUT<11>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_PCOUT<10>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_PCOUT<9>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_PCOUT<8>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_PCOUT<7>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_PCOUT<6>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_PCOUT<5>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_PCOUT<4>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_PCOUT<3>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_PCOUT<2>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_PCOUT<1>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_PCOUT<0>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_M<35>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_M<34>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_M<33>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_M<32>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_M<31>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_M<30>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_M<29>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_M<28>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_M<27>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_M<26>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_M<25>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_M<24>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_M<23>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_M<22>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_M<21>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_M<20>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_M<19>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_M<18>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_M<17>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_M<16>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_M<15>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_M<14>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_M<13>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_M<12>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_M<11>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_M<10>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_M<9>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_M<8>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_M<7>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_M<6>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_M<5>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_M<4>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_M<3>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_M<2>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_M<1>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ad_M<0>_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000004e_O_UNCONNECTED ;
  wire \NLW_blk00000001/blk0000000a_O_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b2_CARRYOUTF_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b2_CARRYOUT_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b2_C<47>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b2_C<46>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b2_C<45>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b2_C<44>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b2_C<43>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b2_C<42>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b2_C<41>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b2_C<40>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b2_C<39>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b2_C<38>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b2_C<37>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b2_C<36>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b2_C<35>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b2_C<34>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b2_C<33>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b2_C<32>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b2_C<31>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b2_C<30>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b2_C<29>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b2_C<28>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b2_C<27>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b2_C<26>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b2_C<25>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b2_C<24>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b2_C<23>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b2_C<22>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b2_C<21>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b2_C<20>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b2_C<19>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b2_C<18>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b2_C<17>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b2_C<16>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b2_C<15>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b2_C<14>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b2_C<13>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b2_C<12>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b2_C<11>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b2_C<10>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b2_C<9>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b2_C<8>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b2_C<7>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b2_C<6>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b2_C<5>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b2_C<4>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b2_C<3>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b2_C<2>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b2_C<1>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b2_C<0>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b2_P<16>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b2_P<15>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b2_P<14>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b2_M<35>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b2_M<34>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b2_M<33>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b2_M<32>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b2_M<31>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b2_M<30>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b2_M<29>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b2_M<28>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b2_M<27>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b2_M<26>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b2_M<25>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b2_M<24>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b2_M<23>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b2_M<22>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b2_M<21>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b2_M<20>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b2_M<19>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b2_M<18>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b2_M<17>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b2_M<16>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b2_M<15>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b2_M<14>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b2_M<13>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b2_M<12>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b2_M<11>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b2_M<10>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b2_M<9>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b2_M<8>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b2_M<7>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b2_M<6>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b2_M<5>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b2_M<4>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b2_M<3>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b2_M<2>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b2_M<1>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b2_M<0>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b1_CARRYOUTF_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b1_CARRYOUT_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b1_BCOUT<17>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b1_BCOUT<16>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b1_BCOUT<15>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b1_BCOUT<14>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b1_BCOUT<13>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b1_BCOUT<12>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b1_BCOUT<11>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b1_BCOUT<10>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b1_BCOUT<9>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b1_BCOUT<8>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b1_BCOUT<7>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b1_BCOUT<6>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b1_BCOUT<5>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b1_BCOUT<4>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b1_BCOUT<3>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b1_BCOUT<2>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b1_BCOUT<1>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b1_BCOUT<0>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b1_P<47>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b1_P<46>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b1_P<45>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b1_P<44>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b1_P<43>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b1_P<42>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b1_P<41>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b1_P<40>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b1_P<39>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b1_P<38>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b1_P<37>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b1_P<36>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b1_P<35>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b1_P<34>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b1_P<33>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b1_P<32>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b1_P<31>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b1_P<30>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b1_P<29>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b1_P<28>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b1_P<27>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b1_P<26>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b1_P<25>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b1_P<24>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b1_P<23>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b1_P<22>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b1_P<21>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b1_P<20>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b1_P<19>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b1_P<18>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b1_P<17>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b1_P<16>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b1_M<35>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b1_M<34>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b1_M<33>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b1_M<32>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b1_M<31>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b1_M<30>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b1_M<29>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b1_M<28>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b1_M<27>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b1_M<26>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b1_M<25>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b1_M<24>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b1_M<23>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b1_M<22>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b1_M<21>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b1_M<20>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b1_M<19>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b1_M<18>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b1_M<17>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b1_M<16>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b1_M<15>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b1_M<14>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b1_M<13>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b1_M<12>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b1_M<11>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b1_M<10>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b1_M<9>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b1_M<8>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b1_M<7>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b1_M<6>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b1_M<5>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b1_M<4>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b1_M<3>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b1_M<2>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b1_M<1>_UNCONNECTED ;
  wire \NLW_blk00000001/blk000000ae/blk000000b1_M<0>_UNCONNECTED ;
  wire [24 : 24] NlwRenamedSignal_m_axis_dout_tdata;
  wire [11 : 0] NlwRenamedSig_OI_m_axis_dout_tdata;
  assign
    m_axis_dout_tdata[31] = NlwRenamedSignal_m_axis_dout_tdata[24],
    m_axis_dout_tdata[30] = NlwRenamedSignal_m_axis_dout_tdata[24],
    m_axis_dout_tdata[29] = NlwRenamedSignal_m_axis_dout_tdata[24],
    m_axis_dout_tdata[28] = NlwRenamedSignal_m_axis_dout_tdata[24],
    m_axis_dout_tdata[27] = NlwRenamedSignal_m_axis_dout_tdata[24],
    m_axis_dout_tdata[26] = NlwRenamedSignal_m_axis_dout_tdata[24],
    m_axis_dout_tdata[25] = NlwRenamedSignal_m_axis_dout_tdata[24],
    m_axis_dout_tdata[24] = NlwRenamedSignal_m_axis_dout_tdata[24],
    m_axis_dout_tdata[11] = NlwRenamedSig_OI_m_axis_dout_tdata[11],
    m_axis_dout_tdata[10] = NlwRenamedSig_OI_m_axis_dout_tdata[10],
    m_axis_dout_tdata[9] = NlwRenamedSig_OI_m_axis_dout_tdata[9],
    m_axis_dout_tdata[8] = NlwRenamedSig_OI_m_axis_dout_tdata[8],
    m_axis_dout_tdata[7] = NlwRenamedSig_OI_m_axis_dout_tdata[7],
    m_axis_dout_tdata[6] = NlwRenamedSig_OI_m_axis_dout_tdata[6],
    m_axis_dout_tdata[5] = NlwRenamedSig_OI_m_axis_dout_tdata[5],
    m_axis_dout_tdata[4] = NlwRenamedSig_OI_m_axis_dout_tdata[4],
    m_axis_dout_tdata[3] = NlwRenamedSig_OI_m_axis_dout_tdata[3],
    m_axis_dout_tdata[2] = NlwRenamedSig_OI_m_axis_dout_tdata[2],
    m_axis_dout_tdata[1] = NlwRenamedSig_OI_m_axis_dout_tdata[1],
    m_axis_dout_tdata[0] = NlwRenamedSig_OI_m_axis_dout_tdata[0],
    s_axis_divisor_tready = NlwRenamedSignal_s_axis_dividend_tready,
    s_axis_dividend_tready = NlwRenamedSignal_s_axis_dividend_tready;
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000004ad  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000005f5 ),
    .Q(m_axis_dout_tvalid)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk000004ac  (
    .A0(\blk00000001/sig0000003a ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000003a ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig0000003b ),
    .Q(\blk00000001/sig000005f5 ),
    .Q15(\NLW_blk00000001/blk000004ac_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000004ab  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000005f4 ),
    .Q(\blk00000001/sig0000009d )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk000004aa  (
    .A0(\blk00000001/sig0000051d ),
    .A1(\blk00000001/sig0000003a ),
    .A2(\blk00000001/sig0000003a ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig00000192 ),
    .Q(\blk00000001/sig000005f4 ),
    .Q15(\NLW_blk00000001/blk000004aa_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000004a9  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000005f3 ),
    .Q(\blk00000001/sig0000003b )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk000004a8  (
    .A0(\blk00000001/sig0000003a ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig0000003c ),
    .Q(\blk00000001/sig000005f3 ),
    .Q15(\NLW_blk00000001/blk000004a8_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000004a7  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000005f2 ),
    .Q(\blk00000001/sig0000007d )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk000004a6  (
    .A0(\blk00000001/sig0000003a ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig000001de ),
    .Q(\blk00000001/sig000005f2 ),
    .Q15(\NLW_blk00000001/blk000004a6_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000004a5  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000005f1 ),
    .Q(\blk00000001/sig0000007e )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk000004a4  (
    .A0(\blk00000001/sig0000003a ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig000001df ),
    .Q(\blk00000001/sig000005f1 ),
    .Q15(\NLW_blk00000001/blk000004a4_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000004a3  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000005f0 ),
    .Q(\blk00000001/sig00000192 )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk000004a2  (
    .A0(\blk00000001/sig0000051d ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig000000f6 ),
    .Q(\blk00000001/sig000005f0 ),
    .Q15(\NLW_blk00000001/blk000004a2_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000004a1  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000005ef ),
    .Q(\blk00000001/sig0000003c )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk000004a0  (
    .A0(\blk00000001/sig0000003a ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000003a ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig0000003d ),
    .Q(\blk00000001/sig000005ef ),
    .Q15(\NLW_blk00000001/blk000004a0_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000049f  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000005ee ),
    .Q(\blk00000001/sig00000546 )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk0000049e  (
    .A0(\blk00000001/sig0000003a ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig0000055c ),
    .Q(\blk00000001/sig000005ee ),
    .Q15(\NLW_blk00000001/blk0000049e_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000049d  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000005ed ),
    .Q(\blk00000001/sig00000547 )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk0000049c  (
    .A0(\blk00000001/sig0000051d ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig00000557 ),
    .Q(\blk00000001/sig000005ed ),
    .Q15(\NLW_blk00000001/blk0000049c_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000049b  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000005ec ),
    .Q(\blk00000001/sig00000548 )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk0000049a  (
    .A0(\blk00000001/sig0000051d ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig00000558 ),
    .Q(\blk00000001/sig000005ec ),
    .Q15(\NLW_blk00000001/blk0000049a_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000499  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000005eb ),
    .Q(\blk00000001/sig00000549 )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk00000498  (
    .A0(\blk00000001/sig0000051d ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig00000559 ),
    .Q(\blk00000001/sig000005eb ),
    .Q15(\NLW_blk00000001/blk00000498_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000497  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000005ea ),
    .Q(\blk00000001/sig0000054a )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk00000496  (
    .A0(\blk00000001/sig0000051d ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig0000055a ),
    .Q(\blk00000001/sig000005ea ),
    .Q15(\NLW_blk00000001/blk00000496_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000495  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000005e9 ),
    .Q(\blk00000001/sig0000054b )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk00000494  (
    .A0(\blk00000001/sig0000051d ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(NlwRenamedSig_OI_m_axis_dout_tdata[0]),
    .Q(\blk00000001/sig000005e9 ),
    .Q15(\NLW_blk00000001/blk00000494_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000493  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000005e8 ),
    .Q(\blk00000001/sig0000054c )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk00000492  (
    .A0(\blk00000001/sig0000051d ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(NlwRenamedSig_OI_m_axis_dout_tdata[1]),
    .Q(\blk00000001/sig000005e8 ),
    .Q15(\NLW_blk00000001/blk00000492_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000491  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000005e7 ),
    .Q(\blk00000001/sig0000054d )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk00000490  (
    .A0(\blk00000001/sig0000051d ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(NlwRenamedSig_OI_m_axis_dout_tdata[2]),
    .Q(\blk00000001/sig000005e7 ),
    .Q15(\NLW_blk00000001/blk00000490_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000048f  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000005e6 ),
    .Q(\blk00000001/sig0000054e )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk0000048e  (
    .A0(\blk00000001/sig0000051d ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(NlwRenamedSig_OI_m_axis_dout_tdata[3]),
    .Q(\blk00000001/sig000005e6 ),
    .Q15(\NLW_blk00000001/blk0000048e_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000048d  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000005e5 ),
    .Q(\blk00000001/sig0000054f )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk0000048c  (
    .A0(\blk00000001/sig0000051d ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(NlwRenamedSig_OI_m_axis_dout_tdata[4]),
    .Q(\blk00000001/sig000005e5 ),
    .Q15(\NLW_blk00000001/blk0000048c_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000048b  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000005e4 ),
    .Q(\blk00000001/sig00000550 )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk0000048a  (
    .A0(\blk00000001/sig0000051d ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(NlwRenamedSig_OI_m_axis_dout_tdata[5]),
    .Q(\blk00000001/sig000005e4 ),
    .Q15(\NLW_blk00000001/blk0000048a_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000489  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000005e3 ),
    .Q(\blk00000001/sig00000551 )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk00000488  (
    .A0(\blk00000001/sig0000051d ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(NlwRenamedSig_OI_m_axis_dout_tdata[6]),
    .Q(\blk00000001/sig000005e3 ),
    .Q15(\NLW_blk00000001/blk00000488_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000487  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000005e2 ),
    .Q(\blk00000001/sig00000552 )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk00000486  (
    .A0(\blk00000001/sig0000051d ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(NlwRenamedSig_OI_m_axis_dout_tdata[7]),
    .Q(\blk00000001/sig000005e2 ),
    .Q15(\NLW_blk00000001/blk00000486_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000485  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000005e1 ),
    .Q(\blk00000001/sig00000553 )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk00000484  (
    .A0(\blk00000001/sig0000051d ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(NlwRenamedSig_OI_m_axis_dout_tdata[8]),
    .Q(\blk00000001/sig000005e1 ),
    .Q15(\NLW_blk00000001/blk00000484_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000483  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000005e0 ),
    .Q(\blk00000001/sig00000555 )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk00000482  (
    .A0(\blk00000001/sig0000051d ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(NlwRenamedSig_OI_m_axis_dout_tdata[10]),
    .Q(\blk00000001/sig000005e0 ),
    .Q15(\NLW_blk00000001/blk00000482_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000481  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000005df ),
    .Q(\blk00000001/sig00000556 )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk00000480  (
    .A0(\blk00000001/sig0000051d ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(NlwRenamedSig_OI_m_axis_dout_tdata[11]),
    .Q(\blk00000001/sig000005df ),
    .Q15(\NLW_blk00000001/blk00000480_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000047f  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000005de ),
    .Q(\blk00000001/sig00000554 )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk0000047e  (
    .A0(\blk00000001/sig0000051d ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(NlwRenamedSig_OI_m_axis_dout_tdata[9]),
    .Q(\blk00000001/sig000005de ),
    .Q15(\NLW_blk00000001/blk0000047e_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000047d  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000005dd ),
    .Q(\blk00000001/sig0000045e )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk0000047c  (
    .A0(\blk00000001/sig0000003a ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig0000044e ),
    .Q(\blk00000001/sig000005dd ),
    .Q15(\NLW_blk00000001/blk0000047c_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000047b  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000005dc ),
    .Q(\blk00000001/sig0000045f )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk0000047a  (
    .A0(\blk00000001/sig0000003a ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig0000044f ),
    .Q(\blk00000001/sig000005dc ),
    .Q15(\NLW_blk00000001/blk0000047a_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000479  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000005db ),
    .Q(\blk00000001/sig00000460 )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk00000478  (
    .A0(\blk00000001/sig0000003a ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig00000450 ),
    .Q(\blk00000001/sig000005db ),
    .Q15(\NLW_blk00000001/blk00000478_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000477  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000005da ),
    .Q(\blk00000001/sig00000461 )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk00000476  (
    .A0(\blk00000001/sig0000003a ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig00000451 ),
    .Q(\blk00000001/sig000005da ),
    .Q15(\NLW_blk00000001/blk00000476_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000475  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000005d9 ),
    .Q(\blk00000001/sig00000462 )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk00000474  (
    .A0(\blk00000001/sig0000003a ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig00000452 ),
    .Q(\blk00000001/sig000005d9 ),
    .Q15(\NLW_blk00000001/blk00000474_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000473  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000005d8 ),
    .Q(\blk00000001/sig00000463 )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk00000472  (
    .A0(\blk00000001/sig0000003a ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig00000453 ),
    .Q(\blk00000001/sig000005d8 ),
    .Q15(\NLW_blk00000001/blk00000472_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000471  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000005d7 ),
    .Q(\blk00000001/sig00000464 )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk00000470  (
    .A0(\blk00000001/sig0000003a ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig00000454 ),
    .Q(\blk00000001/sig000005d7 ),
    .Q15(\NLW_blk00000001/blk00000470_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000046f  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000005d6 ),
    .Q(\blk00000001/sig00000465 )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk0000046e  (
    .A0(\blk00000001/sig0000003a ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig00000455 ),
    .Q(\blk00000001/sig000005d6 ),
    .Q15(\NLW_blk00000001/blk0000046e_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000046d  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000005d5 ),
    .Q(\blk00000001/sig00000466 )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk0000046c  (
    .A0(\blk00000001/sig0000003a ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig00000456 ),
    .Q(\blk00000001/sig000005d5 ),
    .Q15(\NLW_blk00000001/blk0000046c_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000046b  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000005d4 ),
    .Q(\blk00000001/sig00000467 )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk0000046a  (
    .A0(\blk00000001/sig0000003a ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig00000457 ),
    .Q(\blk00000001/sig000005d4 ),
    .Q15(\NLW_blk00000001/blk0000046a_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000469  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000005d3 ),
    .Q(\blk00000001/sig00000468 )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk00000468  (
    .A0(\blk00000001/sig0000003a ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig00000458 ),
    .Q(\blk00000001/sig000005d3 ),
    .Q15(\NLW_blk00000001/blk00000468_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000467  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000005d2 ),
    .Q(\blk00000001/sig00000469 )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk00000466  (
    .A0(\blk00000001/sig0000003a ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig00000459 ),
    .Q(\blk00000001/sig000005d2 ),
    .Q15(\NLW_blk00000001/blk00000466_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000465  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000005d1 ),
    .Q(\blk00000001/sig0000046a )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk00000464  (
    .A0(\blk00000001/sig0000003a ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig0000045a ),
    .Q(\blk00000001/sig000005d1 ),
    .Q15(\NLW_blk00000001/blk00000464_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000463  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000005d0 ),
    .Q(\blk00000001/sig0000046b )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk00000462  (
    .A0(\blk00000001/sig0000003a ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig0000045b ),
    .Q(\blk00000001/sig000005d0 ),
    .Q15(\NLW_blk00000001/blk00000462_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000461  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000005cf ),
    .Q(\blk00000001/sig0000046d )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk00000460  (
    .A0(\blk00000001/sig0000003a ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig0000045d ),
    .Q(\blk00000001/sig000005cf ),
    .Q15(\NLW_blk00000001/blk00000460_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000045f  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000005ce ),
    .Q(\blk00000001/sig000003d7 )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk0000045e  (
    .A0(\blk00000001/sig0000003a ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig000003c7 ),
    .Q(\blk00000001/sig000005ce ),
    .Q15(\NLW_blk00000001/blk0000045e_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000045d  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000005cd ),
    .Q(\blk00000001/sig0000046c )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk0000045c  (
    .A0(\blk00000001/sig0000003a ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig0000045c ),
    .Q(\blk00000001/sig000005cd ),
    .Q15(\NLW_blk00000001/blk0000045c_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000045b  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000005cc ),
    .Q(\blk00000001/sig000003d8 )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk0000045a  (
    .A0(\blk00000001/sig0000003a ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig000003c8 ),
    .Q(\blk00000001/sig000005cc ),
    .Q15(\NLW_blk00000001/blk0000045a_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000459  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000005cb ),
    .Q(\blk00000001/sig000003d9 )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk00000458  (
    .A0(\blk00000001/sig0000003a ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig000003c9 ),
    .Q(\blk00000001/sig000005cb ),
    .Q15(\NLW_blk00000001/blk00000458_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000457  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000005ca ),
    .Q(\blk00000001/sig000003da )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk00000456  (
    .A0(\blk00000001/sig0000003a ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig000003ca ),
    .Q(\blk00000001/sig000005ca ),
    .Q15(\NLW_blk00000001/blk00000456_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000455  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000005c9 ),
    .Q(\blk00000001/sig000003db )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk00000454  (
    .A0(\blk00000001/sig0000003a ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig000003cb ),
    .Q(\blk00000001/sig000005c9 ),
    .Q15(\NLW_blk00000001/blk00000454_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000453  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000005c8 ),
    .Q(\blk00000001/sig000003dc )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk00000452  (
    .A0(\blk00000001/sig0000003a ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig000003cc ),
    .Q(\blk00000001/sig000005c8 ),
    .Q15(\NLW_blk00000001/blk00000452_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000451  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000005c7 ),
    .Q(\blk00000001/sig000003dd )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk00000450  (
    .A0(\blk00000001/sig0000003a ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig000003cd ),
    .Q(\blk00000001/sig000005c7 ),
    .Q15(\NLW_blk00000001/blk00000450_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000044f  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000005c6 ),
    .Q(\blk00000001/sig000003de )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk0000044e  (
    .A0(\blk00000001/sig0000003a ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig000003ce ),
    .Q(\blk00000001/sig000005c6 ),
    .Q15(\NLW_blk00000001/blk0000044e_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000044d  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000005c5 ),
    .Q(\blk00000001/sig000003df )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk0000044c  (
    .A0(\blk00000001/sig0000003a ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig000003cf ),
    .Q(\blk00000001/sig000005c5 ),
    .Q15(\NLW_blk00000001/blk0000044c_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000044b  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000005c4 ),
    .Q(\blk00000001/sig000003e0 )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk0000044a  (
    .A0(\blk00000001/sig0000003a ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig000003d0 ),
    .Q(\blk00000001/sig000005c4 ),
    .Q15(\NLW_blk00000001/blk0000044a_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000449  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000005c3 ),
    .Q(\blk00000001/sig000003e1 )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk00000448  (
    .A0(\blk00000001/sig0000003a ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig000003d1 ),
    .Q(\blk00000001/sig000005c3 ),
    .Q15(\NLW_blk00000001/blk00000448_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000447  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000005c2 ),
    .Q(\blk00000001/sig000003e2 )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk00000446  (
    .A0(\blk00000001/sig0000003a ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig000003d2 ),
    .Q(\blk00000001/sig000005c2 ),
    .Q15(\NLW_blk00000001/blk00000446_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000445  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000005c1 ),
    .Q(\blk00000001/sig000003e3 )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk00000444  (
    .A0(\blk00000001/sig0000003a ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig000003d3 ),
    .Q(\blk00000001/sig000005c1 ),
    .Q15(\NLW_blk00000001/blk00000444_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000443  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000005c0 ),
    .Q(\blk00000001/sig000003e4 )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk00000442  (
    .A0(\blk00000001/sig0000003a ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig000003d4 ),
    .Q(\blk00000001/sig000005c0 ),
    .Q15(\NLW_blk00000001/blk00000442_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000441  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000005bf ),
    .Q(\blk00000001/sig000003e5 )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk00000440  (
    .A0(\blk00000001/sig0000003a ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig000003d5 ),
    .Q(\blk00000001/sig000005bf ),
    .Q15(\NLW_blk00000001/blk00000440_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000043f  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000005be ),
    .Q(\blk00000001/sig0000047e )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk0000043e  (
    .A0(\blk00000001/sig0000051d ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig00000544 ),
    .Q(\blk00000001/sig000005be ),
    .Q15(\NLW_blk00000001/blk0000043e_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000043d  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000005bd ),
    .Q(\blk00000001/sig000004f7 )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk0000043c  (
    .A0(\blk00000001/sig0000003a ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig0000050a ),
    .Q(\blk00000001/sig000005bd ),
    .Q15(\NLW_blk00000001/blk0000043c_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000043b  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000005bc ),
    .Q(\blk00000001/sig000003e6 )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk0000043a  (
    .A0(\blk00000001/sig0000003a ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig000003d6 ),
    .Q(\blk00000001/sig000005bc ),
    .Q15(\NLW_blk00000001/blk0000043a_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000439  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000005bb ),
    .Q(\blk00000001/sig000004f8 )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk00000438  (
    .A0(\blk00000001/sig0000003a ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig0000050b ),
    .Q(\blk00000001/sig000005bb ),
    .Q15(\NLW_blk00000001/blk00000438_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000437  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000005ba ),
    .Q(\blk00000001/sig000004f9 )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk00000436  (
    .A0(\blk00000001/sig0000003a ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig0000050c ),
    .Q(\blk00000001/sig000005ba ),
    .Q15(\NLW_blk00000001/blk00000436_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000435  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000005b9 ),
    .Q(\blk00000001/sig000004fa )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk00000434  (
    .A0(\blk00000001/sig0000003a ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig0000050d ),
    .Q(\blk00000001/sig000005b9 ),
    .Q15(\NLW_blk00000001/blk00000434_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000433  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000005b8 ),
    .Q(\blk00000001/sig000004fb )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk00000432  (
    .A0(\blk00000001/sig0000003a ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig0000050e ),
    .Q(\blk00000001/sig000005b8 ),
    .Q15(\NLW_blk00000001/blk00000432_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000431  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000005b7 ),
    .Q(\blk00000001/sig000004fc )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk00000430  (
    .A0(\blk00000001/sig0000003a ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig0000050f ),
    .Q(\blk00000001/sig000005b7 ),
    .Q15(\NLW_blk00000001/blk00000430_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000042f  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000005b6 ),
    .Q(\blk00000001/sig000004fd )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk0000042e  (
    .A0(\blk00000001/sig0000003a ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig00000510 ),
    .Q(\blk00000001/sig000005b6 ),
    .Q15(\NLW_blk00000001/blk0000042e_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000042d  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000005b5 ),
    .Q(\blk00000001/sig000004fe )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk0000042c  (
    .A0(\blk00000001/sig0000003a ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig00000511 ),
    .Q(\blk00000001/sig000005b5 ),
    .Q15(\NLW_blk00000001/blk0000042c_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000042b  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000005b4 ),
    .Q(\blk00000001/sig000004ff )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk0000042a  (
    .A0(\blk00000001/sig0000003a ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig00000512 ),
    .Q(\blk00000001/sig000005b4 ),
    .Q15(\NLW_blk00000001/blk0000042a_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000429  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000005b3 ),
    .Q(\blk00000001/sig00000500 )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk00000428  (
    .A0(\blk00000001/sig0000003a ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig00000513 ),
    .Q(\blk00000001/sig000005b3 ),
    .Q15(\NLW_blk00000001/blk00000428_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000427  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000005b2 ),
    .Q(\blk00000001/sig00000501 )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk00000426  (
    .A0(\blk00000001/sig0000003a ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig00000514 ),
    .Q(\blk00000001/sig000005b2 ),
    .Q15(\NLW_blk00000001/blk00000426_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000425  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000005b1 ),
    .Q(\blk00000001/sig00000502 )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk00000424  (
    .A0(\blk00000001/sig0000003a ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig00000515 ),
    .Q(\blk00000001/sig000005b1 ),
    .Q15(\NLW_blk00000001/blk00000424_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000423  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000005b0 ),
    .Q(\blk00000001/sig00000503 )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk00000422  (
    .A0(\blk00000001/sig0000003a ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig00000516 ),
    .Q(\blk00000001/sig000005b0 ),
    .Q15(\NLW_blk00000001/blk00000422_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000421  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000005af ),
    .Q(\blk00000001/sig00000504 )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk00000420  (
    .A0(\blk00000001/sig0000003a ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig00000517 ),
    .Q(\blk00000001/sig000005af ),
    .Q15(\NLW_blk00000001/blk00000420_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000041f  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000005ae ),
    .Q(\blk00000001/sig00000505 )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk0000041e  (
    .A0(\blk00000001/sig0000003a ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig00000518 ),
    .Q(\blk00000001/sig000005ae ),
    .Q15(\NLW_blk00000001/blk0000041e_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000041d  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000005ad ),
    .Q(\blk00000001/sig00000507 )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk0000041c  (
    .A0(\blk00000001/sig0000003a ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig0000051a ),
    .Q(\blk00000001/sig000005ad ),
    .Q15(\NLW_blk00000001/blk0000041c_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000041b  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000005ac ),
    .Q(\blk00000001/sig00000508 )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk0000041a  (
    .A0(\blk00000001/sig0000003a ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig0000051b ),
    .Q(\blk00000001/sig000005ac ),
    .Q15(\NLW_blk00000001/blk0000041a_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000419  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000005ab ),
    .Q(\blk00000001/sig00000506 )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk00000418  (
    .A0(\blk00000001/sig0000003a ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig00000519 ),
    .Q(\blk00000001/sig000005ab ),
    .Q15(\NLW_blk00000001/blk00000418_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000417  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000005aa ),
    .Q(\blk00000001/sig00000509 )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk00000416  (
    .A0(\blk00000001/sig0000003a ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig0000051c ),
    .Q(\blk00000001/sig000005aa ),
    .Q15(\NLW_blk00000001/blk00000416_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000415  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000005a9 ),
    .Q(\blk00000001/sig0000003f )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk00000414  (
    .A0(\blk00000001/sig0000051d ),
    .A1(\blk00000001/sig0000003a ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig00000040 ),
    .Q(\blk00000001/sig000005a9 ),
    .Q15(\NLW_blk00000001/blk00000414_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000413  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000005a8 ),
    .Q(\blk00000001/sig0000006a )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk00000412  (
    .A0(\blk00000001/sig0000051d ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig000000b6 ),
    .Q(\blk00000001/sig000005a8 ),
    .Q15(\NLW_blk00000001/blk00000412_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000411  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000005a7 ),
    .Q(\blk00000001/sig0000006b )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk00000410  (
    .A0(\blk00000001/sig0000051d ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig000000b7 ),
    .Q(\blk00000001/sig000005a7 ),
    .Q15(\NLW_blk00000001/blk00000410_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000040f  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000005a6 ),
    .Q(\blk00000001/sig0000006c )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk0000040e  (
    .A0(\blk00000001/sig0000051d ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig000000b8 ),
    .Q(\blk00000001/sig000005a6 ),
    .Q15(\NLW_blk00000001/blk0000040e_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000040d  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000005a5 ),
    .Q(\blk00000001/sig0000006d )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk0000040c  (
    .A0(\blk00000001/sig0000051d ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig000000b9 ),
    .Q(\blk00000001/sig000005a5 ),
    .Q15(\NLW_blk00000001/blk0000040c_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000040b  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000005a4 ),
    .Q(\blk00000001/sig0000006e )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk0000040a  (
    .A0(\blk00000001/sig0000051d ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig000000ba ),
    .Q(\blk00000001/sig000005a4 ),
    .Q15(\NLW_blk00000001/blk0000040a_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000409  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000005a3 ),
    .Q(\blk00000001/sig0000007f )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk00000408  (
    .A0(\blk00000001/sig0000003a ),
    .A1(\blk00000001/sig0000003a ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig000000ac ),
    .Q(\blk00000001/sig000005a3 ),
    .Q15(\NLW_blk00000001/blk00000408_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000407  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000005a2 ),
    .Q(\blk00000001/sig00000080 )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk00000406  (
    .A0(\blk00000001/sig0000003a ),
    .A1(\blk00000001/sig0000003a ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig000000ad ),
    .Q(\blk00000001/sig000005a2 ),
    .Q15(\NLW_blk00000001/blk00000406_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000405  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000005a1 ),
    .Q(\blk00000001/sig00000081 )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk00000404  (
    .A0(\blk00000001/sig0000003a ),
    .A1(\blk00000001/sig0000003a ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig000000ae ),
    .Q(\blk00000001/sig000005a1 ),
    .Q15(\NLW_blk00000001/blk00000404_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000403  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000005a0 ),
    .Q(\blk00000001/sig00000082 )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk00000402  (
    .A0(\blk00000001/sig0000003a ),
    .A1(\blk00000001/sig0000003a ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig000000af ),
    .Q(\blk00000001/sig000005a0 ),
    .Q15(\NLW_blk00000001/blk00000402_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000401  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig0000059f ),
    .Q(\blk00000001/sig00000083 )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk00000400  (
    .A0(\blk00000001/sig0000003a ),
    .A1(\blk00000001/sig0000003a ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig000000b0 ),
    .Q(\blk00000001/sig0000059f ),
    .Q15(\NLW_blk00000001/blk00000400_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000003ff  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig0000059e ),
    .Q(\blk00000001/sig00000085 )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk000003fe  (
    .A0(\blk00000001/sig0000003a ),
    .A1(\blk00000001/sig0000003a ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig000000b2 ),
    .Q(\blk00000001/sig0000059e ),
    .Q15(\NLW_blk00000001/blk000003fe_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000003fd  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig0000059d ),
    .Q(\blk00000001/sig00000086 )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk000003fc  (
    .A0(\blk00000001/sig0000003a ),
    .A1(\blk00000001/sig0000003a ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig000000b3 ),
    .Q(\blk00000001/sig0000059d ),
    .Q15(\NLW_blk00000001/blk000003fc_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000003fb  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig0000059c ),
    .Q(\blk00000001/sig00000084 )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk000003fa  (
    .A0(\blk00000001/sig0000003a ),
    .A1(\blk00000001/sig0000003a ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig000000b1 ),
    .Q(\blk00000001/sig0000059c ),
    .Q15(\NLW_blk00000001/blk000003fa_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000003f9  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig0000059b ),
    .Q(\blk00000001/sig00000087 )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk000003f8  (
    .A0(\blk00000001/sig0000003a ),
    .A1(\blk00000001/sig0000003a ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig000000b4 ),
    .Q(\blk00000001/sig0000059b ),
    .Q15(\NLW_blk00000001/blk000003f8_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000003f7  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig0000059a ),
    .Q(\blk00000001/sig00000088 )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk000003f6  (
    .A0(\blk00000001/sig0000003a ),
    .A1(\blk00000001/sig0000003a ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig000000b5 ),
    .Q(\blk00000001/sig0000059a ),
    .Q15(\NLW_blk00000001/blk000003f6_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000003f5  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000599 ),
    .Q(\blk00000001/sig00000089 )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk000003f4  (
    .A0(\blk00000001/sig0000003a ),
    .A1(\blk00000001/sig0000003a ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig0000003a ),
    .Q(\blk00000001/sig00000599 ),
    .Q15(\NLW_blk00000001/blk000003f4_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000003f3  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000598 ),
    .Q(\blk00000001/sig00000195 )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk000003f2  (
    .A0(\blk00000001/sig0000051d ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig000001da ),
    .Q(\blk00000001/sig00000598 ),
    .Q15(\NLW_blk00000001/blk000003f2_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000003f1  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000597 ),
    .Q(\blk00000001/sig00000196 )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk000003f0  (
    .A0(\blk00000001/sig0000051d ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig000001db ),
    .Q(\blk00000001/sig00000597 ),
    .Q15(\NLW_blk00000001/blk000003f0_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000003ef  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000596 ),
    .Q(\blk00000001/sig00000197 )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk000003ee  (
    .A0(\blk00000001/sig0000051d ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig000001dc ),
    .Q(\blk00000001/sig00000596 ),
    .Q15(\NLW_blk00000001/blk000003ee_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000003ed  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000595 ),
    .Q(\blk00000001/sig00000198 )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk000003ec  (
    .A0(\blk00000001/sig0000051d ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig000001dd ),
    .Q(\blk00000001/sig00000595 ),
    .Q15(\NLW_blk00000001/blk000003ec_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000003eb  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000594 ),
    .Q(\blk00000001/sig00000199 )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk000003ea  (
    .A0(\blk00000001/sig0000051d ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig000001ac ),
    .Q(\blk00000001/sig00000594 ),
    .Q15(\NLW_blk00000001/blk000003ea_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000003e9  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000593 ),
    .Q(\blk00000001/sig0000019a )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk000003e8  (
    .A0(\blk00000001/sig0000051d ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig000001ad ),
    .Q(\blk00000001/sig00000593 ),
    .Q15(\NLW_blk00000001/blk000003e8_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000003e7  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000592 ),
    .Q(\blk00000001/sig0000019b )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk000003e6  (
    .A0(\blk00000001/sig0000051d ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig000001ae ),
    .Q(\blk00000001/sig00000592 ),
    .Q15(\NLW_blk00000001/blk000003e6_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000003e5  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000591 ),
    .Q(\blk00000001/sig0000019c )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk000003e4  (
    .A0(\blk00000001/sig0000051d ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig000001af ),
    .Q(\blk00000001/sig00000591 ),
    .Q15(\NLW_blk00000001/blk000003e4_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000003e3  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000590 ),
    .Q(\blk00000001/sig0000019d )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk000003e2  (
    .A0(\blk00000001/sig0000051d ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig000001b0 ),
    .Q(\blk00000001/sig00000590 ),
    .Q15(\NLW_blk00000001/blk000003e2_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000003e1  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig0000058f ),
    .Q(\blk00000001/sig0000019e )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk000003e0  (
    .A0(\blk00000001/sig0000051d ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig000001b1 ),
    .Q(\blk00000001/sig0000058f ),
    .Q15(\NLW_blk00000001/blk000003e0_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000003df  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig0000058e ),
    .Q(\blk00000001/sig0000019f )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk000003de  (
    .A0(\blk00000001/sig0000051d ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig000001b2 ),
    .Q(\blk00000001/sig0000058e ),
    .Q15(\NLW_blk00000001/blk000003de_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000003dd  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig0000058d ),
    .Q(\blk00000001/sig000001a1 )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk000003dc  (
    .A0(\blk00000001/sig0000051d ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig000001b4 ),
    .Q(\blk00000001/sig0000058d ),
    .Q15(\NLW_blk00000001/blk000003dc_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000003db  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig0000058c ),
    .Q(\blk00000001/sig000001a2 )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk000003da  (
    .A0(\blk00000001/sig0000051d ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig000001b5 ),
    .Q(\blk00000001/sig0000058c ),
    .Q15(\NLW_blk00000001/blk000003da_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000003d9  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig0000058b ),
    .Q(\blk00000001/sig000001a0 )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk000003d8  (
    .A0(\blk00000001/sig0000051d ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig000001b3 ),
    .Q(\blk00000001/sig0000058b ),
    .Q15(\NLW_blk00000001/blk000003d8_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000003d7  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig0000058a ),
    .Q(\blk00000001/sig000001a3 )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk000003d6  (
    .A0(\blk00000001/sig0000051d ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig000001b6 ),
    .Q(\blk00000001/sig0000058a ),
    .Q15(\NLW_blk00000001/blk000003d6_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000003d5  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000589 ),
    .Q(\blk00000001/sig000001a4 )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk000003d4  (
    .A0(\blk00000001/sig0000051d ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig000001b7 ),
    .Q(\blk00000001/sig00000589 ),
    .Q15(\NLW_blk00000001/blk000003d4_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000003d3  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000588 ),
    .Q(\blk00000001/sig000001a5 )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk000003d2  (
    .A0(\blk00000001/sig0000051d ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig000001b8 ),
    .Q(\blk00000001/sig00000588 ),
    .Q15(\NLW_blk00000001/blk000003d2_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000003d1  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000587 ),
    .Q(\blk00000001/sig000001a6 )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk000003d0  (
    .A0(\blk00000001/sig0000051d ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig000001b9 ),
    .Q(\blk00000001/sig00000587 ),
    .Q15(\NLW_blk00000001/blk000003d0_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000003cf  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000586 ),
    .Q(\blk00000001/sig000001a7 )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk000003ce  (
    .A0(\blk00000001/sig0000051d ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig000001ba ),
    .Q(\blk00000001/sig00000586 ),
    .Q15(\NLW_blk00000001/blk000003ce_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000003cd  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000585 ),
    .Q(\blk00000001/sig000001a8 )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk000003cc  (
    .A0(\blk00000001/sig0000051d ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig000001bb ),
    .Q(\blk00000001/sig00000585 ),
    .Q15(\NLW_blk00000001/blk000003cc_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000003cb  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000584 ),
    .Q(\blk00000001/sig000001a9 )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk000003ca  (
    .A0(\blk00000001/sig0000051d ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig000001bc ),
    .Q(\blk00000001/sig00000584 ),
    .Q15(\NLW_blk00000001/blk000003ca_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000003c9  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000583 ),
    .Q(\blk00000001/sig000001aa )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk000003c8  (
    .A0(\blk00000001/sig0000051d ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig000001bd ),
    .Q(\blk00000001/sig00000583 ),
    .Q15(\NLW_blk00000001/blk000003c8_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000003c7  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000582 ),
    .Q(\blk00000001/sig000001de )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk000003c6  (
    .A0(\blk00000001/sig0000051d ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig000000aa ),
    .Q(\blk00000001/sig00000582 ),
    .Q15(\NLW_blk00000001/blk000003c6_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000003c5  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000581 ),
    .Q(\blk00000001/sig000001df )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk000003c4  (
    .A0(\blk00000001/sig0000051d ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig000000ab ),
    .Q(\blk00000001/sig00000581 ),
    .Q15(\NLW_blk00000001/blk000003c4_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000003c3  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000580 ),
    .Q(\blk00000001/sig000001ab )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk000003c2  (
    .A0(\blk00000001/sig0000051d ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig00000194 ),
    .Q(\blk00000001/sig00000580 ),
    .Q15(\NLW_blk00000001/blk000003c2_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000003c1  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig0000057f ),
    .Q(\blk00000001/sig000000cb )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk000003c0  (
    .A0(\blk00000001/sig0000051d ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig000000cf ),
    .Q(\blk00000001/sig0000057f ),
    .Q15(\NLW_blk00000001/blk000003c0_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000003bf  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig0000057e ),
    .Q(\blk00000001/sig000000f6 )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk000003be  (
    .A0(\blk00000001/sig0000003a ),
    .A1(\blk00000001/sig0000003a ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(s_axis_divisor_tdata[12]),
    .Q(\blk00000001/sig0000057e ),
    .Q15(\NLW_blk00000001/blk000003be_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000003bd  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig0000057d ),
    .Q(\blk00000001/sig000000fc )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk000003bc  (
    .A0(\blk00000001/sig0000051d ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig000000c7 ),
    .Q(\blk00000001/sig0000057d ),
    .Q15(\NLW_blk00000001/blk000003bc_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000003bb  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig0000057c ),
    .Q(\blk00000001/sig000000ca )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk000003ba  (
    .A0(\blk00000001/sig0000051d ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig000000ce ),
    .Q(\blk00000001/sig0000057c ),
    .Q15(\NLW_blk00000001/blk000003ba_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000003b9  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig0000057b ),
    .Q(\blk00000001/sig0000009e )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk000003b8  (
    .A0(\blk00000001/sig0000051d ),
    .A1(\blk00000001/sig0000003a ),
    .A2(\blk00000001/sig0000003a ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(s_axis_dividend_tdata[0]),
    .Q(\blk00000001/sig0000057b ),
    .Q15(\NLW_blk00000001/blk000003b8_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000003b7  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig0000057a ),
    .Q(\blk00000001/sig0000009f )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk000003b6  (
    .A0(\blk00000001/sig0000051d ),
    .A1(\blk00000001/sig0000003a ),
    .A2(\blk00000001/sig0000003a ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(s_axis_dividend_tdata[1]),
    .Q(\blk00000001/sig0000057a ),
    .Q15(\NLW_blk00000001/blk000003b6_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000003b5  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000579 ),
    .Q(\blk00000001/sig000000a0 )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk000003b4  (
    .A0(\blk00000001/sig0000051d ),
    .A1(\blk00000001/sig0000003a ),
    .A2(\blk00000001/sig0000003a ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(s_axis_dividend_tdata[2]),
    .Q(\blk00000001/sig00000579 ),
    .Q15(\NLW_blk00000001/blk000003b4_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000003b3  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000578 ),
    .Q(\blk00000001/sig000000a1 )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk000003b2  (
    .A0(\blk00000001/sig0000051d ),
    .A1(\blk00000001/sig0000003a ),
    .A2(\blk00000001/sig0000003a ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(s_axis_dividend_tdata[3]),
    .Q(\blk00000001/sig00000578 ),
    .Q15(\NLW_blk00000001/blk000003b2_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000003b1  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000577 ),
    .Q(\blk00000001/sig000000a2 )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk000003b0  (
    .A0(\blk00000001/sig0000051d ),
    .A1(\blk00000001/sig0000003a ),
    .A2(\blk00000001/sig0000003a ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(s_axis_dividend_tdata[4]),
    .Q(\blk00000001/sig00000577 ),
    .Q15(\NLW_blk00000001/blk000003b0_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000003af  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000576 ),
    .Q(\blk00000001/sig000000a3 )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk000003ae  (
    .A0(\blk00000001/sig0000051d ),
    .A1(\blk00000001/sig0000003a ),
    .A2(\blk00000001/sig0000003a ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(s_axis_dividend_tdata[5]),
    .Q(\blk00000001/sig00000576 ),
    .Q15(\NLW_blk00000001/blk000003ae_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000003ad  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000575 ),
    .Q(\blk00000001/sig000000a4 )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk000003ac  (
    .A0(\blk00000001/sig0000051d ),
    .A1(\blk00000001/sig0000003a ),
    .A2(\blk00000001/sig0000003a ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(s_axis_dividend_tdata[6]),
    .Q(\blk00000001/sig00000575 ),
    .Q15(\NLW_blk00000001/blk000003ac_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000003ab  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000574 ),
    .Q(\blk00000001/sig000000a5 )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk000003aa  (
    .A0(\blk00000001/sig0000051d ),
    .A1(\blk00000001/sig0000003a ),
    .A2(\blk00000001/sig0000003a ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(s_axis_dividend_tdata[7]),
    .Q(\blk00000001/sig00000574 ),
    .Q15(\NLW_blk00000001/blk000003aa_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000003a9  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000573 ),
    .Q(\blk00000001/sig000000a6 )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk000003a8  (
    .A0(\blk00000001/sig0000051d ),
    .A1(\blk00000001/sig0000003a ),
    .A2(\blk00000001/sig0000003a ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(s_axis_dividend_tdata[8]),
    .Q(\blk00000001/sig00000573 ),
    .Q15(\NLW_blk00000001/blk000003a8_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000003a7  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000572 ),
    .Q(\blk00000001/sig000000a7 )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk000003a6  (
    .A0(\blk00000001/sig0000051d ),
    .A1(\blk00000001/sig0000003a ),
    .A2(\blk00000001/sig0000003a ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(s_axis_dividend_tdata[9]),
    .Q(\blk00000001/sig00000572 ),
    .Q15(\NLW_blk00000001/blk000003a6_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000003a5  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000571 ),
    .Q(\blk00000001/sig000000a8 )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk000003a4  (
    .A0(\blk00000001/sig0000051d ),
    .A1(\blk00000001/sig0000003a ),
    .A2(\blk00000001/sig0000003a ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(s_axis_dividend_tdata[10]),
    .Q(\blk00000001/sig00000571 ),
    .Q15(\NLW_blk00000001/blk000003a4_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000003a3  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000570 ),
    .Q(\blk00000001/sig000000a9 )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk000003a2  (
    .A0(\blk00000001/sig0000051d ),
    .A1(\blk00000001/sig0000003a ),
    .A2(\blk00000001/sig0000003a ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(s_axis_dividend_tdata[11]),
    .Q(\blk00000001/sig00000570 ),
    .Q15(\NLW_blk00000001/blk000003a2_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000003a1  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig0000056f ),
    .Q(\blk00000001/sig00000237 )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk000003a0  (
    .A0(\blk00000001/sig0000051d ),
    .A1(\blk00000001/sig0000003a ),
    .A2(\blk00000001/sig0000003a ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(s_axis_dividend_tdata[12]),
    .Q(\blk00000001/sig0000056f ),
    .Q15(\NLW_blk00000001/blk000003a0_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000039f  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig0000056e ),
    .Q(\blk00000001/sig0000003d )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000001/blk0000039e  (
    .A0(\blk00000001/sig0000003a ),
    .A1(\blk00000001/sig0000051d ),
    .A2(\blk00000001/sig0000051d ),
    .A3(\blk00000001/sig0000051d ),
    .CE(\blk00000001/sig0000003a ),
    .CLK(aclk),
    .D(\blk00000001/sig0000003e ),
    .Q(\blk00000001/sig0000056e ),
    .Q15(\NLW_blk00000001/blk0000039e_Q15_UNCONNECTED )
  );
  RAMB16BWER #(
    .INITP_00 ( 256'hAAAAAAAAAAAAAAAAAAAAAAAAAAABFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF ),
    .INITP_01 ( 256'h5555555555555555555555555555555555555555556AAAAAAAAAAAAAAAAAAAAA ),
    .INITP_02 ( 256'h0000000000000000000000000000000000000015555555555555555555555555 ),
    .INITP_03 ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INITP_04 ( 256'h775FD7D777D5FFF77FDFF757D557DD77F77F7FF55F755D5D7F5F75F775D5DD55 ),
    .INITP_05 ( 256'h5F5D5757DDD5DFD577DF5D7D55F75F5F777D55D5DFD7FDFFD775F5FFDDDF5F5F ),
    .INITP_06 ( 256'h75757DD5D5755DFD7FF7557755777D57F777DF57FD57F5D7775FFD77F7DD75DF ),
    .INITP_07 ( 256'h7D7D7DD77755F5DFDD77F5F77D55F7F7F55575755FD7555F7DFD5FDFD5FF5575 ),
    .INIT_00 ( 256'hC3D3C799CB64CF32D303D6D9DAB2DE8FE26FE654EA3CEE29F219F60DFA05FE01 ),
    .INIT_01 ( 256'h894E8CDC906E9403979C9B389ED7A27AA621A9CAAD78B129B4DDB895BC51C010 ),
    .INIT_02 ( 256'h5222557D58DB5C3C5FA16308667369E16D5270C6743D77B87B367EB7823B85C3 ),
    .INIT_03 ( 256'h1E072133246227932AC82DFF3139347637B73AF93E3F418844D448234B754ECA ),
    .INIT_04 ( 256'hECBEEFBFF2C2F5C8F8D0FBDBFEE901F9050C08220B3A0E561174149417B81ADE ),
    .INIT_05 ( 256'hBE0EC0E6C3C1C69EC97ECC61CF45D22CD516D802DAF1DDE2E0D6E3CCE6C5E9C0 ),
    .INIT_06 ( 256'h91C39476972C99E49C9E9F5BA21AA4DBA79EAA64AD2CAFF6B2C3B592B864BB37 ),
    .INIT_07 ( 256'h67AF6A406CD46F697201749B773679D47C747F1781BB8461870A89B58C628F11 ),
    .INIT_08 ( 256'h3FA9421B448E4704497B4BF54E7050ED536D55EE58715AF65D7E60076292651F ),
    .INIT_09 ( 256'h198B1BE01E36208D22E7254227A029FF2C5F2EC23127338D35F5385F3ACB3D39 ),
    .INIT_0A ( 256'hF534F76DF9A7FBE3FE21006102A204E40729096F0BB70E01104C129914E81739 ),
    .INIT_0B ( 256'hD284D4A3D6C4D8E6DB0ADD2FDF56E17FE3A9E5D5E802EA31EC61EE94F0C8F2FD ),
    .INIT_0C ( 256'hB15FB366B56FB779B984BB91BDA0BFB0C1C2C3D5C5E9C7FFCA17CC30CE4AD066 ),
    .INIT_0D ( 256'h91AB939B958E978199769B6D9D649F5DA158A354A551A750A950AB51AD54AF59 ),
    .INIT_0E ( 256'h7350752C770978E87AC77CA97E8B806F8253843A8621880A89F48BE08DCD8FBB ),
    .INIT_0F ( 256'h563A580259CB5B965D625F2F60FD62CD649E667068436A176BED6DC46F9C7175 ),
    .INIT_10 ( 256'h3A533C093DC03F78413142EC44A74664482249E04BA14D624F2450E852AC5472 ),
    .INIT_11 ( 256'h1F8B212F22D5247B262327CC29752B202CCC2E79302731D73387353836EB389E ),
    .INIT_12 ( 256'h05CF076308F80A8F0C260DBE0F5710F1128C142815C6176419031AA41C451DE7 ),
    .INIT_13 ( 256'hED11EE96F01CF1A2F32AF4B2F63CF7C6F951FADEFC6BFDF9FF89011902AA043C ),
    .INIT_14 ( 256'hD543D6B9D830D9A8DB21DC9ADE15DF90E10DE28AE408E588E708E889EA0BEB8D ),
    .INIT_15 ( 256'hBE56BFBEC127C291C3FCC568C6D5C842C9B1CB20CC90CE01CF73D0E5D259D3CD ),
    .INIT_16 ( 256'hA83EA99AAAF6AC53ADB1AF0FB06FB1CFB330B492B5F4B758B8BCBA21BB87BCEE ),
    .INIT_17 ( 256'h92F19440959096E1983299849AD79C2B9D7F9ED4A02AA181A2D8A431A58AA6E4 ),
    .INIT_18 ( 256'h7E637FA780EB8230837584BB8602874A889389DC8B268C718DBC8F08905591A3 ),
    .INIT_19 ( 256'h6A8B6BC36CFC6E366F7070AB71E773247461759F76DD781C795C7A9D7BDE7D20 ),
    .INIT_1A ( 256'h575F588D59BB5AEA5C1A5D4B5E7C5FAD60E062136347647B65B066E6681C6953 ),
    .INIT_1B ( 256'h44D645FA471F4844496A4A904BB74CDF4E074F2F5059518352AE53D955055632 ),
    .INIT_1C ( 256'h32EA3404351F363B3757387439913AAF3BCD3CEC3E0C3F2C404D416E429143B3 ),
    .INIT_1D ( 256'h219122A323B424C725DA26ED280229162A2B2B412C582D6F2E862F9E30B731D0 ),
    .INIT_1E ( 256'h10C611CE12D813E114EC15F71702180E191A1A271B351C431D511E611F702080 ),
    .INIT_1F ( 256'h008101810282038404860588068B078F089309970A9C0BA20CA80DAF0EB60FBD ),
    .INIT_20 ( 256'h03B80378033C030402C8028C0250021401D801980158011C00E000A000600040 ),
    .INIT_21 ( 256'h073406FC06C80694065C062405EC05B405800548050C04D4049C0464042803F0 ),
    .INIT_22 ( 256'h0A680A340A0409D409A00970093C090808D808A40870083C080807D407A0076C ),
    .INIT_23 ( 256'h0D580D2C0D000CD00CA00C740C480C140BE80BBC0B880B580B280AFC0ACC0A98 ),
    .INIT_24 ( 256'h100C0FE40FB80F900F680F380F0C0EE40EBC0E900E600E340E0C0DE00DB00D84 ),
    .INIT_25 ( 256'h128812641240121811EC11C811A411781150112C110010D810B41088105C1034 ),
    .INIT_26 ( 256'h14D814B81490146C144C1424140013DC13B4139013701348132012FC12D812B0 ),
    .INIT_27 ( 256'h16F816D816B81698167416541634161015EC15CC15AC158415641544151C14F8 ),
    .INIT_28 ( 256'h18F418D818B8189818781858183C181C17FC17DC17BC179C177C175C173C171C ),
    .INIT_29 ( 256'h1ACC1AAC1A941A781A581A381A1C1A0419E419C419AC198C196C195019301910 ),
    .INIT_2A ( 256'h1C801C681C4C1C301C141BFC1BE41BC41BA81B901B741B581B3C1B201B001AE8 ),
    .INIT_2B ( 256'h1E181E001DE81DD01DB81D9C1D841D6C1D501D381D201D041CE81CCC1CB81C9C ),
    .INIT_2C ( 256'h1F981F801F681F541F3C1F241F081EF01EDC1EC41EAC1E941E7C1E641E4C1E34 ),
    .INIT_2D ( 256'h20FC20E820D020BC20A42090207C2064204C20342020200C1FF41FDC1FC41FAC ),
    .INIT_2E ( 256'h224C22382220221021F821E421D021BC21A82190217C21682154213C21282110 ),
    .INIT_2F ( 256'h23842374235C234C233C2324231022FC22E822D822C422B0229C22882274225C ),
    .INIT_30 ( 256'h24A8249C24882474246424502440242C241C240823F423E423D023C023AC2394 ),
    .INIT_31 ( 256'h25C025B025A02590257C256C255C2548253825282514250424F424E024D024BC ),
    .INIT_32 ( 256'h26C826B826A4269426882678266426542648263426242614260025F425E425D0 ),
    .INIT_33 ( 256'h27B827AC27A0279027802770276027542744273027242714270426F826E426D4 ),
    .INIT_34 ( 256'h28A4289828882878286C286028502840283028242814280427F827E827DC27CC ),
    .INIT_35 ( 256'h297C2974296829582948293C293029202914290828F828E828DC28D028C028B0 ),
    .INIT_36 ( 256'h2A502A442A382A282A1C2A102A0429F829E829DC29D029C029B429A8299C298C ),
    .INIT_37 ( 256'h2B142B082AFC2AF02AE42AD82ACC2AC02AB42AA42A9C2A902A802A742A682A5C ),
    .INIT_38 ( 256'h2BCC2BC42BB82BAC2BA42B982B882B7C2B742B682B582B502B442B382B2C2B20 ),
    .INIT_39 ( 256'h2C802C742C6C2C602C542C482C3C2C342C282C1C2C142C082BFC2BF02BE42BD8 ),
    .INIT_3A ( 256'h2D282D1C2D142D082CFC2CF42CEC2CE02CD42CC82CC02CB82CA82C9C2C942C8C ),
    .INIT_3B ( 256'h2DC82DBC2DB42DA82DA02D982D882D802D7C2D702D642D582D4C2D482D3C2D30 ),
    .INIT_3C ( 256'h2E602E542E4C2E442E382E302E282E1C2E142E0C2E002DF42DF02DE42DD82DD4 ),
    .INIT_3D ( 256'h2EEC2EE82EE02ED42ECC2EC02EB82EB42EA82E9C2E942E8C2E842E7C2E702E68 ),
    .INIT_3E ( 256'h2F782F702F682F602F542F502F482F3C2F342F2C2F242F1C2F102F082F042EF8 ),
    .INIT_3F ( 256'h2FF82FF42FEC2FE42FDC2FD42FCC2FC42FBC2FB42FAC2FA02F982F942F8C2F80 ),
    .INIT_A ( 36'h000000000 ),
    .INIT_B ( 36'h000000000 ),
    .WRITE_MODE_A ( "WRITE_FIRST" ),
    .WRITE_MODE_B ( "WRITE_FIRST" ),
    .DATA_WIDTH_A ( 18 ),
    .DATA_WIDTH_B ( 18 ),
    .DOA_REG ( 0 ),
    .DOB_REG ( 0 ),
    .EN_RSTRAM_A ( "TRUE" ),
    .EN_RSTRAM_B ( "TRUE" ),
    .RST_PRIORITY_A ( "CE" ),
    .RST_PRIORITY_B ( "CE" ),
    .RSTTYPE ( "SYNC" ),
    .SRVAL_A ( 36'h000000000 ),
    .SRVAL_B ( 36'h000000000 ),
    .SIM_COLLISION_CHECK ( "ALL" ),
    .SIM_DEVICE ( "SPARTAN6" ),
    .INIT_FILE ( "NONE" ))
  \blk00000001/blk0000039d  (
    .REGCEA(\blk00000001/sig0000051d ),
    .CLKA(aclk),
    .ENB(\blk00000001/sig0000003a ),
    .RSTB(\blk00000001/sig0000051d ),
    .CLKB(aclk),
    .REGCEB(\blk00000001/sig0000051d ),
    .RSTA(\blk00000001/sig0000051d ),
    .ENA(\blk00000001/sig0000003a ),
    .DIPA({\NLW_blk00000001/blk0000039d_DIPA<3>_UNCONNECTED , \NLW_blk00000001/blk0000039d_DIPA<2>_UNCONNECTED , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d }),
    .WEA({\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d }),
    .DOA({\NLW_blk00000001/blk0000039d_DOA<31>_UNCONNECTED , \NLW_blk00000001/blk0000039d_DOA<30>_UNCONNECTED ,
\NLW_blk00000001/blk0000039d_DOA<29>_UNCONNECTED , \NLW_blk00000001/blk0000039d_DOA<28>_UNCONNECTED ,
\NLW_blk00000001/blk0000039d_DOA<27>_UNCONNECTED , \NLW_blk00000001/blk0000039d_DOA<26>_UNCONNECTED ,
\NLW_blk00000001/blk0000039d_DOA<25>_UNCONNECTED , \NLW_blk00000001/blk0000039d_DOA<24>_UNCONNECTED ,
\NLW_blk00000001/blk0000039d_DOA<23>_UNCONNECTED , \NLW_blk00000001/blk0000039d_DOA<22>_UNCONNECTED ,
\NLW_blk00000001/blk0000039d_DOA<21>_UNCONNECTED , \NLW_blk00000001/blk0000039d_DOA<20>_UNCONNECTED ,
\NLW_blk00000001/blk0000039d_DOA<19>_UNCONNECTED , \NLW_blk00000001/blk0000039d_DOA<18>_UNCONNECTED ,
\NLW_blk00000001/blk0000039d_DOA<17>_UNCONNECTED , \NLW_blk00000001/blk0000039d_DOA<16>_UNCONNECTED , \blk00000001/sig000001bb ,
\blk00000001/sig000001ba , \blk00000001/sig000001b9 , \blk00000001/sig000001b8 , \blk00000001/sig000001b7 , \blk00000001/sig000001b6 ,
\blk00000001/sig000001b5 , \blk00000001/sig000001b4 , \blk00000001/sig000001b3 , \blk00000001/sig000001b2 , \blk00000001/sig000001b1 ,
\blk00000001/sig000001b0 , \blk00000001/sig000001af , \blk00000001/sig000001ae , \blk00000001/sig000001ad , \blk00000001/sig000001ac }),
    .ADDRA({\blk00000001/sig0000051d , \blk00000001/sig000000b5 , \blk00000001/sig000000b4 , \blk00000001/sig000000b3 , \blk00000001/sig000000b2 ,
\blk00000001/sig000000b1 , \blk00000001/sig000000b0 , \blk00000001/sig000000af , \blk00000001/sig000000ae , \blk00000001/sig000000ad ,
\NLW_blk00000001/blk0000039d_ADDRA<3>_UNCONNECTED , \NLW_blk00000001/blk0000039d_ADDRA<2>_UNCONNECTED ,
\NLW_blk00000001/blk0000039d_ADDRA<1>_UNCONNECTED , \NLW_blk00000001/blk0000039d_ADDRA<0>_UNCONNECTED }),
    .ADDRB({\blk00000001/sig0000003a , \blk00000001/sig000000b5 , \blk00000001/sig000000b4 , \blk00000001/sig000000b3 , \blk00000001/sig000000b2 ,
\blk00000001/sig000000b1 , \blk00000001/sig000000b0 , \blk00000001/sig000000af , \blk00000001/sig000000ae , \blk00000001/sig000000ad ,
\NLW_blk00000001/blk0000039d_ADDRB<3>_UNCONNECTED , \NLW_blk00000001/blk0000039d_ADDRB<2>_UNCONNECTED ,
\NLW_blk00000001/blk0000039d_ADDRB<1>_UNCONNECTED , \NLW_blk00000001/blk0000039d_ADDRB<0>_UNCONNECTED }),
    .DIB({\NLW_blk00000001/blk0000039d_DIB<31>_UNCONNECTED , \NLW_blk00000001/blk0000039d_DIB<30>_UNCONNECTED ,
\NLW_blk00000001/blk0000039d_DIB<29>_UNCONNECTED , \NLW_blk00000001/blk0000039d_DIB<28>_UNCONNECTED ,
\NLW_blk00000001/blk0000039d_DIB<27>_UNCONNECTED , \NLW_blk00000001/blk0000039d_DIB<26>_UNCONNECTED ,
\NLW_blk00000001/blk0000039d_DIB<25>_UNCONNECTED , \NLW_blk00000001/blk0000039d_DIB<24>_UNCONNECTED ,
\NLW_blk00000001/blk0000039d_DIB<23>_UNCONNECTED , \NLW_blk00000001/blk0000039d_DIB<22>_UNCONNECTED ,
\NLW_blk00000001/blk0000039d_DIB<21>_UNCONNECTED , \NLW_blk00000001/blk0000039d_DIB<20>_UNCONNECTED ,
\NLW_blk00000001/blk0000039d_DIB<19>_UNCONNECTED , \NLW_blk00000001/blk0000039d_DIB<18>_UNCONNECTED ,
\NLW_blk00000001/blk0000039d_DIB<17>_UNCONNECTED , \NLW_blk00000001/blk0000039d_DIB<16>_UNCONNECTED , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d }),
    .DOPA({\NLW_blk00000001/blk0000039d_DOPA<3>_UNCONNECTED , \NLW_blk00000001/blk0000039d_DOPA<2>_UNCONNECTED , \blk00000001/sig000001bd ,
\blk00000001/sig000001bc }),
    .DIPB({\NLW_blk00000001/blk0000039d_DIPB<3>_UNCONNECTED , \NLW_blk00000001/blk0000039d_DIPB<2>_UNCONNECTED , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d }),
    .DOPB({\NLW_blk00000001/blk0000039d_DOPB<3>_UNCONNECTED , \NLW_blk00000001/blk0000039d_DOPB<2>_UNCONNECTED , \blk00000001/sig000001dd ,
\blk00000001/sig000001dc }),
    .DOB({\NLW_blk00000001/blk0000039d_DOB<31>_UNCONNECTED , \NLW_blk00000001/blk0000039d_DOB<30>_UNCONNECTED ,
\NLW_blk00000001/blk0000039d_DOB<29>_UNCONNECTED , \NLW_blk00000001/blk0000039d_DOB<28>_UNCONNECTED ,
\NLW_blk00000001/blk0000039d_DOB<27>_UNCONNECTED , \NLW_blk00000001/blk0000039d_DOB<26>_UNCONNECTED ,
\NLW_blk00000001/blk0000039d_DOB<25>_UNCONNECTED , \NLW_blk00000001/blk0000039d_DOB<24>_UNCONNECTED ,
\NLW_blk00000001/blk0000039d_DOB<23>_UNCONNECTED , \NLW_blk00000001/blk0000039d_DOB<22>_UNCONNECTED ,
\NLW_blk00000001/blk0000039d_DOB<21>_UNCONNECTED , \NLW_blk00000001/blk0000039d_DOB<20>_UNCONNECTED ,
\NLW_blk00000001/blk0000039d_DOB<19>_UNCONNECTED , \NLW_blk00000001/blk0000039d_DOB<18>_UNCONNECTED ,
\NLW_blk00000001/blk0000039d_DOB<17>_UNCONNECTED , \NLW_blk00000001/blk0000039d_DOB<16>_UNCONNECTED , \blk00000001/sig000001db ,
\blk00000001/sig000001da , \blk00000001/sig000001d9 , \blk00000001/sig000001d8 , \blk00000001/sig000001d7 , \blk00000001/sig000001d6 ,
\blk00000001/sig000001d5 , \blk00000001/sig000001d4 , \blk00000001/sig000001d3 , \blk00000001/sig000001d2 , \blk00000001/sig000001d1 ,
\blk00000001/sig000001d0 , \blk00000001/sig000001cf , \blk00000001/sig000001ce , \blk00000001/sig000001cd , \blk00000001/sig000001cc }),
    .WEB({\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d }),
    .DIA({\NLW_blk00000001/blk0000039d_DIA<31>_UNCONNECTED , \NLW_blk00000001/blk0000039d_DIA<30>_UNCONNECTED ,
\NLW_blk00000001/blk0000039d_DIA<29>_UNCONNECTED , \NLW_blk00000001/blk0000039d_DIA<28>_UNCONNECTED ,
\NLW_blk00000001/blk0000039d_DIA<27>_UNCONNECTED , \NLW_blk00000001/blk0000039d_DIA<26>_UNCONNECTED ,
\NLW_blk00000001/blk0000039d_DIA<25>_UNCONNECTED , \NLW_blk00000001/blk0000039d_DIA<24>_UNCONNECTED ,
\NLW_blk00000001/blk0000039d_DIA<23>_UNCONNECTED , \NLW_blk00000001/blk0000039d_DIA<22>_UNCONNECTED ,
\NLW_blk00000001/blk0000039d_DIA<21>_UNCONNECTED , \NLW_blk00000001/blk0000039d_DIA<20>_UNCONNECTED ,
\NLW_blk00000001/blk0000039d_DIA<19>_UNCONNECTED , \NLW_blk00000001/blk0000039d_DIA<18>_UNCONNECTED ,
\NLW_blk00000001/blk0000039d_DIA<17>_UNCONNECTED , \NLW_blk00000001/blk0000039d_DIA<16>_UNCONNECTED , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d })
  );
  INV   \blk00000001/blk0000039c  (
    .I(\blk00000001/sig00000040 ),
    .O(\blk00000001/sig0000055b )
  );
  INV   \blk00000001/blk0000039b  (
    .I(\blk00000001/sig0000006e ),
    .O(\blk00000001/sig0000026c )
  );
  INV   \blk00000001/blk0000039a  (
    .I(\blk00000001/sig0000006d ),
    .O(\blk00000001/sig0000026b )
  );
  INV   \blk00000001/blk00000399  (
    .I(\blk00000001/sig0000006c ),
    .O(\blk00000001/sig0000026a )
  );
  INV   \blk00000001/blk00000398  (
    .I(\blk00000001/sig0000006b ),
    .O(\blk00000001/sig00000269 )
  );
  INV   \blk00000001/blk00000397  (
    .I(\blk00000001/sig0000006a ),
    .O(\blk00000001/sig00000268 )
  );
  INV   \blk00000001/blk00000396  (
    .I(\blk00000001/sig000000ac ),
    .O(\blk00000001/sig00000194 )
  );
  INV   \blk00000001/blk00000395  (
    .I(\blk00000001/sig0000003d ),
    .O(NlwRenamedSignal_s_axis_dividend_tready)
  );
  LUT4 #(
    .INIT ( 16'hA280 ))
  \blk00000001/blk00000394  (
    .I0(\blk00000001/sig0000006b ),
    .I1(\blk00000001/sig0000006a ),
    .I2(\blk00000001/sig0000009f ),
    .I3(\blk00000001/sig0000009e ),
    .O(\blk00000001/sig00000229 )
  );
  LUT5 #(
    .INIT ( 32'hFBEA5140 ))
  \blk00000001/blk00000393  (
    .I0(\blk00000001/sig0000006b ),
    .I1(\blk00000001/sig0000006a ),
    .I2(\blk00000001/sig000000a9 ),
    .I3(\blk00000001/sig000000a8 ),
    .I4(\blk00000001/sig00000237 ),
    .O(\blk00000001/sig00000235 )
  );
  LUT3 #(
    .INIT ( 8'h80 ))
  \blk00000001/blk00000392  (
    .I0(\blk00000001/sig0000006b ),
    .I1(\blk00000001/sig0000006a ),
    .I2(\blk00000001/sig0000009e ),
    .O(\blk00000001/sig00000228 )
  );
  LUT4 #(
    .INIT ( 16'h5410 ))
  \blk00000001/blk00000391  (
    .I0(\blk00000001/sig00000256 ),
    .I1(\blk00000001/sig00000258 ),
    .I2(\blk00000001/sig00000260 ),
    .I3(\blk00000001/sig0000025c ),
    .O(\blk00000001/sig00000213 )
  );
  LUT4 #(
    .INIT ( 16'h5410 ))
  \blk00000001/blk00000390  (
    .I0(\blk00000001/sig00000256 ),
    .I1(\blk00000001/sig00000258 ),
    .I2(\blk00000001/sig0000025f ),
    .I3(\blk00000001/sig0000025b ),
    .O(\blk00000001/sig00000212 )
  );
  LUT4 #(
    .INIT ( 16'h5410 ))
  \blk00000001/blk0000038f  (
    .I0(\blk00000001/sig00000256 ),
    .I1(\blk00000001/sig00000258 ),
    .I2(\blk00000001/sig0000025e ),
    .I3(\blk00000001/sig0000025a ),
    .O(\blk00000001/sig00000211 )
  );
  LUT4 #(
    .INIT ( 16'h5410 ))
  \blk00000001/blk0000038e  (
    .I0(\blk00000001/sig00000256 ),
    .I1(\blk00000001/sig00000258 ),
    .I2(\blk00000001/sig0000025d ),
    .I3(\blk00000001/sig00000259 ),
    .O(\blk00000001/sig00000210 )
  );
  LUT3 #(
    .INIT ( 8'h10 ))
  \blk00000001/blk0000038d  (
    .I0(\blk00000001/sig00000256 ),
    .I1(\blk00000001/sig00000258 ),
    .I2(\blk00000001/sig0000025c ),
    .O(\blk00000001/sig0000020f )
  );
  LUT3 #(
    .INIT ( 8'h10 ))
  \blk00000001/blk0000038c  (
    .I0(\blk00000001/sig00000256 ),
    .I1(\blk00000001/sig00000258 ),
    .I2(\blk00000001/sig0000025b ),
    .O(\blk00000001/sig0000020e )
  );
  LUT5 #(
    .INIT ( 32'hFD75A820 ))
  \blk00000001/blk0000038b  (
    .I0(\blk00000001/sig00000256 ),
    .I1(\blk00000001/sig00000258 ),
    .I2(\blk00000001/sig00000267 ),
    .I3(\blk00000001/sig00000263 ),
    .I4(\blk00000001/sig00000227 ),
    .O(\blk00000001/sig00000222 )
  );
  LUT5 #(
    .INIT ( 32'hFD75A820 ))
  \blk00000001/blk0000038a  (
    .I0(\blk00000001/sig00000256 ),
    .I1(\blk00000001/sig00000258 ),
    .I2(\blk00000001/sig00000266 ),
    .I3(\blk00000001/sig00000262 ),
    .I4(\blk00000001/sig00000227 ),
    .O(\blk00000001/sig00000221 )
  );
  LUT5 #(
    .INIT ( 32'hFD75A820 ))
  \blk00000001/blk00000389  (
    .I0(\blk00000001/sig00000256 ),
    .I1(\blk00000001/sig00000258 ),
    .I2(\blk00000001/sig00000265 ),
    .I3(\blk00000001/sig00000261 ),
    .I4(\blk00000001/sig00000227 ),
    .O(\blk00000001/sig00000220 )
  );
  LUT3 #(
    .INIT ( 8'h10 ))
  \blk00000001/blk00000388  (
    .I0(\blk00000001/sig00000256 ),
    .I1(\blk00000001/sig00000258 ),
    .I2(\blk00000001/sig0000025a ),
    .O(\blk00000001/sig0000020d )
  );
  LUT5 #(
    .INIT ( 32'hFD75A820 ))
  \blk00000001/blk00000387  (
    .I0(\blk00000001/sig00000256 ),
    .I1(\blk00000001/sig00000258 ),
    .I2(\blk00000001/sig00000264 ),
    .I3(\blk00000001/sig00000260 ),
    .I4(\blk00000001/sig00000227 ),
    .O(\blk00000001/sig0000021f )
  );
  LUT3 #(
    .INIT ( 8'h10 ))
  \blk00000001/blk00000386  (
    .I0(\blk00000001/sig00000256 ),
    .I1(\blk00000001/sig00000258 ),
    .I2(\blk00000001/sig00000259 ),
    .O(\blk00000001/sig0000020c )
  );
  LUT4 #(
    .INIT ( 16'hABA8 ))
  \blk00000001/blk00000385  (
    .I0(\blk00000001/sig00000237 ),
    .I1(\blk00000001/sig0000006b ),
    .I2(\blk00000001/sig0000006a ),
    .I3(\blk00000001/sig000000a9 ),
    .O(\blk00000001/sig00000236 )
  );
  LUT4 #(
    .INIT ( 16'hEA2A ))
  \blk00000001/blk00000384  (
    .I0(\blk00000001/sig00000227 ),
    .I1(\blk00000001/sig00000256 ),
    .I2(\blk00000001/sig00000258 ),
    .I3(\blk00000001/sig00000267 ),
    .O(\blk00000001/sig00000226 )
  );
  LUT4 #(
    .INIT ( 16'hEA2A ))
  \blk00000001/blk00000383  (
    .I0(\blk00000001/sig00000227 ),
    .I1(\blk00000001/sig00000256 ),
    .I2(\blk00000001/sig00000258 ),
    .I3(\blk00000001/sig00000266 ),
    .O(\blk00000001/sig00000225 )
  );
  LUT4 #(
    .INIT ( 16'hEA2A ))
  \blk00000001/blk00000382  (
    .I0(\blk00000001/sig00000227 ),
    .I1(\blk00000001/sig00000256 ),
    .I2(\blk00000001/sig00000258 ),
    .I3(\blk00000001/sig00000265 ),
    .O(\blk00000001/sig00000224 )
  );
  LUT4 #(
    .INIT ( 16'hEA2A ))
  \blk00000001/blk00000381  (
    .I0(\blk00000001/sig00000227 ),
    .I1(\blk00000001/sig00000256 ),
    .I2(\blk00000001/sig00000258 ),
    .I3(\blk00000001/sig00000264 ),
    .O(\blk00000001/sig00000223 )
  );
  LUT6 #(
    .INIT ( 64'h5410FEBA54105410 ))
  \blk00000001/blk00000380  (
    .I0(\blk00000001/sig000000cf ),
    .I1(\blk00000001/sig00000127 ),
    .I2(\blk00000001/sig000000d8 ),
    .I3(\blk00000001/sig000000d4 ),
    .I4(\blk00000001/sig00000126 ),
    .I5(\blk00000001/sig000000d0 ),
    .O(\blk00000001/sig00000145 )
  );
  LUT6 #(
    .INIT ( 64'h5410FEBA54105410 ))
  \blk00000001/blk0000037f  (
    .I0(\blk00000001/sig000000cf ),
    .I1(\blk00000001/sig00000127 ),
    .I2(\blk00000001/sig000000d9 ),
    .I3(\blk00000001/sig000000d5 ),
    .I4(\blk00000001/sig00000126 ),
    .I5(\blk00000001/sig000000d1 ),
    .O(\blk00000001/sig00000144 )
  );
  LUT6 #(
    .INIT ( 64'h5410FEBA54105410 ))
  \blk00000001/blk0000037e  (
    .I0(\blk00000001/sig000000cf ),
    .I1(\blk00000001/sig00000127 ),
    .I2(\blk00000001/sig000000da ),
    .I3(\blk00000001/sig000000d6 ),
    .I4(\blk00000001/sig00000126 ),
    .I5(\blk00000001/sig000000d2 ),
    .O(\blk00000001/sig00000143 )
  );
  LUT6 #(
    .INIT ( 64'h5410FEBA54105410 ))
  \blk00000001/blk0000037d  (
    .I0(\blk00000001/sig000000cf ),
    .I1(\blk00000001/sig00000127 ),
    .I2(\blk00000001/sig000000db ),
    .I3(\blk00000001/sig000000d7 ),
    .I4(\blk00000001/sig00000126 ),
    .I5(\blk00000001/sig000000d3 ),
    .O(\blk00000001/sig00000142 )
  );
  LUT3 #(
    .INIT ( 8'h10 ))
  \blk00000001/blk0000037c  (
    .I0(\blk00000001/sig000000cf ),
    .I1(\blk00000001/sig00000127 ),
    .I2(\blk00000001/sig000000d0 ),
    .O(\blk00000001/sig0000014d )
  );
  LUT3 #(
    .INIT ( 8'h10 ))
  \blk00000001/blk0000037b  (
    .I0(\blk00000001/sig000000cf ),
    .I1(\blk00000001/sig00000127 ),
    .I2(\blk00000001/sig000000d1 ),
    .O(\blk00000001/sig0000014c )
  );
  LUT3 #(
    .INIT ( 8'h10 ))
  \blk00000001/blk0000037a  (
    .I0(\blk00000001/sig000000cf ),
    .I1(\blk00000001/sig00000127 ),
    .I2(\blk00000001/sig000000d2 ),
    .O(\blk00000001/sig0000014b )
  );
  LUT3 #(
    .INIT ( 8'h10 ))
  \blk00000001/blk00000379  (
    .I0(\blk00000001/sig000000cf ),
    .I1(\blk00000001/sig00000127 ),
    .I2(\blk00000001/sig000000d3 ),
    .O(\blk00000001/sig0000014a )
  );
  LUT4 #(
    .INIT ( 16'h5410 ))
  \blk00000001/blk00000378  (
    .I0(\blk00000001/sig000000cf ),
    .I1(\blk00000001/sig00000127 ),
    .I2(\blk00000001/sig000000d6 ),
    .I3(\blk00000001/sig000000d2 ),
    .O(\blk00000001/sig00000147 )
  );
  LUT4 #(
    .INIT ( 16'h5410 ))
  \blk00000001/blk00000377  (
    .I0(\blk00000001/sig000000cf ),
    .I1(\blk00000001/sig00000127 ),
    .I2(\blk00000001/sig000000d7 ),
    .I3(\blk00000001/sig000000d3 ),
    .O(\blk00000001/sig00000146 )
  );
  LUT4 #(
    .INIT ( 16'h5410 ))
  \blk00000001/blk00000376  (
    .I0(\blk00000001/sig000000cf ),
    .I1(\blk00000001/sig00000127 ),
    .I2(\blk00000001/sig000000d4 ),
    .I3(\blk00000001/sig000000d0 ),
    .O(\blk00000001/sig00000149 )
  );
  LUT4 #(
    .INIT ( 16'h5410 ))
  \blk00000001/blk00000375  (
    .I0(\blk00000001/sig000000cf ),
    .I1(\blk00000001/sig00000127 ),
    .I2(\blk00000001/sig000000d5 ),
    .I3(\blk00000001/sig000000d1 ),
    .O(\blk00000001/sig00000148 )
  );
  LUT4 #(
    .INIT ( 16'hE444 ))
  \blk00000001/blk00000374  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig000004b3 ),
    .I2(\blk00000001/sig0000008a ),
    .I3(\blk00000001/sig00000069 ),
    .O(\blk00000001/sig000002bf )
  );
  LUT4 #(
    .INIT ( 16'hE444 ))
  \blk00000001/blk00000373  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig000004b2 ),
    .I2(\blk00000001/sig0000008a ),
    .I3(\blk00000001/sig00000069 ),
    .O(\blk00000001/sig000002be )
  );
  LUT4 #(
    .INIT ( 16'hE444 ))
  \blk00000001/blk00000372  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig000004b1 ),
    .I2(\blk00000001/sig0000008a ),
    .I3(\blk00000001/sig00000069 ),
    .O(\blk00000001/sig000002bd )
  );
  LUT4 #(
    .INIT ( 16'hE444 ))
  \blk00000001/blk00000371  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig000004b0 ),
    .I2(\blk00000001/sig0000008a ),
    .I3(\blk00000001/sig00000069 ),
    .O(\blk00000001/sig000002bc )
  );
  LUT4 #(
    .INIT ( 16'hE444 ))
  \blk00000001/blk00000370  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig000004af ),
    .I2(\blk00000001/sig0000008a ),
    .I3(\blk00000001/sig00000069 ),
    .O(\blk00000001/sig000002bb )
  );
  LUT4 #(
    .INIT ( 16'hE444 ))
  \blk00000001/blk0000036f  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig000004ae ),
    .I2(\blk00000001/sig0000008a ),
    .I3(\blk00000001/sig00000069 ),
    .O(\blk00000001/sig000002ba )
  );
  LUT4 #(
    .INIT ( 16'hE444 ))
  \blk00000001/blk0000036e  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig000004ad ),
    .I2(\blk00000001/sig0000008a ),
    .I3(\blk00000001/sig00000069 ),
    .O(\blk00000001/sig000002b9 )
  );
  LUT4 #(
    .INIT ( 16'hE444 ))
  \blk00000001/blk0000036d  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig000004ac ),
    .I2(\blk00000001/sig0000008a ),
    .I3(\blk00000001/sig00000069 ),
    .O(\blk00000001/sig000002b8 )
  );
  LUT4 #(
    .INIT ( 16'hE444 ))
  \blk00000001/blk0000036c  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig000004ab ),
    .I2(\blk00000001/sig0000008a ),
    .I3(\blk00000001/sig00000069 ),
    .O(\blk00000001/sig000002b7 )
  );
  LUT4 #(
    .INIT ( 16'hE444 ))
  \blk00000001/blk0000036b  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig000004aa ),
    .I2(\blk00000001/sig0000008a ),
    .I3(\blk00000001/sig00000069 ),
    .O(\blk00000001/sig000002b6 )
  );
  LUT4 #(
    .INIT ( 16'hE444 ))
  \blk00000001/blk0000036a  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig000004a9 ),
    .I2(\blk00000001/sig0000008a ),
    .I3(\blk00000001/sig00000069 ),
    .O(\blk00000001/sig000002b5 )
  );
  LUT4 #(
    .INIT ( 16'hE444 ))
  \blk00000001/blk00000369  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig000004a8 ),
    .I2(\blk00000001/sig0000008a ),
    .I3(\blk00000001/sig00000069 ),
    .O(\blk00000001/sig000002b4 )
  );
  LUT4 #(
    .INIT ( 16'hE444 ))
  \blk00000001/blk00000368  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig000004a7 ),
    .I2(\blk00000001/sig0000008a ),
    .I3(\blk00000001/sig00000069 ),
    .O(\blk00000001/sig000002b3 )
  );
  LUT4 #(
    .INIT ( 16'hE444 ))
  \blk00000001/blk00000367  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig000004a6 ),
    .I2(\blk00000001/sig0000008a ),
    .I3(\blk00000001/sig00000069 ),
    .O(\blk00000001/sig000002b2 )
  );
  LUT4 #(
    .INIT ( 16'hE444 ))
  \blk00000001/blk00000366  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig000004a5 ),
    .I2(\blk00000001/sig0000008a ),
    .I3(\blk00000001/sig00000069 ),
    .O(\blk00000001/sig000002b1 )
  );
  LUT4 #(
    .INIT ( 16'hE444 ))
  \blk00000001/blk00000365  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig000004a4 ),
    .I2(\blk00000001/sig0000008a ),
    .I3(\blk00000001/sig00000069 ),
    .O(\blk00000001/sig000002b0 )
  );
  LUT6 #(
    .INIT ( 64'hFD75EC64B931A820 ))
  \blk00000001/blk00000364  (
    .I0(\blk00000001/sig0000006a ),
    .I1(\blk00000001/sig0000006b ),
    .I2(\blk00000001/sig000000a5 ),
    .I3(\blk00000001/sig000000a7 ),
    .I4(\blk00000001/sig000000a4 ),
    .I5(\blk00000001/sig000000a6 ),
    .O(\blk00000001/sig00000231 )
  );
  LUT6 #(
    .INIT ( 64'hFD75EC64B931A820 ))
  \blk00000001/blk00000363  (
    .I0(\blk00000001/sig0000006a ),
    .I1(\blk00000001/sig0000006b ),
    .I2(\blk00000001/sig000000a4 ),
    .I3(\blk00000001/sig000000a6 ),
    .I4(\blk00000001/sig000000a3 ),
    .I5(\blk00000001/sig000000a5 ),
    .O(\blk00000001/sig00000230 )
  );
  LUT6 #(
    .INIT ( 64'hFD75EC64B931A820 ))
  \blk00000001/blk00000362  (
    .I0(\blk00000001/sig0000006a ),
    .I1(\blk00000001/sig0000006b ),
    .I2(\blk00000001/sig000000a3 ),
    .I3(\blk00000001/sig000000a5 ),
    .I4(\blk00000001/sig000000a2 ),
    .I5(\blk00000001/sig000000a4 ),
    .O(\blk00000001/sig0000022f )
  );
  LUT6 #(
    .INIT ( 64'hFD75EC64B931A820 ))
  \blk00000001/blk00000361  (
    .I0(\blk00000001/sig0000006a ),
    .I1(\blk00000001/sig0000006b ),
    .I2(\blk00000001/sig000000a2 ),
    .I3(\blk00000001/sig000000a4 ),
    .I4(\blk00000001/sig000000a1 ),
    .I5(\blk00000001/sig000000a3 ),
    .O(\blk00000001/sig0000022e )
  );
  LUT6 #(
    .INIT ( 64'hFD75EC64B931A820 ))
  \blk00000001/blk00000360  (
    .I0(\blk00000001/sig0000006a ),
    .I1(\blk00000001/sig0000006b ),
    .I2(\blk00000001/sig000000a1 ),
    .I3(\blk00000001/sig000000a3 ),
    .I4(\blk00000001/sig000000a0 ),
    .I5(\blk00000001/sig000000a2 ),
    .O(\blk00000001/sig0000022d )
  );
  LUT6 #(
    .INIT ( 64'hFD75EC64B931A820 ))
  \blk00000001/blk0000035f  (
    .I0(\blk00000001/sig0000006a ),
    .I1(\blk00000001/sig0000006b ),
    .I2(\blk00000001/sig000000a0 ),
    .I3(\blk00000001/sig000000a2 ),
    .I4(\blk00000001/sig0000009f ),
    .I5(\blk00000001/sig000000a1 ),
    .O(\blk00000001/sig0000022c )
  );
  LUT6 #(
    .INIT ( 64'hFD75EC64B931A820 ))
  \blk00000001/blk0000035e  (
    .I0(\blk00000001/sig0000006a ),
    .I1(\blk00000001/sig0000006b ),
    .I2(\blk00000001/sig0000009f ),
    .I3(\blk00000001/sig000000a1 ),
    .I4(\blk00000001/sig0000009e ),
    .I5(\blk00000001/sig000000a0 ),
    .O(\blk00000001/sig0000022b )
  );
  LUT5 #(
    .INIT ( 32'hEC64A820 ))
  \blk00000001/blk0000035d  (
    .I0(\blk00000001/sig0000006a ),
    .I1(\blk00000001/sig0000006b ),
    .I2(\blk00000001/sig0000009e ),
    .I3(\blk00000001/sig000000a0 ),
    .I4(\blk00000001/sig0000009f ),
    .O(\blk00000001/sig0000022a )
  );
  LUT6 #(
    .INIT ( 64'hFD75EC64B931A820 ))
  \blk00000001/blk0000035c  (
    .I0(\blk00000001/sig0000006a ),
    .I1(\blk00000001/sig0000006b ),
    .I2(\blk00000001/sig000000a8 ),
    .I3(\blk00000001/sig00000237 ),
    .I4(\blk00000001/sig000000a7 ),
    .I5(\blk00000001/sig000000a9 ),
    .O(\blk00000001/sig00000234 )
  );
  LUT6 #(
    .INIT ( 64'hFD75EC64B931A820 ))
  \blk00000001/blk0000035b  (
    .I0(\blk00000001/sig0000006a ),
    .I1(\blk00000001/sig0000006b ),
    .I2(\blk00000001/sig000000a7 ),
    .I3(\blk00000001/sig000000a9 ),
    .I4(\blk00000001/sig000000a6 ),
    .I5(\blk00000001/sig000000a8 ),
    .O(\blk00000001/sig00000233 )
  );
  LUT6 #(
    .INIT ( 64'hFD75EC64B931A820 ))
  \blk00000001/blk0000035a  (
    .I0(\blk00000001/sig0000006a ),
    .I1(\blk00000001/sig0000006b ),
    .I2(\blk00000001/sig000000a6 ),
    .I3(\blk00000001/sig000000a8 ),
    .I4(\blk00000001/sig000000a5 ),
    .I5(\blk00000001/sig000000a7 ),
    .O(\blk00000001/sig00000232 )
  );
  LUT5 #(
    .INIT ( 32'h73625140 ))
  \blk00000001/blk00000359  (
    .I0(\blk00000001/sig00000256 ),
    .I1(\blk00000001/sig00000258 ),
    .I2(\blk00000001/sig0000025e ),
    .I3(\blk00000001/sig00000262 ),
    .I4(\blk00000001/sig0000025a ),
    .O(\blk00000001/sig00000215 )
  );
  LUT5 #(
    .INIT ( 32'h73625140 ))
  \blk00000001/blk00000358  (
    .I0(\blk00000001/sig00000256 ),
    .I1(\blk00000001/sig00000258 ),
    .I2(\blk00000001/sig0000025d ),
    .I3(\blk00000001/sig00000261 ),
    .I4(\blk00000001/sig00000259 ),
    .O(\blk00000001/sig00000214 )
  );
  LUT6 #(
    .INIT ( 64'hFD75EC64B931A820 ))
  \blk00000001/blk00000357  (
    .I0(\blk00000001/sig00000258 ),
    .I1(\blk00000001/sig00000256 ),
    .I2(\blk00000001/sig00000267 ),
    .I3(\blk00000001/sig0000025f ),
    .I4(\blk00000001/sig00000227 ),
    .I5(\blk00000001/sig00000263 ),
    .O(\blk00000001/sig0000021e )
  );
  LUT6 #(
    .INIT ( 64'hFD75EC64B931A820 ))
  \blk00000001/blk00000356  (
    .I0(\blk00000001/sig00000258 ),
    .I1(\blk00000001/sig00000256 ),
    .I2(\blk00000001/sig00000266 ),
    .I3(\blk00000001/sig0000025e ),
    .I4(\blk00000001/sig00000227 ),
    .I5(\blk00000001/sig00000262 ),
    .O(\blk00000001/sig0000021d )
  );
  LUT6 #(
    .INIT ( 64'hFD75EC64B931A820 ))
  \blk00000001/blk00000355  (
    .I0(\blk00000001/sig00000258 ),
    .I1(\blk00000001/sig00000256 ),
    .I2(\blk00000001/sig00000265 ),
    .I3(\blk00000001/sig0000025d ),
    .I4(\blk00000001/sig00000227 ),
    .I5(\blk00000001/sig00000261 ),
    .O(\blk00000001/sig0000021c )
  );
  LUT6 #(
    .INIT ( 64'hFD75EC64B931A820 ))
  \blk00000001/blk00000354  (
    .I0(\blk00000001/sig00000258 ),
    .I1(\blk00000001/sig00000256 ),
    .I2(\blk00000001/sig00000264 ),
    .I3(\blk00000001/sig0000025c ),
    .I4(\blk00000001/sig00000227 ),
    .I5(\blk00000001/sig00000260 ),
    .O(\blk00000001/sig0000021b )
  );
  LUT6 #(
    .INIT ( 64'hFD75EC64B931A820 ))
  \blk00000001/blk00000353  (
    .I0(\blk00000001/sig00000258 ),
    .I1(\blk00000001/sig00000256 ),
    .I2(\blk00000001/sig00000263 ),
    .I3(\blk00000001/sig0000025b ),
    .I4(\blk00000001/sig00000267 ),
    .I5(\blk00000001/sig0000025f ),
    .O(\blk00000001/sig0000021a )
  );
  LUT6 #(
    .INIT ( 64'hFD75EC64B931A820 ))
  \blk00000001/blk00000352  (
    .I0(\blk00000001/sig00000258 ),
    .I1(\blk00000001/sig00000256 ),
    .I2(\blk00000001/sig00000262 ),
    .I3(\blk00000001/sig0000025a ),
    .I4(\blk00000001/sig00000266 ),
    .I5(\blk00000001/sig0000025e ),
    .O(\blk00000001/sig00000219 )
  );
  LUT6 #(
    .INIT ( 64'hFD75EC64B931A820 ))
  \blk00000001/blk00000351  (
    .I0(\blk00000001/sig00000258 ),
    .I1(\blk00000001/sig00000256 ),
    .I2(\blk00000001/sig00000261 ),
    .I3(\blk00000001/sig00000259 ),
    .I4(\blk00000001/sig00000265 ),
    .I5(\blk00000001/sig0000025d ),
    .O(\blk00000001/sig00000218 )
  );
  LUT5 #(
    .INIT ( 32'h73625140 ))
  \blk00000001/blk00000350  (
    .I0(\blk00000001/sig00000256 ),
    .I1(\blk00000001/sig00000258 ),
    .I2(\blk00000001/sig00000260 ),
    .I3(\blk00000001/sig00000264 ),
    .I4(\blk00000001/sig0000025c ),
    .O(\blk00000001/sig00000217 )
  );
  LUT5 #(
    .INIT ( 32'h73625140 ))
  \blk00000001/blk0000034f  (
    .I0(\blk00000001/sig00000256 ),
    .I1(\blk00000001/sig00000258 ),
    .I2(\blk00000001/sig0000025f ),
    .I3(\blk00000001/sig00000263 ),
    .I4(\blk00000001/sig0000025b ),
    .O(\blk00000001/sig00000216 )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk00000001/blk0000034e  (
    .I0(\blk00000001/sig0000015b ),
    .O(\blk00000001/sig0000056d )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk00000001/blk0000034d  (
    .I0(\blk00000001/sig0000015c ),
    .O(\blk00000001/sig0000056c )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk00000001/blk0000034c  (
    .I0(\blk00000001/sig0000015d ),
    .O(\blk00000001/sig0000056b )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk00000001/blk0000034b  (
    .I0(\blk00000001/sig0000015e ),
    .O(\blk00000001/sig0000056a )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk00000001/blk0000034a  (
    .I0(\blk00000001/sig0000015f ),
    .O(\blk00000001/sig00000569 )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk00000001/blk00000349  (
    .I0(\blk00000001/sig00000160 ),
    .O(\blk00000001/sig00000568 )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk00000001/blk00000348  (
    .I0(\blk00000001/sig00000161 ),
    .O(\blk00000001/sig00000567 )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk00000001/blk00000347  (
    .I0(\blk00000001/sig00000162 ),
    .O(\blk00000001/sig00000566 )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk00000001/blk00000346  (
    .I0(\blk00000001/sig00000163 ),
    .O(\blk00000001/sig00000565 )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk00000001/blk00000345  (
    .I0(\blk00000001/sig00000164 ),
    .O(\blk00000001/sig00000564 )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk00000001/blk00000344  (
    .I0(\blk00000001/sig00000165 ),
    .O(\blk00000001/sig00000563 )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk00000001/blk00000343  (
    .I0(\blk00000001/sig00000166 ),
    .O(\blk00000001/sig00000562 )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk00000001/blk00000342  (
    .I0(\blk00000001/sig0000016b ),
    .O(\blk00000001/sig00000561 )
  );
  FD   \blk00000001/blk00000341  (
    .C(aclk),
    .D(\blk00000001/sig000000f7 ),
    .Q(\blk00000001/sig000000b6 )
  );
  FD   \blk00000001/blk00000340  (
    .C(aclk),
    .D(\blk00000001/sig000000f8 ),
    .Q(\blk00000001/sig000000b7 )
  );
  FD   \blk00000001/blk0000033f  (
    .C(aclk),
    .D(\blk00000001/sig000000f9 ),
    .Q(\blk00000001/sig000000b8 )
  );
  FD   \blk00000001/blk0000033e  (
    .C(aclk),
    .D(\blk00000001/sig000000fa ),
    .Q(\blk00000001/sig000000b9 )
  );
  FD   \blk00000001/blk0000033d  (
    .C(aclk),
    .D(\blk00000001/sig000000fb ),
    .Q(\blk00000001/sig000000ba )
  );
  LUT6 #(
    .INIT ( 64'h0404040037373733 ))
  \blk00000001/blk0000033c  (
    .I0(\blk00000001/sig000000d9 ),
    .I1(\blk00000001/sig00000127 ),
    .I2(\blk00000001/sig000000d8 ),
    .I3(\blk00000001/sig000000d6 ),
    .I4(\blk00000001/sig000000d7 ),
    .I5(\blk00000001/sig00000560 ),
    .O(\blk00000001/sig00000130 )
  );
  LUT3 #(
    .INIT ( 8'hF1 ))
  \blk00000001/blk0000033b  (
    .I0(\blk00000001/sig000000db ),
    .I1(\blk00000001/sig000000da ),
    .I2(\blk00000001/sig000000dc ),
    .O(\blk00000001/sig00000560 )
  );
  LUT6 #(
    .INIT ( 64'h2222020077775755 ))
  \blk00000001/blk0000033a  (
    .I0(\blk00000001/sig00000127 ),
    .I1(\blk00000001/sig000000d9 ),
    .I2(\blk00000001/sig000000d7 ),
    .I3(\blk00000001/sig000000d6 ),
    .I4(\blk00000001/sig000000d8 ),
    .I5(\blk00000001/sig0000055f ),
    .O(\blk00000001/sig00000131 )
  );
  LUT3 #(
    .INIT ( 8'h45 ))
  \blk00000001/blk00000339  (
    .I0(\blk00000001/sig000000dc ),
    .I1(\blk00000001/sig000000db ),
    .I2(\blk00000001/sig000000da ),
    .O(\blk00000001/sig0000055f )
  );
  LUT6 #(
    .INIT ( 64'h10111010DCDDDCDC ))
  \blk00000001/blk00000338  (
    .I0(\blk00000001/sig000000d5 ),
    .I1(\blk00000001/sig00000126 ),
    .I2(\blk00000001/sig000000d4 ),
    .I3(\blk00000001/sig000000d3 ),
    .I4(\blk00000001/sig000000d2 ),
    .I5(\blk00000001/sig0000055e ),
    .O(\blk00000001/sig0000012f )
  );
  LUT2 #(
    .INIT ( 4'hB ))
  \blk00000001/blk00000337  (
    .I0(\blk00000001/sig000000d1 ),
    .I1(\blk00000001/sig000000d0 ),
    .O(\blk00000001/sig0000055e )
  );
  LUT6 #(
    .INIT ( 64'h4444441444444444 ))
  \blk00000001/blk00000336  (
    .I0(\blk00000001/sig000000fc ),
    .I1(\blk00000001/sig00000101 ),
    .I2(\blk00000001/sig000000fd ),
    .I3(\blk00000001/sig00000167 ),
    .I4(\blk00000001/sig0000055d ),
    .I5(\blk00000001/sig000000fe ),
    .O(\blk00000001/sig000000fb )
  );
  LUT2 #(
    .INIT ( 4'h7 ))
  \blk00000001/blk00000335  (
    .I0(\blk00000001/sig00000100 ),
    .I1(\blk00000001/sig000000ff ),
    .O(\blk00000001/sig0000055d )
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  \blk00000001/blk00000334  (
    .I0(\blk00000001/sig00000040 ),
    .I1(\blk00000001/sig00000546 ),
    .I2(\blk00000001/sig0000009d ),
    .O(\blk00000001/sig00000545 )
  );
  LUT2 #(
    .INIT ( 4'hB ))
  \blk00000001/blk00000333  (
    .I0(\blk00000001/sig0000009c ),
    .I1(\blk00000001/sig0000003c ),
    .O(\blk00000001/sig0000031c )
  );
  LUT3 #(
    .INIT ( 8'h80 ))
  \blk00000001/blk00000332  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig0000008a ),
    .I2(\blk00000001/sig00000063 ),
    .O(\blk00000001/sig000002aa )
  );
  LUT3 #(
    .INIT ( 8'h80 ))
  \blk00000001/blk00000331  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig0000008a ),
    .I2(\blk00000001/sig00000062 ),
    .O(\blk00000001/sig000002a9 )
  );
  LUT3 #(
    .INIT ( 8'h80 ))
  \blk00000001/blk00000330  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig0000008a ),
    .I2(\blk00000001/sig00000061 ),
    .O(\blk00000001/sig000002a8 )
  );
  LUT3 #(
    .INIT ( 8'h80 ))
  \blk00000001/blk0000032f  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig0000008a ),
    .I2(\blk00000001/sig00000060 ),
    .O(\blk00000001/sig000002a7 )
  );
  LUT3 #(
    .INIT ( 8'h80 ))
  \blk00000001/blk0000032e  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig0000008a ),
    .I2(\blk00000001/sig0000005f ),
    .O(\blk00000001/sig000002a6 )
  );
  LUT3 #(
    .INIT ( 8'h80 ))
  \blk00000001/blk0000032d  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig0000008a ),
    .I2(\blk00000001/sig0000005e ),
    .O(\blk00000001/sig000002a5 )
  );
  LUT3 #(
    .INIT ( 8'h80 ))
  \blk00000001/blk0000032c  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig0000008a ),
    .I2(\blk00000001/sig0000005d ),
    .O(\blk00000001/sig000002a4 )
  );
  LUT3 #(
    .INIT ( 8'h80 ))
  \blk00000001/blk0000032b  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig0000008a ),
    .I2(\blk00000001/sig0000005c ),
    .O(\blk00000001/sig000002a3 )
  );
  LUT3 #(
    .INIT ( 8'h80 ))
  \blk00000001/blk0000032a  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig0000008a ),
    .I2(\blk00000001/sig0000005b ),
    .O(\blk00000001/sig000002a2 )
  );
  LUT3 #(
    .INIT ( 8'h80 ))
  \blk00000001/blk00000329  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig0000008a ),
    .I2(\blk00000001/sig00000068 ),
    .O(\blk00000001/sig000002af )
  );
  LUT3 #(
    .INIT ( 8'h80 ))
  \blk00000001/blk00000328  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig0000008a ),
    .I2(\blk00000001/sig00000067 ),
    .O(\blk00000001/sig000002ae )
  );
  LUT3 #(
    .INIT ( 8'h80 ))
  \blk00000001/blk00000327  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig0000008a ),
    .I2(\blk00000001/sig00000066 ),
    .O(\blk00000001/sig000002ad )
  );
  LUT3 #(
    .INIT ( 8'h80 ))
  \blk00000001/blk00000326  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig0000008a ),
    .I2(\blk00000001/sig00000065 ),
    .O(\blk00000001/sig000002ac )
  );
  LUT3 #(
    .INIT ( 8'h80 ))
  \blk00000001/blk00000325  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig0000008a ),
    .I2(\blk00000001/sig00000064 ),
    .O(\blk00000001/sig000002ab )
  );
  LUT3 #(
    .INIT ( 8'h80 ))
  \blk00000001/blk00000324  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig0000008a ),
    .I2(\blk00000001/sig0000005a ),
    .O(\blk00000001/sig000002a1 )
  );
  LUT2 #(
    .INIT ( 4'h8 ))
  \blk00000001/blk00000323  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig00000053 ),
    .O(\blk00000001/sig000002f5 )
  );
  LUT2 #(
    .INIT ( 4'h8 ))
  \blk00000001/blk00000322  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig00000052 ),
    .O(\blk00000001/sig000002f4 )
  );
  LUT2 #(
    .INIT ( 4'h8 ))
  \blk00000001/blk00000321  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig00000051 ),
    .O(\blk00000001/sig000002f3 )
  );
  LUT2 #(
    .INIT ( 4'h8 ))
  \blk00000001/blk00000320  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig00000059 ),
    .O(\blk00000001/sig000002fb )
  );
  LUT2 #(
    .INIT ( 4'h8 ))
  \blk00000001/blk0000031f  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig00000058 ),
    .O(\blk00000001/sig000002fa )
  );
  LUT2 #(
    .INIT ( 4'h8 ))
  \blk00000001/blk0000031e  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig00000057 ),
    .O(\blk00000001/sig000002f9 )
  );
  LUT2 #(
    .INIT ( 4'h8 ))
  \blk00000001/blk0000031d  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig00000056 ),
    .O(\blk00000001/sig000002f8 )
  );
  LUT2 #(
    .INIT ( 4'h8 ))
  \blk00000001/blk0000031c  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig00000055 ),
    .O(\blk00000001/sig000002f7 )
  );
  LUT2 #(
    .INIT ( 4'h8 ))
  \blk00000001/blk0000031b  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig00000054 ),
    .O(\blk00000001/sig000002f6 )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk0000031a  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig0000034a ),
    .O(\blk00000001/sig00000297 )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk00000319  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig00000349 ),
    .O(\blk00000001/sig00000296 )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk00000318  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig00000348 ),
    .O(\blk00000001/sig00000295 )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk00000317  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig00000347 ),
    .O(\blk00000001/sig00000294 )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk00000316  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig00000346 ),
    .O(\blk00000001/sig00000293 )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk00000315  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig00000345 ),
    .O(\blk00000001/sig00000292 )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk00000314  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig00000344 ),
    .O(\blk00000001/sig00000291 )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk00000313  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig00000343 ),
    .O(\blk00000001/sig00000290 )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk00000312  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig00000342 ),
    .O(\blk00000001/sig0000028f )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk00000311  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig00000353 ),
    .O(\blk00000001/sig000002a0 )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk00000310  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig00000352 ),
    .O(\blk00000001/sig0000029f )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk0000030f  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig00000351 ),
    .O(\blk00000001/sig0000029e )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk0000030e  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig00000350 ),
    .O(\blk00000001/sig0000029d )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk0000030d  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig0000034f ),
    .O(\blk00000001/sig0000029c )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk0000030c  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig0000034e ),
    .O(\blk00000001/sig0000029b )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk0000030b  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig0000034d ),
    .O(\blk00000001/sig0000029a )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk0000030a  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig0000034c ),
    .O(\blk00000001/sig00000299 )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk00000309  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig0000034b ),
    .O(\blk00000001/sig00000298 )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk00000308  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig00000341 ),
    .O(\blk00000001/sig0000028e )
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  \blk00000001/blk00000307  (
    .I0(\blk00000001/sig0000047e ),
    .I1(\blk00000001/sig000003e0 ),
    .I2(\blk00000001/sig00000076 ),
    .O(\blk00000001/sig00000315 )
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  \blk00000001/blk00000306  (
    .I0(\blk00000001/sig0000047e ),
    .I1(\blk00000001/sig000003df ),
    .I2(\blk00000001/sig00000075 ),
    .O(\blk00000001/sig00000314 )
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  \blk00000001/blk00000305  (
    .I0(\blk00000001/sig0000047e ),
    .I1(\blk00000001/sig000003de ),
    .I2(\blk00000001/sig00000074 ),
    .O(\blk00000001/sig00000313 )
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  \blk00000001/blk00000304  (
    .I0(\blk00000001/sig0000047e ),
    .I1(\blk00000001/sig000003dd ),
    .I2(\blk00000001/sig00000073 ),
    .O(\blk00000001/sig00000312 )
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  \blk00000001/blk00000303  (
    .I0(\blk00000001/sig0000047e ),
    .I1(\blk00000001/sig000003dc ),
    .I2(\blk00000001/sig00000072 ),
    .O(\blk00000001/sig00000311 )
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  \blk00000001/blk00000302  (
    .I0(\blk00000001/sig0000047e ),
    .I1(\blk00000001/sig000003db ),
    .I2(\blk00000001/sig00000071 ),
    .O(\blk00000001/sig00000310 )
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  \blk00000001/blk00000301  (
    .I0(\blk00000001/sig0000047e ),
    .I1(\blk00000001/sig000003da ),
    .I2(\blk00000001/sig00000070 ),
    .O(\blk00000001/sig0000030f )
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  \blk00000001/blk00000300  (
    .I0(\blk00000001/sig0000047e ),
    .I1(\blk00000001/sig000003d9 ),
    .I2(\blk00000001/sig0000006f ),
    .O(\blk00000001/sig0000030e )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk000002ff  (
    .I0(\blk00000001/sig0000047e ),
    .I1(\blk00000001/sig000003d8 ),
    .O(\blk00000001/sig0000030d )
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  \blk00000001/blk000002fe  (
    .I0(\blk00000001/sig0000047e ),
    .I1(\blk00000001/sig000003e6 ),
    .I2(\blk00000001/sig0000007c ),
    .O(\blk00000001/sig0000031b )
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  \blk00000001/blk000002fd  (
    .I0(\blk00000001/sig0000047e ),
    .I1(\blk00000001/sig000003e5 ),
    .I2(\blk00000001/sig0000007b ),
    .O(\blk00000001/sig0000031a )
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  \blk00000001/blk000002fc  (
    .I0(\blk00000001/sig0000047e ),
    .I1(\blk00000001/sig000003e4 ),
    .I2(\blk00000001/sig0000007a ),
    .O(\blk00000001/sig00000319 )
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  \blk00000001/blk000002fb  (
    .I0(\blk00000001/sig0000047e ),
    .I1(\blk00000001/sig000003e3 ),
    .I2(\blk00000001/sig00000079 ),
    .O(\blk00000001/sig00000318 )
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  \blk00000001/blk000002fa  (
    .I0(\blk00000001/sig0000047e ),
    .I1(\blk00000001/sig000003e2 ),
    .I2(\blk00000001/sig00000078 ),
    .O(\blk00000001/sig00000317 )
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  \blk00000001/blk000002f9  (
    .I0(\blk00000001/sig0000047e ),
    .I1(\blk00000001/sig000003e1 ),
    .I2(\blk00000001/sig00000077 ),
    .O(\blk00000001/sig00000316 )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk000002f8  (
    .I0(\blk00000001/sig0000047e ),
    .I1(\blk00000001/sig000003d7 ),
    .O(\blk00000001/sig0000030c )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk000002f7  (
    .I0(\blk00000001/sig0000047e ),
    .I1(\blk00000001/sig00000467 ),
    .O(\blk00000001/sig00000305 )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk000002f6  (
    .I0(\blk00000001/sig0000047e ),
    .I1(\blk00000001/sig00000466 ),
    .O(\blk00000001/sig00000304 )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk000002f5  (
    .I0(\blk00000001/sig0000047e ),
    .I1(\blk00000001/sig00000465 ),
    .O(\blk00000001/sig00000303 )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk000002f4  (
    .I0(\blk00000001/sig0000047e ),
    .I1(\blk00000001/sig00000464 ),
    .O(\blk00000001/sig00000302 )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk000002f3  (
    .I0(\blk00000001/sig0000047e ),
    .I1(\blk00000001/sig00000463 ),
    .O(\blk00000001/sig00000301 )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk000002f2  (
    .I0(\blk00000001/sig0000047e ),
    .I1(\blk00000001/sig00000462 ),
    .O(\blk00000001/sig00000300 )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk000002f1  (
    .I0(\blk00000001/sig0000047e ),
    .I1(\blk00000001/sig00000461 ),
    .O(\blk00000001/sig000002ff )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk000002f0  (
    .I0(\blk00000001/sig0000047e ),
    .I1(\blk00000001/sig00000460 ),
    .O(\blk00000001/sig000002fe )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk000002ef  (
    .I0(\blk00000001/sig0000047e ),
    .I1(\blk00000001/sig0000045f ),
    .O(\blk00000001/sig000002fd )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk000002ee  (
    .I0(\blk00000001/sig0000047e ),
    .I1(\blk00000001/sig0000046d ),
    .O(\blk00000001/sig0000030b )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk000002ed  (
    .I0(\blk00000001/sig0000047e ),
    .I1(\blk00000001/sig0000046c ),
    .O(\blk00000001/sig0000030a )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk000002ec  (
    .I0(\blk00000001/sig0000047e ),
    .I1(\blk00000001/sig0000046b ),
    .O(\blk00000001/sig00000309 )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk000002eb  (
    .I0(\blk00000001/sig0000047e ),
    .I1(\blk00000001/sig0000046a ),
    .O(\blk00000001/sig00000308 )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk000002ea  (
    .I0(\blk00000001/sig0000047e ),
    .I1(\blk00000001/sig00000469 ),
    .O(\blk00000001/sig00000307 )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk000002e9  (
    .I0(\blk00000001/sig0000047e ),
    .I1(\blk00000001/sig00000468 ),
    .O(\blk00000001/sig00000306 )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk000002e8  (
    .I0(\blk00000001/sig0000047e ),
    .I1(\blk00000001/sig0000045e ),
    .O(\blk00000001/sig000002fc )
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  \blk00000001/blk000002e7  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig00000500 ),
    .I2(\blk00000001/sig00000093 ),
    .O(\blk00000001/sig00000538 )
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  \blk00000001/blk000002e6  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig000004ff ),
    .I2(\blk00000001/sig00000092 ),
    .O(\blk00000001/sig00000537 )
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  \blk00000001/blk000002e5  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig000004fe ),
    .I2(\blk00000001/sig00000091 ),
    .O(\blk00000001/sig00000536 )
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  \blk00000001/blk000002e4  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig000004fd ),
    .I2(\blk00000001/sig00000090 ),
    .O(\blk00000001/sig00000535 )
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  \blk00000001/blk000002e3  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig000004fc ),
    .I2(\blk00000001/sig0000008f ),
    .O(\blk00000001/sig00000534 )
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  \blk00000001/blk000002e2  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig000004fb ),
    .I2(\blk00000001/sig0000008e ),
    .O(\blk00000001/sig00000533 )
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  \blk00000001/blk000002e1  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig000004fa ),
    .I2(\blk00000001/sig0000008d ),
    .O(\blk00000001/sig00000532 )
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  \blk00000001/blk000002e0  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig000004f9 ),
    .I2(\blk00000001/sig0000008c ),
    .O(\blk00000001/sig00000531 )
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  \blk00000001/blk000002df  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig000004f8 ),
    .I2(\blk00000001/sig0000008b ),
    .O(\blk00000001/sig00000530 )
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  \blk00000001/blk000002de  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig00000509 ),
    .I2(\blk00000001/sig0000009c ),
    .O(\blk00000001/sig00000541 )
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  \blk00000001/blk000002dd  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig00000508 ),
    .I2(\blk00000001/sig0000009b ),
    .O(\blk00000001/sig00000540 )
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  \blk00000001/blk000002dc  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig00000507 ),
    .I2(\blk00000001/sig0000009a ),
    .O(\blk00000001/sig0000053f )
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  \blk00000001/blk000002db  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig00000506 ),
    .I2(\blk00000001/sig00000099 ),
    .O(\blk00000001/sig0000053e )
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  \blk00000001/blk000002da  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig00000505 ),
    .I2(\blk00000001/sig00000098 ),
    .O(\blk00000001/sig0000053d )
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  \blk00000001/blk000002d9  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig00000504 ),
    .I2(\blk00000001/sig00000097 ),
    .O(\blk00000001/sig0000053c )
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  \blk00000001/blk000002d8  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig00000503 ),
    .I2(\blk00000001/sig00000096 ),
    .O(\blk00000001/sig0000053b )
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  \blk00000001/blk000002d7  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig00000502 ),
    .I2(\blk00000001/sig00000095 ),
    .O(\blk00000001/sig0000053a )
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  \blk00000001/blk000002d6  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig00000501 ),
    .I2(\blk00000001/sig00000094 ),
    .O(\blk00000001/sig00000539 )
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  \blk00000001/blk000002d5  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig000004f7 ),
    .I2(\blk00000001/sig0000008a ),
    .O(\blk00000001/sig00000542 )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk000002d4  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig00000456 ),
    .O(\blk00000001/sig000002eb )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk000002d3  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig00000455 ),
    .O(\blk00000001/sig000002ea )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk000002d2  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig00000454 ),
    .O(\blk00000001/sig000002e9 )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk000002d1  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig00000453 ),
    .O(\blk00000001/sig000002e8 )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk000002d0  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig00000452 ),
    .O(\blk00000001/sig000002e7 )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk000002cf  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig00000451 ),
    .O(\blk00000001/sig000002e6 )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk000002ce  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig00000450 ),
    .O(\blk00000001/sig000002e5 )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk000002cd  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig0000044f ),
    .O(\blk00000001/sig000002e4 )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk000002cc  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig0000044e ),
    .O(\blk00000001/sig000002e3 )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk000002cb  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig0000045d ),
    .O(\blk00000001/sig000002f2 )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk000002ca  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig0000045c ),
    .O(\blk00000001/sig000002f1 )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk000002c9  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig0000045b ),
    .O(\blk00000001/sig000002f0 )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk000002c8  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig0000045a ),
    .O(\blk00000001/sig000002ef )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk000002c7  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig00000459 ),
    .O(\blk00000001/sig000002ee )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk000002c6  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig00000458 ),
    .O(\blk00000001/sig000002ed )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk000002c5  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig00000457 ),
    .O(\blk00000001/sig000002ec )
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  \blk00000001/blk000002c4  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig000003cf ),
    .I2(\blk00000001/sig00000062 ),
    .O(\blk00000001/sig000002c8 )
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  \blk00000001/blk000002c3  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig000003ce ),
    .I2(\blk00000001/sig00000061 ),
    .O(\blk00000001/sig000002c7 )
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  \blk00000001/blk000002c2  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig000003cd ),
    .I2(\blk00000001/sig00000060 ),
    .O(\blk00000001/sig000002c6 )
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  \blk00000001/blk000002c1  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig000003cc ),
    .I2(\blk00000001/sig0000005f ),
    .O(\blk00000001/sig000002c5 )
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  \blk00000001/blk000002c0  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig000003cb ),
    .I2(\blk00000001/sig0000005e ),
    .O(\blk00000001/sig000002c4 )
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  \blk00000001/blk000002bf  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig000003ca ),
    .I2(\blk00000001/sig0000005d ),
    .O(\blk00000001/sig000002c3 )
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  \blk00000001/blk000002be  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig000003c9 ),
    .I2(\blk00000001/sig0000005c ),
    .O(\blk00000001/sig000002c2 )
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  \blk00000001/blk000002bd  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig000003c8 ),
    .I2(\blk00000001/sig0000005b ),
    .O(\blk00000001/sig000002c1 )
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  \blk00000001/blk000002bc  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig000003c7 ),
    .I2(\blk00000001/sig0000005a ),
    .O(\blk00000001/sig000002c0 )
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  \blk00000001/blk000002bb  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig000003d6 ),
    .I2(\blk00000001/sig00000069 ),
    .O(\blk00000001/sig000002cf )
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  \blk00000001/blk000002ba  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig000003d5 ),
    .I2(\blk00000001/sig00000068 ),
    .O(\blk00000001/sig000002ce )
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  \blk00000001/blk000002b9  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig000003d4 ),
    .I2(\blk00000001/sig00000067 ),
    .O(\blk00000001/sig000002cd )
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  \blk00000001/blk000002b8  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig000003d3 ),
    .I2(\blk00000001/sig00000066 ),
    .O(\blk00000001/sig000002cc )
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  \blk00000001/blk000002b7  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig000003d2 ),
    .I2(\blk00000001/sig00000065 ),
    .O(\blk00000001/sig000002cb )
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  \blk00000001/blk000002b6  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig000003d1 ),
    .I2(\blk00000001/sig00000064 ),
    .O(\blk00000001/sig000002ca )
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  \blk00000001/blk000002b5  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig000003d0 ),
    .I2(\blk00000001/sig00000063 ),
    .O(\blk00000001/sig000002c9 )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk000002b4  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig0000049b ),
    .O(\blk00000001/sig00000338 )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk000002b3  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig0000049a ),
    .O(\blk00000001/sig00000337 )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk000002b2  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig00000499 ),
    .O(\blk00000001/sig00000336 )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk000002b1  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig00000498 ),
    .O(\blk00000001/sig00000335 )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk000002b0  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig00000497 ),
    .O(\blk00000001/sig00000334 )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk000002af  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig00000496 ),
    .O(\blk00000001/sig00000333 )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk000002ae  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig00000495 ),
    .O(\blk00000001/sig00000332 )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk000002ad  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig00000494 ),
    .O(\blk00000001/sig00000331 )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk000002ac  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig00000493 ),
    .O(\blk00000001/sig00000330 )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk000002ab  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig000004a3 ),
    .O(\blk00000001/sig00000340 )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk000002aa  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig000004a2 ),
    .O(\blk00000001/sig0000033f )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk000002a9  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig000004a1 ),
    .O(\blk00000001/sig0000033e )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk000002a8  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig000004a0 ),
    .O(\blk00000001/sig0000033d )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk000002a7  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig0000049f ),
    .O(\blk00000001/sig0000033c )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk000002a6  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig0000049e ),
    .O(\blk00000001/sig0000033b )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk000002a5  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig0000049d ),
    .O(\blk00000001/sig0000033a )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk000002a4  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig0000049c ),
    .O(\blk00000001/sig00000339 )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk000002a3  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig00000492 ),
    .O(\blk00000001/sig0000032f )
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  \blk00000001/blk000002a2  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig0000004a ),
    .I2(\blk00000001/sig00000094 ),
    .O(\blk00000001/sig00000326 )
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  \blk00000001/blk000002a1  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig00000049 ),
    .I2(\blk00000001/sig00000093 ),
    .O(\blk00000001/sig00000325 )
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  \blk00000001/blk000002a0  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig00000048 ),
    .I2(\blk00000001/sig00000092 ),
    .O(\blk00000001/sig00000324 )
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  \blk00000001/blk0000029f  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig00000047 ),
    .I2(\blk00000001/sig00000091 ),
    .O(\blk00000001/sig00000323 )
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  \blk00000001/blk0000029e  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig00000046 ),
    .I2(\blk00000001/sig00000090 ),
    .O(\blk00000001/sig00000322 )
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  \blk00000001/blk0000029d  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig00000045 ),
    .I2(\blk00000001/sig0000008f ),
    .O(\blk00000001/sig00000321 )
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  \blk00000001/blk0000029c  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig00000044 ),
    .I2(\blk00000001/sig0000008e ),
    .O(\blk00000001/sig00000320 )
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  \blk00000001/blk0000029b  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig00000043 ),
    .I2(\blk00000001/sig0000008d ),
    .O(\blk00000001/sig0000031f )
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  \blk00000001/blk0000029a  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig00000042 ),
    .I2(\blk00000001/sig0000008c ),
    .O(\blk00000001/sig0000031e )
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  \blk00000001/blk00000299  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig00000050 ),
    .I2(\blk00000001/sig0000009c ),
    .O(\blk00000001/sig0000032e )
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  \blk00000001/blk00000298  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig00000050 ),
    .I2(\blk00000001/sig0000009b ),
    .O(\blk00000001/sig0000032d )
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  \blk00000001/blk00000297  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig00000050 ),
    .I2(\blk00000001/sig0000009a ),
    .O(\blk00000001/sig0000032c )
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  \blk00000001/blk00000296  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig0000004f ),
    .I2(\blk00000001/sig00000099 ),
    .O(\blk00000001/sig0000032b )
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  \blk00000001/blk00000295  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig0000004e ),
    .I2(\blk00000001/sig00000098 ),
    .O(\blk00000001/sig0000032a )
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  \blk00000001/blk00000294  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig0000004d ),
    .I2(\blk00000001/sig00000097 ),
    .O(\blk00000001/sig00000329 )
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  \blk00000001/blk00000293  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig0000004c ),
    .I2(\blk00000001/sig00000096 ),
    .O(\blk00000001/sig00000328 )
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  \blk00000001/blk00000292  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig0000004b ),
    .I2(\blk00000001/sig00000095 ),
    .O(\blk00000001/sig00000327 )
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  \blk00000001/blk00000291  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig00000041 ),
    .I2(\blk00000001/sig0000008b ),
    .O(\blk00000001/sig0000031d )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk00000290  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig00000401 ),
    .O(\blk00000001/sig000002d9 )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk0000028f  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig00000400 ),
    .O(\blk00000001/sig000002d8 )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk0000028e  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig000003ff ),
    .O(\blk00000001/sig000002d7 )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk0000028d  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig000003fe ),
    .O(\blk00000001/sig000002d6 )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk0000028c  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig000003fd ),
    .O(\blk00000001/sig000002d5 )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk0000028b  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig000003fc ),
    .O(\blk00000001/sig000002d4 )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk0000028a  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig000003fb ),
    .O(\blk00000001/sig000002d3 )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk00000289  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig000003fa ),
    .O(\blk00000001/sig000002d2 )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk00000288  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig000003f9 ),
    .O(\blk00000001/sig000002d1 )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk00000287  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig0000040a ),
    .O(\blk00000001/sig000002e2 )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk00000286  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig00000409 ),
    .O(\blk00000001/sig000002e1 )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk00000285  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig00000408 ),
    .O(\blk00000001/sig000002e0 )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk00000284  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig00000407 ),
    .O(\blk00000001/sig000002df )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk00000283  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig00000406 ),
    .O(\blk00000001/sig000002de )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk00000282  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig00000405 ),
    .O(\blk00000001/sig000002dd )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk00000281  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig00000404 ),
    .O(\blk00000001/sig000002dc )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk00000280  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig00000403 ),
    .O(\blk00000001/sig000002db )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk0000027f  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig00000402 ),
    .O(\blk00000001/sig000002da )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk0000027e  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig000003f8 ),
    .O(\blk00000001/sig000002d0 )
  );
  LUT3 #(
    .INIT ( 8'h80 ))
  \blk00000001/blk0000027d  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig0000008a ),
    .I2(\blk00000001/sig00000054 ),
    .O(\blk00000001/sig00000288 )
  );
  LUT3 #(
    .INIT ( 8'h80 ))
  \blk00000001/blk0000027c  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig0000008a ),
    .I2(\blk00000001/sig00000053 ),
    .O(\blk00000001/sig00000287 )
  );
  LUT3 #(
    .INIT ( 8'h80 ))
  \blk00000001/blk0000027b  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig0000008a ),
    .I2(\blk00000001/sig00000052 ),
    .O(\blk00000001/sig00000286 )
  );
  LUT3 #(
    .INIT ( 8'h80 ))
  \blk00000001/blk0000027a  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig0000008a ),
    .I2(\blk00000001/sig00000051 ),
    .O(\blk00000001/sig00000285 )
  );
  LUT3 #(
    .INIT ( 8'h80 ))
  \blk00000001/blk00000279  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig0000008a ),
    .I2(\blk00000001/sig00000059 ),
    .O(\blk00000001/sig0000028d )
  );
  LUT3 #(
    .INIT ( 8'h80 ))
  \blk00000001/blk00000278  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig0000008a ),
    .I2(\blk00000001/sig00000058 ),
    .O(\blk00000001/sig0000028c )
  );
  LUT3 #(
    .INIT ( 8'h80 ))
  \blk00000001/blk00000277  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig0000008a ),
    .I2(\blk00000001/sig00000057 ),
    .O(\blk00000001/sig0000028b )
  );
  LUT3 #(
    .INIT ( 8'h80 ))
  \blk00000001/blk00000276  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig0000008a ),
    .I2(\blk00000001/sig00000056 ),
    .O(\blk00000001/sig0000028a )
  );
  LUT3 #(
    .INIT ( 8'h80 ))
  \blk00000001/blk00000275  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig0000008a ),
    .I2(\blk00000001/sig00000055 ),
    .O(\blk00000001/sig00000289 )
  );
  LUT3 #(
    .INIT ( 8'h80 ))
  \blk00000001/blk00000274  (
    .I0(\blk00000001/sig0000003c ),
    .I1(\blk00000001/sig0000008a ),
    .I2(\blk00000001/sig00000069 ),
    .O(\blk00000001/sig00000284 )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk00000273  (
    .I0(\blk00000001/sig00000238 ),
    .I1(\blk00000001/sig00000242 ),
    .O(\blk00000001/sig000001e9 )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk00000272  (
    .I0(\blk00000001/sig00000238 ),
    .I1(\blk00000001/sig00000241 ),
    .O(\blk00000001/sig000001e8 )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk00000271  (
    .I0(\blk00000001/sig00000238 ),
    .I1(\blk00000001/sig00000240 ),
    .O(\blk00000001/sig000001e7 )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk00000270  (
    .I0(\blk00000001/sig00000238 ),
    .I1(\blk00000001/sig0000023f ),
    .O(\blk00000001/sig000001e6 )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk0000026f  (
    .I0(\blk00000001/sig00000238 ),
    .I1(\blk00000001/sig0000023e ),
    .O(\blk00000001/sig000001e5 )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk0000026e  (
    .I0(\blk00000001/sig00000238 ),
    .I1(\blk00000001/sig0000023d ),
    .O(\blk00000001/sig000001e4 )
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  \blk00000001/blk0000026d  (
    .I0(\blk00000001/sig00000238 ),
    .I1(\blk00000001/sig0000020b ),
    .I2(\blk00000001/sig00000253 ),
    .O(\blk00000001/sig0000020a )
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  \blk00000001/blk0000026c  (
    .I0(\blk00000001/sig00000238 ),
    .I1(\blk00000001/sig0000020b ),
    .I2(\blk00000001/sig00000252 ),
    .O(\blk00000001/sig00000209 )
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  \blk00000001/blk0000026b  (
    .I0(\blk00000001/sig00000238 ),
    .I1(\blk00000001/sig0000020b ),
    .I2(\blk00000001/sig00000251 ),
    .O(\blk00000001/sig00000208 )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk0000026a  (
    .I0(\blk00000001/sig00000238 ),
    .I1(\blk00000001/sig0000023c ),
    .O(\blk00000001/sig000001e3 )
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  \blk00000001/blk00000269  (
    .I0(\blk00000001/sig00000238 ),
    .I1(\blk00000001/sig0000020b ),
    .I2(\blk00000001/sig00000250 ),
    .O(\blk00000001/sig00000207 )
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  \blk00000001/blk00000268  (
    .I0(\blk00000001/sig00000238 ),
    .I1(\blk00000001/sig0000020b ),
    .I2(\blk00000001/sig0000024f ),
    .O(\blk00000001/sig00000206 )
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  \blk00000001/blk00000267  (
    .I0(\blk00000001/sig00000238 ),
    .I1(\blk00000001/sig0000020b ),
    .I2(\blk00000001/sig0000024e ),
    .O(\blk00000001/sig00000205 )
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  \blk00000001/blk00000266  (
    .I0(\blk00000001/sig00000238 ),
    .I1(\blk00000001/sig0000020b ),
    .I2(\blk00000001/sig0000024d ),
    .O(\blk00000001/sig00000204 )
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  \blk00000001/blk00000265  (
    .I0(\blk00000001/sig00000238 ),
    .I1(\blk00000001/sig0000020b ),
    .I2(\blk00000001/sig0000024c ),
    .O(\blk00000001/sig00000203 )
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  \blk00000001/blk00000264  (
    .I0(\blk00000001/sig00000238 ),
    .I1(\blk00000001/sig0000020b ),
    .I2(\blk00000001/sig0000024b ),
    .O(\blk00000001/sig00000202 )
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  \blk00000001/blk00000263  (
    .I0(\blk00000001/sig00000238 ),
    .I1(\blk00000001/sig0000020b ),
    .I2(\blk00000001/sig0000024a ),
    .O(\blk00000001/sig00000201 )
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  \blk00000001/blk00000262  (
    .I0(\blk00000001/sig00000238 ),
    .I1(\blk00000001/sig0000020b ),
    .I2(\blk00000001/sig00000249 ),
    .O(\blk00000001/sig00000200 )
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  \blk00000001/blk00000261  (
    .I0(\blk00000001/sig00000238 ),
    .I1(\blk00000001/sig0000020b ),
    .I2(\blk00000001/sig00000248 ),
    .O(\blk00000001/sig000001ff )
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  \blk00000001/blk00000260  (
    .I0(\blk00000001/sig00000238 ),
    .I1(\blk00000001/sig0000020b ),
    .I2(\blk00000001/sig00000247 ),
    .O(\blk00000001/sig000001fe )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk0000025f  (
    .I0(\blk00000001/sig00000238 ),
    .I1(\blk00000001/sig0000023b ),
    .O(\blk00000001/sig000001e2 )
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  \blk00000001/blk0000025e  (
    .I0(\blk00000001/sig00000238 ),
    .I1(\blk00000001/sig0000020b ),
    .I2(\blk00000001/sig00000246 ),
    .O(\blk00000001/sig000001fd )
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  \blk00000001/blk0000025d  (
    .I0(\blk00000001/sig00000238 ),
    .I1(\blk00000001/sig0000020b ),
    .I2(\blk00000001/sig00000245 ),
    .O(\blk00000001/sig000001fc )
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  \blk00000001/blk0000025c  (
    .I0(\blk00000001/sig00000238 ),
    .I1(\blk00000001/sig0000020b ),
    .I2(\blk00000001/sig00000244 ),
    .O(\blk00000001/sig000001fb )
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  \blk00000001/blk0000025b  (
    .I0(\blk00000001/sig00000238 ),
    .I1(\blk00000001/sig00000253 ),
    .I2(\blk00000001/sig00000243 ),
    .O(\blk00000001/sig000001fa )
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  \blk00000001/blk0000025a  (
    .I0(\blk00000001/sig00000238 ),
    .I1(\blk00000001/sig00000252 ),
    .I2(\blk00000001/sig00000242 ),
    .O(\blk00000001/sig000001f9 )
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  \blk00000001/blk00000259  (
    .I0(\blk00000001/sig00000238 ),
    .I1(\blk00000001/sig00000251 ),
    .I2(\blk00000001/sig00000241 ),
    .O(\blk00000001/sig000001f8 )
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  \blk00000001/blk00000258  (
    .I0(\blk00000001/sig00000238 ),
    .I1(\blk00000001/sig00000250 ),
    .I2(\blk00000001/sig00000240 ),
    .O(\blk00000001/sig000001f7 )
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  \blk00000001/blk00000257  (
    .I0(\blk00000001/sig00000238 ),
    .I1(\blk00000001/sig0000024f ),
    .I2(\blk00000001/sig0000023f ),
    .O(\blk00000001/sig000001f6 )
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  \blk00000001/blk00000256  (
    .I0(\blk00000001/sig00000238 ),
    .I1(\blk00000001/sig0000024e ),
    .I2(\blk00000001/sig0000023e ),
    .O(\blk00000001/sig000001f5 )
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  \blk00000001/blk00000255  (
    .I0(\blk00000001/sig00000238 ),
    .I1(\blk00000001/sig0000024d ),
    .I2(\blk00000001/sig0000023d ),
    .O(\blk00000001/sig000001f4 )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk00000254  (
    .I0(\blk00000001/sig00000238 ),
    .I1(\blk00000001/sig0000023a ),
    .O(\blk00000001/sig000001e1 )
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  \blk00000001/blk00000253  (
    .I0(\blk00000001/sig00000238 ),
    .I1(\blk00000001/sig0000024c ),
    .I2(\blk00000001/sig0000023c ),
    .O(\blk00000001/sig000001f3 )
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  \blk00000001/blk00000252  (
    .I0(\blk00000001/sig00000238 ),
    .I1(\blk00000001/sig0000024b ),
    .I2(\blk00000001/sig0000023b ),
    .O(\blk00000001/sig000001f2 )
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  \blk00000001/blk00000251  (
    .I0(\blk00000001/sig00000238 ),
    .I1(\blk00000001/sig0000024a ),
    .I2(\blk00000001/sig0000023a ),
    .O(\blk00000001/sig000001f1 )
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  \blk00000001/blk00000250  (
    .I0(\blk00000001/sig00000238 ),
    .I1(\blk00000001/sig00000249 ),
    .I2(\blk00000001/sig00000239 ),
    .O(\blk00000001/sig000001f0 )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk0000024f  (
    .I0(\blk00000001/sig00000238 ),
    .I1(\blk00000001/sig00000248 ),
    .O(\blk00000001/sig000001ef )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk0000024e  (
    .I0(\blk00000001/sig00000238 ),
    .I1(\blk00000001/sig00000247 ),
    .O(\blk00000001/sig000001ee )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk0000024d  (
    .I0(\blk00000001/sig00000238 ),
    .I1(\blk00000001/sig00000246 ),
    .O(\blk00000001/sig000001ed )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk0000024c  (
    .I0(\blk00000001/sig00000238 ),
    .I1(\blk00000001/sig00000245 ),
    .O(\blk00000001/sig000001ec )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk0000024b  (
    .I0(\blk00000001/sig00000238 ),
    .I1(\blk00000001/sig00000244 ),
    .O(\blk00000001/sig000001eb )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk0000024a  (
    .I0(\blk00000001/sig00000238 ),
    .I1(\blk00000001/sig00000243 ),
    .O(\blk00000001/sig000001ea )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk00000249  (
    .I0(\blk00000001/sig00000238 ),
    .I1(\blk00000001/sig00000239 ),
    .O(\blk00000001/sig000001e0 )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk00000248  (
    .I0(\blk00000001/sig000000fc ),
    .I1(\blk00000001/sig000000c6 ),
    .O(\blk00000001/sig00000191 )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk00000247  (
    .I0(\blk00000001/sig000000fc ),
    .I1(\blk00000001/sig000000c5 ),
    .O(\blk00000001/sig00000190 )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk00000246  (
    .I0(\blk00000001/sig000000fc ),
    .I1(\blk00000001/sig000000c4 ),
    .O(\blk00000001/sig0000018f )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk00000245  (
    .I0(\blk00000001/sig000000fc ),
    .I1(\blk00000001/sig000000c3 ),
    .O(\blk00000001/sig0000018e )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk00000244  (
    .I0(\blk00000001/sig000000fc ),
    .I1(\blk00000001/sig000000c1 ),
    .O(\blk00000001/sig0000018c )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk00000243  (
    .I0(\blk00000001/sig000000fc ),
    .I1(\blk00000001/sig000000c0 ),
    .O(\blk00000001/sig0000018b )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk00000242  (
    .I0(\blk00000001/sig000000fc ),
    .I1(\blk00000001/sig000000c2 ),
    .O(\blk00000001/sig0000018d )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk00000241  (
    .I0(\blk00000001/sig000000fc ),
    .I1(\blk00000001/sig000000bf ),
    .O(\blk00000001/sig0000018a )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk00000240  (
    .I0(\blk00000001/sig000000fc ),
    .I1(\blk00000001/sig000000be ),
    .O(\blk00000001/sig00000189 )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk0000023f  (
    .I0(\blk00000001/sig000000fc ),
    .I1(\blk00000001/sig000000bb ),
    .O(\blk00000001/sig00000186 )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk0000023e  (
    .I0(\blk00000001/sig000000fc ),
    .I1(\blk00000001/sig000000bd ),
    .O(\blk00000001/sig00000188 )
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk00000001/blk0000023d  (
    .I0(\blk00000001/sig000000fc ),
    .I1(\blk00000001/sig000000bc ),
    .O(\blk00000001/sig00000187 )
  );
  LUT2 #(
    .INIT ( 4'h7 ))
  \blk00000001/blk0000023c  (
    .I0(\blk00000001/sig0000016b ),
    .I1(\blk00000001/sig00000161 ),
    .O(\blk00000001/sig0000016a )
  );
  LUT3 #(
    .INIT ( 8'h10 ))
  \blk00000001/blk0000023b  (
    .I0(\blk00000001/sig000000cd ),
    .I1(\blk00000001/sig000000cc ),
    .I2(\blk00000001/sig0000015a ),
    .O(\blk00000001/sig00000140 )
  );
  LUT4 #(
    .INIT ( 16'h5410 ))
  \blk00000001/blk0000023a  (
    .I0(\blk00000001/sig000000cd ),
    .I1(\blk00000001/sig000000cc ),
    .I2(\blk00000001/sig00000159 ),
    .I3(\blk00000001/sig0000015a ),
    .O(\blk00000001/sig0000013f )
  );
  LUT6 #(
    .INIT ( 64'hFD75EC64B931A820 ))
  \blk00000001/blk00000239  (
    .I0(\blk00000001/sig000000cc ),
    .I1(\blk00000001/sig000000cd ),
    .I2(\blk00000001/sig00000150 ),
    .I3(\blk00000001/sig00000152 ),
    .I4(\blk00000001/sig0000014f ),
    .I5(\blk00000001/sig00000151 ),
    .O(\blk00000001/sig00000135 )
  );
  LUT6 #(
    .INIT ( 64'hFD75EC64B931A820 ))
  \blk00000001/blk00000238  (
    .I0(\blk00000001/sig000000cc ),
    .I1(\blk00000001/sig000000cd ),
    .I2(\blk00000001/sig0000014f ),
    .I3(\blk00000001/sig00000151 ),
    .I4(\blk00000001/sig0000014e ),
    .I5(\blk00000001/sig00000150 ),
    .O(\blk00000001/sig00000134 )
  );
  LUT6 #(
    .INIT ( 64'hFD75EC64B931A820 ))
  \blk00000001/blk00000237  (
    .I0(\blk00000001/sig000000cc ),
    .I1(\blk00000001/sig000000cd ),
    .I2(\blk00000001/sig00000151 ),
    .I3(\blk00000001/sig00000153 ),
    .I4(\blk00000001/sig00000150 ),
    .I5(\blk00000001/sig00000152 ),
    .O(\blk00000001/sig00000136 )
  );
  LUT6 #(
    .INIT ( 64'hFD75EC64B931A820 ))
  \blk00000001/blk00000236  (
    .I0(\blk00000001/sig000000cc ),
    .I1(\blk00000001/sig000000cd ),
    .I2(\blk00000001/sig00000152 ),
    .I3(\blk00000001/sig00000154 ),
    .I4(\blk00000001/sig00000151 ),
    .I5(\blk00000001/sig00000153 ),
    .O(\blk00000001/sig00000137 )
  );
  LUT6 #(
    .INIT ( 64'hFD75EC64B931A820 ))
  \blk00000001/blk00000235  (
    .I0(\blk00000001/sig000000cc ),
    .I1(\blk00000001/sig000000cd ),
    .I2(\blk00000001/sig00000153 ),
    .I3(\blk00000001/sig00000155 ),
    .I4(\blk00000001/sig00000152 ),
    .I5(\blk00000001/sig00000154 ),
    .O(\blk00000001/sig00000138 )
  );
  LUT6 #(
    .INIT ( 64'hFD75EC64B931A820 ))
  \blk00000001/blk00000234  (
    .I0(\blk00000001/sig000000cc ),
    .I1(\blk00000001/sig000000cd ),
    .I2(\blk00000001/sig00000154 ),
    .I3(\blk00000001/sig00000156 ),
    .I4(\blk00000001/sig00000153 ),
    .I5(\blk00000001/sig00000155 ),
    .O(\blk00000001/sig00000139 )
  );
  LUT6 #(
    .INIT ( 64'hFD75EC64B931A820 ))
  \blk00000001/blk00000233  (
    .I0(\blk00000001/sig000000cc ),
    .I1(\blk00000001/sig000000cd ),
    .I2(\blk00000001/sig00000155 ),
    .I3(\blk00000001/sig00000157 ),
    .I4(\blk00000001/sig00000154 ),
    .I5(\blk00000001/sig00000156 ),
    .O(\blk00000001/sig0000013a )
  );
  LUT6 #(
    .INIT ( 64'hFD75EC64B931A820 ))
  \blk00000001/blk00000232  (
    .I0(\blk00000001/sig000000cc ),
    .I1(\blk00000001/sig000000cd ),
    .I2(\blk00000001/sig00000158 ),
    .I3(\blk00000001/sig0000015a ),
    .I4(\blk00000001/sig00000157 ),
    .I5(\blk00000001/sig00000159 ),
    .O(\blk00000001/sig0000013d )
  );
  LUT6 #(
    .INIT ( 64'hFD75EC64B931A820 ))
  \blk00000001/blk00000231  (
    .I0(\blk00000001/sig000000cc ),
    .I1(\blk00000001/sig000000cd ),
    .I2(\blk00000001/sig00000156 ),
    .I3(\blk00000001/sig00000158 ),
    .I4(\blk00000001/sig00000155 ),
    .I5(\blk00000001/sig00000157 ),
    .O(\blk00000001/sig0000013b )
  );
  LUT5 #(
    .INIT ( 32'h73625140 ))
  \blk00000001/blk00000230  (
    .I0(\blk00000001/sig000000cd ),
    .I1(\blk00000001/sig000000cc ),
    .I2(\blk00000001/sig00000159 ),
    .I3(\blk00000001/sig00000158 ),
    .I4(\blk00000001/sig0000015a ),
    .O(\blk00000001/sig0000013e )
  );
  LUT6 #(
    .INIT ( 64'hFD75EC64B931A820 ))
  \blk00000001/blk0000022f  (
    .I0(\blk00000001/sig000000cc ),
    .I1(\blk00000001/sig000000cd ),
    .I2(\blk00000001/sig00000157 ),
    .I3(\blk00000001/sig00000159 ),
    .I4(\blk00000001/sig00000156 ),
    .I5(\blk00000001/sig00000158 ),
    .O(\blk00000001/sig0000013c )
  );
  LUT6 #(
    .INIT ( 64'hFD75EC64B931A820 ))
  \blk00000001/blk0000022e  (
    .I0(\blk00000001/sig000000ce ),
    .I1(\blk00000001/sig000000cf ),
    .I2(\blk00000001/sig000000d8 ),
    .I3(\blk00000001/sig000000d0 ),
    .I4(\blk00000001/sig000000dc ),
    .I5(\blk00000001/sig000000d4 ),
    .O(\blk00000001/sig00000141 )
  );
  LUT2 #(
    .INIT ( 4'h8 ))
  \blk00000001/blk0000022d  (
    .I0(\blk00000001/sig00000127 ),
    .I1(\blk00000001/sig000000cf ),
    .O(\blk00000001/sig00000133 )
  );
  LUT2 #(
    .INIT ( 4'h8 ))
  \blk00000001/blk0000022c  (
    .I0(\blk00000001/sig00000126 ),
    .I1(\blk00000001/sig00000125 ),
    .O(\blk00000001/sig00000132 )
  );
  LUT5 #(
    .INIT ( 32'h01010100 ))
  \blk00000001/blk0000022b  (
    .I0(\blk00000001/sig00000126 ),
    .I1(\blk00000001/sig000000d4 ),
    .I2(\blk00000001/sig000000d5 ),
    .I3(\blk00000001/sig000000d2 ),
    .I4(\blk00000001/sig000000d3 ),
    .O(\blk00000001/sig0000012e )
  );
  LUT2 #(
    .INIT ( 4'h1 ))
  \blk00000001/blk0000022a  (
    .I0(\blk00000001/sig000000de ),
    .I1(\blk00000001/sig000000dd ),
    .O(\blk00000001/sig00000124 )
  );
  LUT4 #(
    .INIT ( 16'h0001 ))
  \blk00000001/blk00000229  (
    .I0(\blk00000001/sig000000e0 ),
    .I1(\blk00000001/sig000000df ),
    .I2(\blk00000001/sig000000e2 ),
    .I3(\blk00000001/sig000000e1 ),
    .O(\blk00000001/sig00000123 )
  );
  LUT4 #(
    .INIT ( 16'h0001 ))
  \blk00000001/blk00000228  (
    .I0(\blk00000001/sig000000e6 ),
    .I1(\blk00000001/sig000000e5 ),
    .I2(\blk00000001/sig000000e4 ),
    .I3(\blk00000001/sig000000e3 ),
    .O(\blk00000001/sig00000122 )
  );
  LUT3 #(
    .INIT ( 8'h01 ))
  \blk00000001/blk00000227  (
    .I0(\blk00000001/sig000000e9 ),
    .I1(\blk00000001/sig000000e8 ),
    .I2(\blk00000001/sig000000e7 ),
    .O(\blk00000001/sig00000121 )
  );
  LUT2 #(
    .INIT ( 4'h8 ))
  \blk00000001/blk00000226  (
    .I0(\blk00000001/sig000000cf ),
    .I1(\blk00000001/sig00000125 ),
    .O(\blk00000001/sig00000120 )
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  \blk00000001/blk00000225  (
    .I0(\blk00000001/sig000000cf ),
    .I1(\blk00000001/sig00000127 ),
    .I2(\blk00000001/sig00000126 ),
    .O(\blk00000001/sig000000ce )
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  \blk00000001/blk00000224  (
    .I0(\blk00000001/sig000000c9 ),
    .I1(\blk00000001/sig000000c8 ),
    .O(\blk00000001/sig00000102 )
  );
  LUT3 #(
    .INIT ( 8'h56 ))
  \blk00000001/blk00000223  (
    .I0(\blk00000001/sig000000ca ),
    .I1(\blk00000001/sig000000c9 ),
    .I2(\blk00000001/sig000000c8 ),
    .O(\blk00000001/sig00000103 )
  );
  LUT6 #(
    .INIT ( 64'h5050505014505050 ))
  \blk00000001/blk00000222  (
    .I0(\blk00000001/sig000000fc ),
    .I1(\blk00000001/sig000000ff ),
    .I2(\blk00000001/sig00000100 ),
    .I3(\blk00000001/sig000000fe ),
    .I4(\blk00000001/sig000000fd ),
    .I5(\blk00000001/sig00000167 ),
    .O(\blk00000001/sig000000fa )
  );
  LUT5 #(
    .INIT ( 32'h44441444 ))
  \blk00000001/blk00000221  (
    .I0(\blk00000001/sig000000fc ),
    .I1(\blk00000001/sig000000ff ),
    .I2(\blk00000001/sig000000fe ),
    .I3(\blk00000001/sig000000fd ),
    .I4(\blk00000001/sig00000167 ),
    .O(\blk00000001/sig000000f9 )
  );
  LUT4 #(
    .INIT ( 16'h4414 ))
  \blk00000001/blk00000220  (
    .I0(\blk00000001/sig000000fc ),
    .I1(\blk00000001/sig000000fe ),
    .I2(\blk00000001/sig000000fd ),
    .I3(\blk00000001/sig00000167 ),
    .O(\blk00000001/sig000000f8 )
  );
  LUT3 #(
    .INIT ( 8'h41 ))
  \blk00000001/blk0000021f  (
    .I0(\blk00000001/sig000000fc ),
    .I1(\blk00000001/sig000000fd ),
    .I2(\blk00000001/sig00000167 ),
    .O(\blk00000001/sig000000f7 )
  );
  LUT4 #(
    .INIT ( 16'hFFFE ))
  \blk00000001/blk0000021e  (
    .I0(\blk00000001/sig000000cb ),
    .I1(\blk00000001/sig000000c8 ),
    .I2(\blk00000001/sig000000c9 ),
    .I3(\blk00000001/sig000000ca ),
    .O(\blk00000001/sig00000105 )
  );
  LUT4 #(
    .INIT ( 16'h5556 ))
  \blk00000001/blk0000021d  (
    .I0(\blk00000001/sig000000cb ),
    .I1(\blk00000001/sig000000c8 ),
    .I2(\blk00000001/sig000000c9 ),
    .I3(\blk00000001/sig000000ca ),
    .O(\blk00000001/sig00000104 )
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  \blk00000001/blk0000021c  (
    .I0(s_axis_divisor_tdata[9]),
    .I1(s_axis_divisor_tdata[12]),
    .O(\blk00000001/sig000000f3 )
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  \blk00000001/blk0000021b  (
    .I0(s_axis_divisor_tdata[8]),
    .I1(s_axis_divisor_tdata[12]),
    .O(\blk00000001/sig000000f2 )
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  \blk00000001/blk0000021a  (
    .I0(s_axis_divisor_tdata[7]),
    .I1(s_axis_divisor_tdata[12]),
    .O(\blk00000001/sig000000f1 )
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  \blk00000001/blk00000219  (
    .I0(s_axis_divisor_tdata[6]),
    .I1(s_axis_divisor_tdata[12]),
    .O(\blk00000001/sig000000f0 )
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  \blk00000001/blk00000218  (
    .I0(s_axis_divisor_tdata[5]),
    .I1(s_axis_divisor_tdata[12]),
    .O(\blk00000001/sig000000ef )
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  \blk00000001/blk00000217  (
    .I0(s_axis_divisor_tdata[4]),
    .I1(s_axis_divisor_tdata[12]),
    .O(\blk00000001/sig000000ee )
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  \blk00000001/blk00000216  (
    .I0(s_axis_divisor_tdata[3]),
    .I1(s_axis_divisor_tdata[12]),
    .O(\blk00000001/sig000000ed )
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  \blk00000001/blk00000215  (
    .I0(s_axis_divisor_tdata[2]),
    .I1(s_axis_divisor_tdata[12]),
    .O(\blk00000001/sig000000ec )
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  \blk00000001/blk00000214  (
    .I0(s_axis_divisor_tdata[1]),
    .I1(s_axis_divisor_tdata[12]),
    .O(\blk00000001/sig000000eb )
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  \blk00000001/blk00000213  (
    .I0(s_axis_divisor_tdata[11]),
    .I1(s_axis_divisor_tdata[12]),
    .O(\blk00000001/sig000000f5 )
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  \blk00000001/blk00000212  (
    .I0(s_axis_divisor_tdata[10]),
    .I1(s_axis_divisor_tdata[12]),
    .O(\blk00000001/sig000000f4 )
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  \blk00000001/blk00000211  (
    .I0(s_axis_divisor_tdata[0]),
    .I1(s_axis_divisor_tdata[12]),
    .O(\blk00000001/sig000000ea )
  );
  LUT3 #(
    .INIT ( 8'h40 ))
  \blk00000001/blk00000210  (
    .I0(\blk00000001/sig0000003d ),
    .I1(s_axis_dividend_tvalid),
    .I2(s_axis_divisor_tvalid),
    .O(\blk00000001/sig00000039 )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000020f  (
    .C(aclk),
    .D(\blk00000001/sig00000545 ),
    .Q(\blk00000001/sig0000055c )
  );
  DSP48A1 #(
    .A0REG ( 0 ),
    .A1REG ( 1 ),
    .B0REG ( 0 ),
    .B1REG ( 1 ),
    .CARRYINREG ( 0 ),
    .CARRYINSEL ( "OPMODE5" ),
    .CREG ( 1 ),
    .DREG ( 1 ),
    .MREG ( 0 ),
    .OPMODEREG ( 1 ),
    .PREG ( 1 ),
    .RSTTYPE ( "SYNC" ),
    .CARRYOUTREG ( 0 ))
  \blk00000001/blk0000020e  (
    .CECARRYIN(\blk00000001/sig0000051d ),
    .RSTC(\blk00000001/sig0000051d ),
    .RSTCARRYIN(\blk00000001/sig0000051d ),
    .CED(\blk00000001/sig0000003a ),
    .RSTD(\blk00000001/sig0000051d ),
    .CEOPMODE(\blk00000001/sig0000003a ),
    .CEC(\blk00000001/sig0000003a ),
    .CARRYOUTF(\NLW_blk00000001/blk0000020e_CARRYOUTF_UNCONNECTED ),
    .RSTOPMODE(\blk00000001/sig0000051d ),
    .RSTM(\blk00000001/sig0000051d ),
    .CLK(aclk),
    .RSTB(\blk00000001/sig0000051d ),
    .CEM(\blk00000001/sig0000051d ),
    .CEB(\blk00000001/sig0000003a ),
    .CARRYIN(\blk00000001/sig0000051d ),
    .CEP(\blk00000001/sig0000003a ),
    .CEA(\blk00000001/sig0000003a ),
    .CARRYOUT(\NLW_blk00000001/blk0000020e_CARRYOUT_UNCONNECTED ),
    .RSTA(\blk00000001/sig0000051d ),
    .RSTP(\blk00000001/sig0000051d ),
    .B({\blk00000001/sig00000050 , \blk00000001/sig00000050 , \blk00000001/sig00000050 , \blk00000001/sig0000004f , \blk00000001/sig0000004e ,
\blk00000001/sig0000004d , \blk00000001/sig0000004c , \blk00000001/sig0000004b , \blk00000001/sig0000004a , \blk00000001/sig00000049 ,
\blk00000001/sig00000048 , \blk00000001/sig00000047 , \blk00000001/sig00000046 , \blk00000001/sig00000045 , \blk00000001/sig00000044 ,
\blk00000001/sig00000043 , \blk00000001/sig00000042 , \blk00000001/sig00000041 }),
    .BCOUT({\NLW_blk00000001/blk0000020e_BCOUT<17>_UNCONNECTED , \NLW_blk00000001/blk0000020e_BCOUT<16>_UNCONNECTED ,
\NLW_blk00000001/blk0000020e_BCOUT<15>_UNCONNECTED , \NLW_blk00000001/blk0000020e_BCOUT<14>_UNCONNECTED ,
\NLW_blk00000001/blk0000020e_BCOUT<13>_UNCONNECTED , \NLW_blk00000001/blk0000020e_BCOUT<12>_UNCONNECTED ,
\NLW_blk00000001/blk0000020e_BCOUT<11>_UNCONNECTED , \NLW_blk00000001/blk0000020e_BCOUT<10>_UNCONNECTED ,
\NLW_blk00000001/blk0000020e_BCOUT<9>_UNCONNECTED , \NLW_blk00000001/blk0000020e_BCOUT<8>_UNCONNECTED ,
\NLW_blk00000001/blk0000020e_BCOUT<7>_UNCONNECTED , \NLW_blk00000001/blk0000020e_BCOUT<6>_UNCONNECTED ,
\NLW_blk00000001/blk0000020e_BCOUT<5>_UNCONNECTED , \NLW_blk00000001/blk0000020e_BCOUT<4>_UNCONNECTED ,
\NLW_blk00000001/blk0000020e_BCOUT<3>_UNCONNECTED , \NLW_blk00000001/blk0000020e_BCOUT<2>_UNCONNECTED ,
\NLW_blk00000001/blk0000020e_BCOUT<1>_UNCONNECTED , \NLW_blk00000001/blk0000020e_BCOUT<0>_UNCONNECTED }),
    .PCIN({\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d }),
    .C({\blk00000001/sig00000556 , \blk00000001/sig00000556 , \blk00000001/sig00000556 , \blk00000001/sig00000556 , \blk00000001/sig00000556 ,
\blk00000001/sig00000556 , \blk00000001/sig00000556 , \blk00000001/sig00000556 , \blk00000001/sig00000556 , \blk00000001/sig00000556 ,
\blk00000001/sig00000556 , \blk00000001/sig00000556 , \blk00000001/sig00000556 , \blk00000001/sig00000556 , \blk00000001/sig00000556 ,
\blk00000001/sig00000556 , \blk00000001/sig00000556 , \blk00000001/sig00000556 , \blk00000001/sig00000556 , \blk00000001/sig00000555 ,
\blk00000001/sig00000554 , \blk00000001/sig00000553 , \blk00000001/sig00000552 , \blk00000001/sig00000551 , \blk00000001/sig00000550 ,
\blk00000001/sig0000054f , \blk00000001/sig0000054e , \blk00000001/sig0000054d , \blk00000001/sig0000054c , \blk00000001/sig0000054b ,
\blk00000001/sig0000054a , \blk00000001/sig00000549 , \blk00000001/sig00000548 , \blk00000001/sig00000547 , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000003f ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d }),
    .P({\NLW_blk00000001/blk0000020e_P<47>_UNCONNECTED , \NLW_blk00000001/blk0000020e_P<46>_UNCONNECTED ,
\NLW_blk00000001/blk0000020e_P<45>_UNCONNECTED , \NLW_blk00000001/blk0000020e_P<44>_UNCONNECTED , \NLW_blk00000001/blk0000020e_P<43>_UNCONNECTED ,
\NLW_blk00000001/blk0000020e_P<42>_UNCONNECTED , \NLW_blk00000001/blk0000020e_P<41>_UNCONNECTED , \NLW_blk00000001/blk0000020e_P<40>_UNCONNECTED ,
\NLW_blk00000001/blk0000020e_P<39>_UNCONNECTED , \NLW_blk00000001/blk0000020e_P<38>_UNCONNECTED , \NLW_blk00000001/blk0000020e_P<37>_UNCONNECTED ,
\NLW_blk00000001/blk0000020e_P<36>_UNCONNECTED , \NLW_blk00000001/blk0000020e_P<35>_UNCONNECTED , \NLW_blk00000001/blk0000020e_P<34>_UNCONNECTED ,
\NLW_blk00000001/blk0000020e_P<33>_UNCONNECTED , \NLW_blk00000001/blk0000020e_P<32>_UNCONNECTED , \NLW_blk00000001/blk0000020e_P<31>_UNCONNECTED ,
\NLW_blk00000001/blk0000020e_P<30>_UNCONNECTED , \NLW_blk00000001/blk0000020e_P<29>_UNCONNECTED , NlwRenamedSignal_m_axis_dout_tdata[24],
m_axis_dout_tdata[23], m_axis_dout_tdata[22], m_axis_dout_tdata[21], m_axis_dout_tdata[20], m_axis_dout_tdata[19], m_axis_dout_tdata[18],
m_axis_dout_tdata[17], m_axis_dout_tdata[16], m_axis_dout_tdata[15], m_axis_dout_tdata[14], m_axis_dout_tdata[13], m_axis_dout_tdata[12],
NlwRenamedSig_OI_m_axis_dout_tdata[11], NlwRenamedSig_OI_m_axis_dout_tdata[10], NlwRenamedSig_OI_m_axis_dout_tdata[9],
NlwRenamedSig_OI_m_axis_dout_tdata[8], NlwRenamedSig_OI_m_axis_dout_tdata[7], NlwRenamedSig_OI_m_axis_dout_tdata[6],
NlwRenamedSig_OI_m_axis_dout_tdata[5], NlwRenamedSig_OI_m_axis_dout_tdata[4], NlwRenamedSig_OI_m_axis_dout_tdata[3],
NlwRenamedSig_OI_m_axis_dout_tdata[2], NlwRenamedSig_OI_m_axis_dout_tdata[1], NlwRenamedSig_OI_m_axis_dout_tdata[0], \blk00000001/sig0000055a ,
\blk00000001/sig00000559 , \blk00000001/sig00000558 , \blk00000001/sig00000557 }),
    .OPMODE({\blk00000001/sig00000545 , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000055b ,
\blk00000001/sig0000055b , \blk00000001/sig0000003a , \blk00000001/sig0000003a }),
    .D({\blk00000001/sig00000050 , \blk00000001/sig00000050 , \blk00000001/sig00000050 , \blk00000001/sig00000050 , \blk00000001/sig00000050 ,
\blk00000001/sig00000050 , \blk00000001/sig00000050 , \blk00000001/sig00000050 , \blk00000001/sig00000050 , \blk00000001/sig00000050 ,
\blk00000001/sig00000050 , \blk00000001/sig00000050 , \blk00000001/sig00000050 , \blk00000001/sig00000050 , \blk00000001/sig00000050 ,
\blk00000001/sig00000050 , \blk00000001/sig00000050 , \blk00000001/sig00000050 }),
    .PCOUT({\NLW_blk00000001/blk0000020e_PCOUT<47>_UNCONNECTED , \NLW_blk00000001/blk0000020e_PCOUT<46>_UNCONNECTED ,
\NLW_blk00000001/blk0000020e_PCOUT<45>_UNCONNECTED , \NLW_blk00000001/blk0000020e_PCOUT<44>_UNCONNECTED ,
\NLW_blk00000001/blk0000020e_PCOUT<43>_UNCONNECTED , \NLW_blk00000001/blk0000020e_PCOUT<42>_UNCONNECTED ,
\NLW_blk00000001/blk0000020e_PCOUT<41>_UNCONNECTED , \NLW_blk00000001/blk0000020e_PCOUT<40>_UNCONNECTED ,
\NLW_blk00000001/blk0000020e_PCOUT<39>_UNCONNECTED , \NLW_blk00000001/blk0000020e_PCOUT<38>_UNCONNECTED ,
\NLW_blk00000001/blk0000020e_PCOUT<37>_UNCONNECTED , \NLW_blk00000001/blk0000020e_PCOUT<36>_UNCONNECTED ,
\NLW_blk00000001/blk0000020e_PCOUT<35>_UNCONNECTED , \NLW_blk00000001/blk0000020e_PCOUT<34>_UNCONNECTED ,
\NLW_blk00000001/blk0000020e_PCOUT<33>_UNCONNECTED , \NLW_blk00000001/blk0000020e_PCOUT<32>_UNCONNECTED ,
\NLW_blk00000001/blk0000020e_PCOUT<31>_UNCONNECTED , \NLW_blk00000001/blk0000020e_PCOUT<30>_UNCONNECTED ,
\NLW_blk00000001/blk0000020e_PCOUT<29>_UNCONNECTED , \NLW_blk00000001/blk0000020e_PCOUT<28>_UNCONNECTED ,
\NLW_blk00000001/blk0000020e_PCOUT<27>_UNCONNECTED , \NLW_blk00000001/blk0000020e_PCOUT<26>_UNCONNECTED ,
\NLW_blk00000001/blk0000020e_PCOUT<25>_UNCONNECTED , \NLW_blk00000001/blk0000020e_PCOUT<24>_UNCONNECTED ,
\NLW_blk00000001/blk0000020e_PCOUT<23>_UNCONNECTED , \NLW_blk00000001/blk0000020e_PCOUT<22>_UNCONNECTED ,
\NLW_blk00000001/blk0000020e_PCOUT<21>_UNCONNECTED , \NLW_blk00000001/blk0000020e_PCOUT<20>_UNCONNECTED ,
\NLW_blk00000001/blk0000020e_PCOUT<19>_UNCONNECTED , \NLW_blk00000001/blk0000020e_PCOUT<18>_UNCONNECTED ,
\NLW_blk00000001/blk0000020e_PCOUT<17>_UNCONNECTED , \NLW_blk00000001/blk0000020e_PCOUT<16>_UNCONNECTED ,
\NLW_blk00000001/blk0000020e_PCOUT<15>_UNCONNECTED , \NLW_blk00000001/blk0000020e_PCOUT<14>_UNCONNECTED ,
\NLW_blk00000001/blk0000020e_PCOUT<13>_UNCONNECTED , \NLW_blk00000001/blk0000020e_PCOUT<12>_UNCONNECTED ,
\NLW_blk00000001/blk0000020e_PCOUT<11>_UNCONNECTED , \NLW_blk00000001/blk0000020e_PCOUT<10>_UNCONNECTED ,
\NLW_blk00000001/blk0000020e_PCOUT<9>_UNCONNECTED , \NLW_blk00000001/blk0000020e_PCOUT<8>_UNCONNECTED ,
\NLW_blk00000001/blk0000020e_PCOUT<7>_UNCONNECTED , \NLW_blk00000001/blk0000020e_PCOUT<6>_UNCONNECTED ,
\NLW_blk00000001/blk0000020e_PCOUT<5>_UNCONNECTED , \NLW_blk00000001/blk0000020e_PCOUT<4>_UNCONNECTED ,
\NLW_blk00000001/blk0000020e_PCOUT<3>_UNCONNECTED , \NLW_blk00000001/blk0000020e_PCOUT<2>_UNCONNECTED ,
\NLW_blk00000001/blk0000020e_PCOUT<1>_UNCONNECTED , \NLW_blk00000001/blk0000020e_PCOUT<0>_UNCONNECTED }),
    .A({\blk00000001/sig00000050 , \blk00000001/sig00000050 , \blk00000001/sig00000050 , \blk00000001/sig00000050 , \blk00000001/sig00000050 ,
\blk00000001/sig00000050 , \blk00000001/sig00000050 , \blk00000001/sig00000050 , \blk00000001/sig00000050 , \blk00000001/sig00000050 ,
\blk00000001/sig00000050 , \blk00000001/sig00000050 , \blk00000001/sig00000050 , \blk00000001/sig00000050 , \blk00000001/sig00000050 ,
\blk00000001/sig00000050 , \blk00000001/sig00000050 , \blk00000001/sig00000050 }),
    .M({\NLW_blk00000001/blk0000020e_M<35>_UNCONNECTED , \NLW_blk00000001/blk0000020e_M<34>_UNCONNECTED ,
\NLW_blk00000001/blk0000020e_M<33>_UNCONNECTED , \NLW_blk00000001/blk0000020e_M<32>_UNCONNECTED , \NLW_blk00000001/blk0000020e_M<31>_UNCONNECTED ,
\NLW_blk00000001/blk0000020e_M<30>_UNCONNECTED , \NLW_blk00000001/blk0000020e_M<29>_UNCONNECTED , \NLW_blk00000001/blk0000020e_M<28>_UNCONNECTED ,
\NLW_blk00000001/blk0000020e_M<27>_UNCONNECTED , \NLW_blk00000001/blk0000020e_M<26>_UNCONNECTED , \NLW_blk00000001/blk0000020e_M<25>_UNCONNECTED ,
\NLW_blk00000001/blk0000020e_M<24>_UNCONNECTED , \NLW_blk00000001/blk0000020e_M<23>_UNCONNECTED , \NLW_blk00000001/blk0000020e_M<22>_UNCONNECTED ,
\NLW_blk00000001/blk0000020e_M<21>_UNCONNECTED , \NLW_blk00000001/blk0000020e_M<20>_UNCONNECTED , \NLW_blk00000001/blk0000020e_M<19>_UNCONNECTED ,
\NLW_blk00000001/blk0000020e_M<18>_UNCONNECTED , \NLW_blk00000001/blk0000020e_M<17>_UNCONNECTED , \NLW_blk00000001/blk0000020e_M<16>_UNCONNECTED ,
\NLW_blk00000001/blk0000020e_M<15>_UNCONNECTED , \NLW_blk00000001/blk0000020e_M<14>_UNCONNECTED , \NLW_blk00000001/blk0000020e_M<13>_UNCONNECTED ,
\NLW_blk00000001/blk0000020e_M<12>_UNCONNECTED , \NLW_blk00000001/blk0000020e_M<11>_UNCONNECTED , \NLW_blk00000001/blk0000020e_M<10>_UNCONNECTED ,
\NLW_blk00000001/blk0000020e_M<9>_UNCONNECTED , \NLW_blk00000001/blk0000020e_M<8>_UNCONNECTED , \NLW_blk00000001/blk0000020e_M<7>_UNCONNECTED ,
\NLW_blk00000001/blk0000020e_M<6>_UNCONNECTED , \NLW_blk00000001/blk0000020e_M<5>_UNCONNECTED , \NLW_blk00000001/blk0000020e_M<4>_UNCONNECTED ,
\NLW_blk00000001/blk0000020e_M<3>_UNCONNECTED , \NLW_blk00000001/blk0000020e_M<2>_UNCONNECTED , \NLW_blk00000001/blk0000020e_M<1>_UNCONNECTED ,
\NLW_blk00000001/blk0000020e_M<0>_UNCONNECTED })
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000020d  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000002a1 ),
    .Q(\blk00000001/sig00000397 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000020c  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000002a2 ),
    .Q(\blk00000001/sig00000398 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000020b  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000002a3 ),
    .Q(\blk00000001/sig00000399 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000020a  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000002a4 ),
    .Q(\blk00000001/sig0000039a )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000209  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000002a5 ),
    .Q(\blk00000001/sig0000039b )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000208  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000002a6 ),
    .Q(\blk00000001/sig0000039c )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000207  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000002a7 ),
    .Q(\blk00000001/sig0000039d )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000206  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000002a8 ),
    .Q(\blk00000001/sig0000039e )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000205  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000002a9 ),
    .Q(\blk00000001/sig0000039f )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000204  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000002aa ),
    .Q(\blk00000001/sig000003a0 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000203  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000002ab ),
    .Q(\blk00000001/sig000003a1 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000202  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000002ac ),
    .Q(\blk00000001/sig000003a2 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000201  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000002ad ),
    .Q(\blk00000001/sig000003a3 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000200  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000002ae ),
    .Q(\blk00000001/sig000003a4 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000001ff  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000002af ),
    .Q(\blk00000001/sig000003a5 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000001fe  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000284 ),
    .Q(\blk00000001/sig000003a6 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000001fd  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000284 ),
    .Q(\blk00000001/sig000003a7 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000001fc  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000002b0 ),
    .Q(\blk00000001/sig000003a8 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000001fb  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000002b1 ),
    .Q(\blk00000001/sig000003a9 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000001fa  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000002b2 ),
    .Q(\blk00000001/sig000003aa )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000001f9  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000002b3 ),
    .Q(\blk00000001/sig000003ab )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000001f8  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000002b4 ),
    .Q(\blk00000001/sig000003ac )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000001f7  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000002b5 ),
    .Q(\blk00000001/sig000003ad )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000001f6  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000002b6 ),
    .Q(\blk00000001/sig000003ae )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000001f5  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000002b7 ),
    .Q(\blk00000001/sig000003af )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000001f4  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000002b8 ),
    .Q(\blk00000001/sig000003b0 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000001f3  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000002b9 ),
    .Q(\blk00000001/sig000003b1 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000001f2  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000002ba ),
    .Q(\blk00000001/sig000003b2 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000001f1  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000002bb ),
    .Q(\blk00000001/sig000003b3 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000001f0  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000002bc ),
    .Q(\blk00000001/sig000003b4 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000001ef  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000002bd ),
    .Q(\blk00000001/sig000003b5 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000001ee  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000002be ),
    .Q(\blk00000001/sig000003b6 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000001ed  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000002bf ),
    .Q(\blk00000001/sig000003b7 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000001ec  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000284 ),
    .Q(\blk00000001/sig000003b8 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000001eb  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000284 ),
    .Q(\blk00000001/sig000003b9 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000001ea  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000284 ),
    .Q(\blk00000001/sig000003ba )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000001e9  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000284 ),
    .Q(\blk00000001/sig000003bb )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000001e8  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000284 ),
    .Q(\blk00000001/sig000003bc )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000001e7  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000284 ),
    .Q(\blk00000001/sig000003bd )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000001e6  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000284 ),
    .Q(\blk00000001/sig000003be )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000001e5  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000284 ),
    .Q(\blk00000001/sig000003bf )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000001e4  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000284 ),
    .Q(\blk00000001/sig000003c0 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000001e3  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000284 ),
    .Q(\blk00000001/sig000003c1 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000001e2  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000284 ),
    .Q(\blk00000001/sig000003c2 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000001e1  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000284 ),
    .Q(\blk00000001/sig000003c3 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000001e0  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000284 ),
    .Q(\blk00000001/sig000003c4 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000001df  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000284 ),
    .Q(\blk00000001/sig000003c5 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000001de  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000284 ),
    .Q(\blk00000001/sig000003c6 )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000001dd  (
    .C(aclk),
    .D(\blk00000001/sig0000003c ),
    .Q(\blk00000001/sig00000544 )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000001dc  (
    .C(aclk),
    .D(\blk00000001/sig0000031c ),
    .Q(\blk00000001/sig00000543 )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000001db  (
    .C(aclk),
    .D(\blk00000001/sig00000543 ),
    .Q(\blk00000001/sig00000491 )
  );
  DSP48A1 #(
    .A0REG ( 0 ),
    .A1REG ( 1 ),
    .B0REG ( 0 ),
    .B1REG ( 1 ),
    .CARRYINREG ( 0 ),
    .CARRYINSEL ( "OPMODE5" ),
    .CREG ( 1 ),
    .DREG ( 1 ),
    .MREG ( 1 ),
    .OPMODEREG ( 1 ),
    .PREG ( 1 ),
    .RSTTYPE ( "SYNC" ),
    .CARRYOUTREG ( 0 ))
  \blk00000001/blk000001da  (
    .CECARRYIN(\blk00000001/sig0000051d ),
    .RSTC(\blk00000001/sig0000051d ),
    .RSTCARRYIN(\blk00000001/sig0000051d ),
    .CED(\blk00000001/sig0000003a ),
    .RSTD(\blk00000001/sig0000051d ),
    .CEOPMODE(\blk00000001/sig0000003a ),
    .CEC(\blk00000001/sig0000003a ),
    .CARRYOUTF(\NLW_blk00000001/blk000001da_CARRYOUTF_UNCONNECTED ),
    .RSTOPMODE(\blk00000001/sig0000051d ),
    .RSTM(\blk00000001/sig0000051d ),
    .CLK(aclk),
    .RSTB(\blk00000001/sig0000051d ),
    .CEM(\blk00000001/sig0000003a ),
    .CEB(\blk00000001/sig0000003a ),
    .CARRYIN(\blk00000001/sig0000051d ),
    .CEP(\blk00000001/sig0000003a ),
    .CEA(\blk00000001/sig0000003a ),
    .CARRYOUT(\NLW_blk00000001/blk000001da_CARRYOUT_UNCONNECTED ),
    .RSTA(\blk00000001/sig0000051d ),
    .RSTP(\blk00000001/sig0000051d ),
    .B({\blk00000001/sig000003f7 , \blk00000001/sig000003f6 , \blk00000001/sig000003f5 , \blk00000001/sig000003f4 , \blk00000001/sig000003f3 ,
\blk00000001/sig000003f2 , \blk00000001/sig000003f1 , \blk00000001/sig000003f0 , \blk00000001/sig000003ef , \blk00000001/sig000003ee ,
\blk00000001/sig000003ed , \blk00000001/sig000003ec , \blk00000001/sig000003eb , \blk00000001/sig000003ea , \blk00000001/sig000003e9 ,
\blk00000001/sig000003e8 , \blk00000001/sig000003e7 , \blk00000001/sig0000051d }),
    .BCOUT({\NLW_blk00000001/blk000001da_BCOUT<17>_UNCONNECTED , \NLW_blk00000001/blk000001da_BCOUT<16>_UNCONNECTED ,
\NLW_blk00000001/blk000001da_BCOUT<15>_UNCONNECTED , \NLW_blk00000001/blk000001da_BCOUT<14>_UNCONNECTED ,
\NLW_blk00000001/blk000001da_BCOUT<13>_UNCONNECTED , \NLW_blk00000001/blk000001da_BCOUT<12>_UNCONNECTED ,
\NLW_blk00000001/blk000001da_BCOUT<11>_UNCONNECTED , \NLW_blk00000001/blk000001da_BCOUT<10>_UNCONNECTED ,
\NLW_blk00000001/blk000001da_BCOUT<9>_UNCONNECTED , \NLW_blk00000001/blk000001da_BCOUT<8>_UNCONNECTED ,
\NLW_blk00000001/blk000001da_BCOUT<7>_UNCONNECTED , \NLW_blk00000001/blk000001da_BCOUT<6>_UNCONNECTED ,
\NLW_blk00000001/blk000001da_BCOUT<5>_UNCONNECTED , \NLW_blk00000001/blk000001da_BCOUT<4>_UNCONNECTED ,
\NLW_blk00000001/blk000001da_BCOUT<3>_UNCONNECTED , \NLW_blk00000001/blk000001da_BCOUT<2>_UNCONNECTED ,
\NLW_blk00000001/blk000001da_BCOUT<1>_UNCONNECTED , \NLW_blk00000001/blk000001da_BCOUT<0>_UNCONNECTED }),
    .PCIN({\blk00000001/sig00000383 , \blk00000001/sig00000382 , \blk00000001/sig00000381 , \blk00000001/sig00000380 , \blk00000001/sig0000037f ,
\blk00000001/sig0000037e , \blk00000001/sig0000037d , \blk00000001/sig0000037c , \blk00000001/sig0000037b , \blk00000001/sig0000037a ,
\blk00000001/sig00000379 , \blk00000001/sig00000378 , \blk00000001/sig00000377 , \blk00000001/sig00000376 , \blk00000001/sig00000375 ,
\blk00000001/sig00000374 , \blk00000001/sig00000373 , \blk00000001/sig00000372 , \blk00000001/sig00000371 , \blk00000001/sig00000370 ,
\blk00000001/sig0000036f , \blk00000001/sig0000036e , \blk00000001/sig0000036d , \blk00000001/sig0000036c , \blk00000001/sig0000036b ,
\blk00000001/sig0000036a , \blk00000001/sig00000369 , \blk00000001/sig00000368 , \blk00000001/sig00000367 , \blk00000001/sig00000366 ,
\blk00000001/sig00000365 , \blk00000001/sig00000364 , \blk00000001/sig00000363 , \blk00000001/sig00000362 , \blk00000001/sig00000361 ,
\blk00000001/sig00000360 , \blk00000001/sig0000035f , \blk00000001/sig0000035e , \blk00000001/sig0000035d , \blk00000001/sig0000035c ,
\blk00000001/sig0000035b , \blk00000001/sig0000035a , \blk00000001/sig00000359 , \blk00000001/sig00000358 , \blk00000001/sig00000357 ,
\blk00000001/sig00000356 , \blk00000001/sig00000355 , \blk00000001/sig00000354 }),
    .C({\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d }),
    .P({\blk00000001/sig00000050 , \NLW_blk00000001/blk000001da_P<46>_UNCONNECTED , \NLW_blk00000001/blk000001da_P<45>_UNCONNECTED ,
\NLW_blk00000001/blk000001da_P<44>_UNCONNECTED , \NLW_blk00000001/blk000001da_P<43>_UNCONNECTED , \NLW_blk00000001/blk000001da_P<42>_UNCONNECTED ,
\NLW_blk00000001/blk000001da_P<41>_UNCONNECTED , \NLW_blk00000001/blk000001da_P<40>_UNCONNECTED , \NLW_blk00000001/blk000001da_P<39>_UNCONNECTED ,
\NLW_blk00000001/blk000001da_P<38>_UNCONNECTED , \NLW_blk00000001/blk000001da_P<37>_UNCONNECTED , \NLW_blk00000001/blk000001da_P<36>_UNCONNECTED ,
\NLW_blk00000001/blk000001da_P<35>_UNCONNECTED , \NLW_blk00000001/blk000001da_P<34>_UNCONNECTED , \blk00000001/sig0000004f , \blk00000001/sig0000004e
, \blk00000001/sig0000004d , \blk00000001/sig0000004c , \blk00000001/sig0000004b , \blk00000001/sig0000004a , \blk00000001/sig00000049 ,
\blk00000001/sig00000048 , \blk00000001/sig00000047 , \blk00000001/sig00000046 , \blk00000001/sig00000045 , \blk00000001/sig00000044 ,
\blk00000001/sig00000043 , \blk00000001/sig00000042 , \blk00000001/sig00000041 , \blk00000001/sig00000353 , \blk00000001/sig00000352 ,
\blk00000001/sig00000351 , \blk00000001/sig00000350 , \blk00000001/sig0000034f , \blk00000001/sig0000034e , \blk00000001/sig0000034d ,
\blk00000001/sig0000034c , \blk00000001/sig0000034b , \blk00000001/sig0000034a , \blk00000001/sig00000349 , \blk00000001/sig00000348 ,
\blk00000001/sig00000347 , \blk00000001/sig00000346 , \blk00000001/sig00000345 , \blk00000001/sig00000344 , \blk00000001/sig00000343 ,
\blk00000001/sig00000342 , \blk00000001/sig00000341 }),
    .OPMODE({\blk00000001/sig00000491 , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000003a , \blk00000001/sig0000051d , \blk00000001/sig0000003a }),
    .D({\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d }),
    .PCOUT({\NLW_blk00000001/blk000001da_PCOUT<47>_UNCONNECTED , \NLW_blk00000001/blk000001da_PCOUT<46>_UNCONNECTED ,
\NLW_blk00000001/blk000001da_PCOUT<45>_UNCONNECTED , \NLW_blk00000001/blk000001da_PCOUT<44>_UNCONNECTED ,
\NLW_blk00000001/blk000001da_PCOUT<43>_UNCONNECTED , \NLW_blk00000001/blk000001da_PCOUT<42>_UNCONNECTED ,
\NLW_blk00000001/blk000001da_PCOUT<41>_UNCONNECTED , \NLW_blk00000001/blk000001da_PCOUT<40>_UNCONNECTED ,
\NLW_blk00000001/blk000001da_PCOUT<39>_UNCONNECTED , \NLW_blk00000001/blk000001da_PCOUT<38>_UNCONNECTED ,
\NLW_blk00000001/blk000001da_PCOUT<37>_UNCONNECTED , \NLW_blk00000001/blk000001da_PCOUT<36>_UNCONNECTED ,
\NLW_blk00000001/blk000001da_PCOUT<35>_UNCONNECTED , \NLW_blk00000001/blk000001da_PCOUT<34>_UNCONNECTED ,
\NLW_blk00000001/blk000001da_PCOUT<33>_UNCONNECTED , \NLW_blk00000001/blk000001da_PCOUT<32>_UNCONNECTED ,
\NLW_blk00000001/blk000001da_PCOUT<31>_UNCONNECTED , \NLW_blk00000001/blk000001da_PCOUT<30>_UNCONNECTED ,
\NLW_blk00000001/blk000001da_PCOUT<29>_UNCONNECTED , \NLW_blk00000001/blk000001da_PCOUT<28>_UNCONNECTED ,
\NLW_blk00000001/blk000001da_PCOUT<27>_UNCONNECTED , \NLW_blk00000001/blk000001da_PCOUT<26>_UNCONNECTED ,
\NLW_blk00000001/blk000001da_PCOUT<25>_UNCONNECTED , \NLW_blk00000001/blk000001da_PCOUT<24>_UNCONNECTED ,
\NLW_blk00000001/blk000001da_PCOUT<23>_UNCONNECTED , \NLW_blk00000001/blk000001da_PCOUT<22>_UNCONNECTED ,
\NLW_blk00000001/blk000001da_PCOUT<21>_UNCONNECTED , \NLW_blk00000001/blk000001da_PCOUT<20>_UNCONNECTED ,
\NLW_blk00000001/blk000001da_PCOUT<19>_UNCONNECTED , \NLW_blk00000001/blk000001da_PCOUT<18>_UNCONNECTED ,
\NLW_blk00000001/blk000001da_PCOUT<17>_UNCONNECTED , \NLW_blk00000001/blk000001da_PCOUT<16>_UNCONNECTED ,
\NLW_blk00000001/blk000001da_PCOUT<15>_UNCONNECTED , \NLW_blk00000001/blk000001da_PCOUT<14>_UNCONNECTED ,
\NLW_blk00000001/blk000001da_PCOUT<13>_UNCONNECTED , \NLW_blk00000001/blk000001da_PCOUT<12>_UNCONNECTED ,
\NLW_blk00000001/blk000001da_PCOUT<11>_UNCONNECTED , \NLW_blk00000001/blk000001da_PCOUT<10>_UNCONNECTED ,
\NLW_blk00000001/blk000001da_PCOUT<9>_UNCONNECTED , \NLW_blk00000001/blk000001da_PCOUT<8>_UNCONNECTED ,
\NLW_blk00000001/blk000001da_PCOUT<7>_UNCONNECTED , \NLW_blk00000001/blk000001da_PCOUT<6>_UNCONNECTED ,
\NLW_blk00000001/blk000001da_PCOUT<5>_UNCONNECTED , \NLW_blk00000001/blk000001da_PCOUT<4>_UNCONNECTED ,
\NLW_blk00000001/blk000001da_PCOUT<3>_UNCONNECTED , \NLW_blk00000001/blk000001da_PCOUT<2>_UNCONNECTED ,
\NLW_blk00000001/blk000001da_PCOUT<1>_UNCONNECTED , \NLW_blk00000001/blk000001da_PCOUT<0>_UNCONNECTED }),
    .A({\blk00000001/sig00000490 , \blk00000001/sig0000048f , \blk00000001/sig0000048e , \blk00000001/sig0000048d , \blk00000001/sig0000048c ,
\blk00000001/sig0000048b , \blk00000001/sig0000048a , \blk00000001/sig00000489 , \blk00000001/sig00000488 , \blk00000001/sig00000487 ,
\blk00000001/sig00000486 , \blk00000001/sig00000485 , \blk00000001/sig00000484 , \blk00000001/sig00000483 , \blk00000001/sig00000482 ,
\blk00000001/sig00000481 , \blk00000001/sig00000480 , \blk00000001/sig0000047f }),
    .M({\NLW_blk00000001/blk000001da_M<35>_UNCONNECTED , \NLW_blk00000001/blk000001da_M<34>_UNCONNECTED ,
\NLW_blk00000001/blk000001da_M<33>_UNCONNECTED , \NLW_blk00000001/blk000001da_M<32>_UNCONNECTED , \NLW_blk00000001/blk000001da_M<31>_UNCONNECTED ,
\NLW_blk00000001/blk000001da_M<30>_UNCONNECTED , \NLW_blk00000001/blk000001da_M<29>_UNCONNECTED , \NLW_blk00000001/blk000001da_M<28>_UNCONNECTED ,
\NLW_blk00000001/blk000001da_M<27>_UNCONNECTED , \NLW_blk00000001/blk000001da_M<26>_UNCONNECTED , \NLW_blk00000001/blk000001da_M<25>_UNCONNECTED ,
\NLW_blk00000001/blk000001da_M<24>_UNCONNECTED , \NLW_blk00000001/blk000001da_M<23>_UNCONNECTED , \NLW_blk00000001/blk000001da_M<22>_UNCONNECTED ,
\NLW_blk00000001/blk000001da_M<21>_UNCONNECTED , \NLW_blk00000001/blk000001da_M<20>_UNCONNECTED , \NLW_blk00000001/blk000001da_M<19>_UNCONNECTED ,
\NLW_blk00000001/blk000001da_M<18>_UNCONNECTED , \NLW_blk00000001/blk000001da_M<17>_UNCONNECTED , \NLW_blk00000001/blk000001da_M<16>_UNCONNECTED ,
\NLW_blk00000001/blk000001da_M<15>_UNCONNECTED , \NLW_blk00000001/blk000001da_M<14>_UNCONNECTED , \NLW_blk00000001/blk000001da_M<13>_UNCONNECTED ,
\NLW_blk00000001/blk000001da_M<12>_UNCONNECTED , \NLW_blk00000001/blk000001da_M<11>_UNCONNECTED , \NLW_blk00000001/blk000001da_M<10>_UNCONNECTED ,
\NLW_blk00000001/blk000001da_M<9>_UNCONNECTED , \NLW_blk00000001/blk000001da_M<8>_UNCONNECTED , \NLW_blk00000001/blk000001da_M<7>_UNCONNECTED ,
\NLW_blk00000001/blk000001da_M<6>_UNCONNECTED , \NLW_blk00000001/blk000001da_M<5>_UNCONNECTED , \NLW_blk00000001/blk000001da_M<4>_UNCONNECTED ,
\NLW_blk00000001/blk000001da_M<3>_UNCONNECTED , \NLW_blk00000001/blk000001da_M<2>_UNCONNECTED , \NLW_blk00000001/blk000001da_M<1>_UNCONNECTED ,
\NLW_blk00000001/blk000001da_M<0>_UNCONNECTED })
  );
  DSP48A1 #(
    .A0REG ( 0 ),
    .A1REG ( 1 ),
    .B0REG ( 0 ),
    .B1REG ( 1 ),
    .CARRYINREG ( 0 ),
    .CARRYINSEL ( "OPMODE5" ),
    .CREG ( 1 ),
    .DREG ( 1 ),
    .MREG ( 1 ),
    .OPMODEREG ( 1 ),
    .PREG ( 1 ),
    .RSTTYPE ( "SYNC" ),
    .CARRYOUTREG ( 0 ))
  \blk00000001/blk000001d9  (
    .CECARRYIN(\blk00000001/sig0000051d ),
    .RSTC(\blk00000001/sig0000051d ),
    .RSTCARRYIN(\blk00000001/sig0000051d ),
    .CED(\blk00000001/sig0000003a ),
    .RSTD(\blk00000001/sig0000051d ),
    .CEOPMODE(\blk00000001/sig0000003a ),
    .CEC(\blk00000001/sig0000003a ),
    .CARRYOUTF(\NLW_blk00000001/blk000001d9_CARRYOUTF_UNCONNECTED ),
    .RSTOPMODE(\blk00000001/sig0000051d ),
    .RSTM(\blk00000001/sig0000051d ),
    .CLK(aclk),
    .RSTB(\blk00000001/sig0000051d ),
    .CEM(\blk00000001/sig0000003a ),
    .CEB(\blk00000001/sig0000003a ),
    .CARRYIN(\blk00000001/sig0000051d ),
    .CEP(\blk00000001/sig0000003a ),
    .CEA(\blk00000001/sig0000003a ),
    .CARRYOUT(\NLW_blk00000001/blk000001d9_CARRYOUT_UNCONNECTED ),
    .RSTA(\blk00000001/sig0000051d ),
    .RSTP(\blk00000001/sig0000051d ),
    .B({\blk00000001/sig0000051d , \blk00000001/sig0000047d , \blk00000001/sig0000047c , \blk00000001/sig0000047b , \blk00000001/sig0000047a ,
\blk00000001/sig00000479 , \blk00000001/sig00000478 , \blk00000001/sig00000477 , \blk00000001/sig00000476 , \blk00000001/sig00000475 ,
\blk00000001/sig00000474 , \blk00000001/sig00000473 , \blk00000001/sig00000472 , \blk00000001/sig00000471 , \blk00000001/sig00000470 ,
\blk00000001/sig0000046f , \blk00000001/sig0000046e , \blk00000001/sig0000051d }),
    .BCOUT({\NLW_blk00000001/blk000001d9_BCOUT<17>_UNCONNECTED , \NLW_blk00000001/blk000001d9_BCOUT<16>_UNCONNECTED ,
\NLW_blk00000001/blk000001d9_BCOUT<15>_UNCONNECTED , \NLW_blk00000001/blk000001d9_BCOUT<14>_UNCONNECTED ,
\NLW_blk00000001/blk000001d9_BCOUT<13>_UNCONNECTED , \NLW_blk00000001/blk000001d9_BCOUT<12>_UNCONNECTED ,
\NLW_blk00000001/blk000001d9_BCOUT<11>_UNCONNECTED , \NLW_blk00000001/blk000001d9_BCOUT<10>_UNCONNECTED ,
\NLW_blk00000001/blk000001d9_BCOUT<9>_UNCONNECTED , \NLW_blk00000001/blk000001d9_BCOUT<8>_UNCONNECTED ,
\NLW_blk00000001/blk000001d9_BCOUT<7>_UNCONNECTED , \NLW_blk00000001/blk000001d9_BCOUT<6>_UNCONNECTED ,
\NLW_blk00000001/blk000001d9_BCOUT<5>_UNCONNECTED , \NLW_blk00000001/blk000001d9_BCOUT<4>_UNCONNECTED ,
\NLW_blk00000001/blk000001d9_BCOUT<3>_UNCONNECTED , \NLW_blk00000001/blk000001d9_BCOUT<2>_UNCONNECTED ,
\NLW_blk00000001/blk000001d9_BCOUT<1>_UNCONNECTED , \NLW_blk00000001/blk000001d9_BCOUT<0>_UNCONNECTED }),
    .PCIN({\blk00000001/sig0000043a , \blk00000001/sig00000439 , \blk00000001/sig00000438 , \blk00000001/sig00000437 , \blk00000001/sig00000436 ,
\blk00000001/sig00000435 , \blk00000001/sig00000434 , \blk00000001/sig00000433 , \blk00000001/sig00000432 , \blk00000001/sig00000431 ,
\blk00000001/sig00000430 , \blk00000001/sig0000042f , \blk00000001/sig0000042e , \blk00000001/sig0000042d , \blk00000001/sig0000042c ,
\blk00000001/sig0000042b , \blk00000001/sig0000042a , \blk00000001/sig00000429 , \blk00000001/sig00000428 , \blk00000001/sig00000427 ,
\blk00000001/sig00000426 , \blk00000001/sig00000425 , \blk00000001/sig00000424 , \blk00000001/sig00000423 , \blk00000001/sig00000422 ,
\blk00000001/sig00000421 , \blk00000001/sig00000420 , \blk00000001/sig0000041f , \blk00000001/sig0000041e , \blk00000001/sig0000041d ,
\blk00000001/sig0000041c , \blk00000001/sig0000041b , \blk00000001/sig0000041a , \blk00000001/sig00000419 , \blk00000001/sig00000418 ,
\blk00000001/sig00000417 , \blk00000001/sig00000416 , \blk00000001/sig00000415 , \blk00000001/sig00000414 , \blk00000001/sig00000413 ,
\blk00000001/sig00000412 , \blk00000001/sig00000411 , \blk00000001/sig00000410 , \blk00000001/sig0000040f , \blk00000001/sig0000040e ,
\blk00000001/sig0000040d , \blk00000001/sig0000040c , \blk00000001/sig0000040b }),
    .C({\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d }),
    .P({\NLW_blk00000001/blk000001d9_P<47>_UNCONNECTED , \NLW_blk00000001/blk000001d9_P<46>_UNCONNECTED ,
\NLW_blk00000001/blk000001d9_P<45>_UNCONNECTED , \NLW_blk00000001/blk000001d9_P<44>_UNCONNECTED , \NLW_blk00000001/blk000001d9_P<43>_UNCONNECTED ,
\NLW_blk00000001/blk000001d9_P<42>_UNCONNECTED , \NLW_blk00000001/blk000001d9_P<41>_UNCONNECTED , \NLW_blk00000001/blk000001d9_P<40>_UNCONNECTED ,
\NLW_blk00000001/blk000001d9_P<39>_UNCONNECTED , \NLW_blk00000001/blk000001d9_P<38>_UNCONNECTED , \NLW_blk00000001/blk000001d9_P<37>_UNCONNECTED ,
\NLW_blk00000001/blk000001d9_P<36>_UNCONNECTED , \NLW_blk00000001/blk000001d9_P<35>_UNCONNECTED , \NLW_blk00000001/blk000001d9_P<34>_UNCONNECTED ,
\NLW_blk00000001/blk000001d9_P<33>_UNCONNECTED , \NLW_blk00000001/blk000001d9_P<32>_UNCONNECTED , \NLW_blk00000001/blk000001d9_P<31>_UNCONNECTED ,
\NLW_blk00000001/blk000001d9_P<30>_UNCONNECTED , \NLW_blk00000001/blk000001d9_P<29>_UNCONNECTED , \NLW_blk00000001/blk000001d9_P<28>_UNCONNECTED ,
\NLW_blk00000001/blk000001d9_P<27>_UNCONNECTED , \NLW_blk00000001/blk000001d9_P<26>_UNCONNECTED , \NLW_blk00000001/blk000001d9_P<25>_UNCONNECTED ,
\NLW_blk00000001/blk000001d9_P<24>_UNCONNECTED , \NLW_blk00000001/blk000001d9_P<23>_UNCONNECTED , \NLW_blk00000001/blk000001d9_P<22>_UNCONNECTED ,
\NLW_blk00000001/blk000001d9_P<21>_UNCONNECTED , \NLW_blk00000001/blk000001d9_P<20>_UNCONNECTED , \NLW_blk00000001/blk000001d9_P<19>_UNCONNECTED ,
\blk00000001/sig0000040a , \blk00000001/sig00000409 , \blk00000001/sig00000408 , \blk00000001/sig00000407 , \blk00000001/sig00000406 ,
\blk00000001/sig00000405 , \blk00000001/sig00000404 , \blk00000001/sig00000403 , \blk00000001/sig00000402 , \blk00000001/sig00000401 ,
\blk00000001/sig00000400 , \blk00000001/sig000003ff , \blk00000001/sig000003fe , \blk00000001/sig000003fd , \blk00000001/sig000003fc ,
\blk00000001/sig000003fb , \blk00000001/sig000003fa , \blk00000001/sig000003f9 , \blk00000001/sig000003f8 }),
    .OPMODE({\blk00000001/sig00000491 , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000003a , \blk00000001/sig0000051d , \blk00000001/sig0000003a }),
    .D({\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d }),
    .PCOUT({\NLW_blk00000001/blk000001d9_PCOUT<47>_UNCONNECTED , \NLW_blk00000001/blk000001d9_PCOUT<46>_UNCONNECTED ,
\NLW_blk00000001/blk000001d9_PCOUT<45>_UNCONNECTED , \NLW_blk00000001/blk000001d9_PCOUT<44>_UNCONNECTED ,
\NLW_blk00000001/blk000001d9_PCOUT<43>_UNCONNECTED , \NLW_blk00000001/blk000001d9_PCOUT<42>_UNCONNECTED ,
\NLW_blk00000001/blk000001d9_PCOUT<41>_UNCONNECTED , \NLW_blk00000001/blk000001d9_PCOUT<40>_UNCONNECTED ,
\NLW_blk00000001/blk000001d9_PCOUT<39>_UNCONNECTED , \NLW_blk00000001/blk000001d9_PCOUT<38>_UNCONNECTED ,
\NLW_blk00000001/blk000001d9_PCOUT<37>_UNCONNECTED , \NLW_blk00000001/blk000001d9_PCOUT<36>_UNCONNECTED ,
\NLW_blk00000001/blk000001d9_PCOUT<35>_UNCONNECTED , \NLW_blk00000001/blk000001d9_PCOUT<34>_UNCONNECTED ,
\NLW_blk00000001/blk000001d9_PCOUT<33>_UNCONNECTED , \NLW_blk00000001/blk000001d9_PCOUT<32>_UNCONNECTED ,
\NLW_blk00000001/blk000001d9_PCOUT<31>_UNCONNECTED , \NLW_blk00000001/blk000001d9_PCOUT<30>_UNCONNECTED ,
\NLW_blk00000001/blk000001d9_PCOUT<29>_UNCONNECTED , \NLW_blk00000001/blk000001d9_PCOUT<28>_UNCONNECTED ,
\NLW_blk00000001/blk000001d9_PCOUT<27>_UNCONNECTED , \NLW_blk00000001/blk000001d9_PCOUT<26>_UNCONNECTED ,
\NLW_blk00000001/blk000001d9_PCOUT<25>_UNCONNECTED , \NLW_blk00000001/blk000001d9_PCOUT<24>_UNCONNECTED ,
\NLW_blk00000001/blk000001d9_PCOUT<23>_UNCONNECTED , \NLW_blk00000001/blk000001d9_PCOUT<22>_UNCONNECTED ,
\NLW_blk00000001/blk000001d9_PCOUT<21>_UNCONNECTED , \NLW_blk00000001/blk000001d9_PCOUT<20>_UNCONNECTED ,
\NLW_blk00000001/blk000001d9_PCOUT<19>_UNCONNECTED , \NLW_blk00000001/blk000001d9_PCOUT<18>_UNCONNECTED ,
\NLW_blk00000001/blk000001d9_PCOUT<17>_UNCONNECTED , \NLW_blk00000001/blk000001d9_PCOUT<16>_UNCONNECTED ,
\NLW_blk00000001/blk000001d9_PCOUT<15>_UNCONNECTED , \NLW_blk00000001/blk000001d9_PCOUT<14>_UNCONNECTED ,
\NLW_blk00000001/blk000001d9_PCOUT<13>_UNCONNECTED , \NLW_blk00000001/blk000001d9_PCOUT<12>_UNCONNECTED ,
\NLW_blk00000001/blk000001d9_PCOUT<11>_UNCONNECTED , \NLW_blk00000001/blk000001d9_PCOUT<10>_UNCONNECTED ,
\NLW_blk00000001/blk000001d9_PCOUT<9>_UNCONNECTED , \NLW_blk00000001/blk000001d9_PCOUT<8>_UNCONNECTED ,
\NLW_blk00000001/blk000001d9_PCOUT<7>_UNCONNECTED , \NLW_blk00000001/blk000001d9_PCOUT<6>_UNCONNECTED ,
\NLW_blk00000001/blk000001d9_PCOUT<5>_UNCONNECTED , \NLW_blk00000001/blk000001d9_PCOUT<4>_UNCONNECTED ,
\NLW_blk00000001/blk000001d9_PCOUT<3>_UNCONNECTED , \NLW_blk00000001/blk000001d9_PCOUT<2>_UNCONNECTED ,
\NLW_blk00000001/blk000001d9_PCOUT<1>_UNCONNECTED , \NLW_blk00000001/blk000001d9_PCOUT<0>_UNCONNECTED }),
    .A({\blk00000001/sig00000490 , \blk00000001/sig0000048f , \blk00000001/sig0000048e , \blk00000001/sig0000048d , \blk00000001/sig0000048c ,
\blk00000001/sig0000048b , \blk00000001/sig0000048a , \blk00000001/sig00000489 , \blk00000001/sig00000488 , \blk00000001/sig00000487 ,
\blk00000001/sig00000486 , \blk00000001/sig00000485 , \blk00000001/sig00000484 , \blk00000001/sig00000483 , \blk00000001/sig00000482 ,
\blk00000001/sig00000481 , \blk00000001/sig00000480 , \blk00000001/sig0000047f }),
    .M({\NLW_blk00000001/blk000001d9_M<35>_UNCONNECTED , \NLW_blk00000001/blk000001d9_M<34>_UNCONNECTED ,
\NLW_blk00000001/blk000001d9_M<33>_UNCONNECTED , \NLW_blk00000001/blk000001d9_M<32>_UNCONNECTED , \NLW_blk00000001/blk000001d9_M<31>_UNCONNECTED ,
\NLW_blk00000001/blk000001d9_M<30>_UNCONNECTED , \NLW_blk00000001/blk000001d9_M<29>_UNCONNECTED , \NLW_blk00000001/blk000001d9_M<28>_UNCONNECTED ,
\NLW_blk00000001/blk000001d9_M<27>_UNCONNECTED , \NLW_blk00000001/blk000001d9_M<26>_UNCONNECTED , \NLW_blk00000001/blk000001d9_M<25>_UNCONNECTED ,
\NLW_blk00000001/blk000001d9_M<24>_UNCONNECTED , \NLW_blk00000001/blk000001d9_M<23>_UNCONNECTED , \NLW_blk00000001/blk000001d9_M<22>_UNCONNECTED ,
\NLW_blk00000001/blk000001d9_M<21>_UNCONNECTED , \NLW_blk00000001/blk000001d9_M<20>_UNCONNECTED , \NLW_blk00000001/blk000001d9_M<19>_UNCONNECTED ,
\NLW_blk00000001/blk000001d9_M<18>_UNCONNECTED , \NLW_blk00000001/blk000001d9_M<17>_UNCONNECTED , \NLW_blk00000001/blk000001d9_M<16>_UNCONNECTED ,
\NLW_blk00000001/blk000001d9_M<15>_UNCONNECTED , \NLW_blk00000001/blk000001d9_M<14>_UNCONNECTED , \NLW_blk00000001/blk000001d9_M<13>_UNCONNECTED ,
\NLW_blk00000001/blk000001d9_M<12>_UNCONNECTED , \NLW_blk00000001/blk000001d9_M<11>_UNCONNECTED , \NLW_blk00000001/blk000001d9_M<10>_UNCONNECTED ,
\NLW_blk00000001/blk000001d9_M<9>_UNCONNECTED , \NLW_blk00000001/blk000001d9_M<8>_UNCONNECTED , \NLW_blk00000001/blk000001d9_M<7>_UNCONNECTED ,
\NLW_blk00000001/blk000001d9_M<6>_UNCONNECTED , \NLW_blk00000001/blk000001d9_M<5>_UNCONNECTED , \NLW_blk00000001/blk000001d9_M<4>_UNCONNECTED ,
\NLW_blk00000001/blk000001d9_M<3>_UNCONNECTED , \NLW_blk00000001/blk000001d9_M<2>_UNCONNECTED , \NLW_blk00000001/blk000001d9_M<1>_UNCONNECTED ,
\NLW_blk00000001/blk000001d9_M<0>_UNCONNECTED })
  );
  DSP48A1 #(
    .A0REG ( 0 ),
    .A1REG ( 1 ),
    .B0REG ( 0 ),
    .B1REG ( 1 ),
    .CARRYINREG ( 0 ),
    .CARRYINSEL ( "OPMODE5" ),
    .CREG ( 1 ),
    .DREG ( 1 ),
    .MREG ( 1 ),
    .OPMODEREG ( 1 ),
    .PREG ( 1 ),
    .RSTTYPE ( "SYNC" ),
    .CARRYOUTREG ( 0 ))
  \blk00000001/blk000001d8  (
    .CECARRYIN(\blk00000001/sig0000051d ),
    .RSTC(\blk00000001/sig0000051d ),
    .RSTCARRYIN(\blk00000001/sig0000051d ),
    .CED(\blk00000001/sig0000003a ),
    .RSTD(\blk00000001/sig0000051d ),
    .CEOPMODE(\blk00000001/sig0000003a ),
    .CEC(\blk00000001/sig0000003a ),
    .CARRYOUTF(\NLW_blk00000001/blk000001d8_CARRYOUTF_UNCONNECTED ),
    .RSTOPMODE(\blk00000001/sig0000051d ),
    .RSTM(\blk00000001/sig0000051d ),
    .CLK(aclk),
    .RSTB(\blk00000001/sig0000051d ),
    .CEM(\blk00000001/sig0000003a ),
    .CEB(\blk00000001/sig0000003a ),
    .CARRYIN(\blk00000001/sig0000051d ),
    .CEP(\blk00000001/sig0000003a ),
    .CEA(\blk00000001/sig0000003a ),
    .CARRYOUT(\NLW_blk00000001/blk000001d8_CARRYOUT_UNCONNECTED ),
    .RSTA(\blk00000001/sig0000051d ),
    .RSTP(\blk00000001/sig0000051d ),
    .B({\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig00000526 , \blk00000001/sig00000525 , \blk00000001/sig00000524 ,
\blk00000001/sig00000523 , \blk00000001/sig00000522 , \blk00000001/sig00000521 , \blk00000001/sig00000520 , \blk00000001/sig0000051f ,
\blk00000001/sig0000051e , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d }),
    .BCOUT({\NLW_blk00000001/blk000001d8_BCOUT<17>_UNCONNECTED , \NLW_blk00000001/blk000001d8_BCOUT<16>_UNCONNECTED ,
\NLW_blk00000001/blk000001d8_BCOUT<15>_UNCONNECTED , \NLW_blk00000001/blk000001d8_BCOUT<14>_UNCONNECTED ,
\NLW_blk00000001/blk000001d8_BCOUT<13>_UNCONNECTED , \NLW_blk00000001/blk000001d8_BCOUT<12>_UNCONNECTED ,
\NLW_blk00000001/blk000001d8_BCOUT<11>_UNCONNECTED , \NLW_blk00000001/blk000001d8_BCOUT<10>_UNCONNECTED ,
\NLW_blk00000001/blk000001d8_BCOUT<9>_UNCONNECTED , \NLW_blk00000001/blk000001d8_BCOUT<8>_UNCONNECTED ,
\NLW_blk00000001/blk000001d8_BCOUT<7>_UNCONNECTED , \NLW_blk00000001/blk000001d8_BCOUT<6>_UNCONNECTED ,
\NLW_blk00000001/blk000001d8_BCOUT<5>_UNCONNECTED , \NLW_blk00000001/blk000001d8_BCOUT<4>_UNCONNECTED ,
\NLW_blk00000001/blk000001d8_BCOUT<3>_UNCONNECTED , \NLW_blk00000001/blk000001d8_BCOUT<2>_UNCONNECTED ,
\NLW_blk00000001/blk000001d8_BCOUT<1>_UNCONNECTED , \NLW_blk00000001/blk000001d8_BCOUT<0>_UNCONNECTED }),
    .PCIN({\blk00000001/sig000004e3 , \blk00000001/sig000004e2 , \blk00000001/sig000004e1 , \blk00000001/sig000004e0 , \blk00000001/sig000004df ,
\blk00000001/sig000004de , \blk00000001/sig000004dd , \blk00000001/sig000004dc , \blk00000001/sig000004db , \blk00000001/sig000004da ,
\blk00000001/sig000004d9 , \blk00000001/sig000004d8 , \blk00000001/sig000004d7 , \blk00000001/sig000004d6 , \blk00000001/sig000004d5 ,
\blk00000001/sig000004d4 , \blk00000001/sig000004d3 , \blk00000001/sig000004d2 , \blk00000001/sig000004d1 , \blk00000001/sig000004d0 ,
\blk00000001/sig000004cf , \blk00000001/sig000004ce , \blk00000001/sig000004cd , \blk00000001/sig000004cc , \blk00000001/sig000004cb ,
\blk00000001/sig000004ca , \blk00000001/sig000004c9 , \blk00000001/sig000004c8 , \blk00000001/sig000004c7 , \blk00000001/sig000004c6 ,
\blk00000001/sig000004c5 , \blk00000001/sig000004c4 , \blk00000001/sig000004c3 , \blk00000001/sig000004c2 , \blk00000001/sig000004c1 ,
\blk00000001/sig000004c0 , \blk00000001/sig000004bf , \blk00000001/sig000004be , \blk00000001/sig000004bd , \blk00000001/sig000004bc ,
\blk00000001/sig000004bb , \blk00000001/sig000004ba , \blk00000001/sig000004b9 , \blk00000001/sig000004b8 , \blk00000001/sig000004b7 ,
\blk00000001/sig000004b6 , \blk00000001/sig000004b5 , \blk00000001/sig000004b4 }),
    .C({\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d }),
    .P({\NLW_blk00000001/blk000001d8_P<47>_UNCONNECTED , \NLW_blk00000001/blk000001d8_P<46>_UNCONNECTED ,
\NLW_blk00000001/blk000001d8_P<45>_UNCONNECTED , \NLW_blk00000001/blk000001d8_P<44>_UNCONNECTED , \NLW_blk00000001/blk000001d8_P<43>_UNCONNECTED ,
\NLW_blk00000001/blk000001d8_P<42>_UNCONNECTED , \NLW_blk00000001/blk000001d8_P<41>_UNCONNECTED , \NLW_blk00000001/blk000001d8_P<40>_UNCONNECTED ,
\NLW_blk00000001/blk000001d8_P<39>_UNCONNECTED , \NLW_blk00000001/blk000001d8_P<38>_UNCONNECTED , \NLW_blk00000001/blk000001d8_P<37>_UNCONNECTED ,
\NLW_blk00000001/blk000001d8_P<36>_UNCONNECTED , \NLW_blk00000001/blk000001d8_P<35>_UNCONNECTED , \NLW_blk00000001/blk000001d8_P<34>_UNCONNECTED ,
\blk00000001/sig000004b3 , \blk00000001/sig000004b2 , \blk00000001/sig000004b1 , \blk00000001/sig000004b0 , \blk00000001/sig000004af ,
\blk00000001/sig000004ae , \blk00000001/sig000004ad , \blk00000001/sig000004ac , \blk00000001/sig000004ab , \blk00000001/sig000004aa ,
\blk00000001/sig000004a9 , \blk00000001/sig000004a8 , \blk00000001/sig000004a7 , \blk00000001/sig000004a6 , \blk00000001/sig000004a5 ,
\blk00000001/sig000004a4 , \blk00000001/sig000004a3 , \blk00000001/sig000004a2 , \blk00000001/sig000004a1 , \blk00000001/sig000004a0 ,
\blk00000001/sig0000049f , \blk00000001/sig0000049e , \blk00000001/sig0000049d , \blk00000001/sig0000049c , \blk00000001/sig0000049b ,
\blk00000001/sig0000049a , \blk00000001/sig00000499 , \blk00000001/sig00000498 , \blk00000001/sig00000497 , \blk00000001/sig00000496 ,
\blk00000001/sig00000495 , \blk00000001/sig00000494 , \blk00000001/sig00000493 , \blk00000001/sig00000492 }),
    .OPMODE({\blk00000001/sig000004e4 , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000003a , \blk00000001/sig0000051d , \blk00000001/sig0000003a }),
    .D({\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d }),
    .PCOUT({\NLW_blk00000001/blk000001d8_PCOUT<47>_UNCONNECTED , \NLW_blk00000001/blk000001d8_PCOUT<46>_UNCONNECTED ,
\NLW_blk00000001/blk000001d8_PCOUT<45>_UNCONNECTED , \NLW_blk00000001/blk000001d8_PCOUT<44>_UNCONNECTED ,
\NLW_blk00000001/blk000001d8_PCOUT<43>_UNCONNECTED , \NLW_blk00000001/blk000001d8_PCOUT<42>_UNCONNECTED ,
\NLW_blk00000001/blk000001d8_PCOUT<41>_UNCONNECTED , \NLW_blk00000001/blk000001d8_PCOUT<40>_UNCONNECTED ,
\NLW_blk00000001/blk000001d8_PCOUT<39>_UNCONNECTED , \NLW_blk00000001/blk000001d8_PCOUT<38>_UNCONNECTED ,
\NLW_blk00000001/blk000001d8_PCOUT<37>_UNCONNECTED , \NLW_blk00000001/blk000001d8_PCOUT<36>_UNCONNECTED ,
\NLW_blk00000001/blk000001d8_PCOUT<35>_UNCONNECTED , \NLW_blk00000001/blk000001d8_PCOUT<34>_UNCONNECTED ,
\NLW_blk00000001/blk000001d8_PCOUT<33>_UNCONNECTED , \NLW_blk00000001/blk000001d8_PCOUT<32>_UNCONNECTED ,
\NLW_blk00000001/blk000001d8_PCOUT<31>_UNCONNECTED , \NLW_blk00000001/blk000001d8_PCOUT<30>_UNCONNECTED ,
\NLW_blk00000001/blk000001d8_PCOUT<29>_UNCONNECTED , \NLW_blk00000001/blk000001d8_PCOUT<28>_UNCONNECTED ,
\NLW_blk00000001/blk000001d8_PCOUT<27>_UNCONNECTED , \NLW_blk00000001/blk000001d8_PCOUT<26>_UNCONNECTED ,
\NLW_blk00000001/blk000001d8_PCOUT<25>_UNCONNECTED , \NLW_blk00000001/blk000001d8_PCOUT<24>_UNCONNECTED ,
\NLW_blk00000001/blk000001d8_PCOUT<23>_UNCONNECTED , \NLW_blk00000001/blk000001d8_PCOUT<22>_UNCONNECTED ,
\NLW_blk00000001/blk000001d8_PCOUT<21>_UNCONNECTED , \NLW_blk00000001/blk000001d8_PCOUT<20>_UNCONNECTED ,
\NLW_blk00000001/blk000001d8_PCOUT<19>_UNCONNECTED , \NLW_blk00000001/blk000001d8_PCOUT<18>_UNCONNECTED ,
\NLW_blk00000001/blk000001d8_PCOUT<17>_UNCONNECTED , \NLW_blk00000001/blk000001d8_PCOUT<16>_UNCONNECTED ,
\NLW_blk00000001/blk000001d8_PCOUT<15>_UNCONNECTED , \NLW_blk00000001/blk000001d8_PCOUT<14>_UNCONNECTED ,
\NLW_blk00000001/blk000001d8_PCOUT<13>_UNCONNECTED , \NLW_blk00000001/blk000001d8_PCOUT<12>_UNCONNECTED ,
\NLW_blk00000001/blk000001d8_PCOUT<11>_UNCONNECTED , \NLW_blk00000001/blk000001d8_PCOUT<10>_UNCONNECTED ,
\NLW_blk00000001/blk000001d8_PCOUT<9>_UNCONNECTED , \NLW_blk00000001/blk000001d8_PCOUT<8>_UNCONNECTED ,
\NLW_blk00000001/blk000001d8_PCOUT<7>_UNCONNECTED , \NLW_blk00000001/blk000001d8_PCOUT<6>_UNCONNECTED ,
\NLW_blk00000001/blk000001d8_PCOUT<5>_UNCONNECTED , \NLW_blk00000001/blk000001d8_PCOUT<4>_UNCONNECTED ,
\NLW_blk00000001/blk000001d8_PCOUT<3>_UNCONNECTED , \NLW_blk00000001/blk000001d8_PCOUT<2>_UNCONNECTED ,
\NLW_blk00000001/blk000001d8_PCOUT<1>_UNCONNECTED , \NLW_blk00000001/blk000001d8_PCOUT<0>_UNCONNECTED }),
    .A({\blk00000001/sig0000051c , \blk00000001/sig0000051b , \blk00000001/sig0000051a , \blk00000001/sig00000519 , \blk00000001/sig00000518 ,
\blk00000001/sig00000517 , \blk00000001/sig00000516 , \blk00000001/sig00000515 , \blk00000001/sig00000514 , \blk00000001/sig00000513 ,
\blk00000001/sig00000512 , \blk00000001/sig00000511 , \blk00000001/sig00000510 , \blk00000001/sig0000050f , \blk00000001/sig0000050e ,
\blk00000001/sig0000050d , \blk00000001/sig0000050c , \blk00000001/sig0000050b }),
    .M({\NLW_blk00000001/blk000001d8_M<35>_UNCONNECTED , \NLW_blk00000001/blk000001d8_M<34>_UNCONNECTED ,
\NLW_blk00000001/blk000001d8_M<33>_UNCONNECTED , \NLW_blk00000001/blk000001d8_M<32>_UNCONNECTED , \NLW_blk00000001/blk000001d8_M<31>_UNCONNECTED ,
\NLW_blk00000001/blk000001d8_M<30>_UNCONNECTED , \NLW_blk00000001/blk000001d8_M<29>_UNCONNECTED , \NLW_blk00000001/blk000001d8_M<28>_UNCONNECTED ,
\NLW_blk00000001/blk000001d8_M<27>_UNCONNECTED , \NLW_blk00000001/blk000001d8_M<26>_UNCONNECTED , \NLW_blk00000001/blk000001d8_M<25>_UNCONNECTED ,
\NLW_blk00000001/blk000001d8_M<24>_UNCONNECTED , \NLW_blk00000001/blk000001d8_M<23>_UNCONNECTED , \NLW_blk00000001/blk000001d8_M<22>_UNCONNECTED ,
\NLW_blk00000001/blk000001d8_M<21>_UNCONNECTED , \NLW_blk00000001/blk000001d8_M<20>_UNCONNECTED , \NLW_blk00000001/blk000001d8_M<19>_UNCONNECTED ,
\NLW_blk00000001/blk000001d8_M<18>_UNCONNECTED , \NLW_blk00000001/blk000001d8_M<17>_UNCONNECTED , \NLW_blk00000001/blk000001d8_M<16>_UNCONNECTED ,
\NLW_blk00000001/blk000001d8_M<15>_UNCONNECTED , \NLW_blk00000001/blk000001d8_M<14>_UNCONNECTED , \NLW_blk00000001/blk000001d8_M<13>_UNCONNECTED ,
\NLW_blk00000001/blk000001d8_M<12>_UNCONNECTED , \NLW_blk00000001/blk000001d8_M<11>_UNCONNECTED , \NLW_blk00000001/blk000001d8_M<10>_UNCONNECTED ,
\NLW_blk00000001/blk000001d8_M<9>_UNCONNECTED , \NLW_blk00000001/blk000001d8_M<8>_UNCONNECTED , \NLW_blk00000001/blk000001d8_M<7>_UNCONNECTED ,
\NLW_blk00000001/blk000001d8_M<6>_UNCONNECTED , \NLW_blk00000001/blk000001d8_M<5>_UNCONNECTED , \NLW_blk00000001/blk000001d8_M<4>_UNCONNECTED ,
\NLW_blk00000001/blk000001d8_M<3>_UNCONNECTED , \NLW_blk00000001/blk000001d8_M<2>_UNCONNECTED , \NLW_blk00000001/blk000001d8_M<1>_UNCONNECTED ,
\NLW_blk00000001/blk000001d8_M<0>_UNCONNECTED })
  );
  DSP48A1 #(
    .A0REG ( 0 ),
    .A1REG ( 1 ),
    .B0REG ( 0 ),
    .B1REG ( 1 ),
    .CARRYINREG ( 0 ),
    .CARRYINSEL ( "OPMODE5" ),
    .CREG ( 1 ),
    .DREG ( 1 ),
    .MREG ( 0 ),
    .OPMODEREG ( 1 ),
    .PREG ( 1 ),
    .RSTTYPE ( "SYNC" ),
    .CARRYOUTREG ( 0 ))
  \blk00000001/blk000001d7  (
    .CECARRYIN(\blk00000001/sig0000051d ),
    .RSTC(\blk00000001/sig0000051d ),
    .RSTCARRYIN(\blk00000001/sig0000051d ),
    .CED(\blk00000001/sig0000003a ),
    .RSTD(\blk00000001/sig0000051d ),
    .CEOPMODE(\blk00000001/sig0000003a ),
    .CEC(\blk00000001/sig0000003a ),
    .CARRYOUTF(\NLW_blk00000001/blk000001d7_CARRYOUTF_UNCONNECTED ),
    .RSTOPMODE(\blk00000001/sig0000051d ),
    .RSTM(\blk00000001/sig0000051d ),
    .CLK(aclk),
    .RSTB(\blk00000001/sig0000051d ),
    .CEM(\blk00000001/sig0000051d ),
    .CEB(\blk00000001/sig0000003a ),
    .CARRYIN(\blk00000001/sig0000051d ),
    .CEP(\blk00000001/sig0000003a ),
    .CEA(\blk00000001/sig0000003a ),
    .CARRYOUT(\NLW_blk00000001/blk000001d7_CARRYOUT_UNCONNECTED ),
    .RSTA(\blk00000001/sig0000051d ),
    .RSTP(\blk00000001/sig0000051d ),
    .B({\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000052f , \blk00000001/sig0000052e ,
\blk00000001/sig0000052d , \blk00000001/sig0000052c , \blk00000001/sig0000052b , \blk00000001/sig0000052a , \blk00000001/sig00000529 ,
\blk00000001/sig00000528 , \blk00000001/sig00000527 , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d }),
    .BCOUT({\NLW_blk00000001/blk000001d7_BCOUT<17>_UNCONNECTED , \NLW_blk00000001/blk000001d7_BCOUT<16>_UNCONNECTED ,
\NLW_blk00000001/blk000001d7_BCOUT<15>_UNCONNECTED , \NLW_blk00000001/blk000001d7_BCOUT<14>_UNCONNECTED ,
\NLW_blk00000001/blk000001d7_BCOUT<13>_UNCONNECTED , \NLW_blk00000001/blk000001d7_BCOUT<12>_UNCONNECTED ,
\NLW_blk00000001/blk000001d7_BCOUT<11>_UNCONNECTED , \NLW_blk00000001/blk000001d7_BCOUT<10>_UNCONNECTED ,
\NLW_blk00000001/blk000001d7_BCOUT<9>_UNCONNECTED , \NLW_blk00000001/blk000001d7_BCOUT<8>_UNCONNECTED ,
\NLW_blk00000001/blk000001d7_BCOUT<7>_UNCONNECTED , \NLW_blk00000001/blk000001d7_BCOUT<6>_UNCONNECTED ,
\NLW_blk00000001/blk000001d7_BCOUT<5>_UNCONNECTED , \NLW_blk00000001/blk000001d7_BCOUT<4>_UNCONNECTED ,
\NLW_blk00000001/blk000001d7_BCOUT<3>_UNCONNECTED , \NLW_blk00000001/blk000001d7_BCOUT<2>_UNCONNECTED ,
\NLW_blk00000001/blk000001d7_BCOUT<1>_UNCONNECTED , \NLW_blk00000001/blk000001d7_BCOUT<0>_UNCONNECTED }),
    .PCIN({\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d }),
    .C({\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig000004f6 , \blk00000001/sig000004f5 , \blk00000001/sig000004f4 , \blk00000001/sig000004f3 ,
\blk00000001/sig000004f2 , \blk00000001/sig000004f1 , \blk00000001/sig000004f0 , \blk00000001/sig000004ef , \blk00000001/sig000004ee ,
\blk00000001/sig000004ed , \blk00000001/sig000004ec , \blk00000001/sig000004eb , \blk00000001/sig000004ea , \blk00000001/sig000004e9 ,
\blk00000001/sig000004e8 , \blk00000001/sig000004e7 , \blk00000001/sig000004e6 , \blk00000001/sig000004e5 , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d }),
    .P({\NLW_blk00000001/blk000001d7_P<47>_UNCONNECTED , \NLW_blk00000001/blk000001d7_P<46>_UNCONNECTED ,
\NLW_blk00000001/blk000001d7_P<45>_UNCONNECTED , \NLW_blk00000001/blk000001d7_P<44>_UNCONNECTED , \NLW_blk00000001/blk000001d7_P<43>_UNCONNECTED ,
\NLW_blk00000001/blk000001d7_P<42>_UNCONNECTED , \NLW_blk00000001/blk000001d7_P<41>_UNCONNECTED , \NLW_blk00000001/blk000001d7_P<40>_UNCONNECTED ,
\NLW_blk00000001/blk000001d7_P<39>_UNCONNECTED , \NLW_blk00000001/blk000001d7_P<38>_UNCONNECTED , \NLW_blk00000001/blk000001d7_P<37>_UNCONNECTED ,
\NLW_blk00000001/blk000001d7_P<36>_UNCONNECTED , \NLW_blk00000001/blk000001d7_P<35>_UNCONNECTED , \NLW_blk00000001/blk000001d7_P<34>_UNCONNECTED ,
\NLW_blk00000001/blk000001d7_P<33>_UNCONNECTED , \NLW_blk00000001/blk000001d7_P<32>_UNCONNECTED , \NLW_blk00000001/blk000001d7_P<31>_UNCONNECTED ,
\NLW_blk00000001/blk000001d7_P<30>_UNCONNECTED , \NLW_blk00000001/blk000001d7_P<29>_UNCONNECTED , \NLW_blk00000001/blk000001d7_P<28>_UNCONNECTED ,
\NLW_blk00000001/blk000001d7_P<27>_UNCONNECTED , \NLW_blk00000001/blk000001d7_P<26>_UNCONNECTED , \NLW_blk00000001/blk000001d7_P<25>_UNCONNECTED ,
\NLW_blk00000001/blk000001d7_P<24>_UNCONNECTED , \NLW_blk00000001/blk000001d7_P<23>_UNCONNECTED , \NLW_blk00000001/blk000001d7_P<22>_UNCONNECTED ,
\NLW_blk00000001/blk000001d7_P<21>_UNCONNECTED , \NLW_blk00000001/blk000001d7_P<20>_UNCONNECTED , \NLW_blk00000001/blk000001d7_P<19>_UNCONNECTED ,
\NLW_blk00000001/blk000001d7_P<18>_UNCONNECTED , \NLW_blk00000001/blk000001d7_P<17>_UNCONNECTED , \NLW_blk00000001/blk000001d7_P<16>_UNCONNECTED ,
\NLW_blk00000001/blk000001d7_P<15>_UNCONNECTED , \NLW_blk00000001/blk000001d7_P<14>_UNCONNECTED , \NLW_blk00000001/blk000001d7_P<13>_UNCONNECTED ,
\NLW_blk00000001/blk000001d7_P<12>_UNCONNECTED , \NLW_blk00000001/blk000001d7_P<11>_UNCONNECTED , \NLW_blk00000001/blk000001d7_P<10>_UNCONNECTED ,
\NLW_blk00000001/blk000001d7_P<9>_UNCONNECTED , \NLW_blk00000001/blk000001d7_P<8>_UNCONNECTED , \NLW_blk00000001/blk000001d7_P<7>_UNCONNECTED ,
\NLW_blk00000001/blk000001d7_P<6>_UNCONNECTED , \NLW_blk00000001/blk000001d7_P<5>_UNCONNECTED , \NLW_blk00000001/blk000001d7_P<4>_UNCONNECTED ,
\NLW_blk00000001/blk000001d7_P<3>_UNCONNECTED , \NLW_blk00000001/blk000001d7_P<2>_UNCONNECTED , \NLW_blk00000001/blk000001d7_P<1>_UNCONNECTED ,
\NLW_blk00000001/blk000001d7_P<0>_UNCONNECTED }),
    .OPMODE({\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000003a ,
\blk00000001/sig0000003a , \blk00000001/sig0000003a , \blk00000001/sig0000003a }),
    .D({\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d }),
    .PCOUT({\blk00000001/sig000004e3 , \blk00000001/sig000004e2 , \blk00000001/sig000004e1 , \blk00000001/sig000004e0 , \blk00000001/sig000004df ,
\blk00000001/sig000004de , \blk00000001/sig000004dd , \blk00000001/sig000004dc , \blk00000001/sig000004db , \blk00000001/sig000004da ,
\blk00000001/sig000004d9 , \blk00000001/sig000004d8 , \blk00000001/sig000004d7 , \blk00000001/sig000004d6 , \blk00000001/sig000004d5 ,
\blk00000001/sig000004d4 , \blk00000001/sig000004d3 , \blk00000001/sig000004d2 , \blk00000001/sig000004d1 , \blk00000001/sig000004d0 ,
\blk00000001/sig000004cf , \blk00000001/sig000004ce , \blk00000001/sig000004cd , \blk00000001/sig000004cc , \blk00000001/sig000004cb ,
\blk00000001/sig000004ca , \blk00000001/sig000004c9 , \blk00000001/sig000004c8 , \blk00000001/sig000004c7 , \blk00000001/sig000004c6 ,
\blk00000001/sig000004c5 , \blk00000001/sig000004c4 , \blk00000001/sig000004c3 , \blk00000001/sig000004c2 , \blk00000001/sig000004c1 ,
\blk00000001/sig000004c0 , \blk00000001/sig000004bf , \blk00000001/sig000004be , \blk00000001/sig000004bd , \blk00000001/sig000004bc ,
\blk00000001/sig000004bb , \blk00000001/sig000004ba , \blk00000001/sig000004b9 , \blk00000001/sig000004b8 , \blk00000001/sig000004b7 ,
\blk00000001/sig000004b6 , \blk00000001/sig000004b5 , \blk00000001/sig000004b4 }),
    .A({\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d }),
    .M({\NLW_blk00000001/blk000001d7_M<35>_UNCONNECTED , \NLW_blk00000001/blk000001d7_M<34>_UNCONNECTED ,
\NLW_blk00000001/blk000001d7_M<33>_UNCONNECTED , \NLW_blk00000001/blk000001d7_M<32>_UNCONNECTED , \NLW_blk00000001/blk000001d7_M<31>_UNCONNECTED ,
\NLW_blk00000001/blk000001d7_M<30>_UNCONNECTED , \NLW_blk00000001/blk000001d7_M<29>_UNCONNECTED , \NLW_blk00000001/blk000001d7_M<28>_UNCONNECTED ,
\NLW_blk00000001/blk000001d7_M<27>_UNCONNECTED , \NLW_blk00000001/blk000001d7_M<26>_UNCONNECTED , \NLW_blk00000001/blk000001d7_M<25>_UNCONNECTED ,
\NLW_blk00000001/blk000001d7_M<24>_UNCONNECTED , \NLW_blk00000001/blk000001d7_M<23>_UNCONNECTED , \NLW_blk00000001/blk000001d7_M<22>_UNCONNECTED ,
\NLW_blk00000001/blk000001d7_M<21>_UNCONNECTED , \NLW_blk00000001/blk000001d7_M<20>_UNCONNECTED , \NLW_blk00000001/blk000001d7_M<19>_UNCONNECTED ,
\NLW_blk00000001/blk000001d7_M<18>_UNCONNECTED , \NLW_blk00000001/blk000001d7_M<17>_UNCONNECTED , \NLW_blk00000001/blk000001d7_M<16>_UNCONNECTED ,
\NLW_blk00000001/blk000001d7_M<15>_UNCONNECTED , \NLW_blk00000001/blk000001d7_M<14>_UNCONNECTED , \NLW_blk00000001/blk000001d7_M<13>_UNCONNECTED ,
\NLW_blk00000001/blk000001d7_M<12>_UNCONNECTED , \NLW_blk00000001/blk000001d7_M<11>_UNCONNECTED , \NLW_blk00000001/blk000001d7_M<10>_UNCONNECTED ,
\NLW_blk00000001/blk000001d7_M<9>_UNCONNECTED , \NLW_blk00000001/blk000001d7_M<8>_UNCONNECTED , \NLW_blk00000001/blk000001d7_M<7>_UNCONNECTED ,
\NLW_blk00000001/blk000001d7_M<6>_UNCONNECTED , \NLW_blk00000001/blk000001d7_M<5>_UNCONNECTED , \NLW_blk00000001/blk000001d7_M<4>_UNCONNECTED ,
\NLW_blk00000001/blk000001d7_M<3>_UNCONNECTED , \NLW_blk00000001/blk000001d7_M<2>_UNCONNECTED , \NLW_blk00000001/blk000001d7_M<1>_UNCONNECTED ,
\NLW_blk00000001/blk000001d7_M<0>_UNCONNECTED })
  );
  DSP48A1 #(
    .A0REG ( 0 ),
    .A1REG ( 1 ),
    .B0REG ( 0 ),
    .B1REG ( 1 ),
    .CARRYINREG ( 0 ),
    .CARRYINSEL ( "OPMODE5" ),
    .CREG ( 1 ),
    .DREG ( 1 ),
    .MREG ( 0 ),
    .OPMODEREG ( 1 ),
    .PREG ( 1 ),
    .RSTTYPE ( "SYNC" ),
    .CARRYOUTREG ( 0 ))
  \blk00000001/blk000001d6  (
    .CECARRYIN(\blk00000001/sig0000051d ),
    .RSTC(\blk00000001/sig0000051d ),
    .RSTCARRYIN(\blk00000001/sig0000051d ),
    .CED(\blk00000001/sig0000003a ),
    .RSTD(\blk00000001/sig0000051d ),
    .CEOPMODE(\blk00000001/sig0000003a ),
    .CEC(\blk00000001/sig0000003a ),
    .CARRYOUTF(\NLW_blk00000001/blk000001d6_CARRYOUTF_UNCONNECTED ),
    .RSTOPMODE(\blk00000001/sig0000051d ),
    .RSTM(\blk00000001/sig0000051d ),
    .CLK(aclk),
    .RSTB(\blk00000001/sig0000051d ),
    .CEM(\blk00000001/sig0000051d ),
    .CEB(\blk00000001/sig0000003a ),
    .CARRYIN(\blk00000001/sig0000051d ),
    .CEP(\blk00000001/sig0000003a ),
    .CEA(\blk00000001/sig0000003a ),
    .CARRYOUT(\NLW_blk00000001/blk000001d6_CARRYOUT_UNCONNECTED ),
    .RSTA(\blk00000001/sig0000051d ),
    .RSTP(\blk00000001/sig0000051d ),
    .B({\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d }),
    .BCOUT({\NLW_blk00000001/blk000001d6_BCOUT<17>_UNCONNECTED , \NLW_blk00000001/blk000001d6_BCOUT<16>_UNCONNECTED ,
\NLW_blk00000001/blk000001d6_BCOUT<15>_UNCONNECTED , \NLW_blk00000001/blk000001d6_BCOUT<14>_UNCONNECTED ,
\NLW_blk00000001/blk000001d6_BCOUT<13>_UNCONNECTED , \NLW_blk00000001/blk000001d6_BCOUT<12>_UNCONNECTED ,
\NLW_blk00000001/blk000001d6_BCOUT<11>_UNCONNECTED , \NLW_blk00000001/blk000001d6_BCOUT<10>_UNCONNECTED ,
\NLW_blk00000001/blk000001d6_BCOUT<9>_UNCONNECTED , \NLW_blk00000001/blk000001d6_BCOUT<8>_UNCONNECTED ,
\NLW_blk00000001/blk000001d6_BCOUT<7>_UNCONNECTED , \NLW_blk00000001/blk000001d6_BCOUT<6>_UNCONNECTED ,
\NLW_blk00000001/blk000001d6_BCOUT<5>_UNCONNECTED , \NLW_blk00000001/blk000001d6_BCOUT<4>_UNCONNECTED ,
\NLW_blk00000001/blk000001d6_BCOUT<3>_UNCONNECTED , \NLW_blk00000001/blk000001d6_BCOUT<2>_UNCONNECTED ,
\NLW_blk00000001/blk000001d6_BCOUT<1>_UNCONNECTED , \NLW_blk00000001/blk000001d6_BCOUT<0>_UNCONNECTED }),
    .PCIN({\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d }),
    .C({\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000044d , \blk00000001/sig0000044c , \blk00000001/sig0000044b , \blk00000001/sig0000044a , \blk00000001/sig00000449 ,
\blk00000001/sig00000448 , \blk00000001/sig00000447 , \blk00000001/sig00000446 , \blk00000001/sig00000445 , \blk00000001/sig00000444 ,
\blk00000001/sig00000443 , \blk00000001/sig00000442 , \blk00000001/sig00000441 , \blk00000001/sig00000440 , \blk00000001/sig0000043f ,
\blk00000001/sig0000043e , \blk00000001/sig0000043d , \blk00000001/sig0000043c , \blk00000001/sig0000043b , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d }),
    .P({\NLW_blk00000001/blk000001d6_P<47>_UNCONNECTED , \NLW_blk00000001/blk000001d6_P<46>_UNCONNECTED ,
\NLW_blk00000001/blk000001d6_P<45>_UNCONNECTED , \NLW_blk00000001/blk000001d6_P<44>_UNCONNECTED , \NLW_blk00000001/blk000001d6_P<43>_UNCONNECTED ,
\NLW_blk00000001/blk000001d6_P<42>_UNCONNECTED , \NLW_blk00000001/blk000001d6_P<41>_UNCONNECTED , \NLW_blk00000001/blk000001d6_P<40>_UNCONNECTED ,
\NLW_blk00000001/blk000001d6_P<39>_UNCONNECTED , \NLW_blk00000001/blk000001d6_P<38>_UNCONNECTED , \NLW_blk00000001/blk000001d6_P<37>_UNCONNECTED ,
\NLW_blk00000001/blk000001d6_P<36>_UNCONNECTED , \NLW_blk00000001/blk000001d6_P<35>_UNCONNECTED , \NLW_blk00000001/blk000001d6_P<34>_UNCONNECTED ,
\NLW_blk00000001/blk000001d6_P<33>_UNCONNECTED , \NLW_blk00000001/blk000001d6_P<32>_UNCONNECTED , \NLW_blk00000001/blk000001d6_P<31>_UNCONNECTED ,
\NLW_blk00000001/blk000001d6_P<30>_UNCONNECTED , \NLW_blk00000001/blk000001d6_P<29>_UNCONNECTED , \NLW_blk00000001/blk000001d6_P<28>_UNCONNECTED ,
\NLW_blk00000001/blk000001d6_P<27>_UNCONNECTED , \NLW_blk00000001/blk000001d6_P<26>_UNCONNECTED , \NLW_blk00000001/blk000001d6_P<25>_UNCONNECTED ,
\NLW_blk00000001/blk000001d6_P<24>_UNCONNECTED , \NLW_blk00000001/blk000001d6_P<23>_UNCONNECTED , \NLW_blk00000001/blk000001d6_P<22>_UNCONNECTED ,
\NLW_blk00000001/blk000001d6_P<21>_UNCONNECTED , \NLW_blk00000001/blk000001d6_P<20>_UNCONNECTED , \NLW_blk00000001/blk000001d6_P<19>_UNCONNECTED ,
\NLW_blk00000001/blk000001d6_P<18>_UNCONNECTED , \NLW_blk00000001/blk000001d6_P<17>_UNCONNECTED , \NLW_blk00000001/blk000001d6_P<16>_UNCONNECTED ,
\NLW_blk00000001/blk000001d6_P<15>_UNCONNECTED , \NLW_blk00000001/blk000001d6_P<14>_UNCONNECTED , \NLW_blk00000001/blk000001d6_P<13>_UNCONNECTED ,
\NLW_blk00000001/blk000001d6_P<12>_UNCONNECTED , \NLW_blk00000001/blk000001d6_P<11>_UNCONNECTED , \NLW_blk00000001/blk000001d6_P<10>_UNCONNECTED ,
\NLW_blk00000001/blk000001d6_P<9>_UNCONNECTED , \NLW_blk00000001/blk000001d6_P<8>_UNCONNECTED , \NLW_blk00000001/blk000001d6_P<7>_UNCONNECTED ,
\NLW_blk00000001/blk000001d6_P<6>_UNCONNECTED , \NLW_blk00000001/blk000001d6_P<5>_UNCONNECTED , \NLW_blk00000001/blk000001d6_P<4>_UNCONNECTED ,
\NLW_blk00000001/blk000001d6_P<3>_UNCONNECTED , \NLW_blk00000001/blk000001d6_P<2>_UNCONNECTED , \NLW_blk00000001/blk000001d6_P<1>_UNCONNECTED ,
\NLW_blk00000001/blk000001d6_P<0>_UNCONNECTED }),
    .OPMODE({\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000003a ,
\blk00000001/sig0000003a , \blk00000001/sig0000003a , \blk00000001/sig0000003a }),
    .D({\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d }),
    .PCOUT({\blk00000001/sig0000043a , \blk00000001/sig00000439 , \blk00000001/sig00000438 , \blk00000001/sig00000437 , \blk00000001/sig00000436 ,
\blk00000001/sig00000435 , \blk00000001/sig00000434 , \blk00000001/sig00000433 , \blk00000001/sig00000432 , \blk00000001/sig00000431 ,
\blk00000001/sig00000430 , \blk00000001/sig0000042f , \blk00000001/sig0000042e , \blk00000001/sig0000042d , \blk00000001/sig0000042c ,
\blk00000001/sig0000042b , \blk00000001/sig0000042a , \blk00000001/sig00000429 , \blk00000001/sig00000428 , \blk00000001/sig00000427 ,
\blk00000001/sig00000426 , \blk00000001/sig00000425 , \blk00000001/sig00000424 , \blk00000001/sig00000423 , \blk00000001/sig00000422 ,
\blk00000001/sig00000421 , \blk00000001/sig00000420 , \blk00000001/sig0000041f , \blk00000001/sig0000041e , \blk00000001/sig0000041d ,
\blk00000001/sig0000041c , \blk00000001/sig0000041b , \blk00000001/sig0000041a , \blk00000001/sig00000419 , \blk00000001/sig00000418 ,
\blk00000001/sig00000417 , \blk00000001/sig00000416 , \blk00000001/sig00000415 , \blk00000001/sig00000414 , \blk00000001/sig00000413 ,
\blk00000001/sig00000412 , \blk00000001/sig00000411 , \blk00000001/sig00000410 , \blk00000001/sig0000040f , \blk00000001/sig0000040e ,
\blk00000001/sig0000040d , \blk00000001/sig0000040c , \blk00000001/sig0000040b }),
    .A({\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d }),
    .M({\NLW_blk00000001/blk000001d6_M<35>_UNCONNECTED , \NLW_blk00000001/blk000001d6_M<34>_UNCONNECTED ,
\NLW_blk00000001/blk000001d6_M<33>_UNCONNECTED , \NLW_blk00000001/blk000001d6_M<32>_UNCONNECTED , \NLW_blk00000001/blk000001d6_M<31>_UNCONNECTED ,
\NLW_blk00000001/blk000001d6_M<30>_UNCONNECTED , \NLW_blk00000001/blk000001d6_M<29>_UNCONNECTED , \NLW_blk00000001/blk000001d6_M<28>_UNCONNECTED ,
\NLW_blk00000001/blk000001d6_M<27>_UNCONNECTED , \NLW_blk00000001/blk000001d6_M<26>_UNCONNECTED , \NLW_blk00000001/blk000001d6_M<25>_UNCONNECTED ,
\NLW_blk00000001/blk000001d6_M<24>_UNCONNECTED , \NLW_blk00000001/blk000001d6_M<23>_UNCONNECTED , \NLW_blk00000001/blk000001d6_M<22>_UNCONNECTED ,
\NLW_blk00000001/blk000001d6_M<21>_UNCONNECTED , \NLW_blk00000001/blk000001d6_M<20>_UNCONNECTED , \NLW_blk00000001/blk000001d6_M<19>_UNCONNECTED ,
\NLW_blk00000001/blk000001d6_M<18>_UNCONNECTED , \NLW_blk00000001/blk000001d6_M<17>_UNCONNECTED , \NLW_blk00000001/blk000001d6_M<16>_UNCONNECTED ,
\NLW_blk00000001/blk000001d6_M<15>_UNCONNECTED , \NLW_blk00000001/blk000001d6_M<14>_UNCONNECTED , \NLW_blk00000001/blk000001d6_M<13>_UNCONNECTED ,
\NLW_blk00000001/blk000001d6_M<12>_UNCONNECTED , \NLW_blk00000001/blk000001d6_M<11>_UNCONNECTED , \NLW_blk00000001/blk000001d6_M<10>_UNCONNECTED ,
\NLW_blk00000001/blk000001d6_M<9>_UNCONNECTED , \NLW_blk00000001/blk000001d6_M<8>_UNCONNECTED , \NLW_blk00000001/blk000001d6_M<7>_UNCONNECTED ,
\NLW_blk00000001/blk000001d6_M<6>_UNCONNECTED , \NLW_blk00000001/blk000001d6_M<5>_UNCONNECTED , \NLW_blk00000001/blk000001d6_M<4>_UNCONNECTED ,
\NLW_blk00000001/blk000001d6_M<3>_UNCONNECTED , \NLW_blk00000001/blk000001d6_M<2>_UNCONNECTED , \NLW_blk00000001/blk000001d6_M<1>_UNCONNECTED ,
\NLW_blk00000001/blk000001d6_M<0>_UNCONNECTED })
  );
  DSP48A1 #(
    .A0REG ( 0 ),
    .A1REG ( 1 ),
    .B0REG ( 0 ),
    .B1REG ( 1 ),
    .CARRYINREG ( 0 ),
    .CARRYINSEL ( "OPMODE5" ),
    .CREG ( 1 ),
    .DREG ( 1 ),
    .MREG ( 0 ),
    .OPMODEREG ( 1 ),
    .PREG ( 1 ),
    .RSTTYPE ( "SYNC" ),
    .CARRYOUTREG ( 0 ))
  \blk00000001/blk000001d5  (
    .CECARRYIN(\blk00000001/sig0000051d ),
    .RSTC(\blk00000001/sig0000051d ),
    .RSTCARRYIN(\blk00000001/sig0000051d ),
    .CED(\blk00000001/sig0000003a ),
    .RSTD(\blk00000001/sig0000051d ),
    .CEOPMODE(\blk00000001/sig0000003a ),
    .CEC(\blk00000001/sig0000003a ),
    .CARRYOUTF(\NLW_blk00000001/blk000001d5_CARRYOUTF_UNCONNECTED ),
    .RSTOPMODE(\blk00000001/sig0000051d ),
    .RSTM(\blk00000001/sig0000051d ),
    .CLK(aclk),
    .RSTB(\blk00000001/sig0000051d ),
    .CEM(\blk00000001/sig0000051d ),
    .CEB(\blk00000001/sig0000003a ),
    .CARRYIN(\blk00000001/sig0000051d ),
    .CEP(\blk00000001/sig0000003a ),
    .CEA(\blk00000001/sig0000003a ),
    .CARRYOUT(\NLW_blk00000001/blk000001d5_CARRYOUT_UNCONNECTED ),
    .RSTA(\blk00000001/sig0000051d ),
    .RSTP(\blk00000001/sig0000051d ),
    .B({\blk00000001/sig000003a8 , \blk00000001/sig000003a7 , \blk00000001/sig000003a6 , \blk00000001/sig000003a5 , \blk00000001/sig000003a4 ,
\blk00000001/sig000003a3 , \blk00000001/sig000003a2 , \blk00000001/sig000003a1 , \blk00000001/sig000003a0 , \blk00000001/sig0000039f ,
\blk00000001/sig0000039e , \blk00000001/sig0000039d , \blk00000001/sig0000039c , \blk00000001/sig0000039b , \blk00000001/sig0000039a ,
\blk00000001/sig00000399 , \blk00000001/sig00000398 , \blk00000001/sig00000397 }),
    .BCOUT({\NLW_blk00000001/blk000001d5_BCOUT<17>_UNCONNECTED , \NLW_blk00000001/blk000001d5_BCOUT<16>_UNCONNECTED ,
\NLW_blk00000001/blk000001d5_BCOUT<15>_UNCONNECTED , \NLW_blk00000001/blk000001d5_BCOUT<14>_UNCONNECTED ,
\NLW_blk00000001/blk000001d5_BCOUT<13>_UNCONNECTED , \NLW_blk00000001/blk000001d5_BCOUT<12>_UNCONNECTED ,
\NLW_blk00000001/blk000001d5_BCOUT<11>_UNCONNECTED , \NLW_blk00000001/blk000001d5_BCOUT<10>_UNCONNECTED ,
\NLW_blk00000001/blk000001d5_BCOUT<9>_UNCONNECTED , \NLW_blk00000001/blk000001d5_BCOUT<8>_UNCONNECTED ,
\NLW_blk00000001/blk000001d5_BCOUT<7>_UNCONNECTED , \NLW_blk00000001/blk000001d5_BCOUT<6>_UNCONNECTED ,
\NLW_blk00000001/blk000001d5_BCOUT<5>_UNCONNECTED , \NLW_blk00000001/blk000001d5_BCOUT<4>_UNCONNECTED ,
\NLW_blk00000001/blk000001d5_BCOUT<3>_UNCONNECTED , \NLW_blk00000001/blk000001d5_BCOUT<2>_UNCONNECTED ,
\NLW_blk00000001/blk000001d5_BCOUT<1>_UNCONNECTED , \NLW_blk00000001/blk000001d5_BCOUT<0>_UNCONNECTED }),
    .PCIN({\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d }),
    .C({\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig00000396 , \blk00000001/sig00000395 , \blk00000001/sig00000394 , \blk00000001/sig00000393 , \blk00000001/sig00000392 ,
\blk00000001/sig00000391 , \blk00000001/sig00000390 , \blk00000001/sig0000038f , \blk00000001/sig0000038e , \blk00000001/sig0000038d ,
\blk00000001/sig0000038c , \blk00000001/sig0000038b , \blk00000001/sig0000038a , \blk00000001/sig00000389 , \blk00000001/sig00000388 ,
\blk00000001/sig00000387 , \blk00000001/sig00000386 , \blk00000001/sig00000385 , \blk00000001/sig00000384 , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d }),
    .P({\NLW_blk00000001/blk000001d5_P<47>_UNCONNECTED , \NLW_blk00000001/blk000001d5_P<46>_UNCONNECTED ,
\NLW_blk00000001/blk000001d5_P<45>_UNCONNECTED , \NLW_blk00000001/blk000001d5_P<44>_UNCONNECTED , \NLW_blk00000001/blk000001d5_P<43>_UNCONNECTED ,
\NLW_blk00000001/blk000001d5_P<42>_UNCONNECTED , \NLW_blk00000001/blk000001d5_P<41>_UNCONNECTED , \NLW_blk00000001/blk000001d5_P<40>_UNCONNECTED ,
\NLW_blk00000001/blk000001d5_P<39>_UNCONNECTED , \NLW_blk00000001/blk000001d5_P<38>_UNCONNECTED , \NLW_blk00000001/blk000001d5_P<37>_UNCONNECTED ,
\NLW_blk00000001/blk000001d5_P<36>_UNCONNECTED , \NLW_blk00000001/blk000001d5_P<35>_UNCONNECTED , \NLW_blk00000001/blk000001d5_P<34>_UNCONNECTED ,
\NLW_blk00000001/blk000001d5_P<33>_UNCONNECTED , \NLW_blk00000001/blk000001d5_P<32>_UNCONNECTED , \NLW_blk00000001/blk000001d5_P<31>_UNCONNECTED ,
\NLW_blk00000001/blk000001d5_P<30>_UNCONNECTED , \NLW_blk00000001/blk000001d5_P<29>_UNCONNECTED , \NLW_blk00000001/blk000001d5_P<28>_UNCONNECTED ,
\NLW_blk00000001/blk000001d5_P<27>_UNCONNECTED , \NLW_blk00000001/blk000001d5_P<26>_UNCONNECTED , \NLW_blk00000001/blk000001d5_P<25>_UNCONNECTED ,
\NLW_blk00000001/blk000001d5_P<24>_UNCONNECTED , \NLW_blk00000001/blk000001d5_P<23>_UNCONNECTED , \NLW_blk00000001/blk000001d5_P<22>_UNCONNECTED ,
\NLW_blk00000001/blk000001d5_P<21>_UNCONNECTED , \NLW_blk00000001/blk000001d5_P<20>_UNCONNECTED , \NLW_blk00000001/blk000001d5_P<19>_UNCONNECTED ,
\NLW_blk00000001/blk000001d5_P<18>_UNCONNECTED , \NLW_blk00000001/blk000001d5_P<17>_UNCONNECTED , \NLW_blk00000001/blk000001d5_P<16>_UNCONNECTED ,
\NLW_blk00000001/blk000001d5_P<15>_UNCONNECTED , \NLW_blk00000001/blk000001d5_P<14>_UNCONNECTED , \NLW_blk00000001/blk000001d5_P<13>_UNCONNECTED ,
\NLW_blk00000001/blk000001d5_P<12>_UNCONNECTED , \NLW_blk00000001/blk000001d5_P<11>_UNCONNECTED , \NLW_blk00000001/blk000001d5_P<10>_UNCONNECTED ,
\NLW_blk00000001/blk000001d5_P<9>_UNCONNECTED , \NLW_blk00000001/blk000001d5_P<8>_UNCONNECTED , \NLW_blk00000001/blk000001d5_P<7>_UNCONNECTED ,
\NLW_blk00000001/blk000001d5_P<6>_UNCONNECTED , \NLW_blk00000001/blk000001d5_P<5>_UNCONNECTED , \NLW_blk00000001/blk000001d5_P<4>_UNCONNECTED ,
\NLW_blk00000001/blk000001d5_P<3>_UNCONNECTED , \NLW_blk00000001/blk000001d5_P<2>_UNCONNECTED , \NLW_blk00000001/blk000001d5_P<1>_UNCONNECTED ,
\NLW_blk00000001/blk000001d5_P<0>_UNCONNECTED }),
    .OPMODE({\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000003a ,
\blk00000001/sig0000003a , \blk00000001/sig0000003a , \blk00000001/sig0000003a }),
    .D({\blk00000001/sig000003c6 , \blk00000001/sig000003c6 , \blk00000001/sig000003c6 , \blk00000001/sig000003c6 , \blk00000001/sig000003c6 ,
\blk00000001/sig000003c6 , \blk00000001/sig000003c6 , \blk00000001/sig000003c5 , \blk00000001/sig000003c4 , \blk00000001/sig000003c3 ,
\blk00000001/sig000003c2 , \blk00000001/sig000003c1 , \blk00000001/sig000003c0 , \blk00000001/sig000003bf , \blk00000001/sig000003be ,
\blk00000001/sig000003bd , \blk00000001/sig000003bc , \blk00000001/sig000003bb }),
    .PCOUT({\blk00000001/sig00000383 , \blk00000001/sig00000382 , \blk00000001/sig00000381 , \blk00000001/sig00000380 , \blk00000001/sig0000037f ,
\blk00000001/sig0000037e , \blk00000001/sig0000037d , \blk00000001/sig0000037c , \blk00000001/sig0000037b , \blk00000001/sig0000037a ,
\blk00000001/sig00000379 , \blk00000001/sig00000378 , \blk00000001/sig00000377 , \blk00000001/sig00000376 , \blk00000001/sig00000375 ,
\blk00000001/sig00000374 , \blk00000001/sig00000373 , \blk00000001/sig00000372 , \blk00000001/sig00000371 , \blk00000001/sig00000370 ,
\blk00000001/sig0000036f , \blk00000001/sig0000036e , \blk00000001/sig0000036d , \blk00000001/sig0000036c , \blk00000001/sig0000036b ,
\blk00000001/sig0000036a , \blk00000001/sig00000369 , \blk00000001/sig00000368 , \blk00000001/sig00000367 , \blk00000001/sig00000366 ,
\blk00000001/sig00000365 , \blk00000001/sig00000364 , \blk00000001/sig00000363 , \blk00000001/sig00000362 , \blk00000001/sig00000361 ,
\blk00000001/sig00000360 , \blk00000001/sig0000035f , \blk00000001/sig0000035e , \blk00000001/sig0000035d , \blk00000001/sig0000035c ,
\blk00000001/sig0000035b , \blk00000001/sig0000035a , \blk00000001/sig00000359 , \blk00000001/sig00000358 , \blk00000001/sig00000357 ,
\blk00000001/sig00000356 , \blk00000001/sig00000355 , \blk00000001/sig00000354 }),
    .A({\blk00000001/sig000003ba , \blk00000001/sig000003b9 , \blk00000001/sig000003b8 , \blk00000001/sig000003b7 , \blk00000001/sig000003b6 ,
\blk00000001/sig000003b5 , \blk00000001/sig000003b4 , \blk00000001/sig000003b3 , \blk00000001/sig000003b2 , \blk00000001/sig000003b1 ,
\blk00000001/sig000003b0 , \blk00000001/sig000003af , \blk00000001/sig000003ae , \blk00000001/sig000003ad , \blk00000001/sig000003ac ,
\blk00000001/sig000003ab , \blk00000001/sig000003aa , \blk00000001/sig000003a9 }),
    .M({\NLW_blk00000001/blk000001d5_M<35>_UNCONNECTED , \NLW_blk00000001/blk000001d5_M<34>_UNCONNECTED ,
\NLW_blk00000001/blk000001d5_M<33>_UNCONNECTED , \NLW_blk00000001/blk000001d5_M<32>_UNCONNECTED , \NLW_blk00000001/blk000001d5_M<31>_UNCONNECTED ,
\NLW_blk00000001/blk000001d5_M<30>_UNCONNECTED , \NLW_blk00000001/blk000001d5_M<29>_UNCONNECTED , \NLW_blk00000001/blk000001d5_M<28>_UNCONNECTED ,
\NLW_blk00000001/blk000001d5_M<27>_UNCONNECTED , \NLW_blk00000001/blk000001d5_M<26>_UNCONNECTED , \NLW_blk00000001/blk000001d5_M<25>_UNCONNECTED ,
\NLW_blk00000001/blk000001d5_M<24>_UNCONNECTED , \NLW_blk00000001/blk000001d5_M<23>_UNCONNECTED , \NLW_blk00000001/blk000001d5_M<22>_UNCONNECTED ,
\NLW_blk00000001/blk000001d5_M<21>_UNCONNECTED , \NLW_blk00000001/blk000001d5_M<20>_UNCONNECTED , \NLW_blk00000001/blk000001d5_M<19>_UNCONNECTED ,
\NLW_blk00000001/blk000001d5_M<18>_UNCONNECTED , \NLW_blk00000001/blk000001d5_M<17>_UNCONNECTED , \NLW_blk00000001/blk000001d5_M<16>_UNCONNECTED ,
\NLW_blk00000001/blk000001d5_M<15>_UNCONNECTED , \NLW_blk00000001/blk000001d5_M<14>_UNCONNECTED , \NLW_blk00000001/blk000001d5_M<13>_UNCONNECTED ,
\NLW_blk00000001/blk000001d5_M<12>_UNCONNECTED , \NLW_blk00000001/blk000001d5_M<11>_UNCONNECTED , \NLW_blk00000001/blk000001d5_M<10>_UNCONNECTED ,
\NLW_blk00000001/blk000001d5_M<9>_UNCONNECTED , \NLW_blk00000001/blk000001d5_M<8>_UNCONNECTED , \NLW_blk00000001/blk000001d5_M<7>_UNCONNECTED ,
\NLW_blk00000001/blk000001d5_M<6>_UNCONNECTED , \NLW_blk00000001/blk000001d5_M<5>_UNCONNECTED , \NLW_blk00000001/blk000001d5_M<4>_UNCONNECTED ,
\NLW_blk00000001/blk000001d5_M<3>_UNCONNECTED , \NLW_blk00000001/blk000001d5_M<2>_UNCONNECTED , \NLW_blk00000001/blk000001d5_M<1>_UNCONNECTED ,
\NLW_blk00000001/blk000001d5_M<0>_UNCONNECTED })
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000001d4  (
    .C(aclk),
    .D(\blk00000001/sig0000051c ),
    .Q(\blk00000001/sig000004e4 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000001d3  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig0000032f ),
    .Q(\blk00000001/sig000004e5 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000001d2  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000330 ),
    .Q(\blk00000001/sig000004e6 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000001d1  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000331 ),
    .Q(\blk00000001/sig000004e7 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000001d0  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000332 ),
    .Q(\blk00000001/sig000004e8 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000001cf  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000333 ),
    .Q(\blk00000001/sig000004e9 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000001ce  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000334 ),
    .Q(\blk00000001/sig000004ea )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000001cd  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000335 ),
    .Q(\blk00000001/sig000004eb )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000001cc  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000336 ),
    .Q(\blk00000001/sig000004ec )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000001cb  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000337 ),
    .Q(\blk00000001/sig000004ed )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000001ca  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000338 ),
    .Q(\blk00000001/sig000004ee )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000001c9  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000339 ),
    .Q(\blk00000001/sig000004ef )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000001c8  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig0000033a ),
    .Q(\blk00000001/sig000004f0 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000001c7  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig0000033b ),
    .Q(\blk00000001/sig000004f1 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000001c6  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig0000033c ),
    .Q(\blk00000001/sig000004f2 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000001c5  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig0000033d ),
    .Q(\blk00000001/sig000004f3 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000001c4  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig0000033e ),
    .Q(\blk00000001/sig000004f4 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000001c3  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig0000033f ),
    .Q(\blk00000001/sig000004f5 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000001c2  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000340 ),
    .Q(\blk00000001/sig000004f6 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000001c1  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig0000031d ),
    .Q(\blk00000001/sig0000047f )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000001c0  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig0000031e ),
    .Q(\blk00000001/sig00000480 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000001bf  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig0000031f ),
    .Q(\blk00000001/sig00000481 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000001be  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000320 ),
    .Q(\blk00000001/sig00000482 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000001bd  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000321 ),
    .Q(\blk00000001/sig00000483 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000001bc  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000322 ),
    .Q(\blk00000001/sig00000484 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000001bb  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000323 ),
    .Q(\blk00000001/sig00000485 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000001ba  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000324 ),
    .Q(\blk00000001/sig00000486 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000001b9  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000325 ),
    .Q(\blk00000001/sig00000487 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000001b8  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000326 ),
    .Q(\blk00000001/sig00000488 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000001b7  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000327 ),
    .Q(\blk00000001/sig00000489 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000001b6  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000328 ),
    .Q(\blk00000001/sig0000048a )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000001b5  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000329 ),
    .Q(\blk00000001/sig0000048b )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000001b4  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig0000032a ),
    .Q(\blk00000001/sig0000048c )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000001b3  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig0000032b ),
    .Q(\blk00000001/sig0000048d )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000001b2  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig0000032c ),
    .Q(\blk00000001/sig0000048e )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000001b1  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig0000032d ),
    .Q(\blk00000001/sig0000048f )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000001b0  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig0000032e ),
    .Q(\blk00000001/sig00000490 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000001af  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000002e3 ),
    .Q(\blk00000001/sig0000046e )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000001ae  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000002e4 ),
    .Q(\blk00000001/sig0000046f )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000001ad  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000002e5 ),
    .Q(\blk00000001/sig00000470 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000001ac  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000002e6 ),
    .Q(\blk00000001/sig00000471 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000001ab  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000002e7 ),
    .Q(\blk00000001/sig00000472 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000001aa  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000002e8 ),
    .Q(\blk00000001/sig00000473 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000001a9  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000002e9 ),
    .Q(\blk00000001/sig00000474 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000001a8  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000002ea ),
    .Q(\blk00000001/sig00000475 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000001a7  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000002eb ),
    .Q(\blk00000001/sig00000476 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000001a6  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000002ec ),
    .Q(\blk00000001/sig00000477 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000001a5  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000002ed ),
    .Q(\blk00000001/sig00000478 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000001a4  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000002ee ),
    .Q(\blk00000001/sig00000479 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000001a3  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000002ef ),
    .Q(\blk00000001/sig0000047a )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000001a2  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000002f0 ),
    .Q(\blk00000001/sig0000047b )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000001a1  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000002f1 ),
    .Q(\blk00000001/sig0000047c )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000001a0  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000002f2 ),
    .Q(\blk00000001/sig0000047d )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000019f  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000002c0 ),
    .Q(\blk00000001/sig000003e7 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000019e  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000002c1 ),
    .Q(\blk00000001/sig000003e8 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000019d  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000002c2 ),
    .Q(\blk00000001/sig000003e9 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000019c  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000002c3 ),
    .Q(\blk00000001/sig000003ea )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000019b  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000002c4 ),
    .Q(\blk00000001/sig000003eb )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000019a  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000002c5 ),
    .Q(\blk00000001/sig000003ec )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000199  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000002c6 ),
    .Q(\blk00000001/sig000003ed )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000198  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000002c7 ),
    .Q(\blk00000001/sig000003ee )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000197  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000002c8 ),
    .Q(\blk00000001/sig000003ef )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000196  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000002c9 ),
    .Q(\blk00000001/sig000003f0 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000195  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000002ca ),
    .Q(\blk00000001/sig000003f1 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000194  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000002cb ),
    .Q(\blk00000001/sig000003f2 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000193  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000002cc ),
    .Q(\blk00000001/sig000003f3 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000192  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000002cd ),
    .Q(\blk00000001/sig000003f4 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000191  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000002ce ),
    .Q(\blk00000001/sig000003f5 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000190  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000002cf ),
    .Q(\blk00000001/sig000003f6 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000018f  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000002cf ),
    .Q(\blk00000001/sig000003f7 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000018e  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000542 ),
    .Q(\blk00000001/sig0000050a )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000018d  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000530 ),
    .Q(\blk00000001/sig0000050b )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000018c  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000531 ),
    .Q(\blk00000001/sig0000050c )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000018b  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000532 ),
    .Q(\blk00000001/sig0000050d )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000018a  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000533 ),
    .Q(\blk00000001/sig0000050e )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000189  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000534 ),
    .Q(\blk00000001/sig0000050f )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000188  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000535 ),
    .Q(\blk00000001/sig00000510 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000187  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000536 ),
    .Q(\blk00000001/sig00000511 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000186  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000537 ),
    .Q(\blk00000001/sig00000512 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000185  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000538 ),
    .Q(\blk00000001/sig00000513 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000184  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000539 ),
    .Q(\blk00000001/sig00000514 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000183  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig0000053a ),
    .Q(\blk00000001/sig00000515 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000182  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig0000053b ),
    .Q(\blk00000001/sig00000516 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000181  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig0000053c ),
    .Q(\blk00000001/sig00000517 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000180  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig0000053d ),
    .Q(\blk00000001/sig00000518 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000017f  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig0000053e ),
    .Q(\blk00000001/sig00000519 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000017e  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig0000053f ),
    .Q(\blk00000001/sig0000051a )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000017d  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000540 ),
    .Q(\blk00000001/sig0000051b )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000017c  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000541 ),
    .Q(\blk00000001/sig0000051c )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000017b  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000002d0 ),
    .Q(\blk00000001/sig0000043b )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000017a  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000002d1 ),
    .Q(\blk00000001/sig0000043c )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000179  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000002d2 ),
    .Q(\blk00000001/sig0000043d )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000178  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000002d3 ),
    .Q(\blk00000001/sig0000043e )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000177  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000002d4 ),
    .Q(\blk00000001/sig0000043f )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000176  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000002d5 ),
    .Q(\blk00000001/sig00000440 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000175  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000002d6 ),
    .Q(\blk00000001/sig00000441 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000174  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000002d7 ),
    .Q(\blk00000001/sig00000442 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000173  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000002d8 ),
    .Q(\blk00000001/sig00000443 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000172  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000002d9 ),
    .Q(\blk00000001/sig00000444 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000171  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000002da ),
    .Q(\blk00000001/sig00000445 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000170  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000002db ),
    .Q(\blk00000001/sig00000446 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000016f  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000002dc ),
    .Q(\blk00000001/sig00000447 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000016e  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000002dd ),
    .Q(\blk00000001/sig00000448 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000016d  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000002de ),
    .Q(\blk00000001/sig00000449 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000016c  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000002df ),
    .Q(\blk00000001/sig0000044a )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000016b  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000002e0 ),
    .Q(\blk00000001/sig0000044b )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000016a  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000002e1 ),
    .Q(\blk00000001/sig0000044c )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000169  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000002e2 ),
    .Q(\blk00000001/sig0000044d )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000168  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig0000028e ),
    .Q(\blk00000001/sig00000384 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000167  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig0000028f ),
    .Q(\blk00000001/sig00000385 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000166  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000290 ),
    .Q(\blk00000001/sig00000386 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000165  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000291 ),
    .Q(\blk00000001/sig00000387 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000164  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000292 ),
    .Q(\blk00000001/sig00000388 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000163  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000293 ),
    .Q(\blk00000001/sig00000389 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000162  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000294 ),
    .Q(\blk00000001/sig0000038a )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000161  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000295 ),
    .Q(\blk00000001/sig0000038b )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000160  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000296 ),
    .Q(\blk00000001/sig0000038c )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000015f  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000297 ),
    .Q(\blk00000001/sig0000038d )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000015e  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000298 ),
    .Q(\blk00000001/sig0000038e )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000015d  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000299 ),
    .Q(\blk00000001/sig0000038f )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000015c  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig0000029a ),
    .Q(\blk00000001/sig00000390 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000015b  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig0000029b ),
    .Q(\blk00000001/sig00000391 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000015a  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig0000029c ),
    .Q(\blk00000001/sig00000392 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000159  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig0000029d ),
    .Q(\blk00000001/sig00000393 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000158  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig0000029e ),
    .Q(\blk00000001/sig00000394 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000157  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig0000029f ),
    .Q(\blk00000001/sig00000395 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000156  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000002a0 ),
    .Q(\blk00000001/sig00000396 )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000155  (
    .C(aclk),
    .D(\blk00000001/sig0000003b ),
    .Q(\blk00000001/sig00000040 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000154  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig0000031b ),
    .Q(\blk00000001/sig000003d6 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000153  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig0000031a ),
    .Q(\blk00000001/sig000003d5 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000152  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000319 ),
    .Q(\blk00000001/sig000003d4 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000151  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000318 ),
    .Q(\blk00000001/sig000003d3 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000150  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000317 ),
    .Q(\blk00000001/sig000003d2 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000014f  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000316 ),
    .Q(\blk00000001/sig000003d1 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000014e  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000315 ),
    .Q(\blk00000001/sig000003d0 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000014d  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000314 ),
    .Q(\blk00000001/sig000003cf )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000014c  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000313 ),
    .Q(\blk00000001/sig000003ce )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000014b  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000312 ),
    .Q(\blk00000001/sig000003cd )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000014a  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000311 ),
    .Q(\blk00000001/sig000003cc )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000149  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000310 ),
    .Q(\blk00000001/sig000003cb )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000148  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig0000030f ),
    .Q(\blk00000001/sig000003ca )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000147  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig0000030e ),
    .Q(\blk00000001/sig000003c9 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000146  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig0000030d ),
    .Q(\blk00000001/sig000003c8 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000145  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig0000030c ),
    .Q(\blk00000001/sig000003c7 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000144  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig0000030b ),
    .Q(\blk00000001/sig0000045d )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000143  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig0000030a ),
    .Q(\blk00000001/sig0000045c )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000142  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000309 ),
    .Q(\blk00000001/sig0000045b )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000141  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000308 ),
    .Q(\blk00000001/sig0000045a )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000140  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000307 ),
    .Q(\blk00000001/sig00000459 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000013f  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000306 ),
    .Q(\blk00000001/sig00000458 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000013e  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000305 ),
    .Q(\blk00000001/sig00000457 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000013d  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000304 ),
    .Q(\blk00000001/sig00000456 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000013c  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000303 ),
    .Q(\blk00000001/sig00000455 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000013b  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000302 ),
    .Q(\blk00000001/sig00000454 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000013a  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000301 ),
    .Q(\blk00000001/sig00000453 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000139  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000300 ),
    .Q(\blk00000001/sig00000452 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000138  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000002ff ),
    .Q(\blk00000001/sig00000451 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000137  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000002fe ),
    .Q(\blk00000001/sig00000450 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000136  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000002fd ),
    .Q(\blk00000001/sig0000044f )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000135  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000002fc ),
    .Q(\blk00000001/sig0000044e )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000134  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000002fb ),
    .Q(\blk00000001/sig00000526 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000133  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000002fa ),
    .Q(\blk00000001/sig00000525 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000132  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000002f9 ),
    .Q(\blk00000001/sig00000524 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000131  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000002f8 ),
    .Q(\blk00000001/sig00000523 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000130  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000002f7 ),
    .Q(\blk00000001/sig00000522 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000012f  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000002f6 ),
    .Q(\blk00000001/sig00000521 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000012e  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000002f5 ),
    .Q(\blk00000001/sig00000520 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000012d  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000002f4 ),
    .Q(\blk00000001/sig0000051f )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000012c  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000002f3 ),
    .Q(\blk00000001/sig0000051e )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000012b  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig0000028d ),
    .Q(\blk00000001/sig0000052f )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000012a  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig0000028c ),
    .Q(\blk00000001/sig0000052e )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000129  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig0000028b ),
    .Q(\blk00000001/sig0000052d )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000128  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig0000028a ),
    .Q(\blk00000001/sig0000052c )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000127  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000289 ),
    .Q(\blk00000001/sig0000052b )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000126  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000288 ),
    .Q(\blk00000001/sig0000052a )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000125  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000287 ),
    .Q(\blk00000001/sig00000529 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000124  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000286 ),
    .Q(\blk00000001/sig00000528 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000123  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000285 ),
    .Q(\blk00000001/sig00000527 )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000122  (
    .C(aclk),
    .D(\blk00000001/sig000001e0 ),
    .Q(\blk00000001/sig00000051 )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000121  (
    .C(aclk),
    .D(\blk00000001/sig000001e1 ),
    .Q(\blk00000001/sig00000052 )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000120  (
    .C(aclk),
    .D(\blk00000001/sig000001e2 ),
    .Q(\blk00000001/sig00000053 )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000011f  (
    .C(aclk),
    .D(\blk00000001/sig000001e3 ),
    .Q(\blk00000001/sig00000054 )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000011e  (
    .C(aclk),
    .D(\blk00000001/sig000001e4 ),
    .Q(\blk00000001/sig00000055 )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000011d  (
    .C(aclk),
    .D(\blk00000001/sig000001e5 ),
    .Q(\blk00000001/sig00000056 )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000011c  (
    .C(aclk),
    .D(\blk00000001/sig000001e6 ),
    .Q(\blk00000001/sig00000057 )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000011b  (
    .C(aclk),
    .D(\blk00000001/sig000001e7 ),
    .Q(\blk00000001/sig00000058 )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000011a  (
    .C(aclk),
    .D(\blk00000001/sig000001e8 ),
    .Q(\blk00000001/sig00000059 )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000119  (
    .C(aclk),
    .D(\blk00000001/sig000001e9 ),
    .Q(\blk00000001/sig0000005a )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000118  (
    .C(aclk),
    .D(\blk00000001/sig000001ea ),
    .Q(\blk00000001/sig0000005b )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000117  (
    .C(aclk),
    .D(\blk00000001/sig000001eb ),
    .Q(\blk00000001/sig0000005c )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000116  (
    .C(aclk),
    .D(\blk00000001/sig000001ec ),
    .Q(\blk00000001/sig0000005d )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000115  (
    .C(aclk),
    .D(\blk00000001/sig000001ed ),
    .Q(\blk00000001/sig0000005e )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000114  (
    .C(aclk),
    .D(\blk00000001/sig000001ee ),
    .Q(\blk00000001/sig0000005f )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000113  (
    .C(aclk),
    .D(\blk00000001/sig000001ef ),
    .Q(\blk00000001/sig00000060 )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000112  (
    .C(aclk),
    .D(\blk00000001/sig000001f0 ),
    .Q(\blk00000001/sig00000061 )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000111  (
    .C(aclk),
    .D(\blk00000001/sig000001f1 ),
    .Q(\blk00000001/sig00000062 )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000110  (
    .C(aclk),
    .D(\blk00000001/sig000001f2 ),
    .Q(\blk00000001/sig00000063 )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000010f  (
    .C(aclk),
    .D(\blk00000001/sig000001f3 ),
    .Q(\blk00000001/sig00000064 )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000010e  (
    .C(aclk),
    .D(\blk00000001/sig000001f4 ),
    .Q(\blk00000001/sig00000065 )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000010d  (
    .C(aclk),
    .D(\blk00000001/sig000001f5 ),
    .Q(\blk00000001/sig00000066 )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000010c  (
    .C(aclk),
    .D(\blk00000001/sig000001f6 ),
    .Q(\blk00000001/sig00000067 )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000010b  (
    .C(aclk),
    .D(\blk00000001/sig000001f7 ),
    .Q(\blk00000001/sig00000068 )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000010a  (
    .C(aclk),
    .D(\blk00000001/sig000001f8 ),
    .Q(\blk00000001/sig00000069 )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000109  (
    .C(aclk),
    .D(\blk00000001/sig000001f9 ),
    .Q(\blk00000001/sig00000271 )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000108  (
    .C(aclk),
    .D(\blk00000001/sig000001fa ),
    .Q(\blk00000001/sig00000272 )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000107  (
    .C(aclk),
    .D(\blk00000001/sig000001fb ),
    .Q(\blk00000001/sig00000273 )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000106  (
    .C(aclk),
    .D(\blk00000001/sig000001fc ),
    .Q(\blk00000001/sig00000274 )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000105  (
    .C(aclk),
    .D(\blk00000001/sig000001fd ),
    .Q(\blk00000001/sig00000275 )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000104  (
    .C(aclk),
    .D(\blk00000001/sig000001fe ),
    .Q(\blk00000001/sig00000276 )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000103  (
    .C(aclk),
    .D(\blk00000001/sig000001ff ),
    .Q(\blk00000001/sig00000277 )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000102  (
    .C(aclk),
    .D(\blk00000001/sig00000200 ),
    .Q(\blk00000001/sig00000278 )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000101  (
    .C(aclk),
    .D(\blk00000001/sig00000201 ),
    .Q(\blk00000001/sig00000279 )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000100  (
    .C(aclk),
    .D(\blk00000001/sig00000202 ),
    .Q(\blk00000001/sig0000027a )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000000ff  (
    .C(aclk),
    .D(\blk00000001/sig00000203 ),
    .Q(\blk00000001/sig0000027b )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000000fe  (
    .C(aclk),
    .D(\blk00000001/sig00000204 ),
    .Q(\blk00000001/sig0000027c )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000000fd  (
    .C(aclk),
    .D(\blk00000001/sig00000205 ),
    .Q(\blk00000001/sig0000027d )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000000fc  (
    .C(aclk),
    .D(\blk00000001/sig00000206 ),
    .Q(\blk00000001/sig0000027e )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000000fb  (
    .C(aclk),
    .D(\blk00000001/sig00000207 ),
    .Q(\blk00000001/sig0000027f )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000000fa  (
    .C(aclk),
    .D(\blk00000001/sig00000208 ),
    .Q(\blk00000001/sig00000280 )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000000f9  (
    .C(aclk),
    .D(\blk00000001/sig00000209 ),
    .Q(\blk00000001/sig00000281 )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000000f8  (
    .C(aclk),
    .D(\blk00000001/sig0000020a ),
    .Q(\blk00000001/sig00000282 )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000000f7  (
    .C(aclk),
    .D(\blk00000001/sig0000020b ),
    .Q(\blk00000001/sig00000283 )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000000f6  (
    .C(aclk),
    .D(\blk00000001/sig0000020c ),
    .Q(\blk00000001/sig00000239 )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000000f5  (
    .C(aclk),
    .D(\blk00000001/sig0000020d ),
    .Q(\blk00000001/sig0000023a )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000000f4  (
    .C(aclk),
    .D(\blk00000001/sig0000020e ),
    .Q(\blk00000001/sig0000023b )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000000f3  (
    .C(aclk),
    .D(\blk00000001/sig0000020f ),
    .Q(\blk00000001/sig0000023c )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000000f2  (
    .C(aclk),
    .D(\blk00000001/sig00000210 ),
    .Q(\blk00000001/sig0000023d )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000000f1  (
    .C(aclk),
    .D(\blk00000001/sig00000211 ),
    .Q(\blk00000001/sig0000023e )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000000f0  (
    .C(aclk),
    .D(\blk00000001/sig00000212 ),
    .Q(\blk00000001/sig0000023f )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000000ef  (
    .C(aclk),
    .D(\blk00000001/sig00000213 ),
    .Q(\blk00000001/sig00000240 )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000000ee  (
    .C(aclk),
    .D(\blk00000001/sig00000214 ),
    .Q(\blk00000001/sig00000241 )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000000ed  (
    .C(aclk),
    .D(\blk00000001/sig00000215 ),
    .Q(\blk00000001/sig00000242 )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000000ec  (
    .C(aclk),
    .D(\blk00000001/sig00000216 ),
    .Q(\blk00000001/sig00000243 )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000000eb  (
    .C(aclk),
    .D(\blk00000001/sig00000217 ),
    .Q(\blk00000001/sig00000244 )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000000ea  (
    .C(aclk),
    .D(\blk00000001/sig00000218 ),
    .Q(\blk00000001/sig00000245 )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000000e9  (
    .C(aclk),
    .D(\blk00000001/sig00000219 ),
    .Q(\blk00000001/sig00000246 )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000000e8  (
    .C(aclk),
    .D(\blk00000001/sig0000021a ),
    .Q(\blk00000001/sig00000247 )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000000e7  (
    .C(aclk),
    .D(\blk00000001/sig0000021b ),
    .Q(\blk00000001/sig00000248 )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000000e6  (
    .C(aclk),
    .D(\blk00000001/sig0000021c ),
    .Q(\blk00000001/sig00000249 )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000000e5  (
    .C(aclk),
    .D(\blk00000001/sig0000021d ),
    .Q(\blk00000001/sig0000024a )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000000e4  (
    .C(aclk),
    .D(\blk00000001/sig0000021e ),
    .Q(\blk00000001/sig0000024b )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000000e3  (
    .C(aclk),
    .D(\blk00000001/sig0000021f ),
    .Q(\blk00000001/sig0000024c )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000000e2  (
    .C(aclk),
    .D(\blk00000001/sig00000220 ),
    .Q(\blk00000001/sig0000024d )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000000e1  (
    .C(aclk),
    .D(\blk00000001/sig00000221 ),
    .Q(\blk00000001/sig0000024e )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000000e0  (
    .C(aclk),
    .D(\blk00000001/sig00000222 ),
    .Q(\blk00000001/sig0000024f )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000000df  (
    .C(aclk),
    .D(\blk00000001/sig00000223 ),
    .Q(\blk00000001/sig00000250 )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000000de  (
    .C(aclk),
    .D(\blk00000001/sig00000224 ),
    .Q(\blk00000001/sig00000251 )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000000dd  (
    .C(aclk),
    .D(\blk00000001/sig00000225 ),
    .Q(\blk00000001/sig00000252 )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000000dc  (
    .C(aclk),
    .D(\blk00000001/sig00000226 ),
    .Q(\blk00000001/sig00000253 )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000000db  (
    .C(aclk),
    .D(\blk00000001/sig00000227 ),
    .Q(\blk00000001/sig0000020b )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000000da  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000268 ),
    .Q(\blk00000001/sig00000254 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000000d9  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000269 ),
    .Q(\blk00000001/sig00000255 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000000d8  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig0000026a ),
    .Q(\blk00000001/sig00000258 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000000d7  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig0000026b ),
    .Q(\blk00000001/sig00000256 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000000d6  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig0000026c ),
    .Q(\blk00000001/sig00000257 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000000d5  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000254 ),
    .Q(\blk00000001/sig0000026d )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000000d4  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000255 ),
    .Q(\blk00000001/sig0000026e )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000000d3  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000258 ),
    .Q(\blk00000001/sig0000026f )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000000d2  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000256 ),
    .Q(\blk00000001/sig00000270 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000000d1  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000257 ),
    .Q(\blk00000001/sig00000238 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000000d0  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000228 ),
    .Q(\blk00000001/sig00000259 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000000cf  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000229 ),
    .Q(\blk00000001/sig0000025a )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000000ce  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig0000022a ),
    .Q(\blk00000001/sig0000025b )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000000cd  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig0000022b ),
    .Q(\blk00000001/sig0000025c )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000000cc  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig0000022c ),
    .Q(\blk00000001/sig0000025d )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000000cb  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig0000022d ),
    .Q(\blk00000001/sig0000025e )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000000ca  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig0000022e ),
    .Q(\blk00000001/sig0000025f )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000000c9  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig0000022f ),
    .Q(\blk00000001/sig00000260 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000000c8  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000230 ),
    .Q(\blk00000001/sig00000261 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000000c7  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000231 ),
    .Q(\blk00000001/sig00000262 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000000c6  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000232 ),
    .Q(\blk00000001/sig00000263 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000000c5  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000233 ),
    .Q(\blk00000001/sig00000264 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000000c4  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000234 ),
    .Q(\blk00000001/sig00000265 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000000c3  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000235 ),
    .Q(\blk00000001/sig00000266 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000000c2  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000236 ),
    .Q(\blk00000001/sig00000267 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000000c1  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000237 ),
    .Q(\blk00000001/sig00000227 )
  );
  DSP48A1 #(
    .A0REG ( 0 ),
    .A1REG ( 1 ),
    .B0REG ( 0 ),
    .B1REG ( 1 ),
    .CARRYINREG ( 0 ),
    .CARRYINSEL ( "OPMODE5" ),
    .CREG ( 1 ),
    .DREG ( 1 ),
    .MREG ( 1 ),
    .OPMODEREG ( 1 ),
    .PREG ( 1 ),
    .RSTTYPE ( "SYNC" ),
    .CARRYOUTREG ( 0 ))
  \blk00000001/blk000000ad  (
    .CECARRYIN(\blk00000001/sig0000051d ),
    .RSTC(\blk00000001/sig0000051d ),
    .RSTCARRYIN(\blk00000001/sig0000051d ),
    .CED(\blk00000001/sig0000003a ),
    .RSTD(\blk00000001/sig0000051d ),
    .CEOPMODE(\blk00000001/sig0000003a ),
    .CEC(\blk00000001/sig0000003a ),
    .CARRYOUTF(\NLW_blk00000001/blk000000ad_CARRYOUTF_UNCONNECTED ),
    .RSTOPMODE(\blk00000001/sig0000051d ),
    .RSTM(\blk00000001/sig0000051d ),
    .CLK(aclk),
    .RSTB(\blk00000001/sig0000051d ),
    .CEM(\blk00000001/sig0000003a ),
    .CEB(\blk00000001/sig0000003a ),
    .CARRYIN(\blk00000001/sig0000051d ),
    .CEP(\blk00000001/sig0000003a ),
    .CEA(\blk00000001/sig0000003a ),
    .CARRYOUT(\NLW_blk00000001/blk000000ad_CARRYOUT_UNCONNECTED ),
    .RSTA(\blk00000001/sig0000051d ),
    .RSTP(\blk00000001/sig0000051d ),
    .B({\blk00000001/sig000001ab , \blk00000001/sig000001ab , \blk00000001/sig000001df , \blk00000001/sig000001de , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d }),
    .BCOUT({\NLW_blk00000001/blk000000ad_BCOUT<17>_UNCONNECTED , \NLW_blk00000001/blk000000ad_BCOUT<16>_UNCONNECTED ,
\NLW_blk00000001/blk000000ad_BCOUT<15>_UNCONNECTED , \NLW_blk00000001/blk000000ad_BCOUT<14>_UNCONNECTED ,
\NLW_blk00000001/blk000000ad_BCOUT<13>_UNCONNECTED , \NLW_blk00000001/blk000000ad_BCOUT<12>_UNCONNECTED ,
\NLW_blk00000001/blk000000ad_BCOUT<11>_UNCONNECTED , \NLW_blk00000001/blk000000ad_BCOUT<10>_UNCONNECTED ,
\NLW_blk00000001/blk000000ad_BCOUT<9>_UNCONNECTED , \NLW_blk00000001/blk000000ad_BCOUT<8>_UNCONNECTED ,
\NLW_blk00000001/blk000000ad_BCOUT<7>_UNCONNECTED , \NLW_blk00000001/blk000000ad_BCOUT<6>_UNCONNECTED ,
\NLW_blk00000001/blk000000ad_BCOUT<5>_UNCONNECTED , \NLW_blk00000001/blk000000ad_BCOUT<4>_UNCONNECTED ,
\NLW_blk00000001/blk000000ad_BCOUT<3>_UNCONNECTED , \NLW_blk00000001/blk000000ad_BCOUT<2>_UNCONNECTED ,
\NLW_blk00000001/blk000000ad_BCOUT<1>_UNCONNECTED , \NLW_blk00000001/blk000000ad_BCOUT<0>_UNCONNECTED }),
    .PCIN({\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d }),
    .C({\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000003a , \blk00000001/sig000001aa ,
\blk00000001/sig000001a9 , \blk00000001/sig000001a8 , \blk00000001/sig000001a7 , \blk00000001/sig000001a6 , \blk00000001/sig000001a5 ,
\blk00000001/sig000001a4 , \blk00000001/sig000001a3 , \blk00000001/sig000001a2 , \blk00000001/sig000001a1 , \blk00000001/sig000001a0 ,
\blk00000001/sig0000019f , \blk00000001/sig0000019e , \blk00000001/sig0000019d , \blk00000001/sig0000019c , \blk00000001/sig0000019b ,
\blk00000001/sig0000019a , \blk00000001/sig00000199 , \blk00000001/sig00000198 , \blk00000001/sig00000197 , \blk00000001/sig00000196 ,
\blk00000001/sig00000195 , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d }),
    .P({\NLW_blk00000001/blk000000ad_P<47>_UNCONNECTED , \NLW_blk00000001/blk000000ad_P<46>_UNCONNECTED ,
\NLW_blk00000001/blk000000ad_P<45>_UNCONNECTED , \NLW_blk00000001/blk000000ad_P<44>_UNCONNECTED , \NLW_blk00000001/blk000000ad_P<43>_UNCONNECTED ,
\NLW_blk00000001/blk000000ad_P<42>_UNCONNECTED , \NLW_blk00000001/blk000000ad_P<41>_UNCONNECTED , \blk00000001/sig0000009c , \blk00000001/sig0000009b
, \blk00000001/sig0000009a , \blk00000001/sig00000099 , \blk00000001/sig00000098 , \blk00000001/sig00000097 , \blk00000001/sig00000096 ,
\blk00000001/sig00000095 , \blk00000001/sig00000094 , \blk00000001/sig00000093 , \blk00000001/sig00000092 , \blk00000001/sig00000091 ,
\blk00000001/sig00000090 , \blk00000001/sig0000008f , \blk00000001/sig0000008e , \blk00000001/sig0000008d , \blk00000001/sig0000008c ,
\blk00000001/sig0000008b , \blk00000001/sig0000008a , \NLW_blk00000001/blk000000ad_P<21>_UNCONNECTED , \NLW_blk00000001/blk000000ad_P<20>_UNCONNECTED
, \NLW_blk00000001/blk000000ad_P<19>_UNCONNECTED , \NLW_blk00000001/blk000000ad_P<18>_UNCONNECTED , \NLW_blk00000001/blk000000ad_P<17>_UNCONNECTED ,
\NLW_blk00000001/blk000000ad_P<16>_UNCONNECTED , \NLW_blk00000001/blk000000ad_P<15>_UNCONNECTED , \NLW_blk00000001/blk000000ad_P<14>_UNCONNECTED ,
\NLW_blk00000001/blk000000ad_P<13>_UNCONNECTED , \NLW_blk00000001/blk000000ad_P<12>_UNCONNECTED , \NLW_blk00000001/blk000000ad_P<11>_UNCONNECTED ,
\NLW_blk00000001/blk000000ad_P<10>_UNCONNECTED , \NLW_blk00000001/blk000000ad_P<9>_UNCONNECTED , \NLW_blk00000001/blk000000ad_P<8>_UNCONNECTED ,
\NLW_blk00000001/blk000000ad_P<7>_UNCONNECTED , \NLW_blk00000001/blk000000ad_P<6>_UNCONNECTED , \NLW_blk00000001/blk000000ad_P<5>_UNCONNECTED ,
\NLW_blk00000001/blk000000ad_P<4>_UNCONNECTED , \NLW_blk00000001/blk000000ad_P<3>_UNCONNECTED , \NLW_blk00000001/blk000000ad_P<2>_UNCONNECTED ,
\NLW_blk00000001/blk000000ad_P<1>_UNCONNECTED , \NLW_blk00000001/blk000000ad_P<0>_UNCONNECTED }),
    .OPMODE({\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000003a ,
\blk00000001/sig0000003a , \blk00000001/sig0000051d , \blk00000001/sig0000003a }),
    .D({\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d ,
\blk00000001/sig0000051d , \blk00000001/sig0000051d , \blk00000001/sig0000051d }),
    .PCOUT({\NLW_blk00000001/blk000000ad_PCOUT<47>_UNCONNECTED , \NLW_blk00000001/blk000000ad_PCOUT<46>_UNCONNECTED ,
\NLW_blk00000001/blk000000ad_PCOUT<45>_UNCONNECTED , \NLW_blk00000001/blk000000ad_PCOUT<44>_UNCONNECTED ,
\NLW_blk00000001/blk000000ad_PCOUT<43>_UNCONNECTED , \NLW_blk00000001/blk000000ad_PCOUT<42>_UNCONNECTED ,
\NLW_blk00000001/blk000000ad_PCOUT<41>_UNCONNECTED , \NLW_blk00000001/blk000000ad_PCOUT<40>_UNCONNECTED ,
\NLW_blk00000001/blk000000ad_PCOUT<39>_UNCONNECTED , \NLW_blk00000001/blk000000ad_PCOUT<38>_UNCONNECTED ,
\NLW_blk00000001/blk000000ad_PCOUT<37>_UNCONNECTED , \NLW_blk00000001/blk000000ad_PCOUT<36>_UNCONNECTED ,
\NLW_blk00000001/blk000000ad_PCOUT<35>_UNCONNECTED , \NLW_blk00000001/blk000000ad_PCOUT<34>_UNCONNECTED ,
\NLW_blk00000001/blk000000ad_PCOUT<33>_UNCONNECTED , \NLW_blk00000001/blk000000ad_PCOUT<32>_UNCONNECTED ,
\NLW_blk00000001/blk000000ad_PCOUT<31>_UNCONNECTED , \NLW_blk00000001/blk000000ad_PCOUT<30>_UNCONNECTED ,
\NLW_blk00000001/blk000000ad_PCOUT<29>_UNCONNECTED , \NLW_blk00000001/blk000000ad_PCOUT<28>_UNCONNECTED ,
\NLW_blk00000001/blk000000ad_PCOUT<27>_UNCONNECTED , \NLW_blk00000001/blk000000ad_PCOUT<26>_UNCONNECTED ,
\NLW_blk00000001/blk000000ad_PCOUT<25>_UNCONNECTED , \NLW_blk00000001/blk000000ad_PCOUT<24>_UNCONNECTED ,
\NLW_blk00000001/blk000000ad_PCOUT<23>_UNCONNECTED , \NLW_blk00000001/blk000000ad_PCOUT<22>_UNCONNECTED ,
\NLW_blk00000001/blk000000ad_PCOUT<21>_UNCONNECTED , \NLW_blk00000001/blk000000ad_PCOUT<20>_UNCONNECTED ,
\NLW_blk00000001/blk000000ad_PCOUT<19>_UNCONNECTED , \NLW_blk00000001/blk000000ad_PCOUT<18>_UNCONNECTED ,
\NLW_blk00000001/blk000000ad_PCOUT<17>_UNCONNECTED , \NLW_blk00000001/blk000000ad_PCOUT<16>_UNCONNECTED ,
\NLW_blk00000001/blk000000ad_PCOUT<15>_UNCONNECTED , \NLW_blk00000001/blk000000ad_PCOUT<14>_UNCONNECTED ,
\NLW_blk00000001/blk000000ad_PCOUT<13>_UNCONNECTED , \NLW_blk00000001/blk000000ad_PCOUT<12>_UNCONNECTED ,
\NLW_blk00000001/blk000000ad_PCOUT<11>_UNCONNECTED , \NLW_blk00000001/blk000000ad_PCOUT<10>_UNCONNECTED ,
\NLW_blk00000001/blk000000ad_PCOUT<9>_UNCONNECTED , \NLW_blk00000001/blk000000ad_PCOUT<8>_UNCONNECTED ,
\NLW_blk00000001/blk000000ad_PCOUT<7>_UNCONNECTED , \NLW_blk00000001/blk000000ad_PCOUT<6>_UNCONNECTED ,
\NLW_blk00000001/blk000000ad_PCOUT<5>_UNCONNECTED , \NLW_blk00000001/blk000000ad_PCOUT<4>_UNCONNECTED ,
\NLW_blk00000001/blk000000ad_PCOUT<3>_UNCONNECTED , \NLW_blk00000001/blk000000ad_PCOUT<2>_UNCONNECTED ,
\NLW_blk00000001/blk000000ad_PCOUT<1>_UNCONNECTED , \NLW_blk00000001/blk000000ad_PCOUT<0>_UNCONNECTED }),
    .A({\blk00000001/sig0000003a , \blk00000001/sig0000003a , \blk00000001/sig0000003a , \blk00000001/sig0000003a , \blk00000001/sig000001cb ,
\blk00000001/sig000001ca , \blk00000001/sig000001c9 , \blk00000001/sig000001c8 , \blk00000001/sig000001c7 , \blk00000001/sig000001c6 ,
\blk00000001/sig000001c5 , \blk00000001/sig000001c4 , \blk00000001/sig000001c3 , \blk00000001/sig000001c2 , \blk00000001/sig000001c1 ,
\blk00000001/sig000001c0 , \blk00000001/sig000001bf , \blk00000001/sig000001be }),
    .M({\NLW_blk00000001/blk000000ad_M<35>_UNCONNECTED , \NLW_blk00000001/blk000000ad_M<34>_UNCONNECTED ,
\NLW_blk00000001/blk000000ad_M<33>_UNCONNECTED , \NLW_blk00000001/blk000000ad_M<32>_UNCONNECTED , \NLW_blk00000001/blk000000ad_M<31>_UNCONNECTED ,
\NLW_blk00000001/blk000000ad_M<30>_UNCONNECTED , \NLW_blk00000001/blk000000ad_M<29>_UNCONNECTED , \NLW_blk00000001/blk000000ad_M<28>_UNCONNECTED ,
\NLW_blk00000001/blk000000ad_M<27>_UNCONNECTED , \NLW_blk00000001/blk000000ad_M<26>_UNCONNECTED , \NLW_blk00000001/blk000000ad_M<25>_UNCONNECTED ,
\NLW_blk00000001/blk000000ad_M<24>_UNCONNECTED , \NLW_blk00000001/blk000000ad_M<23>_UNCONNECTED , \NLW_blk00000001/blk000000ad_M<22>_UNCONNECTED ,
\NLW_blk00000001/blk000000ad_M<21>_UNCONNECTED , \NLW_blk00000001/blk000000ad_M<20>_UNCONNECTED , \NLW_blk00000001/blk000000ad_M<19>_UNCONNECTED ,
\NLW_blk00000001/blk000000ad_M<18>_UNCONNECTED , \NLW_blk00000001/blk000000ad_M<17>_UNCONNECTED , \NLW_blk00000001/blk000000ad_M<16>_UNCONNECTED ,
\NLW_blk00000001/blk000000ad_M<15>_UNCONNECTED , \NLW_blk00000001/blk000000ad_M<14>_UNCONNECTED , \NLW_blk00000001/blk000000ad_M<13>_UNCONNECTED ,
\NLW_blk00000001/blk000000ad_M<12>_UNCONNECTED , \NLW_blk00000001/blk000000ad_M<11>_UNCONNECTED , \NLW_blk00000001/blk000000ad_M<10>_UNCONNECTED ,
\NLW_blk00000001/blk000000ad_M<9>_UNCONNECTED , \NLW_blk00000001/blk000000ad_M<8>_UNCONNECTED , \NLW_blk00000001/blk000000ad_M<7>_UNCONNECTED ,
\NLW_blk00000001/blk000000ad_M<6>_UNCONNECTED , \NLW_blk00000001/blk000000ad_M<5>_UNCONNECTED , \NLW_blk00000001/blk000000ad_M<4>_UNCONNECTED ,
\NLW_blk00000001/blk000000ad_M<3>_UNCONNECTED , \NLW_blk00000001/blk000000ad_M<2>_UNCONNECTED , \NLW_blk00000001/blk000000ad_M<1>_UNCONNECTED ,
\NLW_blk00000001/blk000000ad_M<0>_UNCONNECTED })
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000000ac  (
    .C(aclk),
    .D(\blk00000001/sig000001cc ),
    .Q(\blk00000001/sig000001be )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000000ab  (
    .C(aclk),
    .D(\blk00000001/sig000001cd ),
    .Q(\blk00000001/sig000001bf )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000000aa  (
    .C(aclk),
    .D(\blk00000001/sig000001ce ),
    .Q(\blk00000001/sig000001c0 )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000000a9  (
    .C(aclk),
    .D(\blk00000001/sig000001cf ),
    .Q(\blk00000001/sig000001c1 )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000000a8  (
    .C(aclk),
    .D(\blk00000001/sig000001d0 ),
    .Q(\blk00000001/sig000001c2 )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000000a7  (
    .C(aclk),
    .D(\blk00000001/sig000001d1 ),
    .Q(\blk00000001/sig000001c3 )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000000a6  (
    .C(aclk),
    .D(\blk00000001/sig000001d2 ),
    .Q(\blk00000001/sig000001c4 )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000000a5  (
    .C(aclk),
    .D(\blk00000001/sig000001d3 ),
    .Q(\blk00000001/sig000001c5 )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000000a4  (
    .C(aclk),
    .D(\blk00000001/sig000001d4 ),
    .Q(\blk00000001/sig000001c6 )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000000a3  (
    .C(aclk),
    .D(\blk00000001/sig000001d5 ),
    .Q(\blk00000001/sig000001c7 )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000000a2  (
    .C(aclk),
    .D(\blk00000001/sig000001d6 ),
    .Q(\blk00000001/sig000001c8 )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000000a1  (
    .C(aclk),
    .D(\blk00000001/sig000001d7 ),
    .Q(\blk00000001/sig000001c9 )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000000a0  (
    .C(aclk),
    .D(\blk00000001/sig000001d8 ),
    .Q(\blk00000001/sig000001ca )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000009f  (
    .C(aclk),
    .D(\blk00000001/sig000001d9 ),
    .Q(\blk00000001/sig000001cb )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000009e  (
    .C(aclk),
    .D(\blk00000001/sig0000051d ),
    .Q(\blk00000001/sig00000193 )
  );
  FD   \blk00000001/blk0000009d  (
    .C(aclk),
    .D(\blk00000001/sig00000186 ),
    .Q(\blk00000001/sig000000aa )
  );
  FD   \blk00000001/blk0000009c  (
    .C(aclk),
    .D(\blk00000001/sig00000187 ),
    .Q(\blk00000001/sig000000ab )
  );
  FD   \blk00000001/blk0000009b  (
    .C(aclk),
    .D(\blk00000001/sig00000188 ),
    .Q(\blk00000001/sig000000ac )
  );
  FD   \blk00000001/blk0000009a  (
    .C(aclk),
    .D(\blk00000001/sig00000189 ),
    .Q(\blk00000001/sig000000ad )
  );
  FD   \blk00000001/blk00000099  (
    .C(aclk),
    .D(\blk00000001/sig0000018a ),
    .Q(\blk00000001/sig000000ae )
  );
  FD   \blk00000001/blk00000098  (
    .C(aclk),
    .D(\blk00000001/sig0000018b ),
    .Q(\blk00000001/sig000000af )
  );
  FD   \blk00000001/blk00000097  (
    .C(aclk),
    .D(\blk00000001/sig0000018c ),
    .Q(\blk00000001/sig000000b0 )
  );
  FD   \blk00000001/blk00000096  (
    .C(aclk),
    .D(\blk00000001/sig0000018d ),
    .Q(\blk00000001/sig000000b1 )
  );
  FD   \blk00000001/blk00000095  (
    .C(aclk),
    .D(\blk00000001/sig0000018e ),
    .Q(\blk00000001/sig000000b2 )
  );
  FD   \blk00000001/blk00000094  (
    .C(aclk),
    .D(\blk00000001/sig0000018f ),
    .Q(\blk00000001/sig000000b3 )
  );
  FD   \blk00000001/blk00000093  (
    .C(aclk),
    .D(\blk00000001/sig00000190 ),
    .Q(\blk00000001/sig000000b4 )
  );
  FD   \blk00000001/blk00000092  (
    .C(aclk),
    .D(\blk00000001/sig00000191 ),
    .Q(\blk00000001/sig000000b5 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000091  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000184 ),
    .Q(\blk00000001/sig000000c1 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000090  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000182 ),
    .Q(\blk00000001/sig000000c2 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000008f  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000180 ),
    .Q(\blk00000001/sig000000c3 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000008e  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig0000017e ),
    .Q(\blk00000001/sig000000c4 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000008d  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig0000017c ),
    .Q(\blk00000001/sig000000c5 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000008c  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig0000017a ),
    .Q(\blk00000001/sig000000c6 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000008b  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000179 ),
    .Q(\blk00000001/sig00000167 )
  );
  MUXCY   \blk00000001/blk0000008a  (
    .CI(\blk00000001/sig00000168 ),
    .DI(\blk00000001/sig0000051d ),
    .S(\blk00000001/sig0000056d ),
    .O(\blk00000001/sig00000185 )
  );
  XORCY   \blk00000001/blk00000089  (
    .CI(\blk00000001/sig00000168 ),
    .LI(\blk00000001/sig0000056d ),
    .O(\blk00000001/sig00000184 )
  );
  MUXCY   \blk00000001/blk00000088  (
    .CI(\blk00000001/sig00000185 ),
    .DI(\blk00000001/sig0000051d ),
    .S(\blk00000001/sig0000056c ),
    .O(\blk00000001/sig00000183 )
  );
  XORCY   \blk00000001/blk00000087  (
    .CI(\blk00000001/sig00000185 ),
    .LI(\blk00000001/sig0000056c ),
    .O(\blk00000001/sig00000182 )
  );
  MUXCY   \blk00000001/blk00000086  (
    .CI(\blk00000001/sig00000183 ),
    .DI(\blk00000001/sig0000051d ),
    .S(\blk00000001/sig0000056b ),
    .O(\blk00000001/sig00000181 )
  );
  XORCY   \blk00000001/blk00000085  (
    .CI(\blk00000001/sig00000183 ),
    .LI(\blk00000001/sig0000056b ),
    .O(\blk00000001/sig00000180 )
  );
  MUXCY   \blk00000001/blk00000084  (
    .CI(\blk00000001/sig00000181 ),
    .DI(\blk00000001/sig0000051d ),
    .S(\blk00000001/sig0000056a ),
    .O(\blk00000001/sig0000017f )
  );
  XORCY   \blk00000001/blk00000083  (
    .CI(\blk00000001/sig00000181 ),
    .LI(\blk00000001/sig0000056a ),
    .O(\blk00000001/sig0000017e )
  );
  MUXCY   \blk00000001/blk00000082  (
    .CI(\blk00000001/sig0000017f ),
    .DI(\blk00000001/sig0000051d ),
    .S(\blk00000001/sig00000569 ),
    .O(\blk00000001/sig0000017d )
  );
  XORCY   \blk00000001/blk00000081  (
    .CI(\blk00000001/sig0000017f ),
    .LI(\blk00000001/sig00000569 ),
    .O(\blk00000001/sig0000017c )
  );
  MUXCY   \blk00000001/blk00000080  (
    .CI(\blk00000001/sig0000017d ),
    .DI(\blk00000001/sig0000051d ),
    .S(\blk00000001/sig00000568 ),
    .O(\blk00000001/sig0000017b )
  );
  XORCY   \blk00000001/blk0000007f  (
    .CI(\blk00000001/sig0000017d ),
    .LI(\blk00000001/sig00000568 ),
    .O(\blk00000001/sig0000017a )
  );
  XORCY   \blk00000001/blk0000007e  (
    .CI(\blk00000001/sig0000017b ),
    .LI(\blk00000001/sig0000003a ),
    .O(\blk00000001/sig00000179 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000007d  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000177 ),
    .Q(\blk00000001/sig000000bb )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000007c  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000175 ),
    .Q(\blk00000001/sig000000bc )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000007b  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000173 ),
    .Q(\blk00000001/sig000000bd )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000007a  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000171 ),
    .Q(\blk00000001/sig000000be )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000079  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig0000016f ),
    .Q(\blk00000001/sig000000bf )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000078  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig0000016e ),
    .Q(\blk00000001/sig000000c0 )
  );
  MUXCY   \blk00000001/blk00000077  (
    .CI(\blk00000001/sig00000169 ),
    .DI(\blk00000001/sig0000051d ),
    .S(\blk00000001/sig00000567 ),
    .O(\blk00000001/sig00000178 )
  );
  XORCY   \blk00000001/blk00000076  (
    .CI(\blk00000001/sig00000169 ),
    .LI(\blk00000001/sig00000567 ),
    .O(\blk00000001/sig00000177 )
  );
  MUXCY   \blk00000001/blk00000075  (
    .CI(\blk00000001/sig00000178 ),
    .DI(\blk00000001/sig0000051d ),
    .S(\blk00000001/sig00000566 ),
    .O(\blk00000001/sig00000176 )
  );
  XORCY   \blk00000001/blk00000074  (
    .CI(\blk00000001/sig00000178 ),
    .LI(\blk00000001/sig00000566 ),
    .O(\blk00000001/sig00000175 )
  );
  MUXCY   \blk00000001/blk00000073  (
    .CI(\blk00000001/sig00000176 ),
    .DI(\blk00000001/sig0000051d ),
    .S(\blk00000001/sig00000565 ),
    .O(\blk00000001/sig00000174 )
  );
  XORCY   \blk00000001/blk00000072  (
    .CI(\blk00000001/sig00000176 ),
    .LI(\blk00000001/sig00000565 ),
    .O(\blk00000001/sig00000173 )
  );
  MUXCY   \blk00000001/blk00000071  (
    .CI(\blk00000001/sig00000174 ),
    .DI(\blk00000001/sig0000051d ),
    .S(\blk00000001/sig00000564 ),
    .O(\blk00000001/sig00000172 )
  );
  XORCY   \blk00000001/blk00000070  (
    .CI(\blk00000001/sig00000174 ),
    .LI(\blk00000001/sig00000564 ),
    .O(\blk00000001/sig00000171 )
  );
  MUXCY   \blk00000001/blk0000006f  (
    .CI(\blk00000001/sig00000172 ),
    .DI(\blk00000001/sig0000051d ),
    .S(\blk00000001/sig00000563 ),
    .O(\blk00000001/sig00000170 )
  );
  XORCY   \blk00000001/blk0000006e  (
    .CI(\blk00000001/sig00000172 ),
    .LI(\blk00000001/sig00000563 ),
    .O(\blk00000001/sig0000016f )
  );
  MUXCY   \blk00000001/blk0000006d  (
    .CI(\blk00000001/sig00000170 ),
    .DI(\blk00000001/sig0000051d ),
    .S(\blk00000001/sig00000562 ),
    .O(\blk00000001/sig00000168 )
  );
  XORCY   \blk00000001/blk0000006c  (
    .CI(\blk00000001/sig00000170 ),
    .LI(\blk00000001/sig00000562 ),
    .O(\blk00000001/sig0000016e )
  );
  MUXCY   \blk00000001/blk0000006b  (
    .CI(\blk00000001/sig0000003a ),
    .DI(\blk00000001/sig0000051d ),
    .S(\blk00000001/sig00000561 ),
    .O(\blk00000001/sig0000016d )
  );
  MUXCY   \blk00000001/blk0000006a  (
    .CI(\blk00000001/sig0000016d ),
    .DI(\blk00000001/sig0000051d ),
    .S(\blk00000001/sig0000051d ),
    .O(\blk00000001/sig0000016c )
  );
  MUXCY   \blk00000001/blk00000069  (
    .CI(\blk00000001/sig0000016c ),
    .DI(\blk00000001/sig0000003a ),
    .S(\blk00000001/sig0000016a ),
    .O(\blk00000001/sig00000169 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000068  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000140 ),
    .Q(\blk00000001/sig0000016b )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000067  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig0000013f ),
    .Q(\blk00000001/sig00000161 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000066  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig0000013e ),
    .Q(\blk00000001/sig00000162 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000065  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig0000013d ),
    .Q(\blk00000001/sig00000163 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000064  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig0000013c ),
    .Q(\blk00000001/sig00000164 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000063  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig0000013b ),
    .Q(\blk00000001/sig00000165 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000062  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig0000013a ),
    .Q(\blk00000001/sig00000166 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000061  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000139 ),
    .Q(\blk00000001/sig0000015b )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000060  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000138 ),
    .Q(\blk00000001/sig0000015c )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000005f  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000137 ),
    .Q(\blk00000001/sig0000015d )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000005e  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000136 ),
    .Q(\blk00000001/sig0000015e )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000005d  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000135 ),
    .Q(\blk00000001/sig0000015f )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000005c  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000134 ),
    .Q(\blk00000001/sig00000160 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000005b  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig0000014d ),
    .Q(\blk00000001/sig0000015a )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000005a  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig0000014c ),
    .Q(\blk00000001/sig00000159 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000059  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig0000014b ),
    .Q(\blk00000001/sig00000158 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000058  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig0000014a ),
    .Q(\blk00000001/sig00000157 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000057  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000149 ),
    .Q(\blk00000001/sig00000156 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000056  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000148 ),
    .Q(\blk00000001/sig00000155 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000055  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000147 ),
    .Q(\blk00000001/sig00000154 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000054  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000146 ),
    .Q(\blk00000001/sig00000153 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000053  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000145 ),
    .Q(\blk00000001/sig00000152 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000052  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000144 ),
    .Q(\blk00000001/sig00000151 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000051  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000143 ),
    .Q(\blk00000001/sig00000150 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000050  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000142 ),
    .Q(\blk00000001/sig0000014f )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000004f  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000141 ),
    .Q(\blk00000001/sig0000014e )
  );
  MUXF7   \blk00000001/blk0000004e  (
    .I0(\blk00000001/sig00000133 ),
    .I1(\blk00000001/sig00000132 ),
    .S(\blk00000001/sig000000cf ),
    .O(\NLW_blk00000001/blk0000004e_O_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000004d  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000000cd ),
    .Q(\blk00000001/sig000000c9 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000004c  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000000cc ),
    .Q(\blk00000001/sig000000c8 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000004b  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig0000012d ),
    .Q(\blk00000001/sig000000cc )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000004a  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig0000012c ),
    .Q(\blk00000001/sig000000cd )
  );
  MUXF7   \blk00000001/blk00000049  (
    .I0(\blk00000001/sig00000131 ),
    .I1(\blk00000001/sig0000012f ),
    .S(\blk00000001/sig000000cf ),
    .O(\blk00000001/sig0000012d )
  );
  MUXF7   \blk00000001/blk00000048  (
    .I0(\blk00000001/sig00000130 ),
    .I1(\blk00000001/sig0000012e ),
    .S(\blk00000001/sig000000cf ),
    .O(\blk00000001/sig0000012c )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000047  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000120 ),
    .Q(\blk00000001/sig000000c7 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000046  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig0000012b ),
    .Q(\blk00000001/sig00000127 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000045  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig0000012a ),
    .Q(\blk00000001/sig000000cf )
  );
  MUXCY   \blk00000001/blk00000044  (
    .CI(\blk00000001/sig0000003a ),
    .DI(\blk00000001/sig0000051d ),
    .S(\blk00000001/sig00000121 ),
    .O(\blk00000001/sig0000012b )
  );
  MUXCY   \blk00000001/blk00000043  (
    .CI(\blk00000001/sig0000012b ),
    .DI(\blk00000001/sig0000051d ),
    .S(\blk00000001/sig00000122 ),
    .O(\blk00000001/sig0000012a )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000042  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000129 ),
    .Q(\blk00000001/sig00000126 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000041  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000128 ),
    .Q(\blk00000001/sig00000125 )
  );
  MUXCY   \blk00000001/blk00000040  (
    .CI(\blk00000001/sig0000003a ),
    .DI(\blk00000001/sig0000051d ),
    .S(\blk00000001/sig00000123 ),
    .O(\blk00000001/sig00000129 )
  );
  MUXCY   \blk00000001/blk0000003f  (
    .CI(\blk00000001/sig00000129 ),
    .DI(\blk00000001/sig0000051d ),
    .S(\blk00000001/sig00000124 ),
    .O(\blk00000001/sig00000128 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000003e  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000000dd ),
    .Q(\blk00000001/sig000000d0 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000003d  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000000de ),
    .Q(\blk00000001/sig000000d1 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000003c  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000000df ),
    .Q(\blk00000001/sig000000d2 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000003b  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000000e0 ),
    .Q(\blk00000001/sig000000d3 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000003a  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000000e1 ),
    .Q(\blk00000001/sig000000d4 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000039  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000000e2 ),
    .Q(\blk00000001/sig000000d5 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000038  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000000e3 ),
    .Q(\blk00000001/sig000000d6 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000037  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000000e4 ),
    .Q(\blk00000001/sig000000d7 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000036  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000000e5 ),
    .Q(\blk00000001/sig000000d8 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000035  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000000e6 ),
    .Q(\blk00000001/sig000000d9 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000034  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000000e7 ),
    .Q(\blk00000001/sig000000da )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000033  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000000e8 ),
    .Q(\blk00000001/sig000000db )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000032  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000000e9 ),
    .Q(\blk00000001/sig000000dc )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000031  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig0000011e ),
    .Q(\blk00000001/sig000000dd )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000030  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig0000011c ),
    .Q(\blk00000001/sig000000de )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000002f  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig0000011a ),
    .Q(\blk00000001/sig000000df )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000002e  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000118 ),
    .Q(\blk00000001/sig000000e0 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000002d  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000116 ),
    .Q(\blk00000001/sig000000e1 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000002c  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000114 ),
    .Q(\blk00000001/sig000000e2 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000002b  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000112 ),
    .Q(\blk00000001/sig000000e3 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk0000002a  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000110 ),
    .Q(\blk00000001/sig000000e4 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000029  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig0000010e ),
    .Q(\blk00000001/sig000000e5 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000028  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig0000010c ),
    .Q(\blk00000001/sig000000e6 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000027  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig0000010a ),
    .Q(\blk00000001/sig000000e7 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000026  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000108 ),
    .Q(\blk00000001/sig000000e8 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000025  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000106 ),
    .Q(\blk00000001/sig000000e9 )
  );
  MUXCY   \blk00000001/blk00000024  (
    .CI(s_axis_divisor_tdata[12]),
    .DI(\blk00000001/sig0000051d ),
    .S(\blk00000001/sig000000ea ),
    .O(\blk00000001/sig0000011f )
  );
  XORCY   \blk00000001/blk00000023  (
    .CI(s_axis_divisor_tdata[12]),
    .LI(\blk00000001/sig000000ea ),
    .O(\blk00000001/sig0000011e )
  );
  MUXCY   \blk00000001/blk00000022  (
    .CI(\blk00000001/sig0000011f ),
    .DI(\blk00000001/sig0000051d ),
    .S(\blk00000001/sig000000eb ),
    .O(\blk00000001/sig0000011d )
  );
  XORCY   \blk00000001/blk00000021  (
    .CI(\blk00000001/sig0000011f ),
    .LI(\blk00000001/sig000000eb ),
    .O(\blk00000001/sig0000011c )
  );
  MUXCY   \blk00000001/blk00000020  (
    .CI(\blk00000001/sig0000011d ),
    .DI(\blk00000001/sig0000051d ),
    .S(\blk00000001/sig000000ec ),
    .O(\blk00000001/sig0000011b )
  );
  XORCY   \blk00000001/blk0000001f  (
    .CI(\blk00000001/sig0000011d ),
    .LI(\blk00000001/sig000000ec ),
    .O(\blk00000001/sig0000011a )
  );
  MUXCY   \blk00000001/blk0000001e  (
    .CI(\blk00000001/sig0000011b ),
    .DI(\blk00000001/sig0000051d ),
    .S(\blk00000001/sig000000ed ),
    .O(\blk00000001/sig00000119 )
  );
  XORCY   \blk00000001/blk0000001d  (
    .CI(\blk00000001/sig0000011b ),
    .LI(\blk00000001/sig000000ed ),
    .O(\blk00000001/sig00000118 )
  );
  MUXCY   \blk00000001/blk0000001c  (
    .CI(\blk00000001/sig00000119 ),
    .DI(\blk00000001/sig0000051d ),
    .S(\blk00000001/sig000000ee ),
    .O(\blk00000001/sig00000117 )
  );
  XORCY   \blk00000001/blk0000001b  (
    .CI(\blk00000001/sig00000119 ),
    .LI(\blk00000001/sig000000ee ),
    .O(\blk00000001/sig00000116 )
  );
  MUXCY   \blk00000001/blk0000001a  (
    .CI(\blk00000001/sig00000117 ),
    .DI(\blk00000001/sig0000051d ),
    .S(\blk00000001/sig000000ef ),
    .O(\blk00000001/sig00000115 )
  );
  XORCY   \blk00000001/blk00000019  (
    .CI(\blk00000001/sig00000117 ),
    .LI(\blk00000001/sig000000ef ),
    .O(\blk00000001/sig00000114 )
  );
  MUXCY   \blk00000001/blk00000018  (
    .CI(\blk00000001/sig00000115 ),
    .DI(\blk00000001/sig0000051d ),
    .S(\blk00000001/sig000000f0 ),
    .O(\blk00000001/sig00000113 )
  );
  XORCY   \blk00000001/blk00000017  (
    .CI(\blk00000001/sig00000115 ),
    .LI(\blk00000001/sig000000f0 ),
    .O(\blk00000001/sig00000112 )
  );
  MUXCY   \blk00000001/blk00000016  (
    .CI(\blk00000001/sig00000113 ),
    .DI(\blk00000001/sig0000051d ),
    .S(\blk00000001/sig000000f1 ),
    .O(\blk00000001/sig00000111 )
  );
  XORCY   \blk00000001/blk00000015  (
    .CI(\blk00000001/sig00000113 ),
    .LI(\blk00000001/sig000000f1 ),
    .O(\blk00000001/sig00000110 )
  );
  MUXCY   \blk00000001/blk00000014  (
    .CI(\blk00000001/sig00000111 ),
    .DI(\blk00000001/sig0000051d ),
    .S(\blk00000001/sig000000f2 ),
    .O(\blk00000001/sig0000010f )
  );
  XORCY   \blk00000001/blk00000013  (
    .CI(\blk00000001/sig00000111 ),
    .LI(\blk00000001/sig000000f2 ),
    .O(\blk00000001/sig0000010e )
  );
  MUXCY   \blk00000001/blk00000012  (
    .CI(\blk00000001/sig0000010f ),
    .DI(\blk00000001/sig0000051d ),
    .S(\blk00000001/sig000000f3 ),
    .O(\blk00000001/sig0000010d )
  );
  XORCY   \blk00000001/blk00000011  (
    .CI(\blk00000001/sig0000010f ),
    .LI(\blk00000001/sig000000f3 ),
    .O(\blk00000001/sig0000010c )
  );
  MUXCY   \blk00000001/blk00000010  (
    .CI(\blk00000001/sig0000010d ),
    .DI(\blk00000001/sig0000051d ),
    .S(\blk00000001/sig000000f4 ),
    .O(\blk00000001/sig0000010b )
  );
  XORCY   \blk00000001/blk0000000f  (
    .CI(\blk00000001/sig0000010d ),
    .LI(\blk00000001/sig000000f4 ),
    .O(\blk00000001/sig0000010a )
  );
  MUXCY   \blk00000001/blk0000000e  (
    .CI(\blk00000001/sig0000010b ),
    .DI(\blk00000001/sig0000051d ),
    .S(\blk00000001/sig000000f5 ),
    .O(\blk00000001/sig00000109 )
  );
  XORCY   \blk00000001/blk0000000d  (
    .CI(\blk00000001/sig0000010b ),
    .LI(\blk00000001/sig000000f5 ),
    .O(\blk00000001/sig00000108 )
  );
  MUXCY   \blk00000001/blk0000000c  (
    .CI(\blk00000001/sig00000109 ),
    .DI(\blk00000001/sig0000051d ),
    .S(\blk00000001/sig0000051d ),
    .O(\blk00000001/sig00000107 )
  );
  XORCY   \blk00000001/blk0000000b  (
    .CI(\blk00000001/sig00000109 ),
    .LI(\blk00000001/sig0000051d ),
    .O(\blk00000001/sig00000106 )
  );
  XORCY   \blk00000001/blk0000000a  (
    .CI(\blk00000001/sig00000107 ),
    .LI(\blk00000001/sig0000051d ),
    .O(\NLW_blk00000001/blk0000000a_O_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000009  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig000000c8 ),
    .Q(\blk00000001/sig000000fd )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000008  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000102 ),
    .Q(\blk00000001/sig000000fe )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000007  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000103 ),
    .Q(\blk00000001/sig000000ff )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000006  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000104 ),
    .Q(\blk00000001/sig00000100 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000005  (
    .C(aclk),
    .CE(\blk00000001/sig0000003a ),
    .D(\blk00000001/sig00000105 ),
    .Q(\blk00000001/sig00000101 )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk00000004  (
    .C(aclk),
    .D(\blk00000001/sig00000039 ),
    .Q(\blk00000001/sig0000003e )
  );
  GND   \blk00000001/blk00000003  (
    .G(\blk00000001/sig0000051d )
  );
  VCC   \blk00000001/blk00000002  (
    .P(\blk00000001/sig0000003a )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000000ae/blk000000c0  (
    .C(aclk),
    .D(\blk00000001/blk000000ae/sig000006b6 ),
    .Q(\blk00000001/sig0000006f )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000000ae/blk000000bf  (
    .C(aclk),
    .D(\blk00000001/blk000000ae/sig000006b7 ),
    .Q(\blk00000001/sig00000070 )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000000ae/blk000000be  (
    .C(aclk),
    .D(\blk00000001/blk000000ae/sig000006b8 ),
    .Q(\blk00000001/sig00000071 )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000000ae/blk000000bd  (
    .C(aclk),
    .D(\blk00000001/blk000000ae/sig000006b9 ),
    .Q(\blk00000001/sig00000072 )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000000ae/blk000000bc  (
    .C(aclk),
    .D(\blk00000001/blk000000ae/sig000006ba ),
    .Q(\blk00000001/sig00000073 )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000000ae/blk000000bb  (
    .C(aclk),
    .D(\blk00000001/blk000000ae/sig000006bb ),
    .Q(\blk00000001/sig00000074 )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000000ae/blk000000ba  (
    .C(aclk),
    .D(\blk00000001/blk000000ae/sig000006bc ),
    .Q(\blk00000001/sig00000075 )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000000ae/blk000000b9  (
    .C(aclk),
    .D(\blk00000001/blk000000ae/sig000006bd ),
    .Q(\blk00000001/sig00000076 )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000000ae/blk000000b8  (
    .C(aclk),
    .D(\blk00000001/blk000000ae/sig000006be ),
    .Q(\blk00000001/sig00000077 )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000000ae/blk000000b7  (
    .C(aclk),
    .D(\blk00000001/blk000000ae/sig000006bf ),
    .Q(\blk00000001/sig00000078 )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000000ae/blk000000b6  (
    .C(aclk),
    .D(\blk00000001/blk000000ae/sig000006c0 ),
    .Q(\blk00000001/sig00000079 )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000000ae/blk000000b5  (
    .C(aclk),
    .D(\blk00000001/blk000000ae/sig000006c1 ),
    .Q(\blk00000001/sig0000007a )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000000ae/blk000000b4  (
    .C(aclk),
    .D(\blk00000001/blk000000ae/sig000006c2 ),
    .Q(\blk00000001/sig0000007b )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk00000001/blk000000ae/blk000000b3  (
    .C(aclk),
    .D(\blk00000001/blk000000ae/sig000006c3 ),
    .Q(\blk00000001/sig0000007c )
  );
  DSP48A1 #(
    .A0REG ( 0 ),
    .A1REG ( 1 ),
    .B0REG ( 0 ),
    .B1REG ( 1 ),
    .CARRYINREG ( 0 ),
    .CARRYINSEL ( "OPMODE5" ),
    .CREG ( 0 ),
    .DREG ( 0 ),
    .MREG ( 1 ),
    .OPMODEREG ( 0 ),
    .PREG ( 0 ),
    .RSTTYPE ( "SYNC" ),
    .CARRYOUTREG ( 0 ))
  \blk00000001/blk000000ae/blk000000b2  (
    .CECARRYIN(\blk00000001/blk000000ae/sig000006d6 ),
    .RSTC(\blk00000001/blk000000ae/sig000006d6 ),
    .RSTCARRYIN(\blk00000001/blk000000ae/sig000006d6 ),
    .CED(\blk00000001/blk000000ae/sig000006d6 ),
    .RSTD(\blk00000001/blk000000ae/sig000006d6 ),
    .CEOPMODE(\blk00000001/blk000000ae/sig000006d6 ),
    .CEC(\blk00000001/blk000000ae/sig000006d6 ),
    .CARRYOUTF(\NLW_blk00000001/blk000000ae/blk000000b2_CARRYOUTF_UNCONNECTED ),
    .RSTOPMODE(\blk00000001/blk000000ae/sig000006d6 ),
    .RSTM(\blk00000001/blk000000ae/sig000006d6 ),
    .CLK(aclk),
    .RSTB(\blk00000001/blk000000ae/sig000006d6 ),
    .CEM(\blk00000001/blk000000ae/sig00000666 ),
    .CEB(\blk00000001/blk000000ae/sig00000666 ),
    .CARRYIN(\blk00000001/blk000000ae/sig000006d6 ),
    .CEP(\blk00000001/blk000000ae/sig000006d6 ),
    .CEA(\blk00000001/blk000000ae/sig00000666 ),
    .CARRYOUT(\NLW_blk00000001/blk000000ae/blk000000b2_CARRYOUT_UNCONNECTED ),
    .RSTA(\blk00000001/blk000000ae/sig000006d6 ),
    .RSTP(\blk00000001/blk000000ae/sig000006d6 ),
    .B({\blk00000001/blk000000ae/sig000006d6 , \blk00000001/blk000000ae/sig000006d6 , \blk00000001/blk000000ae/sig000006d6 ,
\blk00000001/blk000000ae/sig000006d6 , \blk00000001/sig0000051d , \blk00000001/sig00000089 , \blk00000001/sig00000088 , \blk00000001/sig00000087 ,
\blk00000001/sig00000086 , \blk00000001/sig00000085 , \blk00000001/sig00000084 , \blk00000001/sig00000083 , \blk00000001/sig00000082 ,
\blk00000001/sig00000081 , \blk00000001/sig00000080 , \blk00000001/sig0000007f , \blk00000001/sig0000007e , \blk00000001/sig0000007d }),
    .BCOUT({\blk00000001/blk000000ae/sig000006d5 , \blk00000001/blk000000ae/sig000006d4 , \blk00000001/blk000000ae/sig000006d3 ,
\blk00000001/blk000000ae/sig000006d2 , \blk00000001/blk000000ae/sig000006d1 , \blk00000001/blk000000ae/sig000006d0 ,
\blk00000001/blk000000ae/sig000006cf , \blk00000001/blk000000ae/sig000006ce , \blk00000001/blk000000ae/sig000006cd ,
\blk00000001/blk000000ae/sig000006cc , \blk00000001/blk000000ae/sig000006cb , \blk00000001/blk000000ae/sig000006ca ,
\blk00000001/blk000000ae/sig000006c9 , \blk00000001/blk000000ae/sig000006c8 , \blk00000001/blk000000ae/sig000006c7 ,
\blk00000001/blk000000ae/sig000006c6 , \blk00000001/blk000000ae/sig000006c5 , \blk00000001/blk000000ae/sig000006c4 }),
    .PCIN({\blk00000001/blk000000ae/sig000006d6 , \blk00000001/blk000000ae/sig000006d6 , \blk00000001/blk000000ae/sig000006d6 ,
\blk00000001/blk000000ae/sig000006d6 , \blk00000001/blk000000ae/sig000006d6 , \blk00000001/blk000000ae/sig000006d6 ,
\blk00000001/blk000000ae/sig000006d6 , \blk00000001/blk000000ae/sig000006d6 , \blk00000001/blk000000ae/sig000006d6 ,
\blk00000001/blk000000ae/sig000006d6 , \blk00000001/blk000000ae/sig000006d6 , \blk00000001/blk000000ae/sig000006d6 ,
\blk00000001/blk000000ae/sig000006d6 , \blk00000001/blk000000ae/sig000006d6 , \blk00000001/blk000000ae/sig000006d6 ,
\blk00000001/blk000000ae/sig000006d6 , \blk00000001/blk000000ae/sig000006d6 , \blk00000001/blk000000ae/sig000006d6 ,
\blk00000001/blk000000ae/sig000006d6 , \blk00000001/blk000000ae/sig000006d6 , \blk00000001/blk000000ae/sig000006d6 ,
\blk00000001/blk000000ae/sig000006d6 , \blk00000001/blk000000ae/sig000006d6 , \blk00000001/blk000000ae/sig000006d6 ,
\blk00000001/blk000000ae/sig000006d6 , \blk00000001/blk000000ae/sig000006d6 , \blk00000001/blk000000ae/sig000006d6 ,
\blk00000001/blk000000ae/sig000006d6 , \blk00000001/blk000000ae/sig000006d6 , \blk00000001/blk000000ae/sig000006d6 ,
\blk00000001/blk000000ae/sig000006d6 , \blk00000001/blk000000ae/sig000006d6 , \blk00000001/blk000000ae/sig000006d6 ,
\blk00000001/blk000000ae/sig000006d6 , \blk00000001/blk000000ae/sig000006d6 , \blk00000001/blk000000ae/sig000006d6 ,
\blk00000001/blk000000ae/sig000006d6 , \blk00000001/blk000000ae/sig000006d6 , \blk00000001/blk000000ae/sig000006d6 ,
\blk00000001/blk000000ae/sig000006d6 , \blk00000001/blk000000ae/sig000006d6 , \blk00000001/blk000000ae/sig000006d6 ,
\blk00000001/blk000000ae/sig000006d6 , \blk00000001/blk000000ae/sig000006d6 , \blk00000001/blk000000ae/sig000006d6 ,
\blk00000001/blk000000ae/sig000006d6 , \blk00000001/blk000000ae/sig000006d6 , \blk00000001/blk000000ae/sig000006d6 }),
    .C({\NLW_blk00000001/blk000000ae/blk000000b2_C<47>_UNCONNECTED , \NLW_blk00000001/blk000000ae/blk000000b2_C<46>_UNCONNECTED ,
\NLW_blk00000001/blk000000ae/blk000000b2_C<45>_UNCONNECTED , \NLW_blk00000001/blk000000ae/blk000000b2_C<44>_UNCONNECTED ,
\NLW_blk00000001/blk000000ae/blk000000b2_C<43>_UNCONNECTED , \NLW_blk00000001/blk000000ae/blk000000b2_C<42>_UNCONNECTED ,
\NLW_blk00000001/blk000000ae/blk000000b2_C<41>_UNCONNECTED , \NLW_blk00000001/blk000000ae/blk000000b2_C<40>_UNCONNECTED ,
\NLW_blk00000001/blk000000ae/blk000000b2_C<39>_UNCONNECTED , \NLW_blk00000001/blk000000ae/blk000000b2_C<38>_UNCONNECTED ,
\NLW_blk00000001/blk000000ae/blk000000b2_C<37>_UNCONNECTED , \NLW_blk00000001/blk000000ae/blk000000b2_C<36>_UNCONNECTED ,
\NLW_blk00000001/blk000000ae/blk000000b2_C<35>_UNCONNECTED , \NLW_blk00000001/blk000000ae/blk000000b2_C<34>_UNCONNECTED ,
\NLW_blk00000001/blk000000ae/blk000000b2_C<33>_UNCONNECTED , \NLW_blk00000001/blk000000ae/blk000000b2_C<32>_UNCONNECTED ,
\NLW_blk00000001/blk000000ae/blk000000b2_C<31>_UNCONNECTED , \NLW_blk00000001/blk000000ae/blk000000b2_C<30>_UNCONNECTED ,
\NLW_blk00000001/blk000000ae/blk000000b2_C<29>_UNCONNECTED , \NLW_blk00000001/blk000000ae/blk000000b2_C<28>_UNCONNECTED ,
\NLW_blk00000001/blk000000ae/blk000000b2_C<27>_UNCONNECTED , \NLW_blk00000001/blk000000ae/blk000000b2_C<26>_UNCONNECTED ,
\NLW_blk00000001/blk000000ae/blk000000b2_C<25>_UNCONNECTED , \NLW_blk00000001/blk000000ae/blk000000b2_C<24>_UNCONNECTED ,
\NLW_blk00000001/blk000000ae/blk000000b2_C<23>_UNCONNECTED , \NLW_blk00000001/blk000000ae/blk000000b2_C<22>_UNCONNECTED ,
\NLW_blk00000001/blk000000ae/blk000000b2_C<21>_UNCONNECTED , \NLW_blk00000001/blk000000ae/blk000000b2_C<20>_UNCONNECTED ,
\NLW_blk00000001/blk000000ae/blk000000b2_C<19>_UNCONNECTED , \NLW_blk00000001/blk000000ae/blk000000b2_C<18>_UNCONNECTED ,
\NLW_blk00000001/blk000000ae/blk000000b2_C<17>_UNCONNECTED , \NLW_blk00000001/blk000000ae/blk000000b2_C<16>_UNCONNECTED ,
\NLW_blk00000001/blk000000ae/blk000000b2_C<15>_UNCONNECTED , \NLW_blk00000001/blk000000ae/blk000000b2_C<14>_UNCONNECTED ,
\NLW_blk00000001/blk000000ae/blk000000b2_C<13>_UNCONNECTED , \NLW_blk00000001/blk000000ae/blk000000b2_C<12>_UNCONNECTED ,
\NLW_blk00000001/blk000000ae/blk000000b2_C<11>_UNCONNECTED , \NLW_blk00000001/blk000000ae/blk000000b2_C<10>_UNCONNECTED ,
\NLW_blk00000001/blk000000ae/blk000000b2_C<9>_UNCONNECTED , \NLW_blk00000001/blk000000ae/blk000000b2_C<8>_UNCONNECTED ,
\NLW_blk00000001/blk000000ae/blk000000b2_C<7>_UNCONNECTED , \NLW_blk00000001/blk000000ae/blk000000b2_C<6>_UNCONNECTED ,
\NLW_blk00000001/blk000000ae/blk000000b2_C<5>_UNCONNECTED , \NLW_blk00000001/blk000000ae/blk000000b2_C<4>_UNCONNECTED ,
\NLW_blk00000001/blk000000ae/blk000000b2_C<3>_UNCONNECTED , \NLW_blk00000001/blk000000ae/blk000000b2_C<2>_UNCONNECTED ,
\NLW_blk00000001/blk000000ae/blk000000b2_C<1>_UNCONNECTED , \NLW_blk00000001/blk000000ae/blk000000b2_C<0>_UNCONNECTED }),
    .P({\blk00000001/blk000000ae/sig000006b5 , \blk00000001/blk000000ae/sig000006b4 , \blk00000001/blk000000ae/sig000006b3 ,
\blk00000001/blk000000ae/sig000006b2 , \blk00000001/blk000000ae/sig000006b1 , \blk00000001/blk000000ae/sig000006b0 ,
\blk00000001/blk000000ae/sig000006af , \blk00000001/blk000000ae/sig000006ae , \blk00000001/blk000000ae/sig000006ad ,
\blk00000001/blk000000ae/sig000006ac , \blk00000001/blk000000ae/sig000006ab , \blk00000001/blk000000ae/sig000006aa ,
\blk00000001/blk000000ae/sig000006a9 , \blk00000001/blk000000ae/sig000006a8 , \blk00000001/blk000000ae/sig000006a7 ,
\blk00000001/blk000000ae/sig000006a6 , \blk00000001/blk000000ae/sig000006a5 , \blk00000001/blk000000ae/sig000006a4 ,
\blk00000001/blk000000ae/sig000006a3 , \blk00000001/blk000000ae/sig000006a2 , \blk00000001/blk000000ae/sig000006a1 ,
\blk00000001/blk000000ae/sig000006a0 , \blk00000001/blk000000ae/sig0000069f , \blk00000001/blk000000ae/sig0000069e ,
\blk00000001/blk000000ae/sig0000069d , \blk00000001/blk000000ae/sig0000069c , \blk00000001/blk000000ae/sig0000069b ,
\blk00000001/blk000000ae/sig0000069a , \blk00000001/blk000000ae/sig00000699 , \blk00000001/blk000000ae/sig00000698 ,
\blk00000001/blk000000ae/sig00000697 , \NLW_blk00000001/blk000000ae/blk000000b2_P<16>_UNCONNECTED ,
\NLW_blk00000001/blk000000ae/blk000000b2_P<15>_UNCONNECTED , \NLW_blk00000001/blk000000ae/blk000000b2_P<14>_UNCONNECTED ,
\blk00000001/blk000000ae/sig000006c3 , \blk00000001/blk000000ae/sig000006c2 , \blk00000001/blk000000ae/sig000006c1 ,
\blk00000001/blk000000ae/sig000006c0 , \blk00000001/blk000000ae/sig000006bf , \blk00000001/blk000000ae/sig000006be ,
\blk00000001/blk000000ae/sig000006bd , \blk00000001/blk000000ae/sig000006bc , \blk00000001/blk000000ae/sig000006bb ,
\blk00000001/blk000000ae/sig000006ba , \blk00000001/blk000000ae/sig000006b9 , \blk00000001/blk000000ae/sig000006b8 ,
\blk00000001/blk000000ae/sig000006b7 , \blk00000001/blk000000ae/sig000006b6 }),
    .OPMODE({\blk00000001/blk000000ae/sig000006d6 , \blk00000001/blk000000ae/sig000006d6 , \blk00000001/blk000000ae/sig000006d6 ,
\blk00000001/blk000000ae/sig000006d6 , \blk00000001/blk000000ae/sig000006d6 , \blk00000001/blk000000ae/sig000006d6 ,
\blk00000001/blk000000ae/sig000006d6 , \blk00000001/blk000000ae/sig00000666 }),
    .D({\blk00000001/blk000000ae/sig000006d6 , \blk00000001/blk000000ae/sig000006d6 , \blk00000001/blk000000ae/sig000006d6 ,
\blk00000001/blk000000ae/sig000006d6 , \blk00000001/blk000000ae/sig000006d6 , \blk00000001/blk000000ae/sig000006d6 ,
\blk00000001/blk000000ae/sig000006d6 , \blk00000001/blk000000ae/sig000006d6 , \blk00000001/blk000000ae/sig000006d6 ,
\blk00000001/blk000000ae/sig000006d6 , \blk00000001/blk000000ae/sig000006d6 , \blk00000001/blk000000ae/sig000006d6 ,
\blk00000001/blk000000ae/sig000006d6 , \blk00000001/blk000000ae/sig000006d6 , \blk00000001/blk000000ae/sig000006d6 ,
\blk00000001/blk000000ae/sig000006d6 , \blk00000001/blk000000ae/sig000006d6 , \blk00000001/blk000000ae/sig000006d6 }),
    .PCOUT({\blk00000001/blk000000ae/sig00000696 , \blk00000001/blk000000ae/sig00000695 , \blk00000001/blk000000ae/sig00000694 ,
\blk00000001/blk000000ae/sig00000693 , \blk00000001/blk000000ae/sig00000692 , \blk00000001/blk000000ae/sig00000691 ,
\blk00000001/blk000000ae/sig00000690 , \blk00000001/blk000000ae/sig0000068f , \blk00000001/blk000000ae/sig0000068e ,
\blk00000001/blk000000ae/sig0000068d , \blk00000001/blk000000ae/sig0000068c , \blk00000001/blk000000ae/sig0000068b ,
\blk00000001/blk000000ae/sig0000068a , \blk00000001/blk000000ae/sig00000689 , \blk00000001/blk000000ae/sig00000688 ,
\blk00000001/blk000000ae/sig00000687 , \blk00000001/blk000000ae/sig00000686 , \blk00000001/blk000000ae/sig00000685 ,
\blk00000001/blk000000ae/sig00000684 , \blk00000001/blk000000ae/sig00000683 , \blk00000001/blk000000ae/sig00000682 ,
\blk00000001/blk000000ae/sig00000681 , \blk00000001/blk000000ae/sig00000680 , \blk00000001/blk000000ae/sig0000067f ,
\blk00000001/blk000000ae/sig0000067e , \blk00000001/blk000000ae/sig0000067d , \blk00000001/blk000000ae/sig0000067c ,
\blk00000001/blk000000ae/sig0000067b , \blk00000001/blk000000ae/sig0000067a , \blk00000001/blk000000ae/sig00000679 ,
\blk00000001/blk000000ae/sig00000678 , \blk00000001/blk000000ae/sig00000677 , \blk00000001/blk000000ae/sig00000676 ,
\blk00000001/blk000000ae/sig00000675 , \blk00000001/blk000000ae/sig00000674 , \blk00000001/blk000000ae/sig00000673 ,
\blk00000001/blk000000ae/sig00000672 , \blk00000001/blk000000ae/sig00000671 , \blk00000001/blk000000ae/sig00000670 ,
\blk00000001/blk000000ae/sig0000066f , \blk00000001/blk000000ae/sig0000066e , \blk00000001/blk000000ae/sig0000066d ,
\blk00000001/blk000000ae/sig0000066c , \blk00000001/blk000000ae/sig0000066b , \blk00000001/blk000000ae/sig0000066a ,
\blk00000001/blk000000ae/sig00000669 , \blk00000001/blk000000ae/sig00000668 , \blk00000001/blk000000ae/sig00000667 }),
    .A({\blk00000001/blk000000ae/sig000006d6 , \blk00000001/sig0000009a , \blk00000001/sig00000099 , \blk00000001/sig00000098 ,
\blk00000001/sig00000097 , \blk00000001/sig00000096 , \blk00000001/sig00000095 , \blk00000001/sig00000094 , \blk00000001/sig00000093 ,
\blk00000001/sig00000092 , \blk00000001/sig00000091 , \blk00000001/sig00000090 , \blk00000001/sig0000008f , \blk00000001/sig0000008e ,
\blk00000001/sig0000008d , \blk00000001/sig0000008c , \blk00000001/sig0000008b , \blk00000001/sig0000008a }),
    .M({\NLW_blk00000001/blk000000ae/blk000000b2_M<35>_UNCONNECTED , \NLW_blk00000001/blk000000ae/blk000000b2_M<34>_UNCONNECTED ,
\NLW_blk00000001/blk000000ae/blk000000b2_M<33>_UNCONNECTED , \NLW_blk00000001/blk000000ae/blk000000b2_M<32>_UNCONNECTED ,
\NLW_blk00000001/blk000000ae/blk000000b2_M<31>_UNCONNECTED , \NLW_blk00000001/blk000000ae/blk000000b2_M<30>_UNCONNECTED ,
\NLW_blk00000001/blk000000ae/blk000000b2_M<29>_UNCONNECTED , \NLW_blk00000001/blk000000ae/blk000000b2_M<28>_UNCONNECTED ,
\NLW_blk00000001/blk000000ae/blk000000b2_M<27>_UNCONNECTED , \NLW_blk00000001/blk000000ae/blk000000b2_M<26>_UNCONNECTED ,
\NLW_blk00000001/blk000000ae/blk000000b2_M<25>_UNCONNECTED , \NLW_blk00000001/blk000000ae/blk000000b2_M<24>_UNCONNECTED ,
\NLW_blk00000001/blk000000ae/blk000000b2_M<23>_UNCONNECTED , \NLW_blk00000001/blk000000ae/blk000000b2_M<22>_UNCONNECTED ,
\NLW_blk00000001/blk000000ae/blk000000b2_M<21>_UNCONNECTED , \NLW_blk00000001/blk000000ae/blk000000b2_M<20>_UNCONNECTED ,
\NLW_blk00000001/blk000000ae/blk000000b2_M<19>_UNCONNECTED , \NLW_blk00000001/blk000000ae/blk000000b2_M<18>_UNCONNECTED ,
\NLW_blk00000001/blk000000ae/blk000000b2_M<17>_UNCONNECTED , \NLW_blk00000001/blk000000ae/blk000000b2_M<16>_UNCONNECTED ,
\NLW_blk00000001/blk000000ae/blk000000b2_M<15>_UNCONNECTED , \NLW_blk00000001/blk000000ae/blk000000b2_M<14>_UNCONNECTED ,
\NLW_blk00000001/blk000000ae/blk000000b2_M<13>_UNCONNECTED , \NLW_blk00000001/blk000000ae/blk000000b2_M<12>_UNCONNECTED ,
\NLW_blk00000001/blk000000ae/blk000000b2_M<11>_UNCONNECTED , \NLW_blk00000001/blk000000ae/blk000000b2_M<10>_UNCONNECTED ,
\NLW_blk00000001/blk000000ae/blk000000b2_M<9>_UNCONNECTED , \NLW_blk00000001/blk000000ae/blk000000b2_M<8>_UNCONNECTED ,
\NLW_blk00000001/blk000000ae/blk000000b2_M<7>_UNCONNECTED , \NLW_blk00000001/blk000000ae/blk000000b2_M<6>_UNCONNECTED ,
\NLW_blk00000001/blk000000ae/blk000000b2_M<5>_UNCONNECTED , \NLW_blk00000001/blk000000ae/blk000000b2_M<4>_UNCONNECTED ,
\NLW_blk00000001/blk000000ae/blk000000b2_M<3>_UNCONNECTED , \NLW_blk00000001/blk000000ae/blk000000b2_M<2>_UNCONNECTED ,
\NLW_blk00000001/blk000000ae/blk000000b2_M<1>_UNCONNECTED , \NLW_blk00000001/blk000000ae/blk000000b2_M<0>_UNCONNECTED })
  );
  DSP48A1 #(
    .A0REG ( 1 ),
    .A1REG ( 1 ),
    .B0REG ( 0 ),
    .B1REG ( 1 ),
    .CARRYINREG ( 0 ),
    .CARRYINSEL ( "OPMODE5" ),
    .CREG ( 0 ),
    .DREG ( 0 ),
    .MREG ( 0 ),
    .OPMODEREG ( 0 ),
    .PREG ( 1 ),
    .RSTTYPE ( "SYNC" ),
    .CARRYOUTREG ( 0 ))
  \blk00000001/blk000000ae/blk000000b1  (
    .CECARRYIN(\blk00000001/blk000000ae/sig000006d6 ),
    .RSTC(\blk00000001/blk000000ae/sig000006d6 ),
    .RSTCARRYIN(\blk00000001/blk000000ae/sig000006d6 ),
    .CED(\blk00000001/blk000000ae/sig000006d6 ),
    .RSTD(\blk00000001/blk000000ae/sig000006d6 ),
    .CEOPMODE(\blk00000001/blk000000ae/sig000006d6 ),
    .CEC(\blk00000001/blk000000ae/sig000006d6 ),
    .CARRYOUTF(\NLW_blk00000001/blk000000ae/blk000000b1_CARRYOUTF_UNCONNECTED ),
    .RSTOPMODE(\blk00000001/blk000000ae/sig000006d6 ),
    .RSTM(\blk00000001/blk000000ae/sig000006d6 ),
    .CLK(aclk),
    .RSTB(\blk00000001/blk000000ae/sig000006d6 ),
    .CEM(\blk00000001/blk000000ae/sig000006d6 ),
    .CEB(\blk00000001/blk000000ae/sig00000666 ),
    .CARRYIN(\blk00000001/blk000000ae/sig000006d6 ),
    .CEP(\blk00000001/blk000000ae/sig00000666 ),
    .CEA(\blk00000001/blk000000ae/sig00000666 ),
    .CARRYOUT(\NLW_blk00000001/blk000000ae/blk000000b1_CARRYOUT_UNCONNECTED ),
    .RSTA(\blk00000001/blk000000ae/sig000006d6 ),
    .RSTP(\blk00000001/blk000000ae/sig000006d6 ),
    .B({\blk00000001/blk000000ae/sig000006d5 , \blk00000001/blk000000ae/sig000006d4 , \blk00000001/blk000000ae/sig000006d3 ,
\blk00000001/blk000000ae/sig000006d2 , \blk00000001/blk000000ae/sig000006d1 , \blk00000001/blk000000ae/sig000006d0 ,
\blk00000001/blk000000ae/sig000006cf , \blk00000001/blk000000ae/sig000006ce , \blk00000001/blk000000ae/sig000006cd ,
\blk00000001/blk000000ae/sig000006cc , \blk00000001/blk000000ae/sig000006cb , \blk00000001/blk000000ae/sig000006ca ,
\blk00000001/blk000000ae/sig000006c9 , \blk00000001/blk000000ae/sig000006c8 , \blk00000001/blk000000ae/sig000006c7 ,
\blk00000001/blk000000ae/sig000006c6 , \blk00000001/blk000000ae/sig000006c5 , \blk00000001/blk000000ae/sig000006c4 }),
    .BCOUT({\NLW_blk00000001/blk000000ae/blk000000b1_BCOUT<17>_UNCONNECTED , \NLW_blk00000001/blk000000ae/blk000000b1_BCOUT<16>_UNCONNECTED ,
\NLW_blk00000001/blk000000ae/blk000000b1_BCOUT<15>_UNCONNECTED , \NLW_blk00000001/blk000000ae/blk000000b1_BCOUT<14>_UNCONNECTED ,
\NLW_blk00000001/blk000000ae/blk000000b1_BCOUT<13>_UNCONNECTED , \NLW_blk00000001/blk000000ae/blk000000b1_BCOUT<12>_UNCONNECTED ,
\NLW_blk00000001/blk000000ae/blk000000b1_BCOUT<11>_UNCONNECTED , \NLW_blk00000001/blk000000ae/blk000000b1_BCOUT<10>_UNCONNECTED ,
\NLW_blk00000001/blk000000ae/blk000000b1_BCOUT<9>_UNCONNECTED , \NLW_blk00000001/blk000000ae/blk000000b1_BCOUT<8>_UNCONNECTED ,
\NLW_blk00000001/blk000000ae/blk000000b1_BCOUT<7>_UNCONNECTED , \NLW_blk00000001/blk000000ae/blk000000b1_BCOUT<6>_UNCONNECTED ,
\NLW_blk00000001/blk000000ae/blk000000b1_BCOUT<5>_UNCONNECTED , \NLW_blk00000001/blk000000ae/blk000000b1_BCOUT<4>_UNCONNECTED ,
\NLW_blk00000001/blk000000ae/blk000000b1_BCOUT<3>_UNCONNECTED , \NLW_blk00000001/blk000000ae/blk000000b1_BCOUT<2>_UNCONNECTED ,
\NLW_blk00000001/blk000000ae/blk000000b1_BCOUT<1>_UNCONNECTED , \NLW_blk00000001/blk000000ae/blk000000b1_BCOUT<0>_UNCONNECTED }),
    .PCIN({\blk00000001/blk000000ae/sig00000696 , \blk00000001/blk000000ae/sig00000695 , \blk00000001/blk000000ae/sig00000694 ,
\blk00000001/blk000000ae/sig00000693 , \blk00000001/blk000000ae/sig00000692 , \blk00000001/blk000000ae/sig00000691 ,
\blk00000001/blk000000ae/sig00000690 , \blk00000001/blk000000ae/sig0000068f , \blk00000001/blk000000ae/sig0000068e ,
\blk00000001/blk000000ae/sig0000068d , \blk00000001/blk000000ae/sig0000068c , \blk00000001/blk000000ae/sig0000068b ,
\blk00000001/blk000000ae/sig0000068a , \blk00000001/blk000000ae/sig00000689 , \blk00000001/blk000000ae/sig00000688 ,
\blk00000001/blk000000ae/sig00000687 , \blk00000001/blk000000ae/sig00000686 , \blk00000001/blk000000ae/sig00000685 ,
\blk00000001/blk000000ae/sig00000684 , \blk00000001/blk000000ae/sig00000683 , \blk00000001/blk000000ae/sig00000682 ,
\blk00000001/blk000000ae/sig00000681 , \blk00000001/blk000000ae/sig00000680 , \blk00000001/blk000000ae/sig0000067f ,
\blk00000001/blk000000ae/sig0000067e , \blk00000001/blk000000ae/sig0000067d , \blk00000001/blk000000ae/sig0000067c ,
\blk00000001/blk000000ae/sig0000067b , \blk00000001/blk000000ae/sig0000067a , \blk00000001/blk000000ae/sig00000679 ,
\blk00000001/blk000000ae/sig00000678 , \blk00000001/blk000000ae/sig00000677 , \blk00000001/blk000000ae/sig00000676 ,
\blk00000001/blk000000ae/sig00000675 , \blk00000001/blk000000ae/sig00000674 , \blk00000001/blk000000ae/sig00000673 ,
\blk00000001/blk000000ae/sig00000672 , \blk00000001/blk000000ae/sig00000671 , \blk00000001/blk000000ae/sig00000670 ,
\blk00000001/blk000000ae/sig0000066f , \blk00000001/blk000000ae/sig0000066e , \blk00000001/blk000000ae/sig0000066d ,
\blk00000001/blk000000ae/sig0000066c , \blk00000001/blk000000ae/sig0000066b , \blk00000001/blk000000ae/sig0000066a ,
\blk00000001/blk000000ae/sig00000669 , \blk00000001/blk000000ae/sig00000668 , \blk00000001/blk000000ae/sig00000667 }),
    .C({\blk00000001/blk000000ae/sig000006b5 , \blk00000001/blk000000ae/sig000006b5 , \blk00000001/blk000000ae/sig000006b5 ,
\blk00000001/blk000000ae/sig000006b5 , \blk00000001/blk000000ae/sig000006b5 , \blk00000001/blk000000ae/sig000006b5 ,
\blk00000001/blk000000ae/sig000006b5 , \blk00000001/blk000000ae/sig000006b5 , \blk00000001/blk000000ae/sig000006b5 ,
\blk00000001/blk000000ae/sig000006b5 , \blk00000001/blk000000ae/sig000006b5 , \blk00000001/blk000000ae/sig000006b5 ,
\blk00000001/blk000000ae/sig000006b5 , \blk00000001/blk000000ae/sig000006b5 , \blk00000001/blk000000ae/sig000006b5 ,
\blk00000001/blk000000ae/sig000006b5 , \blk00000001/blk000000ae/sig000006b5 , \blk00000001/blk000000ae/sig000006b5 ,
\blk00000001/blk000000ae/sig000006b4 , \blk00000001/blk000000ae/sig000006b3 , \blk00000001/blk000000ae/sig000006b2 ,
\blk00000001/blk000000ae/sig000006b1 , \blk00000001/blk000000ae/sig000006b0 , \blk00000001/blk000000ae/sig000006af ,
\blk00000001/blk000000ae/sig000006ae , \blk00000001/blk000000ae/sig000006ad , \blk00000001/blk000000ae/sig000006ac ,
\blk00000001/blk000000ae/sig000006ab , \blk00000001/blk000000ae/sig000006aa , \blk00000001/blk000000ae/sig000006a9 ,
\blk00000001/blk000000ae/sig000006a8 , \blk00000001/blk000000ae/sig000006a7 , \blk00000001/blk000000ae/sig000006a6 ,
\blk00000001/blk000000ae/sig000006a5 , \blk00000001/blk000000ae/sig000006a4 , \blk00000001/blk000000ae/sig000006a3 ,
\blk00000001/blk000000ae/sig000006a2 , \blk00000001/blk000000ae/sig000006a1 , \blk00000001/blk000000ae/sig000006a0 ,
\blk00000001/blk000000ae/sig0000069f , \blk00000001/blk000000ae/sig0000069e , \blk00000001/blk000000ae/sig0000069d ,
\blk00000001/blk000000ae/sig0000069c , \blk00000001/blk000000ae/sig0000069b , \blk00000001/blk000000ae/sig0000069a ,
\blk00000001/blk000000ae/sig00000699 , \blk00000001/blk000000ae/sig00000698 , \blk00000001/blk000000ae/sig00000697 }),
    .P({\NLW_blk00000001/blk000000ae/blk000000b1_P<47>_UNCONNECTED , \NLW_blk00000001/blk000000ae/blk000000b1_P<46>_UNCONNECTED ,
\NLW_blk00000001/blk000000ae/blk000000b1_P<45>_UNCONNECTED , \NLW_blk00000001/blk000000ae/blk000000b1_P<44>_UNCONNECTED ,
\NLW_blk00000001/blk000000ae/blk000000b1_P<43>_UNCONNECTED , \NLW_blk00000001/blk000000ae/blk000000b1_P<42>_UNCONNECTED ,
\NLW_blk00000001/blk000000ae/blk000000b1_P<41>_UNCONNECTED , \NLW_blk00000001/blk000000ae/blk000000b1_P<40>_UNCONNECTED ,
\NLW_blk00000001/blk000000ae/blk000000b1_P<39>_UNCONNECTED , \NLW_blk00000001/blk000000ae/blk000000b1_P<38>_UNCONNECTED ,
\NLW_blk00000001/blk000000ae/blk000000b1_P<37>_UNCONNECTED , \NLW_blk00000001/blk000000ae/blk000000b1_P<36>_UNCONNECTED ,
\NLW_blk00000001/blk000000ae/blk000000b1_P<35>_UNCONNECTED , \NLW_blk00000001/blk000000ae/blk000000b1_P<34>_UNCONNECTED ,
\NLW_blk00000001/blk000000ae/blk000000b1_P<33>_UNCONNECTED , \NLW_blk00000001/blk000000ae/blk000000b1_P<32>_UNCONNECTED ,
\NLW_blk00000001/blk000000ae/blk000000b1_P<31>_UNCONNECTED , \NLW_blk00000001/blk000000ae/blk000000b1_P<30>_UNCONNECTED ,
\NLW_blk00000001/blk000000ae/blk000000b1_P<29>_UNCONNECTED , \NLW_blk00000001/blk000000ae/blk000000b1_P<28>_UNCONNECTED ,
\NLW_blk00000001/blk000000ae/blk000000b1_P<27>_UNCONNECTED , \NLW_blk00000001/blk000000ae/blk000000b1_P<26>_UNCONNECTED ,
\NLW_blk00000001/blk000000ae/blk000000b1_P<25>_UNCONNECTED , \NLW_blk00000001/blk000000ae/blk000000b1_P<24>_UNCONNECTED ,
\NLW_blk00000001/blk000000ae/blk000000b1_P<23>_UNCONNECTED , \NLW_blk00000001/blk000000ae/blk000000b1_P<22>_UNCONNECTED ,
\NLW_blk00000001/blk000000ae/blk000000b1_P<21>_UNCONNECTED , \NLW_blk00000001/blk000000ae/blk000000b1_P<20>_UNCONNECTED ,
\NLW_blk00000001/blk000000ae/blk000000b1_P<19>_UNCONNECTED , \NLW_blk00000001/blk000000ae/blk000000b1_P<18>_UNCONNECTED ,
\NLW_blk00000001/blk000000ae/blk000000b1_P<17>_UNCONNECTED , \NLW_blk00000001/blk000000ae/blk000000b1_P<16>_UNCONNECTED ,
\blk00000001/blk000000ae/sig00000618 , \blk00000001/blk000000ae/sig00000619 , \blk00000001/blk000000ae/sig0000061a ,
\blk00000001/blk000000ae/sig0000061b , \blk00000001/blk000000ae/sig0000061c , \blk00000001/blk000000ae/sig0000061d ,
\blk00000001/blk000000ae/sig0000061e , \blk00000001/blk000000ae/sig0000061f , \blk00000001/blk000000ae/sig00000620 ,
\blk00000001/blk000000ae/sig00000621 , \blk00000001/blk000000ae/sig00000622 , \blk00000001/blk000000ae/sig00000623 ,
\blk00000001/blk000000ae/sig00000624 , \blk00000001/blk000000ae/sig00000625 , \blk00000001/blk000000ae/sig00000626 ,
\blk00000001/blk000000ae/sig00000627 }),
    .OPMODE({\blk00000001/blk000000ae/sig000006d6 , \blk00000001/blk000000ae/sig000006d6 , \blk00000001/blk000000ae/sig000006d6 ,
\blk00000001/blk000000ae/sig000006d6 , \blk00000001/blk000000ae/sig00000666 , \blk00000001/blk000000ae/sig00000666 ,
\blk00000001/blk000000ae/sig000006d6 , \blk00000001/blk000000ae/sig00000666 }),
    .D({\blk00000001/blk000000ae/sig000006d6 , \blk00000001/blk000000ae/sig000006d6 , \blk00000001/blk000000ae/sig000006d6 ,
\blk00000001/blk000000ae/sig000006d6 , \blk00000001/blk000000ae/sig000006d6 , \blk00000001/blk000000ae/sig000006d6 ,
\blk00000001/blk000000ae/sig000006d6 , \blk00000001/blk000000ae/sig000006d6 , \blk00000001/blk000000ae/sig000006d6 ,
\blk00000001/blk000000ae/sig000006d6 , \blk00000001/blk000000ae/sig000006d6 , \blk00000001/blk000000ae/sig000006d6 ,
\blk00000001/blk000000ae/sig000006d6 , \blk00000001/blk000000ae/sig000006d6 , \blk00000001/blk000000ae/sig000006d6 ,
\blk00000001/blk000000ae/sig000006d6 , \blk00000001/blk000000ae/sig000006d6 , \blk00000001/blk000000ae/sig000006d6 }),
    .PCOUT({\blk00000001/blk000000ae/sig00000636 , \blk00000001/blk000000ae/sig00000637 , \blk00000001/blk000000ae/sig00000638 ,
\blk00000001/blk000000ae/sig00000639 , \blk00000001/blk000000ae/sig0000063a , \blk00000001/blk000000ae/sig0000063b ,
\blk00000001/blk000000ae/sig0000063c , \blk00000001/blk000000ae/sig0000063d , \blk00000001/blk000000ae/sig0000063e ,
\blk00000001/blk000000ae/sig0000063f , \blk00000001/blk000000ae/sig00000640 , \blk00000001/blk000000ae/sig00000641 ,
\blk00000001/blk000000ae/sig00000642 , \blk00000001/blk000000ae/sig00000643 , \blk00000001/blk000000ae/sig00000644 ,
\blk00000001/blk000000ae/sig00000645 , \blk00000001/blk000000ae/sig00000646 , \blk00000001/blk000000ae/sig00000647 ,
\blk00000001/blk000000ae/sig00000648 , \blk00000001/blk000000ae/sig00000649 , \blk00000001/blk000000ae/sig0000064a ,
\blk00000001/blk000000ae/sig0000064b , \blk00000001/blk000000ae/sig0000064c , \blk00000001/blk000000ae/sig0000064d ,
\blk00000001/blk000000ae/sig0000064e , \blk00000001/blk000000ae/sig0000064f , \blk00000001/blk000000ae/sig00000650 ,
\blk00000001/blk000000ae/sig00000651 , \blk00000001/blk000000ae/sig00000652 , \blk00000001/blk000000ae/sig00000653 ,
\blk00000001/blk000000ae/sig00000654 , \blk00000001/blk000000ae/sig00000655 , \blk00000001/blk000000ae/sig00000656 ,
\blk00000001/blk000000ae/sig00000657 , \blk00000001/blk000000ae/sig00000658 , \blk00000001/blk000000ae/sig00000659 ,
\blk00000001/blk000000ae/sig0000065a , \blk00000001/blk000000ae/sig0000065b , \blk00000001/blk000000ae/sig0000065c ,
\blk00000001/blk000000ae/sig0000065d , \blk00000001/blk000000ae/sig0000065e , \blk00000001/blk000000ae/sig0000065f ,
\blk00000001/blk000000ae/sig00000660 , \blk00000001/blk000000ae/sig00000661 , \blk00000001/blk000000ae/sig00000662 ,
\blk00000001/blk000000ae/sig00000663 , \blk00000001/blk000000ae/sig00000664 , \blk00000001/blk000000ae/sig00000665 }),
    .A({\blk00000001/sig0000009c , \blk00000001/sig0000009c , \blk00000001/sig0000009c , \blk00000001/sig0000009c , \blk00000001/sig0000009c ,
\blk00000001/sig0000009c , \blk00000001/sig0000009c , \blk00000001/sig0000009c , \blk00000001/sig0000009c , \blk00000001/sig0000009c ,
\blk00000001/sig0000009c , \blk00000001/sig0000009c , \blk00000001/sig0000009c , \blk00000001/sig0000009c , \blk00000001/sig0000009c ,
\blk00000001/sig0000009c , \blk00000001/sig0000009c , \blk00000001/sig0000009b }),
    .M({\NLW_blk00000001/blk000000ae/blk000000b1_M<35>_UNCONNECTED , \NLW_blk00000001/blk000000ae/blk000000b1_M<34>_UNCONNECTED ,
\NLW_blk00000001/blk000000ae/blk000000b1_M<33>_UNCONNECTED , \NLW_blk00000001/blk000000ae/blk000000b1_M<32>_UNCONNECTED ,
\NLW_blk00000001/blk000000ae/blk000000b1_M<31>_UNCONNECTED , \NLW_blk00000001/blk000000ae/blk000000b1_M<30>_UNCONNECTED ,
\NLW_blk00000001/blk000000ae/blk000000b1_M<29>_UNCONNECTED , \NLW_blk00000001/blk000000ae/blk000000b1_M<28>_UNCONNECTED ,
\NLW_blk00000001/blk000000ae/blk000000b1_M<27>_UNCONNECTED , \NLW_blk00000001/blk000000ae/blk000000b1_M<26>_UNCONNECTED ,
\NLW_blk00000001/blk000000ae/blk000000b1_M<25>_UNCONNECTED , \NLW_blk00000001/blk000000ae/blk000000b1_M<24>_UNCONNECTED ,
\NLW_blk00000001/blk000000ae/blk000000b1_M<23>_UNCONNECTED , \NLW_blk00000001/blk000000ae/blk000000b1_M<22>_UNCONNECTED ,
\NLW_blk00000001/blk000000ae/blk000000b1_M<21>_UNCONNECTED , \NLW_blk00000001/blk000000ae/blk000000b1_M<20>_UNCONNECTED ,
\NLW_blk00000001/blk000000ae/blk000000b1_M<19>_UNCONNECTED , \NLW_blk00000001/blk000000ae/blk000000b1_M<18>_UNCONNECTED ,
\NLW_blk00000001/blk000000ae/blk000000b1_M<17>_UNCONNECTED , \NLW_blk00000001/blk000000ae/blk000000b1_M<16>_UNCONNECTED ,
\NLW_blk00000001/blk000000ae/blk000000b1_M<15>_UNCONNECTED , \NLW_blk00000001/blk000000ae/blk000000b1_M<14>_UNCONNECTED ,
\NLW_blk00000001/blk000000ae/blk000000b1_M<13>_UNCONNECTED , \NLW_blk00000001/blk000000ae/blk000000b1_M<12>_UNCONNECTED ,
\NLW_blk00000001/blk000000ae/blk000000b1_M<11>_UNCONNECTED , \NLW_blk00000001/blk000000ae/blk000000b1_M<10>_UNCONNECTED ,
\NLW_blk00000001/blk000000ae/blk000000b1_M<9>_UNCONNECTED , \NLW_blk00000001/blk000000ae/blk000000b1_M<8>_UNCONNECTED ,
\NLW_blk00000001/blk000000ae/blk000000b1_M<7>_UNCONNECTED , \NLW_blk00000001/blk000000ae/blk000000b1_M<6>_UNCONNECTED ,
\NLW_blk00000001/blk000000ae/blk000000b1_M<5>_UNCONNECTED , \NLW_blk00000001/blk000000ae/blk000000b1_M<4>_UNCONNECTED ,
\NLW_blk00000001/blk000000ae/blk000000b1_M<3>_UNCONNECTED , \NLW_blk00000001/blk000000ae/blk000000b1_M<2>_UNCONNECTED ,
\NLW_blk00000001/blk000000ae/blk000000b1_M<1>_UNCONNECTED , \NLW_blk00000001/blk000000ae/blk000000b1_M<0>_UNCONNECTED })
  );
  GND   \blk00000001/blk000000ae/blk000000b0  (
    .G(\blk00000001/blk000000ae/sig000006d6 )
  );
  VCC   \blk00000001/blk000000ae/blk000000af  (
    .P(\blk00000001/blk000000ae/sig00000666 )
  );
// synthesis translate_on
endmodule