module ADC_SAR_v3_0_0 (
    vplus,
    vminus,
    soc,
    eoc,
    aclk,
    vdac_ref,
    eos);
    inout       vplus;
    electrical  vplus;
    inout       vminus;
    electrical  vminus;
    input       soc;
    output      eoc;
    input       aclk;
    inout       vdac_ref;
    electrical  vdac_ref;
    output      eos;
          wire [3:0] vp_ctl;
          wire [3:0] vn_ctl;
          wire  Net_381;
    electrical  Net_255;
    electrical  Net_267;
    electrical  Net_210;
    electrical  Net_209;
          wire [11:0] Net_207;
          wire  Net_252;
          wire  Net_205;
          wire  Net_378;
          wire  Net_376;
    electrical  Net_368;
    electrical  Net_235;
    electrical  Net_216;
    electrical  Net_233;
          wire  Net_221;
    electrical  Net_248;
    electrical  Net_257;
    electrical  Net_149;
    electrical  Net_126;
    electrical  Net_215;
          wire  Net_188;
	// cy_analog_virtualmux_3 (cy_analog_virtualmux_v1_0)
	cy_connect_v1_0 cy_analog_virtualmux_3_connect(Net_248, Net_235);
	defparam cy_analog_virtualmux_3_connect.sig_width = 1;
    ZeroTerminal ZeroTerminal_1 (
        .z(vp_ctl[0]));
    ZeroTerminal ZeroTerminal_2 (
        .z(vp_ctl[2]));
    ZeroTerminal ZeroTerminal_3 (
        .z(vn_ctl[1]));
    ZeroTerminal ZeroTerminal_4 (
        .z(vn_ctl[3]));
    ZeroTerminal ZeroTerminal_5 (
        .z(vp_ctl[1]));
    ZeroTerminal ZeroTerminal_6 (
        .z(vp_ctl[3]));
    ZeroTerminal ZeroTerminal_7 (
        .z(vn_ctl[0]));
    ZeroTerminal ZeroTerminal_8 (
        .z(vn_ctl[2]));
	// Clock_VirtualMux_1 (cy_virtualmux_v1_0)
	assign Net_188 = aclk;
    cy_psoc5_sar_v2_0 ADC_SAR (
        .clock(Net_188),
        .sof_udb(soc),
        .clk_udb(),
        .vp_ctl_udb(vp_ctl[3:0]),
        .vn_ctl_udb(vn_ctl[3:0]),
        .vplus(vplus),
        .vminus(Net_126),
        .irq(Net_252),
        .data_out(Net_207[11:0]),
        .eof_udb(eoc),
        .pump_clock(Net_188),
        .ext_pin(Net_215),
        .vrefhi_out(Net_257),
        .vref(Net_248),
        .next_out(eos));
	// cy_analog_virtualmux_2 (cy_analog_virtualmux_v1_0)
	cy_connect_v1_0 cy_analog_virtualmux_2_connect(Net_215, Net_209);
	defparam cy_analog_virtualmux_2_connect.sig_width = 1;
	// cy_analog_virtualmux_1 (cy_analog_virtualmux_v1_0)
	cy_connect_v1_0 cy_analog_virtualmux_1_connect(Net_126, Net_149);
	defparam cy_analog_virtualmux_1_connect.sig_width = 1;
    cy_analog_noconnect_v1_0 noconnect (
        .noconnect(Net_209));
	// cy_analog_virtualmux_4 (cy_analog_virtualmux_v1_0)
	cy_connect_v1_0 cy_analog_virtualmux_4_connect(Net_257, Net_149);
	defparam cy_analog_virtualmux_4_connect.sig_width = 1;
    cy_analog_noconnect_v1_0 cy_analog_noconnect_1 (
        .noconnect(Net_255));
	cy_vref_v1_0
		#(.autoenable(1),
		  .guid("4720866E-BC14-478d-B8A0-3E44F38CADAC"),
		  .name("Vdda/2"))
		vRef_Vdda_1
		 (.vout(Net_235));
    cy_analog_noconnect_v1_0 noconnect_1 (
        .noconnect(Net_368));
    assign Net_221 = Net_376 | Net_381;
    assign Net_381 = 1'h0;
endmodule