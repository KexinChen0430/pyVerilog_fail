module header
	// Internal signals
	// Generated Signal List
		wire		sig_01; // __W_PORT_SIGNAL_MAP_REQ
		wire	[4:0]	sig_02;
		wire		sig_03; // __W_PORT_SIGNAL_MAP_REQ
		wire		sig_04; // __W_PORT_SIGNAL_MAP_REQ
		wire	[3:0]	sig_05; // __W_PORT_SIGNAL_MAP_REQ
		wire	[3:0]	sig_06; // __W_PORT_SIGNAL_MAP_REQ
		wire	[6:0]	sig_14;
		wire	[6:0]	sig_i_ae; // __W_PORT_SIGNAL_MAP_REQ
		wire	[7:0]	sig_o_ae; // __W_PORT_SIGNAL_MAP_REQ
	// End of Generated Signal List
	// %COMPILER_OPTS%
	// Generated Signal Assignments
		assign	p_mix_sig_01_go	=	sig_01;  // __I_O_BIT_PORT
		assign	p_mix_sig_03_go	=	sig_03;  // __I_O_BIT_PORT
		assign	sig_04	=	p_mix_sig_04_gi;  // __I_I_BIT_PORT
		assign	p_mix_sig_05_2_1_go[1:0]	=	sig_05[2:1];  // __I_O_SLICE_PORT
		assign	sig_06	=	p_mix_sig_06_gi;  // __I_I_BUS_PORT
		assign	sig_i_ae	=	p_mix_sig_i_ae_gi;  // __I_I_BUS_PORT
		assign	p_mix_sig_o_ae_go	=	sig_o_ae;  // __I_O_BUS_PORT
	// Generated Instances and Port Mappings
	`ifdef insert_emu_mux_inst_aa
		// Emulator Data Injection Path, generated by MIX
		wire emu_mux_inst_aa = 1'b0;
		wire		sig_04_emux_s;
		wire		sig_04_vc_s;
		assign sig_04_emux_s	= emu_mux_inst_aa ? sig_04_vc_s	: sig_04;
	`endif
		// Generated Instance Port Map for inst_aa
		ent_aa inst_aa (
			.port_aa_1(sig_01),	// Use internally test1Will create p_mix_sig_1_go port
			.port_aa_2(sig_02[0]),	// Use internally test2, no port generated
			.port_aa_3(sig_03),	// Interhierachy link, will create p_mix_sig_3_go
		`ifdef insert_emu_mux_inst_aa
			.port_aa_4(sig_04_emux_s),
		`else
			.port_aa_4(sig_04),	// Interhierachy link, will create p_mix_sig_4_gi
		`endif
			.port_aa_5(sig_05),	// Bus, single bits go to outsideBus, single bits go to outside, will create p_mix_sig_5_2_2_goBu...
			.port_aa_6(sig_06),	// Conflicting definition (X2)
			.sig_07(sig_07),	// Conflicting definition, IN false!
			.sig_08(sig_08),	// VHDL intermediate needed (port name)
			.sig_13(sig_13),	// Create internal signal name
			.sig_14(sig_14)	// Multiline comment 1
		);
		// End of Generated Instance Port Map for inst_aa
	`ifdef insert_emu_mux_inst_ab
		// Emulator Data Injection Path, generated by MIX
		wire emu_mux_inst_ab = 1'b0;
		wire		sig_01_emux_s;
		wire		sig_01_vc_s;
		wire	[4:0]	sig_13_emux_s;
		wire	[4:0]	sig_13_vc_s;
		wire	[6:0]	sig_14_emux_s;
		wire	[6:0]	sig_14_vc_s;
		assign sig_01_emux_s	= emu_mux_inst_ab ? sig_01_vc_s	: sig_01;
		assign sig_13_emux_s	= emu_mux_inst_ab ? sig_13_vc_s	: sig_13;
		assign sig_14_emux_s	= emu_mux_inst_ab ? sig_14_vc_s	: sig_14;
	`endif
		// Generated Instance Port Map for inst_ab
		ent_ab inst_ab (
		`ifdef insert_emu_mux_inst_ab
			.port_ab_1(sig_01_emux_s),
		`else
			.port_ab_1(sig_01),	// Use internally test1Will create p_mix_sig_1_go port
		`endif
			.port_ab_2(sig_02[1]),	// Use internally test2, no port generated
		`ifdef insert_emu_mux_inst_ab
			.sig_13(sig_13_emux_s),
		`else
			.sig_13(sig_13),	// Create internal signal name
		`endif
		`ifdef insert_emu_mux_inst_ab
			.sig_14(sig_14_emux_s)
		`else
			.sig_14(sig_14)	// Multiline comment 1
		`endif
		);
		// End of Generated Instance Port Map for inst_ab
	`ifdef insert_emu_mux_inst_ac
		// Emulator Data Injection Path, generated by MIX
		wire emu_mux_inst_ac = 1'b0;
		wire		sig_02_3_emux_s;
		wire		sig_02_3_vc_s;
		assign sig_02[3]	= emu_mux_inst_ac ? sig_02_3_vc_s	: sig_02_3_emux_s;
	`endif
		// Generated Instance Port Map for inst_ac
		ent_ac inst_ac (
		`ifdef insert_emu_mux_inst_ac
			.port_ac_2(sig_02_3_emux_s)
		`else
			.port_ac_2(sig_02[3])	// Use internally test2, no port generated
		`endif
		);
		// End of Generated Instance Port Map for inst_ac
	`ifdef insert_emu_mux_inst_ad
		// Emulator Data Injection Path, generated by MIX
		wire emu_mux_inst_ad = 1'b0;
		wire		sig_02_4_emux_s;
		wire		sig_02_4_vc_s;
		assign sig_02[4]	= emu_mux_inst_ad ? sig_02_4_vc_s	: sig_02_4_emux_s;
	`endif
		// Generated Instance Port Map for inst_ad
		ent_ad inst_ad (
		`ifdef insert_emu_mux_inst_ad
			.port_ad_2(sig_02_4_emux_s)
		`else
			.port_ad_2(sig_02[4])	// Use internally test2, no port generated
		`endif
		);
		// End of Generated Instance Port Map for inst_ad
	`ifdef insert_emu_mux_inst_ae
		// Emulator Data Injection Path, generated by MIX
		wire emu_mux_inst_ae = 1'b0;
		wire	[1:0]	sig_02_1_0_emux_s;
		wire	[1:0]	sig_02_1_0_vc_s;
		wire	[4:3]	sig_02_4_3_emux_s;
		wire	[4:3]	sig_02_4_3_vc_s;
		wire	[3:0]	sig_05_emux_s;
		wire	[3:0]	sig_05_vc_s;
		wire	[3:0]	sig_06_emux_s;
		wire	[3:0]	sig_06_vc_s;
		wire	[5:0]	sig_07_emux_s;
		wire	[5:0]	sig_07_vc_s;
		wire	[8:2]	sig_08_emux_s;
		wire	[8:2]	sig_08_vc_s;
		wire	[6:0]	sig_i_ae_emux_s;
		wire	[6:0]	sig_i_ae_vc_s;
		assign sig_02_1_0_emux_s	= emu_mux_inst_ae ? sig_02_1_0_vc_s	: sig_02[1:0];
		assign sig_02_4_3_emux_s	= emu_mux_inst_ae ? sig_02_4_3_vc_s	: sig_02[4:3];
		assign sig_05_emux_s	= emu_mux_inst_ae ? sig_05_vc_s	: sig_05;
		assign sig_06_emux_s	= emu_mux_inst_ae ? sig_06_vc_s	: sig_06;
		assign sig_07_emux_s	= emu_mux_inst_ae ? sig_07_vc_s	: sig_07;
		assign sig_08_emux_s	= emu_mux_inst_ae ? sig_08_vc_s	: sig_08;
		assign sig_i_ae_emux_s	= emu_mux_inst_ae ? sig_i_ae_vc_s	: sig_i_ae;
	`endif
		// Generated Instance Port Map for inst_ae
		ent_ae inst_ae (
		`ifdef insert_emu_mux_inst_ae
			.port_ae_2[1:0](sig_02_1_0_emux_s),
		`else
			.port_ae_2[1:0](sig_02[1:0]), 	// Use internally test2, no port generated
		`endif
		`ifdef insert_emu_mux_inst_ae
			.port_ae_2[4:3](sig_02_4_3_emux_s),
		`else
			.port_ae_2[4:3](sig_02[4:3]), 	// Use internally test2, no port generated
		`endif
		`ifdef insert_emu_mux_inst_ae
			.port_ae_5(sig_05_emux_s),
		`else
			.port_ae_5(sig_05),	// Bus, single bits go to outsideBus, single bits go to outside, will create p_mix_sig_5_2_2_goBu...
		`endif
		`ifdef insert_emu_mux_inst_ae
			.port_ae_6(sig_06_emux_s),
		`else
			.port_ae_6(sig_06),	// Conflicting definition (X2)
		`endif
		`ifdef insert_emu_mux_inst_ae
			.sig_07(sig_07_emux_s),
		`else
			.sig_07(sig_07),	// Conflicting definition, IN false!
		`endif
		`ifdef insert_emu_mux_inst_ae
			.sig_08(sig_08_emux_s),
		`else
			.sig_08(sig_08),	// VHDL intermediate needed (port name)
		`endif
		`ifdef insert_emu_mux_inst_ae
			.sig_i_ae(sig_i_ae_emux_s),
		`else
			.sig_i_ae(sig_i_ae),	// Input Bus
		`endif
			.sig_o_ae(sig_o_ae)	// Output Bus
		);
		// End of Generated Instance Port Map for inst_ae
endmodule