module DSP_MULTIPLIER #(
`ifdef XIL_TIMING
  parameter LOC = "UNPLACED",
`endif
  parameter AMULTSEL = "A",
  parameter BMULTSEL = "B",
  parameter USE_MULT = "MULTIPLY"
)(
  output AMULT26,
  output BMULT17,
  output [44:0] U,
  output [44:0] V,
  input [26:0] A2A1,
  input [26:0] AD_DATA,
  input [17:0] B2B1
);
// define constants
  localparam MODULE_NAME = "DSP_MULTIPLIER";
// Parameter encodings and registers
  localparam AMULTSEL_A = 0;
  localparam AMULTSEL_AD = 1;
  localparam BMULTSEL_AD = 1;
  localparam BMULTSEL_B = 0;
  localparam USE_MULT_DYNAMIC = 1;
  localparam USE_MULT_MULTIPLY = 0;
  localparam USE_MULT_NONE = 2;
  reg trig_attr;
// include dynamic registers - XILINX test only
`ifdef XIL_DR
  `include "DSP_MULTIPLIER_dr.v"
`else
  reg [16:1] AMULTSEL_REG = AMULTSEL;
  reg [16:1] BMULTSEL_REG = BMULTSEL;
  reg [64:1] USE_MULT_REG = USE_MULT;
`endif
`ifdef XIL_XECLIB
  wire AMULTSEL_BIN;
  wire BMULTSEL_BIN;
  wire [1:0] USE_MULT_BIN;
`else
  reg AMULTSEL_BIN;
  reg BMULTSEL_BIN;
  reg [1:0] USE_MULT_BIN;
`endif
`ifdef XIL_XECLIB
  reg glblGSR = 1'b0;
`else
  tri0 glblGSR = glbl.GSR;
`endif
`ifndef XIL_XECLIB
  reg attr_test;
  reg attr_err;
initial begin
  trig_attr = 1'b0;
`ifdef XIL_ATTR_TEST
  attr_test = 1'b1;
`else
  attr_test = 1'b0;
`endif
  attr_err = 1'b0;
  #1;
  trig_attr = ~trig_attr;
end
`endif
`ifdef XIL_XECLIB
  assign AMULTSEL_BIN =
    (AMULTSEL_REG == "A") ? AMULTSEL_A :
    (AMULTSEL_REG == "AD") ? AMULTSEL_AD :
     AMULTSEL_A;
  assign BMULTSEL_BIN =
    (BMULTSEL_REG == "B") ? BMULTSEL_B :
    (BMULTSEL_REG == "AD") ? BMULTSEL_AD :
     BMULTSEL_B;
  assign USE_MULT_BIN =
    (USE_MULT_REG == "MULTIPLY") ? USE_MULT_MULTIPLY :
    (USE_MULT_REG == "DYNAMIC") ? USE_MULT_DYNAMIC :
    (USE_MULT_REG == "NONE") ? USE_MULT_NONE :
     USE_MULT_MULTIPLY;
`else
always @(trig_attr) begin
#1;
  AMULTSEL_BIN =
    (AMULTSEL_REG == "A") ? AMULTSEL_A :
    (AMULTSEL_REG == "AD") ? AMULTSEL_AD :
     AMULTSEL_A;
  BMULTSEL_BIN =
    (BMULTSEL_REG == "B") ? BMULTSEL_B :
    (BMULTSEL_REG == "AD") ? BMULTSEL_AD :
     BMULTSEL_B;
  USE_MULT_BIN =
    (USE_MULT_REG == "MULTIPLY") ? USE_MULT_MULTIPLY :
    (USE_MULT_REG == "DYNAMIC") ? USE_MULT_DYNAMIC :
    (USE_MULT_REG == "NONE") ? USE_MULT_NONE :
     USE_MULT_MULTIPLY;
end
`endif
`ifndef XIL_TIMING
  initial begin
    $display("Error: [Unisim %s-100] SIMPRIM primitive is not intended for direct instantiation in RTL or functional netlists. This primitive is only available in the SIMPRIM library for implemented netlists, please ensure you are pointing to the correct library. Instance %m", MODULE_NAME);
    #1 $finish;
  end
`endif
`ifndef XIL_XECLIB
  always @(trig_attr) begin
  #1;
    if ((attr_test == 1'b1) ||
        ((AMULTSEL_REG != "A") &&
         (AMULTSEL_REG != "AD"))) begin
      $display("Error: [Unisim %s-101] AMULTSEL attribute is set to %s.  Legal values for this attribute are A or AD. Instance: %m", MODULE_NAME, AMULTSEL_REG);
      attr_err = 1'b1;
    end
    if ((attr_test == 1'b1) ||
        ((BMULTSEL_REG != "B") &&
         (BMULTSEL_REG != "AD"))) begin
      $display("Error: [Unisim %s-102] BMULTSEL attribute is set to %s.  Legal values for this attribute are B or AD. Instance: %m", MODULE_NAME, BMULTSEL_REG);
      attr_err = 1'b1;
    end
    if ((attr_test == 1'b1) ||
        ((USE_MULT_REG != "MULTIPLY") &&
         (USE_MULT_REG != "DYNAMIC") &&
         (USE_MULT_REG != "NONE"))) begin
      $display("Error: [Unisim %s-103] USE_MULT attribute is set to %s.  Legal values for this attribute are MULTIPLY, DYNAMIC or NONE. Instance: %m", MODULE_NAME, USE_MULT_REG);
      attr_err = 1'b1;
    end
    if (attr_err == 1'b1) #1 $finish;
  end
`endif
// begin behavioral model
  localparam M_WIDTH   = 45;
  reg [17:0] b_mult_mux;
  reg [26:0] a_mult_mux;
  reg [M_WIDTH-1:0] mult;
  reg [M_WIDTH-2:0] ps_u_mask;
  reg [M_WIDTH-2:0] ps_v_mask;
// initialize regs
`ifndef XIL_XECLIB
initial begin
  ps_u_mask = 44'h55555555555;
  ps_v_mask = 44'haaaaaaaaaaa;
end
`endif
always @(*) begin
  if (AMULTSEL_BIN == AMULTSEL_A) a_mult_mux = A2A1;
  else a_mult_mux = AD_DATA;
end
always @(*) begin
  if (BMULTSEL_BIN == BMULTSEL_B) b_mult_mux = B2B1;
  else b_mult_mux = AD_DATA;
end
  assign AMULT26 = a_mult_mux[26];
  assign BMULT17 = b_mult_mux[17];
// U[44],V[44]  11 when mult[44]=0,  10 when mult[44]=1
  assign U = {1'b1,      mult[43:0] & ps_u_mask};
  assign V = {~mult[44], mult[43:0] & ps_v_mask};
always @(*) begin
  if (USE_MULT_BIN == USE_MULT_NONE) mult = 45'b0;
  else mult = ({{18{a_mult_mux[26]}},a_mult_mux} * {{27{b_mult_mux[17]}},b_mult_mux});
end
// end behavioral model
`ifndef XIL_XECLIB
`ifdef XIL_TIMING
  specify
    (A2A1[0] => U[10]) = (0:0:0, 0:0:0);
    (A2A1[0] => U[11]) = (0:0:0, 0:0:0);
    (A2A1[0] => U[12]) = (0:0:0, 0:0:0);
    (A2A1[0] => U[13]) = (0:0:0, 0:0:0);
    (A2A1[0] => U[14]) = (0:0:0, 0:0:0);
    (A2A1[0] => U[15]) = (0:0:0, 0:0:0);
    (A2A1[0] => U[16]) = (0:0:0, 0:0:0);
    (A2A1[0] => U[17]) = (0:0:0, 0:0:0);
    (A2A1[0] => U[18]) = (0:0:0, 0:0:0);
    (A2A1[0] => U[19]) = (0:0:0, 0:0:0);
    (A2A1[0] => U[1]) = (0:0:0, 0:0:0);
    (A2A1[0] => U[20]) = (0:0:0, 0:0:0);
    (A2A1[0] => U[21]) = (0:0:0, 0:0:0);
    (A2A1[0] => U[2]) = (0:0:0, 0:0:0);
    (A2A1[0] => U[3]) = (0:0:0, 0:0:0);
    (A2A1[0] => U[4]) = (0:0:0, 0:0:0);
    (A2A1[0] => U[5]) = (0:0:0, 0:0:0);
    (A2A1[0] => U[6]) = (0:0:0, 0:0:0);
    (A2A1[0] => U[7]) = (0:0:0, 0:0:0);
    (A2A1[0] => U[8]) = (0:0:0, 0:0:0);
    (A2A1[0] => U[9]) = (0:0:0, 0:0:0);
    (A2A1[0] => V[0]) = (0:0:0, 0:0:0);
    (A2A1[0] => V[10]) = (0:0:0, 0:0:0);
    (A2A1[0] => V[11]) = (0:0:0, 0:0:0);
    (A2A1[0] => V[12]) = (0:0:0, 0:0:0);
    (A2A1[0] => V[13]) = (0:0:0, 0:0:0);
    (A2A1[0] => V[14]) = (0:0:0, 0:0:0);
    (A2A1[0] => V[15]) = (0:0:0, 0:0:0);
    (A2A1[0] => V[16]) = (0:0:0, 0:0:0);
    (A2A1[0] => V[17]) = (0:0:0, 0:0:0);
    (A2A1[0] => V[18]) = (0:0:0, 0:0:0);
    (A2A1[0] => V[19]) = (0:0:0, 0:0:0);
    (A2A1[0] => V[20]) = (0:0:0, 0:0:0);
    (A2A1[0] => V[4]) = (0:0:0, 0:0:0);
    (A2A1[0] => V[5]) = (0:0:0, 0:0:0);
    (A2A1[0] => V[6]) = (0:0:0, 0:0:0);
    (A2A1[0] => V[7]) = (0:0:0, 0:0:0);
    (A2A1[0] => V[8]) = (0:0:0, 0:0:0);
    (A2A1[0] => V[9]) = (0:0:0, 0:0:0);
    (A2A1[10] => U[11]) = (0:0:0, 0:0:0);
    (A2A1[10] => U[12]) = (0:0:0, 0:0:0);
    (A2A1[10] => U[13]) = (0:0:0, 0:0:0);
    (A2A1[10] => U[14]) = (0:0:0, 0:0:0);
    (A2A1[10] => U[15]) = (0:0:0, 0:0:0);
    (A2A1[10] => U[16]) = (0:0:0, 0:0:0);
    (A2A1[10] => U[17]) = (0:0:0, 0:0:0);
    (A2A1[10] => U[18]) = (0:0:0, 0:0:0);
    (A2A1[10] => U[19]) = (0:0:0, 0:0:0);
    (A2A1[10] => U[20]) = (0:0:0, 0:0:0);
    (A2A1[10] => U[21]) = (0:0:0, 0:0:0);
    (A2A1[10] => U[22]) = (0:0:0, 0:0:0);
    (A2A1[10] => U[23]) = (0:0:0, 0:0:0);
    (A2A1[10] => U[24]) = (0:0:0, 0:0:0);
    (A2A1[10] => U[25]) = (0:0:0, 0:0:0);
    (A2A1[10] => U[26]) = (0:0:0, 0:0:0);
    (A2A1[10] => U[27]) = (0:0:0, 0:0:0);
    (A2A1[10] => U[28]) = (0:0:0, 0:0:0);
    (A2A1[10] => U[29]) = (0:0:0, 0:0:0);
    (A2A1[10] => U[30]) = (0:0:0, 0:0:0);
    (A2A1[10] => U[31]) = (0:0:0, 0:0:0);
    (A2A1[10] => V[10]) = (0:0:0, 0:0:0);
    (A2A1[10] => V[11]) = (0:0:0, 0:0:0);
    (A2A1[10] => V[12]) = (0:0:0, 0:0:0);
    (A2A1[10] => V[13]) = (0:0:0, 0:0:0);
    (A2A1[10] => V[14]) = (0:0:0, 0:0:0);
    (A2A1[10] => V[15]) = (0:0:0, 0:0:0);
    (A2A1[10] => V[16]) = (0:0:0, 0:0:0);
    (A2A1[10] => V[17]) = (0:0:0, 0:0:0);
    (A2A1[10] => V[18]) = (0:0:0, 0:0:0);
    (A2A1[10] => V[19]) = (0:0:0, 0:0:0);
    (A2A1[10] => V[20]) = (0:0:0, 0:0:0);
    (A2A1[10] => V[21]) = (0:0:0, 0:0:0);
    (A2A1[10] => V[22]) = (0:0:0, 0:0:0);
    (A2A1[10] => V[23]) = (0:0:0, 0:0:0);
    (A2A1[10] => V[24]) = (0:0:0, 0:0:0);
    (A2A1[10] => V[25]) = (0:0:0, 0:0:0);
    (A2A1[10] => V[26]) = (0:0:0, 0:0:0);
    (A2A1[10] => V[27]) = (0:0:0, 0:0:0);
    (A2A1[10] => V[28]) = (0:0:0, 0:0:0);
    (A2A1[10] => V[29]) = (0:0:0, 0:0:0);
    (A2A1[10] => V[30]) = (0:0:0, 0:0:0);
    (A2A1[11] => U[12]) = (0:0:0, 0:0:0);
    (A2A1[11] => U[13]) = (0:0:0, 0:0:0);
    (A2A1[11] => U[14]) = (0:0:0, 0:0:0);
    (A2A1[11] => U[15]) = (0:0:0, 0:0:0);
    (A2A1[11] => U[16]) = (0:0:0, 0:0:0);
    (A2A1[11] => U[17]) = (0:0:0, 0:0:0);
    (A2A1[11] => U[18]) = (0:0:0, 0:0:0);
    (A2A1[11] => U[19]) = (0:0:0, 0:0:0);
    (A2A1[11] => U[20]) = (0:0:0, 0:0:0);
    (A2A1[11] => U[21]) = (0:0:0, 0:0:0);
    (A2A1[11] => U[22]) = (0:0:0, 0:0:0);
    (A2A1[11] => U[23]) = (0:0:0, 0:0:0);
    (A2A1[11] => U[24]) = (0:0:0, 0:0:0);
    (A2A1[11] => U[25]) = (0:0:0, 0:0:0);
    (A2A1[11] => U[26]) = (0:0:0, 0:0:0);
    (A2A1[11] => U[27]) = (0:0:0, 0:0:0);
    (A2A1[11] => U[28]) = (0:0:0, 0:0:0);
    (A2A1[11] => U[29]) = (0:0:0, 0:0:0);
    (A2A1[11] => U[30]) = (0:0:0, 0:0:0);
    (A2A1[11] => U[31]) = (0:0:0, 0:0:0);
    (A2A1[11] => U[32]) = (0:0:0, 0:0:0);
    (A2A1[11] => V[11]) = (0:0:0, 0:0:0);
    (A2A1[11] => V[12]) = (0:0:0, 0:0:0);
    (A2A1[11] => V[13]) = (0:0:0, 0:0:0);
    (A2A1[11] => V[14]) = (0:0:0, 0:0:0);
    (A2A1[11] => V[15]) = (0:0:0, 0:0:0);
    (A2A1[11] => V[16]) = (0:0:0, 0:0:0);
    (A2A1[11] => V[17]) = (0:0:0, 0:0:0);
    (A2A1[11] => V[18]) = (0:0:0, 0:0:0);
    (A2A1[11] => V[19]) = (0:0:0, 0:0:0);
    (A2A1[11] => V[20]) = (0:0:0, 0:0:0);
    (A2A1[11] => V[21]) = (0:0:0, 0:0:0);
    (A2A1[11] => V[22]) = (0:0:0, 0:0:0);
    (A2A1[11] => V[23]) = (0:0:0, 0:0:0);
    (A2A1[11] => V[24]) = (0:0:0, 0:0:0);
    (A2A1[11] => V[25]) = (0:0:0, 0:0:0);
    (A2A1[11] => V[26]) = (0:0:0, 0:0:0);
    (A2A1[11] => V[27]) = (0:0:0, 0:0:0);
    (A2A1[11] => V[28]) = (0:0:0, 0:0:0);
    (A2A1[11] => V[29]) = (0:0:0, 0:0:0);
    (A2A1[11] => V[30]) = (0:0:0, 0:0:0);
    (A2A1[11] => V[31]) = (0:0:0, 0:0:0);
    (A2A1[12] => U[13]) = (0:0:0, 0:0:0);
    (A2A1[12] => U[14]) = (0:0:0, 0:0:0);
    (A2A1[12] => U[15]) = (0:0:0, 0:0:0);
    (A2A1[12] => U[16]) = (0:0:0, 0:0:0);
    (A2A1[12] => U[17]) = (0:0:0, 0:0:0);
    (A2A1[12] => U[18]) = (0:0:0, 0:0:0);
    (A2A1[12] => U[19]) = (0:0:0, 0:0:0);
    (A2A1[12] => U[20]) = (0:0:0, 0:0:0);
    (A2A1[12] => U[21]) = (0:0:0, 0:0:0);
    (A2A1[12] => U[22]) = (0:0:0, 0:0:0);
    (A2A1[12] => U[23]) = (0:0:0, 0:0:0);
    (A2A1[12] => U[24]) = (0:0:0, 0:0:0);
    (A2A1[12] => U[25]) = (0:0:0, 0:0:0);
    (A2A1[12] => U[26]) = (0:0:0, 0:0:0);
    (A2A1[12] => U[27]) = (0:0:0, 0:0:0);
    (A2A1[12] => U[28]) = (0:0:0, 0:0:0);
    (A2A1[12] => U[29]) = (0:0:0, 0:0:0);
    (A2A1[12] => U[30]) = (0:0:0, 0:0:0);
    (A2A1[12] => U[31]) = (0:0:0, 0:0:0);
    (A2A1[12] => U[32]) = (0:0:0, 0:0:0);
    (A2A1[12] => U[33]) = (0:0:0, 0:0:0);
    (A2A1[12] => V[12]) = (0:0:0, 0:0:0);
    (A2A1[12] => V[13]) = (0:0:0, 0:0:0);
    (A2A1[12] => V[14]) = (0:0:0, 0:0:0);
    (A2A1[12] => V[15]) = (0:0:0, 0:0:0);
    (A2A1[12] => V[16]) = (0:0:0, 0:0:0);
    (A2A1[12] => V[17]) = (0:0:0, 0:0:0);
    (A2A1[12] => V[18]) = (0:0:0, 0:0:0);
    (A2A1[12] => V[19]) = (0:0:0, 0:0:0);
    (A2A1[12] => V[20]) = (0:0:0, 0:0:0);
    (A2A1[12] => V[21]) = (0:0:0, 0:0:0);
    (A2A1[12] => V[22]) = (0:0:0, 0:0:0);
    (A2A1[12] => V[23]) = (0:0:0, 0:0:0);
    (A2A1[12] => V[24]) = (0:0:0, 0:0:0);
    (A2A1[12] => V[25]) = (0:0:0, 0:0:0);
    (A2A1[12] => V[26]) = (0:0:0, 0:0:0);
    (A2A1[12] => V[27]) = (0:0:0, 0:0:0);
    (A2A1[12] => V[28]) = (0:0:0, 0:0:0);
    (A2A1[12] => V[29]) = (0:0:0, 0:0:0);
    (A2A1[12] => V[30]) = (0:0:0, 0:0:0);
    (A2A1[12] => V[31]) = (0:0:0, 0:0:0);
    (A2A1[12] => V[32]) = (0:0:0, 0:0:0);
    (A2A1[13] => U[14]) = (0:0:0, 0:0:0);
    (A2A1[13] => U[15]) = (0:0:0, 0:0:0);
    (A2A1[13] => U[16]) = (0:0:0, 0:0:0);
    (A2A1[13] => U[17]) = (0:0:0, 0:0:0);
    (A2A1[13] => U[18]) = (0:0:0, 0:0:0);
    (A2A1[13] => U[19]) = (0:0:0, 0:0:0);
    (A2A1[13] => U[20]) = (0:0:0, 0:0:0);
    (A2A1[13] => U[21]) = (0:0:0, 0:0:0);
    (A2A1[13] => U[22]) = (0:0:0, 0:0:0);
    (A2A1[13] => U[23]) = (0:0:0, 0:0:0);
    (A2A1[13] => U[24]) = (0:0:0, 0:0:0);
    (A2A1[13] => U[25]) = (0:0:0, 0:0:0);
    (A2A1[13] => U[26]) = (0:0:0, 0:0:0);
    (A2A1[13] => U[27]) = (0:0:0, 0:0:0);
    (A2A1[13] => U[28]) = (0:0:0, 0:0:0);
    (A2A1[13] => U[29]) = (0:0:0, 0:0:0);
    (A2A1[13] => U[30]) = (0:0:0, 0:0:0);
    (A2A1[13] => U[31]) = (0:0:0, 0:0:0);
    (A2A1[13] => U[32]) = (0:0:0, 0:0:0);
    (A2A1[13] => U[33]) = (0:0:0, 0:0:0);
    (A2A1[13] => U[34]) = (0:0:0, 0:0:0);
    (A2A1[13] => V[13]) = (0:0:0, 0:0:0);
    (A2A1[13] => V[14]) = (0:0:0, 0:0:0);
    (A2A1[13] => V[15]) = (0:0:0, 0:0:0);
    (A2A1[13] => V[16]) = (0:0:0, 0:0:0);
    (A2A1[13] => V[17]) = (0:0:0, 0:0:0);
    (A2A1[13] => V[18]) = (0:0:0, 0:0:0);
    (A2A1[13] => V[19]) = (0:0:0, 0:0:0);
    (A2A1[13] => V[20]) = (0:0:0, 0:0:0);
    (A2A1[13] => V[21]) = (0:0:0, 0:0:0);
    (A2A1[13] => V[22]) = (0:0:0, 0:0:0);
    (A2A1[13] => V[23]) = (0:0:0, 0:0:0);
    (A2A1[13] => V[24]) = (0:0:0, 0:0:0);
    (A2A1[13] => V[25]) = (0:0:0, 0:0:0);
    (A2A1[13] => V[26]) = (0:0:0, 0:0:0);
    (A2A1[13] => V[27]) = (0:0:0, 0:0:0);
    (A2A1[13] => V[28]) = (0:0:0, 0:0:0);
    (A2A1[13] => V[29]) = (0:0:0, 0:0:0);
    (A2A1[13] => V[30]) = (0:0:0, 0:0:0);
    (A2A1[13] => V[31]) = (0:0:0, 0:0:0);
    (A2A1[13] => V[32]) = (0:0:0, 0:0:0);
    (A2A1[13] => V[33]) = (0:0:0, 0:0:0);
    (A2A1[14] => U[15]) = (0:0:0, 0:0:0);
    (A2A1[14] => U[16]) = (0:0:0, 0:0:0);
    (A2A1[14] => U[17]) = (0:0:0, 0:0:0);
    (A2A1[14] => U[18]) = (0:0:0, 0:0:0);
    (A2A1[14] => U[19]) = (0:0:0, 0:0:0);
    (A2A1[14] => U[20]) = (0:0:0, 0:0:0);
    (A2A1[14] => U[21]) = (0:0:0, 0:0:0);
    (A2A1[14] => U[22]) = (0:0:0, 0:0:0);
    (A2A1[14] => U[23]) = (0:0:0, 0:0:0);
    (A2A1[14] => U[24]) = (0:0:0, 0:0:0);
    (A2A1[14] => U[25]) = (0:0:0, 0:0:0);
    (A2A1[14] => U[26]) = (0:0:0, 0:0:0);
    (A2A1[14] => U[27]) = (0:0:0, 0:0:0);
    (A2A1[14] => U[28]) = (0:0:0, 0:0:0);
    (A2A1[14] => U[29]) = (0:0:0, 0:0:0);
    (A2A1[14] => U[30]) = (0:0:0, 0:0:0);
    (A2A1[14] => U[31]) = (0:0:0, 0:0:0);
    (A2A1[14] => U[32]) = (0:0:0, 0:0:0);
    (A2A1[14] => U[33]) = (0:0:0, 0:0:0);
    (A2A1[14] => U[34]) = (0:0:0, 0:0:0);
    (A2A1[14] => V[14]) = (0:0:0, 0:0:0);
    (A2A1[14] => V[15]) = (0:0:0, 0:0:0);
    (A2A1[14] => V[16]) = (0:0:0, 0:0:0);
    (A2A1[14] => V[17]) = (0:0:0, 0:0:0);
    (A2A1[14] => V[18]) = (0:0:0, 0:0:0);
    (A2A1[14] => V[19]) = (0:0:0, 0:0:0);
    (A2A1[14] => V[20]) = (0:0:0, 0:0:0);
    (A2A1[14] => V[21]) = (0:0:0, 0:0:0);
    (A2A1[14] => V[22]) = (0:0:0, 0:0:0);
    (A2A1[14] => V[23]) = (0:0:0, 0:0:0);
    (A2A1[14] => V[24]) = (0:0:0, 0:0:0);
    (A2A1[14] => V[25]) = (0:0:0, 0:0:0);
    (A2A1[14] => V[26]) = (0:0:0, 0:0:0);
    (A2A1[14] => V[27]) = (0:0:0, 0:0:0);
    (A2A1[14] => V[28]) = (0:0:0, 0:0:0);
    (A2A1[14] => V[29]) = (0:0:0, 0:0:0);
    (A2A1[14] => V[30]) = (0:0:0, 0:0:0);
    (A2A1[14] => V[31]) = (0:0:0, 0:0:0);
    (A2A1[14] => V[32]) = (0:0:0, 0:0:0);
    (A2A1[14] => V[33]) = (0:0:0, 0:0:0);
    (A2A1[15] => U[16]) = (0:0:0, 0:0:0);
    (A2A1[15] => U[17]) = (0:0:0, 0:0:0);
    (A2A1[15] => U[18]) = (0:0:0, 0:0:0);
    (A2A1[15] => U[19]) = (0:0:0, 0:0:0);
    (A2A1[15] => U[20]) = (0:0:0, 0:0:0);
    (A2A1[15] => U[21]) = (0:0:0, 0:0:0);
    (A2A1[15] => U[22]) = (0:0:0, 0:0:0);
    (A2A1[15] => U[23]) = (0:0:0, 0:0:0);
    (A2A1[15] => U[24]) = (0:0:0, 0:0:0);
    (A2A1[15] => U[25]) = (0:0:0, 0:0:0);
    (A2A1[15] => U[26]) = (0:0:0, 0:0:0);
    (A2A1[15] => U[27]) = (0:0:0, 0:0:0);
    (A2A1[15] => U[28]) = (0:0:0, 0:0:0);
    (A2A1[15] => U[29]) = (0:0:0, 0:0:0);
    (A2A1[15] => U[30]) = (0:0:0, 0:0:0);
    (A2A1[15] => U[31]) = (0:0:0, 0:0:0);
    (A2A1[15] => U[32]) = (0:0:0, 0:0:0);
    (A2A1[15] => U[33]) = (0:0:0, 0:0:0);
    (A2A1[15] => U[34]) = (0:0:0, 0:0:0);
    (A2A1[15] => U[35]) = (0:0:0, 0:0:0);
    (A2A1[15] => U[36]) = (0:0:0, 0:0:0);
    (A2A1[15] => V[15]) = (0:0:0, 0:0:0);
    (A2A1[15] => V[16]) = (0:0:0, 0:0:0);
    (A2A1[15] => V[17]) = (0:0:0, 0:0:0);
    (A2A1[15] => V[18]) = (0:0:0, 0:0:0);
    (A2A1[15] => V[19]) = (0:0:0, 0:0:0);
    (A2A1[15] => V[20]) = (0:0:0, 0:0:0);
    (A2A1[15] => V[21]) = (0:0:0, 0:0:0);
    (A2A1[15] => V[22]) = (0:0:0, 0:0:0);
    (A2A1[15] => V[23]) = (0:0:0, 0:0:0);
    (A2A1[15] => V[24]) = (0:0:0, 0:0:0);
    (A2A1[15] => V[25]) = (0:0:0, 0:0:0);
    (A2A1[15] => V[26]) = (0:0:0, 0:0:0);
    (A2A1[15] => V[27]) = (0:0:0, 0:0:0);
    (A2A1[15] => V[28]) = (0:0:0, 0:0:0);
    (A2A1[15] => V[29]) = (0:0:0, 0:0:0);
    (A2A1[15] => V[30]) = (0:0:0, 0:0:0);
    (A2A1[15] => V[31]) = (0:0:0, 0:0:0);
    (A2A1[15] => V[32]) = (0:0:0, 0:0:0);
    (A2A1[15] => V[33]) = (0:0:0, 0:0:0);
    (A2A1[15] => V[34]) = (0:0:0, 0:0:0);
    (A2A1[15] => V[35]) = (0:0:0, 0:0:0);
    (A2A1[16] => U[17]) = (0:0:0, 0:0:0);
    (A2A1[16] => U[18]) = (0:0:0, 0:0:0);
    (A2A1[16] => U[19]) = (0:0:0, 0:0:0);
    (A2A1[16] => U[20]) = (0:0:0, 0:0:0);
    (A2A1[16] => U[21]) = (0:0:0, 0:0:0);
    (A2A1[16] => U[22]) = (0:0:0, 0:0:0);
    (A2A1[16] => U[23]) = (0:0:0, 0:0:0);
    (A2A1[16] => U[24]) = (0:0:0, 0:0:0);
    (A2A1[16] => U[25]) = (0:0:0, 0:0:0);
    (A2A1[16] => U[26]) = (0:0:0, 0:0:0);
    (A2A1[16] => U[27]) = (0:0:0, 0:0:0);
    (A2A1[16] => U[28]) = (0:0:0, 0:0:0);
    (A2A1[16] => U[29]) = (0:0:0, 0:0:0);
    (A2A1[16] => U[30]) = (0:0:0, 0:0:0);
    (A2A1[16] => U[31]) = (0:0:0, 0:0:0);
    (A2A1[16] => U[32]) = (0:0:0, 0:0:0);
    (A2A1[16] => U[33]) = (0:0:0, 0:0:0);
    (A2A1[16] => U[34]) = (0:0:0, 0:0:0);
    (A2A1[16] => U[35]) = (0:0:0, 0:0:0);
    (A2A1[16] => U[36]) = (0:0:0, 0:0:0);
    (A2A1[16] => V[16]) = (0:0:0, 0:0:0);
    (A2A1[16] => V[17]) = (0:0:0, 0:0:0);
    (A2A1[16] => V[18]) = (0:0:0, 0:0:0);
    (A2A1[16] => V[19]) = (0:0:0, 0:0:0);
    (A2A1[16] => V[20]) = (0:0:0, 0:0:0);
    (A2A1[16] => V[21]) = (0:0:0, 0:0:0);
    (A2A1[16] => V[22]) = (0:0:0, 0:0:0);
    (A2A1[16] => V[23]) = (0:0:0, 0:0:0);
    (A2A1[16] => V[24]) = (0:0:0, 0:0:0);
    (A2A1[16] => V[25]) = (0:0:0, 0:0:0);
    (A2A1[16] => V[26]) = (0:0:0, 0:0:0);
    (A2A1[16] => V[27]) = (0:0:0, 0:0:0);
    (A2A1[16] => V[28]) = (0:0:0, 0:0:0);
    (A2A1[16] => V[29]) = (0:0:0, 0:0:0);
    (A2A1[16] => V[30]) = (0:0:0, 0:0:0);
    (A2A1[16] => V[31]) = (0:0:0, 0:0:0);
    (A2A1[16] => V[32]) = (0:0:0, 0:0:0);
    (A2A1[16] => V[33]) = (0:0:0, 0:0:0);
    (A2A1[16] => V[34]) = (0:0:0, 0:0:0);
    (A2A1[16] => V[35]) = (0:0:0, 0:0:0);
    (A2A1[17] => U[18]) = (0:0:0, 0:0:0);
    (A2A1[17] => U[19]) = (0:0:0, 0:0:0);
    (A2A1[17] => U[20]) = (0:0:0, 0:0:0);
    (A2A1[17] => U[21]) = (0:0:0, 0:0:0);
    (A2A1[17] => U[22]) = (0:0:0, 0:0:0);
    (A2A1[17] => U[23]) = (0:0:0, 0:0:0);
    (A2A1[17] => U[24]) = (0:0:0, 0:0:0);
    (A2A1[17] => U[25]) = (0:0:0, 0:0:0);
    (A2A1[17] => U[26]) = (0:0:0, 0:0:0);
    (A2A1[17] => U[27]) = (0:0:0, 0:0:0);
    (A2A1[17] => U[28]) = (0:0:0, 0:0:0);
    (A2A1[17] => U[29]) = (0:0:0, 0:0:0);
    (A2A1[17] => U[30]) = (0:0:0, 0:0:0);
    (A2A1[17] => U[31]) = (0:0:0, 0:0:0);
    (A2A1[17] => U[32]) = (0:0:0, 0:0:0);
    (A2A1[17] => U[33]) = (0:0:0, 0:0:0);
    (A2A1[17] => U[34]) = (0:0:0, 0:0:0);
    (A2A1[17] => U[35]) = (0:0:0, 0:0:0);
    (A2A1[17] => U[36]) = (0:0:0, 0:0:0);
    (A2A1[17] => U[37]) = (0:0:0, 0:0:0);
    (A2A1[17] => V[17]) = (0:0:0, 0:0:0);
    (A2A1[17] => V[18]) = (0:0:0, 0:0:0);
    (A2A1[17] => V[19]) = (0:0:0, 0:0:0);
    (A2A1[17] => V[20]) = (0:0:0, 0:0:0);
    (A2A1[17] => V[21]) = (0:0:0, 0:0:0);
    (A2A1[17] => V[22]) = (0:0:0, 0:0:0);
    (A2A1[17] => V[23]) = (0:0:0, 0:0:0);
    (A2A1[17] => V[24]) = (0:0:0, 0:0:0);
    (A2A1[17] => V[25]) = (0:0:0, 0:0:0);
    (A2A1[17] => V[26]) = (0:0:0, 0:0:0);
    (A2A1[17] => V[27]) = (0:0:0, 0:0:0);
    (A2A1[17] => V[28]) = (0:0:0, 0:0:0);
    (A2A1[17] => V[29]) = (0:0:0, 0:0:0);
    (A2A1[17] => V[30]) = (0:0:0, 0:0:0);
    (A2A1[17] => V[31]) = (0:0:0, 0:0:0);
    (A2A1[17] => V[32]) = (0:0:0, 0:0:0);
    (A2A1[17] => V[33]) = (0:0:0, 0:0:0);
    (A2A1[17] => V[34]) = (0:0:0, 0:0:0);
    (A2A1[17] => V[35]) = (0:0:0, 0:0:0);
    (A2A1[17] => V[36]) = (0:0:0, 0:0:0);
    (A2A1[18] => U[19]) = (0:0:0, 0:0:0);
    (A2A1[18] => U[20]) = (0:0:0, 0:0:0);
    (A2A1[18] => U[21]) = (0:0:0, 0:0:0);
    (A2A1[18] => U[22]) = (0:0:0, 0:0:0);
    (A2A1[18] => U[23]) = (0:0:0, 0:0:0);
    (A2A1[18] => U[24]) = (0:0:0, 0:0:0);
    (A2A1[18] => U[25]) = (0:0:0, 0:0:0);
    (A2A1[18] => U[26]) = (0:0:0, 0:0:0);
    (A2A1[18] => U[27]) = (0:0:0, 0:0:0);
    (A2A1[18] => U[28]) = (0:0:0, 0:0:0);
    (A2A1[18] => U[29]) = (0:0:0, 0:0:0);
    (A2A1[18] => U[30]) = (0:0:0, 0:0:0);
    (A2A1[18] => U[31]) = (0:0:0, 0:0:0);
    (A2A1[18] => U[32]) = (0:0:0, 0:0:0);
    (A2A1[18] => U[33]) = (0:0:0, 0:0:0);
    (A2A1[18] => U[34]) = (0:0:0, 0:0:0);
    (A2A1[18] => U[35]) = (0:0:0, 0:0:0);
    (A2A1[18] => U[36]) = (0:0:0, 0:0:0);
    (A2A1[18] => U[37]) = (0:0:0, 0:0:0);
    (A2A1[18] => U[38]) = (0:0:0, 0:0:0);
    (A2A1[18] => V[18]) = (0:0:0, 0:0:0);
    (A2A1[18] => V[19]) = (0:0:0, 0:0:0);
    (A2A1[18] => V[20]) = (0:0:0, 0:0:0);
    (A2A1[18] => V[21]) = (0:0:0, 0:0:0);
    (A2A1[18] => V[22]) = (0:0:0, 0:0:0);
    (A2A1[18] => V[23]) = (0:0:0, 0:0:0);
    (A2A1[18] => V[24]) = (0:0:0, 0:0:0);
    (A2A1[18] => V[25]) = (0:0:0, 0:0:0);
    (A2A1[18] => V[26]) = (0:0:0, 0:0:0);
    (A2A1[18] => V[27]) = (0:0:0, 0:0:0);
    (A2A1[18] => V[28]) = (0:0:0, 0:0:0);
    (A2A1[18] => V[29]) = (0:0:0, 0:0:0);
    (A2A1[18] => V[30]) = (0:0:0, 0:0:0);
    (A2A1[18] => V[31]) = (0:0:0, 0:0:0);
    (A2A1[18] => V[32]) = (0:0:0, 0:0:0);
    (A2A1[18] => V[33]) = (0:0:0, 0:0:0);
    (A2A1[18] => V[34]) = (0:0:0, 0:0:0);
    (A2A1[18] => V[35]) = (0:0:0, 0:0:0);
    (A2A1[18] => V[36]) = (0:0:0, 0:0:0);
    (A2A1[18] => V[37]) = (0:0:0, 0:0:0);
    (A2A1[19] => U[20]) = (0:0:0, 0:0:0);
    (A2A1[19] => U[21]) = (0:0:0, 0:0:0);
    (A2A1[19] => U[22]) = (0:0:0, 0:0:0);
    (A2A1[19] => U[23]) = (0:0:0, 0:0:0);
    (A2A1[19] => U[24]) = (0:0:0, 0:0:0);
    (A2A1[19] => U[25]) = (0:0:0, 0:0:0);
    (A2A1[19] => U[26]) = (0:0:0, 0:0:0);
    (A2A1[19] => U[27]) = (0:0:0, 0:0:0);
    (A2A1[19] => U[28]) = (0:0:0, 0:0:0);
    (A2A1[19] => U[29]) = (0:0:0, 0:0:0);
    (A2A1[19] => U[30]) = (0:0:0, 0:0:0);
    (A2A1[19] => U[31]) = (0:0:0, 0:0:0);
    (A2A1[19] => U[32]) = (0:0:0, 0:0:0);
    (A2A1[19] => U[33]) = (0:0:0, 0:0:0);
    (A2A1[19] => U[34]) = (0:0:0, 0:0:0);
    (A2A1[19] => U[35]) = (0:0:0, 0:0:0);
    (A2A1[19] => U[36]) = (0:0:0, 0:0:0);
    (A2A1[19] => U[37]) = (0:0:0, 0:0:0);
    (A2A1[19] => U[38]) = (0:0:0, 0:0:0);
    (A2A1[19] => U[39]) = (0:0:0, 0:0:0);
    (A2A1[19] => V[19]) = (0:0:0, 0:0:0);
    (A2A1[19] => V[20]) = (0:0:0, 0:0:0);
    (A2A1[19] => V[21]) = (0:0:0, 0:0:0);
    (A2A1[19] => V[22]) = (0:0:0, 0:0:0);
    (A2A1[19] => V[23]) = (0:0:0, 0:0:0);
    (A2A1[19] => V[24]) = (0:0:0, 0:0:0);
    (A2A1[19] => V[25]) = (0:0:0, 0:0:0);
    (A2A1[19] => V[26]) = (0:0:0, 0:0:0);
    (A2A1[19] => V[27]) = (0:0:0, 0:0:0);
    (A2A1[19] => V[28]) = (0:0:0, 0:0:0);
    (A2A1[19] => V[29]) = (0:0:0, 0:0:0);
    (A2A1[19] => V[30]) = (0:0:0, 0:0:0);
    (A2A1[19] => V[31]) = (0:0:0, 0:0:0);
    (A2A1[19] => V[32]) = (0:0:0, 0:0:0);
    (A2A1[19] => V[33]) = (0:0:0, 0:0:0);
    (A2A1[19] => V[34]) = (0:0:0, 0:0:0);
    (A2A1[19] => V[35]) = (0:0:0, 0:0:0);
    (A2A1[19] => V[36]) = (0:0:0, 0:0:0);
    (A2A1[19] => V[37]) = (0:0:0, 0:0:0);
    (A2A1[19] => V[38]) = (0:0:0, 0:0:0);
    (A2A1[1] => U[10]) = (0:0:0, 0:0:0);
    (A2A1[1] => U[11]) = (0:0:0, 0:0:0);
    (A2A1[1] => U[12]) = (0:0:0, 0:0:0);
    (A2A1[1] => U[13]) = (0:0:0, 0:0:0);
    (A2A1[1] => U[14]) = (0:0:0, 0:0:0);
    (A2A1[1] => U[15]) = (0:0:0, 0:0:0);
    (A2A1[1] => U[16]) = (0:0:0, 0:0:0);
    (A2A1[1] => U[17]) = (0:0:0, 0:0:0);
    (A2A1[1] => U[18]) = (0:0:0, 0:0:0);
    (A2A1[1] => U[19]) = (0:0:0, 0:0:0);
    (A2A1[1] => U[1]) = (0:0:0, 0:0:0);
    (A2A1[1] => U[20]) = (0:0:0, 0:0:0);
    (A2A1[1] => U[21]) = (0:0:0, 0:0:0);
    (A2A1[1] => U[22]) = (0:0:0, 0:0:0);
    (A2A1[1] => U[2]) = (0:0:0, 0:0:0);
    (A2A1[1] => U[3]) = (0:0:0, 0:0:0);
    (A2A1[1] => U[4]) = (0:0:0, 0:0:0);
    (A2A1[1] => U[5]) = (0:0:0, 0:0:0);
    (A2A1[1] => U[6]) = (0:0:0, 0:0:0);
    (A2A1[1] => U[7]) = (0:0:0, 0:0:0);
    (A2A1[1] => U[8]) = (0:0:0, 0:0:0);
    (A2A1[1] => U[9]) = (0:0:0, 0:0:0);
    (A2A1[1] => V[10]) = (0:0:0, 0:0:0);
    (A2A1[1] => V[11]) = (0:0:0, 0:0:0);
    (A2A1[1] => V[12]) = (0:0:0, 0:0:0);
    (A2A1[1] => V[13]) = (0:0:0, 0:0:0);
    (A2A1[1] => V[14]) = (0:0:0, 0:0:0);
    (A2A1[1] => V[15]) = (0:0:0, 0:0:0);
    (A2A1[1] => V[16]) = (0:0:0, 0:0:0);
    (A2A1[1] => V[17]) = (0:0:0, 0:0:0);
    (A2A1[1] => V[18]) = (0:0:0, 0:0:0);
    (A2A1[1] => V[19]) = (0:0:0, 0:0:0);
    (A2A1[1] => V[20]) = (0:0:0, 0:0:0);
    (A2A1[1] => V[21]) = (0:0:0, 0:0:0);
    (A2A1[1] => V[4]) = (0:0:0, 0:0:0);
    (A2A1[1] => V[5]) = (0:0:0, 0:0:0);
    (A2A1[1] => V[6]) = (0:0:0, 0:0:0);
    (A2A1[1] => V[7]) = (0:0:0, 0:0:0);
    (A2A1[1] => V[8]) = (0:0:0, 0:0:0);
    (A2A1[1] => V[9]) = (0:0:0, 0:0:0);
    (A2A1[20] => U[21]) = (0:0:0, 0:0:0);
    (A2A1[20] => U[22]) = (0:0:0, 0:0:0);
    (A2A1[20] => U[23]) = (0:0:0, 0:0:0);
    (A2A1[20] => U[24]) = (0:0:0, 0:0:0);
    (A2A1[20] => U[25]) = (0:0:0, 0:0:0);
    (A2A1[20] => U[26]) = (0:0:0, 0:0:0);
    (A2A1[20] => U[27]) = (0:0:0, 0:0:0);
    (A2A1[20] => U[28]) = (0:0:0, 0:0:0);
    (A2A1[20] => U[29]) = (0:0:0, 0:0:0);
    (A2A1[20] => U[30]) = (0:0:0, 0:0:0);
    (A2A1[20] => U[31]) = (0:0:0, 0:0:0);
    (A2A1[20] => U[32]) = (0:0:0, 0:0:0);
    (A2A1[20] => U[33]) = (0:0:0, 0:0:0);
    (A2A1[20] => U[34]) = (0:0:0, 0:0:0);
    (A2A1[20] => U[35]) = (0:0:0, 0:0:0);
    (A2A1[20] => U[36]) = (0:0:0, 0:0:0);
    (A2A1[20] => U[37]) = (0:0:0, 0:0:0);
    (A2A1[20] => U[38]) = (0:0:0, 0:0:0);
    (A2A1[20] => U[39]) = (0:0:0, 0:0:0);
    (A2A1[20] => V[20]) = (0:0:0, 0:0:0);
    (A2A1[20] => V[21]) = (0:0:0, 0:0:0);
    (A2A1[20] => V[22]) = (0:0:0, 0:0:0);
    (A2A1[20] => V[23]) = (0:0:0, 0:0:0);
    (A2A1[20] => V[24]) = (0:0:0, 0:0:0);
    (A2A1[20] => V[25]) = (0:0:0, 0:0:0);
    (A2A1[20] => V[26]) = (0:0:0, 0:0:0);
    (A2A1[20] => V[27]) = (0:0:0, 0:0:0);
    (A2A1[20] => V[28]) = (0:0:0, 0:0:0);
    (A2A1[20] => V[29]) = (0:0:0, 0:0:0);
    (A2A1[20] => V[30]) = (0:0:0, 0:0:0);
    (A2A1[20] => V[31]) = (0:0:0, 0:0:0);
    (A2A1[20] => V[32]) = (0:0:0, 0:0:0);
    (A2A1[20] => V[33]) = (0:0:0, 0:0:0);
    (A2A1[20] => V[34]) = (0:0:0, 0:0:0);
    (A2A1[20] => V[35]) = (0:0:0, 0:0:0);
    (A2A1[20] => V[36]) = (0:0:0, 0:0:0);
    (A2A1[20] => V[37]) = (0:0:0, 0:0:0);
    (A2A1[20] => V[38]) = (0:0:0, 0:0:0);
    (A2A1[21] => U[22]) = (0:0:0, 0:0:0);
    (A2A1[21] => U[23]) = (0:0:0, 0:0:0);
    (A2A1[21] => U[24]) = (0:0:0, 0:0:0);
    (A2A1[21] => U[25]) = (0:0:0, 0:0:0);
    (A2A1[21] => U[26]) = (0:0:0, 0:0:0);
    (A2A1[21] => U[27]) = (0:0:0, 0:0:0);
    (A2A1[21] => U[28]) = (0:0:0, 0:0:0);
    (A2A1[21] => U[29]) = (0:0:0, 0:0:0);
    (A2A1[21] => U[30]) = (0:0:0, 0:0:0);
    (A2A1[21] => U[31]) = (0:0:0, 0:0:0);
    (A2A1[21] => U[32]) = (0:0:0, 0:0:0);
    (A2A1[21] => U[33]) = (0:0:0, 0:0:0);
    (A2A1[21] => U[34]) = (0:0:0, 0:0:0);
    (A2A1[21] => U[35]) = (0:0:0, 0:0:0);
    (A2A1[21] => U[36]) = (0:0:0, 0:0:0);
    (A2A1[21] => U[37]) = (0:0:0, 0:0:0);
    (A2A1[21] => U[38]) = (0:0:0, 0:0:0);
    (A2A1[21] => U[39]) = (0:0:0, 0:0:0);
    (A2A1[21] => U[40]) = (0:0:0, 0:0:0);
    (A2A1[21] => V[21]) = (0:0:0, 0:0:0);
    (A2A1[21] => V[22]) = (0:0:0, 0:0:0);
    (A2A1[21] => V[23]) = (0:0:0, 0:0:0);
    (A2A1[21] => V[24]) = (0:0:0, 0:0:0);
    (A2A1[21] => V[25]) = (0:0:0, 0:0:0);
    (A2A1[21] => V[26]) = (0:0:0, 0:0:0);
    (A2A1[21] => V[27]) = (0:0:0, 0:0:0);
    (A2A1[21] => V[28]) = (0:0:0, 0:0:0);
    (A2A1[21] => V[29]) = (0:0:0, 0:0:0);
    (A2A1[21] => V[30]) = (0:0:0, 0:0:0);
    (A2A1[21] => V[31]) = (0:0:0, 0:0:0);
    (A2A1[21] => V[32]) = (0:0:0, 0:0:0);
    (A2A1[21] => V[33]) = (0:0:0, 0:0:0);
    (A2A1[21] => V[34]) = (0:0:0, 0:0:0);
    (A2A1[21] => V[35]) = (0:0:0, 0:0:0);
    (A2A1[21] => V[36]) = (0:0:0, 0:0:0);
    (A2A1[21] => V[37]) = (0:0:0, 0:0:0);
    (A2A1[21] => V[38]) = (0:0:0, 0:0:0);
    (A2A1[21] => V[39]) = (0:0:0, 0:0:0);
    (A2A1[22] => U[23]) = (0:0:0, 0:0:0);
    (A2A1[22] => U[24]) = (0:0:0, 0:0:0);
    (A2A1[22] => U[25]) = (0:0:0, 0:0:0);
    (A2A1[22] => U[26]) = (0:0:0, 0:0:0);
    (A2A1[22] => U[27]) = (0:0:0, 0:0:0);
    (A2A1[22] => U[28]) = (0:0:0, 0:0:0);
    (A2A1[22] => U[29]) = (0:0:0, 0:0:0);
    (A2A1[22] => U[30]) = (0:0:0, 0:0:0);
    (A2A1[22] => U[31]) = (0:0:0, 0:0:0);
    (A2A1[22] => U[32]) = (0:0:0, 0:0:0);
    (A2A1[22] => U[33]) = (0:0:0, 0:0:0);
    (A2A1[22] => U[34]) = (0:0:0, 0:0:0);
    (A2A1[22] => U[35]) = (0:0:0, 0:0:0);
    (A2A1[22] => U[36]) = (0:0:0, 0:0:0);
    (A2A1[22] => U[37]) = (0:0:0, 0:0:0);
    (A2A1[22] => U[38]) = (0:0:0, 0:0:0);
    (A2A1[22] => U[39]) = (0:0:0, 0:0:0);
    (A2A1[22] => U[40]) = (0:0:0, 0:0:0);
    (A2A1[22] => U[41]) = (0:0:0, 0:0:0);
    (A2A1[22] => V[22]) = (0:0:0, 0:0:0);
    (A2A1[22] => V[23]) = (0:0:0, 0:0:0);
    (A2A1[22] => V[24]) = (0:0:0, 0:0:0);
    (A2A1[22] => V[25]) = (0:0:0, 0:0:0);
    (A2A1[22] => V[26]) = (0:0:0, 0:0:0);
    (A2A1[22] => V[27]) = (0:0:0, 0:0:0);
    (A2A1[22] => V[28]) = (0:0:0, 0:0:0);
    (A2A1[22] => V[29]) = (0:0:0, 0:0:0);
    (A2A1[22] => V[30]) = (0:0:0, 0:0:0);
    (A2A1[22] => V[31]) = (0:0:0, 0:0:0);
    (A2A1[22] => V[32]) = (0:0:0, 0:0:0);
    (A2A1[22] => V[33]) = (0:0:0, 0:0:0);
    (A2A1[22] => V[34]) = (0:0:0, 0:0:0);
    (A2A1[22] => V[35]) = (0:0:0, 0:0:0);
    (A2A1[22] => V[36]) = (0:0:0, 0:0:0);
    (A2A1[22] => V[37]) = (0:0:0, 0:0:0);
    (A2A1[22] => V[38]) = (0:0:0, 0:0:0);
    (A2A1[22] => V[39]) = (0:0:0, 0:0:0);
    (A2A1[22] => V[40]) = (0:0:0, 0:0:0);
    (A2A1[23] => U[24]) = (0:0:0, 0:0:0);
    (A2A1[23] => U[25]) = (0:0:0, 0:0:0);
    (A2A1[23] => U[26]) = (0:0:0, 0:0:0);
    (A2A1[23] => U[27]) = (0:0:0, 0:0:0);
    (A2A1[23] => U[28]) = (0:0:0, 0:0:0);
    (A2A1[23] => U[29]) = (0:0:0, 0:0:0);
    (A2A1[23] => U[30]) = (0:0:0, 0:0:0);
    (A2A1[23] => U[31]) = (0:0:0, 0:0:0);
    (A2A1[23] => U[32]) = (0:0:0, 0:0:0);
    (A2A1[23] => U[33]) = (0:0:0, 0:0:0);
    (A2A1[23] => U[34]) = (0:0:0, 0:0:0);
    (A2A1[23] => U[35]) = (0:0:0, 0:0:0);
    (A2A1[23] => U[36]) = (0:0:0, 0:0:0);
    (A2A1[23] => U[37]) = (0:0:0, 0:0:0);
    (A2A1[23] => U[38]) = (0:0:0, 0:0:0);
    (A2A1[23] => U[39]) = (0:0:0, 0:0:0);
    (A2A1[23] => U[40]) = (0:0:0, 0:0:0);
    (A2A1[23] => U[41]) = (0:0:0, 0:0:0);
    (A2A1[23] => U[42]) = (0:0:0, 0:0:0);
    (A2A1[23] => V[23]) = (0:0:0, 0:0:0);
    (A2A1[23] => V[24]) = (0:0:0, 0:0:0);
    (A2A1[23] => V[25]) = (0:0:0, 0:0:0);
    (A2A1[23] => V[26]) = (0:0:0, 0:0:0);
    (A2A1[23] => V[27]) = (0:0:0, 0:0:0);
    (A2A1[23] => V[28]) = (0:0:0, 0:0:0);
    (A2A1[23] => V[29]) = (0:0:0, 0:0:0);
    (A2A1[23] => V[30]) = (0:0:0, 0:0:0);
    (A2A1[23] => V[31]) = (0:0:0, 0:0:0);
    (A2A1[23] => V[32]) = (0:0:0, 0:0:0);
    (A2A1[23] => V[33]) = (0:0:0, 0:0:0);
    (A2A1[23] => V[34]) = (0:0:0, 0:0:0);
    (A2A1[23] => V[35]) = (0:0:0, 0:0:0);
    (A2A1[23] => V[36]) = (0:0:0, 0:0:0);
    (A2A1[23] => V[37]) = (0:0:0, 0:0:0);
    (A2A1[23] => V[38]) = (0:0:0, 0:0:0);
    (A2A1[23] => V[39]) = (0:0:0, 0:0:0);
    (A2A1[23] => V[40]) = (0:0:0, 0:0:0);
    (A2A1[23] => V[41]) = (0:0:0, 0:0:0);
    (A2A1[24] => U[25]) = (0:0:0, 0:0:0);
    (A2A1[24] => U[26]) = (0:0:0, 0:0:0);
    (A2A1[24] => U[27]) = (0:0:0, 0:0:0);
    (A2A1[24] => U[28]) = (0:0:0, 0:0:0);
    (A2A1[24] => U[29]) = (0:0:0, 0:0:0);
    (A2A1[24] => U[30]) = (0:0:0, 0:0:0);
    (A2A1[24] => U[31]) = (0:0:0, 0:0:0);
    (A2A1[24] => U[32]) = (0:0:0, 0:0:0);
    (A2A1[24] => U[33]) = (0:0:0, 0:0:0);
    (A2A1[24] => U[34]) = (0:0:0, 0:0:0);
    (A2A1[24] => U[35]) = (0:0:0, 0:0:0);
    (A2A1[24] => U[36]) = (0:0:0, 0:0:0);
    (A2A1[24] => U[37]) = (0:0:0, 0:0:0);
    (A2A1[24] => U[38]) = (0:0:0, 0:0:0);
    (A2A1[24] => U[39]) = (0:0:0, 0:0:0);
    (A2A1[24] => U[40]) = (0:0:0, 0:0:0);
    (A2A1[24] => U[41]) = (0:0:0, 0:0:0);
    (A2A1[24] => U[42]) = (0:0:0, 0:0:0);
    (A2A1[24] => V[24]) = (0:0:0, 0:0:0);
    (A2A1[24] => V[25]) = (0:0:0, 0:0:0);
    (A2A1[24] => V[26]) = (0:0:0, 0:0:0);
    (A2A1[24] => V[27]) = (0:0:0, 0:0:0);
    (A2A1[24] => V[28]) = (0:0:0, 0:0:0);
    (A2A1[24] => V[29]) = (0:0:0, 0:0:0);
    (A2A1[24] => V[30]) = (0:0:0, 0:0:0);
    (A2A1[24] => V[31]) = (0:0:0, 0:0:0);
    (A2A1[24] => V[32]) = (0:0:0, 0:0:0);
    (A2A1[24] => V[33]) = (0:0:0, 0:0:0);
    (A2A1[24] => V[34]) = (0:0:0, 0:0:0);
    (A2A1[24] => V[35]) = (0:0:0, 0:0:0);
    (A2A1[24] => V[36]) = (0:0:0, 0:0:0);
    (A2A1[24] => V[37]) = (0:0:0, 0:0:0);
    (A2A1[24] => V[38]) = (0:0:0, 0:0:0);
    (A2A1[24] => V[39]) = (0:0:0, 0:0:0);
    (A2A1[24] => V[40]) = (0:0:0, 0:0:0);
    (A2A1[24] => V[41]) = (0:0:0, 0:0:0);
    (A2A1[25] => U[26]) = (0:0:0, 0:0:0);
    (A2A1[25] => U[27]) = (0:0:0, 0:0:0);
    (A2A1[25] => U[28]) = (0:0:0, 0:0:0);
    (A2A1[25] => U[29]) = (0:0:0, 0:0:0);
    (A2A1[25] => U[30]) = (0:0:0, 0:0:0);
    (A2A1[25] => U[31]) = (0:0:0, 0:0:0);
    (A2A1[25] => U[32]) = (0:0:0, 0:0:0);
    (A2A1[25] => U[33]) = (0:0:0, 0:0:0);
    (A2A1[25] => U[34]) = (0:0:0, 0:0:0);
    (A2A1[25] => U[35]) = (0:0:0, 0:0:0);
    (A2A1[25] => U[36]) = (0:0:0, 0:0:0);
    (A2A1[25] => U[37]) = (0:0:0, 0:0:0);
    (A2A1[25] => U[38]) = (0:0:0, 0:0:0);
    (A2A1[25] => U[39]) = (0:0:0, 0:0:0);
    (A2A1[25] => U[40]) = (0:0:0, 0:0:0);
    (A2A1[25] => U[41]) = (0:0:0, 0:0:0);
    (A2A1[25] => U[42]) = (0:0:0, 0:0:0);
    (A2A1[25] => U[43]) = (0:0:0, 0:0:0);
    (A2A1[25] => V[25]) = (0:0:0, 0:0:0);
    (A2A1[25] => V[26]) = (0:0:0, 0:0:0);
    (A2A1[25] => V[27]) = (0:0:0, 0:0:0);
    (A2A1[25] => V[28]) = (0:0:0, 0:0:0);
    (A2A1[25] => V[29]) = (0:0:0, 0:0:0);
    (A2A1[25] => V[30]) = (0:0:0, 0:0:0);
    (A2A1[25] => V[31]) = (0:0:0, 0:0:0);
    (A2A1[25] => V[32]) = (0:0:0, 0:0:0);
    (A2A1[25] => V[33]) = (0:0:0, 0:0:0);
    (A2A1[25] => V[34]) = (0:0:0, 0:0:0);
    (A2A1[25] => V[35]) = (0:0:0, 0:0:0);
    (A2A1[25] => V[36]) = (0:0:0, 0:0:0);
    (A2A1[25] => V[37]) = (0:0:0, 0:0:0);
    (A2A1[25] => V[38]) = (0:0:0, 0:0:0);
    (A2A1[25] => V[39]) = (0:0:0, 0:0:0);
    (A2A1[25] => V[40]) = (0:0:0, 0:0:0);
    (A2A1[25] => V[41]) = (0:0:0, 0:0:0);
    (A2A1[25] => V[42]) = (0:0:0, 0:0:0);
    (A2A1[26] => AMULT26) = (0:0:0, 0:0:0);
    (A2A1[26] => U[27]) = (0:0:0, 0:0:0);
    (A2A1[26] => U[28]) = (0:0:0, 0:0:0);
    (A2A1[26] => U[29]) = (0:0:0, 0:0:0);
    (A2A1[26] => U[30]) = (0:0:0, 0:0:0);
    (A2A1[26] => U[31]) = (0:0:0, 0:0:0);
    (A2A1[26] => U[32]) = (0:0:0, 0:0:0);
    (A2A1[26] => U[33]) = (0:0:0, 0:0:0);
    (A2A1[26] => U[34]) = (0:0:0, 0:0:0);
    (A2A1[26] => U[35]) = (0:0:0, 0:0:0);
    (A2A1[26] => U[36]) = (0:0:0, 0:0:0);
    (A2A1[26] => U[37]) = (0:0:0, 0:0:0);
    (A2A1[26] => U[38]) = (0:0:0, 0:0:0);
    (A2A1[26] => U[39]) = (0:0:0, 0:0:0);
    (A2A1[26] => U[40]) = (0:0:0, 0:0:0);
    (A2A1[26] => U[41]) = (0:0:0, 0:0:0);
    (A2A1[26] => U[42]) = (0:0:0, 0:0:0);
    (A2A1[26] => U[43]) = (0:0:0, 0:0:0);
    (A2A1[26] => V[26]) = (0:0:0, 0:0:0);
    (A2A1[26] => V[27]) = (0:0:0, 0:0:0);
    (A2A1[26] => V[28]) = (0:0:0, 0:0:0);
    (A2A1[26] => V[29]) = (0:0:0, 0:0:0);
    (A2A1[26] => V[30]) = (0:0:0, 0:0:0);
    (A2A1[26] => V[31]) = (0:0:0, 0:0:0);
    (A2A1[26] => V[32]) = (0:0:0, 0:0:0);
    (A2A1[26] => V[33]) = (0:0:0, 0:0:0);
    (A2A1[26] => V[34]) = (0:0:0, 0:0:0);
    (A2A1[26] => V[35]) = (0:0:0, 0:0:0);
    (A2A1[26] => V[36]) = (0:0:0, 0:0:0);
    (A2A1[26] => V[37]) = (0:0:0, 0:0:0);
    (A2A1[26] => V[38]) = (0:0:0, 0:0:0);
    (A2A1[26] => V[39]) = (0:0:0, 0:0:0);
    (A2A1[26] => V[40]) = (0:0:0, 0:0:0);
    (A2A1[26] => V[41]) = (0:0:0, 0:0:0);
    (A2A1[26] => V[42]) = (0:0:0, 0:0:0);
    (A2A1[26] => V[43]) = (0:0:0, 0:0:0);
    (A2A1[2] => U[10]) = (0:0:0, 0:0:0);
    (A2A1[2] => U[11]) = (0:0:0, 0:0:0);
    (A2A1[2] => U[12]) = (0:0:0, 0:0:0);
    (A2A1[2] => U[13]) = (0:0:0, 0:0:0);
    (A2A1[2] => U[14]) = (0:0:0, 0:0:0);
    (A2A1[2] => U[15]) = (0:0:0, 0:0:0);
    (A2A1[2] => U[16]) = (0:0:0, 0:0:0);
    (A2A1[2] => U[17]) = (0:0:0, 0:0:0);
    (A2A1[2] => U[18]) = (0:0:0, 0:0:0);
    (A2A1[2] => U[19]) = (0:0:0, 0:0:0);
    (A2A1[2] => U[20]) = (0:0:0, 0:0:0);
    (A2A1[2] => U[21]) = (0:0:0, 0:0:0);
    (A2A1[2] => U[22]) = (0:0:0, 0:0:0);
    (A2A1[2] => U[23]) = (0:0:0, 0:0:0);
    (A2A1[2] => U[2]) = (0:0:0, 0:0:0);
    (A2A1[2] => U[3]) = (0:0:0, 0:0:0);
    (A2A1[2] => U[4]) = (0:0:0, 0:0:0);
    (A2A1[2] => U[5]) = (0:0:0, 0:0:0);
    (A2A1[2] => U[6]) = (0:0:0, 0:0:0);
    (A2A1[2] => U[7]) = (0:0:0, 0:0:0);
    (A2A1[2] => U[8]) = (0:0:0, 0:0:0);
    (A2A1[2] => U[9]) = (0:0:0, 0:0:0);
    (A2A1[2] => V[10]) = (0:0:0, 0:0:0);
    (A2A1[2] => V[11]) = (0:0:0, 0:0:0);
    (A2A1[2] => V[12]) = (0:0:0, 0:0:0);
    (A2A1[2] => V[13]) = (0:0:0, 0:0:0);
    (A2A1[2] => V[14]) = (0:0:0, 0:0:0);
    (A2A1[2] => V[15]) = (0:0:0, 0:0:0);
    (A2A1[2] => V[16]) = (0:0:0, 0:0:0);
    (A2A1[2] => V[17]) = (0:0:0, 0:0:0);
    (A2A1[2] => V[18]) = (0:0:0, 0:0:0);
    (A2A1[2] => V[19]) = (0:0:0, 0:0:0);
    (A2A1[2] => V[20]) = (0:0:0, 0:0:0);
    (A2A1[2] => V[21]) = (0:0:0, 0:0:0);
    (A2A1[2] => V[22]) = (0:0:0, 0:0:0);
    (A2A1[2] => V[4]) = (0:0:0, 0:0:0);
    (A2A1[2] => V[5]) = (0:0:0, 0:0:0);
    (A2A1[2] => V[6]) = (0:0:0, 0:0:0);
    (A2A1[2] => V[7]) = (0:0:0, 0:0:0);
    (A2A1[2] => V[8]) = (0:0:0, 0:0:0);
    (A2A1[2] => V[9]) = (0:0:0, 0:0:0);
    (A2A1[3] => U[10]) = (0:0:0, 0:0:0);
    (A2A1[3] => U[11]) = (0:0:0, 0:0:0);
    (A2A1[3] => U[12]) = (0:0:0, 0:0:0);
    (A2A1[3] => U[13]) = (0:0:0, 0:0:0);
    (A2A1[3] => U[14]) = (0:0:0, 0:0:0);
    (A2A1[3] => U[15]) = (0:0:0, 0:0:0);
    (A2A1[3] => U[16]) = (0:0:0, 0:0:0);
    (A2A1[3] => U[17]) = (0:0:0, 0:0:0);
    (A2A1[3] => U[18]) = (0:0:0, 0:0:0);
    (A2A1[3] => U[19]) = (0:0:0, 0:0:0);
    (A2A1[3] => U[20]) = (0:0:0, 0:0:0);
    (A2A1[3] => U[21]) = (0:0:0, 0:0:0);
    (A2A1[3] => U[22]) = (0:0:0, 0:0:0);
    (A2A1[3] => U[23]) = (0:0:0, 0:0:0);
    (A2A1[3] => U[24]) = (0:0:0, 0:0:0);
    (A2A1[3] => U[3]) = (0:0:0, 0:0:0);
    (A2A1[3] => U[4]) = (0:0:0, 0:0:0);
    (A2A1[3] => U[5]) = (0:0:0, 0:0:0);
    (A2A1[3] => U[6]) = (0:0:0, 0:0:0);
    (A2A1[3] => U[7]) = (0:0:0, 0:0:0);
    (A2A1[3] => U[8]) = (0:0:0, 0:0:0);
    (A2A1[3] => U[9]) = (0:0:0, 0:0:0);
    (A2A1[3] => V[10]) = (0:0:0, 0:0:0);
    (A2A1[3] => V[11]) = (0:0:0, 0:0:0);
    (A2A1[3] => V[12]) = (0:0:0, 0:0:0);
    (A2A1[3] => V[13]) = (0:0:0, 0:0:0);
    (A2A1[3] => V[14]) = (0:0:0, 0:0:0);
    (A2A1[3] => V[15]) = (0:0:0, 0:0:0);
    (A2A1[3] => V[16]) = (0:0:0, 0:0:0);
    (A2A1[3] => V[17]) = (0:0:0, 0:0:0);
    (A2A1[3] => V[18]) = (0:0:0, 0:0:0);
    (A2A1[3] => V[19]) = (0:0:0, 0:0:0);
    (A2A1[3] => V[20]) = (0:0:0, 0:0:0);
    (A2A1[3] => V[21]) = (0:0:0, 0:0:0);
    (A2A1[3] => V[22]) = (0:0:0, 0:0:0);
    (A2A1[3] => V[23]) = (0:0:0, 0:0:0);
    (A2A1[3] => V[4]) = (0:0:0, 0:0:0);
    (A2A1[3] => V[5]) = (0:0:0, 0:0:0);
    (A2A1[3] => V[6]) = (0:0:0, 0:0:0);
    (A2A1[3] => V[7]) = (0:0:0, 0:0:0);
    (A2A1[3] => V[8]) = (0:0:0, 0:0:0);
    (A2A1[3] => V[9]) = (0:0:0, 0:0:0);
    (A2A1[4] => U[10]) = (0:0:0, 0:0:0);
    (A2A1[4] => U[11]) = (0:0:0, 0:0:0);
    (A2A1[4] => U[12]) = (0:0:0, 0:0:0);
    (A2A1[4] => U[13]) = (0:0:0, 0:0:0);
    (A2A1[4] => U[14]) = (0:0:0, 0:0:0);
    (A2A1[4] => U[15]) = (0:0:0, 0:0:0);
    (A2A1[4] => U[16]) = (0:0:0, 0:0:0);
    (A2A1[4] => U[17]) = (0:0:0, 0:0:0);
    (A2A1[4] => U[18]) = (0:0:0, 0:0:0);
    (A2A1[4] => U[19]) = (0:0:0, 0:0:0);
    (A2A1[4] => U[20]) = (0:0:0, 0:0:0);
    (A2A1[4] => U[21]) = (0:0:0, 0:0:0);
    (A2A1[4] => U[22]) = (0:0:0, 0:0:0);
    (A2A1[4] => U[23]) = (0:0:0, 0:0:0);
    (A2A1[4] => U[24]) = (0:0:0, 0:0:0);
    (A2A1[4] => U[25]) = (0:0:0, 0:0:0);
    (A2A1[4] => U[5]) = (0:0:0, 0:0:0);
    (A2A1[4] => U[6]) = (0:0:0, 0:0:0);
    (A2A1[4] => U[7]) = (0:0:0, 0:0:0);
    (A2A1[4] => U[8]) = (0:0:0, 0:0:0);
    (A2A1[4] => U[9]) = (0:0:0, 0:0:0);
    (A2A1[4] => V[10]) = (0:0:0, 0:0:0);
    (A2A1[4] => V[11]) = (0:0:0, 0:0:0);
    (A2A1[4] => V[12]) = (0:0:0, 0:0:0);
    (A2A1[4] => V[13]) = (0:0:0, 0:0:0);
    (A2A1[4] => V[14]) = (0:0:0, 0:0:0);
    (A2A1[4] => V[15]) = (0:0:0, 0:0:0);
    (A2A1[4] => V[16]) = (0:0:0, 0:0:0);
    (A2A1[4] => V[17]) = (0:0:0, 0:0:0);
    (A2A1[4] => V[18]) = (0:0:0, 0:0:0);
    (A2A1[4] => V[19]) = (0:0:0, 0:0:0);
    (A2A1[4] => V[20]) = (0:0:0, 0:0:0);
    (A2A1[4] => V[21]) = (0:0:0, 0:0:0);
    (A2A1[4] => V[22]) = (0:0:0, 0:0:0);
    (A2A1[4] => V[23]) = (0:0:0, 0:0:0);
    (A2A1[4] => V[24]) = (0:0:0, 0:0:0);
    (A2A1[4] => V[4]) = (0:0:0, 0:0:0);
    (A2A1[4] => V[5]) = (0:0:0, 0:0:0);
    (A2A1[4] => V[6]) = (0:0:0, 0:0:0);
    (A2A1[4] => V[7]) = (0:0:0, 0:0:0);
    (A2A1[4] => V[8]) = (0:0:0, 0:0:0);
    (A2A1[4] => V[9]) = (0:0:0, 0:0:0);
    (A2A1[5] => U[10]) = (0:0:0, 0:0:0);
    (A2A1[5] => U[11]) = (0:0:0, 0:0:0);
    (A2A1[5] => U[12]) = (0:0:0, 0:0:0);
    (A2A1[5] => U[13]) = (0:0:0, 0:0:0);
    (A2A1[5] => U[14]) = (0:0:0, 0:0:0);
    (A2A1[5] => U[15]) = (0:0:0, 0:0:0);
    (A2A1[5] => U[16]) = (0:0:0, 0:0:0);
    (A2A1[5] => U[17]) = (0:0:0, 0:0:0);
    (A2A1[5] => U[18]) = (0:0:0, 0:0:0);
    (A2A1[5] => U[19]) = (0:0:0, 0:0:0);
    (A2A1[5] => U[20]) = (0:0:0, 0:0:0);
    (A2A1[5] => U[21]) = (0:0:0, 0:0:0);
    (A2A1[5] => U[22]) = (0:0:0, 0:0:0);
    (A2A1[5] => U[23]) = (0:0:0, 0:0:0);
    (A2A1[5] => U[24]) = (0:0:0, 0:0:0);
    (A2A1[5] => U[25]) = (0:0:0, 0:0:0);
    (A2A1[5] => U[26]) = (0:0:0, 0:0:0);
    (A2A1[5] => U[6]) = (0:0:0, 0:0:0);
    (A2A1[5] => U[7]) = (0:0:0, 0:0:0);
    (A2A1[5] => U[8]) = (0:0:0, 0:0:0);
    (A2A1[5] => U[9]) = (0:0:0, 0:0:0);
    (A2A1[5] => V[10]) = (0:0:0, 0:0:0);
    (A2A1[5] => V[11]) = (0:0:0, 0:0:0);
    (A2A1[5] => V[12]) = (0:0:0, 0:0:0);
    (A2A1[5] => V[13]) = (0:0:0, 0:0:0);
    (A2A1[5] => V[14]) = (0:0:0, 0:0:0);
    (A2A1[5] => V[15]) = (0:0:0, 0:0:0);
    (A2A1[5] => V[16]) = (0:0:0, 0:0:0);
    (A2A1[5] => V[17]) = (0:0:0, 0:0:0);
    (A2A1[5] => V[18]) = (0:0:0, 0:0:0);
    (A2A1[5] => V[19]) = (0:0:0, 0:0:0);
    (A2A1[5] => V[20]) = (0:0:0, 0:0:0);
    (A2A1[5] => V[21]) = (0:0:0, 0:0:0);
    (A2A1[5] => V[22]) = (0:0:0, 0:0:0);
    (A2A1[5] => V[23]) = (0:0:0, 0:0:0);
    (A2A1[5] => V[24]) = (0:0:0, 0:0:0);
    (A2A1[5] => V[25]) = (0:0:0, 0:0:0);
    (A2A1[5] => V[5]) = (0:0:0, 0:0:0);
    (A2A1[5] => V[6]) = (0:0:0, 0:0:0);
    (A2A1[5] => V[7]) = (0:0:0, 0:0:0);
    (A2A1[5] => V[8]) = (0:0:0, 0:0:0);
    (A2A1[5] => V[9]) = (0:0:0, 0:0:0);
    (A2A1[6] => U[10]) = (0:0:0, 0:0:0);
    (A2A1[6] => U[11]) = (0:0:0, 0:0:0);
    (A2A1[6] => U[12]) = (0:0:0, 0:0:0);
    (A2A1[6] => U[13]) = (0:0:0, 0:0:0);
    (A2A1[6] => U[14]) = (0:0:0, 0:0:0);
    (A2A1[6] => U[15]) = (0:0:0, 0:0:0);
    (A2A1[6] => U[16]) = (0:0:0, 0:0:0);
    (A2A1[6] => U[17]) = (0:0:0, 0:0:0);
    (A2A1[6] => U[18]) = (0:0:0, 0:0:0);
    (A2A1[6] => U[19]) = (0:0:0, 0:0:0);
    (A2A1[6] => U[20]) = (0:0:0, 0:0:0);
    (A2A1[6] => U[21]) = (0:0:0, 0:0:0);
    (A2A1[6] => U[22]) = (0:0:0, 0:0:0);
    (A2A1[6] => U[23]) = (0:0:0, 0:0:0);
    (A2A1[6] => U[24]) = (0:0:0, 0:0:0);
    (A2A1[6] => U[25]) = (0:0:0, 0:0:0);
    (A2A1[6] => U[26]) = (0:0:0, 0:0:0);
    (A2A1[6] => U[27]) = (0:0:0, 0:0:0);
    (A2A1[6] => U[7]) = (0:0:0, 0:0:0);
    (A2A1[6] => U[8]) = (0:0:0, 0:0:0);
    (A2A1[6] => U[9]) = (0:0:0, 0:0:0);
    (A2A1[6] => V[10]) = (0:0:0, 0:0:0);
    (A2A1[6] => V[11]) = (0:0:0, 0:0:0);
    (A2A1[6] => V[12]) = (0:0:0, 0:0:0);
    (A2A1[6] => V[13]) = (0:0:0, 0:0:0);
    (A2A1[6] => V[14]) = (0:0:0, 0:0:0);
    (A2A1[6] => V[15]) = (0:0:0, 0:0:0);
    (A2A1[6] => V[16]) = (0:0:0, 0:0:0);
    (A2A1[6] => V[17]) = (0:0:0, 0:0:0);
    (A2A1[6] => V[18]) = (0:0:0, 0:0:0);
    (A2A1[6] => V[19]) = (0:0:0, 0:0:0);
    (A2A1[6] => V[20]) = (0:0:0, 0:0:0);
    (A2A1[6] => V[21]) = (0:0:0, 0:0:0);
    (A2A1[6] => V[22]) = (0:0:0, 0:0:0);
    (A2A1[6] => V[23]) = (0:0:0, 0:0:0);
    (A2A1[6] => V[24]) = (0:0:0, 0:0:0);
    (A2A1[6] => V[25]) = (0:0:0, 0:0:0);
    (A2A1[6] => V[26]) = (0:0:0, 0:0:0);
    (A2A1[6] => V[6]) = (0:0:0, 0:0:0);
    (A2A1[6] => V[7]) = (0:0:0, 0:0:0);
    (A2A1[6] => V[8]) = (0:0:0, 0:0:0);
    (A2A1[6] => V[9]) = (0:0:0, 0:0:0);
    (A2A1[7] => U[10]) = (0:0:0, 0:0:0);
    (A2A1[7] => U[11]) = (0:0:0, 0:0:0);
    (A2A1[7] => U[12]) = (0:0:0, 0:0:0);
    (A2A1[7] => U[13]) = (0:0:0, 0:0:0);
    (A2A1[7] => U[14]) = (0:0:0, 0:0:0);
    (A2A1[7] => U[15]) = (0:0:0, 0:0:0);
    (A2A1[7] => U[16]) = (0:0:0, 0:0:0);
    (A2A1[7] => U[17]) = (0:0:0, 0:0:0);
    (A2A1[7] => U[18]) = (0:0:0, 0:0:0);
    (A2A1[7] => U[19]) = (0:0:0, 0:0:0);
    (A2A1[7] => U[20]) = (0:0:0, 0:0:0);
    (A2A1[7] => U[21]) = (0:0:0, 0:0:0);
    (A2A1[7] => U[22]) = (0:0:0, 0:0:0);
    (A2A1[7] => U[23]) = (0:0:0, 0:0:0);
    (A2A1[7] => U[24]) = (0:0:0, 0:0:0);
    (A2A1[7] => U[25]) = (0:0:0, 0:0:0);
    (A2A1[7] => U[26]) = (0:0:0, 0:0:0);
    (A2A1[7] => U[27]) = (0:0:0, 0:0:0);
    (A2A1[7] => U[28]) = (0:0:0, 0:0:0);
    (A2A1[7] => U[8]) = (0:0:0, 0:0:0);
    (A2A1[7] => U[9]) = (0:0:0, 0:0:0);
    (A2A1[7] => V[10]) = (0:0:0, 0:0:0);
    (A2A1[7] => V[11]) = (0:0:0, 0:0:0);
    (A2A1[7] => V[12]) = (0:0:0, 0:0:0);
    (A2A1[7] => V[13]) = (0:0:0, 0:0:0);
    (A2A1[7] => V[14]) = (0:0:0, 0:0:0);
    (A2A1[7] => V[15]) = (0:0:0, 0:0:0);
    (A2A1[7] => V[16]) = (0:0:0, 0:0:0);
    (A2A1[7] => V[17]) = (0:0:0, 0:0:0);
    (A2A1[7] => V[18]) = (0:0:0, 0:0:0);
    (A2A1[7] => V[19]) = (0:0:0, 0:0:0);
    (A2A1[7] => V[20]) = (0:0:0, 0:0:0);
    (A2A1[7] => V[21]) = (0:0:0, 0:0:0);
    (A2A1[7] => V[22]) = (0:0:0, 0:0:0);
    (A2A1[7] => V[23]) = (0:0:0, 0:0:0);
    (A2A1[7] => V[24]) = (0:0:0, 0:0:0);
    (A2A1[7] => V[25]) = (0:0:0, 0:0:0);
    (A2A1[7] => V[26]) = (0:0:0, 0:0:0);
    (A2A1[7] => V[27]) = (0:0:0, 0:0:0);
    (A2A1[7] => V[7]) = (0:0:0, 0:0:0);
    (A2A1[7] => V[8]) = (0:0:0, 0:0:0);
    (A2A1[7] => V[9]) = (0:0:0, 0:0:0);
    (A2A1[8] => U[10]) = (0:0:0, 0:0:0);
    (A2A1[8] => U[11]) = (0:0:0, 0:0:0);
    (A2A1[8] => U[12]) = (0:0:0, 0:0:0);
    (A2A1[8] => U[13]) = (0:0:0, 0:0:0);
    (A2A1[8] => U[14]) = (0:0:0, 0:0:0);
    (A2A1[8] => U[15]) = (0:0:0, 0:0:0);
    (A2A1[8] => U[16]) = (0:0:0, 0:0:0);
    (A2A1[8] => U[17]) = (0:0:0, 0:0:0);
    (A2A1[8] => U[18]) = (0:0:0, 0:0:0);
    (A2A1[8] => U[19]) = (0:0:0, 0:0:0);
    (A2A1[8] => U[20]) = (0:0:0, 0:0:0);
    (A2A1[8] => U[21]) = (0:0:0, 0:0:0);
    (A2A1[8] => U[22]) = (0:0:0, 0:0:0);
    (A2A1[8] => U[23]) = (0:0:0, 0:0:0);
    (A2A1[8] => U[24]) = (0:0:0, 0:0:0);
    (A2A1[8] => U[25]) = (0:0:0, 0:0:0);
    (A2A1[8] => U[26]) = (0:0:0, 0:0:0);
    (A2A1[8] => U[27]) = (0:0:0, 0:0:0);
    (A2A1[8] => U[28]) = (0:0:0, 0:0:0);
    (A2A1[8] => U[29]) = (0:0:0, 0:0:0);
    (A2A1[8] => U[9]) = (0:0:0, 0:0:0);
    (A2A1[8] => V[10]) = (0:0:0, 0:0:0);
    (A2A1[8] => V[11]) = (0:0:0, 0:0:0);
    (A2A1[8] => V[12]) = (0:0:0, 0:0:0);
    (A2A1[8] => V[13]) = (0:0:0, 0:0:0);
    (A2A1[8] => V[14]) = (0:0:0, 0:0:0);
    (A2A1[8] => V[15]) = (0:0:0, 0:0:0);
    (A2A1[8] => V[16]) = (0:0:0, 0:0:0);
    (A2A1[8] => V[17]) = (0:0:0, 0:0:0);
    (A2A1[8] => V[18]) = (0:0:0, 0:0:0);
    (A2A1[8] => V[19]) = (0:0:0, 0:0:0);
    (A2A1[8] => V[20]) = (0:0:0, 0:0:0);
    (A2A1[8] => V[21]) = (0:0:0, 0:0:0);
    (A2A1[8] => V[22]) = (0:0:0, 0:0:0);
    (A2A1[8] => V[23]) = (0:0:0, 0:0:0);
    (A2A1[8] => V[24]) = (0:0:0, 0:0:0);
    (A2A1[8] => V[25]) = (0:0:0, 0:0:0);
    (A2A1[8] => V[26]) = (0:0:0, 0:0:0);
    (A2A1[8] => V[27]) = (0:0:0, 0:0:0);
    (A2A1[8] => V[28]) = (0:0:0, 0:0:0);
    (A2A1[8] => V[8]) = (0:0:0, 0:0:0);
    (A2A1[8] => V[9]) = (0:0:0, 0:0:0);
    (A2A1[9] => U[10]) = (0:0:0, 0:0:0);
    (A2A1[9] => U[11]) = (0:0:0, 0:0:0);
    (A2A1[9] => U[12]) = (0:0:0, 0:0:0);
    (A2A1[9] => U[13]) = (0:0:0, 0:0:0);
    (A2A1[9] => U[14]) = (0:0:0, 0:0:0);
    (A2A1[9] => U[15]) = (0:0:0, 0:0:0);
    (A2A1[9] => U[16]) = (0:0:0, 0:0:0);
    (A2A1[9] => U[17]) = (0:0:0, 0:0:0);
    (A2A1[9] => U[18]) = (0:0:0, 0:0:0);
    (A2A1[9] => U[19]) = (0:0:0, 0:0:0);
    (A2A1[9] => U[20]) = (0:0:0, 0:0:0);
    (A2A1[9] => U[21]) = (0:0:0, 0:0:0);
    (A2A1[9] => U[22]) = (0:0:0, 0:0:0);
    (A2A1[9] => U[23]) = (0:0:0, 0:0:0);
    (A2A1[9] => U[24]) = (0:0:0, 0:0:0);
    (A2A1[9] => U[25]) = (0:0:0, 0:0:0);
    (A2A1[9] => U[26]) = (0:0:0, 0:0:0);
    (A2A1[9] => U[27]) = (0:0:0, 0:0:0);
    (A2A1[9] => U[28]) = (0:0:0, 0:0:0);
    (A2A1[9] => U[29]) = (0:0:0, 0:0:0);
    (A2A1[9] => U[30]) = (0:0:0, 0:0:0);
    (A2A1[9] => V[10]) = (0:0:0, 0:0:0);
    (A2A1[9] => V[11]) = (0:0:0, 0:0:0);
    (A2A1[9] => V[12]) = (0:0:0, 0:0:0);
    (A2A1[9] => V[13]) = (0:0:0, 0:0:0);
    (A2A1[9] => V[14]) = (0:0:0, 0:0:0);
    (A2A1[9] => V[15]) = (0:0:0, 0:0:0);
    (A2A1[9] => V[16]) = (0:0:0, 0:0:0);
    (A2A1[9] => V[17]) = (0:0:0, 0:0:0);
    (A2A1[9] => V[18]) = (0:0:0, 0:0:0);
    (A2A1[9] => V[19]) = (0:0:0, 0:0:0);
    (A2A1[9] => V[20]) = (0:0:0, 0:0:0);
    (A2A1[9] => V[21]) = (0:0:0, 0:0:0);
    (A2A1[9] => V[22]) = (0:0:0, 0:0:0);
    (A2A1[9] => V[23]) = (0:0:0, 0:0:0);
    (A2A1[9] => V[24]) = (0:0:0, 0:0:0);
    (A2A1[9] => V[25]) = (0:0:0, 0:0:0);
    (A2A1[9] => V[26]) = (0:0:0, 0:0:0);
    (A2A1[9] => V[27]) = (0:0:0, 0:0:0);
    (A2A1[9] => V[28]) = (0:0:0, 0:0:0);
    (A2A1[9] => V[29]) = (0:0:0, 0:0:0);
    (A2A1[9] => V[9]) = (0:0:0, 0:0:0);
    (AD_DATA[0] => U[10]) = (0:0:0, 0:0:0);
    (AD_DATA[0] => U[11]) = (0:0:0, 0:0:0);
    (AD_DATA[0] => U[12]) = (0:0:0, 0:0:0);
    (AD_DATA[0] => U[13]) = (0:0:0, 0:0:0);
    (AD_DATA[0] => U[14]) = (0:0:0, 0:0:0);
    (AD_DATA[0] => U[15]) = (0:0:0, 0:0:0);
    (AD_DATA[0] => U[16]) = (0:0:0, 0:0:0);
    (AD_DATA[0] => U[17]) = (0:0:0, 0:0:0);
    (AD_DATA[0] => U[18]) = (0:0:0, 0:0:0);
    (AD_DATA[0] => U[19]) = (0:0:0, 0:0:0);
    (AD_DATA[0] => U[1]) = (0:0:0, 0:0:0);
    (AD_DATA[0] => U[20]) = (0:0:0, 0:0:0);
    (AD_DATA[0] => U[21]) = (0:0:0, 0:0:0);
    (AD_DATA[0] => U[22]) = (0:0:0, 0:0:0);
    (AD_DATA[0] => U[23]) = (0:0:0, 0:0:0);
    (AD_DATA[0] => U[24]) = (0:0:0, 0:0:0);
    (AD_DATA[0] => U[25]) = (0:0:0, 0:0:0);
    (AD_DATA[0] => U[26]) = (0:0:0, 0:0:0);
    (AD_DATA[0] => U[27]) = (0:0:0, 0:0:0);
    (AD_DATA[0] => U[28]) = (0:0:0, 0:0:0);
    (AD_DATA[0] => U[29]) = (0:0:0, 0:0:0);
    (AD_DATA[0] => U[2]) = (0:0:0, 0:0:0);
    (AD_DATA[0] => U[30]) = (0:0:0, 0:0:0);
    (AD_DATA[0] => U[31]) = (0:0:0, 0:0:0);
    (AD_DATA[0] => U[3]) = (0:0:0, 0:0:0);
    (AD_DATA[0] => U[4]) = (0:0:0, 0:0:0);
    (AD_DATA[0] => U[5]) = (0:0:0, 0:0:0);
    (AD_DATA[0] => U[6]) = (0:0:0, 0:0:0);
    (AD_DATA[0] => U[7]) = (0:0:0, 0:0:0);
    (AD_DATA[0] => U[8]) = (0:0:0, 0:0:0);
    (AD_DATA[0] => U[9]) = (0:0:0, 0:0:0);
    (AD_DATA[0] => V[0]) = (0:0:0, 0:0:0);
    (AD_DATA[0] => V[10]) = (0:0:0, 0:0:0);
    (AD_DATA[0] => V[11]) = (0:0:0, 0:0:0);
    (AD_DATA[0] => V[12]) = (0:0:0, 0:0:0);
    (AD_DATA[0] => V[13]) = (0:0:0, 0:0:0);
    (AD_DATA[0] => V[14]) = (0:0:0, 0:0:0);
    (AD_DATA[0] => V[15]) = (0:0:0, 0:0:0);
    (AD_DATA[0] => V[16]) = (0:0:0, 0:0:0);
    (AD_DATA[0] => V[17]) = (0:0:0, 0:0:0);
    (AD_DATA[0] => V[18]) = (0:0:0, 0:0:0);
    (AD_DATA[0] => V[19]) = (0:0:0, 0:0:0);
    (AD_DATA[0] => V[20]) = (0:0:0, 0:0:0);
    (AD_DATA[0] => V[21]) = (0:0:0, 0:0:0);
    (AD_DATA[0] => V[22]) = (0:0:0, 0:0:0);
    (AD_DATA[0] => V[23]) = (0:0:0, 0:0:0);
    (AD_DATA[0] => V[24]) = (0:0:0, 0:0:0);
    (AD_DATA[0] => V[25]) = (0:0:0, 0:0:0);
    (AD_DATA[0] => V[26]) = (0:0:0, 0:0:0);
    (AD_DATA[0] => V[27]) = (0:0:0, 0:0:0);
    (AD_DATA[0] => V[28]) = (0:0:0, 0:0:0);
    (AD_DATA[0] => V[29]) = (0:0:0, 0:0:0);
    (AD_DATA[0] => V[30]) = (0:0:0, 0:0:0);
    (AD_DATA[0] => V[4]) = (0:0:0, 0:0:0);
    (AD_DATA[0] => V[5]) = (0:0:0, 0:0:0);
    (AD_DATA[0] => V[6]) = (0:0:0, 0:0:0);
    (AD_DATA[0] => V[7]) = (0:0:0, 0:0:0);
    (AD_DATA[0] => V[8]) = (0:0:0, 0:0:0);
    (AD_DATA[0] => V[9]) = (0:0:0, 0:0:0);
    (AD_DATA[10] => U[11]) = (0:0:0, 0:0:0);
    (AD_DATA[10] => U[12]) = (0:0:0, 0:0:0);
    (AD_DATA[10] => U[13]) = (0:0:0, 0:0:0);
    (AD_DATA[10] => U[14]) = (0:0:0, 0:0:0);
    (AD_DATA[10] => U[15]) = (0:0:0, 0:0:0);
    (AD_DATA[10] => U[16]) = (0:0:0, 0:0:0);
    (AD_DATA[10] => U[17]) = (0:0:0, 0:0:0);
    (AD_DATA[10] => U[18]) = (0:0:0, 0:0:0);
    (AD_DATA[10] => U[19]) = (0:0:0, 0:0:0);
    (AD_DATA[10] => U[20]) = (0:0:0, 0:0:0);
    (AD_DATA[10] => U[21]) = (0:0:0, 0:0:0);
    (AD_DATA[10] => U[22]) = (0:0:0, 0:0:0);
    (AD_DATA[10] => U[23]) = (0:0:0, 0:0:0);
    (AD_DATA[10] => U[24]) = (0:0:0, 0:0:0);
    (AD_DATA[10] => U[25]) = (0:0:0, 0:0:0);
    (AD_DATA[10] => U[26]) = (0:0:0, 0:0:0);
    (AD_DATA[10] => U[27]) = (0:0:0, 0:0:0);
    (AD_DATA[10] => U[28]) = (0:0:0, 0:0:0);
    (AD_DATA[10] => U[29]) = (0:0:0, 0:0:0);
    (AD_DATA[10] => U[30]) = (0:0:0, 0:0:0);
    (AD_DATA[10] => U[31]) = (0:0:0, 0:0:0);
    (AD_DATA[10] => U[32]) = (0:0:0, 0:0:0);
    (AD_DATA[10] => U[33]) = (0:0:0, 0:0:0);
    (AD_DATA[10] => U[34]) = (0:0:0, 0:0:0);
    (AD_DATA[10] => U[35]) = (0:0:0, 0:0:0);
    (AD_DATA[10] => U[36]) = (0:0:0, 0:0:0);
    (AD_DATA[10] => U[37]) = (0:0:0, 0:0:0);
    (AD_DATA[10] => U[38]) = (0:0:0, 0:0:0);
    (AD_DATA[10] => U[39]) = (0:0:0, 0:0:0);
    (AD_DATA[10] => U[40]) = (0:0:0, 0:0:0);
    (AD_DATA[10] => V[10]) = (0:0:0, 0:0:0);
    (AD_DATA[10] => V[11]) = (0:0:0, 0:0:0);
    (AD_DATA[10] => V[12]) = (0:0:0, 0:0:0);
    (AD_DATA[10] => V[13]) = (0:0:0, 0:0:0);
    (AD_DATA[10] => V[14]) = (0:0:0, 0:0:0);
    (AD_DATA[10] => V[15]) = (0:0:0, 0:0:0);
    (AD_DATA[10] => V[16]) = (0:0:0, 0:0:0);
    (AD_DATA[10] => V[17]) = (0:0:0, 0:0:0);
    (AD_DATA[10] => V[18]) = (0:0:0, 0:0:0);
    (AD_DATA[10] => V[19]) = (0:0:0, 0:0:0);
    (AD_DATA[10] => V[20]) = (0:0:0, 0:0:0);
    (AD_DATA[10] => V[21]) = (0:0:0, 0:0:0);
    (AD_DATA[10] => V[22]) = (0:0:0, 0:0:0);
    (AD_DATA[10] => V[23]) = (0:0:0, 0:0:0);
    (AD_DATA[10] => V[24]) = (0:0:0, 0:0:0);
    (AD_DATA[10] => V[25]) = (0:0:0, 0:0:0);
    (AD_DATA[10] => V[26]) = (0:0:0, 0:0:0);
    (AD_DATA[10] => V[27]) = (0:0:0, 0:0:0);
    (AD_DATA[10] => V[28]) = (0:0:0, 0:0:0);
    (AD_DATA[10] => V[29]) = (0:0:0, 0:0:0);
    (AD_DATA[10] => V[30]) = (0:0:0, 0:0:0);
    (AD_DATA[10] => V[31]) = (0:0:0, 0:0:0);
    (AD_DATA[10] => V[32]) = (0:0:0, 0:0:0);
    (AD_DATA[10] => V[33]) = (0:0:0, 0:0:0);
    (AD_DATA[10] => V[34]) = (0:0:0, 0:0:0);
    (AD_DATA[10] => V[35]) = (0:0:0, 0:0:0);
    (AD_DATA[10] => V[36]) = (0:0:0, 0:0:0);
    (AD_DATA[10] => V[37]) = (0:0:0, 0:0:0);
    (AD_DATA[10] => V[38]) = (0:0:0, 0:0:0);
    (AD_DATA[10] => V[39]) = (0:0:0, 0:0:0);
    (AD_DATA[11] => U[11]) = (0:0:0, 0:0:0);
    (AD_DATA[11] => U[12]) = (0:0:0, 0:0:0);
    (AD_DATA[11] => U[13]) = (0:0:0, 0:0:0);
    (AD_DATA[11] => U[14]) = (0:0:0, 0:0:0);
    (AD_DATA[11] => U[15]) = (0:0:0, 0:0:0);
    (AD_DATA[11] => U[16]) = (0:0:0, 0:0:0);
    (AD_DATA[11] => U[17]) = (0:0:0, 0:0:0);
    (AD_DATA[11] => U[18]) = (0:0:0, 0:0:0);
    (AD_DATA[11] => U[19]) = (0:0:0, 0:0:0);
    (AD_DATA[11] => U[20]) = (0:0:0, 0:0:0);
    (AD_DATA[11] => U[21]) = (0:0:0, 0:0:0);
    (AD_DATA[11] => U[22]) = (0:0:0, 0:0:0);
    (AD_DATA[11] => U[23]) = (0:0:0, 0:0:0);
    (AD_DATA[11] => U[24]) = (0:0:0, 0:0:0);
    (AD_DATA[11] => U[25]) = (0:0:0, 0:0:0);
    (AD_DATA[11] => U[26]) = (0:0:0, 0:0:0);
    (AD_DATA[11] => U[27]) = (0:0:0, 0:0:0);
    (AD_DATA[11] => U[28]) = (0:0:0, 0:0:0);
    (AD_DATA[11] => U[29]) = (0:0:0, 0:0:0);
    (AD_DATA[11] => U[30]) = (0:0:0, 0:0:0);
    (AD_DATA[11] => U[31]) = (0:0:0, 0:0:0);
    (AD_DATA[11] => U[32]) = (0:0:0, 0:0:0);
    (AD_DATA[11] => U[33]) = (0:0:0, 0:0:0);
    (AD_DATA[11] => U[34]) = (0:0:0, 0:0:0);
    (AD_DATA[11] => U[35]) = (0:0:0, 0:0:0);
    (AD_DATA[11] => U[36]) = (0:0:0, 0:0:0);
    (AD_DATA[11] => U[37]) = (0:0:0, 0:0:0);
    (AD_DATA[11] => U[38]) = (0:0:0, 0:0:0);
    (AD_DATA[11] => U[39]) = (0:0:0, 0:0:0);
    (AD_DATA[11] => U[40]) = (0:0:0, 0:0:0);
    (AD_DATA[11] => U[41]) = (0:0:0, 0:0:0);
    (AD_DATA[11] => V[10]) = (0:0:0, 0:0:0);
    (AD_DATA[11] => V[11]) = (0:0:0, 0:0:0);
    (AD_DATA[11] => V[12]) = (0:0:0, 0:0:0);
    (AD_DATA[11] => V[13]) = (0:0:0, 0:0:0);
    (AD_DATA[11] => V[14]) = (0:0:0, 0:0:0);
    (AD_DATA[11] => V[15]) = (0:0:0, 0:0:0);
    (AD_DATA[11] => V[16]) = (0:0:0, 0:0:0);
    (AD_DATA[11] => V[17]) = (0:0:0, 0:0:0);
    (AD_DATA[11] => V[18]) = (0:0:0, 0:0:0);
    (AD_DATA[11] => V[19]) = (0:0:0, 0:0:0);
    (AD_DATA[11] => V[20]) = (0:0:0, 0:0:0);
    (AD_DATA[11] => V[21]) = (0:0:0, 0:0:0);
    (AD_DATA[11] => V[22]) = (0:0:0, 0:0:0);
    (AD_DATA[11] => V[23]) = (0:0:0, 0:0:0);
    (AD_DATA[11] => V[24]) = (0:0:0, 0:0:0);
    (AD_DATA[11] => V[25]) = (0:0:0, 0:0:0);
    (AD_DATA[11] => V[26]) = (0:0:0, 0:0:0);
    (AD_DATA[11] => V[27]) = (0:0:0, 0:0:0);
    (AD_DATA[11] => V[28]) = (0:0:0, 0:0:0);
    (AD_DATA[11] => V[29]) = (0:0:0, 0:0:0);
    (AD_DATA[11] => V[30]) = (0:0:0, 0:0:0);
    (AD_DATA[11] => V[31]) = (0:0:0, 0:0:0);
    (AD_DATA[11] => V[32]) = (0:0:0, 0:0:0);
    (AD_DATA[11] => V[33]) = (0:0:0, 0:0:0);
    (AD_DATA[11] => V[34]) = (0:0:0, 0:0:0);
    (AD_DATA[11] => V[35]) = (0:0:0, 0:0:0);
    (AD_DATA[11] => V[36]) = (0:0:0, 0:0:0);
    (AD_DATA[11] => V[37]) = (0:0:0, 0:0:0);
    (AD_DATA[11] => V[38]) = (0:0:0, 0:0:0);
    (AD_DATA[11] => V[39]) = (0:0:0, 0:0:0);
    (AD_DATA[11] => V[40]) = (0:0:0, 0:0:0);
    (AD_DATA[12] => U[13]) = (0:0:0, 0:0:0);
    (AD_DATA[12] => U[14]) = (0:0:0, 0:0:0);
    (AD_DATA[12] => U[15]) = (0:0:0, 0:0:0);
    (AD_DATA[12] => U[16]) = (0:0:0, 0:0:0);
    (AD_DATA[12] => U[17]) = (0:0:0, 0:0:0);
    (AD_DATA[12] => U[18]) = (0:0:0, 0:0:0);
    (AD_DATA[12] => U[19]) = (0:0:0, 0:0:0);
    (AD_DATA[12] => U[20]) = (0:0:0, 0:0:0);
    (AD_DATA[12] => U[21]) = (0:0:0, 0:0:0);
    (AD_DATA[12] => U[22]) = (0:0:0, 0:0:0);
    (AD_DATA[12] => U[23]) = (0:0:0, 0:0:0);
    (AD_DATA[12] => U[24]) = (0:0:0, 0:0:0);
    (AD_DATA[12] => U[25]) = (0:0:0, 0:0:0);
    (AD_DATA[12] => U[26]) = (0:0:0, 0:0:0);
    (AD_DATA[12] => U[27]) = (0:0:0, 0:0:0);
    (AD_DATA[12] => U[28]) = (0:0:0, 0:0:0);
    (AD_DATA[12] => U[29]) = (0:0:0, 0:0:0);
    (AD_DATA[12] => U[30]) = (0:0:0, 0:0:0);
    (AD_DATA[12] => U[31]) = (0:0:0, 0:0:0);
    (AD_DATA[12] => U[32]) = (0:0:0, 0:0:0);
    (AD_DATA[12] => U[33]) = (0:0:0, 0:0:0);
    (AD_DATA[12] => U[34]) = (0:0:0, 0:0:0);
    (AD_DATA[12] => U[35]) = (0:0:0, 0:0:0);
    (AD_DATA[12] => U[36]) = (0:0:0, 0:0:0);
    (AD_DATA[12] => U[37]) = (0:0:0, 0:0:0);
    (AD_DATA[12] => U[38]) = (0:0:0, 0:0:0);
    (AD_DATA[12] => U[39]) = (0:0:0, 0:0:0);
    (AD_DATA[12] => U[40]) = (0:0:0, 0:0:0);
    (AD_DATA[12] => U[41]) = (0:0:0, 0:0:0);
    (AD_DATA[12] => V[12]) = (0:0:0, 0:0:0);
    (AD_DATA[12] => V[13]) = (0:0:0, 0:0:0);
    (AD_DATA[12] => V[14]) = (0:0:0, 0:0:0);
    (AD_DATA[12] => V[15]) = (0:0:0, 0:0:0);
    (AD_DATA[12] => V[16]) = (0:0:0, 0:0:0);
    (AD_DATA[12] => V[17]) = (0:0:0, 0:0:0);
    (AD_DATA[12] => V[18]) = (0:0:0, 0:0:0);
    (AD_DATA[12] => V[19]) = (0:0:0, 0:0:0);
    (AD_DATA[12] => V[20]) = (0:0:0, 0:0:0);
    (AD_DATA[12] => V[21]) = (0:0:0, 0:0:0);
    (AD_DATA[12] => V[22]) = (0:0:0, 0:0:0);
    (AD_DATA[12] => V[23]) = (0:0:0, 0:0:0);
    (AD_DATA[12] => V[24]) = (0:0:0, 0:0:0);
    (AD_DATA[12] => V[25]) = (0:0:0, 0:0:0);
    (AD_DATA[12] => V[26]) = (0:0:0, 0:0:0);
    (AD_DATA[12] => V[27]) = (0:0:0, 0:0:0);
    (AD_DATA[12] => V[28]) = (0:0:0, 0:0:0);
    (AD_DATA[12] => V[29]) = (0:0:0, 0:0:0);
    (AD_DATA[12] => V[30]) = (0:0:0, 0:0:0);
    (AD_DATA[12] => V[31]) = (0:0:0, 0:0:0);
    (AD_DATA[12] => V[32]) = (0:0:0, 0:0:0);
    (AD_DATA[12] => V[33]) = (0:0:0, 0:0:0);
    (AD_DATA[12] => V[34]) = (0:0:0, 0:0:0);
    (AD_DATA[12] => V[35]) = (0:0:0, 0:0:0);
    (AD_DATA[12] => V[36]) = (0:0:0, 0:0:0);
    (AD_DATA[12] => V[37]) = (0:0:0, 0:0:0);
    (AD_DATA[12] => V[38]) = (0:0:0, 0:0:0);
    (AD_DATA[12] => V[39]) = (0:0:0, 0:0:0);
    (AD_DATA[12] => V[40]) = (0:0:0, 0:0:0);
    (AD_DATA[13] => U[13]) = (0:0:0, 0:0:0);
    (AD_DATA[13] => U[14]) = (0:0:0, 0:0:0);
    (AD_DATA[13] => U[15]) = (0:0:0, 0:0:0);
    (AD_DATA[13] => U[16]) = (0:0:0, 0:0:0);
    (AD_DATA[13] => U[17]) = (0:0:0, 0:0:0);
    (AD_DATA[13] => U[18]) = (0:0:0, 0:0:0);
    (AD_DATA[13] => U[19]) = (0:0:0, 0:0:0);
    (AD_DATA[13] => U[20]) = (0:0:0, 0:0:0);
    (AD_DATA[13] => U[21]) = (0:0:0, 0:0:0);
    (AD_DATA[13] => U[22]) = (0:0:0, 0:0:0);
    (AD_DATA[13] => U[23]) = (0:0:0, 0:0:0);
    (AD_DATA[13] => U[24]) = (0:0:0, 0:0:0);
    (AD_DATA[13] => U[25]) = (0:0:0, 0:0:0);
    (AD_DATA[13] => U[26]) = (0:0:0, 0:0:0);
    (AD_DATA[13] => U[27]) = (0:0:0, 0:0:0);
    (AD_DATA[13] => U[28]) = (0:0:0, 0:0:0);
    (AD_DATA[13] => U[29]) = (0:0:0, 0:0:0);
    (AD_DATA[13] => U[30]) = (0:0:0, 0:0:0);
    (AD_DATA[13] => U[31]) = (0:0:0, 0:0:0);
    (AD_DATA[13] => U[32]) = (0:0:0, 0:0:0);
    (AD_DATA[13] => U[33]) = (0:0:0, 0:0:0);
    (AD_DATA[13] => U[34]) = (0:0:0, 0:0:0);
    (AD_DATA[13] => U[35]) = (0:0:0, 0:0:0);
    (AD_DATA[13] => U[36]) = (0:0:0, 0:0:0);
    (AD_DATA[13] => U[37]) = (0:0:0, 0:0:0);
    (AD_DATA[13] => U[38]) = (0:0:0, 0:0:0);
    (AD_DATA[13] => U[39]) = (0:0:0, 0:0:0);
    (AD_DATA[13] => U[40]) = (0:0:0, 0:0:0);
    (AD_DATA[13] => U[41]) = (0:0:0, 0:0:0);
    (AD_DATA[13] => U[42]) = (0:0:0, 0:0:0);
    (AD_DATA[13] => V[12]) = (0:0:0, 0:0:0);
    (AD_DATA[13] => V[13]) = (0:0:0, 0:0:0);
    (AD_DATA[13] => V[14]) = (0:0:0, 0:0:0);
    (AD_DATA[13] => V[15]) = (0:0:0, 0:0:0);
    (AD_DATA[13] => V[16]) = (0:0:0, 0:0:0);
    (AD_DATA[13] => V[17]) = (0:0:0, 0:0:0);
    (AD_DATA[13] => V[18]) = (0:0:0, 0:0:0);
    (AD_DATA[13] => V[19]) = (0:0:0, 0:0:0);
    (AD_DATA[13] => V[20]) = (0:0:0, 0:0:0);
    (AD_DATA[13] => V[21]) = (0:0:0, 0:0:0);
    (AD_DATA[13] => V[22]) = (0:0:0, 0:0:0);
    (AD_DATA[13] => V[23]) = (0:0:0, 0:0:0);
    (AD_DATA[13] => V[24]) = (0:0:0, 0:0:0);
    (AD_DATA[13] => V[25]) = (0:0:0, 0:0:0);
    (AD_DATA[13] => V[26]) = (0:0:0, 0:0:0);
    (AD_DATA[13] => V[27]) = (0:0:0, 0:0:0);
    (AD_DATA[13] => V[28]) = (0:0:0, 0:0:0);
    (AD_DATA[13] => V[29]) = (0:0:0, 0:0:0);
    (AD_DATA[13] => V[30]) = (0:0:0, 0:0:0);
    (AD_DATA[13] => V[31]) = (0:0:0, 0:0:0);
    (AD_DATA[13] => V[32]) = (0:0:0, 0:0:0);
    (AD_DATA[13] => V[33]) = (0:0:0, 0:0:0);
    (AD_DATA[13] => V[34]) = (0:0:0, 0:0:0);
    (AD_DATA[13] => V[35]) = (0:0:0, 0:0:0);
    (AD_DATA[13] => V[36]) = (0:0:0, 0:0:0);
    (AD_DATA[13] => V[37]) = (0:0:0, 0:0:0);
    (AD_DATA[13] => V[38]) = (0:0:0, 0:0:0);
    (AD_DATA[13] => V[39]) = (0:0:0, 0:0:0);
    (AD_DATA[13] => V[40]) = (0:0:0, 0:0:0);
    (AD_DATA[13] => V[41]) = (0:0:0, 0:0:0);
    (AD_DATA[14] => U[15]) = (0:0:0, 0:0:0);
    (AD_DATA[14] => U[16]) = (0:0:0, 0:0:0);
    (AD_DATA[14] => U[17]) = (0:0:0, 0:0:0);
    (AD_DATA[14] => U[18]) = (0:0:0, 0:0:0);
    (AD_DATA[14] => U[19]) = (0:0:0, 0:0:0);
    (AD_DATA[14] => U[20]) = (0:0:0, 0:0:0);
    (AD_DATA[14] => U[21]) = (0:0:0, 0:0:0);
    (AD_DATA[14] => U[22]) = (0:0:0, 0:0:0);
    (AD_DATA[14] => U[23]) = (0:0:0, 0:0:0);
    (AD_DATA[14] => U[24]) = (0:0:0, 0:0:0);
    (AD_DATA[14] => U[25]) = (0:0:0, 0:0:0);
    (AD_DATA[14] => U[26]) = (0:0:0, 0:0:0);
    (AD_DATA[14] => U[27]) = (0:0:0, 0:0:0);
    (AD_DATA[14] => U[28]) = (0:0:0, 0:0:0);
    (AD_DATA[14] => U[29]) = (0:0:0, 0:0:0);
    (AD_DATA[14] => U[30]) = (0:0:0, 0:0:0);
    (AD_DATA[14] => U[31]) = (0:0:0, 0:0:0);
    (AD_DATA[14] => U[32]) = (0:0:0, 0:0:0);
    (AD_DATA[14] => U[33]) = (0:0:0, 0:0:0);
    (AD_DATA[14] => U[34]) = (0:0:0, 0:0:0);
    (AD_DATA[14] => U[35]) = (0:0:0, 0:0:0);
    (AD_DATA[14] => U[36]) = (0:0:0, 0:0:0);
    (AD_DATA[14] => U[37]) = (0:0:0, 0:0:0);
    (AD_DATA[14] => U[38]) = (0:0:0, 0:0:0);
    (AD_DATA[14] => U[39]) = (0:0:0, 0:0:0);
    (AD_DATA[14] => U[40]) = (0:0:0, 0:0:0);
    (AD_DATA[14] => U[41]) = (0:0:0, 0:0:0);
    (AD_DATA[14] => U[42]) = (0:0:0, 0:0:0);
    (AD_DATA[14] => V[14]) = (0:0:0, 0:0:0);
    (AD_DATA[14] => V[15]) = (0:0:0, 0:0:0);
    (AD_DATA[14] => V[16]) = (0:0:0, 0:0:0);
    (AD_DATA[14] => V[17]) = (0:0:0, 0:0:0);
    (AD_DATA[14] => V[18]) = (0:0:0, 0:0:0);
    (AD_DATA[14] => V[19]) = (0:0:0, 0:0:0);
    (AD_DATA[14] => V[20]) = (0:0:0, 0:0:0);
    (AD_DATA[14] => V[21]) = (0:0:0, 0:0:0);
    (AD_DATA[14] => V[22]) = (0:0:0, 0:0:0);
    (AD_DATA[14] => V[23]) = (0:0:0, 0:0:0);
    (AD_DATA[14] => V[24]) = (0:0:0, 0:0:0);
    (AD_DATA[14] => V[25]) = (0:0:0, 0:0:0);
    (AD_DATA[14] => V[26]) = (0:0:0, 0:0:0);
    (AD_DATA[14] => V[27]) = (0:0:0, 0:0:0);
    (AD_DATA[14] => V[28]) = (0:0:0, 0:0:0);
    (AD_DATA[14] => V[29]) = (0:0:0, 0:0:0);
    (AD_DATA[14] => V[30]) = (0:0:0, 0:0:0);
    (AD_DATA[14] => V[31]) = (0:0:0, 0:0:0);
    (AD_DATA[14] => V[32]) = (0:0:0, 0:0:0);
    (AD_DATA[14] => V[33]) = (0:0:0, 0:0:0);
    (AD_DATA[14] => V[34]) = (0:0:0, 0:0:0);
    (AD_DATA[14] => V[35]) = (0:0:0, 0:0:0);
    (AD_DATA[14] => V[36]) = (0:0:0, 0:0:0);
    (AD_DATA[14] => V[37]) = (0:0:0, 0:0:0);
    (AD_DATA[14] => V[38]) = (0:0:0, 0:0:0);
    (AD_DATA[14] => V[39]) = (0:0:0, 0:0:0);
    (AD_DATA[14] => V[40]) = (0:0:0, 0:0:0);
    (AD_DATA[14] => V[41]) = (0:0:0, 0:0:0);
    (AD_DATA[15] => U[15]) = (0:0:0, 0:0:0);
    (AD_DATA[15] => U[16]) = (0:0:0, 0:0:0);
    (AD_DATA[15] => U[17]) = (0:0:0, 0:0:0);
    (AD_DATA[15] => U[18]) = (0:0:0, 0:0:0);
    (AD_DATA[15] => U[19]) = (0:0:0, 0:0:0);
    (AD_DATA[15] => U[20]) = (0:0:0, 0:0:0);
    (AD_DATA[15] => U[21]) = (0:0:0, 0:0:0);
    (AD_DATA[15] => U[22]) = (0:0:0, 0:0:0);
    (AD_DATA[15] => U[23]) = (0:0:0, 0:0:0);
    (AD_DATA[15] => U[24]) = (0:0:0, 0:0:0);
    (AD_DATA[15] => U[25]) = (0:0:0, 0:0:0);
    (AD_DATA[15] => U[26]) = (0:0:0, 0:0:0);
    (AD_DATA[15] => U[27]) = (0:0:0, 0:0:0);
    (AD_DATA[15] => U[28]) = (0:0:0, 0:0:0);
    (AD_DATA[15] => U[29]) = (0:0:0, 0:0:0);
    (AD_DATA[15] => U[30]) = (0:0:0, 0:0:0);
    (AD_DATA[15] => U[31]) = (0:0:0, 0:0:0);
    (AD_DATA[15] => U[32]) = (0:0:0, 0:0:0);
    (AD_DATA[15] => U[33]) = (0:0:0, 0:0:0);
    (AD_DATA[15] => U[34]) = (0:0:0, 0:0:0);
    (AD_DATA[15] => U[35]) = (0:0:0, 0:0:0);
    (AD_DATA[15] => U[36]) = (0:0:0, 0:0:0);
    (AD_DATA[15] => U[37]) = (0:0:0, 0:0:0);
    (AD_DATA[15] => U[38]) = (0:0:0, 0:0:0);
    (AD_DATA[15] => U[39]) = (0:0:0, 0:0:0);
    (AD_DATA[15] => U[40]) = (0:0:0, 0:0:0);
    (AD_DATA[15] => U[41]) = (0:0:0, 0:0:0);
    (AD_DATA[15] => U[42]) = (0:0:0, 0:0:0);
    (AD_DATA[15] => U[43]) = (0:0:0, 0:0:0);
    (AD_DATA[15] => V[14]) = (0:0:0, 0:0:0);
    (AD_DATA[15] => V[15]) = (0:0:0, 0:0:0);
    (AD_DATA[15] => V[16]) = (0:0:0, 0:0:0);
    (AD_DATA[15] => V[17]) = (0:0:0, 0:0:0);
    (AD_DATA[15] => V[18]) = (0:0:0, 0:0:0);
    (AD_DATA[15] => V[19]) = (0:0:0, 0:0:0);
    (AD_DATA[15] => V[20]) = (0:0:0, 0:0:0);
    (AD_DATA[15] => V[21]) = (0:0:0, 0:0:0);
    (AD_DATA[15] => V[22]) = (0:0:0, 0:0:0);
    (AD_DATA[15] => V[23]) = (0:0:0, 0:0:0);
    (AD_DATA[15] => V[24]) = (0:0:0, 0:0:0);
    (AD_DATA[15] => V[25]) = (0:0:0, 0:0:0);
    (AD_DATA[15] => V[26]) = (0:0:0, 0:0:0);
    (AD_DATA[15] => V[27]) = (0:0:0, 0:0:0);
    (AD_DATA[15] => V[28]) = (0:0:0, 0:0:0);
    (AD_DATA[15] => V[29]) = (0:0:0, 0:0:0);
    (AD_DATA[15] => V[30]) = (0:0:0, 0:0:0);
    (AD_DATA[15] => V[31]) = (0:0:0, 0:0:0);
    (AD_DATA[15] => V[32]) = (0:0:0, 0:0:0);
    (AD_DATA[15] => V[33]) = (0:0:0, 0:0:0);
    (AD_DATA[15] => V[34]) = (0:0:0, 0:0:0);
    (AD_DATA[15] => V[35]) = (0:0:0, 0:0:0);
    (AD_DATA[15] => V[36]) = (0:0:0, 0:0:0);
    (AD_DATA[15] => V[37]) = (0:0:0, 0:0:0);
    (AD_DATA[15] => V[38]) = (0:0:0, 0:0:0);
    (AD_DATA[15] => V[39]) = (0:0:0, 0:0:0);
    (AD_DATA[15] => V[40]) = (0:0:0, 0:0:0);
    (AD_DATA[15] => V[41]) = (0:0:0, 0:0:0);
    (AD_DATA[15] => V[42]) = (0:0:0, 0:0:0);
    (AD_DATA[15] => V[43]) = (0:0:0, 0:0:0);
    (AD_DATA[16] => U[17]) = (0:0:0, 0:0:0);
    (AD_DATA[16] => U[18]) = (0:0:0, 0:0:0);
    (AD_DATA[16] => U[19]) = (0:0:0, 0:0:0);
    (AD_DATA[16] => U[20]) = (0:0:0, 0:0:0);
    (AD_DATA[16] => U[21]) = (0:0:0, 0:0:0);
    (AD_DATA[16] => U[22]) = (0:0:0, 0:0:0);
    (AD_DATA[16] => U[23]) = (0:0:0, 0:0:0);
    (AD_DATA[16] => U[24]) = (0:0:0, 0:0:0);
    (AD_DATA[16] => U[25]) = (0:0:0, 0:0:0);
    (AD_DATA[16] => U[26]) = (0:0:0, 0:0:0);
    (AD_DATA[16] => U[27]) = (0:0:0, 0:0:0);
    (AD_DATA[16] => U[28]) = (0:0:0, 0:0:0);
    (AD_DATA[16] => U[29]) = (0:0:0, 0:0:0);
    (AD_DATA[16] => U[30]) = (0:0:0, 0:0:0);
    (AD_DATA[16] => U[31]) = (0:0:0, 0:0:0);
    (AD_DATA[16] => U[32]) = (0:0:0, 0:0:0);
    (AD_DATA[16] => U[33]) = (0:0:0, 0:0:0);
    (AD_DATA[16] => U[34]) = (0:0:0, 0:0:0);
    (AD_DATA[16] => U[35]) = (0:0:0, 0:0:0);
    (AD_DATA[16] => U[36]) = (0:0:0, 0:0:0);
    (AD_DATA[16] => U[37]) = (0:0:0, 0:0:0);
    (AD_DATA[16] => U[38]) = (0:0:0, 0:0:0);
    (AD_DATA[16] => U[39]) = (0:0:0, 0:0:0);
    (AD_DATA[16] => U[40]) = (0:0:0, 0:0:0);
    (AD_DATA[16] => U[41]) = (0:0:0, 0:0:0);
    (AD_DATA[16] => U[42]) = (0:0:0, 0:0:0);
    (AD_DATA[16] => U[43]) = (0:0:0, 0:0:0);
    (AD_DATA[16] => V[16]) = (0:0:0, 0:0:0);
    (AD_DATA[16] => V[17]) = (0:0:0, 0:0:0);
    (AD_DATA[16] => V[18]) = (0:0:0, 0:0:0);
    (AD_DATA[16] => V[19]) = (0:0:0, 0:0:0);
    (AD_DATA[16] => V[20]) = (0:0:0, 0:0:0);
    (AD_DATA[16] => V[21]) = (0:0:0, 0:0:0);
    (AD_DATA[16] => V[22]) = (0:0:0, 0:0:0);
    (AD_DATA[16] => V[23]) = (0:0:0, 0:0:0);
    (AD_DATA[16] => V[24]) = (0:0:0, 0:0:0);
    (AD_DATA[16] => V[25]) = (0:0:0, 0:0:0);
    (AD_DATA[16] => V[26]) = (0:0:0, 0:0:0);
    (AD_DATA[16] => V[27]) = (0:0:0, 0:0:0);
    (AD_DATA[16] => V[28]) = (0:0:0, 0:0:0);
    (AD_DATA[16] => V[29]) = (0:0:0, 0:0:0);
    (AD_DATA[16] => V[30]) = (0:0:0, 0:0:0);
    (AD_DATA[16] => V[31]) = (0:0:0, 0:0:0);
    (AD_DATA[16] => V[32]) = (0:0:0, 0:0:0);
    (AD_DATA[16] => V[33]) = (0:0:0, 0:0:0);
    (AD_DATA[16] => V[34]) = (0:0:0, 0:0:0);
    (AD_DATA[16] => V[35]) = (0:0:0, 0:0:0);
    (AD_DATA[16] => V[36]) = (0:0:0, 0:0:0);
    (AD_DATA[16] => V[37]) = (0:0:0, 0:0:0);
    (AD_DATA[16] => V[38]) = (0:0:0, 0:0:0);
    (AD_DATA[16] => V[39]) = (0:0:0, 0:0:0);
    (AD_DATA[16] => V[40]) = (0:0:0, 0:0:0);
    (AD_DATA[16] => V[41]) = (0:0:0, 0:0:0);
    (AD_DATA[16] => V[42]) = (0:0:0, 0:0:0);
    (AD_DATA[16] => V[43]) = (0:0:0, 0:0:0);
    (AD_DATA[17] => BMULT17) = (0:0:0, 0:0:0);
    (AD_DATA[17] => U[17]) = (0:0:0, 0:0:0);
    (AD_DATA[17] => U[18]) = (0:0:0, 0:0:0);
    (AD_DATA[17] => U[19]) = (0:0:0, 0:0:0);
    (AD_DATA[17] => U[20]) = (0:0:0, 0:0:0);
    (AD_DATA[17] => U[21]) = (0:0:0, 0:0:0);
    (AD_DATA[17] => U[22]) = (0:0:0, 0:0:0);
    (AD_DATA[17] => U[23]) = (0:0:0, 0:0:0);
    (AD_DATA[17] => U[24]) = (0:0:0, 0:0:0);
    (AD_DATA[17] => U[25]) = (0:0:0, 0:0:0);
    (AD_DATA[17] => U[26]) = (0:0:0, 0:0:0);
    (AD_DATA[17] => U[27]) = (0:0:0, 0:0:0);
    (AD_DATA[17] => U[28]) = (0:0:0, 0:0:0);
    (AD_DATA[17] => U[29]) = (0:0:0, 0:0:0);
    (AD_DATA[17] => U[30]) = (0:0:0, 0:0:0);
    (AD_DATA[17] => U[31]) = (0:0:0, 0:0:0);
    (AD_DATA[17] => U[32]) = (0:0:0, 0:0:0);
    (AD_DATA[17] => U[33]) = (0:0:0, 0:0:0);
    (AD_DATA[17] => U[34]) = (0:0:0, 0:0:0);
    (AD_DATA[17] => U[35]) = (0:0:0, 0:0:0);
    (AD_DATA[17] => U[36]) = (0:0:0, 0:0:0);
    (AD_DATA[17] => U[37]) = (0:0:0, 0:0:0);
    (AD_DATA[17] => U[38]) = (0:0:0, 0:0:0);
    (AD_DATA[17] => U[39]) = (0:0:0, 0:0:0);
    (AD_DATA[17] => U[40]) = (0:0:0, 0:0:0);
    (AD_DATA[17] => U[41]) = (0:0:0, 0:0:0);
    (AD_DATA[17] => U[42]) = (0:0:0, 0:0:0);
    (AD_DATA[17] => U[43]) = (0:0:0, 0:0:0);
    (AD_DATA[17] => V[16]) = (0:0:0, 0:0:0);
    (AD_DATA[17] => V[17]) = (0:0:0, 0:0:0);
    (AD_DATA[17] => V[18]) = (0:0:0, 0:0:0);
    (AD_DATA[17] => V[19]) = (0:0:0, 0:0:0);
    (AD_DATA[17] => V[20]) = (0:0:0, 0:0:0);
    (AD_DATA[17] => V[21]) = (0:0:0, 0:0:0);
    (AD_DATA[17] => V[22]) = (0:0:0, 0:0:0);
    (AD_DATA[17] => V[23]) = (0:0:0, 0:0:0);
    (AD_DATA[17] => V[24]) = (0:0:0, 0:0:0);
    (AD_DATA[17] => V[25]) = (0:0:0, 0:0:0);
    (AD_DATA[17] => V[26]) = (0:0:0, 0:0:0);
    (AD_DATA[17] => V[27]) = (0:0:0, 0:0:0);
    (AD_DATA[17] => V[28]) = (0:0:0, 0:0:0);
    (AD_DATA[17] => V[29]) = (0:0:0, 0:0:0);
    (AD_DATA[17] => V[30]) = (0:0:0, 0:0:0);
    (AD_DATA[17] => V[31]) = (0:0:0, 0:0:0);
    (AD_DATA[17] => V[32]) = (0:0:0, 0:0:0);
    (AD_DATA[17] => V[33]) = (0:0:0, 0:0:0);
    (AD_DATA[17] => V[34]) = (0:0:0, 0:0:0);
    (AD_DATA[17] => V[35]) = (0:0:0, 0:0:0);
    (AD_DATA[17] => V[36]) = (0:0:0, 0:0:0);
    (AD_DATA[17] => V[37]) = (0:0:0, 0:0:0);
    (AD_DATA[17] => V[38]) = (0:0:0, 0:0:0);
    (AD_DATA[17] => V[39]) = (0:0:0, 0:0:0);
    (AD_DATA[17] => V[40]) = (0:0:0, 0:0:0);
    (AD_DATA[17] => V[41]) = (0:0:0, 0:0:0);
    (AD_DATA[17] => V[42]) = (0:0:0, 0:0:0);
    (AD_DATA[17] => V[43]) = (0:0:0, 0:0:0);
    (AD_DATA[18] => U[19]) = (0:0:0, 0:0:0);
    (AD_DATA[18] => U[20]) = (0:0:0, 0:0:0);
    (AD_DATA[18] => U[21]) = (0:0:0, 0:0:0);
    (AD_DATA[18] => U[22]) = (0:0:0, 0:0:0);
    (AD_DATA[18] => U[23]) = (0:0:0, 0:0:0);
    (AD_DATA[18] => U[24]) = (0:0:0, 0:0:0);
    (AD_DATA[18] => U[25]) = (0:0:0, 0:0:0);
    (AD_DATA[18] => U[26]) = (0:0:0, 0:0:0);
    (AD_DATA[18] => U[27]) = (0:0:0, 0:0:0);
    (AD_DATA[18] => U[28]) = (0:0:0, 0:0:0);
    (AD_DATA[18] => U[29]) = (0:0:0, 0:0:0);
    (AD_DATA[18] => U[30]) = (0:0:0, 0:0:0);
    (AD_DATA[18] => U[31]) = (0:0:0, 0:0:0);
    (AD_DATA[18] => U[32]) = (0:0:0, 0:0:0);
    (AD_DATA[18] => U[33]) = (0:0:0, 0:0:0);
    (AD_DATA[18] => U[34]) = (0:0:0, 0:0:0);
    (AD_DATA[18] => U[35]) = (0:0:0, 0:0:0);
    (AD_DATA[18] => U[36]) = (0:0:0, 0:0:0);
    (AD_DATA[18] => U[37]) = (0:0:0, 0:0:0);
    (AD_DATA[18] => U[38]) = (0:0:0, 0:0:0);
    (AD_DATA[18] => V[18]) = (0:0:0, 0:0:0);
    (AD_DATA[18] => V[19]) = (0:0:0, 0:0:0);
    (AD_DATA[18] => V[20]) = (0:0:0, 0:0:0);
    (AD_DATA[18] => V[21]) = (0:0:0, 0:0:0);
    (AD_DATA[18] => V[22]) = (0:0:0, 0:0:0);
    (AD_DATA[18] => V[23]) = (0:0:0, 0:0:0);
    (AD_DATA[18] => V[24]) = (0:0:0, 0:0:0);
    (AD_DATA[18] => V[25]) = (0:0:0, 0:0:0);
    (AD_DATA[18] => V[26]) = (0:0:0, 0:0:0);
    (AD_DATA[18] => V[27]) = (0:0:0, 0:0:0);
    (AD_DATA[18] => V[28]) = (0:0:0, 0:0:0);
    (AD_DATA[18] => V[29]) = (0:0:0, 0:0:0);
    (AD_DATA[18] => V[30]) = (0:0:0, 0:0:0);
    (AD_DATA[18] => V[31]) = (0:0:0, 0:0:0);
    (AD_DATA[18] => V[32]) = (0:0:0, 0:0:0);
    (AD_DATA[18] => V[33]) = (0:0:0, 0:0:0);
    (AD_DATA[18] => V[34]) = (0:0:0, 0:0:0);
    (AD_DATA[18] => V[35]) = (0:0:0, 0:0:0);
    (AD_DATA[18] => V[36]) = (0:0:0, 0:0:0);
    (AD_DATA[18] => V[37]) = (0:0:0, 0:0:0);
    (AD_DATA[19] => U[20]) = (0:0:0, 0:0:0);
    (AD_DATA[19] => U[21]) = (0:0:0, 0:0:0);
    (AD_DATA[19] => U[22]) = (0:0:0, 0:0:0);
    (AD_DATA[19] => U[23]) = (0:0:0, 0:0:0);
    (AD_DATA[19] => U[24]) = (0:0:0, 0:0:0);
    (AD_DATA[19] => U[25]) = (0:0:0, 0:0:0);
    (AD_DATA[19] => U[26]) = (0:0:0, 0:0:0);
    (AD_DATA[19] => U[27]) = (0:0:0, 0:0:0);
    (AD_DATA[19] => U[28]) = (0:0:0, 0:0:0);
    (AD_DATA[19] => U[29]) = (0:0:0, 0:0:0);
    (AD_DATA[19] => U[30]) = (0:0:0, 0:0:0);
    (AD_DATA[19] => U[31]) = (0:0:0, 0:0:0);
    (AD_DATA[19] => U[32]) = (0:0:0, 0:0:0);
    (AD_DATA[19] => U[33]) = (0:0:0, 0:0:0);
    (AD_DATA[19] => U[34]) = (0:0:0, 0:0:0);
    (AD_DATA[19] => U[35]) = (0:0:0, 0:0:0);
    (AD_DATA[19] => U[36]) = (0:0:0, 0:0:0);
    (AD_DATA[19] => U[37]) = (0:0:0, 0:0:0);
    (AD_DATA[19] => U[38]) = (0:0:0, 0:0:0);
    (AD_DATA[19] => U[39]) = (0:0:0, 0:0:0);
    (AD_DATA[19] => V[19]) = (0:0:0, 0:0:0);
    (AD_DATA[19] => V[20]) = (0:0:0, 0:0:0);
    (AD_DATA[19] => V[21]) = (0:0:0, 0:0:0);
    (AD_DATA[19] => V[22]) = (0:0:0, 0:0:0);
    (AD_DATA[19] => V[23]) = (0:0:0, 0:0:0);
    (AD_DATA[19] => V[24]) = (0:0:0, 0:0:0);
    (AD_DATA[19] => V[25]) = (0:0:0, 0:0:0);
    (AD_DATA[19] => V[26]) = (0:0:0, 0:0:0);
    (AD_DATA[19] => V[27]) = (0:0:0, 0:0:0);
    (AD_DATA[19] => V[28]) = (0:0:0, 0:0:0);
    (AD_DATA[19] => V[29]) = (0:0:0, 0:0:0);
    (AD_DATA[19] => V[30]) = (0:0:0, 0:0:0);
    (AD_DATA[19] => V[31]) = (0:0:0, 0:0:0);
    (AD_DATA[19] => V[32]) = (0:0:0, 0:0:0);
    (AD_DATA[19] => V[33]) = (0:0:0, 0:0:0);
    (AD_DATA[19] => V[34]) = (0:0:0, 0:0:0);
    (AD_DATA[19] => V[35]) = (0:0:0, 0:0:0);
    (AD_DATA[19] => V[36]) = (0:0:0, 0:0:0);
    (AD_DATA[19] => V[37]) = (0:0:0, 0:0:0);
    (AD_DATA[19] => V[38]) = (0:0:0, 0:0:0);
    (AD_DATA[1] => U[0]) = (0:0:0, 0:0:0);
    (AD_DATA[1] => U[10]) = (0:0:0, 0:0:0);
    (AD_DATA[1] => U[11]) = (0:0:0, 0:0:0);
    (AD_DATA[1] => U[12]) = (0:0:0, 0:0:0);
    (AD_DATA[1] => U[13]) = (0:0:0, 0:0:0);
    (AD_DATA[1] => U[14]) = (0:0:0, 0:0:0);
    (AD_DATA[1] => U[15]) = (0:0:0, 0:0:0);
    (AD_DATA[1] => U[16]) = (0:0:0, 0:0:0);
    (AD_DATA[1] => U[17]) = (0:0:0, 0:0:0);
    (AD_DATA[1] => U[18]) = (0:0:0, 0:0:0);
    (AD_DATA[1] => U[19]) = (0:0:0, 0:0:0);
    (AD_DATA[1] => U[1]) = (0:0:0, 0:0:0);
    (AD_DATA[1] => U[20]) = (0:0:0, 0:0:0);
    (AD_DATA[1] => U[21]) = (0:0:0, 0:0:0);
    (AD_DATA[1] => U[22]) = (0:0:0, 0:0:0);
    (AD_DATA[1] => U[23]) = (0:0:0, 0:0:0);
    (AD_DATA[1] => U[24]) = (0:0:0, 0:0:0);
    (AD_DATA[1] => U[25]) = (0:0:0, 0:0:0);
    (AD_DATA[1] => U[26]) = (0:0:0, 0:0:0);
    (AD_DATA[1] => U[27]) = (0:0:0, 0:0:0);
    (AD_DATA[1] => U[28]) = (0:0:0, 0:0:0);
    (AD_DATA[1] => U[29]) = (0:0:0, 0:0:0);
    (AD_DATA[1] => U[2]) = (0:0:0, 0:0:0);
    (AD_DATA[1] => U[30]) = (0:0:0, 0:0:0);
    (AD_DATA[1] => U[31]) = (0:0:0, 0:0:0);
    (AD_DATA[1] => U[32]) = (0:0:0, 0:0:0);
    (AD_DATA[1] => U[33]) = (0:0:0, 0:0:0);
    (AD_DATA[1] => U[3]) = (0:0:0, 0:0:0);
    (AD_DATA[1] => U[4]) = (0:0:0, 0:0:0);
    (AD_DATA[1] => U[5]) = (0:0:0, 0:0:0);
    (AD_DATA[1] => U[6]) = (0:0:0, 0:0:0);
    (AD_DATA[1] => U[7]) = (0:0:0, 0:0:0);
    (AD_DATA[1] => U[8]) = (0:0:0, 0:0:0);
    (AD_DATA[1] => U[9]) = (0:0:0, 0:0:0);
    (AD_DATA[1] => V[0]) = (0:0:0, 0:0:0);
    (AD_DATA[1] => V[10]) = (0:0:0, 0:0:0);
    (AD_DATA[1] => V[11]) = (0:0:0, 0:0:0);
    (AD_DATA[1] => V[12]) = (0:0:0, 0:0:0);
    (AD_DATA[1] => V[13]) = (0:0:0, 0:0:0);
    (AD_DATA[1] => V[14]) = (0:0:0, 0:0:0);
    (AD_DATA[1] => V[15]) = (0:0:0, 0:0:0);
    (AD_DATA[1] => V[16]) = (0:0:0, 0:0:0);
    (AD_DATA[1] => V[17]) = (0:0:0, 0:0:0);
    (AD_DATA[1] => V[18]) = (0:0:0, 0:0:0);
    (AD_DATA[1] => V[19]) = (0:0:0, 0:0:0);
    (AD_DATA[1] => V[20]) = (0:0:0, 0:0:0);
    (AD_DATA[1] => V[21]) = (0:0:0, 0:0:0);
    (AD_DATA[1] => V[22]) = (0:0:0, 0:0:0);
    (AD_DATA[1] => V[23]) = (0:0:0, 0:0:0);
    (AD_DATA[1] => V[24]) = (0:0:0, 0:0:0);
    (AD_DATA[1] => V[25]) = (0:0:0, 0:0:0);
    (AD_DATA[1] => V[26]) = (0:0:0, 0:0:0);
    (AD_DATA[1] => V[27]) = (0:0:0, 0:0:0);
    (AD_DATA[1] => V[28]) = (0:0:0, 0:0:0);
    (AD_DATA[1] => V[29]) = (0:0:0, 0:0:0);
    (AD_DATA[1] => V[30]) = (0:0:0, 0:0:0);
    (AD_DATA[1] => V[31]) = (0:0:0, 0:0:0);
    (AD_DATA[1] => V[32]) = (0:0:0, 0:0:0);
    (AD_DATA[1] => V[4]) = (0:0:0, 0:0:0);
    (AD_DATA[1] => V[5]) = (0:0:0, 0:0:0);
    (AD_DATA[1] => V[6]) = (0:0:0, 0:0:0);
    (AD_DATA[1] => V[7]) = (0:0:0, 0:0:0);
    (AD_DATA[1] => V[8]) = (0:0:0, 0:0:0);
    (AD_DATA[1] => V[9]) = (0:0:0, 0:0:0);
    (AD_DATA[20] => U[21]) = (0:0:0, 0:0:0);
    (AD_DATA[20] => U[22]) = (0:0:0, 0:0:0);
    (AD_DATA[20] => U[23]) = (0:0:0, 0:0:0);
    (AD_DATA[20] => U[24]) = (0:0:0, 0:0:0);
    (AD_DATA[20] => U[25]) = (0:0:0, 0:0:0);
    (AD_DATA[20] => U[26]) = (0:0:0, 0:0:0);
    (AD_DATA[20] => U[27]) = (0:0:0, 0:0:0);
    (AD_DATA[20] => U[28]) = (0:0:0, 0:0:0);
    (AD_DATA[20] => U[29]) = (0:0:0, 0:0:0);
    (AD_DATA[20] => U[30]) = (0:0:0, 0:0:0);
    (AD_DATA[20] => U[31]) = (0:0:0, 0:0:0);
    (AD_DATA[20] => U[32]) = (0:0:0, 0:0:0);
    (AD_DATA[20] => U[33]) = (0:0:0, 0:0:0);
    (AD_DATA[20] => U[34]) = (0:0:0, 0:0:0);
    (AD_DATA[20] => U[35]) = (0:0:0, 0:0:0);
    (AD_DATA[20] => U[36]) = (0:0:0, 0:0:0);
    (AD_DATA[20] => U[37]) = (0:0:0, 0:0:0);
    (AD_DATA[20] => U[38]) = (0:0:0, 0:0:0);
    (AD_DATA[20] => U[39]) = (0:0:0, 0:0:0);
    (AD_DATA[20] => V[20]) = (0:0:0, 0:0:0);
    (AD_DATA[20] => V[21]) = (0:0:0, 0:0:0);
    (AD_DATA[20] => V[22]) = (0:0:0, 0:0:0);
    (AD_DATA[20] => V[23]) = (0:0:0, 0:0:0);
    (AD_DATA[20] => V[24]) = (0:0:0, 0:0:0);
    (AD_DATA[20] => V[25]) = (0:0:0, 0:0:0);
    (AD_DATA[20] => V[26]) = (0:0:0, 0:0:0);
    (AD_DATA[20] => V[27]) = (0:0:0, 0:0:0);
    (AD_DATA[20] => V[28]) = (0:0:0, 0:0:0);
    (AD_DATA[20] => V[29]) = (0:0:0, 0:0:0);
    (AD_DATA[20] => V[30]) = (0:0:0, 0:0:0);
    (AD_DATA[20] => V[31]) = (0:0:0, 0:0:0);
    (AD_DATA[20] => V[32]) = (0:0:0, 0:0:0);
    (AD_DATA[20] => V[33]) = (0:0:0, 0:0:0);
    (AD_DATA[20] => V[34]) = (0:0:0, 0:0:0);
    (AD_DATA[20] => V[35]) = (0:0:0, 0:0:0);
    (AD_DATA[20] => V[36]) = (0:0:0, 0:0:0);
    (AD_DATA[20] => V[37]) = (0:0:0, 0:0:0);
    (AD_DATA[20] => V[38]) = (0:0:0, 0:0:0);
    (AD_DATA[21] => U[22]) = (0:0:0, 0:0:0);
    (AD_DATA[21] => U[23]) = (0:0:0, 0:0:0);
    (AD_DATA[21] => U[24]) = (0:0:0, 0:0:0);
    (AD_DATA[21] => U[25]) = (0:0:0, 0:0:0);
    (AD_DATA[21] => U[26]) = (0:0:0, 0:0:0);
    (AD_DATA[21] => U[27]) = (0:0:0, 0:0:0);
    (AD_DATA[21] => U[28]) = (0:0:0, 0:0:0);
    (AD_DATA[21] => U[29]) = (0:0:0, 0:0:0);
    (AD_DATA[21] => U[30]) = (0:0:0, 0:0:0);
    (AD_DATA[21] => U[31]) = (0:0:0, 0:0:0);
    (AD_DATA[21] => U[32]) = (0:0:0, 0:0:0);
    (AD_DATA[21] => U[33]) = (0:0:0, 0:0:0);
    (AD_DATA[21] => U[34]) = (0:0:0, 0:0:0);
    (AD_DATA[21] => U[35]) = (0:0:0, 0:0:0);
    (AD_DATA[21] => U[36]) = (0:0:0, 0:0:0);
    (AD_DATA[21] => U[37]) = (0:0:0, 0:0:0);
    (AD_DATA[21] => U[38]) = (0:0:0, 0:0:0);
    (AD_DATA[21] => U[39]) = (0:0:0, 0:0:0);
    (AD_DATA[21] => U[40]) = (0:0:0, 0:0:0);
    (AD_DATA[21] => V[21]) = (0:0:0, 0:0:0);
    (AD_DATA[21] => V[22]) = (0:0:0, 0:0:0);
    (AD_DATA[21] => V[23]) = (0:0:0, 0:0:0);
    (AD_DATA[21] => V[24]) = (0:0:0, 0:0:0);
    (AD_DATA[21] => V[25]) = (0:0:0, 0:0:0);
    (AD_DATA[21] => V[26]) = (0:0:0, 0:0:0);
    (AD_DATA[21] => V[27]) = (0:0:0, 0:0:0);
    (AD_DATA[21] => V[28]) = (0:0:0, 0:0:0);
    (AD_DATA[21] => V[29]) = (0:0:0, 0:0:0);
    (AD_DATA[21] => V[30]) = (0:0:0, 0:0:0);
    (AD_DATA[21] => V[31]) = (0:0:0, 0:0:0);
    (AD_DATA[21] => V[32]) = (0:0:0, 0:0:0);
    (AD_DATA[21] => V[33]) = (0:0:0, 0:0:0);
    (AD_DATA[21] => V[34]) = (0:0:0, 0:0:0);
    (AD_DATA[21] => V[35]) = (0:0:0, 0:0:0);
    (AD_DATA[21] => V[36]) = (0:0:0, 0:0:0);
    (AD_DATA[21] => V[37]) = (0:0:0, 0:0:0);
    (AD_DATA[21] => V[38]) = (0:0:0, 0:0:0);
    (AD_DATA[21] => V[39]) = (0:0:0, 0:0:0);
    (AD_DATA[22] => U[23]) = (0:0:0, 0:0:0);
    (AD_DATA[22] => U[24]) = (0:0:0, 0:0:0);
    (AD_DATA[22] => U[25]) = (0:0:0, 0:0:0);
    (AD_DATA[22] => U[26]) = (0:0:0, 0:0:0);
    (AD_DATA[22] => U[27]) = (0:0:0, 0:0:0);
    (AD_DATA[22] => U[28]) = (0:0:0, 0:0:0);
    (AD_DATA[22] => U[29]) = (0:0:0, 0:0:0);
    (AD_DATA[22] => U[30]) = (0:0:0, 0:0:0);
    (AD_DATA[22] => U[31]) = (0:0:0, 0:0:0);
    (AD_DATA[22] => U[32]) = (0:0:0, 0:0:0);
    (AD_DATA[22] => U[33]) = (0:0:0, 0:0:0);
    (AD_DATA[22] => U[34]) = (0:0:0, 0:0:0);
    (AD_DATA[22] => U[35]) = (0:0:0, 0:0:0);
    (AD_DATA[22] => U[36]) = (0:0:0, 0:0:0);
    (AD_DATA[22] => U[37]) = (0:0:0, 0:0:0);
    (AD_DATA[22] => U[38]) = (0:0:0, 0:0:0);
    (AD_DATA[22] => U[39]) = (0:0:0, 0:0:0);
    (AD_DATA[22] => U[40]) = (0:0:0, 0:0:0);
    (AD_DATA[22] => U[41]) = (0:0:0, 0:0:0);
    (AD_DATA[22] => V[22]) = (0:0:0, 0:0:0);
    (AD_DATA[22] => V[23]) = (0:0:0, 0:0:0);
    (AD_DATA[22] => V[24]) = (0:0:0, 0:0:0);
    (AD_DATA[22] => V[25]) = (0:0:0, 0:0:0);
    (AD_DATA[22] => V[26]) = (0:0:0, 0:0:0);
    (AD_DATA[22] => V[27]) = (0:0:0, 0:0:0);
    (AD_DATA[22] => V[28]) = (0:0:0, 0:0:0);
    (AD_DATA[22] => V[29]) = (0:0:0, 0:0:0);
    (AD_DATA[22] => V[30]) = (0:0:0, 0:0:0);
    (AD_DATA[22] => V[31]) = (0:0:0, 0:0:0);
    (AD_DATA[22] => V[32]) = (0:0:0, 0:0:0);
    (AD_DATA[22] => V[33]) = (0:0:0, 0:0:0);
    (AD_DATA[22] => V[34]) = (0:0:0, 0:0:0);
    (AD_DATA[22] => V[35]) = (0:0:0, 0:0:0);
    (AD_DATA[22] => V[36]) = (0:0:0, 0:0:0);
    (AD_DATA[22] => V[37]) = (0:0:0, 0:0:0);
    (AD_DATA[22] => V[38]) = (0:0:0, 0:0:0);
    (AD_DATA[22] => V[39]) = (0:0:0, 0:0:0);
    (AD_DATA[22] => V[40]) = (0:0:0, 0:0:0);
    (AD_DATA[23] => U[24]) = (0:0:0, 0:0:0);
    (AD_DATA[23] => U[25]) = (0:0:0, 0:0:0);
    (AD_DATA[23] => U[26]) = (0:0:0, 0:0:0);
    (AD_DATA[23] => U[27]) = (0:0:0, 0:0:0);
    (AD_DATA[23] => U[28]) = (0:0:0, 0:0:0);
    (AD_DATA[23] => U[29]) = (0:0:0, 0:0:0);
    (AD_DATA[23] => U[30]) = (0:0:0, 0:0:0);
    (AD_DATA[23] => U[31]) = (0:0:0, 0:0:0);
    (AD_DATA[23] => U[32]) = (0:0:0, 0:0:0);
    (AD_DATA[23] => U[33]) = (0:0:0, 0:0:0);
    (AD_DATA[23] => U[34]) = (0:0:0, 0:0:0);
    (AD_DATA[23] => U[35]) = (0:0:0, 0:0:0);
    (AD_DATA[23] => U[36]) = (0:0:0, 0:0:0);
    (AD_DATA[23] => U[37]) = (0:0:0, 0:0:0);
    (AD_DATA[23] => U[38]) = (0:0:0, 0:0:0);
    (AD_DATA[23] => U[39]) = (0:0:0, 0:0:0);
    (AD_DATA[23] => U[40]) = (0:0:0, 0:0:0);
    (AD_DATA[23] => U[41]) = (0:0:0, 0:0:0);
    (AD_DATA[23] => U[42]) = (0:0:0, 0:0:0);
    (AD_DATA[23] => V[23]) = (0:0:0, 0:0:0);
    (AD_DATA[23] => V[24]) = (0:0:0, 0:0:0);
    (AD_DATA[23] => V[25]) = (0:0:0, 0:0:0);
    (AD_DATA[23] => V[26]) = (0:0:0, 0:0:0);
    (AD_DATA[23] => V[27]) = (0:0:0, 0:0:0);
    (AD_DATA[23] => V[28]) = (0:0:0, 0:0:0);
    (AD_DATA[23] => V[29]) = (0:0:0, 0:0:0);
    (AD_DATA[23] => V[30]) = (0:0:0, 0:0:0);
    (AD_DATA[23] => V[31]) = (0:0:0, 0:0:0);
    (AD_DATA[23] => V[32]) = (0:0:0, 0:0:0);
    (AD_DATA[23] => V[33]) = (0:0:0, 0:0:0);
    (AD_DATA[23] => V[34]) = (0:0:0, 0:0:0);
    (AD_DATA[23] => V[35]) = (0:0:0, 0:0:0);
    (AD_DATA[23] => V[36]) = (0:0:0, 0:0:0);
    (AD_DATA[23] => V[37]) = (0:0:0, 0:0:0);
    (AD_DATA[23] => V[38]) = (0:0:0, 0:0:0);
    (AD_DATA[23] => V[39]) = (0:0:0, 0:0:0);
    (AD_DATA[23] => V[40]) = (0:0:0, 0:0:0);
    (AD_DATA[23] => V[41]) = (0:0:0, 0:0:0);
    (AD_DATA[24] => U[25]) = (0:0:0, 0:0:0);
    (AD_DATA[24] => U[26]) = (0:0:0, 0:0:0);
    (AD_DATA[24] => U[27]) = (0:0:0, 0:0:0);
    (AD_DATA[24] => U[28]) = (0:0:0, 0:0:0);
    (AD_DATA[24] => U[29]) = (0:0:0, 0:0:0);
    (AD_DATA[24] => U[30]) = (0:0:0, 0:0:0);
    (AD_DATA[24] => U[31]) = (0:0:0, 0:0:0);
    (AD_DATA[24] => U[32]) = (0:0:0, 0:0:0);
    (AD_DATA[24] => U[33]) = (0:0:0, 0:0:0);
    (AD_DATA[24] => U[34]) = (0:0:0, 0:0:0);
    (AD_DATA[24] => U[35]) = (0:0:0, 0:0:0);
    (AD_DATA[24] => U[36]) = (0:0:0, 0:0:0);
    (AD_DATA[24] => U[37]) = (0:0:0, 0:0:0);
    (AD_DATA[24] => U[38]) = (0:0:0, 0:0:0);
    (AD_DATA[24] => U[39]) = (0:0:0, 0:0:0);
    (AD_DATA[24] => U[40]) = (0:0:0, 0:0:0);
    (AD_DATA[24] => U[41]) = (0:0:0, 0:0:0);
    (AD_DATA[24] => U[42]) = (0:0:0, 0:0:0);
    (AD_DATA[24] => V[24]) = (0:0:0, 0:0:0);
    (AD_DATA[24] => V[25]) = (0:0:0, 0:0:0);
    (AD_DATA[24] => V[26]) = (0:0:0, 0:0:0);
    (AD_DATA[24] => V[27]) = (0:0:0, 0:0:0);
    (AD_DATA[24] => V[28]) = (0:0:0, 0:0:0);
    (AD_DATA[24] => V[29]) = (0:0:0, 0:0:0);
    (AD_DATA[24] => V[30]) = (0:0:0, 0:0:0);
    (AD_DATA[24] => V[31]) = (0:0:0, 0:0:0);
    (AD_DATA[24] => V[32]) = (0:0:0, 0:0:0);
    (AD_DATA[24] => V[33]) = (0:0:0, 0:0:0);
    (AD_DATA[24] => V[34]) = (0:0:0, 0:0:0);
    (AD_DATA[24] => V[35]) = (0:0:0, 0:0:0);
    (AD_DATA[24] => V[36]) = (0:0:0, 0:0:0);
    (AD_DATA[24] => V[37]) = (0:0:0, 0:0:0);
    (AD_DATA[24] => V[38]) = (0:0:0, 0:0:0);
    (AD_DATA[24] => V[39]) = (0:0:0, 0:0:0);
    (AD_DATA[24] => V[40]) = (0:0:0, 0:0:0);
    (AD_DATA[24] => V[41]) = (0:0:0, 0:0:0);
    (AD_DATA[25] => U[26]) = (0:0:0, 0:0:0);
    (AD_DATA[25] => U[27]) = (0:0:0, 0:0:0);
    (AD_DATA[25] => U[28]) = (0:0:0, 0:0:0);
    (AD_DATA[25] => U[29]) = (0:0:0, 0:0:0);
    (AD_DATA[25] => U[30]) = (0:0:0, 0:0:0);
    (AD_DATA[25] => U[31]) = (0:0:0, 0:0:0);
    (AD_DATA[25] => U[32]) = (0:0:0, 0:0:0);
    (AD_DATA[25] => U[33]) = (0:0:0, 0:0:0);
    (AD_DATA[25] => U[34]) = (0:0:0, 0:0:0);
    (AD_DATA[25] => U[35]) = (0:0:0, 0:0:0);
    (AD_DATA[25] => U[36]) = (0:0:0, 0:0:0);
    (AD_DATA[25] => U[37]) = (0:0:0, 0:0:0);
    (AD_DATA[25] => U[38]) = (0:0:0, 0:0:0);
    (AD_DATA[25] => U[39]) = (0:0:0, 0:0:0);
    (AD_DATA[25] => U[40]) = (0:0:0, 0:0:0);
    (AD_DATA[25] => U[41]) = (0:0:0, 0:0:0);
    (AD_DATA[25] => U[42]) = (0:0:0, 0:0:0);
    (AD_DATA[25] => U[43]) = (0:0:0, 0:0:0);
    (AD_DATA[25] => V[25]) = (0:0:0, 0:0:0);
    (AD_DATA[25] => V[26]) = (0:0:0, 0:0:0);
    (AD_DATA[25] => V[27]) = (0:0:0, 0:0:0);
    (AD_DATA[25] => V[28]) = (0:0:0, 0:0:0);
    (AD_DATA[25] => V[29]) = (0:0:0, 0:0:0);
    (AD_DATA[25] => V[30]) = (0:0:0, 0:0:0);
    (AD_DATA[25] => V[31]) = (0:0:0, 0:0:0);
    (AD_DATA[25] => V[32]) = (0:0:0, 0:0:0);
    (AD_DATA[25] => V[33]) = (0:0:0, 0:0:0);
    (AD_DATA[25] => V[34]) = (0:0:0, 0:0:0);
    (AD_DATA[25] => V[35]) = (0:0:0, 0:0:0);
    (AD_DATA[25] => V[36]) = (0:0:0, 0:0:0);
    (AD_DATA[25] => V[37]) = (0:0:0, 0:0:0);
    (AD_DATA[25] => V[38]) = (0:0:0, 0:0:0);
    (AD_DATA[25] => V[39]) = (0:0:0, 0:0:0);
    (AD_DATA[25] => V[40]) = (0:0:0, 0:0:0);
    (AD_DATA[25] => V[41]) = (0:0:0, 0:0:0);
    (AD_DATA[25] => V[42]) = (0:0:0, 0:0:0);
    (AD_DATA[26] => AMULT26) = (0:0:0, 0:0:0);
    (AD_DATA[26] => U[27]) = (0:0:0, 0:0:0);
    (AD_DATA[26] => U[28]) = (0:0:0, 0:0:0);
    (AD_DATA[26] => U[29]) = (0:0:0, 0:0:0);
    (AD_DATA[26] => U[30]) = (0:0:0, 0:0:0);
    (AD_DATA[26] => U[31]) = (0:0:0, 0:0:0);
    (AD_DATA[26] => U[32]) = (0:0:0, 0:0:0);
    (AD_DATA[26] => U[33]) = (0:0:0, 0:0:0);
    (AD_DATA[26] => U[34]) = (0:0:0, 0:0:0);
    (AD_DATA[26] => U[35]) = (0:0:0, 0:0:0);
    (AD_DATA[26] => U[36]) = (0:0:0, 0:0:0);
    (AD_DATA[26] => U[37]) = (0:0:0, 0:0:0);
    (AD_DATA[26] => U[38]) = (0:0:0, 0:0:0);
    (AD_DATA[26] => U[39]) = (0:0:0, 0:0:0);
    (AD_DATA[26] => U[40]) = (0:0:0, 0:0:0);
    (AD_DATA[26] => U[41]) = (0:0:0, 0:0:0);
    (AD_DATA[26] => U[42]) = (0:0:0, 0:0:0);
    (AD_DATA[26] => U[43]) = (0:0:0, 0:0:0);
    (AD_DATA[26] => V[26]) = (0:0:0, 0:0:0);
    (AD_DATA[26] => V[27]) = (0:0:0, 0:0:0);
    (AD_DATA[26] => V[28]) = (0:0:0, 0:0:0);
    (AD_DATA[26] => V[29]) = (0:0:0, 0:0:0);
    (AD_DATA[26] => V[30]) = (0:0:0, 0:0:0);
    (AD_DATA[26] => V[31]) = (0:0:0, 0:0:0);
    (AD_DATA[26] => V[32]) = (0:0:0, 0:0:0);
    (AD_DATA[26] => V[33]) = (0:0:0, 0:0:0);
    (AD_DATA[26] => V[34]) = (0:0:0, 0:0:0);
    (AD_DATA[26] => V[35]) = (0:0:0, 0:0:0);
    (AD_DATA[26] => V[36]) = (0:0:0, 0:0:0);
    (AD_DATA[26] => V[37]) = (0:0:0, 0:0:0);
    (AD_DATA[26] => V[38]) = (0:0:0, 0:0:0);
    (AD_DATA[26] => V[39]) = (0:0:0, 0:0:0);
    (AD_DATA[26] => V[40]) = (0:0:0, 0:0:0);
    (AD_DATA[26] => V[41]) = (0:0:0, 0:0:0);
    (AD_DATA[26] => V[42]) = (0:0:0, 0:0:0);
    (AD_DATA[26] => V[43]) = (0:0:0, 0:0:0);
    (AD_DATA[2] => U[10]) = (0:0:0, 0:0:0);
    (AD_DATA[2] => U[11]) = (0:0:0, 0:0:0);
    (AD_DATA[2] => U[12]) = (0:0:0, 0:0:0);
    (AD_DATA[2] => U[13]) = (0:0:0, 0:0:0);
    (AD_DATA[2] => U[14]) = (0:0:0, 0:0:0);
    (AD_DATA[2] => U[15]) = (0:0:0, 0:0:0);
    (AD_DATA[2] => U[16]) = (0:0:0, 0:0:0);
    (AD_DATA[2] => U[17]) = (0:0:0, 0:0:0);
    (AD_DATA[2] => U[18]) = (0:0:0, 0:0:0);
    (AD_DATA[2] => U[19]) = (0:0:0, 0:0:0);
    (AD_DATA[2] => U[20]) = (0:0:0, 0:0:0);
    (AD_DATA[2] => U[21]) = (0:0:0, 0:0:0);
    (AD_DATA[2] => U[22]) = (0:0:0, 0:0:0);
    (AD_DATA[2] => U[23]) = (0:0:0, 0:0:0);
    (AD_DATA[2] => U[24]) = (0:0:0, 0:0:0);
    (AD_DATA[2] => U[25]) = (0:0:0, 0:0:0);
    (AD_DATA[2] => U[26]) = (0:0:0, 0:0:0);
    (AD_DATA[2] => U[27]) = (0:0:0, 0:0:0);
    (AD_DATA[2] => U[28]) = (0:0:0, 0:0:0);
    (AD_DATA[2] => U[29]) = (0:0:0, 0:0:0);
    (AD_DATA[2] => U[2]) = (0:0:0, 0:0:0);
    (AD_DATA[2] => U[30]) = (0:0:0, 0:0:0);
    (AD_DATA[2] => U[31]) = (0:0:0, 0:0:0);
    (AD_DATA[2] => U[32]) = (0:0:0, 0:0:0);
    (AD_DATA[2] => U[33]) = (0:0:0, 0:0:0);
    (AD_DATA[2] => U[3]) = (0:0:0, 0:0:0);
    (AD_DATA[2] => U[4]) = (0:0:0, 0:0:0);
    (AD_DATA[2] => U[5]) = (0:0:0, 0:0:0);
    (AD_DATA[2] => U[6]) = (0:0:0, 0:0:0);
    (AD_DATA[2] => U[7]) = (0:0:0, 0:0:0);
    (AD_DATA[2] => U[8]) = (0:0:0, 0:0:0);
    (AD_DATA[2] => U[9]) = (0:0:0, 0:0:0);
    (AD_DATA[2] => V[10]) = (0:0:0, 0:0:0);
    (AD_DATA[2] => V[11]) = (0:0:0, 0:0:0);
    (AD_DATA[2] => V[12]) = (0:0:0, 0:0:0);
    (AD_DATA[2] => V[13]) = (0:0:0, 0:0:0);
    (AD_DATA[2] => V[14]) = (0:0:0, 0:0:0);
    (AD_DATA[2] => V[15]) = (0:0:0, 0:0:0);
    (AD_DATA[2] => V[16]) = (0:0:0, 0:0:0);
    (AD_DATA[2] => V[17]) = (0:0:0, 0:0:0);
    (AD_DATA[2] => V[18]) = (0:0:0, 0:0:0);
    (AD_DATA[2] => V[19]) = (0:0:0, 0:0:0);
    (AD_DATA[2] => V[20]) = (0:0:0, 0:0:0);
    (AD_DATA[2] => V[21]) = (0:0:0, 0:0:0);
    (AD_DATA[2] => V[22]) = (0:0:0, 0:0:0);
    (AD_DATA[2] => V[23]) = (0:0:0, 0:0:0);
    (AD_DATA[2] => V[24]) = (0:0:0, 0:0:0);
    (AD_DATA[2] => V[25]) = (0:0:0, 0:0:0);
    (AD_DATA[2] => V[26]) = (0:0:0, 0:0:0);
    (AD_DATA[2] => V[27]) = (0:0:0, 0:0:0);
    (AD_DATA[2] => V[28]) = (0:0:0, 0:0:0);
    (AD_DATA[2] => V[29]) = (0:0:0, 0:0:0);
    (AD_DATA[2] => V[30]) = (0:0:0, 0:0:0);
    (AD_DATA[2] => V[31]) = (0:0:0, 0:0:0);
    (AD_DATA[2] => V[32]) = (0:0:0, 0:0:0);
    (AD_DATA[2] => V[4]) = (0:0:0, 0:0:0);
    (AD_DATA[2] => V[5]) = (0:0:0, 0:0:0);
    (AD_DATA[2] => V[6]) = (0:0:0, 0:0:0);
    (AD_DATA[2] => V[7]) = (0:0:0, 0:0:0);
    (AD_DATA[2] => V[8]) = (0:0:0, 0:0:0);
    (AD_DATA[2] => V[9]) = (0:0:0, 0:0:0);
    (AD_DATA[3] => U[10]) = (0:0:0, 0:0:0);
    (AD_DATA[3] => U[11]) = (0:0:0, 0:0:0);
    (AD_DATA[3] => U[12]) = (0:0:0, 0:0:0);
    (AD_DATA[3] => U[13]) = (0:0:0, 0:0:0);
    (AD_DATA[3] => U[14]) = (0:0:0, 0:0:0);
    (AD_DATA[3] => U[15]) = (0:0:0, 0:0:0);
    (AD_DATA[3] => U[16]) = (0:0:0, 0:0:0);
    (AD_DATA[3] => U[17]) = (0:0:0, 0:0:0);
    (AD_DATA[3] => U[18]) = (0:0:0, 0:0:0);
    (AD_DATA[3] => U[19]) = (0:0:0, 0:0:0);
    (AD_DATA[3] => U[20]) = (0:0:0, 0:0:0);
    (AD_DATA[3] => U[21]) = (0:0:0, 0:0:0);
    (AD_DATA[3] => U[22]) = (0:0:0, 0:0:0);
    (AD_DATA[3] => U[23]) = (0:0:0, 0:0:0);
    (AD_DATA[3] => U[24]) = (0:0:0, 0:0:0);
    (AD_DATA[3] => U[25]) = (0:0:0, 0:0:0);
    (AD_DATA[3] => U[26]) = (0:0:0, 0:0:0);
    (AD_DATA[3] => U[27]) = (0:0:0, 0:0:0);
    (AD_DATA[3] => U[28]) = (0:0:0, 0:0:0);
    (AD_DATA[3] => U[29]) = (0:0:0, 0:0:0);
    (AD_DATA[3] => U[2]) = (0:0:0, 0:0:0);
    (AD_DATA[3] => U[30]) = (0:0:0, 0:0:0);
    (AD_DATA[3] => U[31]) = (0:0:0, 0:0:0);
    (AD_DATA[3] => U[32]) = (0:0:0, 0:0:0);
    (AD_DATA[3] => U[33]) = (0:0:0, 0:0:0);
    (AD_DATA[3] => U[34]) = (0:0:0, 0:0:0);
    (AD_DATA[3] => U[35]) = (0:0:0, 0:0:0);
    (AD_DATA[3] => U[3]) = (0:0:0, 0:0:0);
    (AD_DATA[3] => U[4]) = (0:0:0, 0:0:0);
    (AD_DATA[3] => U[5]) = (0:0:0, 0:0:0);
    (AD_DATA[3] => U[6]) = (0:0:0, 0:0:0);
    (AD_DATA[3] => U[7]) = (0:0:0, 0:0:0);
    (AD_DATA[3] => U[8]) = (0:0:0, 0:0:0);
    (AD_DATA[3] => U[9]) = (0:0:0, 0:0:0);
    (AD_DATA[3] => V[10]) = (0:0:0, 0:0:0);
    (AD_DATA[3] => V[11]) = (0:0:0, 0:0:0);
    (AD_DATA[3] => V[12]) = (0:0:0, 0:0:0);
    (AD_DATA[3] => V[13]) = (0:0:0, 0:0:0);
    (AD_DATA[3] => V[14]) = (0:0:0, 0:0:0);
    (AD_DATA[3] => V[15]) = (0:0:0, 0:0:0);
    (AD_DATA[3] => V[16]) = (0:0:0, 0:0:0);
    (AD_DATA[3] => V[17]) = (0:0:0, 0:0:0);
    (AD_DATA[3] => V[18]) = (0:0:0, 0:0:0);
    (AD_DATA[3] => V[19]) = (0:0:0, 0:0:0);
    (AD_DATA[3] => V[20]) = (0:0:0, 0:0:0);
    (AD_DATA[3] => V[21]) = (0:0:0, 0:0:0);
    (AD_DATA[3] => V[22]) = (0:0:0, 0:0:0);
    (AD_DATA[3] => V[23]) = (0:0:0, 0:0:0);
    (AD_DATA[3] => V[24]) = (0:0:0, 0:0:0);
    (AD_DATA[3] => V[25]) = (0:0:0, 0:0:0);
    (AD_DATA[3] => V[26]) = (0:0:0, 0:0:0);
    (AD_DATA[3] => V[27]) = (0:0:0, 0:0:0);
    (AD_DATA[3] => V[28]) = (0:0:0, 0:0:0);
    (AD_DATA[3] => V[29]) = (0:0:0, 0:0:0);
    (AD_DATA[3] => V[30]) = (0:0:0, 0:0:0);
    (AD_DATA[3] => V[31]) = (0:0:0, 0:0:0);
    (AD_DATA[3] => V[32]) = (0:0:0, 0:0:0);
    (AD_DATA[3] => V[33]) = (0:0:0, 0:0:0);
    (AD_DATA[3] => V[34]) = (0:0:0, 0:0:0);
    (AD_DATA[3] => V[4]) = (0:0:0, 0:0:0);
    (AD_DATA[3] => V[5]) = (0:0:0, 0:0:0);
    (AD_DATA[3] => V[6]) = (0:0:0, 0:0:0);
    (AD_DATA[3] => V[7]) = (0:0:0, 0:0:0);
    (AD_DATA[3] => V[8]) = (0:0:0, 0:0:0);
    (AD_DATA[3] => V[9]) = (0:0:0, 0:0:0);
    (AD_DATA[4] => U[10]) = (0:0:0, 0:0:0);
    (AD_DATA[4] => U[11]) = (0:0:0, 0:0:0);
    (AD_DATA[4] => U[12]) = (0:0:0, 0:0:0);
    (AD_DATA[4] => U[13]) = (0:0:0, 0:0:0);
    (AD_DATA[4] => U[14]) = (0:0:0, 0:0:0);
    (AD_DATA[4] => U[15]) = (0:0:0, 0:0:0);
    (AD_DATA[4] => U[16]) = (0:0:0, 0:0:0);
    (AD_DATA[4] => U[17]) = (0:0:0, 0:0:0);
    (AD_DATA[4] => U[18]) = (0:0:0, 0:0:0);
    (AD_DATA[4] => U[19]) = (0:0:0, 0:0:0);
    (AD_DATA[4] => U[20]) = (0:0:0, 0:0:0);
    (AD_DATA[4] => U[21]) = (0:0:0, 0:0:0);
    (AD_DATA[4] => U[22]) = (0:0:0, 0:0:0);
    (AD_DATA[4] => U[23]) = (0:0:0, 0:0:0);
    (AD_DATA[4] => U[24]) = (0:0:0, 0:0:0);
    (AD_DATA[4] => U[25]) = (0:0:0, 0:0:0);
    (AD_DATA[4] => U[26]) = (0:0:0, 0:0:0);
    (AD_DATA[4] => U[27]) = (0:0:0, 0:0:0);
    (AD_DATA[4] => U[28]) = (0:0:0, 0:0:0);
    (AD_DATA[4] => U[29]) = (0:0:0, 0:0:0);
    (AD_DATA[4] => U[30]) = (0:0:0, 0:0:0);
    (AD_DATA[4] => U[31]) = (0:0:0, 0:0:0);
    (AD_DATA[4] => U[32]) = (0:0:0, 0:0:0);
    (AD_DATA[4] => U[33]) = (0:0:0, 0:0:0);
    (AD_DATA[4] => U[34]) = (0:0:0, 0:0:0);
    (AD_DATA[4] => U[35]) = (0:0:0, 0:0:0);
    (AD_DATA[4] => U[5]) = (0:0:0, 0:0:0);
    (AD_DATA[4] => U[6]) = (0:0:0, 0:0:0);
    (AD_DATA[4] => U[7]) = (0:0:0, 0:0:0);
    (AD_DATA[4] => U[8]) = (0:0:0, 0:0:0);
    (AD_DATA[4] => U[9]) = (0:0:0, 0:0:0);
    (AD_DATA[4] => V[10]) = (0:0:0, 0:0:0);
    (AD_DATA[4] => V[11]) = (0:0:0, 0:0:0);
    (AD_DATA[4] => V[12]) = (0:0:0, 0:0:0);
    (AD_DATA[4] => V[13]) = (0:0:0, 0:0:0);
    (AD_DATA[4] => V[14]) = (0:0:0, 0:0:0);
    (AD_DATA[4] => V[15]) = (0:0:0, 0:0:0);
    (AD_DATA[4] => V[16]) = (0:0:0, 0:0:0);
    (AD_DATA[4] => V[17]) = (0:0:0, 0:0:0);
    (AD_DATA[4] => V[18]) = (0:0:0, 0:0:0);
    (AD_DATA[4] => V[19]) = (0:0:0, 0:0:0);
    (AD_DATA[4] => V[20]) = (0:0:0, 0:0:0);
    (AD_DATA[4] => V[21]) = (0:0:0, 0:0:0);
    (AD_DATA[4] => V[22]) = (0:0:0, 0:0:0);
    (AD_DATA[4] => V[23]) = (0:0:0, 0:0:0);
    (AD_DATA[4] => V[24]) = (0:0:0, 0:0:0);
    (AD_DATA[4] => V[25]) = (0:0:0, 0:0:0);
    (AD_DATA[4] => V[26]) = (0:0:0, 0:0:0);
    (AD_DATA[4] => V[27]) = (0:0:0, 0:0:0);
    (AD_DATA[4] => V[28]) = (0:0:0, 0:0:0);
    (AD_DATA[4] => V[29]) = (0:0:0, 0:0:0);
    (AD_DATA[4] => V[30]) = (0:0:0, 0:0:0);
    (AD_DATA[4] => V[31]) = (0:0:0, 0:0:0);
    (AD_DATA[4] => V[32]) = (0:0:0, 0:0:0);
    (AD_DATA[4] => V[33]) = (0:0:0, 0:0:0);
    (AD_DATA[4] => V[34]) = (0:0:0, 0:0:0);
    (AD_DATA[4] => V[4]) = (0:0:0, 0:0:0);
    (AD_DATA[4] => V[5]) = (0:0:0, 0:0:0);
    (AD_DATA[4] => V[6]) = (0:0:0, 0:0:0);
    (AD_DATA[4] => V[7]) = (0:0:0, 0:0:0);
    (AD_DATA[4] => V[8]) = (0:0:0, 0:0:0);
    (AD_DATA[4] => V[9]) = (0:0:0, 0:0:0);
    (AD_DATA[5] => U[10]) = (0:0:0, 0:0:0);
    (AD_DATA[5] => U[11]) = (0:0:0, 0:0:0);
    (AD_DATA[5] => U[12]) = (0:0:0, 0:0:0);
    (AD_DATA[5] => U[13]) = (0:0:0, 0:0:0);
    (AD_DATA[5] => U[14]) = (0:0:0, 0:0:0);
    (AD_DATA[5] => U[15]) = (0:0:0, 0:0:0);
    (AD_DATA[5] => U[16]) = (0:0:0, 0:0:0);
    (AD_DATA[5] => U[17]) = (0:0:0, 0:0:0);
    (AD_DATA[5] => U[18]) = (0:0:0, 0:0:0);
    (AD_DATA[5] => U[19]) = (0:0:0, 0:0:0);
    (AD_DATA[5] => U[20]) = (0:0:0, 0:0:0);
    (AD_DATA[5] => U[21]) = (0:0:0, 0:0:0);
    (AD_DATA[5] => U[22]) = (0:0:0, 0:0:0);
    (AD_DATA[5] => U[23]) = (0:0:0, 0:0:0);
    (AD_DATA[5] => U[24]) = (0:0:0, 0:0:0);
    (AD_DATA[5] => U[25]) = (0:0:0, 0:0:0);
    (AD_DATA[5] => U[26]) = (0:0:0, 0:0:0);
    (AD_DATA[5] => U[27]) = (0:0:0, 0:0:0);
    (AD_DATA[5] => U[28]) = (0:0:0, 0:0:0);
    (AD_DATA[5] => U[29]) = (0:0:0, 0:0:0);
    (AD_DATA[5] => U[30]) = (0:0:0, 0:0:0);
    (AD_DATA[5] => U[31]) = (0:0:0, 0:0:0);
    (AD_DATA[5] => U[32]) = (0:0:0, 0:0:0);
    (AD_DATA[5] => U[33]) = (0:0:0, 0:0:0);
    (AD_DATA[5] => U[34]) = (0:0:0, 0:0:0);
    (AD_DATA[5] => U[35]) = (0:0:0, 0:0:0);
    (AD_DATA[5] => U[36]) = (0:0:0, 0:0:0);
    (AD_DATA[5] => U[5]) = (0:0:0, 0:0:0);
    (AD_DATA[5] => U[6]) = (0:0:0, 0:0:0);
    (AD_DATA[5] => U[7]) = (0:0:0, 0:0:0);
    (AD_DATA[5] => U[8]) = (0:0:0, 0:0:0);
    (AD_DATA[5] => U[9]) = (0:0:0, 0:0:0);
    (AD_DATA[5] => V[10]) = (0:0:0, 0:0:0);
    (AD_DATA[5] => V[11]) = (0:0:0, 0:0:0);
    (AD_DATA[5] => V[12]) = (0:0:0, 0:0:0);
    (AD_DATA[5] => V[13]) = (0:0:0, 0:0:0);
    (AD_DATA[5] => V[14]) = (0:0:0, 0:0:0);
    (AD_DATA[5] => V[15]) = (0:0:0, 0:0:0);
    (AD_DATA[5] => V[16]) = (0:0:0, 0:0:0);
    (AD_DATA[5] => V[17]) = (0:0:0, 0:0:0);
    (AD_DATA[5] => V[18]) = (0:0:0, 0:0:0);
    (AD_DATA[5] => V[19]) = (0:0:0, 0:0:0);
    (AD_DATA[5] => V[20]) = (0:0:0, 0:0:0);
    (AD_DATA[5] => V[21]) = (0:0:0, 0:0:0);
    (AD_DATA[5] => V[22]) = (0:0:0, 0:0:0);
    (AD_DATA[5] => V[23]) = (0:0:0, 0:0:0);
    (AD_DATA[5] => V[24]) = (0:0:0, 0:0:0);
    (AD_DATA[5] => V[25]) = (0:0:0, 0:0:0);
    (AD_DATA[5] => V[26]) = (0:0:0, 0:0:0);
    (AD_DATA[5] => V[27]) = (0:0:0, 0:0:0);
    (AD_DATA[5] => V[28]) = (0:0:0, 0:0:0);
    (AD_DATA[5] => V[29]) = (0:0:0, 0:0:0);
    (AD_DATA[5] => V[30]) = (0:0:0, 0:0:0);
    (AD_DATA[5] => V[31]) = (0:0:0, 0:0:0);
    (AD_DATA[5] => V[32]) = (0:0:0, 0:0:0);
    (AD_DATA[5] => V[33]) = (0:0:0, 0:0:0);
    (AD_DATA[5] => V[34]) = (0:0:0, 0:0:0);
    (AD_DATA[5] => V[35]) = (0:0:0, 0:0:0);
    (AD_DATA[5] => V[4]) = (0:0:0, 0:0:0);
    (AD_DATA[5] => V[5]) = (0:0:0, 0:0:0);
    (AD_DATA[5] => V[6]) = (0:0:0, 0:0:0);
    (AD_DATA[5] => V[7]) = (0:0:0, 0:0:0);
    (AD_DATA[5] => V[8]) = (0:0:0, 0:0:0);
    (AD_DATA[5] => V[9]) = (0:0:0, 0:0:0);
    (AD_DATA[6] => U[10]) = (0:0:0, 0:0:0);
    (AD_DATA[6] => U[11]) = (0:0:0, 0:0:0);
    (AD_DATA[6] => U[12]) = (0:0:0, 0:0:0);
    (AD_DATA[6] => U[13]) = (0:0:0, 0:0:0);
    (AD_DATA[6] => U[14]) = (0:0:0, 0:0:0);
    (AD_DATA[6] => U[15]) = (0:0:0, 0:0:0);
    (AD_DATA[6] => U[16]) = (0:0:0, 0:0:0);
    (AD_DATA[6] => U[17]) = (0:0:0, 0:0:0);
    (AD_DATA[6] => U[18]) = (0:0:0, 0:0:0);
    (AD_DATA[6] => U[19]) = (0:0:0, 0:0:0);
    (AD_DATA[6] => U[20]) = (0:0:0, 0:0:0);
    (AD_DATA[6] => U[21]) = (0:0:0, 0:0:0);
    (AD_DATA[6] => U[22]) = (0:0:0, 0:0:0);
    (AD_DATA[6] => U[23]) = (0:0:0, 0:0:0);
    (AD_DATA[6] => U[24]) = (0:0:0, 0:0:0);
    (AD_DATA[6] => U[25]) = (0:0:0, 0:0:0);
    (AD_DATA[6] => U[26]) = (0:0:0, 0:0:0);
    (AD_DATA[6] => U[27]) = (0:0:0, 0:0:0);
    (AD_DATA[6] => U[28]) = (0:0:0, 0:0:0);
    (AD_DATA[6] => U[29]) = (0:0:0, 0:0:0);
    (AD_DATA[6] => U[30]) = (0:0:0, 0:0:0);
    (AD_DATA[6] => U[31]) = (0:0:0, 0:0:0);
    (AD_DATA[6] => U[32]) = (0:0:0, 0:0:0);
    (AD_DATA[6] => U[33]) = (0:0:0, 0:0:0);
    (AD_DATA[6] => U[34]) = (0:0:0, 0:0:0);
    (AD_DATA[6] => U[35]) = (0:0:0, 0:0:0);
    (AD_DATA[6] => U[36]) = (0:0:0, 0:0:0);
    (AD_DATA[6] => U[7]) = (0:0:0, 0:0:0);
    (AD_DATA[6] => U[8]) = (0:0:0, 0:0:0);
    (AD_DATA[6] => U[9]) = (0:0:0, 0:0:0);
    (AD_DATA[6] => V[10]) = (0:0:0, 0:0:0);
    (AD_DATA[6] => V[11]) = (0:0:0, 0:0:0);
    (AD_DATA[6] => V[12]) = (0:0:0, 0:0:0);
    (AD_DATA[6] => V[13]) = (0:0:0, 0:0:0);
    (AD_DATA[6] => V[14]) = (0:0:0, 0:0:0);
    (AD_DATA[6] => V[15]) = (0:0:0, 0:0:0);
    (AD_DATA[6] => V[16]) = (0:0:0, 0:0:0);
    (AD_DATA[6] => V[17]) = (0:0:0, 0:0:0);
    (AD_DATA[6] => V[18]) = (0:0:0, 0:0:0);
    (AD_DATA[6] => V[19]) = (0:0:0, 0:0:0);
    (AD_DATA[6] => V[20]) = (0:0:0, 0:0:0);
    (AD_DATA[6] => V[21]) = (0:0:0, 0:0:0);
    (AD_DATA[6] => V[22]) = (0:0:0, 0:0:0);
    (AD_DATA[6] => V[23]) = (0:0:0, 0:0:0);
    (AD_DATA[6] => V[24]) = (0:0:0, 0:0:0);
    (AD_DATA[6] => V[25]) = (0:0:0, 0:0:0);
    (AD_DATA[6] => V[26]) = (0:0:0, 0:0:0);
    (AD_DATA[6] => V[27]) = (0:0:0, 0:0:0);
    (AD_DATA[6] => V[28]) = (0:0:0, 0:0:0);
    (AD_DATA[6] => V[29]) = (0:0:0, 0:0:0);
    (AD_DATA[6] => V[30]) = (0:0:0, 0:0:0);
    (AD_DATA[6] => V[31]) = (0:0:0, 0:0:0);
    (AD_DATA[6] => V[32]) = (0:0:0, 0:0:0);
    (AD_DATA[6] => V[33]) = (0:0:0, 0:0:0);
    (AD_DATA[6] => V[34]) = (0:0:0, 0:0:0);
    (AD_DATA[6] => V[35]) = (0:0:0, 0:0:0);
    (AD_DATA[6] => V[6]) = (0:0:0, 0:0:0);
    (AD_DATA[6] => V[7]) = (0:0:0, 0:0:0);
    (AD_DATA[6] => V[8]) = (0:0:0, 0:0:0);
    (AD_DATA[6] => V[9]) = (0:0:0, 0:0:0);
    (AD_DATA[7] => U[10]) = (0:0:0, 0:0:0);
    (AD_DATA[7] => U[11]) = (0:0:0, 0:0:0);
    (AD_DATA[7] => U[12]) = (0:0:0, 0:0:0);
    (AD_DATA[7] => U[13]) = (0:0:0, 0:0:0);
    (AD_DATA[7] => U[14]) = (0:0:0, 0:0:0);
    (AD_DATA[7] => U[15]) = (0:0:0, 0:0:0);
    (AD_DATA[7] => U[16]) = (0:0:0, 0:0:0);
    (AD_DATA[7] => U[17]) = (0:0:0, 0:0:0);
    (AD_DATA[7] => U[18]) = (0:0:0, 0:0:0);
    (AD_DATA[7] => U[19]) = (0:0:0, 0:0:0);
    (AD_DATA[7] => U[20]) = (0:0:0, 0:0:0);
    (AD_DATA[7] => U[21]) = (0:0:0, 0:0:0);
    (AD_DATA[7] => U[22]) = (0:0:0, 0:0:0);
    (AD_DATA[7] => U[23]) = (0:0:0, 0:0:0);
    (AD_DATA[7] => U[24]) = (0:0:0, 0:0:0);
    (AD_DATA[7] => U[25]) = (0:0:0, 0:0:0);
    (AD_DATA[7] => U[26]) = (0:0:0, 0:0:0);
    (AD_DATA[7] => U[27]) = (0:0:0, 0:0:0);
    (AD_DATA[7] => U[28]) = (0:0:0, 0:0:0);
    (AD_DATA[7] => U[29]) = (0:0:0, 0:0:0);
    (AD_DATA[7] => U[30]) = (0:0:0, 0:0:0);
    (AD_DATA[7] => U[31]) = (0:0:0, 0:0:0);
    (AD_DATA[7] => U[32]) = (0:0:0, 0:0:0);
    (AD_DATA[7] => U[33]) = (0:0:0, 0:0:0);
    (AD_DATA[7] => U[34]) = (0:0:0, 0:0:0);
    (AD_DATA[7] => U[35]) = (0:0:0, 0:0:0);
    (AD_DATA[7] => U[36]) = (0:0:0, 0:0:0);
    (AD_DATA[7] => U[37]) = (0:0:0, 0:0:0);
    (AD_DATA[7] => U[38]) = (0:0:0, 0:0:0);
    (AD_DATA[7] => U[7]) = (0:0:0, 0:0:0);
    (AD_DATA[7] => U[8]) = (0:0:0, 0:0:0);
    (AD_DATA[7] => U[9]) = (0:0:0, 0:0:0);
    (AD_DATA[7] => V[10]) = (0:0:0, 0:0:0);
    (AD_DATA[7] => V[11]) = (0:0:0, 0:0:0);
    (AD_DATA[7] => V[12]) = (0:0:0, 0:0:0);
    (AD_DATA[7] => V[13]) = (0:0:0, 0:0:0);
    (AD_DATA[7] => V[14]) = (0:0:0, 0:0:0);
    (AD_DATA[7] => V[15]) = (0:0:0, 0:0:0);
    (AD_DATA[7] => V[16]) = (0:0:0, 0:0:0);
    (AD_DATA[7] => V[17]) = (0:0:0, 0:0:0);
    (AD_DATA[7] => V[18]) = (0:0:0, 0:0:0);
    (AD_DATA[7] => V[19]) = (0:0:0, 0:0:0);
    (AD_DATA[7] => V[20]) = (0:0:0, 0:0:0);
    (AD_DATA[7] => V[21]) = (0:0:0, 0:0:0);
    (AD_DATA[7] => V[22]) = (0:0:0, 0:0:0);
    (AD_DATA[7] => V[23]) = (0:0:0, 0:0:0);
    (AD_DATA[7] => V[24]) = (0:0:0, 0:0:0);
    (AD_DATA[7] => V[25]) = (0:0:0, 0:0:0);
    (AD_DATA[7] => V[26]) = (0:0:0, 0:0:0);
    (AD_DATA[7] => V[27]) = (0:0:0, 0:0:0);
    (AD_DATA[7] => V[28]) = (0:0:0, 0:0:0);
    (AD_DATA[7] => V[29]) = (0:0:0, 0:0:0);
    (AD_DATA[7] => V[30]) = (0:0:0, 0:0:0);
    (AD_DATA[7] => V[31]) = (0:0:0, 0:0:0);
    (AD_DATA[7] => V[32]) = (0:0:0, 0:0:0);
    (AD_DATA[7] => V[33]) = (0:0:0, 0:0:0);
    (AD_DATA[7] => V[34]) = (0:0:0, 0:0:0);
    (AD_DATA[7] => V[35]) = (0:0:0, 0:0:0);
    (AD_DATA[7] => V[36]) = (0:0:0, 0:0:0);
    (AD_DATA[7] => V[37]) = (0:0:0, 0:0:0);
    (AD_DATA[7] => V[6]) = (0:0:0, 0:0:0);
    (AD_DATA[7] => V[7]) = (0:0:0, 0:0:0);
    (AD_DATA[7] => V[8]) = (0:0:0, 0:0:0);
    (AD_DATA[7] => V[9]) = (0:0:0, 0:0:0);
    (AD_DATA[8] => U[10]) = (0:0:0, 0:0:0);
    (AD_DATA[8] => U[11]) = (0:0:0, 0:0:0);
    (AD_DATA[8] => U[12]) = (0:0:0, 0:0:0);
    (AD_DATA[8] => U[13]) = (0:0:0, 0:0:0);
    (AD_DATA[8] => U[14]) = (0:0:0, 0:0:0);
    (AD_DATA[8] => U[15]) = (0:0:0, 0:0:0);
    (AD_DATA[8] => U[16]) = (0:0:0, 0:0:0);
    (AD_DATA[8] => U[17]) = (0:0:0, 0:0:0);
    (AD_DATA[8] => U[18]) = (0:0:0, 0:0:0);
    (AD_DATA[8] => U[19]) = (0:0:0, 0:0:0);
    (AD_DATA[8] => U[20]) = (0:0:0, 0:0:0);
    (AD_DATA[8] => U[21]) = (0:0:0, 0:0:0);
    (AD_DATA[8] => U[22]) = (0:0:0, 0:0:0);
    (AD_DATA[8] => U[23]) = (0:0:0, 0:0:0);
    (AD_DATA[8] => U[24]) = (0:0:0, 0:0:0);
    (AD_DATA[8] => U[25]) = (0:0:0, 0:0:0);
    (AD_DATA[8] => U[26]) = (0:0:0, 0:0:0);
    (AD_DATA[8] => U[27]) = (0:0:0, 0:0:0);
    (AD_DATA[8] => U[28]) = (0:0:0, 0:0:0);
    (AD_DATA[8] => U[29]) = (0:0:0, 0:0:0);
    (AD_DATA[8] => U[30]) = (0:0:0, 0:0:0);
    (AD_DATA[8] => U[31]) = (0:0:0, 0:0:0);
    (AD_DATA[8] => U[32]) = (0:0:0, 0:0:0);
    (AD_DATA[8] => U[33]) = (0:0:0, 0:0:0);
    (AD_DATA[8] => U[34]) = (0:0:0, 0:0:0);
    (AD_DATA[8] => U[35]) = (0:0:0, 0:0:0);
    (AD_DATA[8] => U[36]) = (0:0:0, 0:0:0);
    (AD_DATA[8] => U[37]) = (0:0:0, 0:0:0);
    (AD_DATA[8] => U[38]) = (0:0:0, 0:0:0);
    (AD_DATA[8] => U[9]) = (0:0:0, 0:0:0);
    (AD_DATA[8] => V[10]) = (0:0:0, 0:0:0);
    (AD_DATA[8] => V[11]) = (0:0:0, 0:0:0);
    (AD_DATA[8] => V[12]) = (0:0:0, 0:0:0);
    (AD_DATA[8] => V[13]) = (0:0:0, 0:0:0);
    (AD_DATA[8] => V[14]) = (0:0:0, 0:0:0);
    (AD_DATA[8] => V[15]) = (0:0:0, 0:0:0);
    (AD_DATA[8] => V[16]) = (0:0:0, 0:0:0);
    (AD_DATA[8] => V[17]) = (0:0:0, 0:0:0);
    (AD_DATA[8] => V[18]) = (0:0:0, 0:0:0);
    (AD_DATA[8] => V[19]) = (0:0:0, 0:0:0);
    (AD_DATA[8] => V[20]) = (0:0:0, 0:0:0);
    (AD_DATA[8] => V[21]) = (0:0:0, 0:0:0);
    (AD_DATA[8] => V[22]) = (0:0:0, 0:0:0);
    (AD_DATA[8] => V[23]) = (0:0:0, 0:0:0);
    (AD_DATA[8] => V[24]) = (0:0:0, 0:0:0);
    (AD_DATA[8] => V[25]) = (0:0:0, 0:0:0);
    (AD_DATA[8] => V[26]) = (0:0:0, 0:0:0);
    (AD_DATA[8] => V[27]) = (0:0:0, 0:0:0);
    (AD_DATA[8] => V[28]) = (0:0:0, 0:0:0);
    (AD_DATA[8] => V[29]) = (0:0:0, 0:0:0);
    (AD_DATA[8] => V[30]) = (0:0:0, 0:0:0);
    (AD_DATA[8] => V[31]) = (0:0:0, 0:0:0);
    (AD_DATA[8] => V[32]) = (0:0:0, 0:0:0);
    (AD_DATA[8] => V[33]) = (0:0:0, 0:0:0);
    (AD_DATA[8] => V[34]) = (0:0:0, 0:0:0);
    (AD_DATA[8] => V[35]) = (0:0:0, 0:0:0);
    (AD_DATA[8] => V[36]) = (0:0:0, 0:0:0);
    (AD_DATA[8] => V[37]) = (0:0:0, 0:0:0);
    (AD_DATA[8] => V[8]) = (0:0:0, 0:0:0);
    (AD_DATA[8] => V[9]) = (0:0:0, 0:0:0);
    (AD_DATA[9] => U[10]) = (0:0:0, 0:0:0);
    (AD_DATA[9] => U[11]) = (0:0:0, 0:0:0);
    (AD_DATA[9] => U[12]) = (0:0:0, 0:0:0);
    (AD_DATA[9] => U[13]) = (0:0:0, 0:0:0);
    (AD_DATA[9] => U[14]) = (0:0:0, 0:0:0);
    (AD_DATA[9] => U[15]) = (0:0:0, 0:0:0);
    (AD_DATA[9] => U[16]) = (0:0:0, 0:0:0);
    (AD_DATA[9] => U[17]) = (0:0:0, 0:0:0);
    (AD_DATA[9] => U[18]) = (0:0:0, 0:0:0);
    (AD_DATA[9] => U[19]) = (0:0:0, 0:0:0);
    (AD_DATA[9] => U[20]) = (0:0:0, 0:0:0);
    (AD_DATA[9] => U[21]) = (0:0:0, 0:0:0);
    (AD_DATA[9] => U[22]) = (0:0:0, 0:0:0);
    (AD_DATA[9] => U[23]) = (0:0:0, 0:0:0);
    (AD_DATA[9] => U[24]) = (0:0:0, 0:0:0);
    (AD_DATA[9] => U[25]) = (0:0:0, 0:0:0);
    (AD_DATA[9] => U[26]) = (0:0:0, 0:0:0);
    (AD_DATA[9] => U[27]) = (0:0:0, 0:0:0);
    (AD_DATA[9] => U[28]) = (0:0:0, 0:0:0);
    (AD_DATA[9] => U[29]) = (0:0:0, 0:0:0);
    (AD_DATA[9] => U[30]) = (0:0:0, 0:0:0);
    (AD_DATA[9] => U[31]) = (0:0:0, 0:0:0);
    (AD_DATA[9] => U[32]) = (0:0:0, 0:0:0);
    (AD_DATA[9] => U[33]) = (0:0:0, 0:0:0);
    (AD_DATA[9] => U[34]) = (0:0:0, 0:0:0);
    (AD_DATA[9] => U[35]) = (0:0:0, 0:0:0);
    (AD_DATA[9] => U[36]) = (0:0:0, 0:0:0);
    (AD_DATA[9] => U[37]) = (0:0:0, 0:0:0);
    (AD_DATA[9] => U[38]) = (0:0:0, 0:0:0);
    (AD_DATA[9] => U[39]) = (0:0:0, 0:0:0);
    (AD_DATA[9] => U[40]) = (0:0:0, 0:0:0);
    (AD_DATA[9] => U[9]) = (0:0:0, 0:0:0);
    (AD_DATA[9] => V[10]) = (0:0:0, 0:0:0);
    (AD_DATA[9] => V[11]) = (0:0:0, 0:0:0);
    (AD_DATA[9] => V[12]) = (0:0:0, 0:0:0);
    (AD_DATA[9] => V[13]) = (0:0:0, 0:0:0);
    (AD_DATA[9] => V[14]) = (0:0:0, 0:0:0);
    (AD_DATA[9] => V[15]) = (0:0:0, 0:0:0);
    (AD_DATA[9] => V[16]) = (0:0:0, 0:0:0);
    (AD_DATA[9] => V[17]) = (0:0:0, 0:0:0);
    (AD_DATA[9] => V[18]) = (0:0:0, 0:0:0);
    (AD_DATA[9] => V[19]) = (0:0:0, 0:0:0);
    (AD_DATA[9] => V[20]) = (0:0:0, 0:0:0);
    (AD_DATA[9] => V[21]) = (0:0:0, 0:0:0);
    (AD_DATA[9] => V[22]) = (0:0:0, 0:0:0);
    (AD_DATA[9] => V[23]) = (0:0:0, 0:0:0);
    (AD_DATA[9] => V[24]) = (0:0:0, 0:0:0);
    (AD_DATA[9] => V[25]) = (0:0:0, 0:0:0);
    (AD_DATA[9] => V[26]) = (0:0:0, 0:0:0);
    (AD_DATA[9] => V[27]) = (0:0:0, 0:0:0);
    (AD_DATA[9] => V[28]) = (0:0:0, 0:0:0);
    (AD_DATA[9] => V[29]) = (0:0:0, 0:0:0);
    (AD_DATA[9] => V[30]) = (0:0:0, 0:0:0);
    (AD_DATA[9] => V[31]) = (0:0:0, 0:0:0);
    (AD_DATA[9] => V[32]) = (0:0:0, 0:0:0);
    (AD_DATA[9] => V[33]) = (0:0:0, 0:0:0);
    (AD_DATA[9] => V[34]) = (0:0:0, 0:0:0);
    (AD_DATA[9] => V[35]) = (0:0:0, 0:0:0);
    (AD_DATA[9] => V[36]) = (0:0:0, 0:0:0);
    (AD_DATA[9] => V[37]) = (0:0:0, 0:0:0);
    (AD_DATA[9] => V[38]) = (0:0:0, 0:0:0);
    (AD_DATA[9] => V[39]) = (0:0:0, 0:0:0);
    (AD_DATA[9] => V[8]) = (0:0:0, 0:0:0);
    (AD_DATA[9] => V[9]) = (0:0:0, 0:0:0);
    (B2B1[0] => U[10]) = (0:0:0, 0:0:0);
    (B2B1[0] => U[11]) = (0:0:0, 0:0:0);
    (B2B1[0] => U[12]) = (0:0:0, 0:0:0);
    (B2B1[0] => U[13]) = (0:0:0, 0:0:0);
    (B2B1[0] => U[14]) = (0:0:0, 0:0:0);
    (B2B1[0] => U[15]) = (0:0:0, 0:0:0);
    (B2B1[0] => U[16]) = (0:0:0, 0:0:0);
    (B2B1[0] => U[17]) = (0:0:0, 0:0:0);
    (B2B1[0] => U[18]) = (0:0:0, 0:0:0);
    (B2B1[0] => U[19]) = (0:0:0, 0:0:0);
    (B2B1[0] => U[1]) = (0:0:0, 0:0:0);
    (B2B1[0] => U[20]) = (0:0:0, 0:0:0);
    (B2B1[0] => U[21]) = (0:0:0, 0:0:0);
    (B2B1[0] => U[22]) = (0:0:0, 0:0:0);
    (B2B1[0] => U[23]) = (0:0:0, 0:0:0);
    (B2B1[0] => U[24]) = (0:0:0, 0:0:0);
    (B2B1[0] => U[25]) = (0:0:0, 0:0:0);
    (B2B1[0] => U[26]) = (0:0:0, 0:0:0);
    (B2B1[0] => U[27]) = (0:0:0, 0:0:0);
    (B2B1[0] => U[28]) = (0:0:0, 0:0:0);
    (B2B1[0] => U[29]) = (0:0:0, 0:0:0);
    (B2B1[0] => U[2]) = (0:0:0, 0:0:0);
    (B2B1[0] => U[30]) = (0:0:0, 0:0:0);
    (B2B1[0] => U[31]) = (0:0:0, 0:0:0);
    (B2B1[0] => U[3]) = (0:0:0, 0:0:0);
    (B2B1[0] => U[4]) = (0:0:0, 0:0:0);
    (B2B1[0] => U[5]) = (0:0:0, 0:0:0);
    (B2B1[0] => U[6]) = (0:0:0, 0:0:0);
    (B2B1[0] => U[7]) = (0:0:0, 0:0:0);
    (B2B1[0] => U[8]) = (0:0:0, 0:0:0);
    (B2B1[0] => U[9]) = (0:0:0, 0:0:0);
    (B2B1[0] => V[0]) = (0:0:0, 0:0:0);
    (B2B1[0] => V[10]) = (0:0:0, 0:0:0);
    (B2B1[0] => V[11]) = (0:0:0, 0:0:0);
    (B2B1[0] => V[12]) = (0:0:0, 0:0:0);
    (B2B1[0] => V[13]) = (0:0:0, 0:0:0);
    (B2B1[0] => V[14]) = (0:0:0, 0:0:0);
    (B2B1[0] => V[15]) = (0:0:0, 0:0:0);
    (B2B1[0] => V[16]) = (0:0:0, 0:0:0);
    (B2B1[0] => V[17]) = (0:0:0, 0:0:0);
    (B2B1[0] => V[18]) = (0:0:0, 0:0:0);
    (B2B1[0] => V[19]) = (0:0:0, 0:0:0);
    (B2B1[0] => V[20]) = (0:0:0, 0:0:0);
    (B2B1[0] => V[21]) = (0:0:0, 0:0:0);
    (B2B1[0] => V[22]) = (0:0:0, 0:0:0);
    (B2B1[0] => V[23]) = (0:0:0, 0:0:0);
    (B2B1[0] => V[24]) = (0:0:0, 0:0:0);
    (B2B1[0] => V[25]) = (0:0:0, 0:0:0);
    (B2B1[0] => V[26]) = (0:0:0, 0:0:0);
    (B2B1[0] => V[27]) = (0:0:0, 0:0:0);
    (B2B1[0] => V[28]) = (0:0:0, 0:0:0);
    (B2B1[0] => V[29]) = (0:0:0, 0:0:0);
    (B2B1[0] => V[30]) = (0:0:0, 0:0:0);
    (B2B1[0] => V[4]) = (0:0:0, 0:0:0);
    (B2B1[0] => V[5]) = (0:0:0, 0:0:0);
    (B2B1[0] => V[6]) = (0:0:0, 0:0:0);
    (B2B1[0] => V[7]) = (0:0:0, 0:0:0);
    (B2B1[0] => V[8]) = (0:0:0, 0:0:0);
    (B2B1[0] => V[9]) = (0:0:0, 0:0:0);
    (B2B1[10] => U[11]) = (0:0:0, 0:0:0);
    (B2B1[10] => U[12]) = (0:0:0, 0:0:0);
    (B2B1[10] => U[13]) = (0:0:0, 0:0:0);
    (B2B1[10] => U[14]) = (0:0:0, 0:0:0);
    (B2B1[10] => U[15]) = (0:0:0, 0:0:0);
    (B2B1[10] => U[16]) = (0:0:0, 0:0:0);
    (B2B1[10] => U[17]) = (0:0:0, 0:0:0);
    (B2B1[10] => U[18]) = (0:0:0, 0:0:0);
    (B2B1[10] => U[19]) = (0:0:0, 0:0:0);
    (B2B1[10] => U[20]) = (0:0:0, 0:0:0);
    (B2B1[10] => U[21]) = (0:0:0, 0:0:0);
    (B2B1[10] => U[22]) = (0:0:0, 0:0:0);
    (B2B1[10] => U[23]) = (0:0:0, 0:0:0);
    (B2B1[10] => U[24]) = (0:0:0, 0:0:0);
    (B2B1[10] => U[25]) = (0:0:0, 0:0:0);
    (B2B1[10] => U[26]) = (0:0:0, 0:0:0);
    (B2B1[10] => U[27]) = (0:0:0, 0:0:0);
    (B2B1[10] => U[28]) = (0:0:0, 0:0:0);
    (B2B1[10] => U[29]) = (0:0:0, 0:0:0);
    (B2B1[10] => U[30]) = (0:0:0, 0:0:0);
    (B2B1[10] => U[31]) = (0:0:0, 0:0:0);
    (B2B1[10] => U[32]) = (0:0:0, 0:0:0);
    (B2B1[10] => U[33]) = (0:0:0, 0:0:0);
    (B2B1[10] => U[34]) = (0:0:0, 0:0:0);
    (B2B1[10] => U[35]) = (0:0:0, 0:0:0);
    (B2B1[10] => U[36]) = (0:0:0, 0:0:0);
    (B2B1[10] => U[37]) = (0:0:0, 0:0:0);
    (B2B1[10] => U[38]) = (0:0:0, 0:0:0);
    (B2B1[10] => U[39]) = (0:0:0, 0:0:0);
    (B2B1[10] => U[40]) = (0:0:0, 0:0:0);
    (B2B1[10] => V[10]) = (0:0:0, 0:0:0);
    (B2B1[10] => V[11]) = (0:0:0, 0:0:0);
    (B2B1[10] => V[12]) = (0:0:0, 0:0:0);
    (B2B1[10] => V[13]) = (0:0:0, 0:0:0);
    (B2B1[10] => V[14]) = (0:0:0, 0:0:0);
    (B2B1[10] => V[15]) = (0:0:0, 0:0:0);
    (B2B1[10] => V[16]) = (0:0:0, 0:0:0);
    (B2B1[10] => V[17]) = (0:0:0, 0:0:0);
    (B2B1[10] => V[18]) = (0:0:0, 0:0:0);
    (B2B1[10] => V[19]) = (0:0:0, 0:0:0);
    (B2B1[10] => V[20]) = (0:0:0, 0:0:0);
    (B2B1[10] => V[21]) = (0:0:0, 0:0:0);
    (B2B1[10] => V[22]) = (0:0:0, 0:0:0);
    (B2B1[10] => V[23]) = (0:0:0, 0:0:0);
    (B2B1[10] => V[24]) = (0:0:0, 0:0:0);
    (B2B1[10] => V[25]) = (0:0:0, 0:0:0);
    (B2B1[10] => V[26]) = (0:0:0, 0:0:0);
    (B2B1[10] => V[27]) = (0:0:0, 0:0:0);
    (B2B1[10] => V[28]) = (0:0:0, 0:0:0);
    (B2B1[10] => V[29]) = (0:0:0, 0:0:0);
    (B2B1[10] => V[30]) = (0:0:0, 0:0:0);
    (B2B1[10] => V[31]) = (0:0:0, 0:0:0);
    (B2B1[10] => V[32]) = (0:0:0, 0:0:0);
    (B2B1[10] => V[33]) = (0:0:0, 0:0:0);
    (B2B1[10] => V[34]) = (0:0:0, 0:0:0);
    (B2B1[10] => V[35]) = (0:0:0, 0:0:0);
    (B2B1[10] => V[36]) = (0:0:0, 0:0:0);
    (B2B1[10] => V[37]) = (0:0:0, 0:0:0);
    (B2B1[10] => V[38]) = (0:0:0, 0:0:0);
    (B2B1[10] => V[39]) = (0:0:0, 0:0:0);
    (B2B1[11] => U[11]) = (0:0:0, 0:0:0);
    (B2B1[11] => U[12]) = (0:0:0, 0:0:0);
    (B2B1[11] => U[13]) = (0:0:0, 0:0:0);
    (B2B1[11] => U[14]) = (0:0:0, 0:0:0);
    (B2B1[11] => U[15]) = (0:0:0, 0:0:0);
    (B2B1[11] => U[16]) = (0:0:0, 0:0:0);
    (B2B1[11] => U[17]) = (0:0:0, 0:0:0);
    (B2B1[11] => U[18]) = (0:0:0, 0:0:0);
    (B2B1[11] => U[19]) = (0:0:0, 0:0:0);
    (B2B1[11] => U[20]) = (0:0:0, 0:0:0);
    (B2B1[11] => U[21]) = (0:0:0, 0:0:0);
    (B2B1[11] => U[22]) = (0:0:0, 0:0:0);
    (B2B1[11] => U[23]) = (0:0:0, 0:0:0);
    (B2B1[11] => U[24]) = (0:0:0, 0:0:0);
    (B2B1[11] => U[25]) = (0:0:0, 0:0:0);
    (B2B1[11] => U[26]) = (0:0:0, 0:0:0);
    (B2B1[11] => U[27]) = (0:0:0, 0:0:0);
    (B2B1[11] => U[28]) = (0:0:0, 0:0:0);
    (B2B1[11] => U[29]) = (0:0:0, 0:0:0);
    (B2B1[11] => U[30]) = (0:0:0, 0:0:0);
    (B2B1[11] => U[31]) = (0:0:0, 0:0:0);
    (B2B1[11] => U[32]) = (0:0:0, 0:0:0);
    (B2B1[11] => U[33]) = (0:0:0, 0:0:0);
    (B2B1[11] => U[34]) = (0:0:0, 0:0:0);
    (B2B1[11] => U[35]) = (0:0:0, 0:0:0);
    (B2B1[11] => U[36]) = (0:0:0, 0:0:0);
    (B2B1[11] => U[37]) = (0:0:0, 0:0:0);
    (B2B1[11] => U[38]) = (0:0:0, 0:0:0);
    (B2B1[11] => U[39]) = (0:0:0, 0:0:0);
    (B2B1[11] => U[40]) = (0:0:0, 0:0:0);
    (B2B1[11] => U[41]) = (0:0:0, 0:0:0);
    (B2B1[11] => V[10]) = (0:0:0, 0:0:0);
    (B2B1[11] => V[11]) = (0:0:0, 0:0:0);
    (B2B1[11] => V[12]) = (0:0:0, 0:0:0);
    (B2B1[11] => V[13]) = (0:0:0, 0:0:0);
    (B2B1[11] => V[14]) = (0:0:0, 0:0:0);
    (B2B1[11] => V[15]) = (0:0:0, 0:0:0);
    (B2B1[11] => V[16]) = (0:0:0, 0:0:0);
    (B2B1[11] => V[17]) = (0:0:0, 0:0:0);
    (B2B1[11] => V[18]) = (0:0:0, 0:0:0);
    (B2B1[11] => V[19]) = (0:0:0, 0:0:0);
    (B2B1[11] => V[20]) = (0:0:0, 0:0:0);
    (B2B1[11] => V[21]) = (0:0:0, 0:0:0);
    (B2B1[11] => V[22]) = (0:0:0, 0:0:0);
    (B2B1[11] => V[23]) = (0:0:0, 0:0:0);
    (B2B1[11] => V[24]) = (0:0:0, 0:0:0);
    (B2B1[11] => V[25]) = (0:0:0, 0:0:0);
    (B2B1[11] => V[26]) = (0:0:0, 0:0:0);
    (B2B1[11] => V[27]) = (0:0:0, 0:0:0);
    (B2B1[11] => V[28]) = (0:0:0, 0:0:0);
    (B2B1[11] => V[29]) = (0:0:0, 0:0:0);
    (B2B1[11] => V[30]) = (0:0:0, 0:0:0);
    (B2B1[11] => V[31]) = (0:0:0, 0:0:0);
    (B2B1[11] => V[32]) = (0:0:0, 0:0:0);
    (B2B1[11] => V[33]) = (0:0:0, 0:0:0);
    (B2B1[11] => V[34]) = (0:0:0, 0:0:0);
    (B2B1[11] => V[35]) = (0:0:0, 0:0:0);
    (B2B1[11] => V[36]) = (0:0:0, 0:0:0);
    (B2B1[11] => V[37]) = (0:0:0, 0:0:0);
    (B2B1[11] => V[38]) = (0:0:0, 0:0:0);
    (B2B1[11] => V[39]) = (0:0:0, 0:0:0);
    (B2B1[11] => V[40]) = (0:0:0, 0:0:0);
    (B2B1[12] => U[13]) = (0:0:0, 0:0:0);
    (B2B1[12] => U[14]) = (0:0:0, 0:0:0);
    (B2B1[12] => U[15]) = (0:0:0, 0:0:0);
    (B2B1[12] => U[16]) = (0:0:0, 0:0:0);
    (B2B1[12] => U[17]) = (0:0:0, 0:0:0);
    (B2B1[12] => U[18]) = (0:0:0, 0:0:0);
    (B2B1[12] => U[19]) = (0:0:0, 0:0:0);
    (B2B1[12] => U[20]) = (0:0:0, 0:0:0);
    (B2B1[12] => U[21]) = (0:0:0, 0:0:0);
    (B2B1[12] => U[22]) = (0:0:0, 0:0:0);
    (B2B1[12] => U[23]) = (0:0:0, 0:0:0);
    (B2B1[12] => U[24]) = (0:0:0, 0:0:0);
    (B2B1[12] => U[25]) = (0:0:0, 0:0:0);
    (B2B1[12] => U[26]) = (0:0:0, 0:0:0);
    (B2B1[12] => U[27]) = (0:0:0, 0:0:0);
    (B2B1[12] => U[28]) = (0:0:0, 0:0:0);
    (B2B1[12] => U[29]) = (0:0:0, 0:0:0);
    (B2B1[12] => U[30]) = (0:0:0, 0:0:0);
    (B2B1[12] => U[31]) = (0:0:0, 0:0:0);
    (B2B1[12] => U[32]) = (0:0:0, 0:0:0);
    (B2B1[12] => U[33]) = (0:0:0, 0:0:0);
    (B2B1[12] => U[34]) = (0:0:0, 0:0:0);
    (B2B1[12] => U[35]) = (0:0:0, 0:0:0);
    (B2B1[12] => U[36]) = (0:0:0, 0:0:0);
    (B2B1[12] => U[37]) = (0:0:0, 0:0:0);
    (B2B1[12] => U[38]) = (0:0:0, 0:0:0);
    (B2B1[12] => U[39]) = (0:0:0, 0:0:0);
    (B2B1[12] => U[40]) = (0:0:0, 0:0:0);
    (B2B1[12] => U[41]) = (0:0:0, 0:0:0);
    (B2B1[12] => V[12]) = (0:0:0, 0:0:0);
    (B2B1[12] => V[13]) = (0:0:0, 0:0:0);
    (B2B1[12] => V[14]) = (0:0:0, 0:0:0);
    (B2B1[12] => V[15]) = (0:0:0, 0:0:0);
    (B2B1[12] => V[16]) = (0:0:0, 0:0:0);
    (B2B1[12] => V[17]) = (0:0:0, 0:0:0);
    (B2B1[12] => V[18]) = (0:0:0, 0:0:0);
    (B2B1[12] => V[19]) = (0:0:0, 0:0:0);
    (B2B1[12] => V[20]) = (0:0:0, 0:0:0);
    (B2B1[12] => V[21]) = (0:0:0, 0:0:0);
    (B2B1[12] => V[22]) = (0:0:0, 0:0:0);
    (B2B1[12] => V[23]) = (0:0:0, 0:0:0);
    (B2B1[12] => V[24]) = (0:0:0, 0:0:0);
    (B2B1[12] => V[25]) = (0:0:0, 0:0:0);
    (B2B1[12] => V[26]) = (0:0:0, 0:0:0);
    (B2B1[12] => V[27]) = (0:0:0, 0:0:0);
    (B2B1[12] => V[28]) = (0:0:0, 0:0:0);
    (B2B1[12] => V[29]) = (0:0:0, 0:0:0);
    (B2B1[12] => V[30]) = (0:0:0, 0:0:0);
    (B2B1[12] => V[31]) = (0:0:0, 0:0:0);
    (B2B1[12] => V[32]) = (0:0:0, 0:0:0);
    (B2B1[12] => V[33]) = (0:0:0, 0:0:0);
    (B2B1[12] => V[34]) = (0:0:0, 0:0:0);
    (B2B1[12] => V[35]) = (0:0:0, 0:0:0);
    (B2B1[12] => V[36]) = (0:0:0, 0:0:0);
    (B2B1[12] => V[37]) = (0:0:0, 0:0:0);
    (B2B1[12] => V[38]) = (0:0:0, 0:0:0);
    (B2B1[12] => V[39]) = (0:0:0, 0:0:0);
    (B2B1[12] => V[40]) = (0:0:0, 0:0:0);
    (B2B1[13] => U[13]) = (0:0:0, 0:0:0);
    (B2B1[13] => U[14]) = (0:0:0, 0:0:0);
    (B2B1[13] => U[15]) = (0:0:0, 0:0:0);
    (B2B1[13] => U[16]) = (0:0:0, 0:0:0);
    (B2B1[13] => U[17]) = (0:0:0, 0:0:0);
    (B2B1[13] => U[18]) = (0:0:0, 0:0:0);
    (B2B1[13] => U[19]) = (0:0:0, 0:0:0);
    (B2B1[13] => U[20]) = (0:0:0, 0:0:0);
    (B2B1[13] => U[21]) = (0:0:0, 0:0:0);
    (B2B1[13] => U[22]) = (0:0:0, 0:0:0);
    (B2B1[13] => U[23]) = (0:0:0, 0:0:0);
    (B2B1[13] => U[24]) = (0:0:0, 0:0:0);
    (B2B1[13] => U[25]) = (0:0:0, 0:0:0);
    (B2B1[13] => U[26]) = (0:0:0, 0:0:0);
    (B2B1[13] => U[27]) = (0:0:0, 0:0:0);
    (B2B1[13] => U[28]) = (0:0:0, 0:0:0);
    (B2B1[13] => U[29]) = (0:0:0, 0:0:0);
    (B2B1[13] => U[30]) = (0:0:0, 0:0:0);
    (B2B1[13] => U[31]) = (0:0:0, 0:0:0);
    (B2B1[13] => U[32]) = (0:0:0, 0:0:0);
    (B2B1[13] => U[33]) = (0:0:0, 0:0:0);
    (B2B1[13] => U[34]) = (0:0:0, 0:0:0);
    (B2B1[13] => U[35]) = (0:0:0, 0:0:0);
    (B2B1[13] => U[36]) = (0:0:0, 0:0:0);
    (B2B1[13] => U[37]) = (0:0:0, 0:0:0);
    (B2B1[13] => U[38]) = (0:0:0, 0:0:0);
    (B2B1[13] => U[39]) = (0:0:0, 0:0:0);
    (B2B1[13] => U[40]) = (0:0:0, 0:0:0);
    (B2B1[13] => U[41]) = (0:0:0, 0:0:0);
    (B2B1[13] => U[42]) = (0:0:0, 0:0:0);
    (B2B1[13] => V[12]) = (0:0:0, 0:0:0);
    (B2B1[13] => V[13]) = (0:0:0, 0:0:0);
    (B2B1[13] => V[14]) = (0:0:0, 0:0:0);
    (B2B1[13] => V[15]) = (0:0:0, 0:0:0);
    (B2B1[13] => V[16]) = (0:0:0, 0:0:0);
    (B2B1[13] => V[17]) = (0:0:0, 0:0:0);
    (B2B1[13] => V[18]) = (0:0:0, 0:0:0);
    (B2B1[13] => V[19]) = (0:0:0, 0:0:0);
    (B2B1[13] => V[20]) = (0:0:0, 0:0:0);
    (B2B1[13] => V[21]) = (0:0:0, 0:0:0);
    (B2B1[13] => V[22]) = (0:0:0, 0:0:0);
    (B2B1[13] => V[23]) = (0:0:0, 0:0:0);
    (B2B1[13] => V[24]) = (0:0:0, 0:0:0);
    (B2B1[13] => V[25]) = (0:0:0, 0:0:0);
    (B2B1[13] => V[26]) = (0:0:0, 0:0:0);
    (B2B1[13] => V[27]) = (0:0:0, 0:0:0);
    (B2B1[13] => V[28]) = (0:0:0, 0:0:0);
    (B2B1[13] => V[29]) = (0:0:0, 0:0:0);
    (B2B1[13] => V[30]) = (0:0:0, 0:0:0);
    (B2B1[13] => V[31]) = (0:0:0, 0:0:0);
    (B2B1[13] => V[32]) = (0:0:0, 0:0:0);
    (B2B1[13] => V[33]) = (0:0:0, 0:0:0);
    (B2B1[13] => V[34]) = (0:0:0, 0:0:0);
    (B2B1[13] => V[35]) = (0:0:0, 0:0:0);
    (B2B1[13] => V[36]) = (0:0:0, 0:0:0);
    (B2B1[13] => V[37]) = (0:0:0, 0:0:0);
    (B2B1[13] => V[38]) = (0:0:0, 0:0:0);
    (B2B1[13] => V[39]) = (0:0:0, 0:0:0);
    (B2B1[13] => V[40]) = (0:0:0, 0:0:0);
    (B2B1[13] => V[41]) = (0:0:0, 0:0:0);
    (B2B1[14] => U[15]) = (0:0:0, 0:0:0);
    (B2B1[14] => U[16]) = (0:0:0, 0:0:0);
    (B2B1[14] => U[17]) = (0:0:0, 0:0:0);
    (B2B1[14] => U[18]) = (0:0:0, 0:0:0);
    (B2B1[14] => U[19]) = (0:0:0, 0:0:0);
    (B2B1[14] => U[20]) = (0:0:0, 0:0:0);
    (B2B1[14] => U[21]) = (0:0:0, 0:0:0);
    (B2B1[14] => U[22]) = (0:0:0, 0:0:0);
    (B2B1[14] => U[23]) = (0:0:0, 0:0:0);
    (B2B1[14] => U[24]) = (0:0:0, 0:0:0);
    (B2B1[14] => U[25]) = (0:0:0, 0:0:0);
    (B2B1[14] => U[26]) = (0:0:0, 0:0:0);
    (B2B1[14] => U[27]) = (0:0:0, 0:0:0);
    (B2B1[14] => U[28]) = (0:0:0, 0:0:0);
    (B2B1[14] => U[29]) = (0:0:0, 0:0:0);
    (B2B1[14] => U[30]) = (0:0:0, 0:0:0);
    (B2B1[14] => U[31]) = (0:0:0, 0:0:0);
    (B2B1[14] => U[32]) = (0:0:0, 0:0:0);
    (B2B1[14] => U[33]) = (0:0:0, 0:0:0);
    (B2B1[14] => U[34]) = (0:0:0, 0:0:0);
    (B2B1[14] => U[35]) = (0:0:0, 0:0:0);
    (B2B1[14] => U[36]) = (0:0:0, 0:0:0);
    (B2B1[14] => U[37]) = (0:0:0, 0:0:0);
    (B2B1[14] => U[38]) = (0:0:0, 0:0:0);
    (B2B1[14] => U[39]) = (0:0:0, 0:0:0);
    (B2B1[14] => U[40]) = (0:0:0, 0:0:0);
    (B2B1[14] => U[41]) = (0:0:0, 0:0:0);
    (B2B1[14] => U[42]) = (0:0:0, 0:0:0);
    (B2B1[14] => V[14]) = (0:0:0, 0:0:0);
    (B2B1[14] => V[15]) = (0:0:0, 0:0:0);
    (B2B1[14] => V[16]) = (0:0:0, 0:0:0);
    (B2B1[14] => V[17]) = (0:0:0, 0:0:0);
    (B2B1[14] => V[18]) = (0:0:0, 0:0:0);
    (B2B1[14] => V[19]) = (0:0:0, 0:0:0);
    (B2B1[14] => V[20]) = (0:0:0, 0:0:0);
    (B2B1[14] => V[21]) = (0:0:0, 0:0:0);
    (B2B1[14] => V[22]) = (0:0:0, 0:0:0);
    (B2B1[14] => V[23]) = (0:0:0, 0:0:0);
    (B2B1[14] => V[24]) = (0:0:0, 0:0:0);
    (B2B1[14] => V[25]) = (0:0:0, 0:0:0);
    (B2B1[14] => V[26]) = (0:0:0, 0:0:0);
    (B2B1[14] => V[27]) = (0:0:0, 0:0:0);
    (B2B1[14] => V[28]) = (0:0:0, 0:0:0);
    (B2B1[14] => V[29]) = (0:0:0, 0:0:0);
    (B2B1[14] => V[30]) = (0:0:0, 0:0:0);
    (B2B1[14] => V[31]) = (0:0:0, 0:0:0);
    (B2B1[14] => V[32]) = (0:0:0, 0:0:0);
    (B2B1[14] => V[33]) = (0:0:0, 0:0:0);
    (B2B1[14] => V[34]) = (0:0:0, 0:0:0);
    (B2B1[14] => V[35]) = (0:0:0, 0:0:0);
    (B2B1[14] => V[36]) = (0:0:0, 0:0:0);
    (B2B1[14] => V[37]) = (0:0:0, 0:0:0);
    (B2B1[14] => V[38]) = (0:0:0, 0:0:0);
    (B2B1[14] => V[39]) = (0:0:0, 0:0:0);
    (B2B1[14] => V[40]) = (0:0:0, 0:0:0);
    (B2B1[14] => V[41]) = (0:0:0, 0:0:0);
    (B2B1[15] => U[15]) = (0:0:0, 0:0:0);
    (B2B1[15] => U[16]) = (0:0:0, 0:0:0);
    (B2B1[15] => U[17]) = (0:0:0, 0:0:0);
    (B2B1[15] => U[18]) = (0:0:0, 0:0:0);
    (B2B1[15] => U[19]) = (0:0:0, 0:0:0);
    (B2B1[15] => U[20]) = (0:0:0, 0:0:0);
    (B2B1[15] => U[21]) = (0:0:0, 0:0:0);
    (B2B1[15] => U[22]) = (0:0:0, 0:0:0);
    (B2B1[15] => U[23]) = (0:0:0, 0:0:0);
    (B2B1[15] => U[24]) = (0:0:0, 0:0:0);
    (B2B1[15] => U[25]) = (0:0:0, 0:0:0);
    (B2B1[15] => U[26]) = (0:0:0, 0:0:0);
    (B2B1[15] => U[27]) = (0:0:0, 0:0:0);
    (B2B1[15] => U[28]) = (0:0:0, 0:0:0);
    (B2B1[15] => U[29]) = (0:0:0, 0:0:0);
    (B2B1[15] => U[30]) = (0:0:0, 0:0:0);
    (B2B1[15] => U[31]) = (0:0:0, 0:0:0);
    (B2B1[15] => U[32]) = (0:0:0, 0:0:0);
    (B2B1[15] => U[33]) = (0:0:0, 0:0:0);
    (B2B1[15] => U[34]) = (0:0:0, 0:0:0);
    (B2B1[15] => U[35]) = (0:0:0, 0:0:0);
    (B2B1[15] => U[36]) = (0:0:0, 0:0:0);
    (B2B1[15] => U[37]) = (0:0:0, 0:0:0);
    (B2B1[15] => U[38]) = (0:0:0, 0:0:0);
    (B2B1[15] => U[39]) = (0:0:0, 0:0:0);
    (B2B1[15] => U[40]) = (0:0:0, 0:0:0);
    (B2B1[15] => U[41]) = (0:0:0, 0:0:0);
    (B2B1[15] => U[42]) = (0:0:0, 0:0:0);
    (B2B1[15] => U[43]) = (0:0:0, 0:0:0);
    (B2B1[15] => V[14]) = (0:0:0, 0:0:0);
    (B2B1[15] => V[15]) = (0:0:0, 0:0:0);
    (B2B1[15] => V[16]) = (0:0:0, 0:0:0);
    (B2B1[15] => V[17]) = (0:0:0, 0:0:0);
    (B2B1[15] => V[18]) = (0:0:0, 0:0:0);
    (B2B1[15] => V[19]) = (0:0:0, 0:0:0);
    (B2B1[15] => V[20]) = (0:0:0, 0:0:0);
    (B2B1[15] => V[21]) = (0:0:0, 0:0:0);
    (B2B1[15] => V[22]) = (0:0:0, 0:0:0);
    (B2B1[15] => V[23]) = (0:0:0, 0:0:0);
    (B2B1[15] => V[24]) = (0:0:0, 0:0:0);
    (B2B1[15] => V[25]) = (0:0:0, 0:0:0);
    (B2B1[15] => V[26]) = (0:0:0, 0:0:0);
    (B2B1[15] => V[27]) = (0:0:0, 0:0:0);
    (B2B1[15] => V[28]) = (0:0:0, 0:0:0);
    (B2B1[15] => V[29]) = (0:0:0, 0:0:0);
    (B2B1[15] => V[30]) = (0:0:0, 0:0:0);
    (B2B1[15] => V[31]) = (0:0:0, 0:0:0);
    (B2B1[15] => V[32]) = (0:0:0, 0:0:0);
    (B2B1[15] => V[33]) = (0:0:0, 0:0:0);
    (B2B1[15] => V[34]) = (0:0:0, 0:0:0);
    (B2B1[15] => V[35]) = (0:0:0, 0:0:0);
    (B2B1[15] => V[36]) = (0:0:0, 0:0:0);
    (B2B1[15] => V[37]) = (0:0:0, 0:0:0);
    (B2B1[15] => V[38]) = (0:0:0, 0:0:0);
    (B2B1[15] => V[39]) = (0:0:0, 0:0:0);
    (B2B1[15] => V[40]) = (0:0:0, 0:0:0);
    (B2B1[15] => V[41]) = (0:0:0, 0:0:0);
    (B2B1[15] => V[42]) = (0:0:0, 0:0:0);
    (B2B1[15] => V[43]) = (0:0:0, 0:0:0);
    (B2B1[16] => U[17]) = (0:0:0, 0:0:0);
    (B2B1[16] => U[18]) = (0:0:0, 0:0:0);
    (B2B1[16] => U[19]) = (0:0:0, 0:0:0);
    (B2B1[16] => U[20]) = (0:0:0, 0:0:0);
    (B2B1[16] => U[21]) = (0:0:0, 0:0:0);
    (B2B1[16] => U[22]) = (0:0:0, 0:0:0);
    (B2B1[16] => U[23]) = (0:0:0, 0:0:0);
    (B2B1[16] => U[24]) = (0:0:0, 0:0:0);
    (B2B1[16] => U[25]) = (0:0:0, 0:0:0);
    (B2B1[16] => U[26]) = (0:0:0, 0:0:0);
    (B2B1[16] => U[27]) = (0:0:0, 0:0:0);
    (B2B1[16] => U[28]) = (0:0:0, 0:0:0);
    (B2B1[16] => U[29]) = (0:0:0, 0:0:0);
    (B2B1[16] => U[30]) = (0:0:0, 0:0:0);
    (B2B1[16] => U[31]) = (0:0:0, 0:0:0);
    (B2B1[16] => U[32]) = (0:0:0, 0:0:0);
    (B2B1[16] => U[33]) = (0:0:0, 0:0:0);
    (B2B1[16] => U[34]) = (0:0:0, 0:0:0);
    (B2B1[16] => U[35]) = (0:0:0, 0:0:0);
    (B2B1[16] => U[36]) = (0:0:0, 0:0:0);
    (B2B1[16] => U[37]) = (0:0:0, 0:0:0);
    (B2B1[16] => U[38]) = (0:0:0, 0:0:0);
    (B2B1[16] => U[39]) = (0:0:0, 0:0:0);
    (B2B1[16] => U[40]) = (0:0:0, 0:0:0);
    (B2B1[16] => U[41]) = (0:0:0, 0:0:0);
    (B2B1[16] => U[42]) = (0:0:0, 0:0:0);
    (B2B1[16] => U[43]) = (0:0:0, 0:0:0);
    (B2B1[16] => V[16]) = (0:0:0, 0:0:0);
    (B2B1[16] => V[17]) = (0:0:0, 0:0:0);
    (B2B1[16] => V[18]) = (0:0:0, 0:0:0);
    (B2B1[16] => V[19]) = (0:0:0, 0:0:0);
    (B2B1[16] => V[20]) = (0:0:0, 0:0:0);
    (B2B1[16] => V[21]) = (0:0:0, 0:0:0);
    (B2B1[16] => V[22]) = (0:0:0, 0:0:0);
    (B2B1[16] => V[23]) = (0:0:0, 0:0:0);
    (B2B1[16] => V[24]) = (0:0:0, 0:0:0);
    (B2B1[16] => V[25]) = (0:0:0, 0:0:0);
    (B2B1[16] => V[26]) = (0:0:0, 0:0:0);
    (B2B1[16] => V[27]) = (0:0:0, 0:0:0);
    (B2B1[16] => V[28]) = (0:0:0, 0:0:0);
    (B2B1[16] => V[29]) = (0:0:0, 0:0:0);
    (B2B1[16] => V[30]) = (0:0:0, 0:0:0);
    (B2B1[16] => V[31]) = (0:0:0, 0:0:0);
    (B2B1[16] => V[32]) = (0:0:0, 0:0:0);
    (B2B1[16] => V[33]) = (0:0:0, 0:0:0);
    (B2B1[16] => V[34]) = (0:0:0, 0:0:0);
    (B2B1[16] => V[35]) = (0:0:0, 0:0:0);
    (B2B1[16] => V[36]) = (0:0:0, 0:0:0);
    (B2B1[16] => V[37]) = (0:0:0, 0:0:0);
    (B2B1[16] => V[38]) = (0:0:0, 0:0:0);
    (B2B1[16] => V[39]) = (0:0:0, 0:0:0);
    (B2B1[16] => V[40]) = (0:0:0, 0:0:0);
    (B2B1[16] => V[41]) = (0:0:0, 0:0:0);
    (B2B1[16] => V[42]) = (0:0:0, 0:0:0);
    (B2B1[16] => V[43]) = (0:0:0, 0:0:0);
    (B2B1[17] => BMULT17) = (0:0:0, 0:0:0);
    (B2B1[17] => U[17]) = (0:0:0, 0:0:0);
    (B2B1[17] => U[18]) = (0:0:0, 0:0:0);
    (B2B1[17] => U[19]) = (0:0:0, 0:0:0);
    (B2B1[17] => U[20]) = (0:0:0, 0:0:0);
    (B2B1[17] => U[21]) = (0:0:0, 0:0:0);
    (B2B1[17] => U[22]) = (0:0:0, 0:0:0);
    (B2B1[17] => U[23]) = (0:0:0, 0:0:0);
    (B2B1[17] => U[24]) = (0:0:0, 0:0:0);
    (B2B1[17] => U[25]) = (0:0:0, 0:0:0);
    (B2B1[17] => U[26]) = (0:0:0, 0:0:0);
    (B2B1[17] => U[27]) = (0:0:0, 0:0:0);
    (B2B1[17] => U[28]) = (0:0:0, 0:0:0);
    (B2B1[17] => U[29]) = (0:0:0, 0:0:0);
    (B2B1[17] => U[30]) = (0:0:0, 0:0:0);
    (B2B1[17] => U[31]) = (0:0:0, 0:0:0);
    (B2B1[17] => U[32]) = (0:0:0, 0:0:0);
    (B2B1[17] => U[33]) = (0:0:0, 0:0:0);
    (B2B1[17] => U[34]) = (0:0:0, 0:0:0);
    (B2B1[17] => U[35]) = (0:0:0, 0:0:0);
    (B2B1[17] => U[36]) = (0:0:0, 0:0:0);
    (B2B1[17] => U[37]) = (0:0:0, 0:0:0);
    (B2B1[17] => U[38]) = (0:0:0, 0:0:0);
    (B2B1[17] => U[39]) = (0:0:0, 0:0:0);
    (B2B1[17] => U[40]) = (0:0:0, 0:0:0);
    (B2B1[17] => U[41]) = (0:0:0, 0:0:0);
    (B2B1[17] => U[42]) = (0:0:0, 0:0:0);
    (B2B1[17] => U[43]) = (0:0:0, 0:0:0);
    (B2B1[17] => V[16]) = (0:0:0, 0:0:0);
    (B2B1[17] => V[17]) = (0:0:0, 0:0:0);
    (B2B1[17] => V[18]) = (0:0:0, 0:0:0);
    (B2B1[17] => V[19]) = (0:0:0, 0:0:0);
    (B2B1[17] => V[20]) = (0:0:0, 0:0:0);
    (B2B1[17] => V[21]) = (0:0:0, 0:0:0);
    (B2B1[17] => V[22]) = (0:0:0, 0:0:0);
    (B2B1[17] => V[23]) = (0:0:0, 0:0:0);
    (B2B1[17] => V[24]) = (0:0:0, 0:0:0);
    (B2B1[17] => V[25]) = (0:0:0, 0:0:0);
    (B2B1[17] => V[26]) = (0:0:0, 0:0:0);
    (B2B1[17] => V[27]) = (0:0:0, 0:0:0);
    (B2B1[17] => V[28]) = (0:0:0, 0:0:0);
    (B2B1[17] => V[29]) = (0:0:0, 0:0:0);
    (B2B1[17] => V[30]) = (0:0:0, 0:0:0);
    (B2B1[17] => V[31]) = (0:0:0, 0:0:0);
    (B2B1[17] => V[32]) = (0:0:0, 0:0:0);
    (B2B1[17] => V[33]) = (0:0:0, 0:0:0);
    (B2B1[17] => V[34]) = (0:0:0, 0:0:0);
    (B2B1[17] => V[35]) = (0:0:0, 0:0:0);
    (B2B1[17] => V[36]) = (0:0:0, 0:0:0);
    (B2B1[17] => V[37]) = (0:0:0, 0:0:0);
    (B2B1[17] => V[38]) = (0:0:0, 0:0:0);
    (B2B1[17] => V[39]) = (0:0:0, 0:0:0);
    (B2B1[17] => V[40]) = (0:0:0, 0:0:0);
    (B2B1[17] => V[41]) = (0:0:0, 0:0:0);
    (B2B1[17] => V[42]) = (0:0:0, 0:0:0);
    (B2B1[17] => V[43]) = (0:0:0, 0:0:0);
    (B2B1[1] => U[0]) = (0:0:0, 0:0:0);
    (B2B1[1] => U[10]) = (0:0:0, 0:0:0);
    (B2B1[1] => U[11]) = (0:0:0, 0:0:0);
    (B2B1[1] => U[12]) = (0:0:0, 0:0:0);
    (B2B1[1] => U[13]) = (0:0:0, 0:0:0);
    (B2B1[1] => U[14]) = (0:0:0, 0:0:0);
    (B2B1[1] => U[15]) = (0:0:0, 0:0:0);
    (B2B1[1] => U[16]) = (0:0:0, 0:0:0);
    (B2B1[1] => U[17]) = (0:0:0, 0:0:0);
    (B2B1[1] => U[18]) = (0:0:0, 0:0:0);
    (B2B1[1] => U[19]) = (0:0:0, 0:0:0);
    (B2B1[1] => U[1]) = (0:0:0, 0:0:0);
    (B2B1[1] => U[20]) = (0:0:0, 0:0:0);
    (B2B1[1] => U[21]) = (0:0:0, 0:0:0);
    (B2B1[1] => U[22]) = (0:0:0, 0:0:0);
    (B2B1[1] => U[23]) = (0:0:0, 0:0:0);
    (B2B1[1] => U[24]) = (0:0:0, 0:0:0);
    (B2B1[1] => U[25]) = (0:0:0, 0:0:0);
    (B2B1[1] => U[26]) = (0:0:0, 0:0:0);
    (B2B1[1] => U[27]) = (0:0:0, 0:0:0);
    (B2B1[1] => U[28]) = (0:0:0, 0:0:0);
    (B2B1[1] => U[29]) = (0:0:0, 0:0:0);
    (B2B1[1] => U[2]) = (0:0:0, 0:0:0);
    (B2B1[1] => U[30]) = (0:0:0, 0:0:0);
    (B2B1[1] => U[31]) = (0:0:0, 0:0:0);
    (B2B1[1] => U[32]) = (0:0:0, 0:0:0);
    (B2B1[1] => U[33]) = (0:0:0, 0:0:0);
    (B2B1[1] => U[3]) = (0:0:0, 0:0:0);
    (B2B1[1] => U[4]) = (0:0:0, 0:0:0);
    (B2B1[1] => U[5]) = (0:0:0, 0:0:0);
    (B2B1[1] => U[6]) = (0:0:0, 0:0:0);
    (B2B1[1] => U[7]) = (0:0:0, 0:0:0);
    (B2B1[1] => U[8]) = (0:0:0, 0:0:0);
    (B2B1[1] => U[9]) = (0:0:0, 0:0:0);
    (B2B1[1] => V[0]) = (0:0:0, 0:0:0);
    (B2B1[1] => V[10]) = (0:0:0, 0:0:0);
    (B2B1[1] => V[11]) = (0:0:0, 0:0:0);
    (B2B1[1] => V[12]) = (0:0:0, 0:0:0);
    (B2B1[1] => V[13]) = (0:0:0, 0:0:0);
    (B2B1[1] => V[14]) = (0:0:0, 0:0:0);
    (B2B1[1] => V[15]) = (0:0:0, 0:0:0);
    (B2B1[1] => V[16]) = (0:0:0, 0:0:0);
    (B2B1[1] => V[17]) = (0:0:0, 0:0:0);
    (B2B1[1] => V[18]) = (0:0:0, 0:0:0);
    (B2B1[1] => V[19]) = (0:0:0, 0:0:0);
    (B2B1[1] => V[20]) = (0:0:0, 0:0:0);
    (B2B1[1] => V[21]) = (0:0:0, 0:0:0);
    (B2B1[1] => V[22]) = (0:0:0, 0:0:0);
    (B2B1[1] => V[23]) = (0:0:0, 0:0:0);
    (B2B1[1] => V[24]) = (0:0:0, 0:0:0);
    (B2B1[1] => V[25]) = (0:0:0, 0:0:0);
    (B2B1[1] => V[26]) = (0:0:0, 0:0:0);
    (B2B1[1] => V[27]) = (0:0:0, 0:0:0);
    (B2B1[1] => V[28]) = (0:0:0, 0:0:0);
    (B2B1[1] => V[29]) = (0:0:0, 0:0:0);
    (B2B1[1] => V[30]) = (0:0:0, 0:0:0);
    (B2B1[1] => V[31]) = (0:0:0, 0:0:0);
    (B2B1[1] => V[32]) = (0:0:0, 0:0:0);
    (B2B1[1] => V[4]) = (0:0:0, 0:0:0);
    (B2B1[1] => V[5]) = (0:0:0, 0:0:0);
    (B2B1[1] => V[6]) = (0:0:0, 0:0:0);
    (B2B1[1] => V[7]) = (0:0:0, 0:0:0);
    (B2B1[1] => V[8]) = (0:0:0, 0:0:0);
    (B2B1[1] => V[9]) = (0:0:0, 0:0:0);
    (B2B1[2] => U[10]) = (0:0:0, 0:0:0);
    (B2B1[2] => U[11]) = (0:0:0, 0:0:0);
    (B2B1[2] => U[12]) = (0:0:0, 0:0:0);
    (B2B1[2] => U[13]) = (0:0:0, 0:0:0);
    (B2B1[2] => U[14]) = (0:0:0, 0:0:0);
    (B2B1[2] => U[15]) = (0:0:0, 0:0:0);
    (B2B1[2] => U[16]) = (0:0:0, 0:0:0);
    (B2B1[2] => U[17]) = (0:0:0, 0:0:0);
    (B2B1[2] => U[18]) = (0:0:0, 0:0:0);
    (B2B1[2] => U[19]) = (0:0:0, 0:0:0);
    (B2B1[2] => U[20]) = (0:0:0, 0:0:0);
    (B2B1[2] => U[21]) = (0:0:0, 0:0:0);
    (B2B1[2] => U[22]) = (0:0:0, 0:0:0);
    (B2B1[2] => U[23]) = (0:0:0, 0:0:0);
    (B2B1[2] => U[24]) = (0:0:0, 0:0:0);
    (B2B1[2] => U[25]) = (0:0:0, 0:0:0);
    (B2B1[2] => U[26]) = (0:0:0, 0:0:0);
    (B2B1[2] => U[27]) = (0:0:0, 0:0:0);
    (B2B1[2] => U[28]) = (0:0:0, 0:0:0);
    (B2B1[2] => U[29]) = (0:0:0, 0:0:0);
    (B2B1[2] => U[2]) = (0:0:0, 0:0:0);
    (B2B1[2] => U[30]) = (0:0:0, 0:0:0);
    (B2B1[2] => U[31]) = (0:0:0, 0:0:0);
    (B2B1[2] => U[32]) = (0:0:0, 0:0:0);
    (B2B1[2] => U[33]) = (0:0:0, 0:0:0);
    (B2B1[2] => U[3]) = (0:0:0, 0:0:0);
    (B2B1[2] => U[4]) = (0:0:0, 0:0:0);
    (B2B1[2] => U[5]) = (0:0:0, 0:0:0);
    (B2B1[2] => U[6]) = (0:0:0, 0:0:0);
    (B2B1[2] => U[7]) = (0:0:0, 0:0:0);
    (B2B1[2] => U[8]) = (0:0:0, 0:0:0);
    (B2B1[2] => U[9]) = (0:0:0, 0:0:0);
    (B2B1[2] => V[10]) = (0:0:0, 0:0:0);
    (B2B1[2] => V[11]) = (0:0:0, 0:0:0);
    (B2B1[2] => V[12]) = (0:0:0, 0:0:0);
    (B2B1[2] => V[13]) = (0:0:0, 0:0:0);
    (B2B1[2] => V[14]) = (0:0:0, 0:0:0);
    (B2B1[2] => V[15]) = (0:0:0, 0:0:0);
    (B2B1[2] => V[16]) = (0:0:0, 0:0:0);
    (B2B1[2] => V[17]) = (0:0:0, 0:0:0);
    (B2B1[2] => V[18]) = (0:0:0, 0:0:0);
    (B2B1[2] => V[19]) = (0:0:0, 0:0:0);
    (B2B1[2] => V[20]) = (0:0:0, 0:0:0);
    (B2B1[2] => V[21]) = (0:0:0, 0:0:0);
    (B2B1[2] => V[22]) = (0:0:0, 0:0:0);
    (B2B1[2] => V[23]) = (0:0:0, 0:0:0);
    (B2B1[2] => V[24]) = (0:0:0, 0:0:0);
    (B2B1[2] => V[25]) = (0:0:0, 0:0:0);
    (B2B1[2] => V[26]) = (0:0:0, 0:0:0);
    (B2B1[2] => V[27]) = (0:0:0, 0:0:0);
    (B2B1[2] => V[28]) = (0:0:0, 0:0:0);
    (B2B1[2] => V[29]) = (0:0:0, 0:0:0);
    (B2B1[2] => V[30]) = (0:0:0, 0:0:0);
    (B2B1[2] => V[31]) = (0:0:0, 0:0:0);
    (B2B1[2] => V[32]) = (0:0:0, 0:0:0);
    (B2B1[2] => V[4]) = (0:0:0, 0:0:0);
    (B2B1[2] => V[5]) = (0:0:0, 0:0:0);
    (B2B1[2] => V[6]) = (0:0:0, 0:0:0);
    (B2B1[2] => V[7]) = (0:0:0, 0:0:0);
    (B2B1[2] => V[8]) = (0:0:0, 0:0:0);
    (B2B1[2] => V[9]) = (0:0:0, 0:0:0);
    (B2B1[3] => U[10]) = (0:0:0, 0:0:0);
    (B2B1[3] => U[11]) = (0:0:0, 0:0:0);
    (B2B1[3] => U[12]) = (0:0:0, 0:0:0);
    (B2B1[3] => U[13]) = (0:0:0, 0:0:0);
    (B2B1[3] => U[14]) = (0:0:0, 0:0:0);
    (B2B1[3] => U[15]) = (0:0:0, 0:0:0);
    (B2B1[3] => U[16]) = (0:0:0, 0:0:0);
    (B2B1[3] => U[17]) = (0:0:0, 0:0:0);
    (B2B1[3] => U[18]) = (0:0:0, 0:0:0);
    (B2B1[3] => U[19]) = (0:0:0, 0:0:0);
    (B2B1[3] => U[20]) = (0:0:0, 0:0:0);
    (B2B1[3] => U[21]) = (0:0:0, 0:0:0);
    (B2B1[3] => U[22]) = (0:0:0, 0:0:0);
    (B2B1[3] => U[23]) = (0:0:0, 0:0:0);
    (B2B1[3] => U[24]) = (0:0:0, 0:0:0);
    (B2B1[3] => U[25]) = (0:0:0, 0:0:0);
    (B2B1[3] => U[26]) = (0:0:0, 0:0:0);
    (B2B1[3] => U[27]) = (0:0:0, 0:0:0);
    (B2B1[3] => U[28]) = (0:0:0, 0:0:0);
    (B2B1[3] => U[29]) = (0:0:0, 0:0:0);
    (B2B1[3] => U[2]) = (0:0:0, 0:0:0);
    (B2B1[3] => U[30]) = (0:0:0, 0:0:0);
    (B2B1[3] => U[31]) = (0:0:0, 0:0:0);
    (B2B1[3] => U[32]) = (0:0:0, 0:0:0);
    (B2B1[3] => U[33]) = (0:0:0, 0:0:0);
    (B2B1[3] => U[34]) = (0:0:0, 0:0:0);
    (B2B1[3] => U[35]) = (0:0:0, 0:0:0);
    (B2B1[3] => U[3]) = (0:0:0, 0:0:0);
    (B2B1[3] => U[4]) = (0:0:0, 0:0:0);
    (B2B1[3] => U[5]) = (0:0:0, 0:0:0);
    (B2B1[3] => U[6]) = (0:0:0, 0:0:0);
    (B2B1[3] => U[7]) = (0:0:0, 0:0:0);
    (B2B1[3] => U[8]) = (0:0:0, 0:0:0);
    (B2B1[3] => U[9]) = (0:0:0, 0:0:0);
    (B2B1[3] => V[10]) = (0:0:0, 0:0:0);
    (B2B1[3] => V[11]) = (0:0:0, 0:0:0);
    (B2B1[3] => V[12]) = (0:0:0, 0:0:0);
    (B2B1[3] => V[13]) = (0:0:0, 0:0:0);
    (B2B1[3] => V[14]) = (0:0:0, 0:0:0);
    (B2B1[3] => V[15]) = (0:0:0, 0:0:0);
    (B2B1[3] => V[16]) = (0:0:0, 0:0:0);
    (B2B1[3] => V[17]) = (0:0:0, 0:0:0);
    (B2B1[3] => V[18]) = (0:0:0, 0:0:0);
    (B2B1[3] => V[19]) = (0:0:0, 0:0:0);
    (B2B1[3] => V[20]) = (0:0:0, 0:0:0);
    (B2B1[3] => V[21]) = (0:0:0, 0:0:0);
    (B2B1[3] => V[22]) = (0:0:0, 0:0:0);
    (B2B1[3] => V[23]) = (0:0:0, 0:0:0);
    (B2B1[3] => V[24]) = (0:0:0, 0:0:0);
    (B2B1[3] => V[25]) = (0:0:0, 0:0:0);
    (B2B1[3] => V[26]) = (0:0:0, 0:0:0);
    (B2B1[3] => V[27]) = (0:0:0, 0:0:0);
    (B2B1[3] => V[28]) = (0:0:0, 0:0:0);
    (B2B1[3] => V[29]) = (0:0:0, 0:0:0);
    (B2B1[3] => V[30]) = (0:0:0, 0:0:0);
    (B2B1[3] => V[31]) = (0:0:0, 0:0:0);
    (B2B1[3] => V[32]) = (0:0:0, 0:0:0);
    (B2B1[3] => V[33]) = (0:0:0, 0:0:0);
    (B2B1[3] => V[34]) = (0:0:0, 0:0:0);
    (B2B1[3] => V[4]) = (0:0:0, 0:0:0);
    (B2B1[3] => V[5]) = (0:0:0, 0:0:0);
    (B2B1[3] => V[6]) = (0:0:0, 0:0:0);
    (B2B1[3] => V[7]) = (0:0:0, 0:0:0);
    (B2B1[3] => V[8]) = (0:0:0, 0:0:0);
    (B2B1[3] => V[9]) = (0:0:0, 0:0:0);
    (B2B1[4] => U[10]) = (0:0:0, 0:0:0);
    (B2B1[4] => U[11]) = (0:0:0, 0:0:0);
    (B2B1[4] => U[12]) = (0:0:0, 0:0:0);
    (B2B1[4] => U[13]) = (0:0:0, 0:0:0);
    (B2B1[4] => U[14]) = (0:0:0, 0:0:0);
    (B2B1[4] => U[15]) = (0:0:0, 0:0:0);
    (B2B1[4] => U[16]) = (0:0:0, 0:0:0);
    (B2B1[4] => U[17]) = (0:0:0, 0:0:0);
    (B2B1[4] => U[18]) = (0:0:0, 0:0:0);
    (B2B1[4] => U[19]) = (0:0:0, 0:0:0);
    (B2B1[4] => U[20]) = (0:0:0, 0:0:0);
    (B2B1[4] => U[21]) = (0:0:0, 0:0:0);
    (B2B1[4] => U[22]) = (0:0:0, 0:0:0);
    (B2B1[4] => U[23]) = (0:0:0, 0:0:0);
    (B2B1[4] => U[24]) = (0:0:0, 0:0:0);
    (B2B1[4] => U[25]) = (0:0:0, 0:0:0);
    (B2B1[4] => U[26]) = (0:0:0, 0:0:0);
    (B2B1[4] => U[27]) = (0:0:0, 0:0:0);
    (B2B1[4] => U[28]) = (0:0:0, 0:0:0);
    (B2B1[4] => U[29]) = (0:0:0, 0:0:0);
    (B2B1[4] => U[30]) = (0:0:0, 0:0:0);
    (B2B1[4] => U[31]) = (0:0:0, 0:0:0);
    (B2B1[4] => U[32]) = (0:0:0, 0:0:0);
    (B2B1[4] => U[33]) = (0:0:0, 0:0:0);
    (B2B1[4] => U[34]) = (0:0:0, 0:0:0);
    (B2B1[4] => U[35]) = (0:0:0, 0:0:0);
    (B2B1[4] => U[5]) = (0:0:0, 0:0:0);
    (B2B1[4] => U[6]) = (0:0:0, 0:0:0);
    (B2B1[4] => U[7]) = (0:0:0, 0:0:0);
    (B2B1[4] => U[8]) = (0:0:0, 0:0:0);
    (B2B1[4] => U[9]) = (0:0:0, 0:0:0);
    (B2B1[4] => V[10]) = (0:0:0, 0:0:0);
    (B2B1[4] => V[11]) = (0:0:0, 0:0:0);
    (B2B1[4] => V[12]) = (0:0:0, 0:0:0);
    (B2B1[4] => V[13]) = (0:0:0, 0:0:0);
    (B2B1[4] => V[14]) = (0:0:0, 0:0:0);
    (B2B1[4] => V[15]) = (0:0:0, 0:0:0);
    (B2B1[4] => V[16]) = (0:0:0, 0:0:0);
    (B2B1[4] => V[17]) = (0:0:0, 0:0:0);
    (B2B1[4] => V[18]) = (0:0:0, 0:0:0);
    (B2B1[4] => V[19]) = (0:0:0, 0:0:0);
    (B2B1[4] => V[20]) = (0:0:0, 0:0:0);
    (B2B1[4] => V[21]) = (0:0:0, 0:0:0);
    (B2B1[4] => V[22]) = (0:0:0, 0:0:0);
    (B2B1[4] => V[23]) = (0:0:0, 0:0:0);
    (B2B1[4] => V[24]) = (0:0:0, 0:0:0);
    (B2B1[4] => V[25]) = (0:0:0, 0:0:0);
    (B2B1[4] => V[26]) = (0:0:0, 0:0:0);
    (B2B1[4] => V[27]) = (0:0:0, 0:0:0);
    (B2B1[4] => V[28]) = (0:0:0, 0:0:0);
    (B2B1[4] => V[29]) = (0:0:0, 0:0:0);
    (B2B1[4] => V[30]) = (0:0:0, 0:0:0);
    (B2B1[4] => V[31]) = (0:0:0, 0:0:0);
    (B2B1[4] => V[32]) = (0:0:0, 0:0:0);
    (B2B1[4] => V[33]) = (0:0:0, 0:0:0);
    (B2B1[4] => V[34]) = (0:0:0, 0:0:0);
    (B2B1[4] => V[4]) = (0:0:0, 0:0:0);
    (B2B1[4] => V[5]) = (0:0:0, 0:0:0);
    (B2B1[4] => V[6]) = (0:0:0, 0:0:0);
    (B2B1[4] => V[7]) = (0:0:0, 0:0:0);
    (B2B1[4] => V[8]) = (0:0:0, 0:0:0);
    (B2B1[4] => V[9]) = (0:0:0, 0:0:0);
    (B2B1[5] => U[10]) = (0:0:0, 0:0:0);
    (B2B1[5] => U[11]) = (0:0:0, 0:0:0);
    (B2B1[5] => U[12]) = (0:0:0, 0:0:0);
    (B2B1[5] => U[13]) = (0:0:0, 0:0:0);
    (B2B1[5] => U[14]) = (0:0:0, 0:0:0);
    (B2B1[5] => U[15]) = (0:0:0, 0:0:0);
    (B2B1[5] => U[16]) = (0:0:0, 0:0:0);
    (B2B1[5] => U[17]) = (0:0:0, 0:0:0);
    (B2B1[5] => U[18]) = (0:0:0, 0:0:0);
    (B2B1[5] => U[19]) = (0:0:0, 0:0:0);
    (B2B1[5] => U[20]) = (0:0:0, 0:0:0);
    (B2B1[5] => U[21]) = (0:0:0, 0:0:0);
    (B2B1[5] => U[22]) = (0:0:0, 0:0:0);
    (B2B1[5] => U[23]) = (0:0:0, 0:0:0);
    (B2B1[5] => U[24]) = (0:0:0, 0:0:0);
    (B2B1[5] => U[25]) = (0:0:0, 0:0:0);
    (B2B1[5] => U[26]) = (0:0:0, 0:0:0);
    (B2B1[5] => U[27]) = (0:0:0, 0:0:0);
    (B2B1[5] => U[28]) = (0:0:0, 0:0:0);
    (B2B1[5] => U[29]) = (0:0:0, 0:0:0);
    (B2B1[5] => U[30]) = (0:0:0, 0:0:0);
    (B2B1[5] => U[31]) = (0:0:0, 0:0:0);
    (B2B1[5] => U[32]) = (0:0:0, 0:0:0);
    (B2B1[5] => U[33]) = (0:0:0, 0:0:0);
    (B2B1[5] => U[34]) = (0:0:0, 0:0:0);
    (B2B1[5] => U[35]) = (0:0:0, 0:0:0);
    (B2B1[5] => U[36]) = (0:0:0, 0:0:0);
    (B2B1[5] => U[5]) = (0:0:0, 0:0:0);
    (B2B1[5] => U[6]) = (0:0:0, 0:0:0);
    (B2B1[5] => U[7]) = (0:0:0, 0:0:0);
    (B2B1[5] => U[8]) = (0:0:0, 0:0:0);
    (B2B1[5] => U[9]) = (0:0:0, 0:0:0);
    (B2B1[5] => V[10]) = (0:0:0, 0:0:0);
    (B2B1[5] => V[11]) = (0:0:0, 0:0:0);
    (B2B1[5] => V[12]) = (0:0:0, 0:0:0);
    (B2B1[5] => V[13]) = (0:0:0, 0:0:0);
    (B2B1[5] => V[14]) = (0:0:0, 0:0:0);
    (B2B1[5] => V[15]) = (0:0:0, 0:0:0);
    (B2B1[5] => V[16]) = (0:0:0, 0:0:0);
    (B2B1[5] => V[17]) = (0:0:0, 0:0:0);
    (B2B1[5] => V[18]) = (0:0:0, 0:0:0);
    (B2B1[5] => V[19]) = (0:0:0, 0:0:0);
    (B2B1[5] => V[20]) = (0:0:0, 0:0:0);
    (B2B1[5] => V[21]) = (0:0:0, 0:0:0);
    (B2B1[5] => V[22]) = (0:0:0, 0:0:0);
    (B2B1[5] => V[23]) = (0:0:0, 0:0:0);
    (B2B1[5] => V[24]) = (0:0:0, 0:0:0);
    (B2B1[5] => V[25]) = (0:0:0, 0:0:0);
    (B2B1[5] => V[26]) = (0:0:0, 0:0:0);
    (B2B1[5] => V[27]) = (0:0:0, 0:0:0);
    (B2B1[5] => V[28]) = (0:0:0, 0:0:0);
    (B2B1[5] => V[29]) = (0:0:0, 0:0:0);
    (B2B1[5] => V[30]) = (0:0:0, 0:0:0);
    (B2B1[5] => V[31]) = (0:0:0, 0:0:0);
    (B2B1[5] => V[32]) = (0:0:0, 0:0:0);
    (B2B1[5] => V[33]) = (0:0:0, 0:0:0);
    (B2B1[5] => V[34]) = (0:0:0, 0:0:0);
    (B2B1[5] => V[35]) = (0:0:0, 0:0:0);
    (B2B1[5] => V[4]) = (0:0:0, 0:0:0);
    (B2B1[5] => V[5]) = (0:0:0, 0:0:0);
    (B2B1[5] => V[6]) = (0:0:0, 0:0:0);
    (B2B1[5] => V[7]) = (0:0:0, 0:0:0);
    (B2B1[5] => V[8]) = (0:0:0, 0:0:0);
    (B2B1[5] => V[9]) = (0:0:0, 0:0:0);
    (B2B1[6] => U[10]) = (0:0:0, 0:0:0);
    (B2B1[6] => U[11]) = (0:0:0, 0:0:0);
    (B2B1[6] => U[12]) = (0:0:0, 0:0:0);
    (B2B1[6] => U[13]) = (0:0:0, 0:0:0);
    (B2B1[6] => U[14]) = (0:0:0, 0:0:0);
    (B2B1[6] => U[15]) = (0:0:0, 0:0:0);
    (B2B1[6] => U[16]) = (0:0:0, 0:0:0);
    (B2B1[6] => U[17]) = (0:0:0, 0:0:0);
    (B2B1[6] => U[18]) = (0:0:0, 0:0:0);
    (B2B1[6] => U[19]) = (0:0:0, 0:0:0);
    (B2B1[6] => U[20]) = (0:0:0, 0:0:0);
    (B2B1[6] => U[21]) = (0:0:0, 0:0:0);
    (B2B1[6] => U[22]) = (0:0:0, 0:0:0);
    (B2B1[6] => U[23]) = (0:0:0, 0:0:0);
    (B2B1[6] => U[24]) = (0:0:0, 0:0:0);
    (B2B1[6] => U[25]) = (0:0:0, 0:0:0);
    (B2B1[6] => U[26]) = (0:0:0, 0:0:0);
    (B2B1[6] => U[27]) = (0:0:0, 0:0:0);
    (B2B1[6] => U[28]) = (0:0:0, 0:0:0);
    (B2B1[6] => U[29]) = (0:0:0, 0:0:0);
    (B2B1[6] => U[30]) = (0:0:0, 0:0:0);
    (B2B1[6] => U[31]) = (0:0:0, 0:0:0);
    (B2B1[6] => U[32]) = (0:0:0, 0:0:0);
    (B2B1[6] => U[33]) = (0:0:0, 0:0:0);
    (B2B1[6] => U[34]) = (0:0:0, 0:0:0);
    (B2B1[6] => U[35]) = (0:0:0, 0:0:0);
    (B2B1[6] => U[36]) = (0:0:0, 0:0:0);
    (B2B1[6] => U[7]) = (0:0:0, 0:0:0);
    (B2B1[6] => U[8]) = (0:0:0, 0:0:0);
    (B2B1[6] => U[9]) = (0:0:0, 0:0:0);
    (B2B1[6] => V[10]) = (0:0:0, 0:0:0);
    (B2B1[6] => V[11]) = (0:0:0, 0:0:0);
    (B2B1[6] => V[12]) = (0:0:0, 0:0:0);
    (B2B1[6] => V[13]) = (0:0:0, 0:0:0);
    (B2B1[6] => V[14]) = (0:0:0, 0:0:0);
    (B2B1[6] => V[15]) = (0:0:0, 0:0:0);
    (B2B1[6] => V[16]) = (0:0:0, 0:0:0);
    (B2B1[6] => V[17]) = (0:0:0, 0:0:0);
    (B2B1[6] => V[18]) = (0:0:0, 0:0:0);
    (B2B1[6] => V[19]) = (0:0:0, 0:0:0);
    (B2B1[6] => V[20]) = (0:0:0, 0:0:0);
    (B2B1[6] => V[21]) = (0:0:0, 0:0:0);
    (B2B1[6] => V[22]) = (0:0:0, 0:0:0);
    (B2B1[6] => V[23]) = (0:0:0, 0:0:0);
    (B2B1[6] => V[24]) = (0:0:0, 0:0:0);
    (B2B1[6] => V[25]) = (0:0:0, 0:0:0);
    (B2B1[6] => V[26]) = (0:0:0, 0:0:0);
    (B2B1[6] => V[27]) = (0:0:0, 0:0:0);
    (B2B1[6] => V[28]) = (0:0:0, 0:0:0);
    (B2B1[6] => V[29]) = (0:0:0, 0:0:0);
    (B2B1[6] => V[30]) = (0:0:0, 0:0:0);
    (B2B1[6] => V[31]) = (0:0:0, 0:0:0);
    (B2B1[6] => V[32]) = (0:0:0, 0:0:0);
    (B2B1[6] => V[33]) = (0:0:0, 0:0:0);
    (B2B1[6] => V[34]) = (0:0:0, 0:0:0);
    (B2B1[6] => V[35]) = (0:0:0, 0:0:0);
    (B2B1[6] => V[6]) = (0:0:0, 0:0:0);
    (B2B1[6] => V[7]) = (0:0:0, 0:0:0);
    (B2B1[6] => V[8]) = (0:0:0, 0:0:0);
    (B2B1[6] => V[9]) = (0:0:0, 0:0:0);
    (B2B1[7] => U[10]) = (0:0:0, 0:0:0);
    (B2B1[7] => U[11]) = (0:0:0, 0:0:0);
    (B2B1[7] => U[12]) = (0:0:0, 0:0:0);
    (B2B1[7] => U[13]) = (0:0:0, 0:0:0);
    (B2B1[7] => U[14]) = (0:0:0, 0:0:0);
    (B2B1[7] => U[15]) = (0:0:0, 0:0:0);
    (B2B1[7] => U[16]) = (0:0:0, 0:0:0);
    (B2B1[7] => U[17]) = (0:0:0, 0:0:0);
    (B2B1[7] => U[18]) = (0:0:0, 0:0:0);
    (B2B1[7] => U[19]) = (0:0:0, 0:0:0);
    (B2B1[7] => U[20]) = (0:0:0, 0:0:0);
    (B2B1[7] => U[21]) = (0:0:0, 0:0:0);
    (B2B1[7] => U[22]) = (0:0:0, 0:0:0);
    (B2B1[7] => U[23]) = (0:0:0, 0:0:0);
    (B2B1[7] => U[24]) = (0:0:0, 0:0:0);
    (B2B1[7] => U[25]) = (0:0:0, 0:0:0);
    (B2B1[7] => U[26]) = (0:0:0, 0:0:0);
    (B2B1[7] => U[27]) = (0:0:0, 0:0:0);
    (B2B1[7] => U[28]) = (0:0:0, 0:0:0);
    (B2B1[7] => U[29]) = (0:0:0, 0:0:0);
    (B2B1[7] => U[30]) = (0:0:0, 0:0:0);
    (B2B1[7] => U[31]) = (0:0:0, 0:0:0);
    (B2B1[7] => U[32]) = (0:0:0, 0:0:0);
    (B2B1[7] => U[33]) = (0:0:0, 0:0:0);
    (B2B1[7] => U[34]) = (0:0:0, 0:0:0);
    (B2B1[7] => U[35]) = (0:0:0, 0:0:0);
    (B2B1[7] => U[36]) = (0:0:0, 0:0:0);
    (B2B1[7] => U[37]) = (0:0:0, 0:0:0);
    (B2B1[7] => U[38]) = (0:0:0, 0:0:0);
    (B2B1[7] => U[7]) = (0:0:0, 0:0:0);
    (B2B1[7] => U[8]) = (0:0:0, 0:0:0);
    (B2B1[7] => U[9]) = (0:0:0, 0:0:0);
    (B2B1[7] => V[10]) = (0:0:0, 0:0:0);
    (B2B1[7] => V[11]) = (0:0:0, 0:0:0);
    (B2B1[7] => V[12]) = (0:0:0, 0:0:0);
    (B2B1[7] => V[13]) = (0:0:0, 0:0:0);
    (B2B1[7] => V[14]) = (0:0:0, 0:0:0);
    (B2B1[7] => V[15]) = (0:0:0, 0:0:0);
    (B2B1[7] => V[16]) = (0:0:0, 0:0:0);
    (B2B1[7] => V[17]) = (0:0:0, 0:0:0);
    (B2B1[7] => V[18]) = (0:0:0, 0:0:0);
    (B2B1[7] => V[19]) = (0:0:0, 0:0:0);
    (B2B1[7] => V[20]) = (0:0:0, 0:0:0);
    (B2B1[7] => V[21]) = (0:0:0, 0:0:0);
    (B2B1[7] => V[22]) = (0:0:0, 0:0:0);
    (B2B1[7] => V[23]) = (0:0:0, 0:0:0);
    (B2B1[7] => V[24]) = (0:0:0, 0:0:0);
    (B2B1[7] => V[25]) = (0:0:0, 0:0:0);
    (B2B1[7] => V[26]) = (0:0:0, 0:0:0);
    (B2B1[7] => V[27]) = (0:0:0, 0:0:0);
    (B2B1[7] => V[28]) = (0:0:0, 0:0:0);
    (B2B1[7] => V[29]) = (0:0:0, 0:0:0);
    (B2B1[7] => V[30]) = (0:0:0, 0:0:0);
    (B2B1[7] => V[31]) = (0:0:0, 0:0:0);
    (B2B1[7] => V[32]) = (0:0:0, 0:0:0);
    (B2B1[7] => V[33]) = (0:0:0, 0:0:0);
    (B2B1[7] => V[34]) = (0:0:0, 0:0:0);
    (B2B1[7] => V[35]) = (0:0:0, 0:0:0);
    (B2B1[7] => V[36]) = (0:0:0, 0:0:0);
    (B2B1[7] => V[37]) = (0:0:0, 0:0:0);
    (B2B1[7] => V[6]) = (0:0:0, 0:0:0);
    (B2B1[7] => V[7]) = (0:0:0, 0:0:0);
    (B2B1[7] => V[8]) = (0:0:0, 0:0:0);
    (B2B1[7] => V[9]) = (0:0:0, 0:0:0);
    (B2B1[8] => U[10]) = (0:0:0, 0:0:0);
    (B2B1[8] => U[11]) = (0:0:0, 0:0:0);
    (B2B1[8] => U[12]) = (0:0:0, 0:0:0);
    (B2B1[8] => U[13]) = (0:0:0, 0:0:0);
    (B2B1[8] => U[14]) = (0:0:0, 0:0:0);
    (B2B1[8] => U[15]) = (0:0:0, 0:0:0);
    (B2B1[8] => U[16]) = (0:0:0, 0:0:0);
    (B2B1[8] => U[17]) = (0:0:0, 0:0:0);
    (B2B1[8] => U[18]) = (0:0:0, 0:0:0);
    (B2B1[8] => U[19]) = (0:0:0, 0:0:0);
    (B2B1[8] => U[20]) = (0:0:0, 0:0:0);
    (B2B1[8] => U[21]) = (0:0:0, 0:0:0);
    (B2B1[8] => U[22]) = (0:0:0, 0:0:0);
    (B2B1[8] => U[23]) = (0:0:0, 0:0:0);
    (B2B1[8] => U[24]) = (0:0:0, 0:0:0);
    (B2B1[8] => U[25]) = (0:0:0, 0:0:0);
    (B2B1[8] => U[26]) = (0:0:0, 0:0:0);
    (B2B1[8] => U[27]) = (0:0:0, 0:0:0);
    (B2B1[8] => U[28]) = (0:0:0, 0:0:0);
    (B2B1[8] => U[29]) = (0:0:0, 0:0:0);
    (B2B1[8] => U[30]) = (0:0:0, 0:0:0);
    (B2B1[8] => U[31]) = (0:0:0, 0:0:0);
    (B2B1[8] => U[32]) = (0:0:0, 0:0:0);
    (B2B1[8] => U[33]) = (0:0:0, 0:0:0);
    (B2B1[8] => U[34]) = (0:0:0, 0:0:0);
    (B2B1[8] => U[35]) = (0:0:0, 0:0:0);
    (B2B1[8] => U[36]) = (0:0:0, 0:0:0);
    (B2B1[8] => U[37]) = (0:0:0, 0:0:0);
    (B2B1[8] => U[38]) = (0:0:0, 0:0:0);
    (B2B1[8] => U[9]) = (0:0:0, 0:0:0);
    (B2B1[8] => V[10]) = (0:0:0, 0:0:0);
    (B2B1[8] => V[11]) = (0:0:0, 0:0:0);
    (B2B1[8] => V[12]) = (0:0:0, 0:0:0);
    (B2B1[8] => V[13]) = (0:0:0, 0:0:0);
    (B2B1[8] => V[14]) = (0:0:0, 0:0:0);
    (B2B1[8] => V[15]) = (0:0:0, 0:0:0);
    (B2B1[8] => V[16]) = (0:0:0, 0:0:0);
    (B2B1[8] => V[17]) = (0:0:0, 0:0:0);
    (B2B1[8] => V[18]) = (0:0:0, 0:0:0);
    (B2B1[8] => V[19]) = (0:0:0, 0:0:0);
    (B2B1[8] => V[20]) = (0:0:0, 0:0:0);
    (B2B1[8] => V[21]) = (0:0:0, 0:0:0);
    (B2B1[8] => V[22]) = (0:0:0, 0:0:0);
    (B2B1[8] => V[23]) = (0:0:0, 0:0:0);
    (B2B1[8] => V[24]) = (0:0:0, 0:0:0);
    (B2B1[8] => V[25]) = (0:0:0, 0:0:0);
    (B2B1[8] => V[26]) = (0:0:0, 0:0:0);
    (B2B1[8] => V[27]) = (0:0:0, 0:0:0);
    (B2B1[8] => V[28]) = (0:0:0, 0:0:0);
    (B2B1[8] => V[29]) = (0:0:0, 0:0:0);
    (B2B1[8] => V[30]) = (0:0:0, 0:0:0);
    (B2B1[8] => V[31]) = (0:0:0, 0:0:0);
    (B2B1[8] => V[32]) = (0:0:0, 0:0:0);
    (B2B1[8] => V[33]) = (0:0:0, 0:0:0);
    (B2B1[8] => V[34]) = (0:0:0, 0:0:0);
    (B2B1[8] => V[35]) = (0:0:0, 0:0:0);
    (B2B1[8] => V[36]) = (0:0:0, 0:0:0);
    (B2B1[8] => V[37]) = (0:0:0, 0:0:0);
    (B2B1[8] => V[8]) = (0:0:0, 0:0:0);
    (B2B1[8] => V[9]) = (0:0:0, 0:0:0);
    (B2B1[9] => U[10]) = (0:0:0, 0:0:0);
    (B2B1[9] => U[11]) = (0:0:0, 0:0:0);
    (B2B1[9] => U[12]) = (0:0:0, 0:0:0);
    (B2B1[9] => U[13]) = (0:0:0, 0:0:0);
    (B2B1[9] => U[14]) = (0:0:0, 0:0:0);
    (B2B1[9] => U[15]) = (0:0:0, 0:0:0);
    (B2B1[9] => U[16]) = (0:0:0, 0:0:0);
    (B2B1[9] => U[17]) = (0:0:0, 0:0:0);
    (B2B1[9] => U[18]) = (0:0:0, 0:0:0);
    (B2B1[9] => U[19]) = (0:0:0, 0:0:0);
    (B2B1[9] => U[20]) = (0:0:0, 0:0:0);
    (B2B1[9] => U[21]) = (0:0:0, 0:0:0);
    (B2B1[9] => U[22]) = (0:0:0, 0:0:0);
    (B2B1[9] => U[23]) = (0:0:0, 0:0:0);
    (B2B1[9] => U[24]) = (0:0:0, 0:0:0);
    (B2B1[9] => U[25]) = (0:0:0, 0:0:0);
    (B2B1[9] => U[26]) = (0:0:0, 0:0:0);
    (B2B1[9] => U[27]) = (0:0:0, 0:0:0);
    (B2B1[9] => U[28]) = (0:0:0, 0:0:0);
    (B2B1[9] => U[29]) = (0:0:0, 0:0:0);
    (B2B1[9] => U[30]) = (0:0:0, 0:0:0);
    (B2B1[9] => U[31]) = (0:0:0, 0:0:0);
    (B2B1[9] => U[32]) = (0:0:0, 0:0:0);
    (B2B1[9] => U[33]) = (0:0:0, 0:0:0);
    (B2B1[9] => U[34]) = (0:0:0, 0:0:0);
    (B2B1[9] => U[35]) = (0:0:0, 0:0:0);
    (B2B1[9] => U[36]) = (0:0:0, 0:0:0);
    (B2B1[9] => U[37]) = (0:0:0, 0:0:0);
    (B2B1[9] => U[38]) = (0:0:0, 0:0:0);
    (B2B1[9] => U[39]) = (0:0:0, 0:0:0);
    (B2B1[9] => U[40]) = (0:0:0, 0:0:0);
    (B2B1[9] => U[9]) = (0:0:0, 0:0:0);
    (B2B1[9] => V[10]) = (0:0:0, 0:0:0);
    (B2B1[9] => V[11]) = (0:0:0, 0:0:0);
    (B2B1[9] => V[12]) = (0:0:0, 0:0:0);
    (B2B1[9] => V[13]) = (0:0:0, 0:0:0);
    (B2B1[9] => V[14]) = (0:0:0, 0:0:0);
    (B2B1[9] => V[15]) = (0:0:0, 0:0:0);
    (B2B1[9] => V[16]) = (0:0:0, 0:0:0);
    (B2B1[9] => V[17]) = (0:0:0, 0:0:0);
    (B2B1[9] => V[18]) = (0:0:0, 0:0:0);
    (B2B1[9] => V[19]) = (0:0:0, 0:0:0);
    (B2B1[9] => V[20]) = (0:0:0, 0:0:0);
    (B2B1[9] => V[21]) = (0:0:0, 0:0:0);
    (B2B1[9] => V[22]) = (0:0:0, 0:0:0);
    (B2B1[9] => V[23]) = (0:0:0, 0:0:0);
    (B2B1[9] => V[24]) = (0:0:0, 0:0:0);
    (B2B1[9] => V[25]) = (0:0:0, 0:0:0);
    (B2B1[9] => V[26]) = (0:0:0, 0:0:0);
    (B2B1[9] => V[27]) = (0:0:0, 0:0:0);
    (B2B1[9] => V[28]) = (0:0:0, 0:0:0);
    (B2B1[9] => V[29]) = (0:0:0, 0:0:0);
    (B2B1[9] => V[30]) = (0:0:0, 0:0:0);
    (B2B1[9] => V[31]) = (0:0:0, 0:0:0);
    (B2B1[9] => V[32]) = (0:0:0, 0:0:0);
    (B2B1[9] => V[33]) = (0:0:0, 0:0:0);
    (B2B1[9] => V[34]) = (0:0:0, 0:0:0);
    (B2B1[9] => V[35]) = (0:0:0, 0:0:0);
    (B2B1[9] => V[36]) = (0:0:0, 0:0:0);
    (B2B1[9] => V[37]) = (0:0:0, 0:0:0);
    (B2B1[9] => V[38]) = (0:0:0, 0:0:0);
    (B2B1[9] => V[39]) = (0:0:0, 0:0:0);
    (B2B1[9] => V[8]) = (0:0:0, 0:0:0);
    (B2B1[9] => V[9]) = (0:0:0, 0:0:0);
    specparam PATHPULSE$ = 0;
  endspecify
`endif
`endif
endmodule