module  pcie_app_7x #(
  parameter C_DATA_WIDTH = 64,            // RX/TX interface data width
  // Do not override parameters below this line
  parameter KEEP_WIDTH = C_DATA_WIDTH / 8,              // TSTRB width
  parameter TCQ        = 1
)(
  input                         user_clk,
  input                         user_reset,
  input                         user_lnk_up,
  // Tx
  //input  [5:0]                  tx_buf_av,
  //input                         tx_cfg_req,
  //input                         tx_err_drop,
  output                        tx_cfg_gnt,
  input                         s_axis_tx_tready,
  output  [C_DATA_WIDTH-1:0]    s_axis_tx_tdata,
  output  [KEEP_WIDTH-1:0]      s_axis_tx_tkeep,
  output  [3:0]                 s_axis_tx_tuser,
  output                        s_axis_tx_tlast,
  output                        s_axis_tx_tvalid,
  // Rx
  output                        rx_np_ok,
  output                        rx_np_req,
  input  [C_DATA_WIDTH-1:0]     m_axis_rx_tdata,
  input  [KEEP_WIDTH-1:0]       m_axis_rx_tkeep,
  input                         m_axis_rx_tlast,
  input                         m_axis_rx_tvalid,
  output                        m_axis_rx_tready,
  input    [21:0]               m_axis_rx_tuser,
  // Flow Control
  //input  [11:0]                 fc_cpld,
  //input  [7:0]                  fc_cplh,
  //input  [11:0]                 fc_npd,
  //input  [7:0]                  fc_nph,
  //input  [11:0]                 fc_pd,
  //input  [7:0]                  fc_ph,
  output [2:0]                  fc_sel,
  // CFG
  output                        cfg_err_cor,
  output                        cfg_err_ur,
  output                        cfg_err_ecrc,
  output                        cfg_err_cpl_timeout,
  output                        cfg_err_cpl_unexpect,
  output                        cfg_err_cpl_abort,
  output                        cfg_err_atomic_egress_blocked,
  output                        cfg_err_internal_cor,
  output                        cfg_err_malformed,
  output                        cfg_err_mc_blocked,
  output                        cfg_err_poisoned,
  output                        cfg_err_norecovery,
  output                        cfg_err_acs,
  output                        cfg_err_internal_uncor,
  output                        cfg_pm_halt_aspm_l0s,
  output                        cfg_pm_halt_aspm_l1,
  output                        cfg_pm_force_state_en,
  output [1:0]                  cfg_pm_force_state,
  output                        cfg_err_posted,
  output                        cfg_err_locked,
  output [47:0]                 cfg_err_tlp_cpl_header,
//  input                         cfg_err_cpl_rdy,
  output                        cfg_interrupt,
//  input                         cfg_interrupt_rdy,
  output                        cfg_interrupt_assert,
  output [7:0]                  cfg_interrupt_di,
//  input  [7:0]                  cfg_interrupt_do,
//  input  [2:0]                  cfg_interrupt_mmenable,
//  input                         cfg_interrupt_msienable,
//  input                         cfg_interrupt_msixenable,
//  input                         cfg_interrupt_msixfm,
  output                        cfg_turnoff_ok,
  input                         cfg_to_turnoff,
  output                        cfg_trn_pending,
  output                        cfg_pm_wake,
  input   [7:0]                 cfg_bus_number,
  input   [4:0]                 cfg_device_number,
  input   [2:0]                 cfg_function_number,
//  input  [15:0]                 cfg_status,
//  input  [15:0]                 cfg_command,
//  input  [15:0]                 cfg_dstatus,
//  input  [15:0]                 cfg_dcommand,
//  input  [15:0]                 cfg_lstatus,
//  input  [15:0]                 cfg_lcommand,
//  input  [15:0]                 cfg_dcommand2,
//  input   [2:0]                 cfg_pcie_link_state,
  output                        cfg_interrupt_stat,
  output  [4:0]                 cfg_pciecap_interrupt_msgnum,
  output  [1:0]                 pl_directed_link_change,
//  input   [5:0]                 pl_ltssm_state,
  output  [1:0]                 pl_directed_link_width,
  output                        pl_directed_link_speed,
  output                        pl_directed_link_auton,
  output                        pl_upstream_prefer_deemph,
//  input   [1:0]                 pl_sel_lnk_width,
//  input                         pl_sel_lnk_rate,
//  input                         pl_link_gen2_cap,
//  input                         pl_link_partner_gen2_supported,
//  input   [2:0]                 pl_initial_link_width,
//  input                         pl_link_upcfg_cap,
//  input   [1:0]                 pl_lane_reversal_mode,
//  input                         pl_received_hot_rst,
  output [127:0]                cfg_err_aer_headerlog,
  output   [4:0]                cfg_aer_interrupt_msgnum,
//  input                         cfg_err_aer_headerlog_set,
//  input                         cfg_aer_ecrc_check_en,
//  input                         cfg_aer_ecrc_gen_en,
  output [31:0]                 cfg_mgmt_di,
  output  [3:0]                 cfg_mgmt_byte_en,
  output  [9:0]                 cfg_mgmt_dwaddr,
  output                        cfg_mgmt_wr_en,
  output                        cfg_mgmt_rd_en,
  output                        cfg_mgmt_wr_readonly,
  output [63:0]                 cfg_dsn
);
  // PCIe Block EP Tieoffs - Example PIO doesn't support the following inputs                                       //
  assign fc_sel = 3'b0;
  assign rx_np_ok = 1'b1;                          // Allow Reception of Non-posted Traffic
  assign rx_np_req = 1'b1;                         // Always request Non-posted Traffic if available
  assign s_axis_tx_tuser[0] = 1'b0;                // Unused for V6
  assign s_axis_tx_tuser[1] = 1'b0;                // Error forward packet
  assign s_axis_tx_tuser[2] = 1'b0;                // Stream packet
  assign tx_cfg_gnt = 1'b1;                        // Always allow transmission of Config traffic within block
  assign cfg_err_cor = 1'b0;                       // Never report Correctable Error
  assign cfg_err_ur = 1'b0;                        // Never report UR
  assign cfg_err_ecrc = 1'b0;                      // Never report ECRC Error
  assign cfg_err_cpl_timeout = 1'b0;               // Never report Completion Timeout
  assign cfg_err_cpl_abort = 1'b0;                 // Never report Completion Abort
  assign cfg_err_cpl_unexpect = 1'b0;              // Never report unexpected completion
  assign cfg_err_posted = 1'b0;                    // Never qualify cfg_err_* inputs
  assign cfg_err_locked = 1'b0;                    // Never qualify cfg_err_ur or cfg_err_cpl_abort
  assign cfg_pm_wake = 1'b0;                       // Never direct the core to send a PM_PME Message
  assign cfg_trn_pending = 1'b0;                   // Never set the transaction pending bit in the Device Status Register
  assign cfg_err_atomic_egress_blocked = 1'b0;     // Never report Atomic TLP blocked
  assign cfg_err_internal_cor = 1'b0;              // Never report internal error occurred
  assign cfg_err_malformed = 1'b0;                 // Never report malformed error
  assign cfg_err_mc_blocked = 1'b0;                // Never report multi-cast TLP blocked
  assign cfg_err_poisoned = 1'b0;                  // Never report poisoned TLP received
  assign cfg_err_norecovery = 1'b0;                // Never qualify cfg_err_poisoned or cfg_err_cpl_timeout
  assign cfg_err_acs = 1'b0;                       // Never report an ACS violation
  assign cfg_err_internal_uncor = 1'b0;            // Never report internal uncorrectable error
  assign cfg_pm_halt_aspm_l0s = 1'b0;              // Allow entry into L0s
  assign cfg_pm_halt_aspm_l1 = 1'b0;               // Allow entry into L1
  assign cfg_pm_force_state_en  = 1'b0;            // Do not qualify cfg_pm_force_state
  assign cfg_pm_force_state  = 2'b00;              // Do not move force core into specific PM state
  assign cfg_err_aer_headerlog = 128'h0;           // Zero out the AER Header Log
  assign cfg_aer_interrupt_msgnum = 5'b00000;      // Zero out the AER Root Error Status Register
  assign cfg_interrupt_stat = 1'b0;                // Never set the Interrupt Status bit
  assign cfg_pciecap_interrupt_msgnum = 5'b00000;  // Zero out Interrupt Message Number
  assign cfg_interrupt_assert = 1'b0;              // Always drive interrupt de-assert
  assign cfg_interrupt = 1'b0;                     // Never drive interrupt by qualifying cfg_interrupt_assert
  assign pl_directed_link_change = 2'b00;          // Never initiate link change
  assign pl_directed_link_width = 2'b00;          // Zero out directed link width
  assign pl_directed_link_speed = 1'b0;            // Zero out directed link speed
  assign pl_directed_link_auton = 1'b0;            // Zero out link autonomous input
  assign pl_upstream_prefer_deemph = 1'b1;         // Zero out preferred de-emphasis of upstream port
  assign cfg_interrupt_di = 8'b0;                  // Do not set interrupt fields
  assign cfg_err_tlp_cpl_header = 48'h0;           // Zero out the header information
  assign cfg_mgmt_di = 32'h0;                      // Zero out CFG MGMT input data bus
  assign cfg_mgmt_byte_en = 4'h0;                  // Zero out CFG MGMT byte enables
  assign cfg_mgmt_dwaddr = 10'h0;                  // Zero out CFG MGMT 10-bit address port
  assign cfg_mgmt_wr_en = 1'b0;                    // Do not write CFG space
  assign cfg_mgmt_rd_en = 1'b0;                    // Do not read CFG space
  assign cfg_mgmt_wr_readonly = 1'b0;              // Never treat RO bit as RW
  assign cfg_dsn = `DSN;  // Assign the input DSN
  // Programmable I/O Module                                                                                        //
  wire [15:0] cfg_completer_id      = { cfg_bus_number, cfg_device_number, cfg_function_number };
//  wire        cfg_bus_mstr_enable   = cfg_command[2];
  reg         s_axis_tx_tready_i ;
  always @(posedge user_clk)
  begin
   if (user_reset)
      s_axis_tx_tready_i <= #TCQ 1'b0;
   else
      s_axis_tx_tready_i <= #TCQ s_axis_tx_tready;
  end
  PIO  #(
    .C_DATA_WIDTH( C_DATA_WIDTH ),
    .KEEP_WIDTH( KEEP_WIDTH ),
    .TCQ( TCQ )
  ) PIO (
    .user_clk ( user_clk ),                         // I
    .user_reset ( user_reset ),                     // I
    .user_lnk_up ( user_lnk_up ),                   // I
    .s_axis_tx_tready ( s_axis_tx_tready_i ),         // I
    .s_axis_tx_tdata ( s_axis_tx_tdata ),           // O
    .s_axis_tx_tkeep ( s_axis_tx_tkeep ),           // O
    .s_axis_tx_tlast ( s_axis_tx_tlast ),           // O
    .s_axis_tx_tvalid ( s_axis_tx_tvalid ),         // O
    .tx_src_dsc ( s_axis_tx_tuser[3] ),             // O
    .m_axis_rx_tdata( m_axis_rx_tdata ),            // I
    .m_axis_rx_tkeep( m_axis_rx_tkeep ),            // I
    .m_axis_rx_tlast( m_axis_rx_tlast ),            // I
    .m_axis_rx_tvalid( m_axis_rx_tvalid ),          // I
    .m_axis_rx_tready( m_axis_rx_tready ),          // O
    .m_axis_rx_tuser ( m_axis_rx_tuser ),           // I
    .cfg_to_turnoff ( cfg_to_turnoff ),             // I
    .cfg_turnoff_ok ( cfg_turnoff_ok ),             // O
    .cfg_completer_id ( cfg_completer_id )          // I [15:0]
  );
endmodule