module circl_b(
        input  wire [6:0] in_addr,
        output reg  [6:0] out_word
       );
always @*
 case( in_addr )
  7'h01: out_word = 7'h0A;
  7'h02: out_word = 7'h12;
  7'h03: out_word = 7'h18;
  7'h04: out_word = 7'h1C;
  7'h05: out_word = 7'h20;
  7'h06: out_word = 7'h23;
  7'h07: out_word = 7'h26;
  7'h08: out_word = 7'h29;
  7'h09: out_word = 7'h2C;
  7'h0A: out_word = 7'h2E;
  7'h0B: out_word = 7'h30;
  7'h0C: out_word = 7'h33;
  7'h0D: out_word = 7'h35;
  7'h0E: out_word = 7'h37;
  7'h0F: out_word = 7'h38;
  7'h10: out_word = 7'h3A;
  7'h11: out_word = 7'h3C;
  7'h12: out_word = 7'h3E;
  7'h13: out_word = 7'h3F;
  7'h14: out_word = 7'h41;
  7'h15: out_word = 7'h42;
  7'h16: out_word = 7'h44;
  7'h17: out_word = 7'h45;
  7'h18: out_word = 7'h46;
  7'h19: out_word = 7'h48;
  7'h1A: out_word = 7'h49;
  7'h1B: out_word = 7'h4A;
  7'h1C: out_word = 7'h4C;
  7'h1D: out_word = 7'h4D;
  7'h1E: out_word = 7'h4E;
  7'h1F: out_word = 7'h4F;
  7'h20: out_word = 7'h50;
  7'h21: out_word = 7'h51;
  7'h22: out_word = 7'h52;
  7'h23: out_word = 7'h53;
  7'h24: out_word = 7'h54;
  7'h25: out_word = 7'h55;
  7'h26: out_word = 7'h56;
  7'h27: out_word = 7'h57;
  7'h28: out_word = 7'h58;
  7'h29: out_word = 7'h59;
  7'h2A: out_word = 7'h5A;
  7'h2B: out_word = 7'h5B;
  7'h2C: out_word = 7'h5C;
  7'h2D: out_word = 7'h5C;
//  7'h2E: out_word = 7'h5D;
//  7'h2F: out_word = 7'h5E;
//  7'h30: out_word = 7'h5F;
//  7'h31: out_word = 7'h5F;
//  7'h32: out_word = 7'h60;
//  7'h33: out_word = 7'h61;
//  7'h34: out_word = 7'h62;
//  7'h35: out_word = 7'h62;
//  7'h36: out_word = 7'h63;
//  7'h37: out_word = 7'h64;
//  7'h38: out_word = 7'h64;
//  7'h39: out_word = 7'h65;
//  7'h3A: out_word = 7'h66;
//  7'h3B: out_word = 7'h66;
//  7'h3C: out_word = 7'h67;
//  7'h3D: out_word = 7'h67;
//  7'h3E: out_word = 7'h68;
//  7'h3F: out_word = 7'h68;
//  7'h40: out_word = 7'h69;
//  7'h41: out_word = 7'h6A;
//  7'h42: out_word = 7'h6A;
//  7'h43: out_word = 7'h6B;
//  7'h44: out_word = 7'h6B;
//  7'h45: out_word = 7'h6C;
//  7'h46: out_word = 7'h6C;
//  7'h47: out_word = 7'h6C;
//  7'h48: out_word = 7'h6D;
//  7'h49: out_word = 7'h6D;
//  7'h4A: out_word = 7'h6E;
  7'h4B: out_word = 7'h6E;
  7'h4C: out_word = 7'h6F;
  7'h4D: out_word = 7'h6F;
  7'h4E: out_word = 7'h6F;
  7'h4F: out_word = 7'h70;
  7'h50: out_word = 7'h70;
  7'h51: out_word = 7'h70;
  7'h52: out_word = 7'h71;
  7'h53: out_word = 7'h71;
  7'h54: out_word = 7'h71;
  7'h55: out_word = 7'h72;
  7'h56: out_word = 7'h72;
  7'h57: out_word = 7'h72;
  7'h58: out_word = 7'h73;
  7'h59: out_word = 7'h73;
  7'h5A: out_word = 7'h73;
  7'h5B: out_word = 7'h73;
  7'h5C: out_word = 7'h74;
  7'h5D: out_word = 7'h74;
  7'h5E: out_word = 7'h74;
  7'h5F: out_word = 7'h74;
  7'h60: out_word = 7'h75;
  7'h61: out_word = 7'h75;
  7'h62: out_word = 7'h75;
  7'h63: out_word = 7'h75;
  7'h64: out_word = 7'h75;
  7'h65: out_word = 7'h75;
  7'h66: out_word = 7'h76;
  7'h67: out_word = 7'h76;
  7'h68: out_word = 7'h76;
  7'h69: out_word = 7'h76;
  7'h6A: out_word = 7'h76;
  7'h6B: out_word = 7'h76;
  7'h6C: out_word = 7'h76;
  7'h6D: out_word = 7'h76;
  7'h6E: out_word = 7'h77;
  7'h6F: out_word = 7'h77;
  7'h70: out_word = 7'h77;
  7'h71: out_word = 7'h77;
  7'h72: out_word = 7'h77;
  7'h73: out_word = 7'h77;
  7'h74: out_word = 7'h77;
  7'h75: out_word = 7'h77;
  7'h76: out_word = 7'h77;
  7'h77: out_word = 7'h77;
  7'h78: out_word = 7'h77;
 default out_word = 7'h00;
 endcase
endmodule