module outputs
  wire [63 : 0] word_fst;
  wire [4 : 0] word_snd;
  wire RDY_server_reset_request_put, RDY_server_reset_response_get, valid;
  // inlined wires
  wire [68 : 0] dw_result$wget;
  wire dw_valid$wget, dw_valid$whas;
  // register requestR
  reg [214 : 0] requestR;
  wire [214 : 0] requestR$D_IN;
  wire requestR$EN;
  // register resultR
  reg [69 : 0] resultR;
  reg [69 : 0] resultR$D_IN;
  wire resultR$EN;
  // register stateR
  reg [1 : 0] stateR;
  reg [1 : 0] stateR$D_IN;
  wire stateR$EN;
  // ports of submodule fpu
  reg [201 : 0] fpu$server_core_request_put;
  wire [69 : 0] fpu$server_core_response_get;
  wire fpu$EN_server_core_request_put,
       fpu$EN_server_core_response_get,
       fpu$EN_server_reset_request_put,
       fpu$EN_server_reset_response_get,
       fpu$RDY_server_core_request_put,
       fpu$RDY_server_core_response_get,
       fpu$RDY_server_reset_request_put,
       fpu$RDY_server_reset_response_get;
  // ports of submodule frmFpuF
  wire frmFpuF$CLR, frmFpuF$DEQ, frmFpuF$D_IN, frmFpuF$ENQ;
  // ports of submodule resetReqsF
  wire resetReqsF$CLR,
       resetReqsF$DEQ,
       resetReqsF$EMPTY_N,
       resetReqsF$ENQ,
       resetReqsF$FULL_N;
  // ports of submodule resetRspsF
  wire resetRspsF$CLR,
       resetRspsF$DEQ,
       resetRspsF$EMPTY_N,
       resetRspsF$ENQ,
       resetRspsF$FULL_N;
  // rule scheduling signals
  wire CAN_FIRE_RL_doFADD_D,
       CAN_FIRE_RL_doFADD_S,
       CAN_FIRE_RL_doFCLASS_D,
       CAN_FIRE_RL_doFCLASS_S,
       CAN_FIRE_RL_doFCVT_D_L,
       CAN_FIRE_RL_doFCVT_D_LU,
       CAN_FIRE_RL_doFCVT_D_S,
       CAN_FIRE_RL_doFCVT_D_W,
       CAN_FIRE_RL_doFCVT_D_WU,
       CAN_FIRE_RL_doFCVT_LU_D,
       CAN_FIRE_RL_doFCVT_LU_S,
       CAN_FIRE_RL_doFCVT_L_D,
       CAN_FIRE_RL_doFCVT_L_S,
       CAN_FIRE_RL_doFCVT_S_D,
       CAN_FIRE_RL_doFCVT_S_L,
       CAN_FIRE_RL_doFCVT_S_LU,
       CAN_FIRE_RL_doFCVT_S_W,
       CAN_FIRE_RL_doFCVT_S_WU,
       CAN_FIRE_RL_doFCVT_WU_D,
       CAN_FIRE_RL_doFCVT_WU_S,
       CAN_FIRE_RL_doFCVT_W_D,
       CAN_FIRE_RL_doFCVT_W_S,
       CAN_FIRE_RL_doFDIV_D,
       CAN_FIRE_RL_doFDIV_S,
       CAN_FIRE_RL_doFEQ_D,
       CAN_FIRE_RL_doFEQ_S,
       CAN_FIRE_RL_doFLE_D,
       CAN_FIRE_RL_doFLE_S,
       CAN_FIRE_RL_doFLT_D,
       CAN_FIRE_RL_doFLT_S,
       CAN_FIRE_RL_doFMADD_D,
       CAN_FIRE_RL_doFMADD_S,
       CAN_FIRE_RL_doFMAX_D,
       CAN_FIRE_RL_doFMAX_S,
       CAN_FIRE_RL_doFMIN_D,
       CAN_FIRE_RL_doFMIN_S,
       CAN_FIRE_RL_doFMSUB_D,
       CAN_FIRE_RL_doFMSUB_S,
       CAN_FIRE_RL_doFMUL_D,
       CAN_FIRE_RL_doFMUL_S,
       CAN_FIRE_RL_doFMV_D_X,
       CAN_FIRE_RL_doFMV_W_X,
       CAN_FIRE_RL_doFMV_X_D,
       CAN_FIRE_RL_doFMV_X_W,
       CAN_FIRE_RL_doFNMADD_D,
       CAN_FIRE_RL_doFNMADD_S,
       CAN_FIRE_RL_doFNMSUB_D,
       CAN_FIRE_RL_doFNMSUB_S,
       CAN_FIRE_RL_doFSGNJN_D,
       CAN_FIRE_RL_doFSGNJN_S,
       CAN_FIRE_RL_doFSGNJX_D,
       CAN_FIRE_RL_doFSGNJX_S,
       CAN_FIRE_RL_doFSGNJ_D,
       CAN_FIRE_RL_doFSGNJ_S,
       CAN_FIRE_RL_doFSQRT_D,
       CAN_FIRE_RL_doFSQRT_S,
       CAN_FIRE_RL_doFSUB_D,
       CAN_FIRE_RL_doFSUB_S,
       CAN_FIRE_RL_rl_drive_fpu_result,
       CAN_FIRE_RL_rl_get_fpu_result,
       CAN_FIRE_RL_rl_reset_begin,
       CAN_FIRE_RL_rl_reset_end,
       CAN_FIRE_req,
       CAN_FIRE_server_reset_request_put,
       CAN_FIRE_server_reset_response_get,
       WILL_FIRE_RL_doFADD_D,
       WILL_FIRE_RL_doFADD_S,
       WILL_FIRE_RL_doFCLASS_D,
       WILL_FIRE_RL_doFCLASS_S,
       WILL_FIRE_RL_doFCVT_D_L,
       WILL_FIRE_RL_doFCVT_D_LU,
       WILL_FIRE_RL_doFCVT_D_S,
       WILL_FIRE_RL_doFCVT_D_W,
       WILL_FIRE_RL_doFCVT_D_WU,
       WILL_FIRE_RL_doFCVT_LU_D,
       WILL_FIRE_RL_doFCVT_LU_S,
       WILL_FIRE_RL_doFCVT_L_D,
       WILL_FIRE_RL_doFCVT_L_S,
       WILL_FIRE_RL_doFCVT_S_D,
       WILL_FIRE_RL_doFCVT_S_L,
       WILL_FIRE_RL_doFCVT_S_LU,
       WILL_FIRE_RL_doFCVT_S_W,
       WILL_FIRE_RL_doFCVT_S_WU,
       WILL_FIRE_RL_doFCVT_WU_D,
       WILL_FIRE_RL_doFCVT_WU_S,
       WILL_FIRE_RL_doFCVT_W_D,
       WILL_FIRE_RL_doFCVT_W_S,
       WILL_FIRE_RL_doFDIV_D,
       WILL_FIRE_RL_doFDIV_S,
       WILL_FIRE_RL_doFEQ_D,
       WILL_FIRE_RL_doFEQ_S,
       WILL_FIRE_RL_doFLE_D,
       WILL_FIRE_RL_doFLE_S,
       WILL_FIRE_RL_doFLT_D,
       WILL_FIRE_RL_doFLT_S,
       WILL_FIRE_RL_doFMADD_D,
       WILL_FIRE_RL_doFMADD_S,
       WILL_FIRE_RL_doFMAX_D,
       WILL_FIRE_RL_doFMAX_S,
       WILL_FIRE_RL_doFMIN_D,
       WILL_FIRE_RL_doFMIN_S,
       WILL_FIRE_RL_doFMSUB_D,
       WILL_FIRE_RL_doFMSUB_S,
       WILL_FIRE_RL_doFMUL_D,
       WILL_FIRE_RL_doFMUL_S,
       WILL_FIRE_RL_doFMV_D_X,
       WILL_FIRE_RL_doFMV_W_X,
       WILL_FIRE_RL_doFMV_X_D,
       WILL_FIRE_RL_doFMV_X_W,
       WILL_FIRE_RL_doFNMADD_D,
       WILL_FIRE_RL_doFNMADD_S,
       WILL_FIRE_RL_doFNMSUB_D,
       WILL_FIRE_RL_doFNMSUB_S,
       WILL_FIRE_RL_doFSGNJN_D,
       WILL_FIRE_RL_doFSGNJN_S,
       WILL_FIRE_RL_doFSGNJX_D,
       WILL_FIRE_RL_doFSGNJX_S,
       WILL_FIRE_RL_doFSGNJ_D,
       WILL_FIRE_RL_doFSGNJ_S,
       WILL_FIRE_RL_doFSQRT_D,
       WILL_FIRE_RL_doFSQRT_S,
       WILL_FIRE_RL_doFSUB_D,
       WILL_FIRE_RL_doFSUB_S,
       WILL_FIRE_RL_rl_drive_fpu_result,
       WILL_FIRE_RL_rl_get_fpu_result,
       WILL_FIRE_RL_rl_reset_begin,
       WILL_FIRE_RL_rl_reset_end,
       WILL_FIRE_req,
       WILL_FIRE_server_reset_request_put,
       WILL_FIRE_server_reset_response_get;
  // inputs to muxes for submodule ports
  wire [214 : 0] MUX_requestR$write_1__VAL_2;
  wire [201 : 0] MUX_fpu$server_core_request_put_1__VAL_1,
		 MUX_fpu$server_core_request_put_1__VAL_10,
		 MUX_fpu$server_core_request_put_1__VAL_11,
		 MUX_fpu$server_core_request_put_1__VAL_12,
		 MUX_fpu$server_core_request_put_1__VAL_13,
		 MUX_fpu$server_core_request_put_1__VAL_14,
		 MUX_fpu$server_core_request_put_1__VAL_15,
		 MUX_fpu$server_core_request_put_1__VAL_16,
		 MUX_fpu$server_core_request_put_1__VAL_17,
		 MUX_fpu$server_core_request_put_1__VAL_18,
		 MUX_fpu$server_core_request_put_1__VAL_2,
		 MUX_fpu$server_core_request_put_1__VAL_3,
		 MUX_fpu$server_core_request_put_1__VAL_4,
		 MUX_fpu$server_core_request_put_1__VAL_5,
		 MUX_fpu$server_core_request_put_1__VAL_6,
		 MUX_fpu$server_core_request_put_1__VAL_7,
		 MUX_fpu$server_core_request_put_1__VAL_8,
		 MUX_fpu$server_core_request_put_1__VAL_9;
  wire [69 : 0] MUX_resultR$write_1__VAL_10,
		MUX_resultR$write_1__VAL_11,
		MUX_resultR$write_1__VAL_12,
		MUX_resultR$write_1__VAL_13,
		MUX_resultR$write_1__VAL_14,
		MUX_resultR$write_1__VAL_15,
		MUX_resultR$write_1__VAL_16,
		MUX_resultR$write_1__VAL_17,
		MUX_resultR$write_1__VAL_18,
		MUX_resultR$write_1__VAL_19,
		MUX_resultR$write_1__VAL_20,
		MUX_resultR$write_1__VAL_21,
		MUX_resultR$write_1__VAL_22,
		MUX_resultR$write_1__VAL_23,
		MUX_resultR$write_1__VAL_24,
		MUX_resultR$write_1__VAL_25,
		MUX_resultR$write_1__VAL_26,
		MUX_resultR$write_1__VAL_27,
		MUX_resultR$write_1__VAL_28,
		MUX_resultR$write_1__VAL_29,
		MUX_resultR$write_1__VAL_3,
		MUX_resultR$write_1__VAL_30,
		MUX_resultR$write_1__VAL_31,
		MUX_resultR$write_1__VAL_32,
		MUX_resultR$write_1__VAL_33,
		MUX_resultR$write_1__VAL_34,
		MUX_resultR$write_1__VAL_35,
		MUX_resultR$write_1__VAL_36,
		MUX_resultR$write_1__VAL_37,
		MUX_resultR$write_1__VAL_38,
		MUX_resultR$write_1__VAL_39,
		MUX_resultR$write_1__VAL_4,
		MUX_resultR$write_1__VAL_40,
		MUX_resultR$write_1__VAL_41,
		MUX_resultR$write_1__VAL_42,
		MUX_resultR$write_1__VAL_43,
		MUX_resultR$write_1__VAL_6,
		MUX_resultR$write_1__VAL_7,
		MUX_resultR$write_1__VAL_8,
		MUX_resultR$write_1__VAL_9;
  wire [68 : 0] MUX_dw_result$wset_1__VAL_1;
  wire MUX_dw_result$wset_1__SEL_1;
  // declarations used by system tasks
  // synopsys translate_off
  reg [31 : 0] v__h1224;
  reg [31 : 0] v__h1777;
  reg [31 : 0] v__h1966;
  reg [31 : 0] v__h2168;
  reg [31 : 0] v__h2418;
  reg [31 : 0] v__h2593;
  reg [31 : 0] v__h2768;
  reg [31 : 0] v__h2950;
  reg [31 : 0] v__h3139;
  reg [31 : 0] v__h3337;
  reg [31 : 0] v__h3520;
  reg [31 : 0] v__h3693;
  reg [31 : 0] v__h3882;
  reg [31 : 0] v__h16640;
  reg [31 : 0] v__h28741;
  reg [31 : 0] v__h35941;
  reg [31 : 0] v__h42829;
  reg [31 : 0] v__h44905;
  reg [31 : 0] v__h45689;
  reg [31 : 0] v__h47303;
  reg [31 : 0] v__h48090;
  reg [31 : 0] v__h50764;
  reg [31 : 0] v__h53335;
  reg [31 : 0] v__h53495;
  reg [31 : 0] v__h53671;
  reg [31 : 0] v__h55194;
  reg [31 : 0] v__h56303;
  reg [31 : 0] v__h57430;
  reg [31 : 0] v__h57911;
  reg [31 : 0] v__h58124;
  reg [31 : 0] v__h58311;
  reg [31 : 0] v__h58491;
  reg [31 : 0] v__h58676;
  reg [31 : 0] v__h58848;
  reg [31 : 0] v__h59020;
  reg [31 : 0] v__h59199;
  reg [31 : 0] v__h59386;
  reg [31 : 0] v__h59583;
  reg [31 : 0] v__h59744;
  reg [31 : 0] v__h59907;
  reg [31 : 0] v__h60075;
  reg [31 : 0] v__h71274;
  reg [31 : 0] v__h82193;
  reg [31 : 0] v__h83807;
  reg [31 : 0] v__h84594;
  reg [31 : 0] v__h97596;
  reg [31 : 0] v__h110093;
  reg [31 : 0] v__h112152;
  reg [31 : 0] v__h112936;
  reg [31 : 0] v__h167802;
  reg [31 : 0] v__h213792;
  reg [31 : 0] v__h218378;
  reg [31 : 0] v__h222864;
  reg [31 : 0] v__h225599;
  reg [31 : 0] v__h227516;
  reg [31 : 0] v__h229453;
  reg [31 : 0] v__h229605;
  reg [31 : 0] v__h229762;
  reg [31 : 0] v__h1218;
  reg [31 : 0] v__h1771;
  reg [31 : 0] v__h1960;
  reg [31 : 0] v__h2162;
  reg [31 : 0] v__h2412;
  reg [31 : 0] v__h2587;
  reg [31 : 0] v__h2762;
  reg [31 : 0] v__h2944;
  reg [31 : 0] v__h3133;
  reg [31 : 0] v__h3331;
  reg [31 : 0] v__h3514;
  reg [31 : 0] v__h3687;
  reg [31 : 0] v__h3876;
  reg [31 : 0] v__h16634;
  reg [31 : 0] v__h28735;
  reg [31 : 0] v__h35935;
  reg [31 : 0] v__h42823;
  reg [31 : 0] v__h44899;
  reg [31 : 0] v__h45683;
  reg [31 : 0] v__h47297;
  reg [31 : 0] v__h48084;
  reg [31 : 0] v__h50758;
  reg [31 : 0] v__h53329;
  reg [31 : 0] v__h53489;
  reg [31 : 0] v__h53665;
  reg [31 : 0] v__h55188;
  reg [31 : 0] v__h56297;
  reg [31 : 0] v__h57424;
  reg [31 : 0] v__h57905;
  reg [31 : 0] v__h58118;
  reg [31 : 0] v__h58305;
  reg [31 : 0] v__h58485;
  reg [31 : 0] v__h58670;
  reg [31 : 0] v__h58842;
  reg [31 : 0] v__h59014;
  reg [31 : 0] v__h59193;
  reg [31 : 0] v__h59380;
  reg [31 : 0] v__h59577;
  reg [31 : 0] v__h59738;
  reg [31 : 0] v__h59901;
  reg [31 : 0] v__h60069;
  reg [31 : 0] v__h71268;
  reg [31 : 0] v__h82187;
  reg [31 : 0] v__h83801;
  reg [31 : 0] v__h84588;
  reg [31 : 0] v__h97590;
  reg [31 : 0] v__h110087;
  reg [31 : 0] v__h112146;
  reg [31 : 0] v__h112930;
  reg [31 : 0] v__h167796;
  reg [31 : 0] v__h213786;
  reg [31 : 0] v__h218372;
  reg [31 : 0] v__h222858;
  reg [31 : 0] v__h225593;
  reg [31 : 0] v__h227510;
  reg [31 : 0] v__h229447;
  reg [31 : 0] v__h229599;
  reg [31 : 0] v__h229756;
  // synopsys translate_on
  // remaining internal signals
  reg [51 : 0] CASE_guard0129_0b0_sfd___39389_BITS_53_TO_2_0b_ETC__q78,
	       CASE_guard0129_0b0_sfd___39389_BITS_53_TO_2_0b_ETC__q79,
	       CASE_guard02175_0b0_theResult___snd11344_BITS__ETC__q175,
	       CASE_guard02175_0b0_theResult___snd11344_BITS__ETC__q176,
	       CASE_guard0346_0b0_sfd___30336_BITS_54_TO_3_0b_ETC__q93,
	       CASE_guard0346_0b0_sfd___30336_BITS_54_TO_3_0b_ETC__q94,
	       CASE_guard08246_0b0_sfd___37286_BITS_63_TO_12__ETC__q113,
	       CASE_guard08246_0b0_sfd___37286_BITS_63_TO_12__ETC__q114,
	       CASE_guard08975_0b0_sfd___37286_BITS_62_TO_11__ETC__q111,
	       CASE_guard08975_0b0_sfd___37286_BITS_62_TO_11__ETC__q112,
	       CASE_guard1075_0b0_sfd___30336_BITS_53_TO_2_0b_ETC__q91,
	       CASE_guard1075_0b0_sfd___30336_BITS_53_TO_2_0b_ETC__q92,
	       CASE_guard5721_0b0_sfd___35005_BITS_63_TO_12_0_ETC__q107,
	       CASE_guard5721_0b0_sfd___35005_BITS_63_TO_12_0_ETC__q108,
	       CASE_guard6451_0b0_sfd___35005_BITS_62_TO_11_0_ETC__q103,
	       CASE_guard6451_0b0_sfd___35005_BITS_62_TO_11_0_ETC__q104,
	       CASE_guard81312_0b0_theResult___snd90457_BITS__ETC__q171,
	       CASE_guard81312_0b0_theResult___snd90457_BITS__ETC__q172,
	       CASE_guard91853_0b0_sfdin01328_BITS_56_TO_5_0b_ETC__q173,
	       CASE_guard91853_0b0_sfdin01328_BITS_56_TO_5_0b_ETC__q174,
	       CASE_guard9399_0b0_sfd___39389_BITS_54_TO_3_0b_ETC__q82,
	       CASE_guard9399_0b0_sfd___39389_BITS_54_TO_3_0b_ETC__q83,
	       CASE_requestR_BITS_194_TO_192_0x1_450359962737_ETC__q7,
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2474,
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2492,
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2661,
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2676,
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d3013,
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d3031,
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d3170,
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d3185,
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d5100,
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d5127,
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d5146;
  reg [22 : 0] CASE_guard1384_0b0_sfd___31374_BITS_31_TO_9_0b_ETC__q64,
	       CASE_guard1384_0b0_sfd___31374_BITS_31_TO_9_0b_ETC__q65,
	       CASE_guard1910_0b0_sfd___31374_BITS_30_TO_8_0b_ETC__q62,
	       CASE_guard1910_0b0_sfd___31374_BITS_30_TO_8_0b_ETC__q63,
	       CASE_guard26038_0b0_sfdin35384_BITS_56_TO_34_0_ETC__q135,
	       CASE_guard26038_0b0_sfdin35384_BITS_56_TO_34_0_ETC__q136,
	       CASE_guard36028_0b0_theResult___snd45260_BITS__ETC__q137,
	       CASE_guard36028_0b0_theResult___snd45260_BITS__ETC__q138,
	       CASE_guard4468_0b0_sfd___34458_BITS_31_TO_9_0b_ETC__q51,
	       CASE_guard4468_0b0_sfd___34458_BITS_31_TO_9_0b_ETC__q52,
	       CASE_guard46250_0b0_sfdin55725_BITS_56_TO_34_0_ETC__q139,
	       CASE_guard46250_0b0_sfdin55725_BITS_56_TO_34_0_ETC__q140,
	       CASE_guard4995_0b0_sfd___34458_BITS_30_TO_8_0b_ETC__q53,
	       CASE_guard4995_0b0_sfd___34458_BITS_30_TO_8_0b_ETC__q54,
	       CASE_guard5015_0b0_sfd___35005_BITS_63_TO_41_0_ETC__q21,
	       CASE_guard5015_0b0_sfd___35005_BITS_63_TO_41_0_ETC__q22,
	       CASE_guard5545_0b0_sfd___35005_BITS_62_TO_40_0_ETC__q23,
	       CASE_guard5545_0b0_sfd___35005_BITS_62_TO_40_0_ETC__q24,
	       CASE_guard56369_0b0_theResult___snd65625_BITS__ETC__q141,
	       CASE_guard56369_0b0_theResult___snd65625_BITS__ETC__q142,
	       CASE_guard7296_0b0_sfd___37286_BITS_63_TO_41_0_ETC__q39,
	       CASE_guard7296_0b0_sfd___37286_BITS_63_TO_41_0_ETC__q40,
	       CASE_guard7822_0b0_sfd___37286_BITS_62_TO_40_0_ETC__q37,
	       CASE_guard7822_0b0_sfd___37286_BITS_62_TO_40_0_ETC__q38,
	       CASE_requestR_BITS_194_TO_192_0x1_8388607_0x2__ETC__q5,
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1073,
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1088,
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1456,
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1474,
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1680,
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1695,
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d4266,
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d4285,
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d4312,
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d4331,
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d588,
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d606;
  reg [10 : 0] CASE_guard0129_0b0_x0144_BITS_10_TO_0_0b1_theR_ETC__q76,
	       CASE_guard0129_0b0_x0144_BITS_10_TO_0_0b1_x014_ETC__q77,
	       CASE_guard02175_0b0_theResult___fst_exp11398_0_ETC__q163,
	       CASE_guard02175_0b0_theResult___fst_exp11398_0_ETC__q164,
	       CASE_guard0346_0b0_0_0b1_0_0b10_out_exp0965_0b_ETC__q86,
	       CASE_guard0346_0b0_0_0b1_theResult___exp0962_0_ETC__q87,
	       CASE_guard08246_0b0_0_0b1_0_0b10_out_exp08865__ETC__q32,
	       CASE_guard08246_0b0_0_0b1_theResult___exp08862_ETC__q33,
	       CASE_guard08975_0b0_x08990_BITS_10_TO_0_0b1_th_ETC__q109,
	       CASE_guard08975_0b0_x08990_BITS_10_TO_0_0b1_x0_ETC__q110,
	       CASE_guard1075_0b0_x1090_BITS_10_TO_0_0b1_theR_ETC__q89,
	       CASE_guard1075_0b0_x1090_BITS_10_TO_0_0b1_x109_ETC__q90,
	       CASE_guard5721_0b0_0_0b1_0_0b10_out_exp6340_0b_ETC__q106,
	       CASE_guard5721_0b0_0_0b1_theResult___exp6337_0_ETC__q105,
	       CASE_guard6451_0b0_x6466_BITS_10_TO_0_0b1_theR_ETC__q101,
	       CASE_guard6451_0b0_x6466_BITS_10_TO_0_0b1_x646_ETC__q102,
	       CASE_guard81312_0b0_theResult___fst_exp90506_0_ETC__q159,
	       CASE_guard81312_0b0_theResult___fst_exp90506_0_ETC__q160,
	       CASE_guard91853_0b0_theResult___fst_exp01334_0_ETC__q161,
	       CASE_guard91853_0b0_theResult___fst_exp01334_0_ETC__q162,
	       CASE_guard9399_0b0_0_0b1_0_0b10_out_exp0018_0b_ETC__q81,
	       CASE_guard9399_0b0_0_0b1_theResult___exp0015_0_ETC__q80,
	       CASE_requestR_BITS_194_TO_192_0x1_2046_0x2_IF__ETC__q6,
	       CASE_requestR_BITS_194_TO_192_0x3_IF_guard0346_ETC__q88,
	       CASE_requestR_BITS_194_TO_192_0x3_IF_guard0824_ETC__q34,
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2422,
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2451,
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2639,
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2961,
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2990,
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d3147,
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d4673,
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d4998,
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d5067;
  reg [7 : 0] CASE_guard1384_0b0_0_0b1_0_0b10_out_exp1800_0b_ETC__q57,
	      CASE_guard1384_0b0_0_0b1_theResult___exp1797_0_ETC__q58,
	      CASE_guard1910_0b0_x1925_BITS_7_TO_0_0b1_theRe_ETC__q60,
	      CASE_guard1910_0b0_x1925_BITS_7_TO_0_0b1_x1925_ETC__q61,
	      CASE_guard26038_0b0_theResult___fst_exp35390_0_ETC__q127,
	      CASE_guard26038_0b0_theResult___fst_exp35390_0_ETC__q128,
	      CASE_guard36028_0b0_theResult___fst_exp45309_0_ETC__q129,
	      CASE_guard36028_0b0_theResult___fst_exp45309_0_ETC__q130,
	      CASE_guard4468_0b0_0_0b1_0_0b10_out_exp4884_0b_ETC__q44,
	      CASE_guard4468_0b0_0_0b1_theResult___exp4881_0_ETC__q43,
	      CASE_guard46250_0b0_theResult___fst_exp55731_0_ETC__q131,
	      CASE_guard46250_0b0_theResult___fst_exp55731_0_ETC__q132,
	      CASE_guard4995_0b0_x5010_BITS_7_TO_0_0b1_theRe_ETC__q49,
	      CASE_guard4995_0b0_x5010_BITS_7_TO_0_0b1_x5010_ETC__q50,
	      CASE_guard5015_0b0_0_0b1_0_0b10_out_exp5434_0b_ETC__q18,
	      CASE_guard5015_0b0_0_0b1_theResult___exp5431_0_ETC__q17,
	      CASE_guard5545_0b0_x5560_BITS_7_TO_0_0b1_theRe_ETC__q19,
	      CASE_guard5545_0b0_x5560_BITS_7_TO_0_0b1_x5560_ETC__q20,
	      CASE_guard56369_0b0_theResult___fst_exp65679_0_ETC__q133,
	      CASE_guard56369_0b0_theResult___fst_exp65679_0_ETC__q134,
	      CASE_guard7296_0b0_0_0b1_0_0b10_out_exp7712_0b_ETC__q29,
	      CASE_guard7296_0b0_0_0b1_theResult___exp7709_0_ETC__q30,
	      CASE_guard7822_0b0_x7837_BITS_7_TO_0_0b1_theRe_ETC__q35,
	      CASE_guard7822_0b0_x7837_BITS_7_TO_0_0b1_x7837_ETC__q36,
	      CASE_requestR_BITS_194_TO_192_0x1_254_0x2_IF_r_ETC__q4,
	      CASE_requestR_BITS_194_TO_192_0x3_IF_guard1384_ETC__q59,
	      CASE_requestR_BITS_194_TO_192_0x3_IF_guard7296_ETC__q31,
	      IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1050,
	      IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1404,
	      IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1433,
	      IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1657,
	      IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d3719,
	      IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d3836,
	      IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d4163,
	      IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d4232,
	      IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d536,
	      IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d565;
  reg [2 : 0] IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d61;
  reg CASE_guard0129_0b0_requestR_BITS_191_TO_128_BI_ETC__q74,
      CASE_guard02175_0b0_requestR_BITS_191_TO_128_B_ETC__q169,
      CASE_guard26038_0b0_requestR_BITS_191_TO_128_B_ETC__q143,
      CASE_guard36028_0b0_requestR_BITS_191_TO_128_B_ETC__q145,
      CASE_guard4468_0b0_requestR_BITS_191_TO_128_BI_ETC__q45,
      CASE_guard46250_0b0_requestR_BITS_191_TO_128_B_ETC__q147,
      CASE_guard4995_0b0_requestR_BITS_191_TO_128_BI_ETC__q47,
      CASE_guard5015_0b0_requestR_BITS_191_TO_128_BI_ETC__q13,
      CASE_guard5545_0b0_requestR_BITS_191_TO_128_BI_ETC__q15,
      CASE_guard56369_0b0_requestR_BITS_191_TO_128_B_ETC__q149,
      CASE_guard5721_0b0_requestR_BITS_191_TO_128_BI_ETC__q97,
      CASE_guard6451_0b0_requestR_BITS_191_TO_128_BI_ETC__q99,
      CASE_guard81312_0b0_requestR_BITS_191_TO_128_B_ETC__q165,
      CASE_guard91853_0b0_requestR_BITS_191_TO_128_B_ETC__q167,
      CASE_guard9399_0b0_requestR_BITS_191_TO_128_BI_ETC__q72,
      CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q100,
      CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q14,
      CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q144,
      CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q146,
      CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q148,
      CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q150,
      CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q16,
      CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q166,
      CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q168,
      CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q170,
      CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q46,
      CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q48,
      CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q73,
      CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q75,
      CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q98;
  wire [117 : 0] IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d3224,
		 b__h110422,
		 x__h111322,
		 x__h112661;
  wire [88 : 0] IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1757,
		b__h43158,
		x__h44058,
		x__h45414;
  wire [85 : 0] IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2731,
		b__h82525,
		x__h83201,
		x__h84319;
  wire [64 : 0] _1_CONCAT_DONTCARE_CONCAT_IF_requestR_3_BIT_214_ETC___d97,
		_theResult_____2__h110357,
		_theResult_____2__h43093,
		out1___1__h111073,
		out1___1__h43809;
  wire [63 : 0] IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3__ETC___d1816,
		IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3__ETC___d1876,
		IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3__ETC___d2111,
		IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3__ETC___d2112,
		IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3__ETC___d2113,
		IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3__ETC___d2128,
		IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3__ETC___d2129,
		IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3__ETC___d2130,
		IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3__ETC___d2206,
		IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3__ETC___d2207,
		IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1745,
		IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1878,
		IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d3220,
		IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d3283,
		IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d3337,
		IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d5333,
		IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d5348,
		IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d5426,
		IF_NEG_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_re_ETC___d1812,
		IF_NEG_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_re_ETC___d1814,
		IF_NEG_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_re_ETC___d1874,
		IF_NEG_SEXT_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d3279,
		IF_NEG_SEXT_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d3281,
		IF_NEG_SEXT_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d3335,
		requestR_BITS_127_TO_64__q3,
		requestR_BITS_191_TO_128__q1,
		requestR_BITS_63_TO_0__q8,
		res___1__h229866,
		res___1__h230304,
		res___1__h230314,
		res___1__h230333,
		res___1__h57534,
		res___1__h57770,
		res___1__h57780,
		res___1__h57799,
		res__h166745,
		res__h212818,
		res__h217300,
		res__h221886,
		res__h224628,
		res__h227363,
		res__h229280,
		res__h230349,
		res__h230541,
		res__h3932,
		res__h48859,
		res__h49096,
		res__h54627,
		res__h56150,
		res__h57259,
		res__h57815,
		sfd___3__h15005,
		sfd___3__h27286,
		sfd__h3990,
		x__h110179,
		x__h112240,
		x__h113022,
		x__h16727,
		x__h167888,
		x__h213882,
		x__h218468,
		x__h222950,
		x__h225685,
		x__h227602,
		x__h229846,
		x__h230460,
		x__h28828,
		x__h3429,
		x__h36028,
		x__h3605,
		x__h3778,
		x__h42915,
		x__h44993,
		x__h45775,
		x__h47391,
		x__h48180,
		x__h50854,
		x__h53419,
		x__h53579,
		x__h53757,
		x__h55280,
		x__h56389,
		x__h57514,
		x__h59668,
		x__h59829,
		x__h59992,
		x__h60162,
		x__h71361,
		x__h82279,
		x__h83895,
		x__h84681,
		x__h97683;
  wire [56 : 0] IF_0_CONCAT_IF_IF_0b0_CONCAT_NOT_IF_requestR_3_ETC__q117,
		IF_0_CONCAT_IF_IF_3074_MINUS_SEXT_IF_IF_reques_ETC__q154,
		IF_0_CONCAT_IF_IF_3970_MINUS_SEXT_IF_requestR__ETC__q122,
		IF_0_CONCAT_IF_IF_IF_requestR_3_BIT_214_4_THEN_ETC__q151,
		IF_0_CONCAT_IF_IF_IF_requestR_3_BIT_214_4_THEN_ETC__q157,
		IF_0_CONCAT_IF_IF_requestR_3_BIT_214_4_THEN_re_ETC__q119,
		IF_0_CONCAT_IF_IF_requestR_3_BIT_214_4_THEN_re_ETC__q125,
		IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1908,
		_0b0_CONCAT_NOT_IF_IF_requestR_3_BIT_214_4_THEN_ETC___d4691,
		_0b0_CONCAT_NOT_IF_requestR_3_BIT_214_4_THEN_re_ETC___d3858,
		_theResult____h126028,
		_theResult____h146240,
		_theResult____h191843,
		_theResult___snd__h135401,
		_theResult___snd__h135412,
		_theResult___snd__h135414,
		_theResult___snd__h135424,
		_theResult___snd__h135430,
		_theResult___snd__h135453,
		_theResult___snd__h145260,
		_theResult___snd__h145262,
		_theResult___snd__h145269,
		_theResult___snd__h145275,
		_theResult___snd__h145298,
		_theResult___snd__h155742,
		_theResult___snd__h155753,
		_theResult___snd__h155755,
		_theResult___snd__h155765,
		_theResult___snd__h155771,
		_theResult___snd__h155794,
		_theResult___snd__h165625,
		_theResult___snd__h165639,
		_theResult___snd__h165645,
		_theResult___snd__h165663,
		_theResult___snd__h190457,
		_theResult___snd__h190459,
		_theResult___snd__h190466,
		_theResult___snd__h190472,
		_theResult___snd__h190495,
		_theResult___snd__h201345,
		_theResult___snd__h201356,
		_theResult___snd__h201358,
		_theResult___snd__h201368,
		_theResult___snd__h201374,
		_theResult___snd__h201397,
		_theResult___snd__h211344,
		_theResult___snd__h211358,
		_theResult___snd__h211364,
		_theResult___snd__h211382,
		b__h46021,
		result__h146853,
		result__h192456,
		sfd__h117253,
		sfdin__h135384,
		sfdin__h155725,
		sfdin__h201328,
		x__h146948,
		x__h192551,
		x__h46697,
		x__h47815;
  wire [54 : 0] sfd___3__h69389, sfd___3__h80336, sfd__h60177, sfd__h71373;
  wire [53 : 0] sfd__h108263,
		sfd__h109005,
		sfd__h190524,
		sfd__h201426,
		sfd__h211417,
		sfd__h69416,
		sfd__h70159,
		sfd__h80363,
		sfd__h81105,
		sfd__h95738,
		sfd__h96481,
		value__h82527;
  wire [51 : 0] IF_IF_IF_IF_3074_MINUS_SEXT_IF_IF_requestR_3_B_ETC___d5121,
		IF_IF_IF_IF_3074_MINUS_SEXT_IF_IF_requestR_3_B_ETC___d5123,
		IF_IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d5094,
		IF_IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d5096,
		IF_IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d5140,
		IF_IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d5142,
		IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d2468,
		IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d2470,
		IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d2486,
		IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d2488,
		IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d3007,
		IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d3009,
		IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d3025,
		IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d3027,
		IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3__ETC___d5153,
		IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2496,
		IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2680,
		_theResult___fst_sfd__h108959,
		_theResult___fst_sfd__h109714,
		_theResult___fst_sfd__h109717,
		_theResult___fst_sfd__h113549,
		_theResult___fst_sfd__h174201,
		_theResult___fst_sfd__h191260,
		_theResult___fst_sfd__h191263,
		_theResult___fst_sfd__h202162,
		_theResult___fst_sfd__h202165,
		_theResult___fst_sfd__h212177,
		_theResult___fst_sfd__h212180,
		_theResult___fst_sfd__h212189,
		_theResult___fst_sfd__h212195,
		_theResult___fst_sfd__h70113,
		_theResult___fst_sfd__h70869,
		_theResult___fst_sfd__h70872,
		_theResult___fst_sfd__h81059,
		_theResult___fst_sfd__h81814,
		_theResult___fst_sfd__h81817,
		_theResult___fst_sfd__h96435,
		_theResult___fst_sfd__h97191,
		_theResult___fst_sfd__h97194,
		_theResult___sfd__h108863,
		_theResult___sfd__h109618,
		_theResult___sfd__h191162,
		_theResult___sfd__h202064,
		_theResult___sfd__h212079,
		_theResult___sfd__h70016,
		_theResult___sfd__h70772,
		_theResult___sfd__h80963,
		_theResult___sfd__h81718,
		_theResult___sfd__h96338,
		_theResult___sfd__h97094,
		_theResult___snd_fst_sfd__h109720,
		_theResult___snd_fst_sfd__h169840,
		_theResult___snd_fst_sfd__h191266,
		_theResult___snd_fst_sfd__h212183,
		_theResult___snd_fst_sfd__h70875,
		_theResult___snd_fst_sfd__h81820,
		_theResult___snd_fst_sfd__h97197,
		out___1_sfd__h167954,
		out_sfd__h108866,
		out_sfd__h109621,
		out_sfd__h191165,
		out_sfd__h202067,
		out_sfd__h212082,
		out_sfd__h70019,
		out_sfd__h70775,
		out_sfd__h80966,
		out_sfd__h81721,
		out_sfd__h96341,
		out_sfd__h97097,
		value__h113092;
  wire [32 : 0] _theResult_____2__h45956,
		_theResult_____2__h82460,
		out1___1__h46448,
		out1___1__h82952;
  wire [31 : 0] IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3__ETC___d1967,
		IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3__ETC___d2022,
		IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3__ETC___d2108,
		IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3__ETC___d2109,
		IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3__ETC___d2123,
		IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3__ETC___d2125,
		IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3__ETC___d2126,
		IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1904,
		IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2024,
		IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2719,
		IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2790,
		IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2851,
		IF_NEG_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_re_ETC___d1963,
		IF_NEG_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_re_ETC___d1965,
		IF_NEG_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_re_ETC___d2020,
		IF_NEG_SEXT_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d2786,
		IF_NEG_SEXT_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d2788,
		IF_NEG_SEXT_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d2849,
		IF_NOT_IF_IF_requestR_3_BIT_214_4_THEN_request_ETC___d2106,
		IF_NOT_IF_IF_requestR_3_BIT_214_4_THEN_request_ETC___d2122,
		IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d48,
		requestR_BITS_191_TO_128_BITS_31_TO_0__q2,
		sfd___3__h34458,
		sfd___3__h41374,
		sfd__h28849,
		x__h166751,
		x__h28834,
		x__h3436,
		x__h3612,
		x__h3785,
		x__h3975,
		x__h45778,
		x__h47394,
		x__h82282,
		x__h83898;
  wire [30 : 0] IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d37;
  wire [24 : 0] sfd__h135482,
		sfd__h145327,
		sfd__h15032,
		sfd__h15575,
		sfd__h155823,
		sfd__h165698,
		sfd__h27313,
		sfd__h27852,
		sfd__h34485,
		sfd__h35025,
		sfd__h41401,
		sfd__h41940,
		value__h43160;
  wire [23 : 0] NEG_SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d2724,
		NEG_SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d2756,
		NEG_SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d2757,
		NEG_SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d2822,
		NEG_SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d3249,
		NEG_SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d3250,
		NEG_SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d3308;
  wire [22 : 0] IF_IF_IF_IF_0b0_CONCAT_NOT_IF_requestR_3_BIT_2_ETC___d4260,
		IF_IF_IF_IF_0b0_CONCAT_NOT_IF_requestR_3_BIT_2_ETC___d4262,
		IF_IF_IF_IF_3970_MINUS_SEXT_IF_requestR_3_BIT__ETC___d4306,
		IF_IF_IF_IF_3970_MINUS_SEXT_IF_requestR_3_BIT__ETC___d4308,
		IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d1450,
		IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d1452,
		IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d1468,
		IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d1470,
		IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d4279,
		IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d4281,
		IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d4325,
		IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d4327,
		IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d582,
		IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d584,
		IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d600,
		IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d602,
		IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d4338,
		_theResult___fst_sfd__h126011,
		_theResult___fst_sfd__h136015,
		_theResult___fst_sfd__h136018,
		_theResult___fst_sfd__h145860,
		_theResult___fst_sfd__h145863,
		_theResult___fst_sfd__h15529,
		_theResult___fst_sfd__h156356,
		_theResult___fst_sfd__h156359,
		_theResult___fst_sfd__h16082,
		_theResult___fst_sfd__h16085,
		_theResult___fst_sfd__h166255,
		_theResult___fst_sfd__h166258,
		_theResult___fst_sfd__h166267,
		_theResult___fst_sfd__h166273,
		_theResult___fst_sfd__h168212,
		_theResult___fst_sfd__h27806,
		_theResult___fst_sfd__h28358,
		_theResult___fst_sfd__h28361,
		_theResult___fst_sfd__h34979,
		_theResult___fst_sfd__h35532,
		_theResult___fst_sfd__h35535,
		_theResult___fst_sfd__h41894,
		_theResult___fst_sfd__h42446,
		_theResult___fst_sfd__h42449,
		_theResult___sfd__h135917,
		_theResult___sfd__h145762,
		_theResult___sfd__h15432,
		_theResult___sfd__h156258,
		_theResult___sfd__h15985,
		_theResult___sfd__h166157,
		_theResult___sfd__h27710,
		_theResult___sfd__h28262,
		_theResult___sfd__h34882,
		_theResult___sfd__h35435,
		_theResult___sfd__h41798,
		_theResult___sfd__h42350,
		_theResult___snd_fst_sfd__h117207,
		_theResult___snd_fst_sfd__h145866,
		_theResult___snd_fst_sfd__h16088,
		_theResult___snd_fst_sfd__h166261,
		_theResult___snd_fst_sfd__h28364,
		_theResult___snd_fst_sfd__h35538,
		_theResult___snd_fst_sfd__h42452,
		out_sfd__h135920,
		out_sfd__h145765,
		out_sfd__h15435,
		out_sfd__h156261,
		out_sfd__h15988,
		out_sfd__h166160,
		out_sfd__h27713,
		out_sfd__h28265,
		out_sfd__h34885,
		out_sfd__h35438,
		out_sfd__h41801,
		out_sfd__h42353,
		sV1_sfd__h1473,
		sV2_sfd__h1598,
		value__h167957;
  wire [19 : 0] NEG_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d1750,
		NEG_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d1782,
		NEG_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d1783,
		NEG_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d1847,
		NEG_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d1933,
		NEG_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d1934,
		NEG_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d1993;
  wire [11 : 0] IF_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_reques_ETC___d5007,
		SEXT_IF_IF_requestR_3_BIT_214_4_THEN_requestR__ETC___d4684,
		SEXT_IF_IF_requestR_3_BIT_214_4_THEN_requestR__ETC__q153,
		SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_3_B_ETC___d3851,
		SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_3_B_ETC__q121,
		_3074_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_ETC___d3420,
		_3074_MINUS_SEXT_IF_IF_requestR_3_BIT_214_4_THE_ETC___d4687,
		_32_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d2342,
		_32_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d2558,
		_3970_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_21_ETC___d4541,
		_3970_MINUS_SEXT_IF_requestR_3_BIT_214_4_THEN_r_ETC___d3854,
		_64_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d2882,
		_64_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d3068,
		x__h108990,
		x__h146981,
		x__h192584,
		x__h70144,
		x__h81090,
		x__h96466;
  wire [10 : 0] IF_IF_IF_IF_3074_MINUS_SEXT_IF_IF_requestR_3_B_ETC___d4992,
		IF_IF_IF_IF_3074_MINUS_SEXT_IF_IF_requestR_3_B_ETC___d4994,
		IF_IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d4667,
		IF_IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d4669,
		IF_IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d5061,
		IF_IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d5063,
		IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d2419,
		IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d2445,
		IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d2447,
		IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d2958,
		IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d2984,
		IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d2986,
		IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2996,
		IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d2722,
		SEXT_IF_IF_requestR_3_BIT_214_4_THEN_requestR__ETC__q156,
		_theResult___exp__h108862,
		_theResult___exp__h109617,
		_theResult___exp__h191161,
		_theResult___exp__h202063,
		_theResult___exp__h212078,
		_theResult___exp__h70015,
		_theResult___exp__h70771,
		_theResult___exp__h80962,
		_theResult___exp__h81717,
		_theResult___exp__h96337,
		_theResult___exp__h97093,
		_theResult___fst_exp__h108958,
		_theResult___fst_exp__h109713,
		_theResult___fst_exp__h109716,
		_theResult___fst_exp__h174200,
		_theResult___fst_exp__h190497,
		_theResult___fst_exp__h190503,
		_theResult___fst_exp__h190506,
		_theResult___fst_exp__h191259,
		_theResult___fst_exp__h191262,
		_theResult___fst_exp__h201334,
		_theResult___fst_exp__h201399,
		_theResult___fst_exp__h201405,
		_theResult___fst_exp__h201408,
		_theResult___fst_exp__h202161,
		_theResult___fst_exp__h202164,
		_theResult___fst_exp__h211350,
		_theResult___fst_exp__h211389,
		_theResult___fst_exp__h211395,
		_theResult___fst_exp__h211398,
		_theResult___fst_exp__h212176,
		_theResult___fst_exp__h212179,
		_theResult___fst_exp__h212188,
		_theResult___fst_exp__h212191,
		_theResult___fst_exp__h70112,
		_theResult___fst_exp__h70868,
		_theResult___fst_exp__h70871,
		_theResult___fst_exp__h81058,
		_theResult___fst_exp__h81813,
		_theResult___fst_exp__h81816,
		_theResult___fst_exp__h96434,
		_theResult___fst_exp__h97190,
		_theResult___fst_exp__h97193,
		_theResult___snd_fst_exp__h109719,
		_theResult___snd_fst_exp__h109722,
		_theResult___snd_fst_exp__h109725,
		_theResult___snd_fst_exp__h191265,
		_theResult___snd_fst_exp__h212182,
		_theResult___snd_fst_exp__h70874,
		_theResult___snd_fst_exp__h70877,
		_theResult___snd_fst_exp__h70880,
		_theResult___snd_fst_exp__h81819,
		_theResult___snd_fst_exp__h81822,
		_theResult___snd_fst_exp__h81825,
		_theResult___snd_fst_exp__h97196,
		_theResult___snd_fst_exp__h97199,
		_theResult___snd_fst_exp__h97202,
		din_inc___2_exp__h109755,
		din_inc___2_exp__h212214,
		din_inc___2_exp__h212244,
		din_inc___2_exp__h212268,
		din_inc___2_exp__h70914,
		din_inc___2_exp__h81855,
		din_inc___2_exp__h97236,
		out_exp__h108865,
		out_exp__h109620,
		out_exp__h191164,
		out_exp__h202066,
		out_exp__h212081,
		out_exp__h70018,
		out_exp__h70774,
		out_exp__h80965,
		out_exp__h81720,
		out_exp__h96340,
		out_exp__h97096,
		x__h167898;
  wire [8 : 0] IF_SEXT_IF_requestR_3_BIT_214_4_THEN_requestR__ETC___d4172,
	       _32_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d1321,
	       _32_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d1577,
	       _64_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d444,
	       _64_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d969,
	       x__h15560,
	       x__h27837,
	       x__h35010,
	       x__h41925;
  wire [7 : 0] IF_IF_IF_IF_0b0_CONCAT_NOT_IF_requestR_3_BIT_2_ETC___d3713,
	       IF_IF_IF_IF_0b0_CONCAT_NOT_IF_requestR_3_BIT_2_ETC___d3715,
	       IF_IF_IF_IF_3970_MINUS_SEXT_IF_requestR_3_BIT__ETC___d4157,
	       IF_IF_IF_IF_3970_MINUS_SEXT_IF_requestR_3_BIT__ETC___d4159,
	       IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d1401,
	       IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d1427,
	       IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d1429,
	       IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d3830,
	       IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d3832,
	       IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d4226,
	       IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d4228,
	       IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d533,
	       IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d559,
	       IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d561,
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1439,
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1748,
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d571,
	       SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_3_B_ETC__q124,
	       _theResult___exp__h135916,
	       _theResult___exp__h145761,
	       _theResult___exp__h15431,
	       _theResult___exp__h156257,
	       _theResult___exp__h15984,
	       _theResult___exp__h166156,
	       _theResult___exp__h27709,
	       _theResult___exp__h28261,
	       _theResult___exp__h34881,
	       _theResult___exp__h35434,
	       _theResult___exp__h41797,
	       _theResult___exp__h42349,
	       _theResult___fst_exp__h126010,
	       _theResult___fst_exp__h135390,
	       _theResult___fst_exp__h135455,
	       _theResult___fst_exp__h135461,
	       _theResult___fst_exp__h135464,
	       _theResult___fst_exp__h136014,
	       _theResult___fst_exp__h136017,
	       _theResult___fst_exp__h145300,
	       _theResult___fst_exp__h145306,
	       _theResult___fst_exp__h145309,
	       _theResult___fst_exp__h145859,
	       _theResult___fst_exp__h145862,
	       _theResult___fst_exp__h15528,
	       _theResult___fst_exp__h155731,
	       _theResult___fst_exp__h155796,
	       _theResult___fst_exp__h155802,
	       _theResult___fst_exp__h155805,
	       _theResult___fst_exp__h156355,
	       _theResult___fst_exp__h156358,
	       _theResult___fst_exp__h16081,
	       _theResult___fst_exp__h16084,
	       _theResult___fst_exp__h165631,
	       _theResult___fst_exp__h165670,
	       _theResult___fst_exp__h165676,
	       _theResult___fst_exp__h165679,
	       _theResult___fst_exp__h166254,
	       _theResult___fst_exp__h166257,
	       _theResult___fst_exp__h166266,
	       _theResult___fst_exp__h166269,
	       _theResult___fst_exp__h27805,
	       _theResult___fst_exp__h28357,
	       _theResult___fst_exp__h28360,
	       _theResult___fst_exp__h34978,
	       _theResult___fst_exp__h35531,
	       _theResult___fst_exp__h35534,
	       _theResult___fst_exp__h41893,
	       _theResult___fst_exp__h42445,
	       _theResult___fst_exp__h42448,
	       _theResult___snd_fst_exp__h145865,
	       _theResult___snd_fst_exp__h16087,
	       _theResult___snd_fst_exp__h16090,
	       _theResult___snd_fst_exp__h16093,
	       _theResult___snd_fst_exp__h166260,
	       _theResult___snd_fst_exp__h28363,
	       _theResult___snd_fst_exp__h28366,
	       _theResult___snd_fst_exp__h28369,
	       _theResult___snd_fst_exp__h35537,
	       _theResult___snd_fst_exp__h35540,
	       _theResult___snd_fst_exp__h35543,
	       _theResult___snd_fst_exp__h42451,
	       _theResult___snd_fst_exp__h42454,
	       _theResult___snd_fst_exp__h42457,
	       din_inc___2_exp__h16127,
	       din_inc___2_exp__h166288,
	       din_inc___2_exp__h166312,
	       din_inc___2_exp__h166342,
	       din_inc___2_exp__h166366,
	       din_inc___2_exp__h28399,
	       din_inc___2_exp__h35577,
	       din_inc___2_exp__h42487,
	       out_exp__h135919,
	       out_exp__h145764,
	       out_exp__h15434,
	       out_exp__h156260,
	       out_exp__h15987,
	       out_exp__h166159,
	       out_exp__h27712,
	       out_exp__h28264,
	       out_exp__h34884,
	       out_exp__h35437,
	       out_exp__h41800,
	       out_exp__h42352,
	       sV1_exp__h1472,
	       sV2_exp__h1597,
	       x__h113032;
  wire [6 : 0] IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3__ETC___d441,
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d966,
	       requestR_BITS_206_TO_200__q177;
  wire [5 : 0] IF_IF_0b0_CONCAT_NOT_IF_requestR_3_BIT_214_4_T_ETC___d3654,
	       IF_IF_3074_MINUS_SEXT_IF_IF_requestR_3_BIT_214_ETC___d4933,
	       IF_IF_3970_MINUS_SEXT_IF_requestR_3_BIT_214_4__ETC___d4098,
	       IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3__ETC___d1318,
	       IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3__ETC___d2339,
	       IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3__ETC___d4613,
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1574,
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2555,
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d3776;
  wire [4 : 0] _0_CONCAT_IF_IF_0b0_CONCAT_NOT_IF_requestR_3_BI_ETC___d4396,
	       _0_CONCAT_IF_IF_3074_MINUS_SEXT_IF_IF_requestR__ETC___d5220,
	       _0_CONCAT_IF_IF_3970_MINUS_SEXT_IF_requestR_3_B_ETC___d4425,
	       _0_CONCAT_IF_IF_IF_requestR_3_BIT_214_4_THEN_re_ETC___d5203,
	       _0_CONCAT_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d4408,
	       fcsr__h3933,
	       x__h109855,
	       x__h111943,
	       x__h112739,
	       x__h166866,
	       x__h212920,
	       x__h217430,
	       x__h227382,
	       x__h28503,
	       x__h35703,
	       x__h42591,
	       x__h44696,
	       x__h45492,
	       x__h47094,
	       x__h47893,
	       x__h50220,
	       x__h56169,
	       x__h71036,
	       x__h81955,
	       x__h83598,
	       x__h84397,
	       x__h97358;
  wire [1 : 0] IF_sfd___30336_BIT_1_THEN_2_ELSE_0__q85,
	       IF_sfd___30336_BIT_2_THEN_2_ELSE_0__q84,
	       IF_sfd___31374_BIT_7_THEN_2_ELSE_0__q56,
	       IF_sfd___31374_BIT_8_THEN_2_ELSE_0__q55,
	       IF_sfd___34458_BIT_7_THEN_2_ELSE_0__q42,
	       IF_sfd___34458_BIT_8_THEN_2_ELSE_0__q41,
	       IF_sfd___35005_BIT_10_THEN_2_ELSE_0__q12,
	       IF_sfd___35005_BIT_11_THEN_2_ELSE_0__q11,
	       IF_sfd___35005_BIT_39_THEN_2_ELSE_0__q10,
	       IF_sfd___35005_BIT_40_THEN_2_ELSE_0__q9,
	       IF_sfd___37286_BIT_10_THEN_2_ELSE_0__q28,
	       IF_sfd___37286_BIT_11_THEN_2_ELSE_0__q27,
	       IF_sfd___37286_BIT_39_THEN_2_ELSE_0__q26,
	       IF_sfd___37286_BIT_40_THEN_2_ELSE_0__q25,
	       IF_sfd___39389_BIT_1_THEN_2_ELSE_0__q71,
	       IF_sfd___39389_BIT_2_THEN_2_ELSE_0__q70,
	       IF_sfdin01328_BIT_4_THEN_2_ELSE_0__q155,
	       IF_sfdin35384_BIT_33_THEN_2_ELSE_0__q118,
	       IF_sfdin55725_BIT_33_THEN_2_ELSE_0__q123,
	       IF_theResult___snd11344_BIT_4_THEN_2_ELSE_0__q158,
	       IF_theResult___snd45260_BIT_33_THEN_2_ELSE_0__q120,
	       IF_theResult___snd65625_BIT_33_THEN_2_ELSE_0__q126,
	       IF_theResult___snd90457_BIT_4_THEN_2_ELSE_0__q152,
	       IF_x11322_BIT_53_THEN_2_ELSE_0__q115,
	       IF_x12661_BIT_53_THEN_2_ELSE_0__q116,
	       IF_x3201_BIT_53_THEN_2_ELSE_0__q95,
	       IF_x4058_BIT_24_THEN_2_ELSE_0__q66,
	       IF_x4319_BIT_53_THEN_2_ELSE_0__q96,
	       IF_x5414_BIT_24_THEN_2_ELSE_0__q67,
	       IF_x6697_BIT_24_THEN_2_ELSE_0__q68,
	       IF_x7815_BIT_24_THEN_2_ELSE_0__q69,
	       guard__h108246,
	       guard__h108975,
	       guard__h110355,
	       guard__h111133,
	       guard__h112440,
	       guard__h126038,
	       guard__h136028,
	       guard__h146250,
	       guard__h15015,
	       guard__h15545,
	       guard__h156369,
	       guard__h181312,
	       guard__h191853,
	       guard__h202175,
	       guard__h27296,
	       guard__h27822,
	       guard__h34468,
	       guard__h34995,
	       guard__h41384,
	       guard__h41910,
	       guard__h43091,
	       guard__h43869,
	       guard__h45193,
	       guard__h45954,
	       guard__h46508,
	       guard__h47594,
	       guard__h69399,
	       guard__h70129,
	       guard__h80346,
	       guard__h81075,
	       guard__h82458,
	       guard__h83012,
	       guard__h84098,
	       guard__h95721,
	       guard__h96451;
  wire IF_3074_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_21_ETC___d4358,
       IF_32_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_2_ETC___d1379,
       IF_32_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_2_ETC___d1529,
       IF_32_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_2_ETC___d2398,
       IF_32_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_2_ETC___d2513,
       IF_32_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214__ETC___d1718,
       IF_32_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214__ETC___d2697,
       IF_64_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_2_ETC___d2937,
       IF_64_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_2_ETC___d3054,
       IF_64_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_2_ETC___d511,
       IF_64_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_2_ETC___d693,
       IF_64_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214__ETC___d1174,
       IF_64_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214__ETC___d3208,
       IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3__ETC___d5188,
       IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3__ETC___d5189,
       IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3__ETC___d5224,
       IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3__ETC___d5227,
       IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3__ETC___d5234,
       IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3__ETC___d5248,
       IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3__ETC___d5260,
       IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3__ETC___d5272,
       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1520,
       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1523,
       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1532,
       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1774,
       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1806,
       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1868,
       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1885,
       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1896,
       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1925,
       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1957,
       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2014,
       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2032,
       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2043,
       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2067,
       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2077,
       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2081,
       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2090,
       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2091,
       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2092,
       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2095,
       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2097,
       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2115,
       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2156,
       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2167,
       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2171,
       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2748,
       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2780,
       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2843,
       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d3045,
       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d3048,
       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d3057,
       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d3241,
       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d3273,
       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d3329,
       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d4378,
       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d4429,
       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d4440,
       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d4456,
       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d4469,
       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d4482,
       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d4617,
       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d5010,
       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d5326,
       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d684,
       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d687,
       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d696,
       IF_NEG_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_re_ETC___d1837,
       IF_NEG_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_re_ETC___d1983,
       IF_NEG_SEXT_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d2812,
       IF_NEG_SEXT_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d3298,
       IF_NOT_32_MINUS_0_CONCAT_IF_IF_IF_requestR_3_B_ETC___d2399,
       IF_NOT_3970_MINUS_0_CONCAT_IF_IF_IF_requestR_3_ETC___d5169,
       IF_NOT_IF_requestR_3_BIT_214_4_THEN_requestR_3_ETC___d2101,
       IF_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_reques_ETC___d5186,
       IF_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_reques_ETC___d5246,
       IF_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_reques_ETC___d5258,
       IF_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_reques_ETC___d5270,
       IF_SEXT_IF_requestR_3_BIT_214_4_THEN_requestR__ETC___d4376,
       IF_SEXT_IF_requestR_3_BIT_214_4_THEN_requestR__ETC___d4454,
       IF_SEXT_IF_requestR_3_BIT_214_4_THEN_requestR__ETC___d4467,
       IF_SEXT_IF_requestR_3_BIT_214_4_THEN_requestR__ETC___d4480,
       IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d1165,
       IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d1168,
       IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d1177,
       IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d1709,
       IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d1712,
       IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d1721,
       IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d2103,
       IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d2169,
       IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d2861,
       IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d2872,
       IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d3199,
       IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d3202,
       IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d3211,
       IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d3346,
       IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d3357,
       IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d5294,
       IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d5302,
       IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d5306,
       IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d5315,
       IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d5317,
       IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d5318,
       IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d5322,
       IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d5323,
       IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d5339,
       IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d5363,
       IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d5373,
       IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d5378,
       NEG_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d1785,
       NEG_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d1849,
       NEG_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d1936,
       NEG_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d1995,
       NEG_SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d2759,
       NEG_SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d2824,
       NEG_SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d3252,
       NEG_SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d3310,
       NOT_3074_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_2_ETC___d4448,
       NOT_3074_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_2_ETC___d4476,
       NOT_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_ETC___d1326,
       NOT_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_ETC___d1826,
       NOT_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_ETC___d1890,
       NOT_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_ETC___d1975,
       NOT_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_ETC___d2037,
       NOT_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_ETC___d2104,
       NOT_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_ETC___d2105,
       NOT_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_ETC___d2166,
       NOT_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_ETC___d2172,
       NOT_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_ETC___d2192,
       NOT_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_ETC___d2887,
       NOT_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_ETC___d449,
       NOT_IF_requestR_3_BIT_214_4_THEN_requestR_3_BI_ETC___d1059,
       NOT_IF_requestR_3_BIT_214_4_THEN_requestR_3_BI_ETC___d1666,
       NOT_IF_requestR_3_BIT_214_4_THEN_requestR_3_BI_ETC___d2801,
       NOT_IF_requestR_3_BIT_214_4_THEN_requestR_3_BI_ETC___d2866,
       NOT_IF_requestR_3_BIT_214_4_THEN_requestR_3_BI_ETC___d3156,
       NOT_IF_requestR_3_BIT_214_4_THEN_requestR_3_BI_ETC___d3290,
       NOT_IF_requestR_3_BIT_214_4_THEN_requestR_3_BI_ETC___d3351,
       NOT_IF_requestR_3_BIT_214_4_THEN_requestR_3_BI_ETC___d5330,
       NOT_IF_requestR_3_BIT_214_4_THEN_requestR_3_BI_ETC___d5374,
       NOT_IF_requestR_3_BIT_214_4_THEN_requestR_3_BI_ETC___d5399,
       NOT_verbosity_ULE_1_6___d27,
       NOT_verbosity_ULE_2_01___d702,
       SEXT_IF_IF_requestR_3_BIT_214_4_THEN_requestR__ETC___d4685,
       SEXT_IF_IF_requestR_3_BIT_214_4_THEN_requestR__ETC___d4686,
       SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_3_B_ETC___d3852,
       SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_3_B_ETC___d3853,
       _0_CONCAT_IF_IF_0b0_CONCAT_NOT_IF_requestR_3_BI_ETC___d3656,
       _0_CONCAT_IF_IF_3074_MINUS_SEXT_IF_IF_requestR__ETC___d4935,
       _0_CONCAT_IF_IF_3970_MINUS_SEXT_IF_requestR_3_B_ETC___d4100,
       _0_CONCAT_IF_IF_IF_requestR_3_BIT_214_4_THEN_re_ETC___d4615,
       _0_CONCAT_IF_IF_IF_requestR_3_BIT_214_4_THEN_re_ETC___d5008,
       _0_CONCAT_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d3778,
       _0_CONCAT_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d4173,
       _3074_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_ETC___d3421,
       _3074_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_ETC___d3422,
       _3074_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_ETC___d4411,
       _3074_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_ETC___d4436,
       _3074_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_ETC___d4463,
       _32_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d1322,
       _32_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d1324,
       _32_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d1327,
       _32_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d2343,
       _32_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d2345,
       _32_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d2347,
       _32_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d1578,
       _32_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d1579,
       _32_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d1580,
       _32_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d2559,
       _32_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d2560,
       _32_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d2561,
       _3970_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_21_ETC___d4542,
       _3970_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_21_ETC___d4543,
       _64_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d2883,
       _64_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d2885,
       _64_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d2888,
       _64_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d445,
       _64_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d447,
       _64_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d450,
       _64_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d3069,
       _64_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d3070,
       _64_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d3071,
       _64_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d970,
       _64_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d971,
       _64_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d972,
       guard__h146848,
       guard__h192451;
  // action method server_reset_request_put
  assign RDY_server_reset_request_put = resetReqsF$FULL_N ;
  assign CAN_FIRE_server_reset_request_put = resetReqsF$FULL_N ;
  assign WILL_FIRE_server_reset_request_put = EN_server_reset_request_put ;
  // action method server_reset_response_get
  assign RDY_server_reset_response_get = resetRspsF$EMPTY_N ;
  assign CAN_FIRE_server_reset_response_get = resetRspsF$EMPTY_N ;
  assign WILL_FIRE_server_reset_response_get = EN_server_reset_response_get ;
  // action method req
  assign CAN_FIRE_req = 1'd1 ;
  assign WILL_FIRE_req = EN_req ;
  // value method valid
  assign valid = dw_valid$whas && dw_valid$wget ;
  // value method word_fst
  assign word_fst = dw_result$wget[68:5] ;
  // value method word_snd
  assign word_snd = dw_result$wget[4:0] ;
  // submodule fpu
  mkFPU fpu(.CLK(CLK),
	    .RST_N(RST_N),
	    .server_core_request_put(fpu$server_core_request_put),
	    .EN_server_core_request_put(fpu$EN_server_core_request_put),
	    .EN_server_core_response_get(fpu$EN_server_core_response_get),
	    .EN_server_reset_request_put(fpu$EN_server_reset_request_put),
	    .EN_server_reset_response_get(fpu$EN_server_reset_response_get),
	    .RDY_server_core_request_put(fpu$RDY_server_core_request_put),
	    .server_core_response_get(fpu$server_core_response_get),
	    .RDY_server_core_response_get(fpu$RDY_server_core_response_get),
	    .RDY_server_reset_request_put(fpu$RDY_server_reset_request_put),
	    .RDY_server_reset_response_get(fpu$RDY_server_reset_response_get));
  // submodule frmFpuF
  FIFO2 #(.width(32'd1), .guarded(1'd1)) frmFpuF(.RST(RST_N),
						 .CLK(CLK),
						 .D_IN(frmFpuF$D_IN),
						 .ENQ(frmFpuF$ENQ),
						 .DEQ(frmFpuF$DEQ),
						 .CLR(frmFpuF$CLR),
						 .D_OUT(),
						 .FULL_N(),
						 .EMPTY_N());
  // submodule resetReqsF
  FIFO20 #(.guarded(1'd1)) resetReqsF(.RST(RST_N),
				      .CLK(CLK),
				      .ENQ(resetReqsF$ENQ),
				      .DEQ(resetReqsF$DEQ),
				      .CLR(resetReqsF$CLR),
				      .FULL_N(resetReqsF$FULL_N),
				      .EMPTY_N(resetReqsF$EMPTY_N));
  // submodule resetRspsF
  FIFO20 #(.guarded(1'd1)) resetRspsF(.RST(RST_N),
				      .CLK(CLK),
				      .ENQ(resetRspsF$ENQ),
				      .DEQ(resetRspsF$DEQ),
				      .CLR(resetRspsF$CLR),
				      .FULL_N(resetRspsF$FULL_N),
				      .EMPTY_N(resetRspsF$EMPTY_N));
  // rule RL_rl_reset_end
  assign CAN_FIRE_RL_rl_reset_end =
	     fpu$RDY_server_reset_response_get && resetRspsF$FULL_N &&
	     stateR == 2'd0 ;
  assign WILL_FIRE_RL_rl_reset_end = CAN_FIRE_RL_rl_reset_end ;
  // rule RL_doFADD_S
  assign CAN_FIRE_RL_doFADD_S =
	     fpu$RDY_server_core_request_put && requestR[214] &&
	     stateR == 2'd1 &&
	     requestR[213:207] == 7'b1010011 &&
	     requestR[206:200] == 7'h0 ;
  assign WILL_FIRE_RL_doFADD_S = CAN_FIRE_RL_doFADD_S ;
  // rule RL_doFSUB_S
  assign CAN_FIRE_RL_doFSUB_S =
	     fpu$RDY_server_core_request_put && requestR[214] &&
	     stateR == 2'd1 &&
	     requestR[213:207] == 7'b1010011 &&
	     requestR[206:200] == 7'h04 ;
  assign WILL_FIRE_RL_doFSUB_S = CAN_FIRE_RL_doFSUB_S ;
  // rule RL_doFMUL_S
  assign CAN_FIRE_RL_doFMUL_S =
	     fpu$RDY_server_core_request_put && requestR[214] &&
	     stateR == 2'd1 &&
	     requestR[213:207] == 7'b1010011 &&
	     requestR[206:200] == 7'h08 ;
  assign WILL_FIRE_RL_doFMUL_S = CAN_FIRE_RL_doFMUL_S ;
  // rule RL_doFMADD_S
  assign CAN_FIRE_RL_doFMADD_S =
	     fpu$RDY_server_core_request_put && requestR[214] &&
	     stateR == 2'd1 &&
	     requestR[213:207] == 7'b1000011 &&
	     requestR_BITS_206_TO_200__q177[1:0] == 2'd0 ;
  assign WILL_FIRE_RL_doFMADD_S = CAN_FIRE_RL_doFMADD_S ;
  // rule RL_doFMSUB_S
  assign CAN_FIRE_RL_doFMSUB_S =
	     fpu$RDY_server_core_request_put && requestR[214] &&
	     stateR == 2'd1 &&
	     requestR[213:207] == 7'b1000111 &&
	     requestR_BITS_206_TO_200__q177[1:0] == 2'd0 ;
  assign WILL_FIRE_RL_doFMSUB_S = CAN_FIRE_RL_doFMSUB_S ;
  // rule RL_doFNMADD_S
  assign CAN_FIRE_RL_doFNMADD_S =
	     fpu$RDY_server_core_request_put && requestR[214] &&
	     stateR == 2'd1 &&
	     requestR[213:207] == 7'b1001111 &&
	     requestR_BITS_206_TO_200__q177[1:0] == 2'd0 ;
  assign WILL_FIRE_RL_doFNMADD_S = CAN_FIRE_RL_doFNMADD_S ;
  // rule RL_doFNMSUB_S
  assign CAN_FIRE_RL_doFNMSUB_S =
	     fpu$RDY_server_core_request_put && requestR[214] &&
	     stateR == 2'd1 &&
	     requestR[213:207] == 7'b1001011 &&
	     requestR_BITS_206_TO_200__q177[1:0] == 2'd0 ;
  assign WILL_FIRE_RL_doFNMSUB_S = CAN_FIRE_RL_doFNMSUB_S ;
  // rule RL_doFDIV_S
  assign CAN_FIRE_RL_doFDIV_S =
	     fpu$RDY_server_core_request_put && requestR[214] &&
	     stateR == 2'd1 &&
	     requestR[213:207] == 7'b1010011 &&
	     requestR[206:200] == 7'h0C ;
  assign WILL_FIRE_RL_doFDIV_S = CAN_FIRE_RL_doFDIV_S ;
  // rule RL_doFSQRT_S
  assign CAN_FIRE_RL_doFSQRT_S =
	     fpu$RDY_server_core_request_put && requestR[214] &&
	     stateR == 2'd1 &&
	     requestR[213:207] == 7'b1010011 &&
	     requestR[206:200] == 7'h2C ;
  assign WILL_FIRE_RL_doFSQRT_S = CAN_FIRE_RL_doFSQRT_S ;
  // rule RL_doFSGNJ_S
  assign CAN_FIRE_RL_doFSGNJ_S =
	     requestR[214] && stateR == 2'd1 &&
	     requestR[213:207] == 7'b1010011 &&
	     requestR[206:200] == 7'h10 &&
	     requestR[194:192] == 3'h0 ;
  assign WILL_FIRE_RL_doFSGNJ_S = CAN_FIRE_RL_doFSGNJ_S ;
  // rule RL_doFSGNJN_S
  assign CAN_FIRE_RL_doFSGNJN_S =
	     requestR[214] && stateR == 2'd1 &&
	     requestR[213:207] == 7'b1010011 &&
	     requestR[206:200] == 7'h10 &&
	     requestR[194:192] == 3'h1 ;
  assign WILL_FIRE_RL_doFSGNJN_S = CAN_FIRE_RL_doFSGNJN_S ;
  // rule RL_doFSGNJX_S
  assign CAN_FIRE_RL_doFSGNJX_S =
	     requestR[214] && stateR == 2'd1 &&
	     requestR[213:207] == 7'b1010011 &&
	     requestR[206:200] == 7'h10 &&
	     requestR[194:192] == 3'h2 ;
  assign WILL_FIRE_RL_doFSGNJX_S = CAN_FIRE_RL_doFSGNJX_S ;
  // rule RL_doFCVT_S_L
  assign CAN_FIRE_RL_doFCVT_S_L =
	     requestR[214] && stateR == 2'd1 &&
	     requestR[213:207] == 7'b1010011 &&
	     requestR[206:200] == 7'h68 &&
	     requestR[199:195] == 5'd2 ;
  assign WILL_FIRE_RL_doFCVT_S_L = CAN_FIRE_RL_doFCVT_S_L ;
  // rule RL_doFCVT_S_LU
  assign CAN_FIRE_RL_doFCVT_S_LU =
	     requestR[214] && stateR == 2'd1 &&
	     requestR[213:207] == 7'b1010011 &&
	     requestR[206:200] == 7'h68 &&
	     requestR[199:195] == 5'd3 ;
  assign WILL_FIRE_RL_doFCVT_S_LU = CAN_FIRE_RL_doFCVT_S_LU ;
  // rule RL_doFCVT_S_W
  assign CAN_FIRE_RL_doFCVT_S_W =
	     requestR[214] && stateR == 2'd1 &&
	     requestR[213:207] == 7'b1010011 &&
	     requestR[206:200] == 7'h68 &&
	     requestR[199:195] == 5'd0 ;
  assign WILL_FIRE_RL_doFCVT_S_W = CAN_FIRE_RL_doFCVT_S_W ;
  // rule RL_doFCVT_S_WU
  assign CAN_FIRE_RL_doFCVT_S_WU =
	     requestR[214] && stateR == 2'd1 &&
	     requestR[213:207] == 7'b1010011 &&
	     requestR[206:200] == 7'h68 &&
	     requestR[199:195] == 5'd1 ;
  assign WILL_FIRE_RL_doFCVT_S_WU = CAN_FIRE_RL_doFCVT_S_WU ;
  // rule RL_doFCVT_L_S
  assign CAN_FIRE_RL_doFCVT_L_S =
	     requestR[214] && stateR == 2'd1 &&
	     requestR[213:207] == 7'b1010011 &&
	     requestR[206:200] == 7'h60 &&
	     requestR[199:195] == 5'd2 ;
  assign WILL_FIRE_RL_doFCVT_L_S = CAN_FIRE_RL_doFCVT_L_S ;
  // rule RL_doFCVT_LU_S
  assign CAN_FIRE_RL_doFCVT_LU_S =
	     requestR[214] && stateR == 2'd1 &&
	     requestR[213:207] == 7'b1010011 &&
	     requestR[206:200] == 7'h60 &&
	     requestR[199:195] == 5'd3 ;
  assign WILL_FIRE_RL_doFCVT_LU_S = CAN_FIRE_RL_doFCVT_LU_S ;
  // rule RL_doFCVT_W_S
  assign CAN_FIRE_RL_doFCVT_W_S =
	     requestR[214] && stateR == 2'd1 &&
	     requestR[213:207] == 7'b1010011 &&
	     requestR[206:200] == 7'h60 &&
	     requestR[199:195] == 5'd0 ;
  assign WILL_FIRE_RL_doFCVT_W_S = CAN_FIRE_RL_doFCVT_W_S ;
  // rule RL_doFCVT_WU_S
  assign CAN_FIRE_RL_doFCVT_WU_S =
	     requestR[214] && stateR == 2'd1 &&
	     requestR[213:207] == 7'b1010011 &&
	     requestR[206:200] == 7'h60 &&
	     requestR[199:195] == 5'd1 ;
  assign WILL_FIRE_RL_doFCVT_WU_S = CAN_FIRE_RL_doFCVT_WU_S ;
  // rule RL_doFMIN_S
  assign CAN_FIRE_RL_doFMIN_S =
	     requestR[214] && stateR == 2'd1 &&
	     requestR[213:207] == 7'b1010011 &&
	     requestR[206:200] == 7'h14 &&
	     requestR[194:192] == 3'h0 ;
  assign WILL_FIRE_RL_doFMIN_S = CAN_FIRE_RL_doFMIN_S ;
  // rule RL_doFMAX_S
  assign CAN_FIRE_RL_doFMAX_S =
	     requestR[214] && stateR == 2'd1 &&
	     requestR[213:207] == 7'b1010011 &&
	     requestR[206:200] == 7'h14 &&
	     requestR[194:192] == 3'h1 ;
  assign WILL_FIRE_RL_doFMAX_S = CAN_FIRE_RL_doFMAX_S ;
  // rule RL_doFMV_W_X
  assign CAN_FIRE_RL_doFMV_W_X =
	     requestR[214] && stateR == 2'd1 &&
	     requestR[213:207] == 7'b1010011 &&
	     requestR[206:200] == 7'h78 &&
	     requestR[194:192] == 3'h0 ;
  assign WILL_FIRE_RL_doFMV_W_X = CAN_FIRE_RL_doFMV_W_X ;
  // rule RL_doFMV_X_W
  assign CAN_FIRE_RL_doFMV_X_W =
	     requestR[214] && stateR == 2'd1 &&
	     requestR[213:207] == 7'b1010011 &&
	     requestR[206:200] == 7'h70 &&
	     requestR[194:192] == 3'h0 ;
  assign WILL_FIRE_RL_doFMV_X_W = CAN_FIRE_RL_doFMV_X_W ;
  // rule RL_doFEQ_S
  assign CAN_FIRE_RL_doFEQ_S =
	     requestR[214] && stateR == 2'd1 &&
	     requestR[213:207] == 7'b1010011 &&
	     requestR[206:200] == 7'h50 &&
	     requestR[194:192] == 3'h2 ;
  assign WILL_FIRE_RL_doFEQ_S = CAN_FIRE_RL_doFEQ_S ;
  // rule RL_doFLT_S
  assign CAN_FIRE_RL_doFLT_S =
	     requestR[214] && stateR == 2'd1 &&
	     requestR[213:207] == 7'b1010011 &&
	     requestR[206:200] == 7'h50 &&
	     requestR[194:192] == 3'h1 ;
  assign WILL_FIRE_RL_doFLT_S = CAN_FIRE_RL_doFLT_S ;
  // rule RL_doFLE_S
  assign CAN_FIRE_RL_doFLE_S =
	     requestR[214] && stateR == 2'd1 &&
	     requestR[213:207] == 7'b1010011 &&
	     requestR[206:200] == 7'h50 &&
	     requestR[194:192] == 3'h0 ;
  assign WILL_FIRE_RL_doFLE_S = CAN_FIRE_RL_doFLE_S ;
  // rule RL_doFCLASS_S
  assign CAN_FIRE_RL_doFCLASS_S =
	     requestR[214] && stateR == 2'd1 &&
	     requestR[213:207] == 7'b1010011 &&
	     requestR[206:200] == 7'h70 &&
	     requestR[194:192] == 3'h1 ;
  assign WILL_FIRE_RL_doFCLASS_S = CAN_FIRE_RL_doFCLASS_S ;
  // rule RL_doFADD_D
  assign CAN_FIRE_RL_doFADD_D =
	     fpu$RDY_server_core_request_put && requestR[214] &&
	     stateR == 2'd1 &&
	     requestR[213:207] == 7'b1010011 &&
	     requestR[206:200] == 7'h01 ;
  assign WILL_FIRE_RL_doFADD_D = CAN_FIRE_RL_doFADD_D ;
  // rule RL_doFSUB_D
  assign CAN_FIRE_RL_doFSUB_D =
	     fpu$RDY_server_core_request_put && requestR[214] &&
	     stateR == 2'd1 &&
	     requestR[213:207] == 7'b1010011 &&
	     requestR[206:200] == 7'h05 ;
  assign WILL_FIRE_RL_doFSUB_D = CAN_FIRE_RL_doFSUB_D ;
  // rule RL_doFMUL_D
  assign CAN_FIRE_RL_doFMUL_D =
	     fpu$RDY_server_core_request_put && requestR[214] &&
	     stateR == 2'd1 &&
	     requestR[213:207] == 7'b1010011 &&
	     requestR[206:200] == 7'h09 ;
  assign WILL_FIRE_RL_doFMUL_D = CAN_FIRE_RL_doFMUL_D ;
  // rule RL_doFMADD_D
  assign CAN_FIRE_RL_doFMADD_D =
	     fpu$RDY_server_core_request_put && requestR[214] &&
	     stateR == 2'd1 &&
	     requestR[213:207] == 7'b1000011 &&
	     requestR_BITS_206_TO_200__q177[1:0] == 2'd1 ;
  assign WILL_FIRE_RL_doFMADD_D = CAN_FIRE_RL_doFMADD_D ;
  // rule RL_doFMSUB_D
  assign CAN_FIRE_RL_doFMSUB_D =
	     fpu$RDY_server_core_request_put && requestR[214] &&
	     stateR == 2'd1 &&
	     requestR[213:207] == 7'b1000111 &&
	     requestR_BITS_206_TO_200__q177[1:0] == 2'd1 ;
  assign WILL_FIRE_RL_doFMSUB_D = CAN_FIRE_RL_doFMSUB_D ;
  // rule RL_doFNMADD_D
  assign CAN_FIRE_RL_doFNMADD_D =
	     fpu$RDY_server_core_request_put && requestR[214] &&
	     stateR == 2'd1 &&
	     requestR[213:207] == 7'b1001111 &&
	     requestR_BITS_206_TO_200__q177[1:0] == 2'd1 ;
  assign WILL_FIRE_RL_doFNMADD_D = CAN_FIRE_RL_doFNMADD_D ;
  // rule RL_doFNMSUB_D
  assign CAN_FIRE_RL_doFNMSUB_D =
	     fpu$RDY_server_core_request_put && requestR[214] &&
	     stateR == 2'd1 &&
	     requestR[213:207] == 7'b1001011 &&
	     requestR_BITS_206_TO_200__q177[1:0] == 2'd1 ;
  assign WILL_FIRE_RL_doFNMSUB_D = CAN_FIRE_RL_doFNMSUB_D ;
  // rule RL_doFDIV_D
  assign CAN_FIRE_RL_doFDIV_D =
	     fpu$RDY_server_core_request_put && requestR[214] &&
	     stateR == 2'd1 &&
	     requestR[213:207] == 7'b1010011 &&
	     requestR[206:200] == 7'h0D ;
  assign WILL_FIRE_RL_doFDIV_D = CAN_FIRE_RL_doFDIV_D ;
  // rule RL_doFSQRT_D
  assign CAN_FIRE_RL_doFSQRT_D =
	     fpu$RDY_server_core_request_put && requestR[214] &&
	     stateR == 2'd1 &&
	     requestR[213:207] == 7'b1010011 &&
	     requestR[206:200] == 7'h2D ;
  assign WILL_FIRE_RL_doFSQRT_D = CAN_FIRE_RL_doFSQRT_D ;
  // rule RL_doFSGNJ_D
  assign CAN_FIRE_RL_doFSGNJ_D =
	     requestR[214] && stateR == 2'd1 &&
	     requestR[213:207] == 7'b1010011 &&
	     requestR[206:200] == 7'h11 &&
	     requestR[194:192] == 3'h0 ;
  assign WILL_FIRE_RL_doFSGNJ_D = CAN_FIRE_RL_doFSGNJ_D ;
  // rule RL_doFSGNJN_D
  assign CAN_FIRE_RL_doFSGNJN_D =
	     requestR[214] && stateR == 2'd1 &&
	     requestR[213:207] == 7'b1010011 &&
	     requestR[206:200] == 7'h11 &&
	     requestR[194:192] == 3'h1 ;
  assign WILL_FIRE_RL_doFSGNJN_D = CAN_FIRE_RL_doFSGNJN_D ;
  // rule RL_doFSGNJX_D
  assign CAN_FIRE_RL_doFSGNJX_D =
	     requestR[214] && stateR == 2'd1 &&
	     requestR[213:207] == 7'b1010011 &&
	     requestR[206:200] == 7'h11 &&
	     requestR[194:192] == 3'h2 ;
  assign WILL_FIRE_RL_doFSGNJX_D = CAN_FIRE_RL_doFSGNJX_D ;
  // rule RL_doFCVT_D_W
  assign CAN_FIRE_RL_doFCVT_D_W =
	     requestR[214] && stateR == 2'd1 &&
	     requestR[213:207] == 7'b1010011 &&
	     requestR[206:200] == 7'h69 &&
	     requestR[199:195] == 5'd0 ;
  assign WILL_FIRE_RL_doFCVT_D_W = CAN_FIRE_RL_doFCVT_D_W ;
  // rule RL_doFCVT_D_WU
  assign CAN_FIRE_RL_doFCVT_D_WU =
	     requestR[214] && stateR == 2'd1 &&
	     requestR[213:207] == 7'b1010011 &&
	     requestR[206:200] == 7'h69 &&
	     requestR[199:195] == 5'd1 ;
  assign WILL_FIRE_RL_doFCVT_D_WU = CAN_FIRE_RL_doFCVT_D_WU ;
  // rule RL_doFCVT_W_D
  assign CAN_FIRE_RL_doFCVT_W_D =
	     requestR[214] && stateR == 2'd1 &&
	     requestR[213:207] == 7'b1010011 &&
	     requestR[206:200] == 7'h61 &&
	     requestR[199:195] == 5'd0 ;
  assign WILL_FIRE_RL_doFCVT_W_D = CAN_FIRE_RL_doFCVT_W_D ;
  // rule RL_doFCVT_WU_D
  assign CAN_FIRE_RL_doFCVT_WU_D =
	     requestR[214] && stateR == 2'd1 &&
	     requestR[213:207] == 7'b1010011 &&
	     requestR[206:200] == 7'h61 &&
	     requestR[199:195] == 5'd1 ;
  assign WILL_FIRE_RL_doFCVT_WU_D = CAN_FIRE_RL_doFCVT_WU_D ;
  // rule RL_doFCVT_D_L
  assign CAN_FIRE_RL_doFCVT_D_L =
	     requestR[214] && stateR == 2'd1 &&
	     requestR[213:207] == 7'b1010011 &&
	     requestR[206:200] == 7'h69 &&
	     requestR[199:195] == 5'd2 ;
  assign WILL_FIRE_RL_doFCVT_D_L = CAN_FIRE_RL_doFCVT_D_L ;
  // rule RL_doFCVT_D_LU
  assign CAN_FIRE_RL_doFCVT_D_LU =
	     requestR[214] && stateR == 2'd1 &&
	     requestR[213:207] == 7'b1010011 &&
	     requestR[206:200] == 7'h69 &&
	     requestR[199:195] == 5'd3 ;
  assign WILL_FIRE_RL_doFCVT_D_LU = CAN_FIRE_RL_doFCVT_D_LU ;
  // rule RL_doFCVT_L_D
  assign CAN_FIRE_RL_doFCVT_L_D =
	     requestR[214] && stateR == 2'd1 &&
	     requestR[213:207] == 7'b1010011 &&
	     requestR[206:200] == 7'h61 &&
	     requestR[199:195] == 5'd2 ;
  assign WILL_FIRE_RL_doFCVT_L_D = CAN_FIRE_RL_doFCVT_L_D ;
  // rule RL_doFCVT_LU_D
  assign CAN_FIRE_RL_doFCVT_LU_D =
	     requestR[214] && stateR == 2'd1 &&
	     requestR[213:207] == 7'b1010011 &&
	     requestR[206:200] == 7'h61 &&
	     requestR[199:195] == 5'd3 ;
  assign WILL_FIRE_RL_doFCVT_LU_D = CAN_FIRE_RL_doFCVT_LU_D ;
  // rule RL_doFCVT_S_D
  assign CAN_FIRE_RL_doFCVT_S_D =
	     requestR[214] && stateR == 2'd1 &&
	     requestR[213:207] == 7'b1010011 &&
	     requestR[206:200] == 7'h20 &&
	     requestR[199:195] == 5'd1 ;
  assign WILL_FIRE_RL_doFCVT_S_D = CAN_FIRE_RL_doFCVT_S_D ;
  // rule RL_doFCVT_D_S
  assign CAN_FIRE_RL_doFCVT_D_S =
	     requestR[214] && stateR == 2'd1 &&
	     requestR[213:207] == 7'b1010011 &&
	     requestR[206:200] == 7'h21 &&
	     requestR[199:195] == 5'd0 ;
  assign WILL_FIRE_RL_doFCVT_D_S = CAN_FIRE_RL_doFCVT_D_S ;
  // rule RL_doFMIN_D
  assign CAN_FIRE_RL_doFMIN_D =
	     requestR[214] && stateR == 2'd1 &&
	     requestR[213:207] == 7'b1010011 &&
	     requestR[206:200] == 7'h15 &&
	     requestR[194:192] == 3'h0 ;
  assign WILL_FIRE_RL_doFMIN_D = CAN_FIRE_RL_doFMIN_D ;
  // rule RL_doFMAX_D
  assign CAN_FIRE_RL_doFMAX_D =
	     requestR[214] && stateR == 2'd1 &&
	     requestR[213:207] == 7'b1010011 &&
	     requestR[206:200] == 7'h15 &&
	     requestR[194:192] == 3'h1 ;
  assign WILL_FIRE_RL_doFMAX_D = CAN_FIRE_RL_doFMAX_D ;
  // rule RL_doFEQ_D
  assign CAN_FIRE_RL_doFEQ_D =
	     requestR[214] && stateR == 2'd1 &&
	     requestR[213:207] == 7'b1010011 &&
	     requestR[206:200] == 7'h51 &&
	     requestR[194:192] == 3'h2 ;
  assign WILL_FIRE_RL_doFEQ_D = CAN_FIRE_RL_doFEQ_D ;
  // rule RL_doFLT_D
  assign CAN_FIRE_RL_doFLT_D =
	     requestR[214] && stateR == 2'd1 &&
	     requestR[213:207] == 7'b1010011 &&
	     requestR[206:200] == 7'h51 &&
	     requestR[194:192] == 3'h1 ;
  assign WILL_FIRE_RL_doFLT_D = CAN_FIRE_RL_doFLT_D ;
  // rule RL_doFLE_D
  assign CAN_FIRE_RL_doFLE_D =
	     requestR[214] && stateR == 2'd1 &&
	     requestR[213:207] == 7'b1010011 &&
	     requestR[206:200] == 7'h51 &&
	     requestR[194:192] == 3'h0 ;
  assign WILL_FIRE_RL_doFLE_D = CAN_FIRE_RL_doFLE_D ;
  // rule RL_doFMV_D_X
  assign CAN_FIRE_RL_doFMV_D_X =
	     requestR[214] && stateR == 2'd1 &&
	     requestR[213:207] == 7'b1010011 &&
	     requestR[206:200] == 7'h79 &&
	     requestR[194:192] == 3'h0 ;
  assign WILL_FIRE_RL_doFMV_D_X = CAN_FIRE_RL_doFMV_D_X ;
  // rule RL_doFMV_X_D
  assign CAN_FIRE_RL_doFMV_X_D =
	     requestR[214] && stateR == 2'd1 &&
	     requestR[213:207] == 7'b1010011 &&
	     requestR[206:200] == 7'h71 &&
	     requestR[194:192] == 3'h0 ;
  assign WILL_FIRE_RL_doFMV_X_D = CAN_FIRE_RL_doFMV_X_D ;
  // rule RL_doFCLASS_D
  assign CAN_FIRE_RL_doFCLASS_D =
	     requestR[214] && stateR == 2'd1 &&
	     requestR[213:207] == 7'b1010011 &&
	     requestR[206:200] == 7'h71 &&
	     requestR[194:192] == 3'h1 ;
  assign WILL_FIRE_RL_doFCLASS_D = CAN_FIRE_RL_doFCLASS_D ;
  // rule RL_rl_get_fpu_result
  assign CAN_FIRE_RL_rl_get_fpu_result = MUX_dw_result$wset_1__SEL_1 ;
  assign WILL_FIRE_RL_rl_get_fpu_result = MUX_dw_result$wset_1__SEL_1 ;
  // rule RL_rl_drive_fpu_result
  assign CAN_FIRE_RL_rl_drive_fpu_result = stateR == 2'd3 ;
  assign WILL_FIRE_RL_rl_drive_fpu_result = stateR == 2'd3 ;
  // rule RL_rl_reset_begin
  assign CAN_FIRE_RL_rl_reset_begin =
	     fpu$RDY_server_reset_request_put && resetReqsF$EMPTY_N ;
  assign WILL_FIRE_RL_rl_reset_begin = CAN_FIRE_RL_rl_reset_begin ;
  // inputs to muxes for submodule ports
  assign MUX_dw_result$wset_1__SEL_1 =
	     fpu$RDY_server_core_response_get && stateR == 2'd2 ;
  assign MUX_dw_result$wset_1__VAL_1 =
	     { x__h230460, fpu$server_core_response_get[4:0] } ;
  assign MUX_fpu$server_core_request_put_1__VAL_1 =
	     { 33'h1AAAAAAAA,
	       requestR_BITS_191_TO_128__q1[63:32] == 32'hFFFFFFFF &&
	       requestR_BITS_191_TO_128__q1[31],
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d37,
	       33'h1AAAAAAAA,
	       IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d48,
	       65'h0AAAAAAAAAAAAAAAA,
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d61,
	       4'd0 } ;
  assign MUX_fpu$server_core_request_put_1__VAL_2 =
	     { 33'h1AAAAAAAA,
	       requestR_BITS_191_TO_128__q1[63:32] == 32'hFFFFFFFF &&
	       requestR_BITS_191_TO_128__q1[31],
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d37,
	       33'h1AAAAAAAA,
	       IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d48,
	       65'h0AAAAAAAAAAAAAAAA,
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d61,
	       4'd1 } ;
  assign MUX_fpu$server_core_request_put_1__VAL_3 =
	     { 33'h1AAAAAAAA,
	       requestR_BITS_191_TO_128__q1[63:32] == 32'hFFFFFFFF &&
	       requestR_BITS_191_TO_128__q1[31],
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d37,
	       33'h1AAAAAAAA,
	       IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d48,
	       65'h0AAAAAAAAAAAAAAAA,
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d61,
	       4'd2 } ;
  assign MUX_fpu$server_core_request_put_1__VAL_4 =
	     { 33'h1AAAAAAAA,
	       requestR_BITS_191_TO_128__q1[63:32] == 32'hFFFFFFFF &&
	       requestR_BITS_191_TO_128__q1[31],
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d37,
	       33'h1AAAAAAAA,
	       IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d48,
	       _1_CONCAT_DONTCARE_CONCAT_IF_requestR_3_BIT_214_ETC___d97,
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d61,
	       4'd5 } ;
  assign MUX_fpu$server_core_request_put_1__VAL_5 =
	     { 33'h1AAAAAAAA,
	       requestR_BITS_191_TO_128__q1[63:32] == 32'hFFFFFFFF &&
	       requestR_BITS_191_TO_128__q1[31],
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d37,
	       33'h1AAAAAAAA,
	       IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d48,
	       _1_CONCAT_DONTCARE_CONCAT_IF_requestR_3_BIT_214_ETC___d97,
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d61,
	       4'd6 } ;
  assign MUX_fpu$server_core_request_put_1__VAL_6 =
	     { 33'h1AAAAAAAA,
	       requestR_BITS_191_TO_128__q1[63:32] == 32'hFFFFFFFF &&
	       requestR_BITS_191_TO_128__q1[31],
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d37,
	       33'h1AAAAAAAA,
	       IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d48,
	       _1_CONCAT_DONTCARE_CONCAT_IF_requestR_3_BIT_214_ETC___d97,
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d61,
	       4'd7 } ;
  assign MUX_fpu$server_core_request_put_1__VAL_7 =
	     { 33'h1AAAAAAAA,
	       requestR_BITS_191_TO_128__q1[63:32] == 32'hFFFFFFFF &&
	       requestR_BITS_191_TO_128__q1[31],
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d37,
	       33'h1AAAAAAAA,
	       IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d48,
	       _1_CONCAT_DONTCARE_CONCAT_IF_requestR_3_BIT_214_ETC___d97,
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d61,
	       4'd8 } ;
  assign MUX_fpu$server_core_request_put_1__VAL_8 =
	     { 33'h1AAAAAAAA,
	       requestR_BITS_191_TO_128__q1[63:32] == 32'hFFFFFFFF &&
	       requestR_BITS_191_TO_128__q1[31],
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d37,
	       33'h1AAAAAAAA,
	       IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d48,
	       65'h0AAAAAAAAAAAAAAAA,
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d61,
	       4'd3 } ;
  assign MUX_fpu$server_core_request_put_1__VAL_9 =
	     { 33'h1AAAAAAAA,
	       requestR_BITS_191_TO_128__q1[63:32] == 32'hFFFFFFFF &&
	       requestR_BITS_191_TO_128__q1[31],
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d37,
	       130'h15555555555555554AAAAAAAAAAAAAAAA,
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d61,
	       4'd4 } ;
  assign MUX_fpu$server_core_request_put_1__VAL_10 =
	     { 1'd0,
	       requestR[191:128],
	       1'd0,
	       requestR[127:64],
	       65'h0AAAAAAAAAAAAAAAA,
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d61,
	       4'd0 } ;
  assign MUX_fpu$server_core_request_put_1__VAL_11 =
	     { 1'd0,
	       requestR[191:128],
	       1'd0,
	       requestR[127:64],
	       65'h0AAAAAAAAAAAAAAAA,
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d61,
	       4'd1 } ;
  assign MUX_fpu$server_core_request_put_1__VAL_12 =
	     { 1'd0,
	       requestR[191:128],
	       1'd0,
	       requestR[127:64],
	       65'h0AAAAAAAAAAAAAAAA,
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d61,
	       4'd2 } ;
  assign MUX_fpu$server_core_request_put_1__VAL_13 =
	     { 1'd0,
	       requestR[191:128],
	       1'd0,
	       requestR[127:64],
	       1'd0,
	       requestR[63:0],
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d61,
	       4'd5 } ;
  assign MUX_fpu$server_core_request_put_1__VAL_14 =
	     { 1'd0,
	       requestR[191:128],
	       1'd0,
	       requestR[127:64],
	       1'd0,
	       requestR[63:0],
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d61,
	       4'd6 } ;
  assign MUX_fpu$server_core_request_put_1__VAL_15 =
	     { 1'd0,
	       requestR[191:128],
	       1'd0,
	       requestR[127:64],
	       1'd0,
	       requestR[63:0],
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d61,
	       4'd7 } ;
  assign MUX_fpu$server_core_request_put_1__VAL_16 =
	     { 1'd0,
	       requestR[191:128],
	       1'd0,
	       requestR[127:64],
	       1'd0,
	       requestR[63:0],
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d61,
	       4'd8 } ;
  assign MUX_fpu$server_core_request_put_1__VAL_17 =
	     { 1'd0,
	       requestR[191:128],
	       1'd0,
	       requestR[127:64],
	       65'h0AAAAAAAAAAAAAAAA,
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d61,
	       4'd3 } ;
  assign MUX_fpu$server_core_request_put_1__VAL_18 =
	     { 1'd0,
	       requestR[191:128],
	       130'h15555555555555554AAAAAAAAAAAAAAAA,
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d61,
	       4'd4 } ;
  assign MUX_requestR$write_1__VAL_2 =
	     { 1'd1,
	       req_opcode,
	       req_f7,
	       req_rs2,
	       req_rm,
	       req_v1,
	       req_v2,
	       req_v3 } ;
  assign MUX_resultR$write_1__VAL_3 =
	     { 1'd1, x__h230460, fpu$server_core_response_get[4:0] } ;
  assign MUX_resultR$write_1__VAL_4 = { 1'd1, x__h229846, 5'd0 } ;
  assign MUX_resultR$write_1__VAL_6 = { 1'd1, requestR[191:128], 5'd0 } ;
  assign MUX_resultR$write_1__VAL_7 = { 1'd1, x__h227602, x__h227382 } ;
  assign MUX_resultR$write_1__VAL_8 = { 1'd1, x__h225685, x__h227382 } ;
  assign MUX_resultR$write_1__VAL_9 = { 1'd1, x__h222950, x__h217430 } ;
  assign MUX_resultR$write_1__VAL_10 = { 1'd1, x__h218468, x__h217430 } ;
  assign MUX_resultR$write_1__VAL_11 = { 1'd1, x__h213882, x__h217430 } ;
  assign MUX_resultR$write_1__VAL_12 = { 1'd1, x__h167888, x__h212920 } ;
  assign MUX_resultR$write_1__VAL_13 = { 1'd1, x__h113022, x__h166866 } ;
  assign MUX_resultR$write_1__VAL_14 = { 1'd1, x__h112240, x__h112739 } ;
  assign MUX_resultR$write_1__VAL_15 = { 1'd1, x__h110179, x__h111943 } ;
  assign MUX_resultR$write_1__VAL_16 = { 1'd1, x__h97683, x__h109855 } ;
  assign MUX_resultR$write_1__VAL_17 = { 1'd1, x__h84681, x__h97358 } ;
  assign MUX_resultR$write_1__VAL_18 = { 1'd1, x__h83895, x__h84397 } ;
  assign MUX_resultR$write_1__VAL_19 = { 1'd1, x__h82279, x__h83598 } ;
  assign MUX_resultR$write_1__VAL_20 = { 1'd1, x__h71361, x__h81955 } ;
  assign MUX_resultR$write_1__VAL_21 = { 1'd1, x__h60162, x__h71036 } ;
  assign MUX_resultR$write_1__VAL_22 = { 1'd1, x__h59992, 5'd0 } ;
  assign MUX_resultR$write_1__VAL_23 = { 1'd1, x__h59829, 5'd0 } ;
  assign MUX_resultR$write_1__VAL_24 = { 1'd1, x__h59668, 5'd0 } ;
  assign MUX_resultR$write_1__VAL_25 = { 1'd1, x__h57514, 5'd0 } ;
  assign MUX_resultR$write_1__VAL_26 = { 1'd1, x__h56389, x__h56169 } ;
  assign MUX_resultR$write_1__VAL_27 = { 1'd1, x__h55280, x__h56169 } ;
  assign MUX_resultR$write_1__VAL_28 = { 1'd1, x__h53757, x__h50220 } ;
  assign MUX_resultR$write_1__VAL_29 = { 1'd1, x__h53579, 5'd0 } ;
  assign MUX_resultR$write_1__VAL_30 = { 1'd1, x__h53419, 5'd0 } ;
  assign MUX_resultR$write_1__VAL_31 = { 1'd1, x__h50854, x__h50220 } ;
  assign MUX_resultR$write_1__VAL_32 = { 1'd1, x__h48180, x__h50220 } ;
  assign MUX_resultR$write_1__VAL_33 = { 1'd1, x__h47391, x__h47893 } ;
  assign MUX_resultR$write_1__VAL_34 = { 1'd1, x__h45775, x__h47094 } ;
  assign MUX_resultR$write_1__VAL_35 = { 1'd1, x__h44993, x__h45492 } ;
  assign MUX_resultR$write_1__VAL_36 = { 1'd1, x__h42915, x__h44696 } ;
  assign MUX_resultR$write_1__VAL_37 = { 1'd1, x__h36028, x__h42591 } ;
  assign MUX_resultR$write_1__VAL_38 = { 1'd1, x__h28828, x__h35703 } ;
  assign MUX_resultR$write_1__VAL_39 = { 1'd1, x__h16727, x__h28503 } ;
  assign MUX_resultR$write_1__VAL_40 = { 1'd1, res__h3932, fcsr__h3933 } ;
  assign MUX_resultR$write_1__VAL_41 = { 1'd1, x__h3778, 5'd0 } ;
  assign MUX_resultR$write_1__VAL_42 = { 1'd1, x__h3605, 5'd0 } ;
  assign MUX_resultR$write_1__VAL_43 = { 1'd1, x__h3429, 5'd0 } ;
  // inlined wires
  assign dw_valid$wget = !WILL_FIRE_RL_rl_drive_fpu_result || resultR[69] ;
  assign dw_valid$whas =
	     WILL_FIRE_RL_rl_drive_fpu_result ||
	     WILL_FIRE_RL_rl_get_fpu_result ;
  assign dw_result$wget =
	     WILL_FIRE_RL_rl_get_fpu_result ?
	       MUX_dw_result$wset_1__VAL_1 :
	       resultR[68:0] ;
  // register requestR
  assign requestR$D_IN =
	     WILL_FIRE_RL_rl_reset_begin ?
	       215'h2AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA :
	       MUX_requestR$write_1__VAL_2 ;
  assign requestR$EN = WILL_FIRE_RL_rl_reset_begin || EN_req ;
  // register resultR
  always@(WILL_FIRE_RL_rl_reset_begin or
	  EN_req or
	  WILL_FIRE_RL_rl_get_fpu_result or
	  MUX_resultR$write_1__VAL_3 or
	  WILL_FIRE_RL_doFCLASS_D or
	  MUX_resultR$write_1__VAL_4 or
	  WILL_FIRE_RL_doFMV_X_D or
	  MUX_resultR$write_1__VAL_6 or
	  WILL_FIRE_RL_doFMV_D_X or
	  WILL_FIRE_RL_doFLE_D or
	  MUX_resultR$write_1__VAL_7 or
	  WILL_FIRE_RL_doFLT_D or
	  MUX_resultR$write_1__VAL_8 or
	  WILL_FIRE_RL_doFEQ_D or
	  MUX_resultR$write_1__VAL_9 or
	  WILL_FIRE_RL_doFMAX_D or
	  MUX_resultR$write_1__VAL_10 or
	  WILL_FIRE_RL_doFMIN_D or
	  MUX_resultR$write_1__VAL_11 or
	  WILL_FIRE_RL_doFCVT_D_S or
	  MUX_resultR$write_1__VAL_12 or
	  WILL_FIRE_RL_doFCVT_S_D or
	  MUX_resultR$write_1__VAL_13 or
	  WILL_FIRE_RL_doFCVT_LU_D or
	  MUX_resultR$write_1__VAL_14 or
	  WILL_FIRE_RL_doFCVT_L_D or
	  MUX_resultR$write_1__VAL_15 or
	  WILL_FIRE_RL_doFCVT_D_LU or
	  MUX_resultR$write_1__VAL_16 or
	  WILL_FIRE_RL_doFCVT_D_L or
	  MUX_resultR$write_1__VAL_17 or
	  WILL_FIRE_RL_doFCVT_WU_D or
	  MUX_resultR$write_1__VAL_18 or
	  WILL_FIRE_RL_doFCVT_W_D or
	  MUX_resultR$write_1__VAL_19 or
	  WILL_FIRE_RL_doFCVT_D_WU or
	  MUX_resultR$write_1__VAL_20 or
	  WILL_FIRE_RL_doFCVT_D_W or
	  MUX_resultR$write_1__VAL_21 or
	  WILL_FIRE_RL_doFSGNJX_D or
	  MUX_resultR$write_1__VAL_22 or
	  WILL_FIRE_RL_doFSGNJN_D or
	  MUX_resultR$write_1__VAL_23 or
	  WILL_FIRE_RL_doFSGNJ_D or
	  MUX_resultR$write_1__VAL_24 or
	  WILL_FIRE_RL_doFCLASS_S or
	  MUX_resultR$write_1__VAL_25 or
	  WILL_FIRE_RL_doFLE_S or
	  MUX_resultR$write_1__VAL_26 or
	  WILL_FIRE_RL_doFLT_S or
	  MUX_resultR$write_1__VAL_27 or
	  WILL_FIRE_RL_doFEQ_S or
	  MUX_resultR$write_1__VAL_28 or
	  WILL_FIRE_RL_doFMV_X_W or
	  MUX_resultR$write_1__VAL_29 or
	  WILL_FIRE_RL_doFMV_W_X or
	  MUX_resultR$write_1__VAL_30 or
	  WILL_FIRE_RL_doFMAX_S or
	  MUX_resultR$write_1__VAL_31 or
	  WILL_FIRE_RL_doFMIN_S or
	  MUX_resultR$write_1__VAL_32 or
	  WILL_FIRE_RL_doFCVT_WU_S or
	  MUX_resultR$write_1__VAL_33 or
	  WILL_FIRE_RL_doFCVT_W_S or
	  MUX_resultR$write_1__VAL_34 or
	  WILL_FIRE_RL_doFCVT_LU_S or
	  MUX_resultR$write_1__VAL_35 or
	  WILL_FIRE_RL_doFCVT_L_S or
	  MUX_resultR$write_1__VAL_36 or
	  WILL_FIRE_RL_doFCVT_S_WU or
	  MUX_resultR$write_1__VAL_37 or
	  WILL_FIRE_RL_doFCVT_S_W or
	  MUX_resultR$write_1__VAL_38 or
	  WILL_FIRE_RL_doFCVT_S_LU or
	  MUX_resultR$write_1__VAL_39 or
	  WILL_FIRE_RL_doFCVT_S_L or
	  MUX_resultR$write_1__VAL_40 or
	  WILL_FIRE_RL_doFSGNJX_S or
	  MUX_resultR$write_1__VAL_41 or
	  WILL_FIRE_RL_doFSGNJN_S or
	  MUX_resultR$write_1__VAL_42 or
	  WILL_FIRE_RL_doFSGNJ_S or MUX_resultR$write_1__VAL_43)
  case (1'b1)
    WILL_FIRE_RL_rl_reset_begin || EN_req:
	resultR$D_IN = 70'h0AAAAAAAAAAAAAAAAA;
    WILL_FIRE_RL_rl_get_fpu_result: resultR$D_IN = MUX_resultR$write_1__VAL_3;
    WILL_FIRE_RL_doFCLASS_D: resultR$D_IN = MUX_resultR$write_1__VAL_4;
    WILL_FIRE_RL_doFMV_X_D: resultR$D_IN = MUX_resultR$write_1__VAL_6;
    WILL_FIRE_RL_doFMV_D_X: resultR$D_IN = MUX_resultR$write_1__VAL_6;
    WILL_FIRE_RL_doFLE_D: resultR$D_IN = MUX_resultR$write_1__VAL_7;
    WILL_FIRE_RL_doFLT_D: resultR$D_IN = MUX_resultR$write_1__VAL_8;
    WILL_FIRE_RL_doFEQ_D: resultR$D_IN = MUX_resultR$write_1__VAL_9;
    WILL_FIRE_RL_doFMAX_D: resultR$D_IN = MUX_resultR$write_1__VAL_10;
    WILL_FIRE_RL_doFMIN_D: resultR$D_IN = MUX_resultR$write_1__VAL_11;
    WILL_FIRE_RL_doFCVT_D_S: resultR$D_IN = MUX_resultR$write_1__VAL_12;
    WILL_FIRE_RL_doFCVT_S_D: resultR$D_IN = MUX_resultR$write_1__VAL_13;
    WILL_FIRE_RL_doFCVT_LU_D: resultR$D_IN = MUX_resultR$write_1__VAL_14;
    WILL_FIRE_RL_doFCVT_L_D: resultR$D_IN = MUX_resultR$write_1__VAL_15;
    WILL_FIRE_RL_doFCVT_D_LU: resultR$D_IN = MUX_resultR$write_1__VAL_16;
    WILL_FIRE_RL_doFCVT_D_L: resultR$D_IN = MUX_resultR$write_1__VAL_17;
    WILL_FIRE_RL_doFCVT_WU_D: resultR$D_IN = MUX_resultR$write_1__VAL_18;
    WILL_FIRE_RL_doFCVT_W_D: resultR$D_IN = MUX_resultR$write_1__VAL_19;
    WILL_FIRE_RL_doFCVT_D_WU: resultR$D_IN = MUX_resultR$write_1__VAL_20;
    WILL_FIRE_RL_doFCVT_D_W: resultR$D_IN = MUX_resultR$write_1__VAL_21;
    WILL_FIRE_RL_doFSGNJX_D: resultR$D_IN = MUX_resultR$write_1__VAL_22;
    WILL_FIRE_RL_doFSGNJN_D: resultR$D_IN = MUX_resultR$write_1__VAL_23;
    WILL_FIRE_RL_doFSGNJ_D: resultR$D_IN = MUX_resultR$write_1__VAL_24;
    WILL_FIRE_RL_doFCLASS_S: resultR$D_IN = MUX_resultR$write_1__VAL_25;
    WILL_FIRE_RL_doFLE_S: resultR$D_IN = MUX_resultR$write_1__VAL_26;
    WILL_FIRE_RL_doFLT_S: resultR$D_IN = MUX_resultR$write_1__VAL_27;
    WILL_FIRE_RL_doFEQ_S: resultR$D_IN = MUX_resultR$write_1__VAL_28;
    WILL_FIRE_RL_doFMV_X_W: resultR$D_IN = MUX_resultR$write_1__VAL_29;
    WILL_FIRE_RL_doFMV_W_X: resultR$D_IN = MUX_resultR$write_1__VAL_30;
    WILL_FIRE_RL_doFMAX_S: resultR$D_IN = MUX_resultR$write_1__VAL_31;
    WILL_FIRE_RL_doFMIN_S: resultR$D_IN = MUX_resultR$write_1__VAL_32;
    WILL_FIRE_RL_doFCVT_WU_S: resultR$D_IN = MUX_resultR$write_1__VAL_33;
    WILL_FIRE_RL_doFCVT_W_S: resultR$D_IN = MUX_resultR$write_1__VAL_34;
    WILL_FIRE_RL_doFCVT_LU_S: resultR$D_IN = MUX_resultR$write_1__VAL_35;
    WILL_FIRE_RL_doFCVT_L_S: resultR$D_IN = MUX_resultR$write_1__VAL_36;
    WILL_FIRE_RL_doFCVT_S_WU: resultR$D_IN = MUX_resultR$write_1__VAL_37;
    WILL_FIRE_RL_doFCVT_S_W: resultR$D_IN = MUX_resultR$write_1__VAL_38;
    WILL_FIRE_RL_doFCVT_S_LU: resultR$D_IN = MUX_resultR$write_1__VAL_39;
    WILL_FIRE_RL_doFCVT_S_L: resultR$D_IN = MUX_resultR$write_1__VAL_40;
    WILL_FIRE_RL_doFSGNJX_S: resultR$D_IN = MUX_resultR$write_1__VAL_41;
    WILL_FIRE_RL_doFSGNJN_S: resultR$D_IN = MUX_resultR$write_1__VAL_42;
    WILL_FIRE_RL_doFSGNJ_S: resultR$D_IN = MUX_resultR$write_1__VAL_43;
    default: resultR$D_IN = 70'h2AAAAAAAAAAAAAAAAA /* unspecified value */ ;
  endcase
  assign resultR$EN =
	     WILL_FIRE_RL_rl_reset_begin || EN_req ||
	     WILL_FIRE_RL_doFMV_X_D ||
	     WILL_FIRE_RL_doFMV_D_X ||
	     WILL_FIRE_RL_doFSGNJ_S ||
	     WILL_FIRE_RL_doFSGNJN_S ||
	     WILL_FIRE_RL_doFSGNJX_S ||
	     WILL_FIRE_RL_doFCVT_S_L ||
	     WILL_FIRE_RL_doFCVT_S_LU ||
	     WILL_FIRE_RL_doFCVT_S_W ||
	     WILL_FIRE_RL_doFCVT_S_WU ||
	     WILL_FIRE_RL_doFCVT_L_S ||
	     WILL_FIRE_RL_doFCVT_LU_S ||
	     WILL_FIRE_RL_doFCVT_W_S ||
	     WILL_FIRE_RL_doFCVT_WU_S ||
	     WILL_FIRE_RL_doFMIN_S ||
	     WILL_FIRE_RL_doFMAX_S ||
	     WILL_FIRE_RL_doFMV_W_X ||
	     WILL_FIRE_RL_doFMV_X_W ||
	     WILL_FIRE_RL_doFEQ_S ||
	     WILL_FIRE_RL_doFLT_S ||
	     WILL_FIRE_RL_doFLE_S ||
	     WILL_FIRE_RL_doFCLASS_S ||
	     WILL_FIRE_RL_doFSGNJ_D ||
	     WILL_FIRE_RL_doFSGNJN_D ||
	     WILL_FIRE_RL_doFSGNJX_D ||
	     WILL_FIRE_RL_doFCVT_D_W ||
	     WILL_FIRE_RL_doFCVT_D_WU ||
	     WILL_FIRE_RL_doFCVT_W_D ||
	     WILL_FIRE_RL_doFCVT_WU_D ||
	     WILL_FIRE_RL_doFCVT_D_L ||
	     WILL_FIRE_RL_doFCVT_D_LU ||
	     WILL_FIRE_RL_doFCVT_L_D ||
	     WILL_FIRE_RL_doFCVT_LU_D ||
	     WILL_FIRE_RL_doFCVT_S_D ||
	     WILL_FIRE_RL_doFCVT_D_S ||
	     WILL_FIRE_RL_doFMIN_D ||
	     WILL_FIRE_RL_doFMAX_D ||
	     WILL_FIRE_RL_doFEQ_D ||
	     WILL_FIRE_RL_doFLT_D ||
	     WILL_FIRE_RL_doFLE_D ||
	     WILL_FIRE_RL_doFCLASS_D ||
	     WILL_FIRE_RL_rl_get_fpu_result ;
  // register stateR
  always@(WILL_FIRE_RL_rl_reset_begin or
	  EN_req or
	  WILL_FIRE_RL_rl_get_fpu_result or
	  WILL_FIRE_RL_doFCLASS_D or
	  WILL_FIRE_RL_doFMV_X_D or
	  WILL_FIRE_RL_doFMV_D_X or
	  WILL_FIRE_RL_doFLE_D or
	  WILL_FIRE_RL_doFLT_D or
	  WILL_FIRE_RL_doFEQ_D or
	  WILL_FIRE_RL_doFMAX_D or
	  WILL_FIRE_RL_doFMIN_D or
	  WILL_FIRE_RL_doFCVT_D_S or
	  WILL_FIRE_RL_doFCVT_S_D or
	  WILL_FIRE_RL_doFCVT_LU_D or
	  WILL_FIRE_RL_doFCVT_L_D or
	  WILL_FIRE_RL_doFCVT_D_LU or
	  WILL_FIRE_RL_doFCVT_D_L or
	  WILL_FIRE_RL_doFCVT_WU_D or
	  WILL_FIRE_RL_doFCVT_W_D or
	  WILL_FIRE_RL_doFCVT_D_WU or
	  WILL_FIRE_RL_doFCVT_D_W or
	  WILL_FIRE_RL_doFSGNJX_D or
	  WILL_FIRE_RL_doFSGNJN_D or
	  WILL_FIRE_RL_doFSGNJ_D or
	  WILL_FIRE_RL_doFSQRT_D or
	  WILL_FIRE_RL_doFDIV_D or
	  WILL_FIRE_RL_doFNMSUB_D or
	  WILL_FIRE_RL_doFNMADD_D or
	  WILL_FIRE_RL_doFMSUB_D or
	  WILL_FIRE_RL_doFMADD_D or
	  WILL_FIRE_RL_doFMUL_D or
	  WILL_FIRE_RL_doFSUB_D or
	  WILL_FIRE_RL_doFADD_D or
	  WILL_FIRE_RL_doFCLASS_S or
	  WILL_FIRE_RL_doFLE_S or
	  WILL_FIRE_RL_doFLT_S or
	  WILL_FIRE_RL_doFEQ_S or
	  WILL_FIRE_RL_doFMV_X_W or
	  WILL_FIRE_RL_doFMV_W_X or
	  WILL_FIRE_RL_doFMAX_S or
	  WILL_FIRE_RL_doFMIN_S or
	  WILL_FIRE_RL_doFCVT_WU_S or
	  WILL_FIRE_RL_doFCVT_W_S or
	  WILL_FIRE_RL_doFCVT_LU_S or
	  WILL_FIRE_RL_doFCVT_L_S or
	  WILL_FIRE_RL_doFCVT_S_WU or
	  WILL_FIRE_RL_doFCVT_S_W or
	  WILL_FIRE_RL_doFCVT_S_LU or
	  WILL_FIRE_RL_doFCVT_S_L or
	  WILL_FIRE_RL_doFSGNJX_S or
	  WILL_FIRE_RL_doFSGNJN_S or
	  WILL_FIRE_RL_doFSGNJ_S or
	  WILL_FIRE_RL_doFSQRT_S or
	  WILL_FIRE_RL_doFDIV_S or
	  WILL_FIRE_RL_doFNMSUB_S or
	  WILL_FIRE_RL_doFNMADD_S or
	  WILL_FIRE_RL_doFMSUB_S or
	  WILL_FIRE_RL_doFMADD_S or
	  WILL_FIRE_RL_doFMUL_S or
	  WILL_FIRE_RL_doFSUB_S or
	  WILL_FIRE_RL_doFADD_S or WILL_FIRE_RL_rl_reset_end)
  case (1'b1)
    WILL_FIRE_RL_rl_reset_begin: stateR$D_IN = 2'd0;
    EN_req: stateR$D_IN = 2'd1;
    WILL_FIRE_RL_rl_get_fpu_result || WILL_FIRE_RL_doFCLASS_D ||
    WILL_FIRE_RL_doFMV_X_D ||
    WILL_FIRE_RL_doFMV_D_X ||
    WILL_FIRE_RL_doFLE_D ||
    WILL_FIRE_RL_doFLT_D ||
    WILL_FIRE_RL_doFEQ_D ||
    WILL_FIRE_RL_doFMAX_D ||
    WILL_FIRE_RL_doFMIN_D ||
    WILL_FIRE_RL_doFCVT_D_S ||
    WILL_FIRE_RL_doFCVT_S_D ||
    WILL_FIRE_RL_doFCVT_LU_D ||
    WILL_FIRE_RL_doFCVT_L_D ||
    WILL_FIRE_RL_doFCVT_D_LU ||
    WILL_FIRE_RL_doFCVT_D_L ||
    WILL_FIRE_RL_doFCVT_WU_D ||
    WILL_FIRE_RL_doFCVT_W_D ||
    WILL_FIRE_RL_doFCVT_D_WU ||
    WILL_FIRE_RL_doFCVT_D_W ||
    WILL_FIRE_RL_doFSGNJX_D ||
    WILL_FIRE_RL_doFSGNJN_D ||
    WILL_FIRE_RL_doFSGNJ_D:
	stateR$D_IN = 2'd3;
    WILL_FIRE_RL_doFSQRT_D || WILL_FIRE_RL_doFDIV_D ||
    WILL_FIRE_RL_doFNMSUB_D ||
    WILL_FIRE_RL_doFNMADD_D ||
    WILL_FIRE_RL_doFMSUB_D ||
    WILL_FIRE_RL_doFMADD_D ||
    WILL_FIRE_RL_doFMUL_D ||
    WILL_FIRE_RL_doFSUB_D ||
    WILL_FIRE_RL_doFADD_D:
	stateR$D_IN = 2'd2;
    WILL_FIRE_RL_doFCLASS_S || WILL_FIRE_RL_doFLE_S || WILL_FIRE_RL_doFLT_S ||
    WILL_FIRE_RL_doFEQ_S ||
    WILL_FIRE_RL_doFMV_X_W ||
    WILL_FIRE_RL_doFMV_W_X ||
    WILL_FIRE_RL_doFMAX_S ||
    WILL_FIRE_RL_doFMIN_S ||
    WILL_FIRE_RL_doFCVT_WU_S ||
    WILL_FIRE_RL_doFCVT_W_S ||
    WILL_FIRE_RL_doFCVT_LU_S ||
    WILL_FIRE_RL_doFCVT_L_S ||
    WILL_FIRE_RL_doFCVT_S_WU ||
    WILL_FIRE_RL_doFCVT_S_W ||
    WILL_FIRE_RL_doFCVT_S_LU ||
    WILL_FIRE_RL_doFCVT_S_L ||
    WILL_FIRE_RL_doFSGNJX_S ||
    WILL_FIRE_RL_doFSGNJN_S ||
    WILL_FIRE_RL_doFSGNJ_S:
	stateR$D_IN = 2'd3;
    WILL_FIRE_RL_doFSQRT_S || WILL_FIRE_RL_doFDIV_S ||
    WILL_FIRE_RL_doFNMSUB_S ||
    WILL_FIRE_RL_doFNMADD_S ||
    WILL_FIRE_RL_doFMSUB_S ||
    WILL_FIRE_RL_doFMADD_S ||
    WILL_FIRE_RL_doFMUL_S ||
    WILL_FIRE_RL_doFSUB_S ||
    WILL_FIRE_RL_doFADD_S:
	stateR$D_IN = 2'd2;
    WILL_FIRE_RL_rl_reset_end: stateR$D_IN = 2'd1;
    default: stateR$D_IN = 2'b10 /* unspecified value */ ;
  endcase
  assign stateR$EN =
	     WILL_FIRE_RL_rl_reset_begin || WILL_FIRE_RL_rl_reset_end ||
	     EN_req ||
	     WILL_FIRE_RL_doFSQRT_D ||
	     WILL_FIRE_RL_doFDIV_D ||
	     WILL_FIRE_RL_doFNMSUB_D ||
	     WILL_FIRE_RL_doFNMADD_D ||
	     WILL_FIRE_RL_doFMSUB_D ||
	     WILL_FIRE_RL_doFMADD_D ||
	     WILL_FIRE_RL_doFMUL_D ||
	     WILL_FIRE_RL_doFSUB_D ||
	     WILL_FIRE_RL_doFADD_D ||
	     WILL_FIRE_RL_doFSQRT_S ||
	     WILL_FIRE_RL_doFDIV_S ||
	     WILL_FIRE_RL_doFNMSUB_S ||
	     WILL_FIRE_RL_doFNMADD_S ||
	     WILL_FIRE_RL_doFMSUB_S ||
	     WILL_FIRE_RL_doFMADD_S ||
	     WILL_FIRE_RL_doFMUL_S ||
	     WILL_FIRE_RL_doFSUB_S ||
	     WILL_FIRE_RL_doFADD_S ||
	     WILL_FIRE_RL_rl_get_fpu_result ||
	     WILL_FIRE_RL_doFCLASS_D ||
	     WILL_FIRE_RL_doFMV_X_D ||
	     WILL_FIRE_RL_doFMV_D_X ||
	     WILL_FIRE_RL_doFLE_D ||
	     WILL_FIRE_RL_doFLT_D ||
	     WILL_FIRE_RL_doFEQ_D ||
	     WILL_FIRE_RL_doFMAX_D ||
	     WILL_FIRE_RL_doFMIN_D ||
	     WILL_FIRE_RL_doFCVT_D_S ||
	     WILL_FIRE_RL_doFCVT_S_D ||
	     WILL_FIRE_RL_doFCVT_LU_D ||
	     WILL_FIRE_RL_doFCVT_L_D ||
	     WILL_FIRE_RL_doFCVT_D_LU ||
	     WILL_FIRE_RL_doFCVT_D_L ||
	     WILL_FIRE_RL_doFCVT_WU_D ||
	     WILL_FIRE_RL_doFCVT_W_D ||
	     WILL_FIRE_RL_doFCVT_D_WU ||
	     WILL_FIRE_RL_doFCVT_D_W ||
	     WILL_FIRE_RL_doFSGNJX_D ||
	     WILL_FIRE_RL_doFSGNJN_D ||
	     WILL_FIRE_RL_doFSGNJ_D ||
	     WILL_FIRE_RL_doFCLASS_S ||
	     WILL_FIRE_RL_doFLE_S ||
	     WILL_FIRE_RL_doFLT_S ||
	     WILL_FIRE_RL_doFEQ_S ||
	     WILL_FIRE_RL_doFMV_X_W ||
	     WILL_FIRE_RL_doFMV_W_X ||
	     WILL_FIRE_RL_doFMAX_S ||
	     WILL_FIRE_RL_doFMIN_S ||
	     WILL_FIRE_RL_doFCVT_WU_S ||
	     WILL_FIRE_RL_doFCVT_W_S ||
	     WILL_FIRE_RL_doFCVT_LU_S ||
	     WILL_FIRE_RL_doFCVT_L_S ||
	     WILL_FIRE_RL_doFCVT_S_WU ||
	     WILL_FIRE_RL_doFCVT_S_W ||
	     WILL_FIRE_RL_doFCVT_S_LU ||
	     WILL_FIRE_RL_doFCVT_S_L ||
	     WILL_FIRE_RL_doFSGNJX_S ||
	     WILL_FIRE_RL_doFSGNJN_S ||
	     WILL_FIRE_RL_doFSGNJ_S ;
  // submodule fpu
  always@(WILL_FIRE_RL_doFADD_S or
	  MUX_fpu$server_core_request_put_1__VAL_1 or
	  WILL_FIRE_RL_doFSUB_S or
	  MUX_fpu$server_core_request_put_1__VAL_2 or
	  WILL_FIRE_RL_doFMUL_S or
	  MUX_fpu$server_core_request_put_1__VAL_3 or
	  WILL_FIRE_RL_doFMADD_S or
	  MUX_fpu$server_core_request_put_1__VAL_4 or
	  WILL_FIRE_RL_doFMSUB_S or
	  MUX_fpu$server_core_request_put_1__VAL_5 or
	  WILL_FIRE_RL_doFNMADD_S or
	  MUX_fpu$server_core_request_put_1__VAL_6 or
	  WILL_FIRE_RL_doFNMSUB_S or
	  MUX_fpu$server_core_request_put_1__VAL_7 or
	  WILL_FIRE_RL_doFDIV_S or
	  MUX_fpu$server_core_request_put_1__VAL_8 or
	  WILL_FIRE_RL_doFSQRT_S or
	  MUX_fpu$server_core_request_put_1__VAL_9 or
	  WILL_FIRE_RL_doFADD_D or
	  MUX_fpu$server_core_request_put_1__VAL_10 or
	  WILL_FIRE_RL_doFSUB_D or
	  MUX_fpu$server_core_request_put_1__VAL_11 or
	  WILL_FIRE_RL_doFMUL_D or
	  MUX_fpu$server_core_request_put_1__VAL_12 or
	  WILL_FIRE_RL_doFMADD_D or
	  MUX_fpu$server_core_request_put_1__VAL_13 or
	  WILL_FIRE_RL_doFMSUB_D or
	  MUX_fpu$server_core_request_put_1__VAL_14 or
	  WILL_FIRE_RL_doFNMADD_D or
	  MUX_fpu$server_core_request_put_1__VAL_15 or
	  WILL_FIRE_RL_doFNMSUB_D or
	  MUX_fpu$server_core_request_put_1__VAL_16 or
	  WILL_FIRE_RL_doFDIV_D or
	  MUX_fpu$server_core_request_put_1__VAL_17 or
	  WILL_FIRE_RL_doFSQRT_D or MUX_fpu$server_core_request_put_1__VAL_18)
  begin
    case (1'b1) // synopsys parallel_case
      WILL_FIRE_RL_doFADD_S:
	  fpu$server_core_request_put =
	      MUX_fpu$server_core_request_put_1__VAL_1;
      WILL_FIRE_RL_doFSUB_S:
	  fpu$server_core_request_put =
	      MUX_fpu$server_core_request_put_1__VAL_2;
      WILL_FIRE_RL_doFMUL_S:
	  fpu$server_core_request_put =
	      MUX_fpu$server_core_request_put_1__VAL_3;
      WILL_FIRE_RL_doFMADD_S:
	  fpu$server_core_request_put =
	      MUX_fpu$server_core_request_put_1__VAL_4;
      WILL_FIRE_RL_doFMSUB_S:
	  fpu$server_core_request_put =
	      MUX_fpu$server_core_request_put_1__VAL_5;
      WILL_FIRE_RL_doFNMADD_S:
	  fpu$server_core_request_put =
	      MUX_fpu$server_core_request_put_1__VAL_6;
      WILL_FIRE_RL_doFNMSUB_S:
	  fpu$server_core_request_put =
	      MUX_fpu$server_core_request_put_1__VAL_7;
      WILL_FIRE_RL_doFDIV_S:
	  fpu$server_core_request_put =
	      MUX_fpu$server_core_request_put_1__VAL_8;
      WILL_FIRE_RL_doFSQRT_S:
	  fpu$server_core_request_put =
	      MUX_fpu$server_core_request_put_1__VAL_9;
      WILL_FIRE_RL_doFADD_D:
	  fpu$server_core_request_put =
	      MUX_fpu$server_core_request_put_1__VAL_10;
      WILL_FIRE_RL_doFSUB_D:
	  fpu$server_core_request_put =
	      MUX_fpu$server_core_request_put_1__VAL_11;
      WILL_FIRE_RL_doFMUL_D:
	  fpu$server_core_request_put =
	      MUX_fpu$server_core_request_put_1__VAL_12;
      WILL_FIRE_RL_doFMADD_D:
	  fpu$server_core_request_put =
	      MUX_fpu$server_core_request_put_1__VAL_13;
      WILL_FIRE_RL_doFMSUB_D:
	  fpu$server_core_request_put =
	      MUX_fpu$server_core_request_put_1__VAL_14;
      WILL_FIRE_RL_doFNMADD_D:
	  fpu$server_core_request_put =
	      MUX_fpu$server_core_request_put_1__VAL_15;
      WILL_FIRE_RL_doFNMSUB_D:
	  fpu$server_core_request_put =
	      MUX_fpu$server_core_request_put_1__VAL_16;
      WILL_FIRE_RL_doFDIV_D:
	  fpu$server_core_request_put =
	      MUX_fpu$server_core_request_put_1__VAL_17;
      WILL_FIRE_RL_doFSQRT_D:
	  fpu$server_core_request_put =
	      MUX_fpu$server_core_request_put_1__VAL_18;
      default: fpu$server_core_request_put =
		   202'h2AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA /* unspecified value */ ;
    endcase
  end
  assign fpu$EN_server_core_request_put =
	     WILL_FIRE_RL_doFADD_S || WILL_FIRE_RL_doFSUB_S ||
	     WILL_FIRE_RL_doFMUL_S ||
	     WILL_FIRE_RL_doFMADD_S ||
	     WILL_FIRE_RL_doFMSUB_S ||
	     WILL_FIRE_RL_doFNMADD_S ||
	     WILL_FIRE_RL_doFNMSUB_S ||
	     WILL_FIRE_RL_doFDIV_S ||
	     WILL_FIRE_RL_doFSQRT_S ||
	     WILL_FIRE_RL_doFADD_D ||
	     WILL_FIRE_RL_doFSUB_D ||
	     WILL_FIRE_RL_doFMUL_D ||
	     WILL_FIRE_RL_doFMADD_D ||
	     WILL_FIRE_RL_doFMSUB_D ||
	     WILL_FIRE_RL_doFNMADD_D ||
	     WILL_FIRE_RL_doFNMSUB_D ||
	     WILL_FIRE_RL_doFDIV_D ||
	     WILL_FIRE_RL_doFSQRT_D ;
  assign fpu$EN_server_core_response_get = MUX_dw_result$wset_1__SEL_1 ;
  assign fpu$EN_server_reset_request_put = CAN_FIRE_RL_rl_reset_begin ;
  assign fpu$EN_server_reset_response_get = CAN_FIRE_RL_rl_reset_end ;
  // submodule frmFpuF
  assign frmFpuF$D_IN = 1'b0 ;
  assign frmFpuF$ENQ = 1'b0 ;
  assign frmFpuF$DEQ = 1'b0 ;
  assign frmFpuF$CLR = CAN_FIRE_RL_rl_reset_begin ;
  // submodule resetReqsF
  assign resetReqsF$ENQ = EN_server_reset_request_put ;
  assign resetReqsF$DEQ =
	     fpu$RDY_server_reset_request_put && resetReqsF$EMPTY_N ;
  assign resetReqsF$CLR = 1'b0 ;
  // submodule resetRspsF
  assign resetRspsF$ENQ =
	     fpu$RDY_server_reset_response_get && resetRspsF$FULL_N &&
	     stateR == 2'd0 ;
  assign resetRspsF$DEQ = EN_server_reset_response_get ;
  assign resetRspsF$CLR = 1'b0 ;
  // remaining internal signals
  assign IF_0_CONCAT_IF_IF_0b0_CONCAT_NOT_IF_requestR_3_ETC__q117 =
	     _0_CONCAT_IF_IF_0b0_CONCAT_NOT_IF_requestR_3_BI_ETC___d3656 ?
	       _theResult___snd__h135453 :
	       _theResult____h126028 ;
  assign IF_0_CONCAT_IF_IF_3074_MINUS_SEXT_IF_IF_reques_ETC__q154 =
	     _0_CONCAT_IF_IF_3074_MINUS_SEXT_IF_IF_requestR__ETC___d4935 ?
	       _theResult___snd__h201397 :
	       _theResult____h191843 ;
  assign IF_0_CONCAT_IF_IF_3970_MINUS_SEXT_IF_requestR__ETC__q122 =
	     _0_CONCAT_IF_IF_3970_MINUS_SEXT_IF_requestR_3_B_ETC___d4100 ?
	       _theResult___snd__h155794 :
	       _theResult____h146240 ;
  assign IF_0_CONCAT_IF_IF_IF_requestR_3_BIT_214_4_THEN_ETC__q151 =
	     _0_CONCAT_IF_IF_IF_requestR_3_BIT_214_4_THEN_re_ETC___d4615 ?
	       _theResult___snd__h190495 :
	       57'd0 ;
  assign IF_0_CONCAT_IF_IF_IF_requestR_3_BIT_214_4_THEN_ETC__q157 =
	     _0_CONCAT_IF_IF_IF_requestR_3_BIT_214_4_THEN_re_ETC___d5008 ?
	       _theResult___snd__h190495 :
	       _theResult___snd__h211382 ;
  assign IF_0_CONCAT_IF_IF_requestR_3_BIT_214_4_THEN_re_ETC__q119 =
	     _0_CONCAT_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d3778 ?
	       _theResult___snd__h145298 :
	       57'd0 ;
  assign IF_0_CONCAT_IF_IF_requestR_3_BIT_214_4_THEN_re_ETC__q125 =
	     _0_CONCAT_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d4173 ?
	       _theResult___snd__h145298 :
	       _theResult___snd__h165663 ;
  assign IF_3074_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_21_ETC___d4358 =
	     _3074_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_ETC___d3422 ?
	       ((_theResult___fst_exp__h135390 == 8'd255) ?
		  requestR_BITS_191_TO_128__q1[63] :
		  ((requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
		    requestR[194:192] != 3'h3 &&
		    requestR[194:192] != 3'h4) ?
		     CASE_guard26038_0b0_requestR_BITS_191_TO_128_B_ETC__q143 :
		     CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q144)) :
	       ((_theResult___fst_exp__h145309 == 8'd255) ?
		  requestR_BITS_191_TO_128__q1[63] :
		  ((requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
		    requestR[194:192] != 3'h3 &&
		    requestR[194:192] != 3'h4) ?
		     CASE_guard36028_0b0_requestR_BITS_191_TO_128_B_ETC__q145 :
		     CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q146)) ;
  assign IF_32_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_2_ETC___d1379 =
	     _32_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d1327 ?
	       ((requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
		 requestR[194:192] != 3'h3 &&
		 requestR[194:192] != 3'h4) ?
		  CASE_guard4468_0b0_requestR_BITS_191_TO_128_BI_ETC__q45 :
		  CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q46) :
	       ((x__h35010[7:0] == 8'd255) ?
		  requestR_BITS_191_TO_128__q1[31] :
		  ((requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
		    requestR[194:192] != 3'h3 &&
		    requestR[194:192] != 3'h4) ?
		     CASE_guard4995_0b0_requestR_BITS_191_TO_128_BI_ETC__q47 :
		     CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q48)) ;
  assign IF_32_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_2_ETC___d1529 =
	     _32_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d1327 ?
	       guard__h34468 != 2'b0 :
	       x__h35010[7:0] != 8'd255 && guard__h34995 != 2'b0 ;
  assign IF_32_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_2_ETC___d2398 =
	     _32_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d2347 ?
	       ((requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
		 requestR[194:192] != 3'h3 &&
		 requestR[194:192] != 3'h4) ?
		  CASE_guard9399_0b0_requestR_BITS_191_TO_128_BI_ETC__q72 :
		  CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q73) :
	       ((x__h70144[10:0] == 11'd2047) ?
		  requestR_BITS_191_TO_128__q1[31] :
		  ((requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
		    requestR[194:192] != 3'h3 &&
		    requestR[194:192] != 3'h4) ?
		     CASE_guard0129_0b0_requestR_BITS_191_TO_128_BI_ETC__q74 :
		     CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q75)) ;
  assign IF_32_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_2_ETC___d2513 =
	     _32_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d2347 ?
	       guard__h69399 != 2'b0 :
	       x__h70144[10:0] != 11'd2047 && guard__h70129 != 2'b0 ;
  assign IF_32_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214__ETC___d1718 =
	     _32_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d1580 ?
	       guard__h41384 != 2'b0 :
	       x__h41925[7:0] != 8'd255 && guard__h41910 != 2'b0 ;
  assign IF_32_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214__ETC___d2697 =
	     _32_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d2561 ?
	       guard__h80346 != 2'b0 :
	       x__h81090[10:0] != 11'd2047 && guard__h81075 != 2'b0 ;
  assign IF_64_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_2_ETC___d2937 =
	     _64_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d2888 ?
	       ((requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
		 requestR[194:192] != 3'h3 &&
		 requestR[194:192] != 3'h4) ?
		  CASE_guard5721_0b0_requestR_BITS_191_TO_128_BI_ETC__q97 :
		  CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q98) :
	       ((x__h96466[10:0] == 11'd2047) ?
		  requestR_BITS_191_TO_128__q1[63] :
		  ((requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
		    requestR[194:192] != 3'h3 &&
		    requestR[194:192] != 3'h4) ?
		     CASE_guard6451_0b0_requestR_BITS_191_TO_128_BI_ETC__q99 :
		     CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q100)) ;
  assign IF_64_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_2_ETC___d3054 =
	     _64_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d2888 ?
	       guard__h95721 != 2'b0 :
	       x__h96466[10:0] != 11'd2047 && guard__h96451 != 2'b0 ;
  assign IF_64_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_2_ETC___d511 =
	     _64_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d450 ?
	       ((requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
		 requestR[194:192] != 3'h3 &&
		 requestR[194:192] != 3'h4) ?
		  CASE_guard5015_0b0_requestR_BITS_191_TO_128_BI_ETC__q13 :
		  CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q14) :
	       ((x__h15560[7:0] == 8'd255) ?
		  requestR_BITS_191_TO_128__q1[63] :
		  ((requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
		    requestR[194:192] != 3'h3 &&
		    requestR[194:192] != 3'h4) ?
		     CASE_guard5545_0b0_requestR_BITS_191_TO_128_BI_ETC__q15 :
		     CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q16)) ;
  assign IF_64_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_2_ETC___d693 =
	     _64_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d450 ?
	       guard__h15015 != 2'b0 :
	       x__h15560[7:0] != 8'd255 && guard__h15545 != 2'b0 ;
  assign IF_64_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214__ETC___d1174 =
	     _64_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d972 ?
	       guard__h27296 != 2'b0 :
	       x__h27837[7:0] != 8'd255 && guard__h27822 != 2'b0 ;
  assign IF_64_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214__ETC___d3208 =
	     _64_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d3071 ?
	       guard__h108246 != 2'b0 :
	       x__h108990[10:0] != 11'd2047 && guard__h108975 != 2'b0 ;
  assign IF_IF_0b0_CONCAT_NOT_IF_requestR_3_BIT_214_4_T_ETC___d3654 =
	     (_theResult____h126028[56] ?
		6'd0 :
		(_theResult____h126028[55] ?
		   6'd1 :
		   (_theResult____h126028[54] ?
		      6'd2 :
		      (_theResult____h126028[53] ?
			 6'd3 :
			 (_theResult____h126028[52] ?
			    6'd4 :
			    (_theResult____h126028[51] ?
			       6'd5 :
			       (_theResult____h126028[50] ?
				  6'd6 :
				  (_theResult____h126028[49] ?
				     6'd7 :
				     (_theResult____h126028[48] ?
					6'd8 :
					(_theResult____h126028[47] ?
					   6'd9 :
					   (_theResult____h126028[46] ?
					      6'd10 :
					      (_theResult____h126028[45] ?
						 6'd11 :
						 (_theResult____h126028[44] ?
						    6'd12 :
						    (_theResult____h126028[43] ?
						       6'd13 :
						       (_theResult____h126028[42] ?
							  6'd14 :
							  (_theResult____h126028[41] ?
							     6'd15 :
							     (_theResult____h126028[40] ?
								6'd16 :
								(_theResult____h126028[39] ?
								   6'd17 :
								   (_theResult____h126028[38] ?
								      6'd18 :
								      (_theResult____h126028[37] ?
									 6'd19 :
									 (_theResult____h126028[36] ?
									    6'd20 :
									    (_theResult____h126028[35] ?
									       6'd21 :
									       (_theResult____h126028[34] ?
										  6'd22 :
										  (_theResult____h126028[33] ?
										     6'd23 :
										     (_theResult____h126028[32] ?
											6'd24 :
											(_theResult____h126028[31] ?
											   6'd25 :
											   (_theResult____h126028[30] ?
											      6'd26 :
											      (_theResult____h126028[29] ?
												 6'd27 :
												 (_theResult____h126028[28] ?
												    6'd28 :
												    (_theResult____h126028[27] ?
												       6'd29 :
												       (_theResult____h126028[26] ?
													  6'd30 :
													  (_theResult____h126028[25] ?
													     6'd31 :
													     (_theResult____h126028[24] ?
														6'd32 :
														(_theResult____h126028[23] ?
														   6'd33 :
														   (_theResult____h126028[22] ?
														      6'd34 :
														      (_theResult____h126028[21] ?
															 6'd35 :
															 (_theResult____h126028[20] ?
															    6'd36 :
															    (_theResult____h126028[19] ?
															       6'd37 :
															       (_theResult____h126028[18] ?
																  6'd38 :
																  (_theResult____h126028[17] ?
																     6'd39 :
																     (_theResult____h126028[16] ?
																	6'd40 :
																	(_theResult____h126028[15] ?
																	   6'd41 :
																	   (_theResult____h126028[14] ?
																	      6'd42 :
																	      (_theResult____h126028[13] ?
																		 6'd43 :
																		 (_theResult____h126028[12] ?
																		    6'd44 :
																		    (_theResult____h126028[11] ?
																		       6'd45 :
																		       (_theResult____h126028[10] ?
																			  6'd46 :
																			  (_theResult____h126028[9] ?
																			     6'd47 :
																			     (_theResult____h126028[8] ?
																				6'd48 :
																				(_theResult____h126028[7] ?
																				   6'd49 :
																				   (_theResult____h126028[6] ?
																				      6'd50 :
																				      (_theResult____h126028[5] ?
																					 6'd51 :
																					 (_theResult____h126028[4] ?
																					    6'd52 :
																					    (_theResult____h126028[3] ?
																					       6'd53 :
																					       (_theResult____h126028[2] ?
																						  6'd54 :
																						  (_theResult____h126028[1] ?
																						     6'd55 :
																						     (_theResult____h126028[0] ?
																							6'd56 :
																							6'd57))))))))))))))))))))))))))))))))))))))))))))))))))))))))) -
	     6'd1 ;
  assign IF_IF_3074_MINUS_SEXT_IF_IF_requestR_3_BIT_214_ETC___d4933 =
	     (_theResult____h191843[56] ?
		6'd0 :
		(_theResult____h191843[55] ?
		   6'd1 :
		   (_theResult____h191843[54] ?
		      6'd2 :
		      (_theResult____h191843[53] ?
			 6'd3 :
			 (_theResult____h191843[52] ?
			    6'd4 :
			    (_theResult____h191843[51] ?
			       6'd5 :
			       (_theResult____h191843[50] ?
				  6'd6 :
				  (_theResult____h191843[49] ?
				     6'd7 :
				     (_theResult____h191843[48] ?
					6'd8 :
					(_theResult____h191843[47] ?
					   6'd9 :
					   (_theResult____h191843[46] ?
					      6'd10 :
					      (_theResult____h191843[45] ?
						 6'd11 :
						 (_theResult____h191843[44] ?
						    6'd12 :
						    (_theResult____h191843[43] ?
						       6'd13 :
						       (_theResult____h191843[42] ?
							  6'd14 :
							  (_theResult____h191843[41] ?
							     6'd15 :
							     (_theResult____h191843[40] ?
								6'd16 :
								(_theResult____h191843[39] ?
								   6'd17 :
								   (_theResult____h191843[38] ?
								      6'd18 :
								      (_theResult____h191843[37] ?
									 6'd19 :
									 (_theResult____h191843[36] ?
									    6'd20 :
									    (_theResult____h191843[35] ?
									       6'd21 :
									       (_theResult____h191843[34] ?
										  6'd22 :
										  (_theResult____h191843[33] ?
										     6'd23 :
										     (_theResult____h191843[32] ?
											6'd24 :
											(_theResult____h191843[31] ?
											   6'd25 :
											   (_theResult____h191843[30] ?
											      6'd26 :
											      (_theResult____h191843[29] ?
												 6'd27 :
												 (_theResult____h191843[28] ?
												    6'd28 :
												    (_theResult____h191843[27] ?
												       6'd29 :
												       (_theResult____h191843[26] ?
													  6'd30 :
													  (_theResult____h191843[25] ?
													     6'd31 :
													     (_theResult____h191843[24] ?
														6'd32 :
														(_theResult____h191843[23] ?
														   6'd33 :
														   (_theResult____h191843[22] ?
														      6'd34 :
														      (_theResult____h191843[21] ?
															 6'd35 :
															 (_theResult____h191843[20] ?
															    6'd36 :
															    (_theResult____h191843[19] ?
															       6'd37 :
															       (_theResult____h191843[18] ?
																  6'd38 :
																  (_theResult____h191843[17] ?
																     6'd39 :
																     (_theResult____h191843[16] ?
																	6'd40 :
																	(_theResult____h191843[15] ?
																	   6'd41 :
																	   (_theResult____h191843[14] ?
																	      6'd42 :
																	      (_theResult____h191843[13] ?
																		 6'd43 :
																		 (_theResult____h191843[12] ?
																		    6'd44 :
																		    (_theResult____h191843[11] ?
																		       6'd45 :
																		       (_theResult____h191843[10] ?
																			  6'd46 :
																			  (_theResult____h191843[9] ?
																			     6'd47 :
																			     (_theResult____h191843[8] ?
																				6'd48 :
																				(_theResult____h191843[7] ?
																				   6'd49 :
																				   (_theResult____h191843[6] ?
																				      6'd50 :
																				      (_theResult____h191843[5] ?
																					 6'd51 :
																					 (_theResult____h191843[4] ?
																					    6'd52 :
																					    (_theResult____h191843[3] ?
																					       6'd53 :
																					       (_theResult____h191843[2] ?
																						  6'd54 :
																						  (_theResult____h191843[1] ?
																						     6'd55 :
																						     (_theResult____h191843[0] ?
																							6'd56 :
																							6'd57))))))))))))))))))))))))))))))))))))))))))))))))))))))))) -
	     6'd1 ;
  assign IF_IF_3970_MINUS_SEXT_IF_requestR_3_BIT_214_4__ETC___d4098 =
	     (_theResult____h146240[56] ?
		6'd0 :
		(_theResult____h146240[55] ?
		   6'd1 :
		   (_theResult____h146240[54] ?
		      6'd2 :
		      (_theResult____h146240[53] ?
			 6'd3 :
			 (_theResult____h146240[52] ?
			    6'd4 :
			    (_theResult____h146240[51] ?
			       6'd5 :
			       (_theResult____h146240[50] ?
				  6'd6 :
				  (_theResult____h146240[49] ?
				     6'd7 :
				     (_theResult____h146240[48] ?
					6'd8 :
					(_theResult____h146240[47] ?
					   6'd9 :
					   (_theResult____h146240[46] ?
					      6'd10 :
					      (_theResult____h146240[45] ?
						 6'd11 :
						 (_theResult____h146240[44] ?
						    6'd12 :
						    (_theResult____h146240[43] ?
						       6'd13 :
						       (_theResult____h146240[42] ?
							  6'd14 :
							  (_theResult____h146240[41] ?
							     6'd15 :
							     (_theResult____h146240[40] ?
								6'd16 :
								(_theResult____h146240[39] ?
								   6'd17 :
								   (_theResult____h146240[38] ?
								      6'd18 :
								      (_theResult____h146240[37] ?
									 6'd19 :
									 (_theResult____h146240[36] ?
									    6'd20 :
									    (_theResult____h146240[35] ?
									       6'd21 :
									       (_theResult____h146240[34] ?
										  6'd22 :
										  (_theResult____h146240[33] ?
										     6'd23 :
										     (_theResult____h146240[32] ?
											6'd24 :
											(_theResult____h146240[31] ?
											   6'd25 :
											   (_theResult____h146240[30] ?
											      6'd26 :
											      (_theResult____h146240[29] ?
												 6'd27 :
												 (_theResult____h146240[28] ?
												    6'd28 :
												    (_theResult____h146240[27] ?
												       6'd29 :
												       (_theResult____h146240[26] ?
													  6'd30 :
													  (_theResult____h146240[25] ?
													     6'd31 :
													     (_theResult____h146240[24] ?
														6'd32 :
														(_theResult____h146240[23] ?
														   6'd33 :
														   (_theResult____h146240[22] ?
														      6'd34 :
														      (_theResult____h146240[21] ?
															 6'd35 :
															 (_theResult____h146240[20] ?
															    6'd36 :
															    (_theResult____h146240[19] ?
															       6'd37 :
															       (_theResult____h146240[18] ?
																  6'd38 :
																  (_theResult____h146240[17] ?
																     6'd39 :
																     (_theResult____h146240[16] ?
																	6'd40 :
																	(_theResult____h146240[15] ?
																	   6'd41 :
																	   (_theResult____h146240[14] ?
																	      6'd42 :
																	      (_theResult____h146240[13] ?
																		 6'd43 :
																		 (_theResult____h146240[12] ?
																		    6'd44 :
																		    (_theResult____h146240[11] ?
																		       6'd45 :
																		       (_theResult____h146240[10] ?
																			  6'd46 :
																			  (_theResult____h146240[9] ?
																			     6'd47 :
																			     (_theResult____h146240[8] ?
																				6'd48 :
																				(_theResult____h146240[7] ?
																				   6'd49 :
																				   (_theResult____h146240[6] ?
																				      6'd50 :
																				      (_theResult____h146240[5] ?
																					 6'd51 :
																					 (_theResult____h146240[4] ?
																					    6'd52 :
																					    (_theResult____h146240[3] ?
																					       6'd53 :
																					       (_theResult____h146240[2] ?
																						  6'd54 :
																						  (_theResult____h146240[1] ?
																						     6'd55 :
																						     (_theResult____h146240[0] ?
																							6'd56 :
																							6'd57))))))))))))))))))))))))))))))))))))))))))))))))))))))))) -
	     6'd1 ;
  assign IF_IF_IF_IF_0b0_CONCAT_NOT_IF_requestR_3_BIT_2_ETC___d3713 =
	     (guard__h126038 == 2'b0 || requestR_BITS_191_TO_128__q1[63]) ?
	       _theResult___fst_exp__h135390 :
	       _theResult___exp__h135916 ;
  assign IF_IF_IF_IF_0b0_CONCAT_NOT_IF_requestR_3_BIT_2_ETC___d3715 =
	     (guard__h126038 == 2'b0) ?
	       _theResult___fst_exp__h135390 :
	       (requestR_BITS_191_TO_128__q1[63] ?
		  _theResult___exp__h135916 :
		  _theResult___fst_exp__h135390) ;
  assign IF_IF_IF_IF_0b0_CONCAT_NOT_IF_requestR_3_BIT_2_ETC___d4260 =
	     (guard__h126038 == 2'b0 || requestR_BITS_191_TO_128__q1[63]) ?
	       sfdin__h135384[56:34] :
	       _theResult___sfd__h135917 ;
  assign IF_IF_IF_IF_0b0_CONCAT_NOT_IF_requestR_3_BIT_2_ETC___d4262 =
	     (guard__h126038 == 2'b0) ?
	       sfdin__h135384[56:34] :
	       (requestR_BITS_191_TO_128__q1[63] ?
		  _theResult___sfd__h135917 :
		  sfdin__h135384[56:34]) ;
  assign IF_IF_IF_IF_3074_MINUS_SEXT_IF_IF_requestR_3_B_ETC___d4992 =
	     (guard__h191853 == 2'b0 ||
	      requestR_BITS_191_TO_128__q1[63:32] == 32'hFFFFFFFF &&
	      requestR_BITS_191_TO_128__q1[31]) ?
	       _theResult___fst_exp__h201334 :
	       _theResult___exp__h202063 ;
  assign IF_IF_IF_IF_3074_MINUS_SEXT_IF_IF_requestR_3_B_ETC___d4994 =
	     (guard__h191853 == 2'b0) ?
	       _theResult___fst_exp__h201334 :
	       ((requestR_BITS_191_TO_128__q1[63:32] == 32'hFFFFFFFF &&
		 requestR_BITS_191_TO_128__q1[31]) ?
		  _theResult___exp__h202063 :
		  _theResult___fst_exp__h201334) ;
  assign IF_IF_IF_IF_3074_MINUS_SEXT_IF_IF_requestR_3_B_ETC___d5121 =
	     (guard__h191853 == 2'b0 ||
	      requestR_BITS_191_TO_128__q1[63:32] == 32'hFFFFFFFF &&
	      requestR_BITS_191_TO_128__q1[31]) ?
	       sfdin__h201328[56:5] :
	       _theResult___sfd__h202064 ;
  assign IF_IF_IF_IF_3074_MINUS_SEXT_IF_IF_requestR_3_B_ETC___d5123 =
	     (guard__h191853 == 2'b0) ?
	       sfdin__h201328[56:5] :
	       ((requestR_BITS_191_TO_128__q1[63:32] == 32'hFFFFFFFF &&
		 requestR_BITS_191_TO_128__q1[31]) ?
		  _theResult___sfd__h202064 :
		  sfdin__h201328[56:5]) ;
  assign IF_IF_IF_IF_3970_MINUS_SEXT_IF_requestR_3_BIT__ETC___d4157 =
	     (guard__h146250 == 2'b0 || requestR_BITS_191_TO_128__q1[63]) ?
	       _theResult___fst_exp__h155731 :
	       _theResult___exp__h156257 ;
  assign IF_IF_IF_IF_3970_MINUS_SEXT_IF_requestR_3_BIT__ETC___d4159 =
	     (guard__h146250 == 2'b0) ?
	       _theResult___fst_exp__h155731 :
	       (requestR_BITS_191_TO_128__q1[63] ?
		  _theResult___exp__h156257 :
		  _theResult___fst_exp__h155731) ;
  assign IF_IF_IF_IF_3970_MINUS_SEXT_IF_requestR_3_BIT__ETC___d4306 =
	     (guard__h146250 == 2'b0 || requestR_BITS_191_TO_128__q1[63]) ?
	       sfdin__h155725[56:34] :
	       _theResult___sfd__h156258 ;
  assign IF_IF_IF_IF_3970_MINUS_SEXT_IF_requestR_3_BIT__ETC___d4308 =
	     (guard__h146250 == 2'b0) ?
	       sfdin__h155725[56:34] :
	       (requestR_BITS_191_TO_128__q1[63] ?
		  _theResult___sfd__h156258 :
		  sfdin__h155725[56:34]) ;
  assign IF_IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d4667 =
	     (guard__h181312 == 2'b0 ||
	      requestR_BITS_191_TO_128__q1[63:32] == 32'hFFFFFFFF &&
	      requestR_BITS_191_TO_128__q1[31]) ?
	       _theResult___fst_exp__h190506 :
	       _theResult___exp__h191161 ;
  assign IF_IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d4669 =
	     (guard__h181312 == 2'b0) ?
	       _theResult___fst_exp__h190506 :
	       ((requestR_BITS_191_TO_128__q1[63:32] == 32'hFFFFFFFF &&
		 requestR_BITS_191_TO_128__q1[31]) ?
		  _theResult___exp__h191161 :
		  _theResult___fst_exp__h190506) ;
  assign IF_IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d5061 =
	     (guard__h202175 == 2'b0 ||
	      requestR_BITS_191_TO_128__q1[63:32] == 32'hFFFFFFFF &&
	      requestR_BITS_191_TO_128__q1[31]) ?
	       _theResult___fst_exp__h211398 :
	       _theResult___exp__h212078 ;
  assign IF_IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d5063 =
	     (guard__h202175 == 2'b0) ?
	       _theResult___fst_exp__h211398 :
	       ((requestR_BITS_191_TO_128__q1[63:32] == 32'hFFFFFFFF &&
		 requestR_BITS_191_TO_128__q1[31]) ?
		  _theResult___exp__h212078 :
		  _theResult___fst_exp__h211398) ;
  assign IF_IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d5094 =
	     (guard__h181312 == 2'b0 ||
	      requestR_BITS_191_TO_128__q1[63:32] == 32'hFFFFFFFF &&
	      requestR_BITS_191_TO_128__q1[31]) ?
	       _theResult___snd__h190457[56:5] :
	       _theResult___sfd__h191162 ;
  assign IF_IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d5096 =
	     (guard__h181312 == 2'b0) ?
	       _theResult___snd__h190457[56:5] :
	       ((requestR_BITS_191_TO_128__q1[63:32] == 32'hFFFFFFFF &&
		 requestR_BITS_191_TO_128__q1[31]) ?
		  _theResult___sfd__h191162 :
		  _theResult___snd__h190457[56:5]) ;
  assign IF_IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d5140 =
	     (guard__h202175 == 2'b0 ||
	      requestR_BITS_191_TO_128__q1[63:32] == 32'hFFFFFFFF &&
	      requestR_BITS_191_TO_128__q1[31]) ?
	       _theResult___snd__h211344[56:5] :
	       _theResult___sfd__h212079 ;
  assign IF_IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d5142 =
	     (guard__h202175 == 2'b0) ?
	       _theResult___snd__h211344[56:5] :
	       ((requestR_BITS_191_TO_128__q1[63:32] == 32'hFFFFFFFF &&
		 requestR_BITS_191_TO_128__q1[31]) ?
		  _theResult___sfd__h212079 :
		  _theResult___snd__h211344[56:5]) ;
  assign IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d1401 =
	     (guard__h34468 == 2'b0) ?
	       8'd0 :
	       (requestR_BITS_191_TO_128__q1[31] ?
		  _theResult___exp__h34881 :
		  8'd0) ;
  assign IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d1427 =
	     (guard__h34995 == 2'b0 || requestR_BITS_191_TO_128__q1[31]) ?
	       x__h35010[7:0] :
	       _theResult___exp__h35434 ;
  assign IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d1429 =
	     (guard__h34995 == 2'b0) ?
	       x__h35010[7:0] :
	       (requestR_BITS_191_TO_128__q1[31] ?
		  _theResult___exp__h35434 :
		  x__h35010[7:0]) ;
  assign IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d1450 =
	     (guard__h34468 == 2'b0 || requestR_BITS_191_TO_128__q1[31]) ?
	       sfd___3__h34458[31:9] :
	       _theResult___sfd__h34882 ;
  assign IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d1452 =
	     (guard__h34468 == 2'b0) ?
	       sfd___3__h34458[31:9] :
	       (requestR_BITS_191_TO_128__q1[31] ?
		  _theResult___sfd__h34882 :
		  sfd___3__h34458[31:9]) ;
  assign IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d1468 =
	     (guard__h34995 == 2'b0 || requestR_BITS_191_TO_128__q1[31]) ?
	       sfd___3__h34458[30:8] :
	       _theResult___sfd__h35435 ;
  assign IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d1470 =
	     (guard__h34995 == 2'b0) ?
	       sfd___3__h34458[30:8] :
	       (requestR_BITS_191_TO_128__q1[31] ?
		  _theResult___sfd__h35435 :
		  sfd___3__h34458[30:8]) ;
  assign IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d2419 =
	     (guard__h69399 == 2'b0) ?
	       11'd0 :
	       (requestR_BITS_191_TO_128__q1[31] ?
		  _theResult___exp__h70015 :
		  11'd0) ;
  assign IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d2445 =
	     (guard__h70129 == 2'b0 || requestR_BITS_191_TO_128__q1[31]) ?
	       x__h70144[10:0] :
	       _theResult___exp__h70771 ;
  assign IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d2447 =
	     (guard__h70129 == 2'b0) ?
	       x__h70144[10:0] :
	       (requestR_BITS_191_TO_128__q1[31] ?
		  _theResult___exp__h70771 :
		  x__h70144[10:0]) ;
  assign IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d2468 =
	     (guard__h69399 == 2'b0 || requestR_BITS_191_TO_128__q1[31]) ?
	       sfd___3__h69389[54:3] :
	       _theResult___sfd__h70016 ;
  assign IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d2470 =
	     (guard__h69399 == 2'b0) ?
	       sfd___3__h69389[54:3] :
	       (requestR_BITS_191_TO_128__q1[31] ?
		  _theResult___sfd__h70016 :
		  sfd___3__h69389[54:3]) ;
  assign IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d2486 =
	     (guard__h70129 == 2'b0 || requestR_BITS_191_TO_128__q1[31]) ?
	       sfd___3__h69389[53:2] :
	       _theResult___sfd__h70772 ;
  assign IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d2488 =
	     (guard__h70129 == 2'b0) ?
	       sfd___3__h69389[53:2] :
	       (requestR_BITS_191_TO_128__q1[31] ?
		  _theResult___sfd__h70772 :
		  sfd___3__h69389[53:2]) ;
  assign IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d2958 =
	     (guard__h95721 == 2'b0) ?
	       11'd0 :
	       (requestR_BITS_191_TO_128__q1[63] ?
		  _theResult___exp__h96337 :
		  11'd0) ;
  assign IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d2984 =
	     (guard__h96451 == 2'b0 || requestR_BITS_191_TO_128__q1[63]) ?
	       x__h96466[10:0] :
	       _theResult___exp__h97093 ;
  assign IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d2986 =
	     (guard__h96451 == 2'b0) ?
	       x__h96466[10:0] :
	       (requestR_BITS_191_TO_128__q1[63] ?
		  _theResult___exp__h97093 :
		  x__h96466[10:0]) ;
  assign IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d3007 =
	     (guard__h95721 == 2'b0 || requestR_BITS_191_TO_128__q1[63]) ?
	       sfd___3__h15005[63:12] :
	       _theResult___sfd__h96338 ;
  assign IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d3009 =
	     (guard__h95721 == 2'b0) ?
	       sfd___3__h15005[63:12] :
	       (requestR_BITS_191_TO_128__q1[63] ?
		  _theResult___sfd__h96338 :
		  sfd___3__h15005[63:12]) ;
  assign IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d3025 =
	     (guard__h96451 == 2'b0 || requestR_BITS_191_TO_128__q1[63]) ?
	       sfd___3__h15005[62:11] :
	       _theResult___sfd__h97094 ;
  assign IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d3027 =
	     (guard__h96451 == 2'b0) ?
	       sfd___3__h15005[62:11] :
	       (requestR_BITS_191_TO_128__q1[63] ?
		  _theResult___sfd__h97094 :
		  sfd___3__h15005[62:11]) ;
  assign IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d3830 =
	     (guard__h136028 == 2'b0 || requestR_BITS_191_TO_128__q1[63]) ?
	       _theResult___fst_exp__h145309 :
	       _theResult___exp__h145761 ;
  assign IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d3832 =
	     (guard__h136028 == 2'b0) ?
	       _theResult___fst_exp__h145309 :
	       (requestR_BITS_191_TO_128__q1[63] ?
		  _theResult___exp__h145761 :
		  _theResult___fst_exp__h145309) ;
  assign IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d4226 =
	     (guard__h156369 == 2'b0 || requestR_BITS_191_TO_128__q1[63]) ?
	       _theResult___fst_exp__h165679 :
	       _theResult___exp__h166156 ;
  assign IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d4228 =
	     (guard__h156369 == 2'b0) ?
	       _theResult___fst_exp__h165679 :
	       (requestR_BITS_191_TO_128__q1[63] ?
		  _theResult___exp__h166156 :
		  _theResult___fst_exp__h165679) ;
  assign IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d4279 =
	     (guard__h136028 == 2'b0 || requestR_BITS_191_TO_128__q1[63]) ?
	       _theResult___snd__h145260[56:34] :
	       _theResult___sfd__h145762 ;
  assign IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d4281 =
	     (guard__h136028 == 2'b0) ?
	       _theResult___snd__h145260[56:34] :
	       (requestR_BITS_191_TO_128__q1[63] ?
		  _theResult___sfd__h145762 :
		  _theResult___snd__h145260[56:34]) ;
  assign IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d4325 =
	     (guard__h156369 == 2'b0 || requestR_BITS_191_TO_128__q1[63]) ?
	       _theResult___snd__h165625[56:34] :
	       _theResult___sfd__h166157 ;
  assign IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d4327 =
	     (guard__h156369 == 2'b0) ?
	       _theResult___snd__h165625[56:34] :
	       (requestR_BITS_191_TO_128__q1[63] ?
		  _theResult___sfd__h166157 :
		  _theResult___snd__h165625[56:34]) ;
  assign IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d533 =
	     (guard__h15015 == 2'b0) ?
	       8'd0 :
	       (requestR_BITS_191_TO_128__q1[63] ?
		  _theResult___exp__h15431 :
		  8'd0) ;
  assign IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d559 =
	     (guard__h15545 == 2'b0 || requestR_BITS_191_TO_128__q1[63]) ?
	       x__h15560[7:0] :
	       _theResult___exp__h15984 ;
  assign IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d561 =
	     (guard__h15545 == 2'b0) ?
	       x__h15560[7:0] :
	       (requestR_BITS_191_TO_128__q1[63] ?
		  _theResult___exp__h15984 :
		  x__h15560[7:0]) ;
  assign IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d582 =
	     (guard__h15015 == 2'b0 || requestR_BITS_191_TO_128__q1[63]) ?
	       sfd___3__h15005[63:41] :
	       _theResult___sfd__h15432 ;
  assign IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d584 =
	     (guard__h15015 == 2'b0) ?
	       sfd___3__h15005[63:41] :
	       (requestR_BITS_191_TO_128__q1[63] ?
		  _theResult___sfd__h15432 :
		  sfd___3__h15005[63:41]) ;
  assign IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d600 =
	     (guard__h15545 == 2'b0 || requestR_BITS_191_TO_128__q1[63]) ?
	       sfd___3__h15005[62:40] :
	       _theResult___sfd__h15985 ;
  assign IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d602 =
	     (guard__h15545 == 2'b0) ?
	       sfd___3__h15005[62:40] :
	       (requestR_BITS_191_TO_128__q1[63] ?
		  _theResult___sfd__h15985 :
		  sfd___3__h15005[62:40]) ;
  assign IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3__ETC___d1318 =
	     sfd__h28849[31] ?
	       6'd0 :
	       (sfd__h28849[30] ?
		  6'd1 :
		  (sfd__h28849[29] ?
		     6'd2 :
		     (sfd__h28849[28] ?
			6'd3 :
			(sfd__h28849[27] ?
			   6'd4 :
			   (sfd__h28849[26] ?
			      6'd5 :
			      (sfd__h28849[25] ?
				 6'd6 :
				 (sfd__h28849[24] ?
				    6'd7 :
				    (sfd__h28849[23] ?
				       6'd8 :
				       (sfd__h28849[22] ?
					  6'd9 :
					  (sfd__h28849[21] ?
					     6'd10 :
					     (sfd__h28849[20] ?
						6'd11 :
						(sfd__h28849[19] ?
						   6'd12 :
						   (sfd__h28849[18] ?
						      6'd13 :
						      (sfd__h28849[17] ?
							 6'd14 :
							 (sfd__h28849[16] ?
							    6'd15 :
							    (sfd__h28849[15] ?
							       6'd16 :
							       (sfd__h28849[14] ?
								  6'd17 :
								  (sfd__h28849[13] ?
								     6'd18 :
								     (sfd__h28849[12] ?
									6'd19 :
									(sfd__h28849[11] ?
									   6'd20 :
									   (sfd__h28849[10] ?
									      6'd21 :
									      (sfd__h28849[9] ?
										 6'd22 :
										 (sfd__h28849[8] ?
										    6'd23 :
										    (sfd__h28849[7] ?
										       6'd24 :
										       (sfd__h28849[6] ?
											  6'd25 :
											  (sfd__h28849[5] ?
											     6'd26 :
											     (sfd__h28849[4] ?
												6'd27 :
												(sfd__h28849[3] ?
												   6'd28 :
												   (sfd__h28849[2] ?
												      6'd29 :
												      (sfd__h28849[1] ?
													 6'd30 :
													 (sfd__h28849[0] ?
													    6'd31 :
													    6'd32))))))))))))))))))))))))))))))) ;
  assign IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3__ETC___d1816 =
	     (sV1_exp__h1472 == 8'd255 && sV1_sfd__h1473 == 23'd0) ?
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1745 :
	       ((sV1_exp__h1472 == 8'd0 && sV1_sfd__h1473 == 23'd0) ?
		  64'd0 :
		  IF_NEG_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_re_ETC___d1814) ;
  assign IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3__ETC___d1876 =
	     (sV1_exp__h1472 == 8'd0 && sV1_sfd__h1473 == 23'd0) ?
	       64'd0 :
	       (NEG_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d1847[19] ?
		  64'hFFFFFFFFFFFFFFFF :
		  IF_NEG_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_re_ETC___d1874) ;
  assign IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3__ETC___d1967 =
	     (sV1_exp__h1472 == 8'd255 && sV1_sfd__h1473 == 23'd0) ?
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1904 :
	       ((sV1_exp__h1472 == 8'd0 && sV1_sfd__h1473 == 23'd0) ?
		  32'd0 :
		  IF_NEG_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_re_ETC___d1965) ;
  assign IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3__ETC___d2022 =
	     (sV1_exp__h1472 == 8'd0 && sV1_sfd__h1473 == 23'd0) ?
	       32'd0 :
	       (NEG_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d1993[19] ?
		  32'hFFFFFFFF :
		  IF_NEG_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_re_ETC___d2020) ;
  assign IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3__ETC___d2108 =
	     (sV2_exp__h1597 == 8'd255 && sV2_sfd__h1598[22] ||
	      IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2077) ?
	       { requestR_BITS_191_TO_128__q1[63:32] == 32'hFFFFFFFF &&
		 requestR_BITS_191_TO_128__q1[31],
		 IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d37 } :
	       (IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2081 ?
		  IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d48 :
		  IF_NOT_IF_IF_requestR_3_BIT_214_4_THEN_request_ETC___d2106) ;
  assign IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3__ETC___d2109 =
	     (sV1_exp__h1472 == 8'd255 && sV1_sfd__h1473[22]) ?
	       IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d48 :
	       IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3__ETC___d2108 ;
  assign IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3__ETC___d2111 =
	     (sV1_exp__h1472 == 8'd255 && sV1_sfd__h1473[22] &&
	      sV2_exp__h1597 == 8'd255 &&
	      sV2_sfd__h1598[22]) ?
	       64'hFFFFFFFF7FC00000 :
	       { 32'hFFFFFFFF,
		 IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3__ETC___d2109 } ;
  assign IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3__ETC___d2112 =
	     (sV2_exp__h1597 == 8'd255 && sV2_sfd__h1598 != 23'd0 &&
	      !sV2_sfd__h1598[22]) ?
	       res__h49096 :
	       IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3__ETC___d2111 ;
  assign IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3__ETC___d2113 =
	     (sV1_exp__h1472 == 8'd255 && sV1_sfd__h1473 != 23'd0 &&
	      !sV1_sfd__h1473[22]) ?
	       res__h48859 :
	       IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3__ETC___d2112 ;
  assign IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3__ETC___d2123 =
	     IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2081 ?
	       { requestR_BITS_191_TO_128__q1[63:32] == 32'hFFFFFFFF &&
		 requestR_BITS_191_TO_128__q1[31],
		 IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d37 } :
	       IF_NOT_IF_IF_requestR_3_BIT_214_4_THEN_request_ETC___d2122 ;
  assign IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3__ETC___d2125 =
	     (sV2_exp__h1597 == 8'd255 && sV2_sfd__h1598[22]) ?
	       { requestR_BITS_191_TO_128__q1[63:32] == 32'hFFFFFFFF &&
		 requestR_BITS_191_TO_128__q1[31],
		 IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d37 } :
	       (IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2077 ?
		  IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d48 :
		  IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3__ETC___d2123) ;
  assign IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3__ETC___d2126 =
	     (sV1_exp__h1472 == 8'd255 && sV1_sfd__h1473[22]) ?
	       IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d48 :
	       IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3__ETC___d2125 ;
  assign IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3__ETC___d2128 =
	     (sV1_exp__h1472 == 8'd255 && sV1_sfd__h1473[22] &&
	      sV2_exp__h1597 == 8'd255 &&
	      sV2_sfd__h1598[22]) ?
	       64'hFFFFFFFF7FC00000 :
	       { 32'hFFFFFFFF,
		 IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3__ETC___d2126 } ;
  assign IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3__ETC___d2129 =
	     (sV2_exp__h1597 == 8'd255 && sV2_sfd__h1598 != 23'd0 &&
	      !sV2_sfd__h1598[22]) ?
	       res__h49096 :
	       IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3__ETC___d2128 ;
  assign IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3__ETC___d2130 =
	     (sV1_exp__h1472 == 8'd255 && sV1_sfd__h1473 != 23'd0 &&
	      !sV1_sfd__h1473[22]) ?
	       res__h48859 :
	       IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3__ETC___d2129 ;
  assign IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3__ETC___d2206 =
	     (sV1_exp__h1472 == 8'd0 && sV1_sfd__h1473 == 23'd0) ?
	       res___1__h57780 :
	       ((sV1_exp__h1472 == 8'd0) ? res___1__h57799 : res__h57815) ;
  assign IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3__ETC___d2207 =
	     (sV1_exp__h1472 == 8'd255 && sV1_sfd__h1473 == 23'd0) ?
	       res___1__h57770 :
	       IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3__ETC___d2206 ;
  assign IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3__ETC___d2339 =
	     sfd__h28849[31] ?
	       6'd0 :
	       (sfd__h28849[30] ?
		  6'd1 :
		  (sfd__h28849[29] ?
		     6'd2 :
		     (sfd__h28849[28] ?
			6'd3 :
			(sfd__h28849[27] ?
			   6'd4 :
			   (sfd__h28849[26] ?
			      6'd5 :
			      (sfd__h28849[25] ?
				 6'd6 :
				 (sfd__h28849[24] ?
				    6'd7 :
				    (sfd__h28849[23] ?
				       6'd8 :
				       (sfd__h28849[22] ?
					  6'd9 :
					  (sfd__h28849[21] ?
					     6'd10 :
					     (sfd__h28849[20] ?
						6'd11 :
						(sfd__h28849[19] ?
						   6'd12 :
						   (sfd__h28849[18] ?
						      6'd13 :
						      (sfd__h28849[17] ?
							 6'd14 :
							 (sfd__h28849[16] ?
							    6'd15 :
							    (sfd__h28849[15] ?
							       6'd16 :
							       (sfd__h28849[14] ?
								  6'd17 :
								  (sfd__h28849[13] ?
								     6'd18 :
								     (sfd__h28849[12] ?
									6'd19 :
									(sfd__h28849[11] ?
									   6'd20 :
									   (sfd__h28849[10] ?
									      6'd21 :
									      (sfd__h28849[9] ?
										 6'd22 :
										 (sfd__h28849[8] ?
										    6'd23 :
										    (sfd__h28849[7] ?
										       6'd24 :
										       (sfd__h28849[6] ?
											  6'd25 :
											  (sfd__h28849[5] ?
											     6'd26 :
											     (sfd__h28849[4] ?
												6'd27 :
												(sfd__h28849[3] ?
												   6'd28 :
												   (sfd__h28849[2] ?
												      6'd29 :
												      (sfd__h28849[1] ?
													 6'd30 :
													 (sfd__h28849[0] ?
													    6'd31 :
													    6'd55))))))))))))))))))))))))))))))) ;
  assign IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3__ETC___d441 =
	     sfd__h3990[63] ?
	       7'd0 :
	       (sfd__h3990[62] ?
		  7'd1 :
		  (sfd__h3990[61] ?
		     7'd2 :
		     (sfd__h3990[60] ?
			7'd3 :
			(sfd__h3990[59] ?
			   7'd4 :
			   (sfd__h3990[58] ?
			      7'd5 :
			      (sfd__h3990[57] ?
				 7'd6 :
				 (sfd__h3990[56] ?
				    7'd7 :
				    (sfd__h3990[55] ?
				       7'd8 :
				       (sfd__h3990[54] ?
					  7'd9 :
					  (sfd__h3990[53] ?
					     7'd10 :
					     (sfd__h3990[52] ?
						7'd11 :
						(sfd__h3990[51] ?
						   7'd12 :
						   (sfd__h3990[50] ?
						      7'd13 :
						      (sfd__h3990[49] ?
							 7'd14 :
							 (sfd__h3990[48] ?
							    7'd15 :
							    (sfd__h3990[47] ?
							       7'd16 :
							       (sfd__h3990[46] ?
								  7'd17 :
								  (sfd__h3990[45] ?
								     7'd18 :
								     (sfd__h3990[44] ?
									7'd19 :
									(sfd__h3990[43] ?
									   7'd20 :
									   (sfd__h3990[42] ?
									      7'd21 :
									      (sfd__h3990[41] ?
										 7'd22 :
										 (sfd__h3990[40] ?
										    7'd23 :
										    (sfd__h3990[39] ?
										       7'd24 :
										       (sfd__h3990[38] ?
											  7'd25 :
											  (sfd__h3990[37] ?
											     7'd26 :
											     (sfd__h3990[36] ?
												7'd27 :
												(sfd__h3990[35] ?
												   7'd28 :
												   (sfd__h3990[34] ?
												      7'd29 :
												      (sfd__h3990[33] ?
													 7'd30 :
													 (sfd__h3990[32] ?
													    7'd31 :
													    (sfd__h3990[31] ?
													       7'd32 :
													       (sfd__h3990[30] ?
														  7'd33 :
														  (sfd__h3990[29] ?
														     7'd34 :
														     (sfd__h3990[28] ?
															7'd35 :
															(sfd__h3990[27] ?
															   7'd36 :
															   (sfd__h3990[26] ?
															      7'd37 :
															      (sfd__h3990[25] ?
																 7'd38 :
																 (sfd__h3990[24] ?
																    7'd39 :
																    (sfd__h3990[23] ?
																       7'd40 :
																       (sfd__h3990[22] ?
																	  7'd41 :
																	  (sfd__h3990[21] ?
																	     7'd42 :
																	     (sfd__h3990[20] ?
																		7'd43 :
																		(sfd__h3990[19] ?
																		   7'd44 :
																		   (sfd__h3990[18] ?
																		      7'd45 :
																		      (sfd__h3990[17] ?
																			 7'd46 :
																			 (sfd__h3990[16] ?
																			    7'd47 :
																			    (sfd__h3990[15] ?
																			       7'd48 :
																			       (sfd__h3990[14] ?
																				  7'd49 :
																				  (sfd__h3990[13] ?
																				     7'd50 :
																				     (sfd__h3990[12] ?
																					7'd51 :
																					(sfd__h3990[11] ?
																					   7'd52 :
																					   (sfd__h3990[10] ?
																					      7'd53 :
																					      (sfd__h3990[9] ?
																						 7'd54 :
																						 (sfd__h3990[8] ?
																						    7'd55 :
																						    (sfd__h3990[7] ?
																						       7'd56 :
																						       (sfd__h3990[6] ?
																							  7'd57 :
																							  (sfd__h3990[5] ?
																							     7'd58 :
																							     (sfd__h3990[4] ?
																								7'd59 :
																								(sfd__h3990[3] ?
																								   7'd60 :
																								   (sfd__h3990[2] ?
																								      7'd61 :
																								      (sfd__h3990[1] ?
																									 7'd62 :
																									 (sfd__h3990[0] ?
																									    7'd63 :
																									    7'd64))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) ;
  assign IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3__ETC___d4613 =
	     ((sV1_exp__h1472 == 8'd0) ?
		(sV1_sfd__h1473[22] ?
		   6'd2 :
		   (sV1_sfd__h1473[21] ?
		      6'd3 :
		      (sV1_sfd__h1473[20] ?
			 6'd4 :
			 (sV1_sfd__h1473[19] ?
			    6'd5 :
			    (sV1_sfd__h1473[18] ?
			       6'd6 :
			       (sV1_sfd__h1473[17] ?
				  6'd7 :
				  (sV1_sfd__h1473[16] ?
				     6'd8 :
				     (sV1_sfd__h1473[15] ?
					6'd9 :
					(sV1_sfd__h1473[14] ?
					   6'd10 :
					   (sV1_sfd__h1473[13] ?
					      6'd11 :
					      (sV1_sfd__h1473[12] ?
						 6'd12 :
						 (sV1_sfd__h1473[11] ?
						    6'd13 :
						    (sV1_sfd__h1473[10] ?
						       6'd14 :
						       (sV1_sfd__h1473[9] ?
							  6'd15 :
							  (sV1_sfd__h1473[8] ?
							     6'd16 :
							     (sV1_sfd__h1473[7] ?
								6'd17 :
								(sV1_sfd__h1473[6] ?
								   6'd18 :
								   (sV1_sfd__h1473[5] ?
								      6'd19 :
								      (sV1_sfd__h1473[4] ?
									 6'd20 :
									 (sV1_sfd__h1473[3] ?
									    6'd21 :
									    (sV1_sfd__h1473[2] ?
									       6'd22 :
									       (sV1_sfd__h1473[1] ?
										  6'd23 :
										  (sV1_sfd__h1473[0] ?
										     6'd24 :
										     6'd57))))))))))))))))))))))) :
		6'd1) -
	     6'd1 ;
  assign IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3__ETC___d5153 =
	     (sV1_exp__h1472 == 8'd255 && sV1_sfd__h1473 != 23'd0) ?
	       _theResult___snd_fst_sfd__h169840 :
	       _theResult___fst_sfd__h212195 ;
  assign IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3__ETC___d5188 =
	     (sV1_exp__h1472 == 8'd0) ?
	       IF_NOT_3970_MINUS_0_CONCAT_IF_IF_IF_requestR_3_ETC___d5169 :
	       (SEXT_IF_IF_requestR_3_BIT_214_4_THEN_requestR__ETC___d4685 ?
		  IF_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_reques_ETC___d5186 :
		  requestR_BITS_191_TO_128__q1[63:32] == 32'hFFFFFFFF &&
		  requestR_BITS_191_TO_128__q1[31]) ;
  assign IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3__ETC___d5189 =
	     (sV1_exp__h1472 == 8'd255 && sV1_sfd__h1473 != 23'd0 ||
	      (sV1_exp__h1472 == 8'd255 || sV1_exp__h1472 == 8'd0) &&
	      sV1_sfd__h1473 == 23'd0) ?
	       requestR_BITS_191_TO_128__q1[63:32] == 32'hFFFFFFFF &&
	       requestR_BITS_191_TO_128__q1[31] :
	       IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3__ETC___d5188 ;
  assign IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3__ETC___d5224 =
	     (sV1_exp__h1472 == 8'd0) ?
	       _3970_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_21_ETC___d4542 &&
	       !_3970_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_21_ETC___d4543 &&
	       _0_CONCAT_IF_IF_IF_requestR_3_BIT_214_4_THEN_re_ETC___d5203[4] :
	       SEXT_IF_IF_requestR_3_BIT_214_4_THEN_requestR__ETC___d4685 &&
	       SEXT_IF_IF_requestR_3_BIT_214_4_THEN_requestR__ETC___d4686 &&
	       _0_CONCAT_IF_IF_3074_MINUS_SEXT_IF_IF_requestR__ETC___d5220[4] ;
  assign IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3__ETC___d5227 =
	     (sV1_exp__h1472 == 8'd255 && sV1_sfd__h1473 != 23'd0) ?
	       sV1_exp__h1472 == 8'd255 && sV1_sfd__h1473 != 23'd0 &&
	       !sV1_sfd__h1473[22] :
	       (sV1_exp__h1472 != 8'd255 || sV1_sfd__h1473 != 23'd0) &&
	       (sV1_exp__h1472 != 8'd0 || sV1_sfd__h1473 != 23'd0) &&
	       IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3__ETC___d5224 ;
  assign IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3__ETC___d5234 =
	     (sV1_exp__h1472 == 8'd0) ?
	       _3970_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_21_ETC___d4542 &&
	       !_3970_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_21_ETC___d4543 &&
	       _0_CONCAT_IF_IF_IF_requestR_3_BIT_214_4_THEN_re_ETC___d5203[3] :
	       SEXT_IF_IF_requestR_3_BIT_214_4_THEN_requestR__ETC___d4685 &&
	       SEXT_IF_IF_requestR_3_BIT_214_4_THEN_requestR__ETC___d4686 &&
	       _0_CONCAT_IF_IF_3074_MINUS_SEXT_IF_IF_requestR__ETC___d5220[3] ;
  assign IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3__ETC___d5248 =
	     (sV1_exp__h1472 == 8'd0) ?
	       !_3970_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_21_ETC___d4542 ||
	       !_3970_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_21_ETC___d4543 &&
	       _0_CONCAT_IF_IF_IF_requestR_3_BIT_214_4_THEN_re_ETC___d5203[2] :
	       !SEXT_IF_IF_requestR_3_BIT_214_4_THEN_requestR__ETC___d4685 ||
	       IF_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_reques_ETC___d5246 ;
  assign IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3__ETC___d5260 =
	     (sV1_exp__h1472 == 8'd0) ?
	       _3970_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_21_ETC___d4542 &&
	       (_3970_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_21_ETC___d4543 ||
		_0_CONCAT_IF_IF_IF_requestR_3_BIT_214_4_THEN_re_ETC___d5203[1]) :
	       SEXT_IF_IF_requestR_3_BIT_214_4_THEN_requestR__ETC___d4685 &&
	       IF_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_reques_ETC___d5258 ;
  assign IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3__ETC___d5272 =
	     (sV1_exp__h1472 == 8'd0) ?
	       !_3970_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_21_ETC___d4542 ||
	       !_3970_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_21_ETC___d4543 &&
	       _0_CONCAT_IF_IF_IF_requestR_3_BIT_214_4_THEN_re_ETC___d5203[0] :
	       !SEXT_IF_IF_requestR_3_BIT_214_4_THEN_requestR__ETC___d4685 ||
	       IF_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_reques_ETC___d5270 ;
  assign IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1439 =
	     (requestR_BITS_191_TO_128__q1[31:0] == 32'd0 ||
	      !sfd__h28849[31] && !sfd__h28849[30] && !sfd__h28849[29] &&
	      !sfd__h28849[28] &&
	      !sfd__h28849[27] &&
	      !sfd__h28849[26] &&
	      !sfd__h28849[25] &&
	      !sfd__h28849[24] &&
	      !sfd__h28849[23] &&
	      !sfd__h28849[22] &&
	      !sfd__h28849[21] &&
	      !sfd__h28849[20] &&
	      !sfd__h28849[19] &&
	      !sfd__h28849[18] &&
	      !sfd__h28849[17] &&
	      !sfd__h28849[16] &&
	      !sfd__h28849[15] &&
	      !sfd__h28849[14] &&
	      !sfd__h28849[13] &&
	      !sfd__h28849[12] &&
	      !sfd__h28849[11] &&
	      !sfd__h28849[10] &&
	      !sfd__h28849[9] &&
	      !sfd__h28849[8] &&
	      !sfd__h28849[7] &&
	      !sfd__h28849[6] &&
	      !sfd__h28849[5] &&
	      !sfd__h28849[4] &&
	      !sfd__h28849[3] &&
	      !sfd__h28849[2] &&
	      !sfd__h28849[1] &&
	      !sfd__h28849[0]) ?
	       8'd0 :
	       _theResult___snd_fst_exp__h35543 ;
  assign IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1520 =
	     (sfd__h28849[31] || sfd__h28849[30] || sfd__h28849[29] ||
	      sfd__h28849[28] ||
	      sfd__h28849[27] ||
	      sfd__h28849[26] ||
	      sfd__h28849[25] ||
	      sfd__h28849[24] ||
	      sfd__h28849[23] ||
	      sfd__h28849[22] ||
	      sfd__h28849[21] ||
	      sfd__h28849[20] ||
	      sfd__h28849[19] ||
	      sfd__h28849[18] ||
	      sfd__h28849[17] ||
	      sfd__h28849[16] ||
	      sfd__h28849[15] ||
	      sfd__h28849[14] ||
	      sfd__h28849[13] ||
	      sfd__h28849[12] ||
	      sfd__h28849[11] ||
	      sfd__h28849[10] ||
	      sfd__h28849[9] ||
	      sfd__h28849[8] ||
	      sfd__h28849[7] ||
	      sfd__h28849[6] ||
	      sfd__h28849[5] ||
	      sfd__h28849[4] ||
	      sfd__h28849[3] ||
	      sfd__h28849[2] ||
	      sfd__h28849[1] ||
	      sfd__h28849[0]) &&
	     (!_32_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d1322 ||
	      !_32_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d1324 &&
	      !_32_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d1327 &&
	      _theResult___fst_exp__h35534 == 8'd255 &&
	      _theResult___fst_sfd__h35535 == 23'd0) ;
  assign IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1523 =
	     (sfd__h28849[31] || sfd__h28849[30] || sfd__h28849[29] ||
	      sfd__h28849[28] ||
	      sfd__h28849[27] ||
	      sfd__h28849[26] ||
	      sfd__h28849[25] ||
	      sfd__h28849[24] ||
	      sfd__h28849[23] ||
	      sfd__h28849[22] ||
	      sfd__h28849[21] ||
	      sfd__h28849[20] ||
	      sfd__h28849[19] ||
	      sfd__h28849[18] ||
	      sfd__h28849[17] ||
	      sfd__h28849[16] ||
	      sfd__h28849[15] ||
	      sfd__h28849[14] ||
	      sfd__h28849[13] ||
	      sfd__h28849[12] ||
	      sfd__h28849[11] ||
	      sfd__h28849[10] ||
	      sfd__h28849[9] ||
	      sfd__h28849[8] ||
	      sfd__h28849[7] ||
	      sfd__h28849[6] ||
	      sfd__h28849[5] ||
	      sfd__h28849[4] ||
	      sfd__h28849[3] ||
	      sfd__h28849[2] ||
	      sfd__h28849[1] ||
	      sfd__h28849[0]) &&
	     _32_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d1322 &&
	     _32_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d1324 ;
  assign IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1532 =
	     (sfd__h28849[31] || sfd__h28849[30] || sfd__h28849[29] ||
	      sfd__h28849[28] ||
	      sfd__h28849[27] ||
	      sfd__h28849[26] ||
	      sfd__h28849[25] ||
	      sfd__h28849[24] ||
	      sfd__h28849[23] ||
	      sfd__h28849[22] ||
	      sfd__h28849[21] ||
	      sfd__h28849[20] ||
	      sfd__h28849[19] ||
	      sfd__h28849[18] ||
	      sfd__h28849[17] ||
	      sfd__h28849[16] ||
	      sfd__h28849[15] ||
	      sfd__h28849[14] ||
	      sfd__h28849[13] ||
	      sfd__h28849[12] ||
	      sfd__h28849[11] ||
	      sfd__h28849[10] ||
	      sfd__h28849[9] ||
	      sfd__h28849[8] ||
	      sfd__h28849[7] ||
	      sfd__h28849[6] ||
	      sfd__h28849[5] ||
	      sfd__h28849[4] ||
	      sfd__h28849[3] ||
	      sfd__h28849[2] ||
	      sfd__h28849[1] ||
	      sfd__h28849[0]) &&
	     _32_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d1322 &&
	     !_32_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d1324 &&
	     IF_32_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_2_ETC___d1529 ;
  assign IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1574 =
	     requestR_BITS_191_TO_128__q1[31] ?
	       6'd0 :
	       (requestR_BITS_191_TO_128__q1[30] ?
		  6'd1 :
		  (requestR_BITS_191_TO_128__q1[29] ?
		     6'd2 :
		     (requestR_BITS_191_TO_128__q1[28] ?
			6'd3 :
			(requestR_BITS_191_TO_128__q1[27] ?
			   6'd4 :
			   (requestR_BITS_191_TO_128__q1[26] ?
			      6'd5 :
			      (requestR_BITS_191_TO_128__q1[25] ?
				 6'd6 :
				 (requestR_BITS_191_TO_128__q1[24] ?
				    6'd7 :
				    (requestR_BITS_191_TO_128__q1[23] ?
				       6'd8 :
				       (requestR_BITS_191_TO_128__q1[22] ?
					  6'd9 :
					  (requestR_BITS_191_TO_128__q1[21] ?
					     6'd10 :
					     (requestR_BITS_191_TO_128__q1[20] ?
						6'd11 :
						(requestR_BITS_191_TO_128__q1[19] ?
						   6'd12 :
						   (requestR_BITS_191_TO_128__q1[18] ?
						      6'd13 :
						      (requestR_BITS_191_TO_128__q1[17] ?
							 6'd14 :
							 (requestR_BITS_191_TO_128__q1[16] ?
							    6'd15 :
							    (requestR_BITS_191_TO_128__q1[15] ?
							       6'd16 :
							       (requestR_BITS_191_TO_128__q1[14] ?
								  6'd17 :
								  (requestR_BITS_191_TO_128__q1[13] ?
								     6'd18 :
								     (requestR_BITS_191_TO_128__q1[12] ?
									6'd19 :
									(requestR_BITS_191_TO_128__q1[11] ?
									   6'd20 :
									   (requestR_BITS_191_TO_128__q1[10] ?
									      6'd21 :
									      (requestR_BITS_191_TO_128__q1[9] ?
										 6'd22 :
										 (requestR_BITS_191_TO_128__q1[8] ?
										    6'd23 :
										    (requestR_BITS_191_TO_128__q1[7] ?
										       6'd24 :
										       (requestR_BITS_191_TO_128__q1[6] ?
											  6'd25 :
											  (requestR_BITS_191_TO_128__q1[5] ?
											     6'd26 :
											     (requestR_BITS_191_TO_128__q1[4] ?
												6'd27 :
												(requestR_BITS_191_TO_128__q1[3] ?
												   6'd28 :
												   (requestR_BITS_191_TO_128__q1[2] ?
												      6'd29 :
												      (requestR_BITS_191_TO_128__q1[1] ?
													 6'd30 :
													 (requestR_BITS_191_TO_128__q1[0] ?
													    6'd31 :
													    6'd32))))))))))))))))))))))))))))))) ;
  assign IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1745 =
	     (requestR_BITS_191_TO_128__q1[63:32] == 32'hFFFFFFFF &&
	      requestR_BITS_191_TO_128__q1[31]) ?
	       64'h8000000000000000 :
	       64'h7FFFFFFFFFFFFFFF ;
  assign IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1748 =
	     sV1_exp__h1472 - 8'd127 ;
  assign IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1757 =
	     (requestR_BITS_191_TO_128__q1[63:32] == 32'hFFFFFFFF &&
	      requestR_BITS_191_TO_128__q1[31]) ?
	       -b__h43158 :
	       b__h43158 ;
  assign IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1774 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       ((guard__h43091 == 2'b10) ?
		  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1757[24] :
		  guard__h43091 == 2'b11) :
	       ((requestR[194:192] == 3'h3) ?
		  guard__h43091 != 2'd0 :
		  requestR[194:192] == 3'h1 &&
		  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1757[88] &&
		  guard__h43091 != 2'd0) ;
  assign IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1806 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       ((guard__h43869 == 2'b10) ?
		  x__h44058[25] :
		  guard__h43869 == 2'b11) :
	       ((requestR[194:192] == 3'h3) ?
		  guard__h43869 != 2'd0 :
		  requestR[194:192] == 3'h1 && x__h44058[88] &&
		  guard__h43869 != 2'd0) ;
  assign IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1868 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       ((guard__h45193 == 2'b10) ?
		  x__h45414[25] :
		  guard__h45193 == 2'b11) :
	       requestR[194:192] == 3'h3 && guard__h45193 != 2'd0 ;
  assign IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1878 =
	     (requestR_BITS_191_TO_128__q1[63:32] == 32'hFFFFFFFF &&
	      requestR_BITS_191_TO_128__q1[31]) ?
	       64'd0 :
	       ((sV1_exp__h1472 == 8'd255 && sV1_sfd__h1473 == 23'd0) ?
		  64'hFFFFFFFFFFFFFFFF :
		  IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3__ETC___d1876) ;
  assign IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1885 =
	     sV1_exp__h1472 == 8'd255 && sV1_sfd__h1473 != 23'd0 ||
	     sV1_exp__h1472 == 8'd255 && sV1_sfd__h1473 == 23'd0 ||
	     (sV1_exp__h1472 != 8'd0 || sV1_sfd__h1473 != 23'd0) &&
	     (NEG_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d1847[19] ||
	      NEG_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d1849 &&
	      IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1868 &&
	      x__h45414[88:25] == 64'hFFFFFFFFFFFFFFFF) ;
  assign IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1896 =
	     { IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1885,
	       3'd0,
	       (sV1_exp__h1472 != 8'd255 || sV1_sfd__h1473 == 23'd0) &&
	       (sV1_exp__h1472 != 8'd255 || sV1_sfd__h1473 != 23'd0) &&
	       NOT_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_ETC___d1890 } ==
	     5'd0 ||
	     IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1885 ;
  assign IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1904 =
	     (requestR_BITS_191_TO_128__q1[63:32] == 32'hFFFFFFFF &&
	      requestR_BITS_191_TO_128__q1[31]) ?
	       32'h80000000 :
	       32'h7FFFFFFF ;
  assign IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1908 =
	     (requestR_BITS_191_TO_128__q1[63:32] == 32'hFFFFFFFF &&
	      requestR_BITS_191_TO_128__q1[31]) ?
	       -b__h46021 :
	       b__h46021 ;
  assign IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1925 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       ((guard__h45954 == 2'b10) ?
		  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1908[24] :
		  guard__h45954 == 2'b11) :
	       ((requestR[194:192] == 3'h3) ?
		  guard__h45954 != 2'd0 :
		  requestR[194:192] == 3'h1 &&
		  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1908[56] &&
		  guard__h45954 != 2'd0) ;
  assign IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1957 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       ((guard__h46508 == 2'b10) ?
		  x__h46697[25] :
		  guard__h46508 == 2'b11) :
	       ((requestR[194:192] == 3'h3) ?
		  guard__h46508 != 2'd0 :
		  requestR[194:192] == 3'h1 && x__h46697[56] &&
		  guard__h46508 != 2'd0) ;
  assign IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2014 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       ((guard__h47594 == 2'b10) ?
		  x__h47815[25] :
		  guard__h47594 == 2'b11) :
	       requestR[194:192] == 3'h3 && guard__h47594 != 2'd0 ;
  assign IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2024 =
	     (requestR_BITS_191_TO_128__q1[63:32] == 32'hFFFFFFFF &&
	      requestR_BITS_191_TO_128__q1[31]) ?
	       32'd0 :
	       ((sV1_exp__h1472 == 8'd255 && sV1_sfd__h1473 == 23'd0) ?
		  32'hFFFFFFFF :
		  IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3__ETC___d2022) ;
  assign IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2032 =
	     sV1_exp__h1472 == 8'd255 && sV1_sfd__h1473 != 23'd0 ||
	     sV1_exp__h1472 == 8'd255 && sV1_sfd__h1473 == 23'd0 ||
	     (sV1_exp__h1472 != 8'd0 || sV1_sfd__h1473 != 23'd0) &&
	     (NEG_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d1993[19] ||
	      NEG_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d1995 &&
	      IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2014 &&
	      x__h47815[56:25] == 32'hFFFFFFFF) ;
  assign IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2043 =
	     { IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2032,
	       3'd0,
	       (sV1_exp__h1472 != 8'd255 || sV1_sfd__h1473 == 23'd0) &&
	       (sV1_exp__h1472 != 8'd255 || sV1_sfd__h1473 != 23'd0) &&
	       NOT_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_ETC___d2037 } ==
	     5'd0 ||
	     IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2032 ;
  assign IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2067 =
	     sV1_exp__h1472 == 8'd255 && sV1_sfd__h1473 != 23'd0 &&
	     !sV1_sfd__h1473[22] &&
	     sV2_exp__h1597 == 8'd255 &&
	     sV2_sfd__h1598 != 23'd0 &&
	     !sV2_sfd__h1598[22] ;
  assign IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2077 =
	     sV1_exp__h1472 == 8'd0 && sV1_sfd__h1473 == 23'd0 &&
	     requestR_BITS_191_TO_128__q1[63:32] == 32'hFFFFFFFF &&
	     requestR_BITS_191_TO_128__q1[31] &&
	     sV2_exp__h1597 == 8'd0 &&
	     sV2_sfd__h1598 == 23'd0 &&
	     (requestR_BITS_127_TO_64__q3[63:32] != 32'hFFFFFFFF ||
	      !requestR_BITS_127_TO_64__q3[31]) ;
  assign IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2081 =
	     sV2_exp__h1597 == 8'd0 && sV2_sfd__h1598 == 23'd0 &&
	     requestR_BITS_127_TO_64__q3[63:32] == 32'hFFFFFFFF &&
	     requestR_BITS_127_TO_64__q3[31] &&
	     sV1_exp__h1472 == 8'd0 &&
	     sV1_sfd__h1473 == 23'd0 &&
	     (requestR_BITS_191_TO_128__q1[63:32] != 32'hFFFFFFFF ||
	      !requestR_BITS_191_TO_128__q1[31]) ;
  assign IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2090 =
	     sV1_exp__h1472 < sV2_exp__h1597 ;
  assign IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2091 =
	     sV1_exp__h1472 == sV2_exp__h1597 ;
  assign IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2092 =
	     sV1_sfd__h1473 < sV2_sfd__h1598 ;
  assign IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2095 =
	     sV1_exp__h1472 <= sV2_exp__h1597 ;
  assign IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2097 =
	     sV1_sfd__h1473 <= sV2_sfd__h1598 ;
  assign IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2115 =
	     sV1_exp__h1472 == 8'd255 && sV1_sfd__h1473 != 23'd0 &&
	     !sV1_sfd__h1473[22] ||
	     sV2_exp__h1597 == 8'd255 && sV2_sfd__h1598 != 23'd0 &&
	     !sV2_sfd__h1598[22] ;
  assign IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2156 =
	     IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2115 ||
	     sV1_exp__h1472 == 8'd255 && sV1_sfd__h1473[22] ||
	     sV2_exp__h1597 == 8'd255 && sV2_sfd__h1598[22] ;
  assign IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2167 =
	     IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2095 &&
	     (!IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2091 ||
	      IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2097) &&
	     !IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2090 &&
	     (!IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2091 ||
	      !IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2092) ;
  assign IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2171 =
	     sV1_exp__h1472 == 8'd0 && sV1_sfd__h1473 == 23'd0 &&
	     sV2_exp__h1597 == 8'd0 &&
	     sV2_sfd__h1598 == 23'd0 ||
	     (requestR_BITS_191_TO_128__q1[63:32] != 32'hFFFFFFFF ||
	      !requestR_BITS_191_TO_128__q1[31] ||
	      requestR_BITS_127_TO_64__q3[63:32] == 32'hFFFFFFFF &&
	      requestR_BITS_127_TO_64__q3[31]) &&
	     IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d2169 ;
  assign IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2496 =
	     (requestR_BITS_191_TO_128__q1[31:0] == 32'd0 ||
	      !_32_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d2343 ||
	      _32_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d2345) ?
	       52'd0 :
	       _theResult___snd_fst_sfd__h70875 ;
  assign IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2555 =
	     requestR_BITS_191_TO_128__q1[31] ?
	       6'd0 :
	       (requestR_BITS_191_TO_128__q1[30] ?
		  6'd1 :
		  (requestR_BITS_191_TO_128__q1[29] ?
		     6'd2 :
		     (requestR_BITS_191_TO_128__q1[28] ?
			6'd3 :
			(requestR_BITS_191_TO_128__q1[27] ?
			   6'd4 :
			   (requestR_BITS_191_TO_128__q1[26] ?
			      6'd5 :
			      (requestR_BITS_191_TO_128__q1[25] ?
				 6'd6 :
				 (requestR_BITS_191_TO_128__q1[24] ?
				    6'd7 :
				    (requestR_BITS_191_TO_128__q1[23] ?
				       6'd8 :
				       (requestR_BITS_191_TO_128__q1[22] ?
					  6'd9 :
					  (requestR_BITS_191_TO_128__q1[21] ?
					     6'd10 :
					     (requestR_BITS_191_TO_128__q1[20] ?
						6'd11 :
						(requestR_BITS_191_TO_128__q1[19] ?
						   6'd12 :
						   (requestR_BITS_191_TO_128__q1[18] ?
						      6'd13 :
						      (requestR_BITS_191_TO_128__q1[17] ?
							 6'd14 :
							 (requestR_BITS_191_TO_128__q1[16] ?
							    6'd15 :
							    (requestR_BITS_191_TO_128__q1[15] ?
							       6'd16 :
							       (requestR_BITS_191_TO_128__q1[14] ?
								  6'd17 :
								  (requestR_BITS_191_TO_128__q1[13] ?
								     6'd18 :
								     (requestR_BITS_191_TO_128__q1[12] ?
									6'd19 :
									(requestR_BITS_191_TO_128__q1[11] ?
									   6'd20 :
									   (requestR_BITS_191_TO_128__q1[10] ?
									      6'd21 :
									      (requestR_BITS_191_TO_128__q1[9] ?
										 6'd22 :
										 (requestR_BITS_191_TO_128__q1[8] ?
										    6'd23 :
										    (requestR_BITS_191_TO_128__q1[7] ?
										       6'd24 :
										       (requestR_BITS_191_TO_128__q1[6] ?
											  6'd25 :
											  (requestR_BITS_191_TO_128__q1[5] ?
											     6'd26 :
											     (requestR_BITS_191_TO_128__q1[4] ?
												6'd27 :
												(requestR_BITS_191_TO_128__q1[3] ?
												   6'd28 :
												   (requestR_BITS_191_TO_128__q1[2] ?
												      6'd29 :
												      (requestR_BITS_191_TO_128__q1[1] ?
													 6'd30 :
													 (requestR_BITS_191_TO_128__q1[0] ?
													    6'd31 :
													    6'd55))))))))))))))))))))))))))))))) ;
  assign IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2680 =
	     (requestR_BITS_191_TO_128__q1[31:0] == 32'd0 ||
	      !_32_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d2559 ||
	      _32_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d2560) ?
	       52'd0 :
	       _theResult___snd_fst_sfd__h81820 ;
  assign IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2719 =
	     requestR_BITS_191_TO_128__q1[63] ? 32'h80000000 : 32'h7FFFFFFF ;
  assign IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2731 =
	     requestR_BITS_191_TO_128__q1[63] ? -b__h82525 : b__h82525 ;
  assign IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2748 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       ((guard__h82458 == 2'b10) ?
		  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2731[53] :
		  guard__h82458 == 2'b11) :
	       ((requestR[194:192] == 3'h3) ?
		  guard__h82458 != 2'd0 :
		  requestR[194:192] == 3'h1 &&
		  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2731[85] &&
		  guard__h82458 != 2'd0) ;
  assign IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2780 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       ((guard__h83012 == 2'b10) ?
		  x__h83201[54] :
		  guard__h83012 == 2'b11) :
	       ((requestR[194:192] == 3'h3) ?
		  guard__h83012 != 2'd0 :
		  requestR[194:192] == 3'h1 && x__h83201[85] &&
		  guard__h83012 != 2'd0) ;
  assign IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2790 =
	     (requestR_BITS_191_TO_128__q1[62:52] == 11'd2047 &&
	      requestR_BITS_191_TO_128__q1[51:0] == 52'd0) ?
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2719 :
	       ((requestR_BITS_191_TO_128__q1[62:52] == 11'd0 &&
		 requestR_BITS_191_TO_128__q1[51:0] == 52'd0) ?
		  32'd0 :
		  IF_NEG_SEXT_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d2788) ;
  assign IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2843 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       ((guard__h84098 == 2'b10) ?
		  x__h84319[54] :
		  guard__h84098 == 2'b11) :
	       requestR[194:192] == 3'h3 && guard__h84098 != 2'd0 ;
  assign IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2851 =
	     (requestR_BITS_191_TO_128__q1[62:52] == 11'd0 &&
	      requestR_BITS_191_TO_128__q1[51:0] == 52'd0) ?
	       32'd0 :
	       (NEG_SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d2822[23] ?
		  32'hFFFFFFFF :
		  IF_NEG_SEXT_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d2849) ;
  assign IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2996 =
	     (requestR[191:128] == 64'd0 ||
	      !sfd__h3990[63] && !sfd__h3990[62] && !sfd__h3990[61] &&
	      !sfd__h3990[60] &&
	      !sfd__h3990[59] &&
	      !sfd__h3990[58] &&
	      !sfd__h3990[57] &&
	      !sfd__h3990[56] &&
	      !sfd__h3990[55] &&
	      !sfd__h3990[54] &&
	      !sfd__h3990[53] &&
	      !sfd__h3990[52] &&
	      !sfd__h3990[51] &&
	      !sfd__h3990[50] &&
	      !sfd__h3990[49] &&
	      !sfd__h3990[48] &&
	      !sfd__h3990[47] &&
	      !sfd__h3990[46] &&
	      !sfd__h3990[45] &&
	      !sfd__h3990[44] &&
	      !sfd__h3990[43] &&
	      !sfd__h3990[42] &&
	      !sfd__h3990[41] &&
	      !sfd__h3990[40] &&
	      !sfd__h3990[39] &&
	      !sfd__h3990[38] &&
	      !sfd__h3990[37] &&
	      !sfd__h3990[36] &&
	      !sfd__h3990[35] &&
	      !sfd__h3990[34] &&
	      !sfd__h3990[33] &&
	      !sfd__h3990[32] &&
	      !sfd__h3990[31] &&
	      !sfd__h3990[30] &&
	      !sfd__h3990[29] &&
	      !sfd__h3990[28] &&
	      !sfd__h3990[27] &&
	      !sfd__h3990[26] &&
	      !sfd__h3990[25] &&
	      !sfd__h3990[24] &&
	      !sfd__h3990[23] &&
	      !sfd__h3990[22] &&
	      !sfd__h3990[21] &&
	      !sfd__h3990[20] &&
	      !sfd__h3990[19] &&
	      !sfd__h3990[18] &&
	      !sfd__h3990[17] &&
	      !sfd__h3990[16] &&
	      !sfd__h3990[15] &&
	      !sfd__h3990[14] &&
	      !sfd__h3990[13] &&
	      !sfd__h3990[12] &&
	      !sfd__h3990[11] &&
	      !sfd__h3990[10] &&
	      !sfd__h3990[9] &&
	      !sfd__h3990[8] &&
	      !sfd__h3990[7] &&
	      !sfd__h3990[6] &&
	      !sfd__h3990[5] &&
	      !sfd__h3990[4] &&
	      !sfd__h3990[3] &&
	      !sfd__h3990[2] &&
	      !sfd__h3990[1] &&
	      !sfd__h3990[0]) ?
	       11'd0 :
	       _theResult___snd_fst_exp__h97202 ;
  assign IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d3045 =
	     (sfd__h3990[63] || sfd__h3990[62] || sfd__h3990[61] ||
	      sfd__h3990[60] ||
	      sfd__h3990[59] ||
	      sfd__h3990[58] ||
	      sfd__h3990[57] ||
	      sfd__h3990[56] ||
	      sfd__h3990[55] ||
	      sfd__h3990[54] ||
	      sfd__h3990[53] ||
	      sfd__h3990[52] ||
	      sfd__h3990[51] ||
	      sfd__h3990[50] ||
	      sfd__h3990[49] ||
	      sfd__h3990[48] ||
	      sfd__h3990[47] ||
	      sfd__h3990[46] ||
	      sfd__h3990[45] ||
	      sfd__h3990[44] ||
	      sfd__h3990[43] ||
	      sfd__h3990[42] ||
	      sfd__h3990[41] ||
	      sfd__h3990[40] ||
	      sfd__h3990[39] ||
	      sfd__h3990[38] ||
	      sfd__h3990[37] ||
	      sfd__h3990[36] ||
	      sfd__h3990[35] ||
	      sfd__h3990[34] ||
	      sfd__h3990[33] ||
	      sfd__h3990[32] ||
	      sfd__h3990[31] ||
	      sfd__h3990[30] ||
	      sfd__h3990[29] ||
	      sfd__h3990[28] ||
	      sfd__h3990[27] ||
	      sfd__h3990[26] ||
	      sfd__h3990[25] ||
	      sfd__h3990[24] ||
	      sfd__h3990[23] ||
	      sfd__h3990[22] ||
	      sfd__h3990[21] ||
	      sfd__h3990[20] ||
	      sfd__h3990[19] ||
	      sfd__h3990[18] ||
	      sfd__h3990[17] ||
	      sfd__h3990[16] ||
	      sfd__h3990[15] ||
	      sfd__h3990[14] ||
	      sfd__h3990[13] ||
	      sfd__h3990[12] ||
	      sfd__h3990[11] ||
	      sfd__h3990[10] ||
	      sfd__h3990[9] ||
	      sfd__h3990[8] ||
	      sfd__h3990[7] ||
	      sfd__h3990[6] ||
	      sfd__h3990[5] ||
	      sfd__h3990[4] ||
	      sfd__h3990[3] ||
	      sfd__h3990[2] ||
	      sfd__h3990[1] ||
	      sfd__h3990[0]) &&
	     (!_64_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d2883 ||
	      !_64_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d2885 &&
	      !_64_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d2888 &&
	      _theResult___fst_exp__h97193 == 11'd2047 &&
	      _theResult___fst_sfd__h97194 == 52'd0) ;
  assign IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d3048 =
	     (sfd__h3990[63] || sfd__h3990[62] || sfd__h3990[61] ||
	      sfd__h3990[60] ||
	      sfd__h3990[59] ||
	      sfd__h3990[58] ||
	      sfd__h3990[57] ||
	      sfd__h3990[56] ||
	      sfd__h3990[55] ||
	      sfd__h3990[54] ||
	      sfd__h3990[53] ||
	      sfd__h3990[52] ||
	      sfd__h3990[51] ||
	      sfd__h3990[50] ||
	      sfd__h3990[49] ||
	      sfd__h3990[48] ||
	      sfd__h3990[47] ||
	      sfd__h3990[46] ||
	      sfd__h3990[45] ||
	      sfd__h3990[44] ||
	      sfd__h3990[43] ||
	      sfd__h3990[42] ||
	      sfd__h3990[41] ||
	      sfd__h3990[40] ||
	      sfd__h3990[39] ||
	      sfd__h3990[38] ||
	      sfd__h3990[37] ||
	      sfd__h3990[36] ||
	      sfd__h3990[35] ||
	      sfd__h3990[34] ||
	      sfd__h3990[33] ||
	      sfd__h3990[32] ||
	      sfd__h3990[31] ||
	      sfd__h3990[30] ||
	      sfd__h3990[29] ||
	      sfd__h3990[28] ||
	      sfd__h3990[27] ||
	      sfd__h3990[26] ||
	      sfd__h3990[25] ||
	      sfd__h3990[24] ||
	      sfd__h3990[23] ||
	      sfd__h3990[22] ||
	      sfd__h3990[21] ||
	      sfd__h3990[20] ||
	      sfd__h3990[19] ||
	      sfd__h3990[18] ||
	      sfd__h3990[17] ||
	      sfd__h3990[16] ||
	      sfd__h3990[15] ||
	      sfd__h3990[14] ||
	      sfd__h3990[13] ||
	      sfd__h3990[12] ||
	      sfd__h3990[11] ||
	      sfd__h3990[10] ||
	      sfd__h3990[9] ||
	      sfd__h3990[8] ||
	      sfd__h3990[7] ||
	      sfd__h3990[6] ||
	      sfd__h3990[5] ||
	      sfd__h3990[4] ||
	      sfd__h3990[3] ||
	      sfd__h3990[2] ||
	      sfd__h3990[1] ||
	      sfd__h3990[0]) &&
	     _64_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d2883 &&
	     _64_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d2885 ;
  assign IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d3057 =
	     (sfd__h3990[63] || sfd__h3990[62] || sfd__h3990[61] ||
	      sfd__h3990[60] ||
	      sfd__h3990[59] ||
	      sfd__h3990[58] ||
	      sfd__h3990[57] ||
	      sfd__h3990[56] ||
	      sfd__h3990[55] ||
	      sfd__h3990[54] ||
	      sfd__h3990[53] ||
	      sfd__h3990[52] ||
	      sfd__h3990[51] ||
	      sfd__h3990[50] ||
	      sfd__h3990[49] ||
	      sfd__h3990[48] ||
	      sfd__h3990[47] ||
	      sfd__h3990[46] ||
	      sfd__h3990[45] ||
	      sfd__h3990[44] ||
	      sfd__h3990[43] ||
	      sfd__h3990[42] ||
	      sfd__h3990[41] ||
	      sfd__h3990[40] ||
	      sfd__h3990[39] ||
	      sfd__h3990[38] ||
	      sfd__h3990[37] ||
	      sfd__h3990[36] ||
	      sfd__h3990[35] ||
	      sfd__h3990[34] ||
	      sfd__h3990[33] ||
	      sfd__h3990[32] ||
	      sfd__h3990[31] ||
	      sfd__h3990[30] ||
	      sfd__h3990[29] ||
	      sfd__h3990[28] ||
	      sfd__h3990[27] ||
	      sfd__h3990[26] ||
	      sfd__h3990[25] ||
	      sfd__h3990[24] ||
	      sfd__h3990[23] ||
	      sfd__h3990[22] ||
	      sfd__h3990[21] ||
	      sfd__h3990[20] ||
	      sfd__h3990[19] ||
	      sfd__h3990[18] ||
	      sfd__h3990[17] ||
	      sfd__h3990[16] ||
	      sfd__h3990[15] ||
	      sfd__h3990[14] ||
	      sfd__h3990[13] ||
	      sfd__h3990[12] ||
	      sfd__h3990[11] ||
	      sfd__h3990[10] ||
	      sfd__h3990[9] ||
	      sfd__h3990[8] ||
	      sfd__h3990[7] ||
	      sfd__h3990[6] ||
	      sfd__h3990[5] ||
	      sfd__h3990[4] ||
	      sfd__h3990[3] ||
	      sfd__h3990[2] ||
	      sfd__h3990[1] ||
	      sfd__h3990[0]) &&
	     _64_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d2883 &&
	     !_64_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d2885 &&
	     IF_64_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_2_ETC___d3054 ;
  assign IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d3220 =
	     requestR_BITS_191_TO_128__q1[63] ?
	       64'h8000000000000000 :
	       64'h7FFFFFFFFFFFFFFF ;
  assign IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d3224 =
	     requestR_BITS_191_TO_128__q1[63] ? -b__h110422 : b__h110422 ;
  assign IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d3241 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       ((guard__h110355 == 2'b10) ?
		  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d3224[53] :
		  guard__h110355 == 2'b11) :
	       ((requestR[194:192] == 3'h3) ?
		  guard__h110355 != 2'd0 :
		  requestR[194:192] == 3'h1 &&
		  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d3224[117] &&
		  guard__h110355 != 2'd0) ;
  assign IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d3273 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       ((guard__h111133 == 2'b10) ?
		  x__h111322[54] :
		  guard__h111133 == 2'b11) :
	       ((requestR[194:192] == 3'h3) ?
		  guard__h111133 != 2'd0 :
		  requestR[194:192] == 3'h1 && x__h111322[117] &&
		  guard__h111133 != 2'd0) ;
  assign IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d3283 =
	     (requestR_BITS_191_TO_128__q1[62:52] == 11'd2047 &&
	      requestR_BITS_191_TO_128__q1[51:0] == 52'd0) ?
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d3220 :
	       ((requestR_BITS_191_TO_128__q1[62:52] == 11'd0 &&
		 requestR_BITS_191_TO_128__q1[51:0] == 52'd0) ?
		  64'd0 :
		  IF_NEG_SEXT_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d3281) ;
  assign IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d3329 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       ((guard__h112440 == 2'b10) ?
		  x__h112661[54] :
		  guard__h112440 == 2'b11) :
	       requestR[194:192] == 3'h3 && guard__h112440 != 2'd0 ;
  assign IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d3337 =
	     (requestR_BITS_191_TO_128__q1[62:52] == 11'd0 &&
	      requestR_BITS_191_TO_128__q1[51:0] == 52'd0) ?
	       64'd0 :
	       (NEG_SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d3308[23] ?
		  64'hFFFFFFFFFFFFFFFF :
		  IF_NEG_SEXT_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d3335) ;
  assign IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d37 =
	     (requestR_BITS_191_TO_128__q1[63:32] == 32'hFFFFFFFF) ?
	       requestR_BITS_191_TO_128__q1[30:0] :
	       31'h7FC00000 ;
  assign IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d3776 =
	     ((requestR_BITS_191_TO_128__q1[62:52] == 11'd0) ?
		(requestR_BITS_191_TO_128__q1[51] ?
		   6'd2 :
		   (requestR_BITS_191_TO_128__q1[50] ?
		      6'd3 :
		      (requestR_BITS_191_TO_128__q1[49] ?
			 6'd4 :
			 (requestR_BITS_191_TO_128__q1[48] ?
			    6'd5 :
			    (requestR_BITS_191_TO_128__q1[47] ?
			       6'd6 :
			       (requestR_BITS_191_TO_128__q1[46] ?
				  6'd7 :
				  (requestR_BITS_191_TO_128__q1[45] ?
				     6'd8 :
				     (requestR_BITS_191_TO_128__q1[44] ?
					6'd9 :
					(requestR_BITS_191_TO_128__q1[43] ?
					   6'd10 :
					   (requestR_BITS_191_TO_128__q1[42] ?
					      6'd11 :
					      (requestR_BITS_191_TO_128__q1[41] ?
						 6'd12 :
						 (requestR_BITS_191_TO_128__q1[40] ?
						    6'd13 :
						    (requestR_BITS_191_TO_128__q1[39] ?
						       6'd14 :
						       (requestR_BITS_191_TO_128__q1[38] ?
							  6'd15 :
							  (requestR_BITS_191_TO_128__q1[37] ?
							     6'd16 :
							     (requestR_BITS_191_TO_128__q1[36] ?
								6'd17 :
								(requestR_BITS_191_TO_128__q1[35] ?
								   6'd18 :
								   (requestR_BITS_191_TO_128__q1[34] ?
								      6'd19 :
								      (requestR_BITS_191_TO_128__q1[33] ?
									 6'd20 :
									 (requestR_BITS_191_TO_128__q1[32] ?
									    6'd21 :
									    (requestR_BITS_191_TO_128__q1[31] ?
									       6'd22 :
									       (requestR_BITS_191_TO_128__q1[30] ?
										  6'd23 :
										  (requestR_BITS_191_TO_128__q1[29] ?
										     6'd24 :
										     (requestR_BITS_191_TO_128__q1[28] ?
											6'd25 :
											(requestR_BITS_191_TO_128__q1[27] ?
											   6'd26 :
											   (requestR_BITS_191_TO_128__q1[26] ?
											      6'd27 :
											      (requestR_BITS_191_TO_128__q1[25] ?
												 6'd28 :
												 (requestR_BITS_191_TO_128__q1[24] ?
												    6'd29 :
												    (requestR_BITS_191_TO_128__q1[23] ?
												       6'd30 :
												       (requestR_BITS_191_TO_128__q1[22] ?
													  6'd31 :
													  (requestR_BITS_191_TO_128__q1[21] ?
													     6'd32 :
													     (requestR_BITS_191_TO_128__q1[20] ?
														6'd33 :
														(requestR_BITS_191_TO_128__q1[19] ?
														   6'd34 :
														   (requestR_BITS_191_TO_128__q1[18] ?
														      6'd35 :
														      (requestR_BITS_191_TO_128__q1[17] ?
															 6'd36 :
															 (requestR_BITS_191_TO_128__q1[16] ?
															    6'd37 :
															    (requestR_BITS_191_TO_128__q1[15] ?
															       6'd38 :
															       (requestR_BITS_191_TO_128__q1[14] ?
																  6'd39 :
																  (requestR_BITS_191_TO_128__q1[13] ?
																     6'd40 :
																     (requestR_BITS_191_TO_128__q1[12] ?
																	6'd41 :
																	(requestR_BITS_191_TO_128__q1[11] ?
																	   6'd42 :
																	   (requestR_BITS_191_TO_128__q1[10] ?
																	      6'd43 :
																	      (requestR_BITS_191_TO_128__q1[9] ?
																		 6'd44 :
																		 (requestR_BITS_191_TO_128__q1[8] ?
																		    6'd45 :
																		    (requestR_BITS_191_TO_128__q1[7] ?
																		       6'd46 :
																		       (requestR_BITS_191_TO_128__q1[6] ?
																			  6'd47 :
																			  (requestR_BITS_191_TO_128__q1[5] ?
																			     6'd48 :
																			     (requestR_BITS_191_TO_128__q1[4] ?
																				6'd49 :
																				(requestR_BITS_191_TO_128__q1[3] ?
																				   6'd50 :
																				   (requestR_BITS_191_TO_128__q1[2] ?
																				      6'd51 :
																				      (requestR_BITS_191_TO_128__q1[1] ?
																					 6'd52 :
																					 (requestR_BITS_191_TO_128__q1[0] ?
																					    6'd53 :
																					    6'd57)))))))))))))))))))))))))))))))))))))))))))))))))))) :
		6'd1) -
	     6'd1 ;
  assign IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d4338 =
	     (requestR_BITS_191_TO_128__q1[62:52] == 11'd2047 &&
	      requestR_BITS_191_TO_128__q1[51:0] != 52'd0) ?
	       _theResult___snd_fst_sfd__h117207 :
	       _theResult___fst_sfd__h166273 ;
  assign IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d4378 =
	     (requestR_BITS_191_TO_128__q1[62:52] == 11'd0) ?
	       (_3074_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_ETC___d3421 ?
		  IF_3074_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_21_ETC___d4358 :
		  requestR_BITS_191_TO_128__q1[63]) :
	       (SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_3_B_ETC___d3852 ?
		  IF_SEXT_IF_requestR_3_BIT_214_4_THEN_requestR__ETC___d4376 :
		  requestR_BITS_191_TO_128__q1[63]) ;
  assign IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d4429 =
	     (requestR_BITS_191_TO_128__q1[62:52] == 11'd0) ?
	       _3074_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_ETC___d4411 :
	       SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_3_B_ETC___d3852 &&
	       SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_3_B_ETC___d3853 &&
	       _0_CONCAT_IF_IF_3970_MINUS_SEXT_IF_requestR_3_B_ETC___d4425[4] ;
  assign IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d4440 =
	     (requestR_BITS_191_TO_128__q1[62:52] == 11'd0) ?
	       _3074_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_ETC___d4436 :
	       SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_3_B_ETC___d3852 &&
	       SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_3_B_ETC___d3853 &&
	       _0_CONCAT_IF_IF_3970_MINUS_SEXT_IF_requestR_3_B_ETC___d4425[3] ;
  assign IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d4456 =
	     (requestR_BITS_191_TO_128__q1[62:52] == 11'd0) ?
	       NOT_3074_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_2_ETC___d4448 :
	       !SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_3_B_ETC___d3852 ||
	       IF_SEXT_IF_requestR_3_BIT_214_4_THEN_requestR__ETC___d4454 ;
  assign IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d4469 =
	     (requestR_BITS_191_TO_128__q1[62:52] == 11'd0) ?
	       _3074_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_ETC___d4463 :
	       SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_3_B_ETC___d3852 &&
	       IF_SEXT_IF_requestR_3_BIT_214_4_THEN_requestR__ETC___d4467 ;
  assign IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d4482 =
	     (requestR_BITS_191_TO_128__q1[62:52] == 11'd0) ?
	       NOT_3074_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_2_ETC___d4476 :
	       !SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_3_B_ETC___d3852 ||
	       IF_SEXT_IF_requestR_3_BIT_214_4_THEN_requestR__ETC___d4480 ;
  assign IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d4617 =
	     sV1_exp__h1472 == 8'd0 && !sV1_sfd__h1473[22] &&
	     !sV1_sfd__h1473[21] &&
	     !sV1_sfd__h1473[20] &&
	     !sV1_sfd__h1473[19] &&
	     !sV1_sfd__h1473[18] &&
	     !sV1_sfd__h1473[17] &&
	     !sV1_sfd__h1473[16] &&
	     !sV1_sfd__h1473[15] &&
	     !sV1_sfd__h1473[14] &&
	     !sV1_sfd__h1473[13] &&
	     !sV1_sfd__h1473[12] &&
	     !sV1_sfd__h1473[11] &&
	     !sV1_sfd__h1473[10] &&
	     !sV1_sfd__h1473[9] &&
	     !sV1_sfd__h1473[8] &&
	     !sV1_sfd__h1473[7] &&
	     !sV1_sfd__h1473[6] &&
	     !sV1_sfd__h1473[5] &&
	     !sV1_sfd__h1473[4] &&
	     !sV1_sfd__h1473[3] &&
	     !sV1_sfd__h1473[2] &&
	     !sV1_sfd__h1473[1] &&
	     !sV1_sfd__h1473[0] ||
	     !_0_CONCAT_IF_IF_IF_requestR_3_BIT_214_4_THEN_re_ETC___d4615 ;
  assign IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d5010 =
	     sV1_exp__h1472 == 8'd0 && !sV1_sfd__h1473[22] &&
	     !sV1_sfd__h1473[21] &&
	     !sV1_sfd__h1473[20] &&
	     !sV1_sfd__h1473[19] &&
	     !sV1_sfd__h1473[18] &&
	     !sV1_sfd__h1473[17] &&
	     !sV1_sfd__h1473[16] &&
	     !sV1_sfd__h1473[15] &&
	     !sV1_sfd__h1473[14] &&
	     !sV1_sfd__h1473[13] &&
	     !sV1_sfd__h1473[12] &&
	     !sV1_sfd__h1473[11] &&
	     !sV1_sfd__h1473[10] &&
	     !sV1_sfd__h1473[9] &&
	     !sV1_sfd__h1473[8] &&
	     !sV1_sfd__h1473[7] &&
	     !sV1_sfd__h1473[6] &&
	     !sV1_sfd__h1473[5] &&
	     !sV1_sfd__h1473[4] &&
	     !sV1_sfd__h1473[3] &&
	     !sV1_sfd__h1473[2] &&
	     !sV1_sfd__h1473[1] &&
	     !sV1_sfd__h1473[0] ||
	     !_0_CONCAT_IF_IF_IF_requestR_3_BIT_214_4_THEN_re_ETC___d5008 ;
  assign IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d5326 =
	     requestR_BITS_191_TO_128__q1[63] ?
	       !IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d5315 ||
	       IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d5317 &&
	       !IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d5318 :
	       IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d5322 ||
	       IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d5317 &&
	       IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d5323 ;
  assign IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d5333 =
	     (requestR_BITS_127_TO_64__q3[62:52] == 11'd2047 &&
	      requestR_BITS_127_TO_64__q3[51] ||
	      IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d5302) ?
	       requestR[191:128] :
	       (IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d5306 ?
		  requestR[127:64] :
		  res__h217300) ;
  assign IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d5348 =
	     IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d5302 ?
	       requestR[127:64] :
	       (IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d5306 ?
		  requestR[191:128] :
		  res__h221886) ;
  assign IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d5426 =
	     (requestR_BITS_191_TO_128__q1[62:52] == 11'd0 &&
	      requestR_BITS_191_TO_128__q1[51:0] == 52'd0) ?
	       res___1__h230314 :
	       ((requestR_BITS_191_TO_128__q1[62:52] == 11'd0) ?
		  res___1__h230333 :
		  res__h230349) ;
  assign IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d571 =
	     (requestR[191:128] == 64'd0 ||
	      !sfd__h3990[63] && !sfd__h3990[62] && !sfd__h3990[61] &&
	      !sfd__h3990[60] &&
	      !sfd__h3990[59] &&
	      !sfd__h3990[58] &&
	      !sfd__h3990[57] &&
	      !sfd__h3990[56] &&
	      !sfd__h3990[55] &&
	      !sfd__h3990[54] &&
	      !sfd__h3990[53] &&
	      !sfd__h3990[52] &&
	      !sfd__h3990[51] &&
	      !sfd__h3990[50] &&
	      !sfd__h3990[49] &&
	      !sfd__h3990[48] &&
	      !sfd__h3990[47] &&
	      !sfd__h3990[46] &&
	      !sfd__h3990[45] &&
	      !sfd__h3990[44] &&
	      !sfd__h3990[43] &&
	      !sfd__h3990[42] &&
	      !sfd__h3990[41] &&
	      !sfd__h3990[40] &&
	      !sfd__h3990[39] &&
	      !sfd__h3990[38] &&
	      !sfd__h3990[37] &&
	      !sfd__h3990[36] &&
	      !sfd__h3990[35] &&
	      !sfd__h3990[34] &&
	      !sfd__h3990[33] &&
	      !sfd__h3990[32] &&
	      !sfd__h3990[31] &&
	      !sfd__h3990[30] &&
	      !sfd__h3990[29] &&
	      !sfd__h3990[28] &&
	      !sfd__h3990[27] &&
	      !sfd__h3990[26] &&
	      !sfd__h3990[25] &&
	      !sfd__h3990[24] &&
	      !sfd__h3990[23] &&
	      !sfd__h3990[22] &&
	      !sfd__h3990[21] &&
	      !sfd__h3990[20] &&
	      !sfd__h3990[19] &&
	      !sfd__h3990[18] &&
	      !sfd__h3990[17] &&
	      !sfd__h3990[16] &&
	      !sfd__h3990[15] &&
	      !sfd__h3990[14] &&
	      !sfd__h3990[13] &&
	      !sfd__h3990[12] &&
	      !sfd__h3990[11] &&
	      !sfd__h3990[10] &&
	      !sfd__h3990[9] &&
	      !sfd__h3990[8] &&
	      !sfd__h3990[7] &&
	      !sfd__h3990[6] &&
	      !sfd__h3990[5] &&
	      !sfd__h3990[4] &&
	      !sfd__h3990[3] &&
	      !sfd__h3990[2] &&
	      !sfd__h3990[1] &&
	      !sfd__h3990[0]) ?
	       8'd0 :
	       _theResult___snd_fst_exp__h16093 ;
  assign IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d684 =
	     (sfd__h3990[63] || sfd__h3990[62] || sfd__h3990[61] ||
	      sfd__h3990[60] ||
	      sfd__h3990[59] ||
	      sfd__h3990[58] ||
	      sfd__h3990[57] ||
	      sfd__h3990[56] ||
	      sfd__h3990[55] ||
	      sfd__h3990[54] ||
	      sfd__h3990[53] ||
	      sfd__h3990[52] ||
	      sfd__h3990[51] ||
	      sfd__h3990[50] ||
	      sfd__h3990[49] ||
	      sfd__h3990[48] ||
	      sfd__h3990[47] ||
	      sfd__h3990[46] ||
	      sfd__h3990[45] ||
	      sfd__h3990[44] ||
	      sfd__h3990[43] ||
	      sfd__h3990[42] ||
	      sfd__h3990[41] ||
	      sfd__h3990[40] ||
	      sfd__h3990[39] ||
	      sfd__h3990[38] ||
	      sfd__h3990[37] ||
	      sfd__h3990[36] ||
	      sfd__h3990[35] ||
	      sfd__h3990[34] ||
	      sfd__h3990[33] ||
	      sfd__h3990[32] ||
	      sfd__h3990[31] ||
	      sfd__h3990[30] ||
	      sfd__h3990[29] ||
	      sfd__h3990[28] ||
	      sfd__h3990[27] ||
	      sfd__h3990[26] ||
	      sfd__h3990[25] ||
	      sfd__h3990[24] ||
	      sfd__h3990[23] ||
	      sfd__h3990[22] ||
	      sfd__h3990[21] ||
	      sfd__h3990[20] ||
	      sfd__h3990[19] ||
	      sfd__h3990[18] ||
	      sfd__h3990[17] ||
	      sfd__h3990[16] ||
	      sfd__h3990[15] ||
	      sfd__h3990[14] ||
	      sfd__h3990[13] ||
	      sfd__h3990[12] ||
	      sfd__h3990[11] ||
	      sfd__h3990[10] ||
	      sfd__h3990[9] ||
	      sfd__h3990[8] ||
	      sfd__h3990[7] ||
	      sfd__h3990[6] ||
	      sfd__h3990[5] ||
	      sfd__h3990[4] ||
	      sfd__h3990[3] ||
	      sfd__h3990[2] ||
	      sfd__h3990[1] ||
	      sfd__h3990[0]) &&
	     (!_64_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d445 ||
	      !_64_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d447 &&
	      !_64_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d450 &&
	      _theResult___fst_exp__h16084 == 8'd255 &&
	      _theResult___fst_sfd__h16085 == 23'd0) ;
  assign IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d687 =
	     (sfd__h3990[63] || sfd__h3990[62] || sfd__h3990[61] ||
	      sfd__h3990[60] ||
	      sfd__h3990[59] ||
	      sfd__h3990[58] ||
	      sfd__h3990[57] ||
	      sfd__h3990[56] ||
	      sfd__h3990[55] ||
	      sfd__h3990[54] ||
	      sfd__h3990[53] ||
	      sfd__h3990[52] ||
	      sfd__h3990[51] ||
	      sfd__h3990[50] ||
	      sfd__h3990[49] ||
	      sfd__h3990[48] ||
	      sfd__h3990[47] ||
	      sfd__h3990[46] ||
	      sfd__h3990[45] ||
	      sfd__h3990[44] ||
	      sfd__h3990[43] ||
	      sfd__h3990[42] ||
	      sfd__h3990[41] ||
	      sfd__h3990[40] ||
	      sfd__h3990[39] ||
	      sfd__h3990[38] ||
	      sfd__h3990[37] ||
	      sfd__h3990[36] ||
	      sfd__h3990[35] ||
	      sfd__h3990[34] ||
	      sfd__h3990[33] ||
	      sfd__h3990[32] ||
	      sfd__h3990[31] ||
	      sfd__h3990[30] ||
	      sfd__h3990[29] ||
	      sfd__h3990[28] ||
	      sfd__h3990[27] ||
	      sfd__h3990[26] ||
	      sfd__h3990[25] ||
	      sfd__h3990[24] ||
	      sfd__h3990[23] ||
	      sfd__h3990[22] ||
	      sfd__h3990[21] ||
	      sfd__h3990[20] ||
	      sfd__h3990[19] ||
	      sfd__h3990[18] ||
	      sfd__h3990[17] ||
	      sfd__h3990[16] ||
	      sfd__h3990[15] ||
	      sfd__h3990[14] ||
	      sfd__h3990[13] ||
	      sfd__h3990[12] ||
	      sfd__h3990[11] ||
	      sfd__h3990[10] ||
	      sfd__h3990[9] ||
	      sfd__h3990[8] ||
	      sfd__h3990[7] ||
	      sfd__h3990[6] ||
	      sfd__h3990[5] ||
	      sfd__h3990[4] ||
	      sfd__h3990[3] ||
	      sfd__h3990[2] ||
	      sfd__h3990[1] ||
	      sfd__h3990[0]) &&
	     _64_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d445 &&
	     _64_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d447 ;
  assign IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d696 =
	     (sfd__h3990[63] || sfd__h3990[62] || sfd__h3990[61] ||
	      sfd__h3990[60] ||
	      sfd__h3990[59] ||
	      sfd__h3990[58] ||
	      sfd__h3990[57] ||
	      sfd__h3990[56] ||
	      sfd__h3990[55] ||
	      sfd__h3990[54] ||
	      sfd__h3990[53] ||
	      sfd__h3990[52] ||
	      sfd__h3990[51] ||
	      sfd__h3990[50] ||
	      sfd__h3990[49] ||
	      sfd__h3990[48] ||
	      sfd__h3990[47] ||
	      sfd__h3990[46] ||
	      sfd__h3990[45] ||
	      sfd__h3990[44] ||
	      sfd__h3990[43] ||
	      sfd__h3990[42] ||
	      sfd__h3990[41] ||
	      sfd__h3990[40] ||
	      sfd__h3990[39] ||
	      sfd__h3990[38] ||
	      sfd__h3990[37] ||
	      sfd__h3990[36] ||
	      sfd__h3990[35] ||
	      sfd__h3990[34] ||
	      sfd__h3990[33] ||
	      sfd__h3990[32] ||
	      sfd__h3990[31] ||
	      sfd__h3990[30] ||
	      sfd__h3990[29] ||
	      sfd__h3990[28] ||
	      sfd__h3990[27] ||
	      sfd__h3990[26] ||
	      sfd__h3990[25] ||
	      sfd__h3990[24] ||
	      sfd__h3990[23] ||
	      sfd__h3990[22] ||
	      sfd__h3990[21] ||
	      sfd__h3990[20] ||
	      sfd__h3990[19] ||
	      sfd__h3990[18] ||
	      sfd__h3990[17] ||
	      sfd__h3990[16] ||
	      sfd__h3990[15] ||
	      sfd__h3990[14] ||
	      sfd__h3990[13] ||
	      sfd__h3990[12] ||
	      sfd__h3990[11] ||
	      sfd__h3990[10] ||
	      sfd__h3990[9] ||
	      sfd__h3990[8] ||
	      sfd__h3990[7] ||
	      sfd__h3990[6] ||
	      sfd__h3990[5] ||
	      sfd__h3990[4] ||
	      sfd__h3990[3] ||
	      sfd__h3990[2] ||
	      sfd__h3990[1] ||
	      sfd__h3990[0]) &&
	     _64_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d445 &&
	     !_64_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d447 &&
	     IF_64_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_2_ETC___d693 ;
  assign IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d966 =
	     requestR_BITS_191_TO_128__q1[63] ?
	       7'd0 :
	       (requestR_BITS_191_TO_128__q1[62] ?
		  7'd1 :
		  (requestR_BITS_191_TO_128__q1[61] ?
		     7'd2 :
		     (requestR_BITS_191_TO_128__q1[60] ?
			7'd3 :
			(requestR_BITS_191_TO_128__q1[59] ?
			   7'd4 :
			   (requestR_BITS_191_TO_128__q1[58] ?
			      7'd5 :
			      (requestR_BITS_191_TO_128__q1[57] ?
				 7'd6 :
				 (requestR_BITS_191_TO_128__q1[56] ?
				    7'd7 :
				    (requestR_BITS_191_TO_128__q1[55] ?
				       7'd8 :
				       (requestR_BITS_191_TO_128__q1[54] ?
					  7'd9 :
					  (requestR_BITS_191_TO_128__q1[53] ?
					     7'd10 :
					     (requestR_BITS_191_TO_128__q1[52] ?
						7'd11 :
						(requestR_BITS_191_TO_128__q1[51] ?
						   7'd12 :
						   (requestR_BITS_191_TO_128__q1[50] ?
						      7'd13 :
						      (requestR_BITS_191_TO_128__q1[49] ?
							 7'd14 :
							 (requestR_BITS_191_TO_128__q1[48] ?
							    7'd15 :
							    (requestR_BITS_191_TO_128__q1[47] ?
							       7'd16 :
							       (requestR_BITS_191_TO_128__q1[46] ?
								  7'd17 :
								  (requestR_BITS_191_TO_128__q1[45] ?
								     7'd18 :
								     (requestR_BITS_191_TO_128__q1[44] ?
									7'd19 :
									(requestR_BITS_191_TO_128__q1[43] ?
									   7'd20 :
									   (requestR_BITS_191_TO_128__q1[42] ?
									      7'd21 :
									      (requestR_BITS_191_TO_128__q1[41] ?
										 7'd22 :
										 (requestR_BITS_191_TO_128__q1[40] ?
										    7'd23 :
										    (requestR_BITS_191_TO_128__q1[39] ?
										       7'd24 :
										       (requestR_BITS_191_TO_128__q1[38] ?
											  7'd25 :
											  (requestR_BITS_191_TO_128__q1[37] ?
											     7'd26 :
											     (requestR_BITS_191_TO_128__q1[36] ?
												7'd27 :
												(requestR_BITS_191_TO_128__q1[35] ?
												   7'd28 :
												   (requestR_BITS_191_TO_128__q1[34] ?
												      7'd29 :
												      (requestR_BITS_191_TO_128__q1[33] ?
													 7'd30 :
													 (requestR_BITS_191_TO_128__q1[32] ?
													    7'd31 :
													    (requestR_BITS_191_TO_128__q1[31] ?
													       7'd32 :
													       (requestR_BITS_191_TO_128__q1[30] ?
														  7'd33 :
														  (requestR_BITS_191_TO_128__q1[29] ?
														     7'd34 :
														     (requestR_BITS_191_TO_128__q1[28] ?
															7'd35 :
															(requestR_BITS_191_TO_128__q1[27] ?
															   7'd36 :
															   (requestR_BITS_191_TO_128__q1[26] ?
															      7'd37 :
															      (requestR_BITS_191_TO_128__q1[25] ?
																 7'd38 :
																 (requestR_BITS_191_TO_128__q1[24] ?
																    7'd39 :
																    (requestR_BITS_191_TO_128__q1[23] ?
																       7'd40 :
																       (requestR_BITS_191_TO_128__q1[22] ?
																	  7'd41 :
																	  (requestR_BITS_191_TO_128__q1[21] ?
																	     7'd42 :
																	     (requestR_BITS_191_TO_128__q1[20] ?
																		7'd43 :
																		(requestR_BITS_191_TO_128__q1[19] ?
																		   7'd44 :
																		   (requestR_BITS_191_TO_128__q1[18] ?
																		      7'd45 :
																		      (requestR_BITS_191_TO_128__q1[17] ?
																			 7'd46 :
																			 (requestR_BITS_191_TO_128__q1[16] ?
																			    7'd47 :
																			    (requestR_BITS_191_TO_128__q1[15] ?
																			       7'd48 :
																			       (requestR_BITS_191_TO_128__q1[14] ?
																				  7'd49 :
																				  (requestR_BITS_191_TO_128__q1[13] ?
																				     7'd50 :
																				     (requestR_BITS_191_TO_128__q1[12] ?
																					7'd51 :
																					(requestR_BITS_191_TO_128__q1[11] ?
																					   7'd52 :
																					   (requestR_BITS_191_TO_128__q1[10] ?
																					      7'd53 :
																					      (requestR_BITS_191_TO_128__q1[9] ?
																						 7'd54 :
																						 (requestR_BITS_191_TO_128__q1[8] ?
																						    7'd55 :
																						    (requestR_BITS_191_TO_128__q1[7] ?
																						       7'd56 :
																						       (requestR_BITS_191_TO_128__q1[6] ?
																							  7'd57 :
																							  (requestR_BITS_191_TO_128__q1[5] ?
																							     7'd58 :
																							     (requestR_BITS_191_TO_128__q1[4] ?
																								7'd59 :
																								(requestR_BITS_191_TO_128__q1[3] ?
																								   7'd60 :
																								   (requestR_BITS_191_TO_128__q1[2] ?
																								      7'd61 :
																								      (requestR_BITS_191_TO_128__q1[1] ?
																									 7'd62 :
																									 (requestR_BITS_191_TO_128__q1[0] ?
																									    7'd63 :
																									    7'd64))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))) ;
  assign IF_NEG_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_re_ETC___d1812 =
	     NEG_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d1785 ?
	       (IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1806 ?
		  ((x__h44058[88:25] == 64'h7FFFFFFFFFFFFFFF) ?
		     x__h44058[88:25] :
		     x__h44058[88:25] + 64'd1) :
		  x__h44058[88:25]) :
	       64'd0 ;
  assign IF_NEG_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_re_ETC___d1814 =
	     (NEG_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d1750 ==
	      20'd1048513) ?
	       ((_theResult_____2__h43093[64:63] == 2'b11) ?
		  _theResult_____2__h43093[63:0] :
		  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1745) :
	       (NEG_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d1783[19] ?
		  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1745 :
		  IF_NEG_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_re_ETC___d1812) ;
  assign IF_NEG_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_re_ETC___d1837 =
	     (NEG_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d1750 ==
	      20'd1048513) ?
	       _theResult_____2__h43093[64:63] == 2'b11 &&
	       guard__h43091 != 2'd0 :
	       !NEG_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d1783[19] &&
	       (!NEG_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d1785 ||
		guard__h43869 != 2'd0) ;
  assign IF_NEG_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_re_ETC___d1874 =
	     NEG_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d1849 ?
	       (IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1868 ?
		  ((x__h45414[88:25] == 64'hFFFFFFFFFFFFFFFF) ?
		     x__h45414[88:25] :
		     x__h45414[88:25] + 64'd1) :
		  x__h45414[88:25]) :
	       64'd0 ;
  assign IF_NEG_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_re_ETC___d1963 =
	     NEG_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d1936 ?
	       (IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1957 ?
		  ((x__h46697[56:25] == 32'h7FFFFFFF) ?
		     x__h46697[56:25] :
		     x__h46697[56:25] + 32'd1) :
		  x__h46697[56:25]) :
	       32'd0 ;
  assign IF_NEG_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_re_ETC___d1965 =
	     (NEG_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d1750 ==
	      20'd1048545) ?
	       ((_theResult_____2__h45956[32:31] == 2'b11) ?
		  _theResult_____2__h45956[31:0] :
		  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1904) :
	       (NEG_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d1934[19] ?
		  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1904 :
		  IF_NEG_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_re_ETC___d1963) ;
  assign IF_NEG_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_re_ETC___d1983 =
	     (NEG_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d1750 ==
	      20'd1048545) ?
	       _theResult_____2__h45956[32:31] == 2'b11 &&
	       guard__h45954 != 2'd0 :
	       !NEG_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d1934[19] &&
	       (!NEG_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d1936 ||
		guard__h46508 != 2'd0) ;
  assign IF_NEG_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_re_ETC___d2020 =
	     NEG_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d1995 ?
	       (IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2014 ?
		  ((x__h47815[56:25] == 32'hFFFFFFFF) ?
		     x__h47815[56:25] :
		     x__h47815[56:25] + 32'd1) :
		  x__h47815[56:25]) :
	       32'd0 ;
  assign IF_NEG_SEXT_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d2786 =
	     NEG_SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d2759 ?
	       (IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2780 ?
		  ((x__h83201[85:54] == 32'h7FFFFFFF) ?
		     x__h83201[85:54] :
		     x__h83201[85:54] + 32'd1) :
		  x__h83201[85:54]) :
	       32'd0 ;
  assign IF_NEG_SEXT_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d2788 =
	     (NEG_SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d2724 ==
	      24'd16777185) ?
	       ((_theResult_____2__h82460[32:31] == 2'b11) ?
		  _theResult_____2__h82460[31:0] :
		  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2719) :
	       (NEG_SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d2757[23] ?
		  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2719 :
		  IF_NEG_SEXT_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d2786) ;
  assign IF_NEG_SEXT_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d2812 =
	     (NEG_SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d2724 ==
	      24'd16777185) ?
	       _theResult_____2__h82460[32:31] == 2'b11 &&
	       guard__h82458 != 2'd0 :
	       !NEG_SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d2757[23] &&
	       (!NEG_SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d2759 ||
		guard__h83012 != 2'd0) ;
  assign IF_NEG_SEXT_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d2849 =
	     NEG_SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d2824 ?
	       (IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2843 ?
		  ((x__h84319[85:54] == 32'hFFFFFFFF) ?
		     x__h84319[85:54] :
		     x__h84319[85:54] + 32'd1) :
		  x__h84319[85:54]) :
	       32'd0 ;
  assign IF_NEG_SEXT_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d3279 =
	     NEG_SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d3252 ?
	       (IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d3273 ?
		  ((x__h111322[117:54] == 64'h7FFFFFFFFFFFFFFF) ?
		     x__h111322[117:54] :
		     x__h111322[117:54] + 64'd1) :
		  x__h111322[117:54]) :
	       64'd0 ;
  assign IF_NEG_SEXT_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d3281 =
	     (NEG_SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d2724 ==
	      24'd16777153) ?
	       ((_theResult_____2__h110357[64:63] == 2'b11) ?
		  _theResult_____2__h110357[63:0] :
		  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d3220) :
	       (NEG_SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d3250[23] ?
		  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d3220 :
		  IF_NEG_SEXT_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d3279) ;
  assign IF_NEG_SEXT_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d3298 =
	     (NEG_SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d2724 ==
	      24'd16777153) ?
	       _theResult_____2__h110357[64:63] == 2'b11 &&
	       guard__h110355 != 2'd0 :
	       !NEG_SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d3250[23] &&
	       (!NEG_SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d3252 ||
		guard__h111133 != 2'd0) ;
  assign IF_NEG_SEXT_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d3335 =
	     NEG_SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d3310 ?
	       (IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d3329 ?
		  ((x__h112661[117:54] == 64'hFFFFFFFFFFFFFFFF) ?
		     x__h112661[117:54] :
		     x__h112661[117:54] + 64'd1) :
		  x__h112661[117:54]) :
	       64'd0 ;
  assign IF_NOT_32_MINUS_0_CONCAT_IF_IF_IF_requestR_3_B_ETC___d2399 =
	     (!_32_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d2343 ||
	      _32_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d2345) ?
	       requestR_BITS_191_TO_128__q1[31] :
	       IF_32_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_2_ETC___d2398 ;
  assign IF_NOT_3970_MINUS_0_CONCAT_IF_IF_IF_requestR_3_ETC___d5169 =
	     (!_3970_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_21_ETC___d4542 ||
	      _3970_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_21_ETC___d4543 ||
	      _theResult___fst_exp__h190506 == 11'd2047) ?
	       requestR_BITS_191_TO_128__q1[63:32] == 32'hFFFFFFFF &&
	       requestR_BITS_191_TO_128__q1[31] :
	       ((requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
		 requestR[194:192] != 3'h3 &&
		 requestR[194:192] != 3'h4) ?
		  CASE_guard81312_0b0_requestR_BITS_191_TO_128_B_ETC__q165 :
		  CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q166) ;
  assign IF_NOT_IF_IF_requestR_3_BIT_214_4_THEN_request_ETC___d2106 =
	     NOT_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_ETC___d2105 ?
	       { requestR_BITS_191_TO_128__q1[63:32] == 32'hFFFFFFFF &&
		 requestR_BITS_191_TO_128__q1[31],
		 IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d37 } :
	       IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d48 ;
  assign IF_NOT_IF_IF_requestR_3_BIT_214_4_THEN_request_ETC___d2122 =
	     NOT_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_ETC___d2105 ?
	       IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d48 :
	       { requestR_BITS_191_TO_128__q1[63:32] == 32'hFFFFFFFF &&
		 requestR_BITS_191_TO_128__q1[31],
		 IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d37 } ;
  assign IF_NOT_IF_requestR_3_BIT_214_4_THEN_requestR_3_ETC___d2101 =
	     (requestR_BITS_191_TO_128__q1[63:32] != 32'hFFFFFFFF ||
	      !requestR_BITS_191_TO_128__q1[31]) ?
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2090 ||
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2091 &&
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2092 :
	       !IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2095 ||
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2091 &&
	       !IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2097 ;
  assign IF_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_reques_ETC___d5007 =
	     ((SEXT_IF_IF_requestR_3_BIT_214_4_THEN_requestR__ETC__q153[10:0] ==
	       11'd0) ?
		12'd3074 :
		{ SEXT_IF_IF_requestR_3_BIT_214_4_THEN_requestR__ETC__q156[10],
		  SEXT_IF_IF_requestR_3_BIT_214_4_THEN_requestR__ETC__q156 }) -
	     12'd3074 ;
  assign IF_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_reques_ETC___d5186 =
	     SEXT_IF_IF_requestR_3_BIT_214_4_THEN_requestR__ETC___d4686 ?
	       ((_theResult___fst_exp__h201334 == 11'd2047) ?
		  requestR_BITS_191_TO_128__q1[63:32] == 32'hFFFFFFFF &&
		  requestR_BITS_191_TO_128__q1[31] :
		  ((requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
		    requestR[194:192] != 3'h3 &&
		    requestR[194:192] != 3'h4) ?
		     CASE_guard91853_0b0_requestR_BITS_191_TO_128_B_ETC__q167 :
		     CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q168)) :
	       ((_theResult___fst_exp__h211398 == 11'd2047) ?
		  requestR_BITS_191_TO_128__q1[63:32] == 32'hFFFFFFFF &&
		  requestR_BITS_191_TO_128__q1[31] :
		  ((requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
		    requestR[194:192] != 3'h3 &&
		    requestR[194:192] != 3'h4) ?
		     CASE_guard02175_0b0_requestR_BITS_191_TO_128_B_ETC__q169 :
		     CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q170)) ;
  assign IF_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_reques_ETC___d5246 =
	     SEXT_IF_IF_requestR_3_BIT_214_4_THEN_requestR__ETC___d4686 ?
	       _0_CONCAT_IF_IF_3074_MINUS_SEXT_IF_IF_requestR__ETC___d5220[2] :
	       _theResult___fst_exp__h212179 == 11'd2047 &&
	       _theResult___fst_sfd__h212180 == 52'd0 ;
  assign IF_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_reques_ETC___d5258 =
	     SEXT_IF_IF_requestR_3_BIT_214_4_THEN_requestR__ETC___d4686 ?
	       _0_CONCAT_IF_IF_3074_MINUS_SEXT_IF_IF_requestR__ETC___d5220[1] :
	       _theResult___fst_exp__h211398 == 11'd0 &&
	       guard__h202175 != 2'b0 ;
  assign IF_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_reques_ETC___d5270 =
	     SEXT_IF_IF_requestR_3_BIT_214_4_THEN_requestR__ETC___d4686 ?
	       _0_CONCAT_IF_IF_3074_MINUS_SEXT_IF_IF_requestR__ETC___d5220[0] :
	       _theResult___fst_exp__h211398 != 11'd2047 &&
	       guard__h202175 != 2'b0 ;
  assign IF_SEXT_IF_requestR_3_BIT_214_4_THEN_requestR__ETC___d4172 =
	     ((SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_3_B_ETC__q121[7:0] ==
	       8'd0) ?
		9'd386 :
		{ SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_3_B_ETC__q124[7],
		  SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_3_B_ETC__q124 }) -
	     9'd386 ;
  assign IF_SEXT_IF_requestR_3_BIT_214_4_THEN_requestR__ETC___d4376 =
	     SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_3_B_ETC___d3853 ?
	       ((_theResult___fst_exp__h155731 == 8'd255) ?
		  requestR_BITS_191_TO_128__q1[63] :
		  ((requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
		    requestR[194:192] != 3'h3 &&
		    requestR[194:192] != 3'h4) ?
		     CASE_guard46250_0b0_requestR_BITS_191_TO_128_B_ETC__q147 :
		     CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q148)) :
	       ((_theResult___fst_exp__h165679 == 8'd255) ?
		  requestR_BITS_191_TO_128__q1[63] :
		  ((requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
		    requestR[194:192] != 3'h3 &&
		    requestR[194:192] != 3'h4) ?
		     CASE_guard56369_0b0_requestR_BITS_191_TO_128_B_ETC__q149 :
		     CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q150)) ;
  assign IF_SEXT_IF_requestR_3_BIT_214_4_THEN_requestR__ETC___d4454 =
	     SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_3_B_ETC___d3853 ?
	       _0_CONCAT_IF_IF_3970_MINUS_SEXT_IF_requestR_3_B_ETC___d4425[2] :
	       _theResult___fst_exp__h166257 == 8'd255 &&
	       _theResult___fst_sfd__h166258 == 23'd0 ;
  assign IF_SEXT_IF_requestR_3_BIT_214_4_THEN_requestR__ETC___d4467 =
	     SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_3_B_ETC___d3853 ?
	       _0_CONCAT_IF_IF_3970_MINUS_SEXT_IF_requestR_3_B_ETC___d4425[1] :
	       _theResult___fst_exp__h165679 == 8'd0 &&
	       guard__h156369 != 2'b0 ;
  assign IF_SEXT_IF_requestR_3_BIT_214_4_THEN_requestR__ETC___d4480 =
	     SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_3_B_ETC___d3853 ?
	       _0_CONCAT_IF_IF_3970_MINUS_SEXT_IF_requestR_3_B_ETC___d4425[0] :
	       _theResult___fst_exp__h165679 != 8'd255 &&
	       guard__h156369 != 2'b0 ;
  assign IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d1165 =
	     (requestR_BITS_191_TO_128__q1[63] ||
	      requestR_BITS_191_TO_128__q1[62] ||
	      requestR_BITS_191_TO_128__q1[61] ||
	      requestR_BITS_191_TO_128__q1[60] ||
	      requestR_BITS_191_TO_128__q1[59] ||
	      requestR_BITS_191_TO_128__q1[58] ||
	      requestR_BITS_191_TO_128__q1[57] ||
	      requestR_BITS_191_TO_128__q1[56] ||
	      requestR_BITS_191_TO_128__q1[55] ||
	      requestR_BITS_191_TO_128__q1[54] ||
	      requestR_BITS_191_TO_128__q1[53] ||
	      requestR_BITS_191_TO_128__q1[52] ||
	      requestR_BITS_191_TO_128__q1[51] ||
	      requestR_BITS_191_TO_128__q1[50] ||
	      requestR_BITS_191_TO_128__q1[49] ||
	      requestR_BITS_191_TO_128__q1[48] ||
	      requestR_BITS_191_TO_128__q1[47] ||
	      requestR_BITS_191_TO_128__q1[46] ||
	      requestR_BITS_191_TO_128__q1[45] ||
	      requestR_BITS_191_TO_128__q1[44] ||
	      requestR_BITS_191_TO_128__q1[43] ||
	      requestR_BITS_191_TO_128__q1[42] ||
	      requestR_BITS_191_TO_128__q1[41] ||
	      requestR_BITS_191_TO_128__q1[40] ||
	      requestR_BITS_191_TO_128__q1[39] ||
	      requestR_BITS_191_TO_128__q1[38] ||
	      requestR_BITS_191_TO_128__q1[37] ||
	      requestR_BITS_191_TO_128__q1[36] ||
	      requestR_BITS_191_TO_128__q1[35] ||
	      requestR_BITS_191_TO_128__q1[34] ||
	      requestR_BITS_191_TO_128__q1[33] ||
	      requestR_BITS_191_TO_128__q1[32] ||
	      requestR_BITS_191_TO_128__q1[31] ||
	      requestR_BITS_191_TO_128__q1[30] ||
	      requestR_BITS_191_TO_128__q1[29] ||
	      requestR_BITS_191_TO_128__q1[28] ||
	      requestR_BITS_191_TO_128__q1[27] ||
	      requestR_BITS_191_TO_128__q1[26] ||
	      requestR_BITS_191_TO_128__q1[25] ||
	      requestR_BITS_191_TO_128__q1[24] ||
	      requestR_BITS_191_TO_128__q1[23] ||
	      requestR_BITS_191_TO_128__q1[22] ||
	      requestR_BITS_191_TO_128__q1[21] ||
	      requestR_BITS_191_TO_128__q1[20] ||
	      requestR_BITS_191_TO_128__q1[19] ||
	      requestR_BITS_191_TO_128__q1[18] ||
	      requestR_BITS_191_TO_128__q1[17] ||
	      requestR_BITS_191_TO_128__q1[16] ||
	      requestR_BITS_191_TO_128__q1[15] ||
	      requestR_BITS_191_TO_128__q1[14] ||
	      requestR_BITS_191_TO_128__q1[13] ||
	      requestR_BITS_191_TO_128__q1[12] ||
	      requestR_BITS_191_TO_128__q1[11] ||
	      requestR_BITS_191_TO_128__q1[10] ||
	      requestR_BITS_191_TO_128__q1[9] ||
	      requestR_BITS_191_TO_128__q1[8] ||
	      requestR_BITS_191_TO_128__q1[7] ||
	      requestR_BITS_191_TO_128__q1[6] ||
	      requestR_BITS_191_TO_128__q1[5] ||
	      requestR_BITS_191_TO_128__q1[4] ||
	      requestR_BITS_191_TO_128__q1[3] ||
	      requestR_BITS_191_TO_128__q1[2] ||
	      requestR_BITS_191_TO_128__q1[1] ||
	      requestR_BITS_191_TO_128__q1[0]) &&
	     (!_64_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d970 ||
	      !_64_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d971 &&
	      !_64_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d972 &&
	      _theResult___fst_exp__h28360 == 8'd255 &&
	      _theResult___fst_sfd__h28361 == 23'd0) ;
  assign IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d1168 =
	     (requestR_BITS_191_TO_128__q1[63] ||
	      requestR_BITS_191_TO_128__q1[62] ||
	      requestR_BITS_191_TO_128__q1[61] ||
	      requestR_BITS_191_TO_128__q1[60] ||
	      requestR_BITS_191_TO_128__q1[59] ||
	      requestR_BITS_191_TO_128__q1[58] ||
	      requestR_BITS_191_TO_128__q1[57] ||
	      requestR_BITS_191_TO_128__q1[56] ||
	      requestR_BITS_191_TO_128__q1[55] ||
	      requestR_BITS_191_TO_128__q1[54] ||
	      requestR_BITS_191_TO_128__q1[53] ||
	      requestR_BITS_191_TO_128__q1[52] ||
	      requestR_BITS_191_TO_128__q1[51] ||
	      requestR_BITS_191_TO_128__q1[50] ||
	      requestR_BITS_191_TO_128__q1[49] ||
	      requestR_BITS_191_TO_128__q1[48] ||
	      requestR_BITS_191_TO_128__q1[47] ||
	      requestR_BITS_191_TO_128__q1[46] ||
	      requestR_BITS_191_TO_128__q1[45] ||
	      requestR_BITS_191_TO_128__q1[44] ||
	      requestR_BITS_191_TO_128__q1[43] ||
	      requestR_BITS_191_TO_128__q1[42] ||
	      requestR_BITS_191_TO_128__q1[41] ||
	      requestR_BITS_191_TO_128__q1[40] ||
	      requestR_BITS_191_TO_128__q1[39] ||
	      requestR_BITS_191_TO_128__q1[38] ||
	      requestR_BITS_191_TO_128__q1[37] ||
	      requestR_BITS_191_TO_128__q1[36] ||
	      requestR_BITS_191_TO_128__q1[35] ||
	      requestR_BITS_191_TO_128__q1[34] ||
	      requestR_BITS_191_TO_128__q1[33] ||
	      requestR_BITS_191_TO_128__q1[32] ||
	      requestR_BITS_191_TO_128__q1[31] ||
	      requestR_BITS_191_TO_128__q1[30] ||
	      requestR_BITS_191_TO_128__q1[29] ||
	      requestR_BITS_191_TO_128__q1[28] ||
	      requestR_BITS_191_TO_128__q1[27] ||
	      requestR_BITS_191_TO_128__q1[26] ||
	      requestR_BITS_191_TO_128__q1[25] ||
	      requestR_BITS_191_TO_128__q1[24] ||
	      requestR_BITS_191_TO_128__q1[23] ||
	      requestR_BITS_191_TO_128__q1[22] ||
	      requestR_BITS_191_TO_128__q1[21] ||
	      requestR_BITS_191_TO_128__q1[20] ||
	      requestR_BITS_191_TO_128__q1[19] ||
	      requestR_BITS_191_TO_128__q1[18] ||
	      requestR_BITS_191_TO_128__q1[17] ||
	      requestR_BITS_191_TO_128__q1[16] ||
	      requestR_BITS_191_TO_128__q1[15] ||
	      requestR_BITS_191_TO_128__q1[14] ||
	      requestR_BITS_191_TO_128__q1[13] ||
	      requestR_BITS_191_TO_128__q1[12] ||
	      requestR_BITS_191_TO_128__q1[11] ||
	      requestR_BITS_191_TO_128__q1[10] ||
	      requestR_BITS_191_TO_128__q1[9] ||
	      requestR_BITS_191_TO_128__q1[8] ||
	      requestR_BITS_191_TO_128__q1[7] ||
	      requestR_BITS_191_TO_128__q1[6] ||
	      requestR_BITS_191_TO_128__q1[5] ||
	      requestR_BITS_191_TO_128__q1[4] ||
	      requestR_BITS_191_TO_128__q1[3] ||
	      requestR_BITS_191_TO_128__q1[2] ||
	      requestR_BITS_191_TO_128__q1[1] ||
	      requestR_BITS_191_TO_128__q1[0]) &&
	     _64_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d970 &&
	     _64_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d971 ;
  assign IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d1177 =
	     (requestR_BITS_191_TO_128__q1[63] ||
	      requestR_BITS_191_TO_128__q1[62] ||
	      requestR_BITS_191_TO_128__q1[61] ||
	      requestR_BITS_191_TO_128__q1[60] ||
	      requestR_BITS_191_TO_128__q1[59] ||
	      requestR_BITS_191_TO_128__q1[58] ||
	      requestR_BITS_191_TO_128__q1[57] ||
	      requestR_BITS_191_TO_128__q1[56] ||
	      requestR_BITS_191_TO_128__q1[55] ||
	      requestR_BITS_191_TO_128__q1[54] ||
	      requestR_BITS_191_TO_128__q1[53] ||
	      requestR_BITS_191_TO_128__q1[52] ||
	      requestR_BITS_191_TO_128__q1[51] ||
	      requestR_BITS_191_TO_128__q1[50] ||
	      requestR_BITS_191_TO_128__q1[49] ||
	      requestR_BITS_191_TO_128__q1[48] ||
	      requestR_BITS_191_TO_128__q1[47] ||
	      requestR_BITS_191_TO_128__q1[46] ||
	      requestR_BITS_191_TO_128__q1[45] ||
	      requestR_BITS_191_TO_128__q1[44] ||
	      requestR_BITS_191_TO_128__q1[43] ||
	      requestR_BITS_191_TO_128__q1[42] ||
	      requestR_BITS_191_TO_128__q1[41] ||
	      requestR_BITS_191_TO_128__q1[40] ||
	      requestR_BITS_191_TO_128__q1[39] ||
	      requestR_BITS_191_TO_128__q1[38] ||
	      requestR_BITS_191_TO_128__q1[37] ||
	      requestR_BITS_191_TO_128__q1[36] ||
	      requestR_BITS_191_TO_128__q1[35] ||
	      requestR_BITS_191_TO_128__q1[34] ||
	      requestR_BITS_191_TO_128__q1[33] ||
	      requestR_BITS_191_TO_128__q1[32] ||
	      requestR_BITS_191_TO_128__q1[31] ||
	      requestR_BITS_191_TO_128__q1[30] ||
	      requestR_BITS_191_TO_128__q1[29] ||
	      requestR_BITS_191_TO_128__q1[28] ||
	      requestR_BITS_191_TO_128__q1[27] ||
	      requestR_BITS_191_TO_128__q1[26] ||
	      requestR_BITS_191_TO_128__q1[25] ||
	      requestR_BITS_191_TO_128__q1[24] ||
	      requestR_BITS_191_TO_128__q1[23] ||
	      requestR_BITS_191_TO_128__q1[22] ||
	      requestR_BITS_191_TO_128__q1[21] ||
	      requestR_BITS_191_TO_128__q1[20] ||
	      requestR_BITS_191_TO_128__q1[19] ||
	      requestR_BITS_191_TO_128__q1[18] ||
	      requestR_BITS_191_TO_128__q1[17] ||
	      requestR_BITS_191_TO_128__q1[16] ||
	      requestR_BITS_191_TO_128__q1[15] ||
	      requestR_BITS_191_TO_128__q1[14] ||
	      requestR_BITS_191_TO_128__q1[13] ||
	      requestR_BITS_191_TO_128__q1[12] ||
	      requestR_BITS_191_TO_128__q1[11] ||
	      requestR_BITS_191_TO_128__q1[10] ||
	      requestR_BITS_191_TO_128__q1[9] ||
	      requestR_BITS_191_TO_128__q1[8] ||
	      requestR_BITS_191_TO_128__q1[7] ||
	      requestR_BITS_191_TO_128__q1[6] ||
	      requestR_BITS_191_TO_128__q1[5] ||
	      requestR_BITS_191_TO_128__q1[4] ||
	      requestR_BITS_191_TO_128__q1[3] ||
	      requestR_BITS_191_TO_128__q1[2] ||
	      requestR_BITS_191_TO_128__q1[1] ||
	      requestR_BITS_191_TO_128__q1[0]) &&
	     _64_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d970 &&
	     !_64_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d971 &&
	     IF_64_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214__ETC___d1174 ;
  assign IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d1709 =
	     (requestR_BITS_191_TO_128__q1[31] ||
	      requestR_BITS_191_TO_128__q1[30] ||
	      requestR_BITS_191_TO_128__q1[29] ||
	      requestR_BITS_191_TO_128__q1[28] ||
	      requestR_BITS_191_TO_128__q1[27] ||
	      requestR_BITS_191_TO_128__q1[26] ||
	      requestR_BITS_191_TO_128__q1[25] ||
	      requestR_BITS_191_TO_128__q1[24] ||
	      requestR_BITS_191_TO_128__q1[23] ||
	      requestR_BITS_191_TO_128__q1[22] ||
	      requestR_BITS_191_TO_128__q1[21] ||
	      requestR_BITS_191_TO_128__q1[20] ||
	      requestR_BITS_191_TO_128__q1[19] ||
	      requestR_BITS_191_TO_128__q1[18] ||
	      requestR_BITS_191_TO_128__q1[17] ||
	      requestR_BITS_191_TO_128__q1[16] ||
	      requestR_BITS_191_TO_128__q1[15] ||
	      requestR_BITS_191_TO_128__q1[14] ||
	      requestR_BITS_191_TO_128__q1[13] ||
	      requestR_BITS_191_TO_128__q1[12] ||
	      requestR_BITS_191_TO_128__q1[11] ||
	      requestR_BITS_191_TO_128__q1[10] ||
	      requestR_BITS_191_TO_128__q1[9] ||
	      requestR_BITS_191_TO_128__q1[8] ||
	      requestR_BITS_191_TO_128__q1[7] ||
	      requestR_BITS_191_TO_128__q1[6] ||
	      requestR_BITS_191_TO_128__q1[5] ||
	      requestR_BITS_191_TO_128__q1[4] ||
	      requestR_BITS_191_TO_128__q1[3] ||
	      requestR_BITS_191_TO_128__q1[2] ||
	      requestR_BITS_191_TO_128__q1[1] ||
	      requestR_BITS_191_TO_128__q1[0]) &&
	     (!_32_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d1578 ||
	      !_32_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d1579 &&
	      !_32_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d1580 &&
	      _theResult___fst_exp__h42448 == 8'd255 &&
	      _theResult___fst_sfd__h42449 == 23'd0) ;
  assign IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d1712 =
	     (requestR_BITS_191_TO_128__q1[31] ||
	      requestR_BITS_191_TO_128__q1[30] ||
	      requestR_BITS_191_TO_128__q1[29] ||
	      requestR_BITS_191_TO_128__q1[28] ||
	      requestR_BITS_191_TO_128__q1[27] ||
	      requestR_BITS_191_TO_128__q1[26] ||
	      requestR_BITS_191_TO_128__q1[25] ||
	      requestR_BITS_191_TO_128__q1[24] ||
	      requestR_BITS_191_TO_128__q1[23] ||
	      requestR_BITS_191_TO_128__q1[22] ||
	      requestR_BITS_191_TO_128__q1[21] ||
	      requestR_BITS_191_TO_128__q1[20] ||
	      requestR_BITS_191_TO_128__q1[19] ||
	      requestR_BITS_191_TO_128__q1[18] ||
	      requestR_BITS_191_TO_128__q1[17] ||
	      requestR_BITS_191_TO_128__q1[16] ||
	      requestR_BITS_191_TO_128__q1[15] ||
	      requestR_BITS_191_TO_128__q1[14] ||
	      requestR_BITS_191_TO_128__q1[13] ||
	      requestR_BITS_191_TO_128__q1[12] ||
	      requestR_BITS_191_TO_128__q1[11] ||
	      requestR_BITS_191_TO_128__q1[10] ||
	      requestR_BITS_191_TO_128__q1[9] ||
	      requestR_BITS_191_TO_128__q1[8] ||
	      requestR_BITS_191_TO_128__q1[7] ||
	      requestR_BITS_191_TO_128__q1[6] ||
	      requestR_BITS_191_TO_128__q1[5] ||
	      requestR_BITS_191_TO_128__q1[4] ||
	      requestR_BITS_191_TO_128__q1[3] ||
	      requestR_BITS_191_TO_128__q1[2] ||
	      requestR_BITS_191_TO_128__q1[1] ||
	      requestR_BITS_191_TO_128__q1[0]) &&
	     _32_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d1578 &&
	     _32_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d1579 ;
  assign IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d1721 =
	     (requestR_BITS_191_TO_128__q1[31] ||
	      requestR_BITS_191_TO_128__q1[30] ||
	      requestR_BITS_191_TO_128__q1[29] ||
	      requestR_BITS_191_TO_128__q1[28] ||
	      requestR_BITS_191_TO_128__q1[27] ||
	      requestR_BITS_191_TO_128__q1[26] ||
	      requestR_BITS_191_TO_128__q1[25] ||
	      requestR_BITS_191_TO_128__q1[24] ||
	      requestR_BITS_191_TO_128__q1[23] ||
	      requestR_BITS_191_TO_128__q1[22] ||
	      requestR_BITS_191_TO_128__q1[21] ||
	      requestR_BITS_191_TO_128__q1[20] ||
	      requestR_BITS_191_TO_128__q1[19] ||
	      requestR_BITS_191_TO_128__q1[18] ||
	      requestR_BITS_191_TO_128__q1[17] ||
	      requestR_BITS_191_TO_128__q1[16] ||
	      requestR_BITS_191_TO_128__q1[15] ||
	      requestR_BITS_191_TO_128__q1[14] ||
	      requestR_BITS_191_TO_128__q1[13] ||
	      requestR_BITS_191_TO_128__q1[12] ||
	      requestR_BITS_191_TO_128__q1[11] ||
	      requestR_BITS_191_TO_128__q1[10] ||
	      requestR_BITS_191_TO_128__q1[9] ||
	      requestR_BITS_191_TO_128__q1[8] ||
	      requestR_BITS_191_TO_128__q1[7] ||
	      requestR_BITS_191_TO_128__q1[6] ||
	      requestR_BITS_191_TO_128__q1[5] ||
	      requestR_BITS_191_TO_128__q1[4] ||
	      requestR_BITS_191_TO_128__q1[3] ||
	      requestR_BITS_191_TO_128__q1[2] ||
	      requestR_BITS_191_TO_128__q1[1] ||
	      requestR_BITS_191_TO_128__q1[0]) &&
	     _32_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d1578 &&
	     !_32_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d1579 &&
	     IF_32_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214__ETC___d1718 ;
  assign IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d2103 =
	     requestR_BITS_191_TO_128__q1[63:32] == 32'hFFFFFFFF &&
	     requestR_BITS_191_TO_128__q1[31] &&
	     (requestR_BITS_127_TO_64__q3[63:32] != 32'hFFFFFFFF ||
	      !requestR_BITS_127_TO_64__q3[31]) ||
	     (requestR_BITS_191_TO_128__q1[63:32] == 32'hFFFFFFFF &&
	      requestR_BITS_191_TO_128__q1[31] ||
	      requestR_BITS_127_TO_64__q3[63:32] != 32'hFFFFFFFF ||
	      !requestR_BITS_127_TO_64__q3[31]) &&
	     IF_NOT_IF_requestR_3_BIT_214_4_THEN_requestR_3_ETC___d2101 ;
  assign IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d2169 =
	     (requestR_BITS_191_TO_128__q1[63:32] == 32'hFFFFFFFF &&
	      requestR_BITS_191_TO_128__q1[31] ||
	      requestR_BITS_127_TO_64__q3[63:32] != 32'hFFFFFFFF ||
	      !requestR_BITS_127_TO_64__q3[31]) &&
	     ((requestR_BITS_191_TO_128__q1[63:32] != 32'hFFFFFFFF ||
	       !requestR_BITS_191_TO_128__q1[31]) ?
		NOT_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_ETC___d2166 :
		IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2167) ;
  assign IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d2722 =
	     requestR_BITS_191_TO_128__q1[62:52] - 11'd1023 ;
  assign IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d2861 =
	     requestR_BITS_191_TO_128__q1[62:52] == 11'd2047 &&
	     requestR_BITS_191_TO_128__q1[51:0] != 52'd0 ||
	     requestR_BITS_191_TO_128__q1[62:52] == 11'd2047 &&
	     requestR_BITS_191_TO_128__q1[51:0] == 52'd0 ||
	     (requestR_BITS_191_TO_128__q1[62:52] != 11'd0 ||
	      requestR_BITS_191_TO_128__q1[51:0] != 52'd0) &&
	     (NEG_SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d2822[23] ||
	      NEG_SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d2824 &&
	      IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2843 &&
	      x__h84319[85:54] == 32'hFFFFFFFF) ;
  assign IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d2872 =
	     { IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d2861,
	       3'd0,
	       (requestR_BITS_191_TO_128__q1[62:52] != 11'd2047 ||
		requestR_BITS_191_TO_128__q1[51:0] == 52'd0) &&
	       (requestR_BITS_191_TO_128__q1[62:52] != 11'd2047 ||
		requestR_BITS_191_TO_128__q1[51:0] != 52'd0) &&
	       NOT_IF_requestR_3_BIT_214_4_THEN_requestR_3_BI_ETC___d2866 } ==
	     5'd0 ||
	     IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d2861 ;
  assign IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d3199 =
	     (requestR_BITS_191_TO_128__q1[63] ||
	      requestR_BITS_191_TO_128__q1[62] ||
	      requestR_BITS_191_TO_128__q1[61] ||
	      requestR_BITS_191_TO_128__q1[60] ||
	      requestR_BITS_191_TO_128__q1[59] ||
	      requestR_BITS_191_TO_128__q1[58] ||
	      requestR_BITS_191_TO_128__q1[57] ||
	      requestR_BITS_191_TO_128__q1[56] ||
	      requestR_BITS_191_TO_128__q1[55] ||
	      requestR_BITS_191_TO_128__q1[54] ||
	      requestR_BITS_191_TO_128__q1[53] ||
	      requestR_BITS_191_TO_128__q1[52] ||
	      requestR_BITS_191_TO_128__q1[51] ||
	      requestR_BITS_191_TO_128__q1[50] ||
	      requestR_BITS_191_TO_128__q1[49] ||
	      requestR_BITS_191_TO_128__q1[48] ||
	      requestR_BITS_191_TO_128__q1[47] ||
	      requestR_BITS_191_TO_128__q1[46] ||
	      requestR_BITS_191_TO_128__q1[45] ||
	      requestR_BITS_191_TO_128__q1[44] ||
	      requestR_BITS_191_TO_128__q1[43] ||
	      requestR_BITS_191_TO_128__q1[42] ||
	      requestR_BITS_191_TO_128__q1[41] ||
	      requestR_BITS_191_TO_128__q1[40] ||
	      requestR_BITS_191_TO_128__q1[39] ||
	      requestR_BITS_191_TO_128__q1[38] ||
	      requestR_BITS_191_TO_128__q1[37] ||
	      requestR_BITS_191_TO_128__q1[36] ||
	      requestR_BITS_191_TO_128__q1[35] ||
	      requestR_BITS_191_TO_128__q1[34] ||
	      requestR_BITS_191_TO_128__q1[33] ||
	      requestR_BITS_191_TO_128__q1[32] ||
	      requestR_BITS_191_TO_128__q1[31] ||
	      requestR_BITS_191_TO_128__q1[30] ||
	      requestR_BITS_191_TO_128__q1[29] ||
	      requestR_BITS_191_TO_128__q1[28] ||
	      requestR_BITS_191_TO_128__q1[27] ||
	      requestR_BITS_191_TO_128__q1[26] ||
	      requestR_BITS_191_TO_128__q1[25] ||
	      requestR_BITS_191_TO_128__q1[24] ||
	      requestR_BITS_191_TO_128__q1[23] ||
	      requestR_BITS_191_TO_128__q1[22] ||
	      requestR_BITS_191_TO_128__q1[21] ||
	      requestR_BITS_191_TO_128__q1[20] ||
	      requestR_BITS_191_TO_128__q1[19] ||
	      requestR_BITS_191_TO_128__q1[18] ||
	      requestR_BITS_191_TO_128__q1[17] ||
	      requestR_BITS_191_TO_128__q1[16] ||
	      requestR_BITS_191_TO_128__q1[15] ||
	      requestR_BITS_191_TO_128__q1[14] ||
	      requestR_BITS_191_TO_128__q1[13] ||
	      requestR_BITS_191_TO_128__q1[12] ||
	      requestR_BITS_191_TO_128__q1[11] ||
	      requestR_BITS_191_TO_128__q1[10] ||
	      requestR_BITS_191_TO_128__q1[9] ||
	      requestR_BITS_191_TO_128__q1[8] ||
	      requestR_BITS_191_TO_128__q1[7] ||
	      requestR_BITS_191_TO_128__q1[6] ||
	      requestR_BITS_191_TO_128__q1[5] ||
	      requestR_BITS_191_TO_128__q1[4] ||
	      requestR_BITS_191_TO_128__q1[3] ||
	      requestR_BITS_191_TO_128__q1[2] ||
	      requestR_BITS_191_TO_128__q1[1] ||
	      requestR_BITS_191_TO_128__q1[0]) &&
	     (!_64_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d3069 ||
	      !_64_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d3070 &&
	      !_64_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d3071 &&
	      _theResult___fst_exp__h109716 == 11'd2047 &&
	      _theResult___fst_sfd__h109717 == 52'd0) ;
  assign IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d3202 =
	     (requestR_BITS_191_TO_128__q1[63] ||
	      requestR_BITS_191_TO_128__q1[62] ||
	      requestR_BITS_191_TO_128__q1[61] ||
	      requestR_BITS_191_TO_128__q1[60] ||
	      requestR_BITS_191_TO_128__q1[59] ||
	      requestR_BITS_191_TO_128__q1[58] ||
	      requestR_BITS_191_TO_128__q1[57] ||
	      requestR_BITS_191_TO_128__q1[56] ||
	      requestR_BITS_191_TO_128__q1[55] ||
	      requestR_BITS_191_TO_128__q1[54] ||
	      requestR_BITS_191_TO_128__q1[53] ||
	      requestR_BITS_191_TO_128__q1[52] ||
	      requestR_BITS_191_TO_128__q1[51] ||
	      requestR_BITS_191_TO_128__q1[50] ||
	      requestR_BITS_191_TO_128__q1[49] ||
	      requestR_BITS_191_TO_128__q1[48] ||
	      requestR_BITS_191_TO_128__q1[47] ||
	      requestR_BITS_191_TO_128__q1[46] ||
	      requestR_BITS_191_TO_128__q1[45] ||
	      requestR_BITS_191_TO_128__q1[44] ||
	      requestR_BITS_191_TO_128__q1[43] ||
	      requestR_BITS_191_TO_128__q1[42] ||
	      requestR_BITS_191_TO_128__q1[41] ||
	      requestR_BITS_191_TO_128__q1[40] ||
	      requestR_BITS_191_TO_128__q1[39] ||
	      requestR_BITS_191_TO_128__q1[38] ||
	      requestR_BITS_191_TO_128__q1[37] ||
	      requestR_BITS_191_TO_128__q1[36] ||
	      requestR_BITS_191_TO_128__q1[35] ||
	      requestR_BITS_191_TO_128__q1[34] ||
	      requestR_BITS_191_TO_128__q1[33] ||
	      requestR_BITS_191_TO_128__q1[32] ||
	      requestR_BITS_191_TO_128__q1[31] ||
	      requestR_BITS_191_TO_128__q1[30] ||
	      requestR_BITS_191_TO_128__q1[29] ||
	      requestR_BITS_191_TO_128__q1[28] ||
	      requestR_BITS_191_TO_128__q1[27] ||
	      requestR_BITS_191_TO_128__q1[26] ||
	      requestR_BITS_191_TO_128__q1[25] ||
	      requestR_BITS_191_TO_128__q1[24] ||
	      requestR_BITS_191_TO_128__q1[23] ||
	      requestR_BITS_191_TO_128__q1[22] ||
	      requestR_BITS_191_TO_128__q1[21] ||
	      requestR_BITS_191_TO_128__q1[20] ||
	      requestR_BITS_191_TO_128__q1[19] ||
	      requestR_BITS_191_TO_128__q1[18] ||
	      requestR_BITS_191_TO_128__q1[17] ||
	      requestR_BITS_191_TO_128__q1[16] ||
	      requestR_BITS_191_TO_128__q1[15] ||
	      requestR_BITS_191_TO_128__q1[14] ||
	      requestR_BITS_191_TO_128__q1[13] ||
	      requestR_BITS_191_TO_128__q1[12] ||
	      requestR_BITS_191_TO_128__q1[11] ||
	      requestR_BITS_191_TO_128__q1[10] ||
	      requestR_BITS_191_TO_128__q1[9] ||
	      requestR_BITS_191_TO_128__q1[8] ||
	      requestR_BITS_191_TO_128__q1[7] ||
	      requestR_BITS_191_TO_128__q1[6] ||
	      requestR_BITS_191_TO_128__q1[5] ||
	      requestR_BITS_191_TO_128__q1[4] ||
	      requestR_BITS_191_TO_128__q1[3] ||
	      requestR_BITS_191_TO_128__q1[2] ||
	      requestR_BITS_191_TO_128__q1[1] ||
	      requestR_BITS_191_TO_128__q1[0]) &&
	     _64_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d3069 &&
	     _64_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d3070 ;
  assign IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d3211 =
	     (requestR_BITS_191_TO_128__q1[63] ||
	      requestR_BITS_191_TO_128__q1[62] ||
	      requestR_BITS_191_TO_128__q1[61] ||
	      requestR_BITS_191_TO_128__q1[60] ||
	      requestR_BITS_191_TO_128__q1[59] ||
	      requestR_BITS_191_TO_128__q1[58] ||
	      requestR_BITS_191_TO_128__q1[57] ||
	      requestR_BITS_191_TO_128__q1[56] ||
	      requestR_BITS_191_TO_128__q1[55] ||
	      requestR_BITS_191_TO_128__q1[54] ||
	      requestR_BITS_191_TO_128__q1[53] ||
	      requestR_BITS_191_TO_128__q1[52] ||
	      requestR_BITS_191_TO_128__q1[51] ||
	      requestR_BITS_191_TO_128__q1[50] ||
	      requestR_BITS_191_TO_128__q1[49] ||
	      requestR_BITS_191_TO_128__q1[48] ||
	      requestR_BITS_191_TO_128__q1[47] ||
	      requestR_BITS_191_TO_128__q1[46] ||
	      requestR_BITS_191_TO_128__q1[45] ||
	      requestR_BITS_191_TO_128__q1[44] ||
	      requestR_BITS_191_TO_128__q1[43] ||
	      requestR_BITS_191_TO_128__q1[42] ||
	      requestR_BITS_191_TO_128__q1[41] ||
	      requestR_BITS_191_TO_128__q1[40] ||
	      requestR_BITS_191_TO_128__q1[39] ||
	      requestR_BITS_191_TO_128__q1[38] ||
	      requestR_BITS_191_TO_128__q1[37] ||
	      requestR_BITS_191_TO_128__q1[36] ||
	      requestR_BITS_191_TO_128__q1[35] ||
	      requestR_BITS_191_TO_128__q1[34] ||
	      requestR_BITS_191_TO_128__q1[33] ||
	      requestR_BITS_191_TO_128__q1[32] ||
	      requestR_BITS_191_TO_128__q1[31] ||
	      requestR_BITS_191_TO_128__q1[30] ||
	      requestR_BITS_191_TO_128__q1[29] ||
	      requestR_BITS_191_TO_128__q1[28] ||
	      requestR_BITS_191_TO_128__q1[27] ||
	      requestR_BITS_191_TO_128__q1[26] ||
	      requestR_BITS_191_TO_128__q1[25] ||
	      requestR_BITS_191_TO_128__q1[24] ||
	      requestR_BITS_191_TO_128__q1[23] ||
	      requestR_BITS_191_TO_128__q1[22] ||
	      requestR_BITS_191_TO_128__q1[21] ||
	      requestR_BITS_191_TO_128__q1[20] ||
	      requestR_BITS_191_TO_128__q1[19] ||
	      requestR_BITS_191_TO_128__q1[18] ||
	      requestR_BITS_191_TO_128__q1[17] ||
	      requestR_BITS_191_TO_128__q1[16] ||
	      requestR_BITS_191_TO_128__q1[15] ||
	      requestR_BITS_191_TO_128__q1[14] ||
	      requestR_BITS_191_TO_128__q1[13] ||
	      requestR_BITS_191_TO_128__q1[12] ||
	      requestR_BITS_191_TO_128__q1[11] ||
	      requestR_BITS_191_TO_128__q1[10] ||
	      requestR_BITS_191_TO_128__q1[9] ||
	      requestR_BITS_191_TO_128__q1[8] ||
	      requestR_BITS_191_TO_128__q1[7] ||
	      requestR_BITS_191_TO_128__q1[6] ||
	      requestR_BITS_191_TO_128__q1[5] ||
	      requestR_BITS_191_TO_128__q1[4] ||
	      requestR_BITS_191_TO_128__q1[3] ||
	      requestR_BITS_191_TO_128__q1[2] ||
	      requestR_BITS_191_TO_128__q1[1] ||
	      requestR_BITS_191_TO_128__q1[0]) &&
	     _64_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d3069 &&
	     !_64_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d3070 &&
	     IF_64_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214__ETC___d3208 ;
  assign IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d3346 =
	     requestR_BITS_191_TO_128__q1[62:52] == 11'd2047 &&
	     requestR_BITS_191_TO_128__q1[51:0] != 52'd0 ||
	     requestR_BITS_191_TO_128__q1[62:52] == 11'd2047 &&
	     requestR_BITS_191_TO_128__q1[51:0] == 52'd0 ||
	     (requestR_BITS_191_TO_128__q1[62:52] != 11'd0 ||
	      requestR_BITS_191_TO_128__q1[51:0] != 52'd0) &&
	     (NEG_SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d3308[23] ||
	      NEG_SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d3310 &&
	      IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d3329 &&
	      x__h112661[117:54] == 64'hFFFFFFFFFFFFFFFF) ;
  assign IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d3357 =
	     { IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d3346,
	       3'd0,
	       (requestR_BITS_191_TO_128__q1[62:52] != 11'd2047 ||
		requestR_BITS_191_TO_128__q1[51:0] == 52'd0) &&
	       (requestR_BITS_191_TO_128__q1[62:52] != 11'd2047 ||
		requestR_BITS_191_TO_128__q1[51:0] != 52'd0) &&
	       NOT_IF_requestR_3_BIT_214_4_THEN_requestR_3_BI_ETC___d3351 } ==
	     5'd0 ||
	     IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d3346 ;
  assign IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d48 =
	     { requestR_BITS_127_TO_64__q3[63:32] == 32'hFFFFFFFF &&
	       requestR_BITS_127_TO_64__q3[31],
	       (requestR_BITS_127_TO_64__q3[63:32] == 32'hFFFFFFFF) ?
		 requestR_BITS_127_TO_64__q3[30:0] :
		 31'h7FC00000 } ;
  assign IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d5294 =
	     requestR_BITS_191_TO_128__q1[62:52] == 11'd2047 &&
	     requestR_BITS_191_TO_128__q1[51:0] != 52'd0 &&
	     !requestR_BITS_191_TO_128__q1[51] &&
	     requestR_BITS_127_TO_64__q3[62:52] == 11'd2047 &&
	     requestR_BITS_127_TO_64__q3[51:0] != 52'd0 &&
	     !requestR_BITS_127_TO_64__q3[51] ;
  assign IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d5302 =
	     requestR_BITS_191_TO_128__q1[62:52] == 11'd0 &&
	     requestR_BITS_191_TO_128__q1[51:0] == 52'd0 &&
	     requestR_BITS_191_TO_128__q1[63] &&
	     requestR_BITS_127_TO_64__q3[62:52] == 11'd0 &&
	     requestR_BITS_127_TO_64__q3[51:0] == 52'd0 &&
	     !requestR_BITS_127_TO_64__q3[63] ;
  assign IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d5306 =
	     requestR_BITS_127_TO_64__q3[62:52] == 11'd0 &&
	     requestR_BITS_127_TO_64__q3[51:0] == 52'd0 &&
	     requestR_BITS_127_TO_64__q3[63] &&
	     requestR_BITS_191_TO_128__q1[62:52] == 11'd0 &&
	     requestR_BITS_191_TO_128__q1[51:0] == 52'd0 &&
	     !requestR_BITS_191_TO_128__q1[63] ;
  assign IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d5315 =
	     requestR_BITS_191_TO_128__q1[62:52] <=
	     requestR_BITS_127_TO_64__q3[62:52] ;
  assign IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d5317 =
	     requestR_BITS_191_TO_128__q1[62:52] ==
	     requestR_BITS_127_TO_64__q3[62:52] ;
  assign IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d5318 =
	     requestR_BITS_191_TO_128__q1[51:0] <=
	     requestR_BITS_127_TO_64__q3[51:0] ;
  assign IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d5322 =
	     requestR_BITS_191_TO_128__q1[62:52] <
	     requestR_BITS_127_TO_64__q3[62:52] ;
  assign IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d5323 =
	     requestR_BITS_191_TO_128__q1[51:0] <
	     requestR_BITS_127_TO_64__q3[51:0] ;
  assign IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d5339 =
	     requestR_BITS_191_TO_128__q1[62:52] == 11'd2047 &&
	     requestR_BITS_191_TO_128__q1[51:0] != 52'd0 &&
	     !requestR_BITS_191_TO_128__q1[51] ||
	     requestR_BITS_127_TO_64__q3[62:52] == 11'd2047 &&
	     requestR_BITS_127_TO_64__q3[51:0] != 52'd0 &&
	     !requestR_BITS_127_TO_64__q3[51] ;
  assign IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d5363 =
	     IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d5339 ||
	     requestR_BITS_191_TO_128__q1[62:52] == 11'd2047 &&
	     requestR_BITS_191_TO_128__q1[51] ||
	     requestR_BITS_127_TO_64__q3[62:52] == 11'd2047 &&
	     requestR_BITS_127_TO_64__q3[51] ;
  assign IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d5373 =
	     IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d5315 &&
	     (!IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d5317 ||
	      IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d5318) &&
	     !IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d5322 &&
	     (!IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d5317 ||
	      !IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d5323) ;
  assign IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d5378 =
	     requestR_BITS_191_TO_128__q1[62:52] == 11'd0 &&
	     requestR_BITS_191_TO_128__q1[51:0] == 52'd0 &&
	     requestR_BITS_127_TO_64__q3[62:52] == 11'd0 &&
	     requestR_BITS_127_TO_64__q3[51:0] == 52'd0 ||
	     (!requestR_BITS_191_TO_128__q1[63] ||
	      requestR_BITS_127_TO_64__q3[63]) &&
	     (requestR_BITS_191_TO_128__q1[63] ||
	      !requestR_BITS_127_TO_64__q3[63]) &&
	     (requestR_BITS_191_TO_128__q1[63] ?
		IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d5373 :
		NOT_IF_requestR_3_BIT_214_4_THEN_requestR_3_BI_ETC___d5374) ;
  assign IF_sfd___30336_BIT_1_THEN_2_ELSE_0__q85 =
	     sfd___3__h80336[1] ? 2'd2 : 2'd0 ;
  assign IF_sfd___30336_BIT_2_THEN_2_ELSE_0__q84 =
	     sfd___3__h80336[2] ? 2'd2 : 2'd0 ;
  assign IF_sfd___31374_BIT_7_THEN_2_ELSE_0__q56 =
	     sfd___3__h41374[7] ? 2'd2 : 2'd0 ;
  assign IF_sfd___31374_BIT_8_THEN_2_ELSE_0__q55 =
	     sfd___3__h41374[8] ? 2'd2 : 2'd0 ;
  assign IF_sfd___34458_BIT_7_THEN_2_ELSE_0__q42 =
	     sfd___3__h34458[7] ? 2'd2 : 2'd0 ;
  assign IF_sfd___34458_BIT_8_THEN_2_ELSE_0__q41 =
	     sfd___3__h34458[8] ? 2'd2 : 2'd0 ;
  assign IF_sfd___35005_BIT_10_THEN_2_ELSE_0__q12 =
	     sfd___3__h15005[10] ? 2'd2 : 2'd0 ;
  assign IF_sfd___35005_BIT_11_THEN_2_ELSE_0__q11 =
	     sfd___3__h15005[11] ? 2'd2 : 2'd0 ;
  assign IF_sfd___35005_BIT_39_THEN_2_ELSE_0__q10 =
	     sfd___3__h15005[39] ? 2'd2 : 2'd0 ;
  assign IF_sfd___35005_BIT_40_THEN_2_ELSE_0__q9 =
	     sfd___3__h15005[40] ? 2'd2 : 2'd0 ;
  assign IF_sfd___37286_BIT_10_THEN_2_ELSE_0__q28 =
	     sfd___3__h27286[10] ? 2'd2 : 2'd0 ;
  assign IF_sfd___37286_BIT_11_THEN_2_ELSE_0__q27 =
	     sfd___3__h27286[11] ? 2'd2 : 2'd0 ;
  assign IF_sfd___37286_BIT_39_THEN_2_ELSE_0__q26 =
	     sfd___3__h27286[39] ? 2'd2 : 2'd0 ;
  assign IF_sfd___37286_BIT_40_THEN_2_ELSE_0__q25 =
	     sfd___3__h27286[40] ? 2'd2 : 2'd0 ;
  assign IF_sfd___39389_BIT_1_THEN_2_ELSE_0__q71 =
	     sfd___3__h69389[1] ? 2'd2 : 2'd0 ;
  assign IF_sfd___39389_BIT_2_THEN_2_ELSE_0__q70 =
	     sfd___3__h69389[2] ? 2'd2 : 2'd0 ;
  assign IF_sfdin01328_BIT_4_THEN_2_ELSE_0__q155 =
	     sfdin__h201328[4] ? 2'd2 : 2'd0 ;
  assign IF_sfdin35384_BIT_33_THEN_2_ELSE_0__q118 =
	     sfdin__h135384[33] ? 2'd2 : 2'd0 ;
  assign IF_sfdin55725_BIT_33_THEN_2_ELSE_0__q123 =
	     sfdin__h155725[33] ? 2'd2 : 2'd0 ;
  assign IF_theResult___snd11344_BIT_4_THEN_2_ELSE_0__q158 =
	     _theResult___snd__h211344[4] ? 2'd2 : 2'd0 ;
  assign IF_theResult___snd45260_BIT_33_THEN_2_ELSE_0__q120 =
	     _theResult___snd__h145260[33] ? 2'd2 : 2'd0 ;
  assign IF_theResult___snd65625_BIT_33_THEN_2_ELSE_0__q126 =
	     _theResult___snd__h165625[33] ? 2'd2 : 2'd0 ;
  assign IF_theResult___snd90457_BIT_4_THEN_2_ELSE_0__q152 =
	     _theResult___snd__h190457[4] ? 2'd2 : 2'd0 ;
  assign IF_x11322_BIT_53_THEN_2_ELSE_0__q115 = x__h111322[53] ? 2'd2 : 2'd0 ;
  assign IF_x12661_BIT_53_THEN_2_ELSE_0__q116 = x__h112661[53] ? 2'd2 : 2'd0 ;
  assign IF_x3201_BIT_53_THEN_2_ELSE_0__q95 = x__h83201[53] ? 2'd2 : 2'd0 ;
  assign IF_x4058_BIT_24_THEN_2_ELSE_0__q66 = x__h44058[24] ? 2'd2 : 2'd0 ;
  assign IF_x4319_BIT_53_THEN_2_ELSE_0__q96 = x__h84319[53] ? 2'd2 : 2'd0 ;
  assign IF_x5414_BIT_24_THEN_2_ELSE_0__q67 = x__h45414[24] ? 2'd2 : 2'd0 ;
  assign IF_x6697_BIT_24_THEN_2_ELSE_0__q68 = x__h46697[24] ? 2'd2 : 2'd0 ;
  assign IF_x7815_BIT_24_THEN_2_ELSE_0__q69 = x__h47815[24] ? 2'd2 : 2'd0 ;
  assign NEG_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d1750 =
	     -{ {12{IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1748[7]}},
		IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1748 } ;
  assign NEG_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d1782 =
	     NEG_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d1750 +
	     20'd64 ;
  assign NEG_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d1783 =
	     NEG_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d1782 -
	     20'd2 ;
  assign NEG_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d1785 =
	     (NEG_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d1783 ^
	      20'h80000) <=
	     20'd524352 ;
  assign NEG_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d1847 =
	     NEG_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d1782 -
	     20'd1 ;
  assign NEG_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d1849 =
	     (NEG_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d1847 ^
	      20'h80000) <=
	     20'd524352 ;
  assign NEG_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d1933 =
	     NEG_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d1750 +
	     20'd32 ;
  assign NEG_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d1934 =
	     NEG_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d1933 -
	     20'd2 ;
  assign NEG_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d1936 =
	     (NEG_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d1934 ^
	      20'h80000) <=
	     20'd524320 ;
  assign NEG_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d1993 =
	     NEG_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d1933 -
	     20'd1 ;
  assign NEG_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d1995 =
	     (NEG_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d1993 ^
	      20'h80000) <=
	     20'd524320 ;
  assign NEG_SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d2724 =
	     -{ {13{IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d2722[10]}},
		IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d2722 } ;
  assign NEG_SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d2756 =
	     NEG_SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d2724 +
	     24'd32 ;
  assign NEG_SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d2757 =
	     NEG_SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d2756 -
	     24'd2 ;
  assign NEG_SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d2759 =
	     (NEG_SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d2757 ^
	      24'h800000) <=
	     24'd8388640 ;
  assign NEG_SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d2822 =
	     NEG_SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d2756 -
	     24'd1 ;
  assign NEG_SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d2824 =
	     (NEG_SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d2822 ^
	      24'h800000) <=
	     24'd8388640 ;
  assign NEG_SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d3249 =
	     NEG_SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d2724 +
	     24'd64 ;
  assign NEG_SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d3250 =
	     NEG_SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d3249 -
	     24'd2 ;
  assign NEG_SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d3252 =
	     (NEG_SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d3250 ^
	      24'h800000) <=
	     24'd8388672 ;
  assign NEG_SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d3308 =
	     NEG_SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d3249 -
	     24'd1 ;
  assign NEG_SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d3310 =
	     (NEG_SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d3308 ^
	      24'h800000) <=
	     24'd8388672 ;
  assign NOT_3074_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_2_ETC___d4448 =
	     !_3074_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_ETC___d3421 ||
	     (_3074_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_ETC___d3422 ?
		_0_CONCAT_IF_IF_0b0_CONCAT_NOT_IF_requestR_3_BI_ETC___d4396[2] :
		_0_CONCAT_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d4408[2]) ;
  assign NOT_3074_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_2_ETC___d4476 =
	     !_3074_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_ETC___d3421 ||
	     (_3074_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_ETC___d3422 ?
		_0_CONCAT_IF_IF_0b0_CONCAT_NOT_IF_requestR_3_BI_ETC___d4396[0] :
		_0_CONCAT_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d4408[0]) ;
  assign NOT_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_ETC___d1326 =
	     !sfd__h28849[31] && !sfd__h28849[30] && !sfd__h28849[29] &&
	     !sfd__h28849[28] &&
	     !sfd__h28849[27] &&
	     !sfd__h28849[26] &&
	     !sfd__h28849[25] &&
	     !sfd__h28849[24] &&
	     !sfd__h28849[23] &&
	     !sfd__h28849[22] &&
	     !sfd__h28849[21] &&
	     !sfd__h28849[20] &&
	     !sfd__h28849[19] &&
	     !sfd__h28849[18] &&
	     !sfd__h28849[17] &&
	     !sfd__h28849[16] &&
	     !sfd__h28849[15] &&
	     !sfd__h28849[14] &&
	     !sfd__h28849[13] &&
	     !sfd__h28849[12] &&
	     !sfd__h28849[11] &&
	     !sfd__h28849[10] &&
	     !sfd__h28849[9] &&
	     !sfd__h28849[8] &&
	     !sfd__h28849[7] &&
	     !sfd__h28849[6] &&
	     !sfd__h28849[5] &&
	     !sfd__h28849[4] &&
	     !sfd__h28849[3] &&
	     !sfd__h28849[2] &&
	     !sfd__h28849[1] &&
	     !sfd__h28849[0] ||
	     !_32_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d1322 ||
	     _32_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d1324 ;
  assign NOT_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_ETC___d1826 =
	     (sV1_exp__h1472 != 8'd0 || sV1_sfd__h1473 != 23'd0) &&
	     ((NEG_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d1750 ==
	       20'd1048513) ?
		_theResult_____2__h43093[64:63] != 2'b11 :
		NEG_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d1783[19] ||
		NEG_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d1785 &&
		IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1806 &&
		x__h44058[88:25] == 64'h7FFFFFFFFFFFFFFF) ;
  assign NOT_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_ETC___d1890 =
	     (sV1_exp__h1472 != 8'd0 || sV1_sfd__h1473 != 23'd0) &&
	     !NEG_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d1847[19] &&
	     (!NEG_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d1849 ||
	      guard__h45193 != 2'd0) ;
  assign NOT_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_ETC___d1975 =
	     (sV1_exp__h1472 != 8'd0 || sV1_sfd__h1473 != 23'd0) &&
	     ((NEG_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d1750 ==
	       20'd1048545) ?
		_theResult_____2__h45956[32:31] != 2'b11 :
		NEG_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d1934[19] ||
		NEG_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d1936 &&
		IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1957 &&
		x__h46697[56:25] == 32'h7FFFFFFF) ;
  assign NOT_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_ETC___d2037 =
	     (sV1_exp__h1472 != 8'd0 || sV1_sfd__h1473 != 23'd0) &&
	     !NEG_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d1993[19] &&
	     (!NEG_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d1995 ||
	      guard__h47594 != 2'd0) ;
  assign NOT_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_ETC___d2104 =
	     (sV1_exp__h1472 != 8'd0 || sV1_sfd__h1473 != 23'd0 ||
	      sV2_exp__h1597 != 8'd0 ||
	      sV2_sfd__h1598 != 23'd0) &&
	     IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d2103 ;
  assign NOT_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_ETC___d2105 =
	     (sV1_exp__h1472 != 8'd255 || sV1_sfd__h1473 == 23'd0) &&
	     (sV2_exp__h1597 != 8'd255 || sV2_sfd__h1598 == 23'd0) &&
	     NOT_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_ETC___d2104 ;
  assign NOT_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_ETC___d2166 =
	     !IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2090 &&
	     (!IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2091 ||
	      !IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2092) &&
	     IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2095 &&
	     (!IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2091 ||
	      IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2097) ;
  assign NOT_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_ETC___d2172 =
	     (sV1_exp__h1472 != 8'd255 || sV1_sfd__h1473 == 23'd0) &&
	     (sV2_exp__h1597 != 8'd255 || sV2_sfd__h1598 == 23'd0) &&
	     IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2171 ;
  assign NOT_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_ETC___d2192 =
	     (sV1_exp__h1472 != 8'd255 || sV1_sfd__h1473 == 23'd0) &&
	     (sV2_exp__h1597 != 8'd255 || sV2_sfd__h1598 == 23'd0) &&
	     (IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d2103 ||
	      IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2171) ;
  assign NOT_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_ETC___d2887 =
	     !sfd__h3990[63] && !sfd__h3990[62] && !sfd__h3990[61] &&
	     !sfd__h3990[60] &&
	     !sfd__h3990[59] &&
	     !sfd__h3990[58] &&
	     !sfd__h3990[57] &&
	     !sfd__h3990[56] &&
	     !sfd__h3990[55] &&
	     !sfd__h3990[54] &&
	     !sfd__h3990[53] &&
	     !sfd__h3990[52] &&
	     !sfd__h3990[51] &&
	     !sfd__h3990[50] &&
	     !sfd__h3990[49] &&
	     !sfd__h3990[48] &&
	     !sfd__h3990[47] &&
	     !sfd__h3990[46] &&
	     !sfd__h3990[45] &&
	     !sfd__h3990[44] &&
	     !sfd__h3990[43] &&
	     !sfd__h3990[42] &&
	     !sfd__h3990[41] &&
	     !sfd__h3990[40] &&
	     !sfd__h3990[39] &&
	     !sfd__h3990[38] &&
	     !sfd__h3990[37] &&
	     !sfd__h3990[36] &&
	     !sfd__h3990[35] &&
	     !sfd__h3990[34] &&
	     !sfd__h3990[33] &&
	     !sfd__h3990[32] &&
	     !sfd__h3990[31] &&
	     !sfd__h3990[30] &&
	     !sfd__h3990[29] &&
	     !sfd__h3990[28] &&
	     !sfd__h3990[27] &&
	     !sfd__h3990[26] &&
	     !sfd__h3990[25] &&
	     !sfd__h3990[24] &&
	     !sfd__h3990[23] &&
	     !sfd__h3990[22] &&
	     !sfd__h3990[21] &&
	     !sfd__h3990[20] &&
	     !sfd__h3990[19] &&
	     !sfd__h3990[18] &&
	     !sfd__h3990[17] &&
	     !sfd__h3990[16] &&
	     !sfd__h3990[15] &&
	     !sfd__h3990[14] &&
	     !sfd__h3990[13] &&
	     !sfd__h3990[12] &&
	     !sfd__h3990[11] &&
	     !sfd__h3990[10] &&
	     !sfd__h3990[9] &&
	     !sfd__h3990[8] &&
	     !sfd__h3990[7] &&
	     !sfd__h3990[6] &&
	     !sfd__h3990[5] &&
	     !sfd__h3990[4] &&
	     !sfd__h3990[3] &&
	     !sfd__h3990[2] &&
	     !sfd__h3990[1] &&
	     !sfd__h3990[0] ||
	     !_64_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d2883 ||
	     _64_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d2885 ;
  assign NOT_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_ETC___d449 =
	     !sfd__h3990[63] && !sfd__h3990[62] && !sfd__h3990[61] &&
	     !sfd__h3990[60] &&
	     !sfd__h3990[59] &&
	     !sfd__h3990[58] &&
	     !sfd__h3990[57] &&
	     !sfd__h3990[56] &&
	     !sfd__h3990[55] &&
	     !sfd__h3990[54] &&
	     !sfd__h3990[53] &&
	     !sfd__h3990[52] &&
	     !sfd__h3990[51] &&
	     !sfd__h3990[50] &&
	     !sfd__h3990[49] &&
	     !sfd__h3990[48] &&
	     !sfd__h3990[47] &&
	     !sfd__h3990[46] &&
	     !sfd__h3990[45] &&
	     !sfd__h3990[44] &&
	     !sfd__h3990[43] &&
	     !sfd__h3990[42] &&
	     !sfd__h3990[41] &&
	     !sfd__h3990[40] &&
	     !sfd__h3990[39] &&
	     !sfd__h3990[38] &&
	     !sfd__h3990[37] &&
	     !sfd__h3990[36] &&
	     !sfd__h3990[35] &&
	     !sfd__h3990[34] &&
	     !sfd__h3990[33] &&
	     !sfd__h3990[32] &&
	     !sfd__h3990[31] &&
	     !sfd__h3990[30] &&
	     !sfd__h3990[29] &&
	     !sfd__h3990[28] &&
	     !sfd__h3990[27] &&
	     !sfd__h3990[26] &&
	     !sfd__h3990[25] &&
	     !sfd__h3990[24] &&
	     !sfd__h3990[23] &&
	     !sfd__h3990[22] &&
	     !sfd__h3990[21] &&
	     !sfd__h3990[20] &&
	     !sfd__h3990[19] &&
	     !sfd__h3990[18] &&
	     !sfd__h3990[17] &&
	     !sfd__h3990[16] &&
	     !sfd__h3990[15] &&
	     !sfd__h3990[14] &&
	     !sfd__h3990[13] &&
	     !sfd__h3990[12] &&
	     !sfd__h3990[11] &&
	     !sfd__h3990[10] &&
	     !sfd__h3990[9] &&
	     !sfd__h3990[8] &&
	     !sfd__h3990[7] &&
	     !sfd__h3990[6] &&
	     !sfd__h3990[5] &&
	     !sfd__h3990[4] &&
	     !sfd__h3990[3] &&
	     !sfd__h3990[2] &&
	     !sfd__h3990[1] &&
	     !sfd__h3990[0] ||
	     !_64_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d445 ||
	     _64_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d447 ;
  assign NOT_IF_requestR_3_BIT_214_4_THEN_requestR_3_BI_ETC___d1059 =
	     !requestR_BITS_191_TO_128__q1[63] &&
	     !requestR_BITS_191_TO_128__q1[62] &&
	     !requestR_BITS_191_TO_128__q1[61] &&
	     !requestR_BITS_191_TO_128__q1[60] &&
	     !requestR_BITS_191_TO_128__q1[59] &&
	     !requestR_BITS_191_TO_128__q1[58] &&
	     !requestR_BITS_191_TO_128__q1[57] &&
	     !requestR_BITS_191_TO_128__q1[56] &&
	     !requestR_BITS_191_TO_128__q1[55] &&
	     !requestR_BITS_191_TO_128__q1[54] &&
	     !requestR_BITS_191_TO_128__q1[53] &&
	     !requestR_BITS_191_TO_128__q1[52] &&
	     !requestR_BITS_191_TO_128__q1[51] &&
	     !requestR_BITS_191_TO_128__q1[50] &&
	     !requestR_BITS_191_TO_128__q1[49] &&
	     !requestR_BITS_191_TO_128__q1[48] &&
	     !requestR_BITS_191_TO_128__q1[47] &&
	     !requestR_BITS_191_TO_128__q1[46] &&
	     !requestR_BITS_191_TO_128__q1[45] &&
	     !requestR_BITS_191_TO_128__q1[44] &&
	     !requestR_BITS_191_TO_128__q1[43] &&
	     !requestR_BITS_191_TO_128__q1[42] &&
	     !requestR_BITS_191_TO_128__q1[41] &&
	     !requestR_BITS_191_TO_128__q1[40] &&
	     !requestR_BITS_191_TO_128__q1[39] &&
	     !requestR_BITS_191_TO_128__q1[38] &&
	     !requestR_BITS_191_TO_128__q1[37] &&
	     !requestR_BITS_191_TO_128__q1[36] &&
	     !requestR_BITS_191_TO_128__q1[35] &&
	     !requestR_BITS_191_TO_128__q1[34] &&
	     !requestR_BITS_191_TO_128__q1[33] &&
	     !requestR_BITS_191_TO_128__q1[32] &&
	     !requestR_BITS_191_TO_128__q1[31] &&
	     !requestR_BITS_191_TO_128__q1[30] &&
	     !requestR_BITS_191_TO_128__q1[29] &&
	     !requestR_BITS_191_TO_128__q1[28] &&
	     !requestR_BITS_191_TO_128__q1[27] &&
	     !requestR_BITS_191_TO_128__q1[26] &&
	     !requestR_BITS_191_TO_128__q1[25] &&
	     !requestR_BITS_191_TO_128__q1[24] &&
	     !requestR_BITS_191_TO_128__q1[23] &&
	     !requestR_BITS_191_TO_128__q1[22] &&
	     !requestR_BITS_191_TO_128__q1[21] &&
	     !requestR_BITS_191_TO_128__q1[20] &&
	     !requestR_BITS_191_TO_128__q1[19] &&
	     !requestR_BITS_191_TO_128__q1[18] &&
	     !requestR_BITS_191_TO_128__q1[17] &&
	     !requestR_BITS_191_TO_128__q1[16] &&
	     !requestR_BITS_191_TO_128__q1[15] &&
	     !requestR_BITS_191_TO_128__q1[14] &&
	     !requestR_BITS_191_TO_128__q1[13] &&
	     !requestR_BITS_191_TO_128__q1[12] &&
	     !requestR_BITS_191_TO_128__q1[11] &&
	     !requestR_BITS_191_TO_128__q1[10] &&
	     !requestR_BITS_191_TO_128__q1[9] &&
	     !requestR_BITS_191_TO_128__q1[8] &&
	     !requestR_BITS_191_TO_128__q1[7] &&
	     !requestR_BITS_191_TO_128__q1[6] &&
	     !requestR_BITS_191_TO_128__q1[5] &&
	     !requestR_BITS_191_TO_128__q1[4] &&
	     !requestR_BITS_191_TO_128__q1[3] &&
	     !requestR_BITS_191_TO_128__q1[2] &&
	     !requestR_BITS_191_TO_128__q1[1] &&
	     !requestR_BITS_191_TO_128__q1[0] ||
	     !_64_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d970 ||
	     _64_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d971 ;
  assign NOT_IF_requestR_3_BIT_214_4_THEN_requestR_3_BI_ETC___d1666 =
	     !requestR_BITS_191_TO_128__q1[31] &&
	     !requestR_BITS_191_TO_128__q1[30] &&
	     !requestR_BITS_191_TO_128__q1[29] &&
	     !requestR_BITS_191_TO_128__q1[28] &&
	     !requestR_BITS_191_TO_128__q1[27] &&
	     !requestR_BITS_191_TO_128__q1[26] &&
	     !requestR_BITS_191_TO_128__q1[25] &&
	     !requestR_BITS_191_TO_128__q1[24] &&
	     !requestR_BITS_191_TO_128__q1[23] &&
	     !requestR_BITS_191_TO_128__q1[22] &&
	     !requestR_BITS_191_TO_128__q1[21] &&
	     !requestR_BITS_191_TO_128__q1[20] &&
	     !requestR_BITS_191_TO_128__q1[19] &&
	     !requestR_BITS_191_TO_128__q1[18] &&
	     !requestR_BITS_191_TO_128__q1[17] &&
	     !requestR_BITS_191_TO_128__q1[16] &&
	     !requestR_BITS_191_TO_128__q1[15] &&
	     !requestR_BITS_191_TO_128__q1[14] &&
	     !requestR_BITS_191_TO_128__q1[13] &&
	     !requestR_BITS_191_TO_128__q1[12] &&
	     !requestR_BITS_191_TO_128__q1[11] &&
	     !requestR_BITS_191_TO_128__q1[10] &&
	     !requestR_BITS_191_TO_128__q1[9] &&
	     !requestR_BITS_191_TO_128__q1[8] &&
	     !requestR_BITS_191_TO_128__q1[7] &&
	     !requestR_BITS_191_TO_128__q1[6] &&
	     !requestR_BITS_191_TO_128__q1[5] &&
	     !requestR_BITS_191_TO_128__q1[4] &&
	     !requestR_BITS_191_TO_128__q1[3] &&
	     !requestR_BITS_191_TO_128__q1[2] &&
	     !requestR_BITS_191_TO_128__q1[1] &&
	     !requestR_BITS_191_TO_128__q1[0] ||
	     !_32_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d1578 ||
	     _32_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d1579 ;
  assign NOT_IF_requestR_3_BIT_214_4_THEN_requestR_3_BI_ETC___d2801 =
	     (requestR_BITS_191_TO_128__q1[62:52] != 11'd0 ||
	      requestR_BITS_191_TO_128__q1[51:0] != 52'd0) &&
	     ((NEG_SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d2724 ==
	       24'd16777185) ?
		_theResult_____2__h82460[32:31] != 2'b11 :
		NEG_SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d2757[23] ||
		NEG_SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d2759 &&
		IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2780 &&
		x__h83201[85:54] == 32'h7FFFFFFF) ;
  assign NOT_IF_requestR_3_BIT_214_4_THEN_requestR_3_BI_ETC___d2866 =
	     (requestR_BITS_191_TO_128__q1[62:52] != 11'd0 ||
	      requestR_BITS_191_TO_128__q1[51:0] != 52'd0) &&
	     !NEG_SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d2822[23] &&
	     (!NEG_SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d2824 ||
	      guard__h84098 != 2'd0) ;
  assign NOT_IF_requestR_3_BIT_214_4_THEN_requestR_3_BI_ETC___d3156 =
	     !requestR_BITS_191_TO_128__q1[63] &&
	     !requestR_BITS_191_TO_128__q1[62] &&
	     !requestR_BITS_191_TO_128__q1[61] &&
	     !requestR_BITS_191_TO_128__q1[60] &&
	     !requestR_BITS_191_TO_128__q1[59] &&
	     !requestR_BITS_191_TO_128__q1[58] &&
	     !requestR_BITS_191_TO_128__q1[57] &&
	     !requestR_BITS_191_TO_128__q1[56] &&
	     !requestR_BITS_191_TO_128__q1[55] &&
	     !requestR_BITS_191_TO_128__q1[54] &&
	     !requestR_BITS_191_TO_128__q1[53] &&
	     !requestR_BITS_191_TO_128__q1[52] &&
	     !requestR_BITS_191_TO_128__q1[51] &&
	     !requestR_BITS_191_TO_128__q1[50] &&
	     !requestR_BITS_191_TO_128__q1[49] &&
	     !requestR_BITS_191_TO_128__q1[48] &&
	     !requestR_BITS_191_TO_128__q1[47] &&
	     !requestR_BITS_191_TO_128__q1[46] &&
	     !requestR_BITS_191_TO_128__q1[45] &&
	     !requestR_BITS_191_TO_128__q1[44] &&
	     !requestR_BITS_191_TO_128__q1[43] &&
	     !requestR_BITS_191_TO_128__q1[42] &&
	     !requestR_BITS_191_TO_128__q1[41] &&
	     !requestR_BITS_191_TO_128__q1[40] &&
	     !requestR_BITS_191_TO_128__q1[39] &&
	     !requestR_BITS_191_TO_128__q1[38] &&
	     !requestR_BITS_191_TO_128__q1[37] &&
	     !requestR_BITS_191_TO_128__q1[36] &&
	     !requestR_BITS_191_TO_128__q1[35] &&
	     !requestR_BITS_191_TO_128__q1[34] &&
	     !requestR_BITS_191_TO_128__q1[33] &&
	     !requestR_BITS_191_TO_128__q1[32] &&
	     !requestR_BITS_191_TO_128__q1[31] &&
	     !requestR_BITS_191_TO_128__q1[30] &&
	     !requestR_BITS_191_TO_128__q1[29] &&
	     !requestR_BITS_191_TO_128__q1[28] &&
	     !requestR_BITS_191_TO_128__q1[27] &&
	     !requestR_BITS_191_TO_128__q1[26] &&
	     !requestR_BITS_191_TO_128__q1[25] &&
	     !requestR_BITS_191_TO_128__q1[24] &&
	     !requestR_BITS_191_TO_128__q1[23] &&
	     !requestR_BITS_191_TO_128__q1[22] &&
	     !requestR_BITS_191_TO_128__q1[21] &&
	     !requestR_BITS_191_TO_128__q1[20] &&
	     !requestR_BITS_191_TO_128__q1[19] &&
	     !requestR_BITS_191_TO_128__q1[18] &&
	     !requestR_BITS_191_TO_128__q1[17] &&
	     !requestR_BITS_191_TO_128__q1[16] &&
	     !requestR_BITS_191_TO_128__q1[15] &&
	     !requestR_BITS_191_TO_128__q1[14] &&
	     !requestR_BITS_191_TO_128__q1[13] &&
	     !requestR_BITS_191_TO_128__q1[12] &&
	     !requestR_BITS_191_TO_128__q1[11] &&
	     !requestR_BITS_191_TO_128__q1[10] &&
	     !requestR_BITS_191_TO_128__q1[9] &&
	     !requestR_BITS_191_TO_128__q1[8] &&
	     !requestR_BITS_191_TO_128__q1[7] &&
	     !requestR_BITS_191_TO_128__q1[6] &&
	     !requestR_BITS_191_TO_128__q1[5] &&
	     !requestR_BITS_191_TO_128__q1[4] &&
	     !requestR_BITS_191_TO_128__q1[3] &&
	     !requestR_BITS_191_TO_128__q1[2] &&
	     !requestR_BITS_191_TO_128__q1[1] &&
	     !requestR_BITS_191_TO_128__q1[0] ||
	     !_64_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d3069 ||
	     _64_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d3070 ;
  assign NOT_IF_requestR_3_BIT_214_4_THEN_requestR_3_BI_ETC___d3290 =
	     (requestR_BITS_191_TO_128__q1[62:52] != 11'd0 ||
	      requestR_BITS_191_TO_128__q1[51:0] != 52'd0) &&
	     ((NEG_SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d2724 ==
	       24'd16777153) ?
		_theResult_____2__h110357[64:63] != 2'b11 :
		NEG_SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d3250[23] ||
		NEG_SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d3252 &&
		IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d3273 &&
		x__h111322[117:54] == 64'h7FFFFFFFFFFFFFFF) ;
  assign NOT_IF_requestR_3_BIT_214_4_THEN_requestR_3_BI_ETC___d3351 =
	     (requestR_BITS_191_TO_128__q1[62:52] != 11'd0 ||
	      requestR_BITS_191_TO_128__q1[51:0] != 52'd0) &&
	     !NEG_SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d3308[23] &&
	     (!NEG_SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d3310 ||
	      guard__h112440 != 2'd0) ;
  assign NOT_IF_requestR_3_BIT_214_4_THEN_requestR_3_BI_ETC___d5330 =
	     (requestR_BITS_191_TO_128__q1[62:52] != 11'd2047 ||
	      requestR_BITS_191_TO_128__q1[51:0] == 52'd0) &&
	     (requestR_BITS_127_TO_64__q3[62:52] != 11'd2047 ||
	      requestR_BITS_127_TO_64__q3[51:0] == 52'd0) &&
	     (requestR_BITS_191_TO_128__q1[62:52] != 11'd0 ||
	      requestR_BITS_191_TO_128__q1[51:0] != 52'd0 ||
	      requestR_BITS_127_TO_64__q3[62:52] != 11'd0 ||
	      requestR_BITS_127_TO_64__q3[51:0] != 52'd0) &&
	     (requestR_BITS_191_TO_128__q1[63] &&
	      !requestR_BITS_127_TO_64__q3[63] ||
	      (requestR_BITS_191_TO_128__q1[63] ||
	       !requestR_BITS_127_TO_64__q3[63]) &&
	      IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d5326) ;
  assign NOT_IF_requestR_3_BIT_214_4_THEN_requestR_3_BI_ETC___d5374 =
	     !IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d5322 &&
	     (!IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d5317 ||
	      !IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d5323) &&
	     IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d5315 &&
	     (!IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d5317 ||
	      IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d5318) ;
  assign NOT_IF_requestR_3_BIT_214_4_THEN_requestR_3_BI_ETC___d5399 =
	     (requestR_BITS_191_TO_128__q1[62:52] != 11'd2047 ||
	      requestR_BITS_191_TO_128__q1[51:0] == 52'd0) &&
	     (requestR_BITS_127_TO_64__q3[62:52] != 11'd2047 ||
	      requestR_BITS_127_TO_64__q3[51:0] == 52'd0) &&
	     (requestR_BITS_191_TO_128__q1[63] &&
	      !requestR_BITS_127_TO_64__q3[63] ||
	      (requestR_BITS_191_TO_128__q1[63] ||
	       !requestR_BITS_127_TO_64__q3[63]) &&
	      IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d5326 ||
	      IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d5378) ;
  assign NOT_verbosity_ULE_1_6___d27 = verbosity > 4'd1 ;
  assign NOT_verbosity_ULE_2_01___d702 = verbosity > 4'd2 ;
  assign SEXT_IF_IF_requestR_3_BIT_214_4_THEN_requestR__ETC___d4684 =
	     { {4{IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1748[7]}},
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1748 } ;
  assign SEXT_IF_IF_requestR_3_BIT_214_4_THEN_requestR__ETC___d4685 =
	     (SEXT_IF_IF_requestR_3_BIT_214_4_THEN_requestR__ETC___d4684 ^
	      12'h800) <=
	     12'd3071 ;
  assign SEXT_IF_IF_requestR_3_BIT_214_4_THEN_requestR__ETC___d4686 =
	     (SEXT_IF_IF_requestR_3_BIT_214_4_THEN_requestR__ETC___d4684 ^
	      12'h800) <
	     12'd1026 ;
  assign SEXT_IF_IF_requestR_3_BIT_214_4_THEN_requestR__ETC__q153 =
	     SEXT_IF_IF_requestR_3_BIT_214_4_THEN_requestR__ETC___d4684 +
	     12'd1023 ;
  assign SEXT_IF_IF_requestR_3_BIT_214_4_THEN_requestR__ETC__q156 =
	     SEXT_IF_IF_requestR_3_BIT_214_4_THEN_requestR__ETC__q153[10:0] -
	     11'd1023 ;
  assign SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_3_B_ETC___d3851 =
	     { IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d2722[10],
	       IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d2722 } ;
  assign SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_3_B_ETC___d3852 =
	     (SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_3_B_ETC___d3851 ^
	      12'h800) <=
	     12'd2175 ;
  assign SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_3_B_ETC___d3853 =
	     (SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_3_B_ETC___d3851 ^
	      12'h800) <
	     12'd1922 ;
  assign SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_3_B_ETC__q121 =
	     SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_3_B_ETC___d3851 +
	     12'd127 ;
  assign SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_3_B_ETC__q124 =
	     SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_3_B_ETC__q121[7:0] -
	     8'd127 ;
  assign _0_CONCAT_IF_IF_0b0_CONCAT_NOT_IF_requestR_3_BI_ETC___d3656 =
	     ({ 3'd0,
		IF_IF_0b0_CONCAT_NOT_IF_requestR_3_BIT_214_4_T_ETC___d3654 } ^
	      9'h100) <=
	     9'd256 ;
  assign _0_CONCAT_IF_IF_0b0_CONCAT_NOT_IF_requestR_3_BI_ETC___d4396 =
	     { 3'd0,
	       _theResult___fst_exp__h135390 == 8'd0 &&
	       (sfdin__h135384[56:34] == 23'd0 || guard__h126038 != 2'b0),
	       1'd0 } |
	     { 2'd0,
	       _theResult___fst_exp__h136017 == 8'd255 &&
	       _theResult___fst_sfd__h136018 == 23'd0,
	       1'd0,
	       _theResult___fst_exp__h135390 != 8'd255 &&
	       guard__h126038 != 2'b0 } ;
  assign _0_CONCAT_IF_IF_3074_MINUS_SEXT_IF_IF_requestR__ETC___d4935 =
	     ({ 6'd0,
		IF_IF_3074_MINUS_SEXT_IF_IF_requestR_3_BIT_214_ETC___d4933 } ^
	      12'h800) <=
	     12'd2048 ;
  assign _0_CONCAT_IF_IF_3074_MINUS_SEXT_IF_IF_requestR__ETC___d5220 =
	     { 3'd0,
	       _theResult___fst_exp__h201334 == 11'd0 &&
	       (sfdin__h201328[56:5] == 52'd0 || guard__h191853 != 2'b0),
	       1'd0 } |
	     { 2'd0,
	       _theResult___fst_exp__h202164 == 11'd2047 &&
	       _theResult___fst_sfd__h202165 == 52'd0,
	       1'd0,
	       _theResult___fst_exp__h201334 != 11'd2047 &&
	       guard__h191853 != 2'b0 } ;
  assign _0_CONCAT_IF_IF_3970_MINUS_SEXT_IF_requestR_3_B_ETC___d4100 =
	     ({ 3'd0,
		IF_IF_3970_MINUS_SEXT_IF_requestR_3_BIT_214_4__ETC___d4098 } ^
	      9'h100) <=
	     9'd256 ;
  assign _0_CONCAT_IF_IF_3970_MINUS_SEXT_IF_requestR_3_B_ETC___d4425 =
	     { 3'd0,
	       _theResult___fst_exp__h155731 == 8'd0 &&
	       (sfdin__h155725[56:34] == 23'd0 || guard__h146250 != 2'b0),
	       1'd0 } |
	     { 2'd0,
	       _theResult___fst_exp__h156358 == 8'd255 &&
	       _theResult___fst_sfd__h156359 == 23'd0,
	       1'd0,
	       _theResult___fst_exp__h155731 != 8'd255 &&
	       guard__h146250 != 2'b0 } ;
  assign _0_CONCAT_IF_IF_IF_requestR_3_BIT_214_4_THEN_re_ETC___d4615 =
	     ({ 6'd0,
		IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3__ETC___d4613 } ^
	      12'h800) <=
	     12'd2944 ;
  assign _0_CONCAT_IF_IF_IF_requestR_3_BIT_214_4_THEN_re_ETC___d5008 =
	     ({ 6'd0,
		IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3__ETC___d4613 } ^
	      12'h800) <=
	     (IF_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_reques_ETC___d5007 ^
	      12'h800) ;
  assign _0_CONCAT_IF_IF_IF_requestR_3_BIT_214_4_THEN_re_ETC___d5203 =
	     { 3'd0,
	       _theResult___fst_exp__h190506 == 11'd0 &&
	       guard__h181312 != 2'b0,
	       1'd0 } |
	     { 2'd0,
	       _theResult___fst_exp__h191262 == 11'd2047 &&
	       _theResult___fst_sfd__h191263 == 52'd0,
	       1'd0,
	       _theResult___fst_exp__h190506 != 11'd2047 &&
	       guard__h181312 != 2'b0 } ;
  assign _0_CONCAT_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d3778 =
	     ({ 3'd0,
		IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d3776 } ^
	      9'h100) <=
	     9'd384 ;
  assign _0_CONCAT_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d4173 =
	     ({ 3'd0,
		IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d3776 } ^
	      9'h100) <=
	     (IF_SEXT_IF_requestR_3_BIT_214_4_THEN_requestR__ETC___d4172 ^
	      9'h100) ;
  assign _0_CONCAT_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d4408 =
	     { 3'd0,
	       _theResult___fst_exp__h145309 == 8'd0 &&
	       guard__h136028 != 2'b0,
	       1'd0 } |
	     { 2'd0,
	       _theResult___fst_exp__h145862 == 8'd255 &&
	       _theResult___fst_sfd__h145863 == 23'd0,
	       1'd0,
	       _theResult___fst_exp__h145309 != 8'd255 &&
	       guard__h136028 != 2'b0 } ;
  assign _0b0_CONCAT_NOT_IF_IF_requestR_3_BIT_214_4_THEN_ETC___d4691 =
	     b__h46021 >>
	     _3074_MINUS_SEXT_IF_IF_requestR_3_BIT_214_4_THE_ETC___d4687 ;
  assign _0b0_CONCAT_NOT_IF_requestR_3_BIT_214_4_THEN_re_ETC___d3858 =
	     sfd__h117253 >>
	     _3970_MINUS_SEXT_IF_requestR_3_BIT_214_4_THEN_r_ETC___d3854 ;
  assign _1_CONCAT_DONTCARE_CONCAT_IF_requestR_3_BIT_214_ETC___d97 =
	     { 33'h1AAAAAAAA,
	       requestR_BITS_63_TO_0__q8[63:32] == 32'hFFFFFFFF &&
	       requestR_BITS_63_TO_0__q8[31],
	       (requestR_BITS_63_TO_0__q8[63:32] == 32'hFFFFFFFF) ?
		 requestR_BITS_63_TO_0__q8[30:0] :
		 31'h7FC00000 } ;
  assign _3074_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_ETC___d3420 =
	     12'd3074 -
	     { 6'd0,
	       requestR_BITS_191_TO_128__q1[51] ?
		 6'd0 :
		 (requestR_BITS_191_TO_128__q1[50] ?
		    6'd1 :
		    (requestR_BITS_191_TO_128__q1[49] ?
		       6'd2 :
		       (requestR_BITS_191_TO_128__q1[48] ?
			  6'd3 :
			  (requestR_BITS_191_TO_128__q1[47] ?
			     6'd4 :
			     (requestR_BITS_191_TO_128__q1[46] ?
				6'd5 :
				(requestR_BITS_191_TO_128__q1[45] ?
				   6'd6 :
				   (requestR_BITS_191_TO_128__q1[44] ?
				      6'd7 :
				      (requestR_BITS_191_TO_128__q1[43] ?
					 6'd8 :
					 (requestR_BITS_191_TO_128__q1[42] ?
					    6'd9 :
					    (requestR_BITS_191_TO_128__q1[41] ?
					       6'd10 :
					       (requestR_BITS_191_TO_128__q1[40] ?
						  6'd11 :
						  (requestR_BITS_191_TO_128__q1[39] ?
						     6'd12 :
						     (requestR_BITS_191_TO_128__q1[38] ?
							6'd13 :
							(requestR_BITS_191_TO_128__q1[37] ?
							   6'd14 :
							   (requestR_BITS_191_TO_128__q1[36] ?
							      6'd15 :
							      (requestR_BITS_191_TO_128__q1[35] ?
								 6'd16 :
								 (requestR_BITS_191_TO_128__q1[34] ?
								    6'd17 :
								    (requestR_BITS_191_TO_128__q1[33] ?
								       6'd18 :
								       (requestR_BITS_191_TO_128__q1[32] ?
									  6'd19 :
									  (requestR_BITS_191_TO_128__q1[31] ?
									     6'd20 :
									     (requestR_BITS_191_TO_128__q1[30] ?
										6'd21 :
										(requestR_BITS_191_TO_128__q1[29] ?
										   6'd22 :
										   (requestR_BITS_191_TO_128__q1[28] ?
										      6'd23 :
										      (requestR_BITS_191_TO_128__q1[27] ?
											 6'd24 :
											 (requestR_BITS_191_TO_128__q1[26] ?
											    6'd25 :
											    (requestR_BITS_191_TO_128__q1[25] ?
											       6'd26 :
											       (requestR_BITS_191_TO_128__q1[24] ?
												  6'd27 :
												  (requestR_BITS_191_TO_128__q1[23] ?
												     6'd28 :
												     (requestR_BITS_191_TO_128__q1[22] ?
													6'd29 :
													(requestR_BITS_191_TO_128__q1[21] ?
													   6'd30 :
													   (requestR_BITS_191_TO_128__q1[20] ?
													      6'd31 :
													      (requestR_BITS_191_TO_128__q1[19] ?
														 6'd32 :
														 (requestR_BITS_191_TO_128__q1[18] ?
														    6'd33 :
														    (requestR_BITS_191_TO_128__q1[17] ?
														       6'd34 :
														       (requestR_BITS_191_TO_128__q1[16] ?
															  6'd35 :
															  (requestR_BITS_191_TO_128__q1[15] ?
															     6'd36 :
															     (requestR_BITS_191_TO_128__q1[14] ?
																6'd37 :
																(requestR_BITS_191_TO_128__q1[13] ?
																   6'd38 :
																   (requestR_BITS_191_TO_128__q1[12] ?
																      6'd39 :
																      (requestR_BITS_191_TO_128__q1[11] ?
																	 6'd40 :
																	 (requestR_BITS_191_TO_128__q1[10] ?
																	    6'd41 :
																	    (requestR_BITS_191_TO_128__q1[9] ?
																	       6'd42 :
																	       (requestR_BITS_191_TO_128__q1[8] ?
																		  6'd43 :
																		  (requestR_BITS_191_TO_128__q1[7] ?
																		     6'd44 :
																		     (requestR_BITS_191_TO_128__q1[6] ?
																			6'd45 :
																			(requestR_BITS_191_TO_128__q1[5] ?
																			   6'd46 :
																			   (requestR_BITS_191_TO_128__q1[4] ?
																			      6'd47 :
																			      (requestR_BITS_191_TO_128__q1[3] ?
																				 6'd48 :
																				 (requestR_BITS_191_TO_128__q1[2] ?
																				    6'd49 :
																				    (requestR_BITS_191_TO_128__q1[1] ?
																				       6'd50 :
																				       (requestR_BITS_191_TO_128__q1[0] ?
																					  6'd51 :
																					  6'd52))))))))))))))))))))))))))))))))))))))))))))))))))) } ;
  assign _3074_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_ETC___d3421 =
	     (_3074_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_ETC___d3420 ^
	      12'h800) <=
	     12'd2175 ;
  assign _3074_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_ETC___d3422 =
	     (_3074_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_ETC___d3420 ^
	      12'h800) <
	     12'd1922 ;
  assign _3074_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_ETC___d4411 =
	     _3074_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_ETC___d3421 &&
	     (_3074_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_ETC___d3422 ?
		_0_CONCAT_IF_IF_0b0_CONCAT_NOT_IF_requestR_3_BI_ETC___d4396[4] :
		_0_CONCAT_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d4408[4]) ;
  assign _3074_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_ETC___d4436 =
	     _3074_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_ETC___d3421 &&
	     (_3074_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_ETC___d3422 ?
		_0_CONCAT_IF_IF_0b0_CONCAT_NOT_IF_requestR_3_BI_ETC___d4396[3] :
		_0_CONCAT_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d4408[3]) ;
  assign _3074_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_ETC___d4463 =
	     _3074_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_ETC___d3421 &&
	     (_3074_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_ETC___d3422 ?
		_0_CONCAT_IF_IF_0b0_CONCAT_NOT_IF_requestR_3_BI_ETC___d4396[1] :
		_0_CONCAT_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d4408[1]) ;
  assign _3074_MINUS_SEXT_IF_IF_requestR_3_BIT_214_4_THE_ETC___d4687 =
	     12'd3074 -
	     SEXT_IF_IF_requestR_3_BIT_214_4_THEN_requestR__ETC___d4684 ;
  assign _32_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d1321 =
	     (9'd32 -
	      { 3'd0,
		IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3__ETC___d1318 }) -
	     9'd1 ;
  assign _32_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d1322 =
	     (_32_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d1321 ^
	      9'h100) <=
	     9'd383 ;
  assign _32_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d1324 =
	     (_32_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d1321 ^
	      9'h100) <
	     9'd107 ;
  assign _32_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d1327 =
	     (_32_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d1321 ^
	      9'h100) <
	     9'd130 ;
  assign _32_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d2342 =
	     (12'd32 -
	      { 6'd0,
		IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3__ETC___d2339 }) -
	     12'd1 ;
  assign _32_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d2343 =
	     (_32_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d2342 ^
	      12'h800) <=
	     12'd3071 ;
  assign _32_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d2345 =
	     (_32_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d2342 ^
	      12'h800) <
	     12'd974 ;
  assign _32_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d2347 =
	     (_32_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d2342 ^
	      12'h800) <
	     12'd1026 ;
  assign _32_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d1577 =
	     (9'd32 -
	      { 3'd0,
		IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1574 }) -
	     9'd1 ;
  assign _32_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d1578 =
	     (_32_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d1577 ^
	      9'h100) <=
	     9'd383 ;
  assign _32_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d1579 =
	     (_32_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d1577 ^
	      9'h100) <
	     9'd107 ;
  assign _32_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d1580 =
	     (_32_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d1577 ^
	      9'h100) <
	     9'd130 ;
  assign _32_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d2558 =
	     (12'd32 -
	      { 6'd0,
		IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2555 }) -
	     12'd1 ;
  assign _32_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d2559 =
	     (_32_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d2558 ^
	      12'h800) <=
	     12'd3071 ;
  assign _32_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d2560 =
	     (_32_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d2558 ^
	      12'h800) <
	     12'd974 ;
  assign _32_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d2561 =
	     (_32_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d2558 ^
	      12'h800) <
	     12'd1026 ;
  assign _3970_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_21_ETC___d4541 =
	     12'd3970 -
	     { 7'd0,
	       sV1_sfd__h1473[22] ?
		 5'd0 :
		 (sV1_sfd__h1473[21] ?
		    5'd1 :
		    (sV1_sfd__h1473[20] ?
		       5'd2 :
		       (sV1_sfd__h1473[19] ?
			  5'd3 :
			  (sV1_sfd__h1473[18] ?
			     5'd4 :
			     (sV1_sfd__h1473[17] ?
				5'd5 :
				(sV1_sfd__h1473[16] ?
				   5'd6 :
				   (sV1_sfd__h1473[15] ?
				      5'd7 :
				      (sV1_sfd__h1473[14] ?
					 5'd8 :
					 (sV1_sfd__h1473[13] ?
					    5'd9 :
					    (sV1_sfd__h1473[12] ?
					       5'd10 :
					       (sV1_sfd__h1473[11] ?
						  5'd11 :
						  (sV1_sfd__h1473[10] ?
						     5'd12 :
						     (sV1_sfd__h1473[9] ?
							5'd13 :
							(sV1_sfd__h1473[8] ?
							   5'd14 :
							   (sV1_sfd__h1473[7] ?
							      5'd15 :
							      (sV1_sfd__h1473[6] ?
								 5'd16 :
								 (sV1_sfd__h1473[5] ?
								    5'd17 :
								    (sV1_sfd__h1473[4] ?
								       5'd18 :
								       (sV1_sfd__h1473[3] ?
									  5'd19 :
									  (sV1_sfd__h1473[2] ?
									     5'd20 :
									     (sV1_sfd__h1473[1] ?
										5'd21 :
										(sV1_sfd__h1473[0] ?
										   5'd22 :
										   5'd23)))))))))))))))))))))) } ;
  assign _3970_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_21_ETC___d4542 =
	     (_3970_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_21_ETC___d4541 ^
	      12'h800) <=
	     12'd3071 ;
  assign _3970_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_21_ETC___d4543 =
	     (_3970_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_21_ETC___d4541 ^
	      12'h800) <
	     12'd1026 ;
  assign _3970_MINUS_SEXT_IF_requestR_3_BIT_214_4_THEN_r_ETC___d3854 =
	     12'd3970 -
	     SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_3_B_ETC___d3851 ;
  assign _64_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d2882 =
	     (12'd64 -
	      { 5'd0,
		IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3__ETC___d441 }) -
	     12'd1 ;
  assign _64_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d2883 =
	     (_64_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d2882 ^
	      12'h800) <=
	     12'd3071 ;
  assign _64_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d2885 =
	     (_64_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d2882 ^
	      12'h800) <
	     12'd974 ;
  assign _64_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d2888 =
	     (_64_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d2882 ^
	      12'h800) <
	     12'd1026 ;
  assign _64_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d444 =
	     (9'd64 -
	      { 2'd0,
		IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3__ETC___d441 }) -
	     9'd1 ;
  assign _64_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d445 =
	     (_64_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d444 ^
	      9'h100) <=
	     9'd383 ;
  assign _64_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d447 =
	     (_64_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d444 ^
	      9'h100) <
	     9'd107 ;
  assign _64_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d450 =
	     (_64_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d444 ^
	      9'h100) <
	     9'd130 ;
  assign _64_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d3068 =
	     (12'd64 -
	      { 5'd0,
		IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d966 }) -
	     12'd1 ;
  assign _64_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d3069 =
	     (_64_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d3068 ^
	      12'h800) <=
	     12'd3071 ;
  assign _64_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d3070 =
	     (_64_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d3068 ^
	      12'h800) <
	     12'd974 ;
  assign _64_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d3071 =
	     (_64_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d3068 ^
	      12'h800) <
	     12'd1026 ;
  assign _64_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d969 =
	     (9'd64 -
	      { 2'd0,
		IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d966 }) -
	     9'd1 ;
  assign _64_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d970 =
	     (_64_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d969 ^
	      9'h100) <=
	     9'd383 ;
  assign _64_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d971 =
	     (_64_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d969 ^
	      9'h100) <
	     9'd107 ;
  assign _64_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d972 =
	     (_64_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d969 ^
	      9'h100) <
	     9'd130 ;
  assign _theResult_____2__h110357 =
	     IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d3241 ?
	       out1___1__h111073 :
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d3224[117:53] ;
  assign _theResult_____2__h43093 =
	     IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1774 ?
	       out1___1__h43809 :
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1757[88:24] ;
  assign _theResult_____2__h45956 =
	     IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1925 ?
	       out1___1__h46448 :
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1908[56:24] ;
  assign _theResult_____2__h82460 =
	     IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2748 ?
	       out1___1__h82952 :
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2731[85:53] ;
  assign _theResult____h126028 =
	     (value__h82527 == 54'd0) ? sfd__h117253 : 57'd1 ;
  assign _theResult____h146240 =
	     ((_3970_MINUS_SEXT_IF_requestR_3_BIT_214_4_THEN_r_ETC___d3854 ^
	       12'h800) <
	      12'd2105) ?
	       result__h146853 :
	       _theResult____h126028 ;
  assign _theResult____h191843 =
	     ((_3074_MINUS_SEXT_IF_IF_requestR_3_BIT_214_4_THE_ETC___d4687 ^
	       12'h800) <
	      12'd2105) ?
	       result__h192456 :
	       ((value__h43160 == 25'd0) ? b__h46021 : 57'd1) ;
  assign _theResult___exp__h108862 =
	     (sfd__h108263[53] || sfd__h108263[53:52] == 2'b01) ?
	       11'd1 :
	       11'd0 ;
  assign _theResult___exp__h109617 =
	     sfd__h109005[53] ?
	       ((x__h108990[10:0] == 11'd2046) ?
		  11'd2047 :
		  din_inc___2_exp__h109755) :
	       ((x__h108990[10:0] == 11'd0 && sfd__h109005[53:52] == 2'b01) ?
		  11'd1 :
		  x__h108990[10:0]) ;
  assign _theResult___exp__h135916 =
	     sfd__h135482[24] ?
	       ((_theResult___fst_exp__h135390 == 8'd254) ?
		  8'd255 :
		  din_inc___2_exp__h166288) :
	       ((_theResult___fst_exp__h135390 == 8'd0 &&
		 sfd__h135482[24:23] == 2'b01) ?
		  8'd1 :
		  _theResult___fst_exp__h135390) ;
  assign _theResult___exp__h145761 =
	     sfd__h145327[24] ?
	       ((_theResult___fst_exp__h145309 == 8'd254) ?
		  8'd255 :
		  din_inc___2_exp__h166312) :
	       ((_theResult___fst_exp__h145309 == 8'd0 &&
		 sfd__h145327[24:23] == 2'b01) ?
		  8'd1 :
		  _theResult___fst_exp__h145309) ;
  assign _theResult___exp__h15431 =
	     (sfd__h15032[24] || sfd__h15032[24:23] == 2'b01) ? 8'd1 : 8'd0 ;
  assign _theResult___exp__h156257 =
	     sfd__h155823[24] ?
	       ((_theResult___fst_exp__h155731 == 8'd254) ?
		  8'd255 :
		  din_inc___2_exp__h166342) :
	       ((_theResult___fst_exp__h155731 == 8'd0 &&
		 sfd__h155823[24:23] == 2'b01) ?
		  8'd1 :
		  _theResult___fst_exp__h155731) ;
  assign _theResult___exp__h15984 =
	     sfd__h15575[24] ?
	       ((x__h15560[7:0] == 8'd254) ?
		  8'd255 :
		  din_inc___2_exp__h16127) :
	       ((x__h15560[7:0] == 8'd0 && sfd__h15575[24:23] == 2'b01) ?
		  8'd1 :
		  x__h15560[7:0]) ;
  assign _theResult___exp__h166156 =
	     sfd__h165698[24] ?
	       ((_theResult___fst_exp__h165679 == 8'd254) ?
		  8'd255 :
		  din_inc___2_exp__h166366) :
	       ((_theResult___fst_exp__h165679 == 8'd0 &&
		 sfd__h165698[24:23] == 2'b01) ?
		  8'd1 :
		  _theResult___fst_exp__h165679) ;
  assign _theResult___exp__h191161 =
	     sfd__h190524[53] ?
	       ((_theResult___fst_exp__h190506 == 11'd2046) ?
		  11'd2047 :
		  din_inc___2_exp__h212214) :
	       ((_theResult___fst_exp__h190506 == 11'd0 &&
		 sfd__h190524[53:52] == 2'b01) ?
		  11'd1 :
		  _theResult___fst_exp__h190506) ;
  assign _theResult___exp__h202063 =
	     sfd__h201426[53] ?
	       ((_theResult___fst_exp__h201334 == 11'd2046) ?
		  11'd2047 :
		  din_inc___2_exp__h212244) :
	       ((_theResult___fst_exp__h201334 == 11'd0 &&
		 sfd__h201426[53:52] == 2'b01) ?
		  11'd1 :
		  _theResult___fst_exp__h201334) ;
  assign _theResult___exp__h212078 =
	     sfd__h211417[53] ?
	       ((_theResult___fst_exp__h211398 == 11'd2046) ?
		  11'd2047 :
		  din_inc___2_exp__h212268) :
	       ((_theResult___fst_exp__h211398 == 11'd0 &&
		 sfd__h211417[53:52] == 2'b01) ?
		  11'd1 :
		  _theResult___fst_exp__h211398) ;
  assign _theResult___exp__h27709 =
	     (sfd__h27313[24] || sfd__h27313[24:23] == 2'b01) ? 8'd1 : 8'd0 ;
  assign _theResult___exp__h28261 =
	     sfd__h27852[24] ?
	       ((x__h27837[7:0] == 8'd254) ?
		  8'd255 :
		  din_inc___2_exp__h28399) :
	       ((x__h27837[7:0] == 8'd0 && sfd__h27852[24:23] == 2'b01) ?
		  8'd1 :
		  x__h27837[7:0]) ;
  assign _theResult___exp__h34881 =
	     (sfd__h34485[24] || sfd__h34485[24:23] == 2'b01) ? 8'd1 : 8'd0 ;
  assign _theResult___exp__h35434 =
	     sfd__h35025[24] ?
	       ((x__h35010[7:0] == 8'd254) ?
		  8'd255 :
		  din_inc___2_exp__h35577) :
	       ((x__h35010[7:0] == 8'd0 && sfd__h35025[24:23] == 2'b01) ?
		  8'd1 :
		  x__h35010[7:0]) ;
  assign _theResult___exp__h41797 =
	     (sfd__h41401[24] || sfd__h41401[24:23] == 2'b01) ? 8'd1 : 8'd0 ;
  assign _theResult___exp__h42349 =
	     sfd__h41940[24] ?
	       ((x__h41925[7:0] == 8'd254) ?
		  8'd255 :
		  din_inc___2_exp__h42487) :
	       ((x__h41925[7:0] == 8'd0 && sfd__h41940[24:23] == 2'b01) ?
		  8'd1 :
		  x__h41925[7:0]) ;
  assign _theResult___exp__h70015 =
	     (sfd__h69416[53] || sfd__h69416[53:52] == 2'b01) ?
	       11'd1 :
	       11'd0 ;
  assign _theResult___exp__h70771 =
	     sfd__h70159[53] ?
	       ((x__h70144[10:0] == 11'd2046) ?
		  11'd2047 :
		  din_inc___2_exp__h70914) :
	       ((x__h70144[10:0] == 11'd0 && sfd__h70159[53:52] == 2'b01) ?
		  11'd1 :
		  x__h70144[10:0]) ;
  assign _theResult___exp__h80962 =
	     (sfd__h80363[53] || sfd__h80363[53:52] == 2'b01) ?
	       11'd1 :
	       11'd0 ;
  assign _theResult___exp__h81717 =
	     sfd__h81105[53] ?
	       ((x__h81090[10:0] == 11'd2046) ?
		  11'd2047 :
		  din_inc___2_exp__h81855) :
	       ((x__h81090[10:0] == 11'd0 && sfd__h81105[53:52] == 2'b01) ?
		  11'd1 :
		  x__h81090[10:0]) ;
  assign _theResult___exp__h96337 =
	     (sfd__h95738[53] || sfd__h95738[53:52] == 2'b01) ?
	       11'd1 :
	       11'd0 ;
  assign _theResult___exp__h97093 =
	     sfd__h96481[53] ?
	       ((x__h96466[10:0] == 11'd2046) ?
		  11'd2047 :
		  din_inc___2_exp__h97236) :
	       ((x__h96466[10:0] == 11'd0 && sfd__h96481[53:52] == 2'b01) ?
		  11'd1 :
		  x__h96466[10:0]) ;
  assign _theResult___fst_exp__h108958 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       CASE_guard08246_0b0_0_0b1_0_0b10_out_exp08865__ETC__q32 :
	       CASE_requestR_BITS_194_TO_192_0x3_IF_guard0824_ETC__q34 ;
  assign _theResult___fst_exp__h109713 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       CASE_guard08975_0b0_x08990_BITS_10_TO_0_0b1_x0_ETC__q110 :
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d3147 ;
  assign _theResult___fst_exp__h109716 =
	     (x__h108990[10:0] == 11'd2047) ?
	       x__h108990[10:0] :
	       _theResult___fst_exp__h109713 ;
  assign _theResult___fst_exp__h126010 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3) ?
	       8'd255 :
	       CASE_requestR_BITS_194_TO_192_0x1_254_0x2_IF_r_ETC__q4 ;
  assign _theResult___fst_exp__h135390 =
	     _theResult____h126028[56] ?
	       8'd2 :
	       _theResult___fst_exp__h135464 ;
  assign _theResult___fst_exp__h135455 =
	     8'd0 -
	     { 2'd0,
	       IF_IF_0b0_CONCAT_NOT_IF_requestR_3_BIT_214_4_T_ETC___d3654 } ;
  assign _theResult___fst_exp__h135461 =
	     (!_theResult____h126028[56] && !_theResult____h126028[55] &&
	      !_theResult____h126028[54] &&
	      !_theResult____h126028[53] &&
	      !_theResult____h126028[52] &&
	      !_theResult____h126028[51] &&
	      !_theResult____h126028[50] &&
	      !_theResult____h126028[49] &&
	      !_theResult____h126028[48] &&
	      !_theResult____h126028[47] &&
	      !_theResult____h126028[46] &&
	      !_theResult____h126028[45] &&
	      !_theResult____h126028[44] &&
	      !_theResult____h126028[43] &&
	      !_theResult____h126028[42] &&
	      !_theResult____h126028[41] &&
	      !_theResult____h126028[40] &&
	      !_theResult____h126028[39] &&
	      !_theResult____h126028[38] &&
	      !_theResult____h126028[37] &&
	      !_theResult____h126028[36] &&
	      !_theResult____h126028[35] &&
	      !_theResult____h126028[34] &&
	      !_theResult____h126028[33] &&
	      !_theResult____h126028[32] &&
	      !_theResult____h126028[31] &&
	      !_theResult____h126028[30] &&
	      !_theResult____h126028[29] &&
	      !_theResult____h126028[28] &&
	      !_theResult____h126028[27] &&
	      !_theResult____h126028[26] &&
	      !_theResult____h126028[25] &&
	      !_theResult____h126028[24] &&
	      !_theResult____h126028[23] &&
	      !_theResult____h126028[22] &&
	      !_theResult____h126028[21] &&
	      !_theResult____h126028[20] &&
	      !_theResult____h126028[19] &&
	      !_theResult____h126028[18] &&
	      !_theResult____h126028[17] &&
	      !_theResult____h126028[16] &&
	      !_theResult____h126028[15] &&
	      !_theResult____h126028[14] &&
	      !_theResult____h126028[13] &&
	      !_theResult____h126028[12] &&
	      !_theResult____h126028[11] &&
	      !_theResult____h126028[10] &&
	      !_theResult____h126028[9] &&
	      !_theResult____h126028[8] &&
	      !_theResult____h126028[7] &&
	      !_theResult____h126028[6] &&
	      !_theResult____h126028[5] &&
	      !_theResult____h126028[4] &&
	      !_theResult____h126028[3] &&
	      !_theResult____h126028[2] &&
	      !_theResult____h126028[1] &&
	      !_theResult____h126028[0] ||
	      !_0_CONCAT_IF_IF_0b0_CONCAT_NOT_IF_requestR_3_BI_ETC___d3656) ?
	       8'd0 :
	       _theResult___fst_exp__h135455 ;
  assign _theResult___fst_exp__h135464 =
	     (!_theResult____h126028[56] && _theResult____h126028[55]) ?
	       8'd1 :
	       _theResult___fst_exp__h135461 ;
  assign _theResult___fst_exp__h136014 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       CASE_guard26038_0b0_theResult___fst_exp35390_0_ETC__q128 :
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d3719 ;
  assign _theResult___fst_exp__h136017 =
	     (_theResult___fst_exp__h135390 == 8'd255) ?
	       _theResult___fst_exp__h135390 :
	       _theResult___fst_exp__h136014 ;
  assign _theResult___fst_exp__h145300 =
	     8'd129 -
	     { 2'd0,
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d3776 } ;
  assign _theResult___fst_exp__h145306 =
	     (requestR_BITS_191_TO_128__q1[62:52] == 11'd0 &&
	      !requestR_BITS_191_TO_128__q1[51] &&
	      !requestR_BITS_191_TO_128__q1[50] &&
	      !requestR_BITS_191_TO_128__q1[49] &&
	      !requestR_BITS_191_TO_128__q1[48] &&
	      !requestR_BITS_191_TO_128__q1[47] &&
	      !requestR_BITS_191_TO_128__q1[46] &&
	      !requestR_BITS_191_TO_128__q1[45] &&
	      !requestR_BITS_191_TO_128__q1[44] &&
	      !requestR_BITS_191_TO_128__q1[43] &&
	      !requestR_BITS_191_TO_128__q1[42] &&
	      !requestR_BITS_191_TO_128__q1[41] &&
	      !requestR_BITS_191_TO_128__q1[40] &&
	      !requestR_BITS_191_TO_128__q1[39] &&
	      !requestR_BITS_191_TO_128__q1[38] &&
	      !requestR_BITS_191_TO_128__q1[37] &&
	      !requestR_BITS_191_TO_128__q1[36] &&
	      !requestR_BITS_191_TO_128__q1[35] &&
	      !requestR_BITS_191_TO_128__q1[34] &&
	      !requestR_BITS_191_TO_128__q1[33] &&
	      !requestR_BITS_191_TO_128__q1[32] &&
	      !requestR_BITS_191_TO_128__q1[31] &&
	      !requestR_BITS_191_TO_128__q1[30] &&
	      !requestR_BITS_191_TO_128__q1[29] &&
	      !requestR_BITS_191_TO_128__q1[28] &&
	      !requestR_BITS_191_TO_128__q1[27] &&
	      !requestR_BITS_191_TO_128__q1[26] &&
	      !requestR_BITS_191_TO_128__q1[25] &&
	      !requestR_BITS_191_TO_128__q1[24] &&
	      !requestR_BITS_191_TO_128__q1[23] &&
	      !requestR_BITS_191_TO_128__q1[22] &&
	      !requestR_BITS_191_TO_128__q1[21] &&
	      !requestR_BITS_191_TO_128__q1[20] &&
	      !requestR_BITS_191_TO_128__q1[19] &&
	      !requestR_BITS_191_TO_128__q1[18] &&
	      !requestR_BITS_191_TO_128__q1[17] &&
	      !requestR_BITS_191_TO_128__q1[16] &&
	      !requestR_BITS_191_TO_128__q1[15] &&
	      !requestR_BITS_191_TO_128__q1[14] &&
	      !requestR_BITS_191_TO_128__q1[13] &&
	      !requestR_BITS_191_TO_128__q1[12] &&
	      !requestR_BITS_191_TO_128__q1[11] &&
	      !requestR_BITS_191_TO_128__q1[10] &&
	      !requestR_BITS_191_TO_128__q1[9] &&
	      !requestR_BITS_191_TO_128__q1[8] &&
	      !requestR_BITS_191_TO_128__q1[7] &&
	      !requestR_BITS_191_TO_128__q1[6] &&
	      !requestR_BITS_191_TO_128__q1[5] &&
	      !requestR_BITS_191_TO_128__q1[4] &&
	      !requestR_BITS_191_TO_128__q1[3] &&
	      !requestR_BITS_191_TO_128__q1[2] &&
	      !requestR_BITS_191_TO_128__q1[1] &&
	      !requestR_BITS_191_TO_128__q1[0] ||
	      !_0_CONCAT_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d3778) ?
	       8'd0 :
	       _theResult___fst_exp__h145300 ;
  assign _theResult___fst_exp__h145309 =
	     (requestR_BITS_191_TO_128__q1[62:52] == 11'd0) ?
	       _theResult___fst_exp__h145306 :
	       8'd129 ;
  assign _theResult___fst_exp__h145859 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       CASE_guard36028_0b0_theResult___fst_exp45309_0_ETC__q130 :
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d3836 ;
  assign _theResult___fst_exp__h145862 =
	     (_theResult___fst_exp__h145309 == 8'd255) ?
	       _theResult___fst_exp__h145309 :
	       _theResult___fst_exp__h145859 ;
  assign _theResult___fst_exp__h15528 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       CASE_guard5015_0b0_0_0b1_0_0b10_out_exp5434_0b_ETC__q18 :
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d536 ;
  assign _theResult___fst_exp__h155731 =
	     _theResult____h146240[56] ?
	       8'd2 :
	       _theResult___fst_exp__h155805 ;
  assign _theResult___fst_exp__h155796 =
	     8'd0 -
	     { 2'd0,
	       IF_IF_3970_MINUS_SEXT_IF_requestR_3_BIT_214_4__ETC___d4098 } ;
  assign _theResult___fst_exp__h155802 =
	     (!_theResult____h146240[56] && !_theResult____h146240[55] &&
	      !_theResult____h146240[54] &&
	      !_theResult____h146240[53] &&
	      !_theResult____h146240[52] &&
	      !_theResult____h146240[51] &&
	      !_theResult____h146240[50] &&
	      !_theResult____h146240[49] &&
	      !_theResult____h146240[48] &&
	      !_theResult____h146240[47] &&
	      !_theResult____h146240[46] &&
	      !_theResult____h146240[45] &&
	      !_theResult____h146240[44] &&
	      !_theResult____h146240[43] &&
	      !_theResult____h146240[42] &&
	      !_theResult____h146240[41] &&
	      !_theResult____h146240[40] &&
	      !_theResult____h146240[39] &&
	      !_theResult____h146240[38] &&
	      !_theResult____h146240[37] &&
	      !_theResult____h146240[36] &&
	      !_theResult____h146240[35] &&
	      !_theResult____h146240[34] &&
	      !_theResult____h146240[33] &&
	      !_theResult____h146240[32] &&
	      !_theResult____h146240[31] &&
	      !_theResult____h146240[30] &&
	      !_theResult____h146240[29] &&
	      !_theResult____h146240[28] &&
	      !_theResult____h146240[27] &&
	      !_theResult____h146240[26] &&
	      !_theResult____h146240[25] &&
	      !_theResult____h146240[24] &&
	      !_theResult____h146240[23] &&
	      !_theResult____h146240[22] &&
	      !_theResult____h146240[21] &&
	      !_theResult____h146240[20] &&
	      !_theResult____h146240[19] &&
	      !_theResult____h146240[18] &&
	      !_theResult____h146240[17] &&
	      !_theResult____h146240[16] &&
	      !_theResult____h146240[15] &&
	      !_theResult____h146240[14] &&
	      !_theResult____h146240[13] &&
	      !_theResult____h146240[12] &&
	      !_theResult____h146240[11] &&
	      !_theResult____h146240[10] &&
	      !_theResult____h146240[9] &&
	      !_theResult____h146240[8] &&
	      !_theResult____h146240[7] &&
	      !_theResult____h146240[6] &&
	      !_theResult____h146240[5] &&
	      !_theResult____h146240[4] &&
	      !_theResult____h146240[3] &&
	      !_theResult____h146240[2] &&
	      !_theResult____h146240[1] &&
	      !_theResult____h146240[0] ||
	      !_0_CONCAT_IF_IF_3970_MINUS_SEXT_IF_requestR_3_B_ETC___d4100) ?
	       8'd0 :
	       _theResult___fst_exp__h155796 ;
  assign _theResult___fst_exp__h155805 =
	     (!_theResult____h146240[56] && _theResult____h146240[55]) ?
	       8'd1 :
	       _theResult___fst_exp__h155802 ;
  assign _theResult___fst_exp__h156355 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       CASE_guard46250_0b0_theResult___fst_exp55731_0_ETC__q132 :
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d4163 ;
  assign _theResult___fst_exp__h156358 =
	     (_theResult___fst_exp__h155731 == 8'd255) ?
	       _theResult___fst_exp__h155731 :
	       _theResult___fst_exp__h156355 ;
  assign _theResult___fst_exp__h16081 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       CASE_guard5545_0b0_x5560_BITS_7_TO_0_0b1_x5560_ETC__q20 :
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d565 ;
  assign _theResult___fst_exp__h16084 =
	     (x__h15560[7:0] == 8'd255) ?
	       x__h15560[7:0] :
	       _theResult___fst_exp__h16081 ;
  assign _theResult___fst_exp__h165631 =
	     (SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_3_B_ETC__q121[7:0] ==
	      8'd0) ?
	       8'd1 :
	       SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_3_B_ETC__q121[7:0] ;
  assign _theResult___fst_exp__h165670 =
	     SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_3_B_ETC__q121[7:0] -
	     { 2'd0,
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d3776 } ;
  assign _theResult___fst_exp__h165676 =
	     (requestR_BITS_191_TO_128__q1[62:52] == 11'd0 &&
	      !requestR_BITS_191_TO_128__q1[51] &&
	      !requestR_BITS_191_TO_128__q1[50] &&
	      !requestR_BITS_191_TO_128__q1[49] &&
	      !requestR_BITS_191_TO_128__q1[48] &&
	      !requestR_BITS_191_TO_128__q1[47] &&
	      !requestR_BITS_191_TO_128__q1[46] &&
	      !requestR_BITS_191_TO_128__q1[45] &&
	      !requestR_BITS_191_TO_128__q1[44] &&
	      !requestR_BITS_191_TO_128__q1[43] &&
	      !requestR_BITS_191_TO_128__q1[42] &&
	      !requestR_BITS_191_TO_128__q1[41] &&
	      !requestR_BITS_191_TO_128__q1[40] &&
	      !requestR_BITS_191_TO_128__q1[39] &&
	      !requestR_BITS_191_TO_128__q1[38] &&
	      !requestR_BITS_191_TO_128__q1[37] &&
	      !requestR_BITS_191_TO_128__q1[36] &&
	      !requestR_BITS_191_TO_128__q1[35] &&
	      !requestR_BITS_191_TO_128__q1[34] &&
	      !requestR_BITS_191_TO_128__q1[33] &&
	      !requestR_BITS_191_TO_128__q1[32] &&
	      !requestR_BITS_191_TO_128__q1[31] &&
	      !requestR_BITS_191_TO_128__q1[30] &&
	      !requestR_BITS_191_TO_128__q1[29] &&
	      !requestR_BITS_191_TO_128__q1[28] &&
	      !requestR_BITS_191_TO_128__q1[27] &&
	      !requestR_BITS_191_TO_128__q1[26] &&
	      !requestR_BITS_191_TO_128__q1[25] &&
	      !requestR_BITS_191_TO_128__q1[24] &&
	      !requestR_BITS_191_TO_128__q1[23] &&
	      !requestR_BITS_191_TO_128__q1[22] &&
	      !requestR_BITS_191_TO_128__q1[21] &&
	      !requestR_BITS_191_TO_128__q1[20] &&
	      !requestR_BITS_191_TO_128__q1[19] &&
	      !requestR_BITS_191_TO_128__q1[18] &&
	      !requestR_BITS_191_TO_128__q1[17] &&
	      !requestR_BITS_191_TO_128__q1[16] &&
	      !requestR_BITS_191_TO_128__q1[15] &&
	      !requestR_BITS_191_TO_128__q1[14] &&
	      !requestR_BITS_191_TO_128__q1[13] &&
	      !requestR_BITS_191_TO_128__q1[12] &&
	      !requestR_BITS_191_TO_128__q1[11] &&
	      !requestR_BITS_191_TO_128__q1[10] &&
	      !requestR_BITS_191_TO_128__q1[9] &&
	      !requestR_BITS_191_TO_128__q1[8] &&
	      !requestR_BITS_191_TO_128__q1[7] &&
	      !requestR_BITS_191_TO_128__q1[6] &&
	      !requestR_BITS_191_TO_128__q1[5] &&
	      !requestR_BITS_191_TO_128__q1[4] &&
	      !requestR_BITS_191_TO_128__q1[3] &&
	      !requestR_BITS_191_TO_128__q1[2] &&
	      !requestR_BITS_191_TO_128__q1[1] &&
	      !requestR_BITS_191_TO_128__q1[0] ||
	      !_0_CONCAT_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d4173) ?
	       8'd0 :
	       _theResult___fst_exp__h165670 ;
  assign _theResult___fst_exp__h165679 =
	     (requestR_BITS_191_TO_128__q1[62:52] == 11'd0) ?
	       _theResult___fst_exp__h165676 :
	       _theResult___fst_exp__h165631 ;
  assign _theResult___fst_exp__h166254 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       CASE_guard56369_0b0_theResult___fst_exp65679_0_ETC__q134 :
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d4232 ;
  assign _theResult___fst_exp__h166257 =
	     (_theResult___fst_exp__h165679 == 8'd255) ?
	       _theResult___fst_exp__h165679 :
	       _theResult___fst_exp__h166254 ;
  assign _theResult___fst_exp__h166266 =
	     (requestR_BITS_191_TO_128__q1[62:52] == 11'd0) ?
	       (_3074_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_ETC___d3421 ?
		  _theResult___snd_fst_exp__h145865 :
		  _theResult___fst_exp__h126010) :
	       (SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_3_B_ETC___d3852 ?
		  _theResult___snd_fst_exp__h166260 :
		  _theResult___fst_exp__h126010) ;
  assign _theResult___fst_exp__h166269 =
	     (requestR_BITS_191_TO_128__q1[62:52] == 11'd0 &&
	      requestR_BITS_191_TO_128__q1[51:0] == 52'd0) ?
	       8'd0 :
	       _theResult___fst_exp__h166266 ;
  assign _theResult___fst_exp__h174200 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3) ?
	       11'd2047 :
	       CASE_requestR_BITS_194_TO_192_0x1_2046_0x2_IF__ETC__q6 ;
  assign _theResult___fst_exp__h190497 =
	     11'd897 -
	     { 5'd0,
	       IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3__ETC___d4613 } ;
  assign _theResult___fst_exp__h190503 =
	     IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d4617 ?
	       11'd0 :
	       _theResult___fst_exp__h190497 ;
  assign _theResult___fst_exp__h190506 =
	     (sV1_exp__h1472 == 8'd0) ?
	       _theResult___fst_exp__h190503 :
	       11'd897 ;
  assign _theResult___fst_exp__h191259 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       CASE_guard81312_0b0_theResult___fst_exp90506_0_ETC__q160 :
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d4673 ;
  assign _theResult___fst_exp__h191262 =
	     (_theResult___fst_exp__h190506 == 11'd2047) ?
	       _theResult___fst_exp__h190506 :
	       _theResult___fst_exp__h191259 ;
  assign _theResult___fst_exp__h201334 =
	     _theResult____h191843[56] ?
	       11'd2 :
	       _theResult___fst_exp__h201408 ;
  assign _theResult___fst_exp__h201399 =
	     11'd0 -
	     { 5'd0,
	       IF_IF_3074_MINUS_SEXT_IF_IF_requestR_3_BIT_214_ETC___d4933 } ;
  assign _theResult___fst_exp__h201405 =
	     (!_theResult____h191843[56] && !_theResult____h191843[55] &&
	      !_theResult____h191843[54] &&
	      !_theResult____h191843[53] &&
	      !_theResult____h191843[52] &&
	      !_theResult____h191843[51] &&
	      !_theResult____h191843[50] &&
	      !_theResult____h191843[49] &&
	      !_theResult____h191843[48] &&
	      !_theResult____h191843[47] &&
	      !_theResult____h191843[46] &&
	      !_theResult____h191843[45] &&
	      !_theResult____h191843[44] &&
	      !_theResult____h191843[43] &&
	      !_theResult____h191843[42] &&
	      !_theResult____h191843[41] &&
	      !_theResult____h191843[40] &&
	      !_theResult____h191843[39] &&
	      !_theResult____h191843[38] &&
	      !_theResult____h191843[37] &&
	      !_theResult____h191843[36] &&
	      !_theResult____h191843[35] &&
	      !_theResult____h191843[34] &&
	      !_theResult____h191843[33] &&
	      !_theResult____h191843[32] &&
	      !_theResult____h191843[31] &&
	      !_theResult____h191843[30] &&
	      !_theResult____h191843[29] &&
	      !_theResult____h191843[28] &&
	      !_theResult____h191843[27] &&
	      !_theResult____h191843[26] &&
	      !_theResult____h191843[25] &&
	      !_theResult____h191843[24] &&
	      !_theResult____h191843[23] &&
	      !_theResult____h191843[22] &&
	      !_theResult____h191843[21] &&
	      !_theResult____h191843[20] &&
	      !_theResult____h191843[19] &&
	      !_theResult____h191843[18] &&
	      !_theResult____h191843[17] &&
	      !_theResult____h191843[16] &&
	      !_theResult____h191843[15] &&
	      !_theResult____h191843[14] &&
	      !_theResult____h191843[13] &&
	      !_theResult____h191843[12] &&
	      !_theResult____h191843[11] &&
	      !_theResult____h191843[10] &&
	      !_theResult____h191843[9] &&
	      !_theResult____h191843[8] &&
	      !_theResult____h191843[7] &&
	      !_theResult____h191843[6] &&
	      !_theResult____h191843[5] &&
	      !_theResult____h191843[4] &&
	      !_theResult____h191843[3] &&
	      !_theResult____h191843[2] &&
	      !_theResult____h191843[1] &&
	      !_theResult____h191843[0] ||
	      !_0_CONCAT_IF_IF_3074_MINUS_SEXT_IF_IF_requestR__ETC___d4935) ?
	       11'd0 :
	       _theResult___fst_exp__h201399 ;
  assign _theResult___fst_exp__h201408 =
	     (!_theResult____h191843[56] && _theResult____h191843[55]) ?
	       11'd1 :
	       _theResult___fst_exp__h201405 ;
  assign _theResult___fst_exp__h202161 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       CASE_guard91853_0b0_theResult___fst_exp01334_0_ETC__q162 :
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d4998 ;
  assign _theResult___fst_exp__h202164 =
	     (_theResult___fst_exp__h201334 == 11'd2047) ?
	       _theResult___fst_exp__h201334 :
	       _theResult___fst_exp__h202161 ;
  assign _theResult___fst_exp__h211350 =
	     (SEXT_IF_IF_requestR_3_BIT_214_4_THEN_requestR__ETC__q153[10:0] ==
	      11'd0) ?
	       11'd1 :
	       SEXT_IF_IF_requestR_3_BIT_214_4_THEN_requestR__ETC__q153[10:0] ;
  assign _theResult___fst_exp__h211389 =
	     SEXT_IF_IF_requestR_3_BIT_214_4_THEN_requestR__ETC__q153[10:0] -
	     { 5'd0,
	       IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3__ETC___d4613 } ;
  assign _theResult___fst_exp__h211395 =
	     IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d5010 ?
	       11'd0 :
	       _theResult___fst_exp__h211389 ;
  assign _theResult___fst_exp__h211398 =
	     (sV1_exp__h1472 == 8'd0) ?
	       _theResult___fst_exp__h211395 :
	       _theResult___fst_exp__h211350 ;
  assign _theResult___fst_exp__h212176 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       CASE_guard02175_0b0_theResult___fst_exp11398_0_ETC__q164 :
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d5067 ;
  assign _theResult___fst_exp__h212179 =
	     (_theResult___fst_exp__h211398 == 11'd2047) ?
	       _theResult___fst_exp__h211398 :
	       _theResult___fst_exp__h212176 ;
  assign _theResult___fst_exp__h212188 =
	     (sV1_exp__h1472 == 8'd0) ?
	       (_3970_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_21_ETC___d4542 ?
		  _theResult___snd_fst_exp__h191265 :
		  _theResult___fst_exp__h174200) :
	       (SEXT_IF_IF_requestR_3_BIT_214_4_THEN_requestR__ETC___d4685 ?
		  _theResult___snd_fst_exp__h212182 :
		  _theResult___fst_exp__h174200) ;
  assign _theResult___fst_exp__h212191 =
	     (sV1_exp__h1472 == 8'd0 && sV1_sfd__h1473 == 23'd0) ?
	       11'd0 :
	       _theResult___fst_exp__h212188 ;
  assign _theResult___fst_exp__h27805 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       CASE_guard7296_0b0_0_0b1_0_0b10_out_exp7712_0b_ETC__q29 :
	       CASE_requestR_BITS_194_TO_192_0x3_IF_guard7296_ETC__q31 ;
  assign _theResult___fst_exp__h28357 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       CASE_guard7822_0b0_x7837_BITS_7_TO_0_0b1_x7837_ETC__q36 :
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1050 ;
  assign _theResult___fst_exp__h28360 =
	     (x__h27837[7:0] == 8'd255) ?
	       x__h27837[7:0] :
	       _theResult___fst_exp__h28357 ;
  assign _theResult___fst_exp__h34978 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       CASE_guard4468_0b0_0_0b1_0_0b10_out_exp4884_0b_ETC__q44 :
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1404 ;
  assign _theResult___fst_exp__h35531 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       CASE_guard4995_0b0_x5010_BITS_7_TO_0_0b1_x5010_ETC__q50 :
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1433 ;
  assign _theResult___fst_exp__h35534 =
	     (x__h35010[7:0] == 8'd255) ?
	       x__h35010[7:0] :
	       _theResult___fst_exp__h35531 ;
  assign _theResult___fst_exp__h41893 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       CASE_guard1384_0b0_0_0b1_0_0b10_out_exp1800_0b_ETC__q57 :
	       CASE_requestR_BITS_194_TO_192_0x3_IF_guard1384_ETC__q59 ;
  assign _theResult___fst_exp__h42445 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       CASE_guard1910_0b0_x1925_BITS_7_TO_0_0b1_x1925_ETC__q61 :
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1657 ;
  assign _theResult___fst_exp__h42448 =
	     (x__h41925[7:0] == 8'd255) ?
	       x__h41925[7:0] :
	       _theResult___fst_exp__h42445 ;
  assign _theResult___fst_exp__h70112 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       CASE_guard9399_0b0_0_0b1_0_0b10_out_exp0018_0b_ETC__q81 :
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2422 ;
  assign _theResult___fst_exp__h70868 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       CASE_guard0129_0b0_x0144_BITS_10_TO_0_0b1_x014_ETC__q77 :
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2451 ;
  assign _theResult___fst_exp__h70871 =
	     (x__h70144[10:0] == 11'd2047) ?
	       x__h70144[10:0] :
	       _theResult___fst_exp__h70868 ;
  assign _theResult___fst_exp__h81058 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       CASE_guard0346_0b0_0_0b1_0_0b10_out_exp0965_0b_ETC__q86 :
	       CASE_requestR_BITS_194_TO_192_0x3_IF_guard0346_ETC__q88 ;
  assign _theResult___fst_exp__h81813 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       CASE_guard1075_0b0_x1090_BITS_10_TO_0_0b1_x109_ETC__q90 :
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2639 ;
  assign _theResult___fst_exp__h81816 =
	     (x__h81090[10:0] == 11'd2047) ?
	       x__h81090[10:0] :
	       _theResult___fst_exp__h81813 ;
  assign _theResult___fst_exp__h96434 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       CASE_guard5721_0b0_0_0b1_0_0b10_out_exp6340_0b_ETC__q106 :
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2961 ;
  assign _theResult___fst_exp__h97190 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       CASE_guard6451_0b0_x6466_BITS_10_TO_0_0b1_x646_ETC__q102 :
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2990 ;
  assign _theResult___fst_exp__h97193 =
	     (x__h96466[10:0] == 11'd2047) ?
	       x__h96466[10:0] :
	       _theResult___fst_exp__h97190 ;
  assign _theResult___fst_sfd__h108959 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       CASE_guard08246_0b0_sfd___37286_BITS_63_TO_12__ETC__q114 :
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d3170 ;
  assign _theResult___fst_sfd__h109714 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       CASE_guard08975_0b0_sfd___37286_BITS_62_TO_11__ETC__q112 :
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d3185 ;
  assign _theResult___fst_sfd__h109717 =
	     (x__h108990[10:0] == 11'd2047) ?
	       sfd___3__h27286[62:11] :
	       _theResult___fst_sfd__h109714 ;
  assign _theResult___fst_sfd__h113549 =
	     { 1'd1, requestR_BITS_191_TO_128__q1[50:0] } ;
  assign _theResult___fst_sfd__h126011 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3) ?
	       23'd0 :
	       CASE_requestR_BITS_194_TO_192_0x1_8388607_0x2__ETC__q5 ;
  assign _theResult___fst_sfd__h136015 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       CASE_guard26038_0b0_sfdin35384_BITS_56_TO_34_0_ETC__q136 :
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d4266 ;
  assign _theResult___fst_sfd__h136018 =
	     (_theResult___fst_exp__h135390 == 8'd255) ?
	       sfdin__h135384[56:34] :
	       _theResult___fst_sfd__h136015 ;
  assign _theResult___fst_sfd__h145860 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       CASE_guard36028_0b0_theResult___snd45260_BITS__ETC__q138 :
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d4285 ;
  assign _theResult___fst_sfd__h145863 =
	     (_theResult___fst_exp__h145309 == 8'd255) ?
	       _theResult___snd__h145260[56:34] :
	       _theResult___fst_sfd__h145860 ;
  assign _theResult___fst_sfd__h15529 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       CASE_guard5015_0b0_sfd___35005_BITS_63_TO_41_0_ETC__q22 :
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d588 ;
  assign _theResult___fst_sfd__h156356 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       CASE_guard46250_0b0_sfdin55725_BITS_56_TO_34_0_ETC__q140 :
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d4312 ;
  assign _theResult___fst_sfd__h156359 =
	     (_theResult___fst_exp__h155731 == 8'd255) ?
	       sfdin__h155725[56:34] :
	       _theResult___fst_sfd__h156356 ;
  assign _theResult___fst_sfd__h16082 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       CASE_guard5545_0b0_sfd___35005_BITS_62_TO_40_0_ETC__q24 :
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d606 ;
  assign _theResult___fst_sfd__h16085 =
	     (x__h15560[7:0] == 8'd255) ?
	       sfd___3__h15005[62:40] :
	       _theResult___fst_sfd__h16082 ;
  assign _theResult___fst_sfd__h166255 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       CASE_guard56369_0b0_theResult___snd65625_BITS__ETC__q142 :
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d4331 ;
  assign _theResult___fst_sfd__h166258 =
	     (_theResult___fst_exp__h165679 == 8'd255) ?
	       _theResult___snd__h165625[56:34] :
	       _theResult___fst_sfd__h166255 ;
  assign _theResult___fst_sfd__h166267 =
	     (requestR_BITS_191_TO_128__q1[62:52] == 11'd0) ?
	       (_3074_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_ETC___d3421 ?
		  _theResult___snd_fst_sfd__h145866 :
		  _theResult___fst_sfd__h126011) :
	       (SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_3_B_ETC___d3852 ?
		  _theResult___snd_fst_sfd__h166261 :
		  _theResult___fst_sfd__h126011) ;
  assign _theResult___fst_sfd__h166273 =
	     ((requestR_BITS_191_TO_128__q1[62:52] == 11'd2047 ||
	       requestR_BITS_191_TO_128__q1[62:52] == 11'd0) &&
	      requestR_BITS_191_TO_128__q1[51:0] == 52'd0) ?
	       23'd0 :
	       _theResult___fst_sfd__h166267 ;
  assign _theResult___fst_sfd__h168212 = { 1'd1, sV1_sfd__h1473[21:0] } ;
  assign _theResult___fst_sfd__h174201 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3) ?
	       52'd0 :
	       CASE_requestR_BITS_194_TO_192_0x1_450359962737_ETC__q7 ;
  assign _theResult___fst_sfd__h191260 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       CASE_guard81312_0b0_theResult___snd90457_BITS__ETC__q172 :
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d5100 ;
  assign _theResult___fst_sfd__h191263 =
	     (_theResult___fst_exp__h190506 == 11'd2047) ?
	       _theResult___snd__h190457[56:5] :
	       _theResult___fst_sfd__h191260 ;
  assign _theResult___fst_sfd__h202162 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       CASE_guard91853_0b0_sfdin01328_BITS_56_TO_5_0b_ETC__q174 :
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d5127 ;
  assign _theResult___fst_sfd__h202165 =
	     (_theResult___fst_exp__h201334 == 11'd2047) ?
	       sfdin__h201328[56:5] :
	       _theResult___fst_sfd__h202162 ;
  assign _theResult___fst_sfd__h212177 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       CASE_guard02175_0b0_theResult___snd11344_BITS__ETC__q176 :
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d5146 ;
  assign _theResult___fst_sfd__h212180 =
	     (_theResult___fst_exp__h211398 == 11'd2047) ?
	       _theResult___snd__h211344[56:5] :
	       _theResult___fst_sfd__h212177 ;
  assign _theResult___fst_sfd__h212189 =
	     (sV1_exp__h1472 == 8'd0) ?
	       (_3970_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_21_ETC___d4542 ?
		  _theResult___snd_fst_sfd__h191266 :
		  _theResult___fst_sfd__h174201) :
	       (SEXT_IF_IF_requestR_3_BIT_214_4_THEN_requestR__ETC___d4685 ?
		  _theResult___snd_fst_sfd__h212183 :
		  _theResult___fst_sfd__h174201) ;
  assign _theResult___fst_sfd__h212195 =
	     ((sV1_exp__h1472 == 8'd255 || sV1_exp__h1472 == 8'd0) &&
	      sV1_sfd__h1473 == 23'd0) ?
	       52'd0 :
	       _theResult___fst_sfd__h212189 ;
  assign _theResult___fst_sfd__h27806 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       CASE_guard7296_0b0_sfd___37286_BITS_63_TO_41_0_ETC__q40 :
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1073 ;
  assign _theResult___fst_sfd__h28358 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       CASE_guard7822_0b0_sfd___37286_BITS_62_TO_40_0_ETC__q38 :
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1088 ;
  assign _theResult___fst_sfd__h28361 =
	     (x__h27837[7:0] == 8'd255) ?
	       sfd___3__h27286[62:40] :
	       _theResult___fst_sfd__h28358 ;
  assign _theResult___fst_sfd__h34979 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       CASE_guard4468_0b0_sfd___34458_BITS_31_TO_9_0b_ETC__q52 :
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1456 ;
  assign _theResult___fst_sfd__h35532 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       CASE_guard4995_0b0_sfd___34458_BITS_30_TO_8_0b_ETC__q54 :
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1474 ;
  assign _theResult___fst_sfd__h35535 =
	     (x__h35010[7:0] == 8'd255) ?
	       sfd___3__h34458[30:8] :
	       _theResult___fst_sfd__h35532 ;
  assign _theResult___fst_sfd__h41894 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       CASE_guard1384_0b0_sfd___31374_BITS_31_TO_9_0b_ETC__q65 :
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1680 ;
  assign _theResult___fst_sfd__h42446 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       CASE_guard1910_0b0_sfd___31374_BITS_30_TO_8_0b_ETC__q63 :
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1695 ;
  assign _theResult___fst_sfd__h42449 =
	     (x__h41925[7:0] == 8'd255) ?
	       sfd___3__h41374[30:8] :
	       _theResult___fst_sfd__h42446 ;
  assign _theResult___fst_sfd__h70113 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       CASE_guard9399_0b0_sfd___39389_BITS_54_TO_3_0b_ETC__q83 :
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2474 ;
  assign _theResult___fst_sfd__h70869 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       CASE_guard0129_0b0_sfd___39389_BITS_53_TO_2_0b_ETC__q79 :
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2492 ;
  assign _theResult___fst_sfd__h70872 =
	     (x__h70144[10:0] == 11'd2047) ?
	       sfd___3__h69389[53:2] :
	       _theResult___fst_sfd__h70869 ;
  assign _theResult___fst_sfd__h81059 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       CASE_guard0346_0b0_sfd___30336_BITS_54_TO_3_0b_ETC__q94 :
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2661 ;
  assign _theResult___fst_sfd__h81814 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       CASE_guard1075_0b0_sfd___30336_BITS_53_TO_2_0b_ETC__q92 :
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2676 ;
  assign _theResult___fst_sfd__h81817 =
	     (x__h81090[10:0] == 11'd2047) ?
	       sfd___3__h80336[53:2] :
	       _theResult___fst_sfd__h81814 ;
  assign _theResult___fst_sfd__h96435 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       CASE_guard5721_0b0_sfd___35005_BITS_63_TO_12_0_ETC__q108 :
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d3013 ;
  assign _theResult___fst_sfd__h97191 =
	     (requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	      requestR[194:192] != 3'h3 &&
	      requestR[194:192] != 3'h4) ?
	       CASE_guard6451_0b0_sfd___35005_BITS_62_TO_11_0_ETC__q104 :
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d3031 ;
  assign _theResult___fst_sfd__h97194 =
	     (x__h96466[10:0] == 11'd2047) ?
	       sfd___3__h15005[62:11] :
	       _theResult___fst_sfd__h97191 ;
  assign _theResult___sfd__h108863 =
	     sfd__h108263[53] ? sfd__h108263[52:1] : sfd__h108263[51:0] ;
  assign _theResult___sfd__h109618 =
	     sfd__h109005[53] ?
	       ((x__h108990[10:0] == 11'd2046) ? 52'd0 : sfd__h109005[52:1]) :
	       sfd__h109005[51:0] ;
  assign _theResult___sfd__h135917 =
	     sfd__h135482[24] ?
	       ((_theResult___fst_exp__h135390 == 8'd254) ?
		  23'd0 :
		  sfd__h135482[23:1]) :
	       sfd__h135482[22:0] ;
  assign _theResult___sfd__h145762 =
	     sfd__h145327[24] ?
	       ((_theResult___fst_exp__h145309 == 8'd254) ?
		  23'd0 :
		  sfd__h145327[23:1]) :
	       sfd__h145327[22:0] ;
  assign _theResult___sfd__h15432 =
	     sfd__h15032[24] ? sfd__h15032[23:1] : sfd__h15032[22:0] ;
  assign _theResult___sfd__h156258 =
	     sfd__h155823[24] ?
	       ((_theResult___fst_exp__h155731 == 8'd254) ?
		  23'd0 :
		  sfd__h155823[23:1]) :
	       sfd__h155823[22:0] ;
  assign _theResult___sfd__h15985 =
	     sfd__h15575[24] ?
	       ((x__h15560[7:0] == 8'd254) ? 23'd0 : sfd__h15575[23:1]) :
	       sfd__h15575[22:0] ;
  assign _theResult___sfd__h166157 =
	     sfd__h165698[24] ?
	       ((_theResult___fst_exp__h165679 == 8'd254) ?
		  23'd0 :
		  sfd__h165698[23:1]) :
	       sfd__h165698[22:0] ;
  assign _theResult___sfd__h191162 =
	     sfd__h190524[53] ?
	       ((_theResult___fst_exp__h190506 == 11'd2046) ?
		  52'd0 :
		  sfd__h190524[52:1]) :
	       sfd__h190524[51:0] ;
  assign _theResult___sfd__h202064 =
	     sfd__h201426[53] ?
	       ((_theResult___fst_exp__h201334 == 11'd2046) ?
		  52'd0 :
		  sfd__h201426[52:1]) :
	       sfd__h201426[51:0] ;
  assign _theResult___sfd__h212079 =
	     sfd__h211417[53] ?
	       ((_theResult___fst_exp__h211398 == 11'd2046) ?
		  52'd0 :
		  sfd__h211417[52:1]) :
	       sfd__h211417[51:0] ;
  assign _theResult___sfd__h27710 =
	     sfd__h27313[24] ? sfd__h27313[23:1] : sfd__h27313[22:0] ;
  assign _theResult___sfd__h28262 =
	     sfd__h27852[24] ?
	       ((x__h27837[7:0] == 8'd254) ? 23'd0 : sfd__h27852[23:1]) :
	       sfd__h27852[22:0] ;
  assign _theResult___sfd__h34882 =
	     sfd__h34485[24] ? sfd__h34485[23:1] : sfd__h34485[22:0] ;
  assign _theResult___sfd__h35435 =
	     sfd__h35025[24] ?
	       ((x__h35010[7:0] == 8'd254) ? 23'd0 : sfd__h35025[23:1]) :
	       sfd__h35025[22:0] ;
  assign _theResult___sfd__h41798 =
	     sfd__h41401[24] ? sfd__h41401[23:1] : sfd__h41401[22:0] ;
  assign _theResult___sfd__h42350 =
	     sfd__h41940[24] ?
	       ((x__h41925[7:0] == 8'd254) ? 23'd0 : sfd__h41940[23:1]) :
	       sfd__h41940[22:0] ;
  assign _theResult___sfd__h70016 =
	     sfd__h69416[53] ? sfd__h69416[52:1] : sfd__h69416[51:0] ;
  assign _theResult___sfd__h70772 =
	     sfd__h70159[53] ?
	       ((x__h70144[10:0] == 11'd2046) ? 52'd0 : sfd__h70159[52:1]) :
	       sfd__h70159[51:0] ;
  assign _theResult___sfd__h80963 =
	     sfd__h80363[53] ? sfd__h80363[52:1] : sfd__h80363[51:0] ;
  assign _theResult___sfd__h81718 =
	     sfd__h81105[53] ?
	       ((x__h81090[10:0] == 11'd2046) ? 52'd0 : sfd__h81105[52:1]) :
	       sfd__h81105[51:0] ;
  assign _theResult___sfd__h96338 =
	     sfd__h95738[53] ? sfd__h95738[52:1] : sfd__h95738[51:0] ;
  assign _theResult___sfd__h97094 =
	     sfd__h96481[53] ?
	       ((x__h96466[10:0] == 11'd2046) ? 52'd0 : sfd__h96481[52:1]) :
	       sfd__h96481[51:0] ;
  assign _theResult___snd__h135401 = { _theResult____h126028[55:0], 1'd0 } ;
  assign _theResult___snd__h135412 =
	     (!_theResult____h126028[56] && _theResult____h126028[55]) ?
	       _theResult___snd__h135414 :
	       _theResult___snd__h135424 ;
  assign _theResult___snd__h135414 = { _theResult____h126028[54:0], 2'd0 } ;
  assign _theResult___snd__h135424 =
	     (!_theResult____h126028[56] && !_theResult____h126028[55] &&
	      !_theResult____h126028[54] &&
	      !_theResult____h126028[53] &&
	      !_theResult____h126028[52] &&
	      !_theResult____h126028[51] &&
	      !_theResult____h126028[50] &&
	      !_theResult____h126028[49] &&
	      !_theResult____h126028[48] &&
	      !_theResult____h126028[47] &&
	      !_theResult____h126028[46] &&
	      !_theResult____h126028[45] &&
	      !_theResult____h126028[44] &&
	      !_theResult____h126028[43] &&
	      !_theResult____h126028[42] &&
	      !_theResult____h126028[41] &&
	      !_theResult____h126028[40] &&
	      !_theResult____h126028[39] &&
	      !_theResult____h126028[38] &&
	      !_theResult____h126028[37] &&
	      !_theResult____h126028[36] &&
	      !_theResult____h126028[35] &&
	      !_theResult____h126028[34] &&
	      !_theResult____h126028[33] &&
	      !_theResult____h126028[32] &&
	      !_theResult____h126028[31] &&
	      !_theResult____h126028[30] &&
	      !_theResult____h126028[29] &&
	      !_theResult____h126028[28] &&
	      !_theResult____h126028[27] &&
	      !_theResult____h126028[26] &&
	      !_theResult____h126028[25] &&
	      !_theResult____h126028[24] &&
	      !_theResult____h126028[23] &&
	      !_theResult____h126028[22] &&
	      !_theResult____h126028[21] &&
	      !_theResult____h126028[20] &&
	      !_theResult____h126028[19] &&
	      !_theResult____h126028[18] &&
	      !_theResult____h126028[17] &&
	      !_theResult____h126028[16] &&
	      !_theResult____h126028[15] &&
	      !_theResult____h126028[14] &&
	      !_theResult____h126028[13] &&
	      !_theResult____h126028[12] &&
	      !_theResult____h126028[11] &&
	      !_theResult____h126028[10] &&
	      !_theResult____h126028[9] &&
	      !_theResult____h126028[8] &&
	      !_theResult____h126028[7] &&
	      !_theResult____h126028[6] &&
	      !_theResult____h126028[5] &&
	      !_theResult____h126028[4] &&
	      !_theResult____h126028[3] &&
	      !_theResult____h126028[2] &&
	      !_theResult____h126028[1] &&
	      !_theResult____h126028[0]) ?
	       _theResult____h126028 :
	       _theResult___snd__h135430 ;
  assign _theResult___snd__h135430 =
	     { IF_0_CONCAT_IF_IF_0b0_CONCAT_NOT_IF_requestR_3_ETC__q117[54:0],
	       2'd0 } ;
  assign _theResult___snd__h135453 =
	     _theResult____h126028 <<
	     IF_IF_0b0_CONCAT_NOT_IF_requestR_3_BIT_214_4_T_ETC___d3654 ;
  assign _theResult___snd__h145260 =
	     (requestR_BITS_191_TO_128__q1[62:52] == 11'd0) ?
	       _theResult___snd__h145269 :
	       _theResult___snd__h145262 ;
  assign _theResult___snd__h145262 =
	     { requestR_BITS_191_TO_128__q1[51:0], 5'd0 } ;
  assign _theResult___snd__h145269 =
	     (requestR_BITS_191_TO_128__q1[62:52] == 11'd0 &&
	      !requestR_BITS_191_TO_128__q1[51] &&
	      !requestR_BITS_191_TO_128__q1[50] &&
	      !requestR_BITS_191_TO_128__q1[49] &&
	      !requestR_BITS_191_TO_128__q1[48] &&
	      !requestR_BITS_191_TO_128__q1[47] &&
	      !requestR_BITS_191_TO_128__q1[46] &&
	      !requestR_BITS_191_TO_128__q1[45] &&
	      !requestR_BITS_191_TO_128__q1[44] &&
	      !requestR_BITS_191_TO_128__q1[43] &&
	      !requestR_BITS_191_TO_128__q1[42] &&
	      !requestR_BITS_191_TO_128__q1[41] &&
	      !requestR_BITS_191_TO_128__q1[40] &&
	      !requestR_BITS_191_TO_128__q1[39] &&
	      !requestR_BITS_191_TO_128__q1[38] &&
	      !requestR_BITS_191_TO_128__q1[37] &&
	      !requestR_BITS_191_TO_128__q1[36] &&
	      !requestR_BITS_191_TO_128__q1[35] &&
	      !requestR_BITS_191_TO_128__q1[34] &&
	      !requestR_BITS_191_TO_128__q1[33] &&
	      !requestR_BITS_191_TO_128__q1[32] &&
	      !requestR_BITS_191_TO_128__q1[31] &&
	      !requestR_BITS_191_TO_128__q1[30] &&
	      !requestR_BITS_191_TO_128__q1[29] &&
	      !requestR_BITS_191_TO_128__q1[28] &&
	      !requestR_BITS_191_TO_128__q1[27] &&
	      !requestR_BITS_191_TO_128__q1[26] &&
	      !requestR_BITS_191_TO_128__q1[25] &&
	      !requestR_BITS_191_TO_128__q1[24] &&
	      !requestR_BITS_191_TO_128__q1[23] &&
	      !requestR_BITS_191_TO_128__q1[22] &&
	      !requestR_BITS_191_TO_128__q1[21] &&
	      !requestR_BITS_191_TO_128__q1[20] &&
	      !requestR_BITS_191_TO_128__q1[19] &&
	      !requestR_BITS_191_TO_128__q1[18] &&
	      !requestR_BITS_191_TO_128__q1[17] &&
	      !requestR_BITS_191_TO_128__q1[16] &&
	      !requestR_BITS_191_TO_128__q1[15] &&
	      !requestR_BITS_191_TO_128__q1[14] &&
	      !requestR_BITS_191_TO_128__q1[13] &&
	      !requestR_BITS_191_TO_128__q1[12] &&
	      !requestR_BITS_191_TO_128__q1[11] &&
	      !requestR_BITS_191_TO_128__q1[10] &&
	      !requestR_BITS_191_TO_128__q1[9] &&
	      !requestR_BITS_191_TO_128__q1[8] &&
	      !requestR_BITS_191_TO_128__q1[7] &&
	      !requestR_BITS_191_TO_128__q1[6] &&
	      !requestR_BITS_191_TO_128__q1[5] &&
	      !requestR_BITS_191_TO_128__q1[4] &&
	      !requestR_BITS_191_TO_128__q1[3] &&
	      !requestR_BITS_191_TO_128__q1[2] &&
	      !requestR_BITS_191_TO_128__q1[1] &&
	      !requestR_BITS_191_TO_128__q1[0]) ?
	       sfd__h117253 :
	       _theResult___snd__h145275 ;
  assign _theResult___snd__h145275 =
	     { IF_0_CONCAT_IF_IF_requestR_3_BIT_214_4_THEN_re_ETC__q119[54:0],
	       2'd0 } ;
  assign _theResult___snd__h145298 =
	     sfd__h117253 <<
	     IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d3776 ;
  assign _theResult___snd__h155742 = { _theResult____h146240[55:0], 1'd0 } ;
  assign _theResult___snd__h155753 =
	     (!_theResult____h146240[56] && _theResult____h146240[55]) ?
	       _theResult___snd__h155755 :
	       _theResult___snd__h155765 ;
  assign _theResult___snd__h155755 = { _theResult____h146240[54:0], 2'd0 } ;
  assign _theResult___snd__h155765 =
	     (!_theResult____h146240[56] && !_theResult____h146240[55] &&
	      !_theResult____h146240[54] &&
	      !_theResult____h146240[53] &&
	      !_theResult____h146240[52] &&
	      !_theResult____h146240[51] &&
	      !_theResult____h146240[50] &&
	      !_theResult____h146240[49] &&
	      !_theResult____h146240[48] &&
	      !_theResult____h146240[47] &&
	      !_theResult____h146240[46] &&
	      !_theResult____h146240[45] &&
	      !_theResult____h146240[44] &&
	      !_theResult____h146240[43] &&
	      !_theResult____h146240[42] &&
	      !_theResult____h146240[41] &&
	      !_theResult____h146240[40] &&
	      !_theResult____h146240[39] &&
	      !_theResult____h146240[38] &&
	      !_theResult____h146240[37] &&
	      !_theResult____h146240[36] &&
	      !_theResult____h146240[35] &&
	      !_theResult____h146240[34] &&
	      !_theResult____h146240[33] &&
	      !_theResult____h146240[32] &&
	      !_theResult____h146240[31] &&
	      !_theResult____h146240[30] &&
	      !_theResult____h146240[29] &&
	      !_theResult____h146240[28] &&
	      !_theResult____h146240[27] &&
	      !_theResult____h146240[26] &&
	      !_theResult____h146240[25] &&
	      !_theResult____h146240[24] &&
	      !_theResult____h146240[23] &&
	      !_theResult____h146240[22] &&
	      !_theResult____h146240[21] &&
	      !_theResult____h146240[20] &&
	      !_theResult____h146240[19] &&
	      !_theResult____h146240[18] &&
	      !_theResult____h146240[17] &&
	      !_theResult____h146240[16] &&
	      !_theResult____h146240[15] &&
	      !_theResult____h146240[14] &&
	      !_theResult____h146240[13] &&
	      !_theResult____h146240[12] &&
	      !_theResult____h146240[11] &&
	      !_theResult____h146240[10] &&
	      !_theResult____h146240[9] &&
	      !_theResult____h146240[8] &&
	      !_theResult____h146240[7] &&
	      !_theResult____h146240[6] &&
	      !_theResult____h146240[5] &&
	      !_theResult____h146240[4] &&
	      !_theResult____h146240[3] &&
	      !_theResult____h146240[2] &&
	      !_theResult____h146240[1] &&
	      !_theResult____h146240[0]) ?
	       _theResult____h146240 :
	       _theResult___snd__h155771 ;
  assign _theResult___snd__h155771 =
	     { IF_0_CONCAT_IF_IF_3970_MINUS_SEXT_IF_requestR__ETC__q122[54:0],
	       2'd0 } ;
  assign _theResult___snd__h155794 =
	     _theResult____h146240 <<
	     IF_IF_3970_MINUS_SEXT_IF_requestR_3_BIT_214_4__ETC___d4098 ;
  assign _theResult___snd__h165625 =
	     (requestR_BITS_191_TO_128__q1[62:52] == 11'd0) ?
	       _theResult___snd__h165639 :
	       _theResult___snd__h145262 ;
  assign _theResult___snd__h165639 =
	     (requestR_BITS_191_TO_128__q1[62:52] == 11'd0 &&
	      !requestR_BITS_191_TO_128__q1[51] &&
	      !requestR_BITS_191_TO_128__q1[50] &&
	      !requestR_BITS_191_TO_128__q1[49] &&
	      !requestR_BITS_191_TO_128__q1[48] &&
	      !requestR_BITS_191_TO_128__q1[47] &&
	      !requestR_BITS_191_TO_128__q1[46] &&
	      !requestR_BITS_191_TO_128__q1[45] &&
	      !requestR_BITS_191_TO_128__q1[44] &&
	      !requestR_BITS_191_TO_128__q1[43] &&
	      !requestR_BITS_191_TO_128__q1[42] &&
	      !requestR_BITS_191_TO_128__q1[41] &&
	      !requestR_BITS_191_TO_128__q1[40] &&
	      !requestR_BITS_191_TO_128__q1[39] &&
	      !requestR_BITS_191_TO_128__q1[38] &&
	      !requestR_BITS_191_TO_128__q1[37] &&
	      !requestR_BITS_191_TO_128__q1[36] &&
	      !requestR_BITS_191_TO_128__q1[35] &&
	      !requestR_BITS_191_TO_128__q1[34] &&
	      !requestR_BITS_191_TO_128__q1[33] &&
	      !requestR_BITS_191_TO_128__q1[32] &&
	      !requestR_BITS_191_TO_128__q1[31] &&
	      !requestR_BITS_191_TO_128__q1[30] &&
	      !requestR_BITS_191_TO_128__q1[29] &&
	      !requestR_BITS_191_TO_128__q1[28] &&
	      !requestR_BITS_191_TO_128__q1[27] &&
	      !requestR_BITS_191_TO_128__q1[26] &&
	      !requestR_BITS_191_TO_128__q1[25] &&
	      !requestR_BITS_191_TO_128__q1[24] &&
	      !requestR_BITS_191_TO_128__q1[23] &&
	      !requestR_BITS_191_TO_128__q1[22] &&
	      !requestR_BITS_191_TO_128__q1[21] &&
	      !requestR_BITS_191_TO_128__q1[20] &&
	      !requestR_BITS_191_TO_128__q1[19] &&
	      !requestR_BITS_191_TO_128__q1[18] &&
	      !requestR_BITS_191_TO_128__q1[17] &&
	      !requestR_BITS_191_TO_128__q1[16] &&
	      !requestR_BITS_191_TO_128__q1[15] &&
	      !requestR_BITS_191_TO_128__q1[14] &&
	      !requestR_BITS_191_TO_128__q1[13] &&
	      !requestR_BITS_191_TO_128__q1[12] &&
	      !requestR_BITS_191_TO_128__q1[11] &&
	      !requestR_BITS_191_TO_128__q1[10] &&
	      !requestR_BITS_191_TO_128__q1[9] &&
	      !requestR_BITS_191_TO_128__q1[8] &&
	      !requestR_BITS_191_TO_128__q1[7] &&
	      !requestR_BITS_191_TO_128__q1[6] &&
	      !requestR_BITS_191_TO_128__q1[5] &&
	      !requestR_BITS_191_TO_128__q1[4] &&
	      !requestR_BITS_191_TO_128__q1[3] &&
	      !requestR_BITS_191_TO_128__q1[2] &&
	      !requestR_BITS_191_TO_128__q1[1] &&
	      !requestR_BITS_191_TO_128__q1[0]) ?
	       sfd__h117253 :
	       _theResult___snd__h165645 ;
  assign _theResult___snd__h165645 =
	     { IF_0_CONCAT_IF_IF_requestR_3_BIT_214_4_THEN_re_ETC__q125[54:0],
	       2'd0 } ;
  assign _theResult___snd__h165663 =
	     sfd__h117253 <<
	     IF_SEXT_IF_requestR_3_BIT_214_4_THEN_requestR__ETC___d4172 ;
  assign _theResult___snd__h190457 =
	     (sV1_exp__h1472 == 8'd0) ?
	       _theResult___snd__h190466 :
	       _theResult___snd__h190459 ;
  assign _theResult___snd__h190459 = { sV1_sfd__h1473, 34'd0 } ;
  assign _theResult___snd__h190466 =
	     (sV1_exp__h1472 == 8'd0 && !sV1_sfd__h1473[22] &&
	      !sV1_sfd__h1473[21] &&
	      !sV1_sfd__h1473[20] &&
	      !sV1_sfd__h1473[19] &&
	      !sV1_sfd__h1473[18] &&
	      !sV1_sfd__h1473[17] &&
	      !sV1_sfd__h1473[16] &&
	      !sV1_sfd__h1473[15] &&
	      !sV1_sfd__h1473[14] &&
	      !sV1_sfd__h1473[13] &&
	      !sV1_sfd__h1473[12] &&
	      !sV1_sfd__h1473[11] &&
	      !sV1_sfd__h1473[10] &&
	      !sV1_sfd__h1473[9] &&
	      !sV1_sfd__h1473[8] &&
	      !sV1_sfd__h1473[7] &&
	      !sV1_sfd__h1473[6] &&
	      !sV1_sfd__h1473[5] &&
	      !sV1_sfd__h1473[4] &&
	      !sV1_sfd__h1473[3] &&
	      !sV1_sfd__h1473[2] &&
	      !sV1_sfd__h1473[1] &&
	      !sV1_sfd__h1473[0]) ?
	       b__h46021 :
	       _theResult___snd__h190472 ;
  assign _theResult___snd__h190472 =
	     { IF_0_CONCAT_IF_IF_IF_requestR_3_BIT_214_4_THEN_ETC__q151[54:0],
	       2'd0 } ;
  assign _theResult___snd__h190495 =
	     b__h46021 <<
	     IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3__ETC___d4613 ;
  assign _theResult___snd__h201345 = { _theResult____h191843[55:0], 1'd0 } ;
  assign _theResult___snd__h201356 =
	     (!_theResult____h191843[56] && _theResult____h191843[55]) ?
	       _theResult___snd__h201358 :
	       _theResult___snd__h201368 ;
  assign _theResult___snd__h201358 = { _theResult____h191843[54:0], 2'd0 } ;
  assign _theResult___snd__h201368 =
	     (!_theResult____h191843[56] && !_theResult____h191843[55] &&
	      !_theResult____h191843[54] &&
	      !_theResult____h191843[53] &&
	      !_theResult____h191843[52] &&
	      !_theResult____h191843[51] &&
	      !_theResult____h191843[50] &&
	      !_theResult____h191843[49] &&
	      !_theResult____h191843[48] &&
	      !_theResult____h191843[47] &&
	      !_theResult____h191843[46] &&
	      !_theResult____h191843[45] &&
	      !_theResult____h191843[44] &&
	      !_theResult____h191843[43] &&
	      !_theResult____h191843[42] &&
	      !_theResult____h191843[41] &&
	      !_theResult____h191843[40] &&
	      !_theResult____h191843[39] &&
	      !_theResult____h191843[38] &&
	      !_theResult____h191843[37] &&
	      !_theResult____h191843[36] &&
	      !_theResult____h191843[35] &&
	      !_theResult____h191843[34] &&
	      !_theResult____h191843[33] &&
	      !_theResult____h191843[32] &&
	      !_theResult____h191843[31] &&
	      !_theResult____h191843[30] &&
	      !_theResult____h191843[29] &&
	      !_theResult____h191843[28] &&
	      !_theResult____h191843[27] &&
	      !_theResult____h191843[26] &&
	      !_theResult____h191843[25] &&
	      !_theResult____h191843[24] &&
	      !_theResult____h191843[23] &&
	      !_theResult____h191843[22] &&
	      !_theResult____h191843[21] &&
	      !_theResult____h191843[20] &&
	      !_theResult____h191843[19] &&
	      !_theResult____h191843[18] &&
	      !_theResult____h191843[17] &&
	      !_theResult____h191843[16] &&
	      !_theResult____h191843[15] &&
	      !_theResult____h191843[14] &&
	      !_theResult____h191843[13] &&
	      !_theResult____h191843[12] &&
	      !_theResult____h191843[11] &&
	      !_theResult____h191843[10] &&
	      !_theResult____h191843[9] &&
	      !_theResult____h191843[8] &&
	      !_theResult____h191843[7] &&
	      !_theResult____h191843[6] &&
	      !_theResult____h191843[5] &&
	      !_theResult____h191843[4] &&
	      !_theResult____h191843[3] &&
	      !_theResult____h191843[2] &&
	      !_theResult____h191843[1] &&
	      !_theResult____h191843[0]) ?
	       _theResult____h191843 :
	       _theResult___snd__h201374 ;
  assign _theResult___snd__h201374 =
	     { IF_0_CONCAT_IF_IF_3074_MINUS_SEXT_IF_IF_reques_ETC__q154[54:0],
	       2'd0 } ;
  assign _theResult___snd__h201397 =
	     _theResult____h191843 <<
	     IF_IF_3074_MINUS_SEXT_IF_IF_requestR_3_BIT_214_ETC___d4933 ;
  assign _theResult___snd__h211344 =
	     (sV1_exp__h1472 == 8'd0) ?
	       _theResult___snd__h211358 :
	       _theResult___snd__h190459 ;
  assign _theResult___snd__h211358 =
	     (sV1_exp__h1472 == 8'd0 && !sV1_sfd__h1473[22] &&
	      !sV1_sfd__h1473[21] &&
	      !sV1_sfd__h1473[20] &&
	      !sV1_sfd__h1473[19] &&
	      !sV1_sfd__h1473[18] &&
	      !sV1_sfd__h1473[17] &&
	      !sV1_sfd__h1473[16] &&
	      !sV1_sfd__h1473[15] &&
	      !sV1_sfd__h1473[14] &&
	      !sV1_sfd__h1473[13] &&
	      !sV1_sfd__h1473[12] &&
	      !sV1_sfd__h1473[11] &&
	      !sV1_sfd__h1473[10] &&
	      !sV1_sfd__h1473[9] &&
	      !sV1_sfd__h1473[8] &&
	      !sV1_sfd__h1473[7] &&
	      !sV1_sfd__h1473[6] &&
	      !sV1_sfd__h1473[5] &&
	      !sV1_sfd__h1473[4] &&
	      !sV1_sfd__h1473[3] &&
	      !sV1_sfd__h1473[2] &&
	      !sV1_sfd__h1473[1] &&
	      !sV1_sfd__h1473[0]) ?
	       b__h46021 :
	       _theResult___snd__h211364 ;
  assign _theResult___snd__h211364 =
	     { IF_0_CONCAT_IF_IF_IF_requestR_3_BIT_214_4_THEN_ETC__q157[54:0],
	       2'd0 } ;
  assign _theResult___snd__h211382 =
	     b__h46021 <<
	     IF_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_reques_ETC___d5007 ;
  assign _theResult___snd_fst_exp__h109719 =
	     _64_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d3071 ?
	       _theResult___fst_exp__h108958 :
	       _theResult___fst_exp__h109716 ;
  assign _theResult___snd_fst_exp__h109722 =
	     _64_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d3070 ?
	       11'd0 :
	       _theResult___snd_fst_exp__h109719 ;
  assign _theResult___snd_fst_exp__h109725 =
	     _64_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d3069 ?
	       _theResult___snd_fst_exp__h109722 :
	       11'd2047 ;
  assign _theResult___snd_fst_exp__h145865 =
	     _3074_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_ETC___d3422 ?
	       _theResult___fst_exp__h136017 :
	       _theResult___fst_exp__h145862 ;
  assign _theResult___snd_fst_exp__h16087 =
	     _64_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d450 ?
	       _theResult___fst_exp__h15528 :
	       _theResult___fst_exp__h16084 ;
  assign _theResult___snd_fst_exp__h16090 =
	     _64_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d447 ?
	       8'd0 :
	       _theResult___snd_fst_exp__h16087 ;
  assign _theResult___snd_fst_exp__h16093 =
	     _64_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d445 ?
	       _theResult___snd_fst_exp__h16090 :
	       8'd255 ;
  assign _theResult___snd_fst_exp__h166260 =
	     SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_3_B_ETC___d3853 ?
	       _theResult___fst_exp__h156358 :
	       _theResult___fst_exp__h166257 ;
  assign _theResult___snd_fst_exp__h191265 =
	     _3970_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_21_ETC___d4543 ?
	       11'd0 :
	       _theResult___fst_exp__h191262 ;
  assign _theResult___snd_fst_exp__h212182 =
	     SEXT_IF_IF_requestR_3_BIT_214_4_THEN_requestR__ETC___d4686 ?
	       _theResult___fst_exp__h202164 :
	       _theResult___fst_exp__h212179 ;
  assign _theResult___snd_fst_exp__h28363 =
	     _64_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d972 ?
	       _theResult___fst_exp__h27805 :
	       _theResult___fst_exp__h28360 ;
  assign _theResult___snd_fst_exp__h28366 =
	     _64_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d971 ?
	       8'd0 :
	       _theResult___snd_fst_exp__h28363 ;
  assign _theResult___snd_fst_exp__h28369 =
	     _64_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d970 ?
	       _theResult___snd_fst_exp__h28366 :
	       8'd255 ;
  assign _theResult___snd_fst_exp__h35537 =
	     _32_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d1327 ?
	       _theResult___fst_exp__h34978 :
	       _theResult___fst_exp__h35534 ;
  assign _theResult___snd_fst_exp__h35540 =
	     _32_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d1324 ?
	       8'd0 :
	       _theResult___snd_fst_exp__h35537 ;
  assign _theResult___snd_fst_exp__h35543 =
	     _32_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d1322 ?
	       _theResult___snd_fst_exp__h35540 :
	       8'd255 ;
  assign _theResult___snd_fst_exp__h42451 =
	     _32_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d1580 ?
	       _theResult___fst_exp__h41893 :
	       _theResult___fst_exp__h42448 ;
  assign _theResult___snd_fst_exp__h42454 =
	     _32_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d1579 ?
	       8'd0 :
	       _theResult___snd_fst_exp__h42451 ;
  assign _theResult___snd_fst_exp__h42457 =
	     _32_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d1578 ?
	       _theResult___snd_fst_exp__h42454 :
	       8'd255 ;
  assign _theResult___snd_fst_exp__h70874 =
	     _32_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d2347 ?
	       _theResult___fst_exp__h70112 :
	       _theResult___fst_exp__h70871 ;
  assign _theResult___snd_fst_exp__h70877 =
	     _32_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d2345 ?
	       11'd0 :
	       _theResult___snd_fst_exp__h70874 ;
  assign _theResult___snd_fst_exp__h70880 =
	     _32_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d2343 ?
	       _theResult___snd_fst_exp__h70877 :
	       11'd2047 ;
  assign _theResult___snd_fst_exp__h81819 =
	     _32_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d2561 ?
	       _theResult___fst_exp__h81058 :
	       _theResult___fst_exp__h81816 ;
  assign _theResult___snd_fst_exp__h81822 =
	     _32_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d2560 ?
	       11'd0 :
	       _theResult___snd_fst_exp__h81819 ;
  assign _theResult___snd_fst_exp__h81825 =
	     _32_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d2559 ?
	       _theResult___snd_fst_exp__h81822 :
	       11'd2047 ;
  assign _theResult___snd_fst_exp__h97196 =
	     _64_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d2888 ?
	       _theResult___fst_exp__h96434 :
	       _theResult___fst_exp__h97193 ;
  assign _theResult___snd_fst_exp__h97199 =
	     _64_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d2885 ?
	       11'd0 :
	       _theResult___snd_fst_exp__h97196 ;
  assign _theResult___snd_fst_exp__h97202 =
	     _64_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d2883 ?
	       _theResult___snd_fst_exp__h97199 :
	       11'd2047 ;
  assign _theResult___snd_fst_sfd__h109720 =
	     _64_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d3071 ?
	       _theResult___fst_sfd__h108959 :
	       _theResult___fst_sfd__h109717 ;
  assign _theResult___snd_fst_sfd__h117207 =
	     (value__h113092[51:29] == 23'd0) ?
	       23'd2097152 :
	       value__h113092[51:29] ;
  assign _theResult___snd_fst_sfd__h145866 =
	     _3074_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_ETC___d3422 ?
	       _theResult___fst_sfd__h136018 :
	       _theResult___fst_sfd__h145863 ;
  assign _theResult___snd_fst_sfd__h16088 =
	     _64_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d450 ?
	       _theResult___fst_sfd__h15529 :
	       _theResult___fst_sfd__h16085 ;
  assign _theResult___snd_fst_sfd__h166261 =
	     SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_3_B_ETC___d3853 ?
	       _theResult___fst_sfd__h156359 :
	       _theResult___fst_sfd__h166258 ;
  assign _theResult___snd_fst_sfd__h169840 =
	     (value__h167957 == 23'd0) ?
	       52'h4000000000000 :
	       out___1_sfd__h167954 ;
  assign _theResult___snd_fst_sfd__h191266 =
	     _3970_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_21_ETC___d4543 ?
	       52'd0 :
	       _theResult___fst_sfd__h191263 ;
  assign _theResult___snd_fst_sfd__h212183 =
	     SEXT_IF_IF_requestR_3_BIT_214_4_THEN_requestR__ETC___d4686 ?
	       _theResult___fst_sfd__h202165 :
	       _theResult___fst_sfd__h212180 ;
  assign _theResult___snd_fst_sfd__h28364 =
	     _64_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d972 ?
	       _theResult___fst_sfd__h27806 :
	       _theResult___fst_sfd__h28361 ;
  assign _theResult___snd_fst_sfd__h35538 =
	     _32_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d1327 ?
	       _theResult___fst_sfd__h34979 :
	       _theResult___fst_sfd__h35535 ;
  assign _theResult___snd_fst_sfd__h42452 =
	     _32_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d1580 ?
	       _theResult___fst_sfd__h41894 :
	       _theResult___fst_sfd__h42449 ;
  assign _theResult___snd_fst_sfd__h70875 =
	     _32_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d2347 ?
	       _theResult___fst_sfd__h70113 :
	       _theResult___fst_sfd__h70872 ;
  assign _theResult___snd_fst_sfd__h81820 =
	     _32_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d2561 ?
	       _theResult___fst_sfd__h81059 :
	       _theResult___fst_sfd__h81817 ;
  assign _theResult___snd_fst_sfd__h97197 =
	     _64_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d2888 ?
	       _theResult___fst_sfd__h96435 :
	       _theResult___fst_sfd__h97194 ;
  assign b__h110422 = { value__h82527, 64'd0 } ;
  assign b__h43158 = { value__h43160, 64'd0 } ;
  assign b__h46021 = { value__h43160, 32'd0 } ;
  assign b__h82525 = { value__h82527, 32'd0 } ;
  assign din_inc___2_exp__h109755 = x__h108990[10:0] + 11'd1 ;
  assign din_inc___2_exp__h16127 = x__h15560[7:0] + 8'd1 ;
  assign din_inc___2_exp__h166288 = _theResult___fst_exp__h135390 + 8'd1 ;
  assign din_inc___2_exp__h166312 = _theResult___fst_exp__h145309 + 8'd1 ;
  assign din_inc___2_exp__h166342 = _theResult___fst_exp__h155731 + 8'd1 ;
  assign din_inc___2_exp__h166366 = _theResult___fst_exp__h165679 + 8'd1 ;
  assign din_inc___2_exp__h212214 = _theResult___fst_exp__h190506 + 11'd1 ;
  assign din_inc___2_exp__h212244 = _theResult___fst_exp__h201334 + 11'd1 ;
  assign din_inc___2_exp__h212268 = _theResult___fst_exp__h211398 + 11'd1 ;
  assign din_inc___2_exp__h28399 = x__h27837[7:0] + 8'd1 ;
  assign din_inc___2_exp__h35577 = x__h35010[7:0] + 8'd1 ;
  assign din_inc___2_exp__h42487 = x__h41925[7:0] + 8'd1 ;
  assign din_inc___2_exp__h70914 = x__h70144[10:0] + 11'd1 ;
  assign din_inc___2_exp__h81855 = x__h81090[10:0] + 11'd1 ;
  assign din_inc___2_exp__h97236 = x__h96466[10:0] + 11'd1 ;
  assign fcsr__h3933 =
	     { 2'd0,
	       requestR[191:128] != 64'd0 &&
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d684,
	       requestR[191:128] != 64'd0 &&
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d687,
	       requestR[191:128] != 64'd0 &&
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d696 } ;
  assign guard__h108246 =
	     { IF_sfd___37286_BIT_11_THEN_2_ELSE_0__q27[1],
	       { sfd___3__h27286[10:0], 52'd0 } != 63'd0 } ;
  assign guard__h108975 =
	     { IF_sfd___37286_BIT_10_THEN_2_ELSE_0__q28[1],
	       { sfd___3__h27286[9:0], 53'd0 } != 63'd0 } ;
  assign guard__h110355 =
	     { IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d3224[52],
	       { IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d3224[51:0],
		 65'd0 } !=
	       117'd0 } ;
  assign guard__h111133 =
	     { IF_x11322_BIT_53_THEN_2_ELSE_0__q115[1],
	       { x__h111322[52:0], 64'd0 } != 117'd0 } ;
  assign guard__h112440 =
	     { IF_x12661_BIT_53_THEN_2_ELSE_0__q116[1],
	       { x__h112661[52:0], 64'd0 } != 117'd0 } ;
  assign guard__h126038 =
	     { IF_sfdin35384_BIT_33_THEN_2_ELSE_0__q118[1],
	       { sfdin__h135384[32:0], 23'd0 } != 56'd0 } ;
  assign guard__h136028 =
	     { IF_theResult___snd45260_BIT_33_THEN_2_ELSE_0__q120[1],
	       { _theResult___snd__h145260[32:0], 23'd0 } != 56'd0 } ;
  assign guard__h146250 =
	     { IF_sfdin55725_BIT_33_THEN_2_ELSE_0__q123[1],
	       { sfdin__h155725[32:0], 23'd0 } != 56'd0 } ;
  assign guard__h146848 = x__h146948 != 57'd0 ;
  assign guard__h15015 =
	     { IF_sfd___35005_BIT_40_THEN_2_ELSE_0__q9[1],
	       { sfd___3__h15005[39:0], 23'd0 } != 63'd0 } ;
  assign guard__h15545 =
	     { IF_sfd___35005_BIT_39_THEN_2_ELSE_0__q10[1],
	       { sfd___3__h15005[38:0], 24'd0 } != 63'd0 } ;
  assign guard__h156369 =
	     { IF_theResult___snd65625_BIT_33_THEN_2_ELSE_0__q126[1],
	       { _theResult___snd__h165625[32:0], 23'd0 } != 56'd0 } ;
  assign guard__h181312 =
	     { IF_theResult___snd90457_BIT_4_THEN_2_ELSE_0__q152[1],
	       { _theResult___snd__h190457[3:0], 52'd0 } != 56'd0 } ;
  assign guard__h191853 =
	     { IF_sfdin01328_BIT_4_THEN_2_ELSE_0__q155[1],
	       { sfdin__h201328[3:0], 52'd0 } != 56'd0 } ;
  assign guard__h192451 = x__h192551 != 57'd0 ;
  assign guard__h202175 =
	     { IF_theResult___snd11344_BIT_4_THEN_2_ELSE_0__q158[1],
	       { _theResult___snd__h211344[3:0], 52'd0 } != 56'd0 } ;
  assign guard__h27296 =
	     { IF_sfd___37286_BIT_40_THEN_2_ELSE_0__q25[1],
	       { sfd___3__h27286[39:0], 23'd0 } != 63'd0 } ;
  assign guard__h27822 =
	     { IF_sfd___37286_BIT_39_THEN_2_ELSE_0__q26[1],
	       { sfd___3__h27286[38:0], 24'd0 } != 63'd0 } ;
  assign guard__h34468 =
	     { IF_sfd___34458_BIT_8_THEN_2_ELSE_0__q41[1],
	       { sfd___3__h34458[7:0], 23'd0 } != 31'd0 } ;
  assign guard__h34995 =
	     { IF_sfd___34458_BIT_7_THEN_2_ELSE_0__q42[1],
	       { sfd___3__h34458[6:0], 24'd0 } != 31'd0 } ;
  assign guard__h41384 =
	     { IF_sfd___31374_BIT_8_THEN_2_ELSE_0__q55[1],
	       { sfd___3__h41374[7:0], 23'd0 } != 31'd0 } ;
  assign guard__h41910 =
	     { IF_sfd___31374_BIT_7_THEN_2_ELSE_0__q56[1],
	       { sfd___3__h41374[6:0], 24'd0 } != 31'd0 } ;
  assign guard__h43091 =
	     { IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1757[23],
	       { IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1757[22:0],
		 65'd0 } !=
	       88'd0 } ;
  assign guard__h43869 =
	     { IF_x4058_BIT_24_THEN_2_ELSE_0__q66[1],
	       { x__h44058[23:0], 64'd0 } != 88'd0 } ;
  assign guard__h45193 =
	     { IF_x5414_BIT_24_THEN_2_ELSE_0__q67[1],
	       { x__h45414[23:0], 64'd0 } != 88'd0 } ;
  assign guard__h45954 =
	     { IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1908[23],
	       { IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1908[22:0],
		 33'd0 } !=
	       56'd0 } ;
  assign guard__h46508 =
	     { IF_x6697_BIT_24_THEN_2_ELSE_0__q68[1],
	       { x__h46697[23:0], 32'd0 } != 56'd0 } ;
  assign guard__h47594 =
	     { IF_x7815_BIT_24_THEN_2_ELSE_0__q69[1],
	       { x__h47815[23:0], 32'd0 } != 56'd0 } ;
  assign guard__h69399 =
	     { IF_sfd___39389_BIT_2_THEN_2_ELSE_0__q70[1],
	       { sfd___3__h69389[1:0], 52'd0 } != 54'd0 } ;
  assign guard__h70129 =
	     { IF_sfd___39389_BIT_1_THEN_2_ELSE_0__q71[1],
	       { sfd___3__h69389[0], 53'd0 } != 54'd0 } ;
  assign guard__h80346 =
	     { IF_sfd___30336_BIT_2_THEN_2_ELSE_0__q84[1],
	       { sfd___3__h80336[1:0], 52'd0 } != 54'd0 } ;
  assign guard__h81075 =
	     { IF_sfd___30336_BIT_1_THEN_2_ELSE_0__q85[1],
	       { sfd___3__h80336[0], 53'd0 } != 54'd0 } ;
  assign guard__h82458 =
	     { IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2731[52],
	       { IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2731[51:0],
		 33'd0 } !=
	       85'd0 } ;
  assign guard__h83012 =
	     { IF_x3201_BIT_53_THEN_2_ELSE_0__q95[1],
	       { x__h83201[52:0], 32'd0 } != 85'd0 } ;
  assign guard__h84098 =
	     { IF_x4319_BIT_53_THEN_2_ELSE_0__q96[1],
	       { x__h84319[52:0], 32'd0 } != 85'd0 } ;
  assign guard__h95721 =
	     { IF_sfd___35005_BIT_11_THEN_2_ELSE_0__q11[1],
	       { sfd___3__h15005[10:0], 52'd0 } != 63'd0 } ;
  assign guard__h96451 =
	     { IF_sfd___35005_BIT_10_THEN_2_ELSE_0__q12[1],
	       { sfd___3__h15005[9:0], 53'd0 } != 63'd0 } ;
  assign out1___1__h111073 =
	     IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d3224[117:53] +
	     65'd1 ;
  assign out1___1__h43809 =
	     IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1757[88:24] +
	     65'd1 ;
  assign out1___1__h46448 =
	     IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1908[56:24] +
	     33'd1 ;
  assign out1___1__h82952 =
	     IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2731[85:53] +
	     33'd1 ;
  assign out___1_sfd__h167954 = { value__h167957, 29'd0 } ;
  assign out_exp__h108865 =
	     sfd___3__h27286[12] ? _theResult___exp__h108862 : 11'd0 ;
  assign out_exp__h109620 =
	     sfd___3__h27286[11] ?
	       _theResult___exp__h109617 :
	       x__h108990[10:0] ;
  assign out_exp__h135919 =
	     sfdin__h135384[34] ?
	       _theResult___exp__h135916 :
	       _theResult___fst_exp__h135390 ;
  assign out_exp__h145764 =
	     _theResult___snd__h145260[34] ?
	       _theResult___exp__h145761 :
	       _theResult___fst_exp__h145309 ;
  assign out_exp__h15434 =
	     sfd___3__h15005[41] ? _theResult___exp__h15431 : 8'd0 ;
  assign out_exp__h156260 =
	     sfdin__h155725[34] ?
	       _theResult___exp__h156257 :
	       _theResult___fst_exp__h155731 ;
  assign out_exp__h15987 =
	     sfd___3__h15005[40] ? _theResult___exp__h15984 : x__h15560[7:0] ;
  assign out_exp__h166159 =
	     _theResult___snd__h165625[34] ?
	       _theResult___exp__h166156 :
	       _theResult___fst_exp__h165679 ;
  assign out_exp__h191164 =
	     _theResult___snd__h190457[5] ?
	       _theResult___exp__h191161 :
	       _theResult___fst_exp__h190506 ;
  assign out_exp__h202066 =
	     sfdin__h201328[5] ?
	       _theResult___exp__h202063 :
	       _theResult___fst_exp__h201334 ;
  assign out_exp__h212081 =
	     _theResult___snd__h211344[5] ?
	       _theResult___exp__h212078 :
	       _theResult___fst_exp__h211398 ;
  assign out_exp__h27712 =
	     sfd___3__h27286[41] ? _theResult___exp__h27709 : 8'd0 ;
  assign out_exp__h28264 =
	     sfd___3__h27286[40] ? _theResult___exp__h28261 : x__h27837[7:0] ;
  assign out_exp__h34884 =
	     sfd___3__h34458[9] ? _theResult___exp__h34881 : 8'd0 ;
  assign out_exp__h35437 =
	     sfd___3__h34458[8] ? _theResult___exp__h35434 : x__h35010[7:0] ;
  assign out_exp__h41800 =
	     sfd___3__h41374[9] ? _theResult___exp__h41797 : 8'd0 ;
  assign out_exp__h42352 =
	     sfd___3__h41374[8] ? _theResult___exp__h42349 : x__h41925[7:0] ;
  assign out_exp__h70018 =
	     sfd___3__h69389[3] ? _theResult___exp__h70015 : 11'd0 ;
  assign out_exp__h70774 =
	     sfd___3__h69389[2] ? _theResult___exp__h70771 : x__h70144[10:0] ;
  assign out_exp__h80965 =
	     sfd___3__h80336[3] ? _theResult___exp__h80962 : 11'd0 ;
  assign out_exp__h81720 =
	     sfd___3__h80336[2] ? _theResult___exp__h81717 : x__h81090[10:0] ;
  assign out_exp__h96340 =
	     sfd___3__h15005[12] ? _theResult___exp__h96337 : 11'd0 ;
  assign out_exp__h97096 =
	     sfd___3__h15005[11] ?
	       _theResult___exp__h97093 :
	       x__h96466[10:0] ;
  assign out_sfd__h108866 =
	     sfd___3__h27286[12] ?
	       _theResult___sfd__h108863 :
	       sfd___3__h27286[63:12] ;
  assign out_sfd__h109621 =
	     sfd___3__h27286[11] ?
	       _theResult___sfd__h109618 :
	       sfd___3__h27286[62:11] ;
  assign out_sfd__h135920 =
	     sfdin__h135384[34] ?
	       _theResult___sfd__h135917 :
	       sfdin__h135384[56:34] ;
  assign out_sfd__h145765 =
	     _theResult___snd__h145260[34] ?
	       _theResult___sfd__h145762 :
	       _theResult___snd__h145260[56:34] ;
  assign out_sfd__h15435 =
	     sfd___3__h15005[41] ?
	       _theResult___sfd__h15432 :
	       sfd___3__h15005[63:41] ;
  assign out_sfd__h156261 =
	     sfdin__h155725[34] ?
	       _theResult___sfd__h156258 :
	       sfdin__h155725[56:34] ;
  assign out_sfd__h15988 =
	     sfd___3__h15005[40] ?
	       _theResult___sfd__h15985 :
	       sfd___3__h15005[62:40] ;
  assign out_sfd__h166160 =
	     _theResult___snd__h165625[34] ?
	       _theResult___sfd__h166157 :
	       _theResult___snd__h165625[56:34] ;
  assign out_sfd__h191165 =
	     _theResult___snd__h190457[5] ?
	       _theResult___sfd__h191162 :
	       _theResult___snd__h190457[56:5] ;
  assign out_sfd__h202067 =
	     sfdin__h201328[5] ?
	       _theResult___sfd__h202064 :
	       sfdin__h201328[56:5] ;
  assign out_sfd__h212082 =
	     _theResult___snd__h211344[5] ?
	       _theResult___sfd__h212079 :
	       _theResult___snd__h211344[56:5] ;
  assign out_sfd__h27713 =
	     sfd___3__h27286[41] ?
	       _theResult___sfd__h27710 :
	       sfd___3__h27286[63:41] ;
  assign out_sfd__h28265 =
	     sfd___3__h27286[40] ?
	       _theResult___sfd__h28262 :
	       sfd___3__h27286[62:40] ;
  assign out_sfd__h34885 =
	     sfd___3__h34458[9] ?
	       _theResult___sfd__h34882 :
	       sfd___3__h34458[31:9] ;
  assign out_sfd__h35438 =
	     sfd___3__h34458[8] ?
	       _theResult___sfd__h35435 :
	       sfd___3__h34458[30:8] ;
  assign out_sfd__h41801 =
	     sfd___3__h41374[9] ?
	       _theResult___sfd__h41798 :
	       sfd___3__h41374[31:9] ;
  assign out_sfd__h42353 =
	     sfd___3__h41374[8] ?
	       _theResult___sfd__h42350 :
	       sfd___3__h41374[30:8] ;
  assign out_sfd__h70019 =
	     sfd___3__h69389[3] ?
	       _theResult___sfd__h70016 :
	       sfd___3__h69389[54:3] ;
  assign out_sfd__h70775 =
	     sfd___3__h69389[2] ?
	       _theResult___sfd__h70772 :
	       sfd___3__h69389[53:2] ;
  assign out_sfd__h80966 =
	     sfd___3__h80336[3] ?
	       _theResult___sfd__h80963 :
	       sfd___3__h80336[54:3] ;
  assign out_sfd__h81721 =
	     sfd___3__h80336[2] ?
	       _theResult___sfd__h81718 :
	       sfd___3__h80336[53:2] ;
  assign out_sfd__h96341 =
	     sfd___3__h15005[12] ?
	       _theResult___sfd__h96338 :
	       sfd___3__h15005[63:12] ;
  assign out_sfd__h97097 =
	     sfd___3__h15005[11] ?
	       _theResult___sfd__h97094 :
	       sfd___3__h15005[62:11] ;
  assign requestR_BITS_127_TO_64__q3 = requestR[127:64] ;
  assign requestR_BITS_191_TO_128_BITS_31_TO_0__q2 =
	     requestR_BITS_191_TO_128__q1[31:0] ;
  assign requestR_BITS_191_TO_128__q1 = requestR[191:128] ;
  assign requestR_BITS_206_TO_200__q177 = requestR[206:200] ;
  assign requestR_BITS_63_TO_0__q8 = requestR[63:0] ;
  assign res___1__h229866 =
	     (requestR_BITS_191_TO_128__q1[62:52] == 11'd2047 &&
	      requestR_BITS_191_TO_128__q1[51]) ?
	       64'd512 :
	       64'd256 ;
  assign res___1__h230304 =
	     requestR_BITS_191_TO_128__q1[63] ? 64'd1 : 64'd128 ;
  assign res___1__h230314 =
	     requestR_BITS_191_TO_128__q1[63] ? 64'd8 : 64'd16 ;
  assign res___1__h230333 =
	     requestR_BITS_191_TO_128__q1[63] ? 64'd4 : 64'd32 ;
  assign res___1__h57534 =
	     (sV1_exp__h1472 == 8'd255 && sV1_sfd__h1473[22]) ?
	       64'd512 :
	       64'd256 ;
  assign res___1__h57770 =
	     (requestR_BITS_191_TO_128__q1[63:32] == 32'hFFFFFFFF &&
	      requestR_BITS_191_TO_128__q1[31]) ?
	       64'd1 :
	       64'd128 ;
  assign res___1__h57780 =
	     (requestR_BITS_191_TO_128__q1[63:32] == 32'hFFFFFFFF &&
	      requestR_BITS_191_TO_128__q1[31]) ?
	       64'd8 :
	       64'd16 ;
  assign res___1__h57799 =
	     (requestR_BITS_191_TO_128__q1[63:32] == 32'hFFFFFFFF &&
	      requestR_BITS_191_TO_128__q1[31]) ?
	       64'd4 :
	       64'd32 ;
  assign res__h166745 = { 32'hFFFFFFFF, x__h166751 } ;
  assign res__h212818 =
	     { IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3__ETC___d5189,
	       x__h167898,
	       IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3__ETC___d5153 } ;
  assign res__h217300 =
	     NOT_IF_requestR_3_BIT_214_4_THEN_requestR_3_BI_ETC___d5330 ?
	       requestR[191:128] :
	       requestR[127:64] ;
  assign res__h221886 =
	     NOT_IF_requestR_3_BIT_214_4_THEN_requestR_3_BI_ETC___d5330 ?
	       requestR[127:64] :
	       requestR[191:128] ;
  assign res__h224628 =
	     ((requestR_BITS_191_TO_128__q1[62:52] != 11'd2047 ||
	       requestR_BITS_191_TO_128__q1[51:0] == 52'd0) &&
	      (requestR_BITS_127_TO_64__q3[62:52] != 11'd2047 ||
	       requestR_BITS_127_TO_64__q3[51:0] == 52'd0) &&
	      IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d5378) ?
	       64'd1 :
	       64'd0 ;
  assign res__h227363 =
	     NOT_IF_requestR_3_BIT_214_4_THEN_requestR_3_BI_ETC___d5330 ?
	       64'd1 :
	       64'd0 ;
  assign res__h229280 =
	     NOT_IF_requestR_3_BIT_214_4_THEN_requestR_3_BI_ETC___d5399 ?
	       64'd1 :
	       64'd0 ;
  assign res__h230349 = requestR_BITS_191_TO_128__q1[63] ? 64'd2 : 64'd64 ;
  assign res__h230541 = { 32'hFFFFFFFF, fpu$server_core_response_get[36:5] } ;
  assign res__h3932 = { 32'hFFFFFFFF, x__h3975 } ;
  assign res__h48859 =
	     { 32'hFFFFFFFF,
	       IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d48 } ;
  assign res__h49096 =
	     { 32'hFFFFFFFF,
	       requestR_BITS_191_TO_128__q1[63:32] == 32'hFFFFFFFF &&
	       requestR_BITS_191_TO_128__q1[31],
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d37 } ;
  assign res__h54627 =
	     NOT_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_ETC___d2172 ?
	       64'd1 :
	       64'd0 ;
  assign res__h56150 =
	     NOT_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_ETC___d2105 ?
	       64'd1 :
	       64'd0 ;
  assign res__h57259 =
	     NOT_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_ETC___d2192 ?
	       64'd1 :
	       64'd0 ;
  assign res__h57815 =
	     (requestR_BITS_191_TO_128__q1[63:32] == 32'hFFFFFFFF &&
	      requestR_BITS_191_TO_128__q1[31]) ?
	       64'd2 :
	       64'd64 ;
  assign result__h146853 =
	     { _0b0_CONCAT_NOT_IF_requestR_3_BIT_214_4_THEN_re_ETC___d3858[56:1],
	       _0b0_CONCAT_NOT_IF_requestR_3_BIT_214_4_THEN_re_ETC___d3858[0] |
	       guard__h146848 } ;
  assign result__h192456 =
	     { _0b0_CONCAT_NOT_IF_IF_requestR_3_BIT_214_4_THEN_ETC___d4691[56:1],
	       _0b0_CONCAT_NOT_IF_IF_requestR_3_BIT_214_4_THEN_ETC___d4691[0] |
	       guard__h192451 } ;
  assign sV1_exp__h1472 =
	     (requestR_BITS_191_TO_128__q1[63:32] == 32'hFFFFFFFF) ?
	       requestR_BITS_191_TO_128__q1[30:23] :
	       8'd255 ;
  assign sV1_sfd__h1473 =
	     (requestR_BITS_191_TO_128__q1[63:32] == 32'hFFFFFFFF) ?
	       requestR_BITS_191_TO_128__q1[22:0] :
	       23'd4194304 ;
  assign sV2_exp__h1597 =
	     (requestR_BITS_127_TO_64__q3[63:32] == 32'hFFFFFFFF) ?
	       requestR_BITS_127_TO_64__q3[30:23] :
	       8'd255 ;
  assign sV2_sfd__h1598 =
	     (requestR_BITS_127_TO_64__q3[63:32] == 32'hFFFFFFFF) ?
	       requestR_BITS_127_TO_64__q3[22:0] :
	       23'd4194304 ;
  assign sfd___3__h15005 =
	     sfd__h3990 <<
	     IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3__ETC___d441 ;
  assign sfd___3__h27286 =
	     requestR[191:128] <<
	     IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d966 ;
  assign sfd___3__h34458 =
	     sfd__h28849 <<
	     IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3__ETC___d1318 ;
  assign sfd___3__h41374 =
	     requestR_BITS_191_TO_128__q1[31:0] <<
	     IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1574 ;
  assign sfd___3__h69389 =
	     sfd__h60177 <<
	     IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3__ETC___d2339 ;
  assign sfd___3__h80336 =
	     sfd__h71373 <<
	     IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2555 ;
  assign sfd__h108263 = { 2'd0, sfd___3__h27286[63:12] } + 54'd1 ;
  assign sfd__h109005 =
	     { 1'b0, x__h108990[10:0] != 11'd0, sfd___3__h27286[62:11] } +
	     54'd1 ;
  assign sfd__h117253 = { value__h82527, 3'd0 } ;
  assign sfd__h135482 =
	     { 1'b0,
	       _theResult___fst_exp__h135390 != 8'd0,
	       sfdin__h135384[56:34] } +
	     25'd1 ;
  assign sfd__h145327 =
	     { 1'b0,
	       _theResult___fst_exp__h145309 != 8'd0,
	       _theResult___snd__h145260[56:34] } +
	     25'd1 ;
  assign sfd__h15032 = { 2'd0, sfd___3__h15005[63:41] } + 25'd1 ;
  assign sfd__h15575 =
	     { 1'b0, x__h15560[7:0] != 8'd0, sfd___3__h15005[62:40] } +
	     25'd1 ;
  assign sfd__h155823 =
	     { 1'b0,
	       _theResult___fst_exp__h155731 != 8'd0,
	       sfdin__h155725[56:34] } +
	     25'd1 ;
  assign sfd__h165698 =
	     { 1'b0,
	       _theResult___fst_exp__h165679 != 8'd0,
	       _theResult___snd__h165625[56:34] } +
	     25'd1 ;
  assign sfd__h190524 =
	     { 1'b0,
	       _theResult___fst_exp__h190506 != 11'd0,
	       _theResult___snd__h190457[56:5] } +
	     54'd1 ;
  assign sfd__h201426 =
	     { 1'b0,
	       _theResult___fst_exp__h201334 != 11'd0,
	       sfdin__h201328[56:5] } +
	     54'd1 ;
  assign sfd__h211417 =
	     { 1'b0,
	       _theResult___fst_exp__h211398 != 11'd0,
	       _theResult___snd__h211344[56:5] } +
	     54'd1 ;
  assign sfd__h27313 = { 2'd0, sfd___3__h27286[63:41] } + 25'd1 ;
  assign sfd__h27852 =
	     { 1'b0, x__h27837[7:0] != 8'd0, sfd___3__h27286[62:40] } +
	     25'd1 ;
  assign sfd__h28849 =
	     requestR_BITS_191_TO_128__q1[31] ?
	       -requestR_BITS_191_TO_128__q1[31:0] :
	       requestR_BITS_191_TO_128__q1[31:0] ;
  assign sfd__h34485 = { 2'd0, sfd___3__h34458[31:9] } + 25'd1 ;
  assign sfd__h35025 =
	     { 1'b0, x__h35010[7:0] != 8'd0, sfd___3__h34458[30:8] } + 25'd1 ;
  assign sfd__h3990 =
	     requestR_BITS_191_TO_128__q1[63] ?
	       -requestR[191:128] :
	       requestR[191:128] ;
  assign sfd__h41401 = { 2'd0, sfd___3__h41374[31:9] } + 25'd1 ;
  assign sfd__h41940 =
	     { 1'b0, x__h41925[7:0] != 8'd0, sfd___3__h41374[30:8] } + 25'd1 ;
  assign sfd__h60177 = { sfd__h28849, 23'd0 } ;
  assign sfd__h69416 = { 2'd0, sfd___3__h69389[54:3] } + 54'd1 ;
  assign sfd__h70159 =
	     { 1'b0, x__h70144[10:0] != 11'd0, sfd___3__h69389[53:2] } +
	     54'd1 ;
  assign sfd__h71373 = { requestR_BITS_191_TO_128__q1[31:0], 23'd0 } ;
  assign sfd__h80363 = { 2'd0, sfd___3__h80336[54:3] } + 54'd1 ;
  assign sfd__h81105 =
	     { 1'b0, x__h81090[10:0] != 11'd0, sfd___3__h80336[53:2] } +
	     54'd1 ;
  assign sfd__h95738 = { 2'd0, sfd___3__h15005[63:12] } + 54'd1 ;
  assign sfd__h96481 =
	     { 1'b0, x__h96466[10:0] != 11'd0, sfd___3__h15005[62:11] } +
	     54'd1 ;
  assign sfdin__h135384 =
	     _theResult____h126028[56] ?
	       _theResult___snd__h135401 :
	       _theResult___snd__h135412 ;
  assign sfdin__h155725 =
	     _theResult____h146240[56] ?
	       _theResult___snd__h155742 :
	       _theResult___snd__h155753 ;
  assign sfdin__h201328 =
	     _theResult____h191843[56] ?
	       _theResult___snd__h201345 :
	       _theResult___snd__h201356 ;
  assign value__h113092 =
	     (requestR_BITS_191_TO_128__q1[62:52] == 11'd2047 &&
	      requestR_BITS_191_TO_128__q1[51:0] != 52'd0 &&
	      !requestR_BITS_191_TO_128__q1[51]) ?
	       _theResult___fst_sfd__h113549 :
	       requestR_BITS_191_TO_128__q1[51:0] ;
  assign value__h167957 =
	     (sV1_exp__h1472 == 8'd255 && sV1_sfd__h1473 != 23'd0 &&
	      !sV1_sfd__h1473[22]) ?
	       _theResult___fst_sfd__h168212 :
	       sV1_sfd__h1473 ;
  assign value__h43160 = { 1'b0, sV1_exp__h1472 != 8'd0, sV1_sfd__h1473 } ;
  assign value__h82527 =
	     { 1'b0,
	       requestR_BITS_191_TO_128__q1[62:52] != 11'd0,
	       requestR_BITS_191_TO_128__q1[51:0] } ;
  assign x__h108990 =
	     _64_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d3068 +
	     12'd1023 ;
  assign x__h109855 =
	     { 2'd0,
	       requestR[191:128] != 64'd0 &&
	       IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d3199,
	       requestR[191:128] != 64'd0 &&
	       IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d3202,
	       requestR[191:128] != 64'd0 &&
	       IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d3211 } ;
  assign x__h110179 =
	     (requestR_BITS_191_TO_128__q1[62:52] == 11'd2047 &&
	      requestR_BITS_191_TO_128__q1[51:0] != 52'd0 ||
	      !requestR_BITS_191_TO_128__q1[63] &&
	      requestR_BITS_191_TO_128__q1[62:52] == 11'd2047 &&
	      requestR_BITS_191_TO_128__q1[51:0] == 52'd0) ?
	       64'h7FFFFFFFFFFFFFFF :
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d3283 ;
  assign x__h111322 =
	     IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d3224 >>
	     NEG_SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d3250 |
	     ~(118'h3FFFFFFFFFFFFFFFFFFFFFFFFFFFFF >>
	       NEG_SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d3250) &
	     {118{IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d3224[117]}} ;
  assign x__h111943 =
	     { requestR_BITS_191_TO_128__q1[62:52] == 11'd2047 &&
	       requestR_BITS_191_TO_128__q1[51:0] != 52'd0 ||
	       requestR_BITS_191_TO_128__q1[62:52] == 11'd2047 &&
	       requestR_BITS_191_TO_128__q1[51:0] == 52'd0 ||
	       NOT_IF_requestR_3_BIT_214_4_THEN_requestR_3_BI_ETC___d3290,
	       3'd0,
	       (requestR_BITS_191_TO_128__q1[62:52] != 11'd2047 ||
		requestR_BITS_191_TO_128__q1[51:0] == 52'd0) &&
	       (requestR_BITS_191_TO_128__q1[62:52] != 11'd2047 ||
		requestR_BITS_191_TO_128__q1[51:0] != 52'd0) &&
	       (requestR_BITS_191_TO_128__q1[62:52] != 11'd0 ||
		requestR_BITS_191_TO_128__q1[51:0] != 52'd0) &&
	       IF_NEG_SEXT_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d3298 } ;
  assign x__h112240 =
	     (requestR_BITS_191_TO_128__q1[62:52] == 11'd2047 &&
	      requestR_BITS_191_TO_128__q1[51:0] != 52'd0 ||
	      !requestR_BITS_191_TO_128__q1[63] &&
	      requestR_BITS_191_TO_128__q1[62:52] == 11'd2047 &&
	      requestR_BITS_191_TO_128__q1[51:0] == 52'd0) ?
	       64'hFFFFFFFFFFFFFFFF :
	       (requestR_BITS_191_TO_128__q1[63] ?
		  64'd0 :
		  ((requestR_BITS_191_TO_128__q1[62:52] == 11'd2047 &&
		    requestR_BITS_191_TO_128__q1[51:0] == 52'd0) ?
		     64'hFFFFFFFFFFFFFFFF :
		     IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d3337)) ;
  assign x__h112661 =
	     { requestR_BITS_191_TO_128__q1[62:52] != 11'd0,
	       requestR_BITS_191_TO_128__q1[51:0],
	       65'd0 } >>
	     NEG_SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d3308 ;
  assign x__h112739 =
	     { requestR_BITS_191_TO_128__q1[63] ?
		 IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d3357 :
		 IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d3346,
	       3'd0,
	       (requestR_BITS_191_TO_128__q1[62:52] != 11'd2047 ||
		requestR_BITS_191_TO_128__q1[51:0] == 52'd0) &&
	       (requestR_BITS_191_TO_128__q1[62:52] != 11'd2047 ||
		requestR_BITS_191_TO_128__q1[51:0] != 52'd0) &&
	       NOT_IF_requestR_3_BIT_214_4_THEN_requestR_3_BI_ETC___d3351 } ;
  assign x__h113022 =
	     (x__h113032 == 8'd255 &&
	      IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d4338[22]) ?
	       64'hFFFFFFFF7FC00000 :
	       res__h166745 ;
  assign x__h113032 =
	     (requestR_BITS_191_TO_128__q1[62:52] == 11'd2047) ?
	       8'd255 :
	       _theResult___fst_exp__h166269 ;
  assign x__h146948 = sfd__h117253 << x__h146981 ;
  assign x__h146981 =
	     12'd57 -
	     _3970_MINUS_SEXT_IF_requestR_3_BIT_214_4_THEN_r_ETC___d3854 ;
  assign x__h15560 =
	     _64_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d444 +
	     9'd127 ;
  assign x__h166751 =
	     { (requestR_BITS_191_TO_128__q1[62:52] == 11'd2047 &&
		requestR_BITS_191_TO_128__q1[51:0] != 52'd0 ||
		(requestR_BITS_191_TO_128__q1[62:52] == 11'd2047 ||
		 requestR_BITS_191_TO_128__q1[62:52] == 11'd0) &&
		requestR_BITS_191_TO_128__q1[51:0] == 52'd0) ?
		 requestR_BITS_191_TO_128__q1[63] :
		 IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d4378,
	       x__h113032,
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d4338 } ;
  assign x__h166866 =
	     { (requestR_BITS_191_TO_128__q1[62:52] == 11'd2047 &&
		requestR_BITS_191_TO_128__q1[51:0] != 52'd0) ?
		 requestR_BITS_191_TO_128__q1[62:52] == 11'd2047 &&
		 requestR_BITS_191_TO_128__q1[51:0] != 52'd0 &&
		 !requestR_BITS_191_TO_128__q1[51] :
		 (requestR_BITS_191_TO_128__q1[62:52] != 11'd2047 ||
		  requestR_BITS_191_TO_128__q1[51:0] != 52'd0) &&
		 (requestR_BITS_191_TO_128__q1[62:52] != 11'd0 ||
		  requestR_BITS_191_TO_128__q1[51:0] != 52'd0) &&
		 IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d4429,
	       (requestR_BITS_191_TO_128__q1[62:52] != 11'd2047 ||
		requestR_BITS_191_TO_128__q1[51:0] == 52'd0) &&
	       (requestR_BITS_191_TO_128__q1[62:52] != 11'd2047 ||
		requestR_BITS_191_TO_128__q1[51:0] != 52'd0) &&
	       (requestR_BITS_191_TO_128__q1[62:52] != 11'd0 ||
		requestR_BITS_191_TO_128__q1[51:0] != 52'd0) &&
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d4440,
	       (requestR_BITS_191_TO_128__q1[62:52] != 11'd2047 ||
		requestR_BITS_191_TO_128__q1[51:0] == 52'd0) &&
	       (requestR_BITS_191_TO_128__q1[62:52] != 11'd2047 ||
		requestR_BITS_191_TO_128__q1[51:0] != 52'd0) &&
	       (requestR_BITS_191_TO_128__q1[62:52] != 11'd0 ||
		requestR_BITS_191_TO_128__q1[51:0] != 52'd0) &&
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d4456,
	       (requestR_BITS_191_TO_128__q1[62:52] != 11'd2047 ||
		requestR_BITS_191_TO_128__q1[51:0] == 52'd0) &&
	       (requestR_BITS_191_TO_128__q1[62:52] != 11'd2047 ||
		requestR_BITS_191_TO_128__q1[51:0] != 52'd0) &&
	       (requestR_BITS_191_TO_128__q1[62:52] != 11'd0 ||
		requestR_BITS_191_TO_128__q1[51:0] != 52'd0) &&
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d4469,
	       (requestR_BITS_191_TO_128__q1[62:52] != 11'd2047 ||
		requestR_BITS_191_TO_128__q1[51:0] == 52'd0) &&
	       (requestR_BITS_191_TO_128__q1[62:52] != 11'd2047 ||
		requestR_BITS_191_TO_128__q1[51:0] != 52'd0) &&
	       (requestR_BITS_191_TO_128__q1[62:52] != 11'd0 ||
		requestR_BITS_191_TO_128__q1[51:0] != 52'd0) &&
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d4482 } ;
  assign x__h16727 =
	     { 33'h1FFFFFFFE,
	       (requestR[191:128] == 64'd0) ?
		 8'd0 :
		 _theResult___snd_fst_exp__h28369,
	       (requestR[191:128] == 64'd0 ||
		NOT_IF_requestR_3_BIT_214_4_THEN_requestR_3_BI_ETC___d1059) ?
		 23'd0 :
		 _theResult___snd_fst_sfd__h28364 } ;
  assign x__h167888 =
	     (x__h167898 == 11'd2047 &&
	      IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3__ETC___d5153[51]) ?
	       64'h7FF8000000000000 :
	       res__h212818 ;
  assign x__h167898 =
	     (sV1_exp__h1472 == 8'd255) ?
	       11'd2047 :
	       _theResult___fst_exp__h212191 ;
  assign x__h192551 = b__h46021 << x__h192584 ;
  assign x__h192584 =
	     12'd57 -
	     _3074_MINUS_SEXT_IF_IF_requestR_3_BIT_214_4_THE_ETC___d4687 ;
  assign x__h212920 =
	     { IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3__ETC___d5227,
	       (sV1_exp__h1472 != 8'd255 || sV1_sfd__h1473 == 23'd0) &&
	       (sV1_exp__h1472 != 8'd255 || sV1_sfd__h1473 != 23'd0) &&
	       (sV1_exp__h1472 != 8'd0 || sV1_sfd__h1473 != 23'd0) &&
	       IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3__ETC___d5234,
	       (sV1_exp__h1472 != 8'd255 || sV1_sfd__h1473 == 23'd0) &&
	       (sV1_exp__h1472 != 8'd255 || sV1_sfd__h1473 != 23'd0) &&
	       (sV1_exp__h1472 != 8'd0 || sV1_sfd__h1473 != 23'd0) &&
	       IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3__ETC___d5248,
	       (sV1_exp__h1472 != 8'd255 || sV1_sfd__h1473 == 23'd0) &&
	       (sV1_exp__h1472 != 8'd255 || sV1_sfd__h1473 != 23'd0) &&
	       (sV1_exp__h1472 != 8'd0 || sV1_sfd__h1473 != 23'd0) &&
	       IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3__ETC___d5260,
	       (sV1_exp__h1472 != 8'd255 || sV1_sfd__h1473 == 23'd0) &&
	       (sV1_exp__h1472 != 8'd255 || sV1_sfd__h1473 != 23'd0) &&
	       (sV1_exp__h1472 != 8'd0 || sV1_sfd__h1473 != 23'd0) &&
	       IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3__ETC___d5272 } ;
  assign x__h213882 =
	     IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d5294 ?
	       64'h7FF8000000000000 :
	       ((requestR_BITS_191_TO_128__q1[62:52] == 11'd2047 &&
		 requestR_BITS_191_TO_128__q1[51:0] != 52'd0 &&
		 !requestR_BITS_191_TO_128__q1[51]) ?
		  requestR[127:64] :
		  ((requestR_BITS_127_TO_64__q3[62:52] == 11'd2047 &&
		    requestR_BITS_127_TO_64__q3[51:0] != 52'd0 &&
		    !requestR_BITS_127_TO_64__q3[51]) ?
		     requestR[191:128] :
		     ((requestR_BITS_191_TO_128__q1[62:52] == 11'd2047 &&
		       requestR_BITS_191_TO_128__q1[51] &&
		       requestR_BITS_127_TO_64__q3[62:52] == 11'd2047 &&
		       requestR_BITS_127_TO_64__q3[51]) ?
			64'h7FF8000000000000 :
			((requestR_BITS_191_TO_128__q1[62:52] == 11'd2047 &&
			  requestR_BITS_191_TO_128__q1[51]) ?
			   requestR[127:64] :
			   IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d5333)))) ;
  assign x__h217430 =
	     { IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d5339,
	       4'd0 } ;
  assign x__h218468 =
	     IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d5294 ?
	       64'h7FF8000000000000 :
	       ((requestR_BITS_191_TO_128__q1[62:52] == 11'd2047 &&
		 requestR_BITS_191_TO_128__q1[51:0] != 52'd0 &&
		 !requestR_BITS_191_TO_128__q1[51]) ?
		  requestR[127:64] :
		  ((requestR_BITS_127_TO_64__q3[62:52] == 11'd2047 &&
		    requestR_BITS_127_TO_64__q3[51:0] != 52'd0 &&
		    !requestR_BITS_127_TO_64__q3[51]) ?
		     requestR[191:128] :
		     ((requestR_BITS_191_TO_128__q1[62:52] == 11'd2047 &&
		       requestR_BITS_191_TO_128__q1[51] &&
		       requestR_BITS_127_TO_64__q3[62:52] == 11'd2047 &&
		       requestR_BITS_127_TO_64__q3[51]) ?
			64'h7FF8000000000000 :
			((requestR_BITS_191_TO_128__q1[62:52] == 11'd2047 &&
			  requestR_BITS_191_TO_128__q1[51]) ?
			   requestR[127:64] :
			   ((requestR_BITS_127_TO_64__q3[62:52] == 11'd2047 &&
			     requestR_BITS_127_TO_64__q3[51]) ?
			      requestR[191:128] :
			      IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d5348))))) ;
  assign x__h222950 =
	     IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d5363 ?
	       64'd0 :
	       res__h224628 ;
  assign x__h225685 =
	     IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d5363 ?
	       64'd0 :
	       res__h227363 ;
  assign x__h227382 =
	     { requestR_BITS_191_TO_128__q1[62:52] == 11'd2047 &&
	       requestR_BITS_191_TO_128__q1[51:0] != 52'd0 ||
	       requestR_BITS_127_TO_64__q3[62:52] == 11'd2047 &&
	       requestR_BITS_127_TO_64__q3[51:0] != 52'd0,
	       4'd0 } ;
  assign x__h227602 =
	     IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d5363 ?
	       64'd0 :
	       res__h229280 ;
  assign x__h229846 =
	     (requestR_BITS_191_TO_128__q1[62:52] == 11'd2047 &&
	      requestR_BITS_191_TO_128__q1[51:0] != 52'd0) ?
	       res___1__h229866 :
	       ((requestR_BITS_191_TO_128__q1[62:52] == 11'd2047 &&
		 requestR_BITS_191_TO_128__q1[51:0] == 52'd0) ?
		  res___1__h230304 :
		  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d5426) ;
  assign x__h230460 =
	     fpu$server_core_response_get[69] ?
	       ((fpu$server_core_response_get[35:28] == 8'd255 &&
		 fpu$server_core_response_get[27:5] != 23'd0) ?
		  64'hFFFFFFFF7FC00000 :
		  res__h230541) :
	       ((fpu$server_core_response_get[67:57] == 11'd2047 &&
		 fpu$server_core_response_get[56:5] != 52'd0) ?
		  64'h7FF8000000000000 :
		  fpu$server_core_response_get[68:5]) ;
  assign x__h27837 =
	     _64_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d969 +
	     9'd127 ;
  assign x__h28503 =
	     { 2'd0,
	       requestR[191:128] != 64'd0 &&
	       IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d1165,
	       requestR[191:128] != 64'd0 &&
	       IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d1168,
	       requestR[191:128] != 64'd0 &&
	       IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d1177 } ;
  assign x__h28828 = { 32'hFFFFFFFF, x__h28834 } ;
  assign x__h28834 =
	     { requestR_BITS_191_TO_128__q1[31:0] != 32'd0 &&
	       (NOT_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_ETC___d1326 ?
		  requestR_BITS_191_TO_128__q1[31] :
		  IF_32_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_2_ETC___d1379),
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1439,
	       (requestR_BITS_191_TO_128__q1[31:0] == 32'd0 ||
		NOT_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_ETC___d1326) ?
		 23'd0 :
		 _theResult___snd_fst_sfd__h35538 } ;
  assign x__h3429 = { 32'hFFFFFFFF, x__h3436 } ;
  assign x__h3436 =
	     { requestR_BITS_127_TO_64__q3[63:32] == 32'hFFFFFFFF &&
	       requestR_BITS_127_TO_64__q3[31],
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d37 } ;
  assign x__h35010 =
	     _32_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d1321 +
	     9'd127 ;
  assign x__h35703 =
	     { 2'd0,
	       requestR_BITS_191_TO_128__q1[31:0] != 32'd0 &&
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1520,
	       requestR_BITS_191_TO_128__q1[31:0] != 32'd0 &&
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1523,
	       requestR_BITS_191_TO_128__q1[31:0] != 32'd0 &&
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1532 } ;
  assign x__h36028 =
	     { 33'h1FFFFFFFE,
	       (requestR_BITS_191_TO_128__q1[31:0] == 32'd0) ?
		 8'd0 :
		 _theResult___snd_fst_exp__h42457,
	       (requestR_BITS_191_TO_128__q1[31:0] == 32'd0 ||
		NOT_IF_requestR_3_BIT_214_4_THEN_requestR_3_BI_ETC___d1666) ?
		 23'd0 :
		 _theResult___snd_fst_sfd__h42452 } ;
  assign x__h3605 = { 32'hFFFFFFFF, x__h3612 } ;
  assign x__h3612 =
	     { requestR_BITS_127_TO_64__q3[63:32] != 32'hFFFFFFFF ||
	       !requestR_BITS_127_TO_64__q3[31],
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d37 } ;
  assign x__h3778 = { 32'hFFFFFFFF, x__h3785 } ;
  assign x__h3785 =
	     { (requestR_BITS_191_TO_128__q1[63:32] == 32'hFFFFFFFF &&
		requestR_BITS_191_TO_128__q1[31]) !=
	       (requestR_BITS_127_TO_64__q3[63:32] == 32'hFFFFFFFF &&
		requestR_BITS_127_TO_64__q3[31]),
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d37 } ;
  assign x__h3975 =
	     { requestR[191:128] != 64'd0 &&
	       (NOT_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_ETC___d449 ?
		  requestR_BITS_191_TO_128__q1[63] :
		  IF_64_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_2_ETC___d511),
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d571,
	       (requestR[191:128] == 64'd0 ||
		NOT_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_ETC___d449) ?
		 23'd0 :
		 _theResult___snd_fst_sfd__h16088 } ;
  assign x__h41925 =
	     _32_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d1577 +
	     9'd127 ;
  assign x__h42591 =
	     { 2'd0,
	       requestR_BITS_191_TO_128__q1[31:0] != 32'd0 &&
	       IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d1709,
	       requestR_BITS_191_TO_128__q1[31:0] != 32'd0 &&
	       IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d1712,
	       requestR_BITS_191_TO_128__q1[31:0] != 32'd0 &&
	       IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d1721 } ;
  assign x__h42915 =
	     (sV1_exp__h1472 == 8'd255 && sV1_sfd__h1473 != 23'd0 ||
	      (requestR_BITS_191_TO_128__q1[63:32] != 32'hFFFFFFFF ||
	       !requestR_BITS_191_TO_128__q1[31]) &&
	      sV1_exp__h1472 == 8'd255 &&
	      sV1_sfd__h1473 == 23'd0) ?
	       64'h7FFFFFFFFFFFFFFF :
	       IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3__ETC___d1816 ;
  assign x__h44058 =
	     IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1757 >>
	     NEG_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d1783 |
	     ~(89'h1FFFFFFFFFFFFFFFFFFFFFF >>
	       NEG_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d1783) &
	     {89{IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1757[88]}} ;
  assign x__h44696 =
	     { sV1_exp__h1472 == 8'd255 && sV1_sfd__h1473 != 23'd0 ||
	       sV1_exp__h1472 == 8'd255 && sV1_sfd__h1473 == 23'd0 ||
	       NOT_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_ETC___d1826,
	       3'd0,
	       (sV1_exp__h1472 != 8'd255 || sV1_sfd__h1473 == 23'd0) &&
	       (sV1_exp__h1472 != 8'd255 || sV1_sfd__h1473 != 23'd0) &&
	       (sV1_exp__h1472 != 8'd0 || sV1_sfd__h1473 != 23'd0) &&
	       IF_NEG_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_re_ETC___d1837 } ;
  assign x__h44993 =
	     (sV1_exp__h1472 == 8'd255 && sV1_sfd__h1473 != 23'd0 ||
	      (requestR_BITS_191_TO_128__q1[63:32] != 32'hFFFFFFFF ||
	       !requestR_BITS_191_TO_128__q1[31]) &&
	      sV1_exp__h1472 == 8'd255 &&
	      sV1_sfd__h1473 == 23'd0) ?
	       64'hFFFFFFFFFFFFFFFF :
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1878 ;
  assign x__h45414 =
	     { sV1_exp__h1472 != 8'd0, sV1_sfd__h1473, 65'd0 } >>
	     NEG_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d1847 ;
  assign x__h45492 =
	     { (requestR_BITS_191_TO_128__q1[63:32] == 32'hFFFFFFFF &&
		requestR_BITS_191_TO_128__q1[31]) ?
		 IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1896 :
		 IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1885,
	       3'd0,
	       (sV1_exp__h1472 != 8'd255 || sV1_sfd__h1473 == 23'd0) &&
	       (sV1_exp__h1472 != 8'd255 || sV1_sfd__h1473 != 23'd0) &&
	       NOT_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_ETC___d1890 } ;
  assign x__h45775 = { {32{x__h45778[31]}}, x__h45778 } ;
  assign x__h45778 =
	     (sV1_exp__h1472 == 8'd255 && sV1_sfd__h1473 != 23'd0 ||
	      (requestR_BITS_191_TO_128__q1[63:32] != 32'hFFFFFFFF ||
	       !requestR_BITS_191_TO_128__q1[31]) &&
	      sV1_exp__h1472 == 8'd255 &&
	      sV1_sfd__h1473 == 23'd0) ?
	       32'h7FFFFFFF :
	       IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3__ETC___d1967 ;
  assign x__h46697 =
	     IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1908 >>
	     NEG_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d1934 |
	     ~(57'h1FFFFFFFFFFFFFF >>
	       NEG_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d1934) &
	     {57{IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1908[56]}} ;
  assign x__h47094 =
	     { sV1_exp__h1472 == 8'd255 && sV1_sfd__h1473 != 23'd0 ||
	       sV1_exp__h1472 == 8'd255 && sV1_sfd__h1473 == 23'd0 ||
	       NOT_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_ETC___d1975,
	       3'd0,
	       (sV1_exp__h1472 != 8'd255 || sV1_sfd__h1473 == 23'd0) &&
	       (sV1_exp__h1472 != 8'd255 || sV1_sfd__h1473 != 23'd0) &&
	       (sV1_exp__h1472 != 8'd0 || sV1_sfd__h1473 != 23'd0) &&
	       IF_NEG_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_re_ETC___d1983 } ;
  assign x__h47391 = { {32{x__h47394[31]}}, x__h47394 } ;
  assign x__h47394 =
	     (sV1_exp__h1472 == 8'd255 && sV1_sfd__h1473 != 23'd0 ||
	      (requestR_BITS_191_TO_128__q1[63:32] != 32'hFFFFFFFF ||
	       !requestR_BITS_191_TO_128__q1[31]) &&
	      sV1_exp__h1472 == 8'd255 &&
	      sV1_sfd__h1473 == 23'd0) ?
	       32'hFFFFFFFF :
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2024 ;
  assign x__h47815 =
	     { sV1_exp__h1472 != 8'd0, sV1_sfd__h1473, 33'd0 } >>
	     NEG_SEXT_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d1993 ;
  assign x__h47893 =
	     { (requestR_BITS_191_TO_128__q1[63:32] == 32'hFFFFFFFF &&
		requestR_BITS_191_TO_128__q1[31]) ?
		 IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2043 :
		 IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2032,
	       3'd0,
	       (sV1_exp__h1472 != 8'd255 || sV1_sfd__h1473 == 23'd0) &&
	       (sV1_exp__h1472 != 8'd255 || sV1_sfd__h1473 != 23'd0) &&
	       NOT_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_ETC___d2037 } ;
  assign x__h48180 =
	     IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2067 ?
	       64'hFFFFFFFF7FC00000 :
	       IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3__ETC___d2113 ;
  assign x__h50220 =
	     { IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2115,
	       4'd0 } ;
  assign x__h50854 =
	     IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2067 ?
	       64'hFFFFFFFF7FC00000 :
	       IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3__ETC___d2130 ;
  assign x__h53419 = { 32'hFFFFFFFF, requestR_BITS_191_TO_128__q1[31:0] } ;
  assign x__h53579 =
	     { {32{requestR_BITS_191_TO_128_BITS_31_TO_0__q2[31]}},
	       requestR_BITS_191_TO_128_BITS_31_TO_0__q2 } ;
  assign x__h53757 =
	     IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2156 ?
	       64'd0 :
	       res__h54627 ;
  assign x__h55280 =
	     IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2156 ?
	       64'd0 :
	       res__h56150 ;
  assign x__h56169 =
	     { sV1_exp__h1472 == 8'd255 && sV1_sfd__h1473 != 23'd0 ||
	       sV2_exp__h1597 == 8'd255 && sV2_sfd__h1598 != 23'd0,
	       4'd0 } ;
  assign x__h56389 =
	     IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2156 ?
	       64'd0 :
	       res__h57259 ;
  assign x__h57514 =
	     (sV1_exp__h1472 == 8'd255 && sV1_sfd__h1473 != 23'd0) ?
	       res___1__h57534 :
	       IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3__ETC___d2207 ;
  assign x__h59668 =
	     { requestR_BITS_127_TO_64__q3[63],
	       requestR_BITS_191_TO_128__q1[62:0] } ;
  assign x__h59829 =
	     { !requestR_BITS_127_TO_64__q3[63],
	       requestR_BITS_191_TO_128__q1[62:0] } ;
  assign x__h59992 =
	     { requestR_BITS_191_TO_128__q1[63] !=
	       requestR_BITS_127_TO_64__q3[63],
	       requestR_BITS_191_TO_128__q1[62:0] } ;
  assign x__h60162 =
	     { requestR_BITS_191_TO_128__q1[31:0] != 32'd0 &&
	       IF_NOT_32_MINUS_0_CONCAT_IF_IF_IF_requestR_3_B_ETC___d2399,
	       (requestR_BITS_191_TO_128__q1[31:0] == 32'd0) ?
		 11'd0 :
		 _theResult___snd_fst_exp__h70880,
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2496 } ;
  assign x__h70144 =
	     _32_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d2342 +
	     12'd1023 ;
  assign x__h71036 =
	     { 2'd0,
	       requestR_BITS_191_TO_128__q1[31:0] != 32'd0 &&
	       (!_32_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d2343 ||
		!_32_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d2345 &&
		!_32_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d2347 &&
		_theResult___fst_exp__h70871 == 11'd2047 &&
		_theResult___fst_sfd__h70872 == 52'd0),
	       requestR_BITS_191_TO_128__q1[31:0] != 32'd0 &&
	       _32_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d2343 &&
	       _32_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d2345,
	       requestR_BITS_191_TO_128__q1[31:0] != 32'd0 &&
	       _32_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d2343 &&
	       !_32_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d2345 &&
	       IF_32_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_2_ETC___d2513 } ;
  assign x__h71361 =
	     { 1'd0,
	       (requestR_BITS_191_TO_128__q1[31:0] == 32'd0) ?
		 11'd0 :
		 _theResult___snd_fst_exp__h81825,
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2680 } ;
  assign x__h81090 =
	     _32_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d2558 +
	     12'd1023 ;
  assign x__h81955 =
	     { 2'd0,
	       requestR_BITS_191_TO_128__q1[31:0] != 32'd0 &&
	       (!_32_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d2559 ||
		!_32_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d2560 &&
		!_32_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d2561 &&
		_theResult___fst_exp__h81816 == 11'd2047 &&
		_theResult___fst_sfd__h81817 == 52'd0),
	       requestR_BITS_191_TO_128__q1[31:0] != 32'd0 &&
	       _32_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d2559 &&
	       _32_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d2560,
	       requestR_BITS_191_TO_128__q1[31:0] != 32'd0 &&
	       _32_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d2559 &&
	       !_32_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214_4_T_ETC___d2560 &&
	       IF_32_MINUS_0_CONCAT_IF_IF_requestR_3_BIT_214__ETC___d2697 } ;
  assign x__h82279 = { {32{x__h82282[31]}}, x__h82282 } ;
  assign x__h82282 =
	     (requestR_BITS_191_TO_128__q1[62:52] == 11'd2047 &&
	      requestR_BITS_191_TO_128__q1[51:0] != 52'd0 ||
	      !requestR_BITS_191_TO_128__q1[63] &&
	      requestR_BITS_191_TO_128__q1[62:52] == 11'd2047 &&
	      requestR_BITS_191_TO_128__q1[51:0] == 52'd0) ?
	       32'h7FFFFFFF :
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2790 ;
  assign x__h83201 =
	     IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2731 >>
	     NEG_SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d2757 |
	     ~(86'h3FFFFFFFFFFFFFFFFFFFFF >>
	       NEG_SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d2757) &
	     {86{IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2731[85]}} ;
  assign x__h83598 =
	     { requestR_BITS_191_TO_128__q1[62:52] == 11'd2047 &&
	       requestR_BITS_191_TO_128__q1[51:0] != 52'd0 ||
	       requestR_BITS_191_TO_128__q1[62:52] == 11'd2047 &&
	       requestR_BITS_191_TO_128__q1[51:0] == 52'd0 ||
	       NOT_IF_requestR_3_BIT_214_4_THEN_requestR_3_BI_ETC___d2801,
	       3'd0,
	       (requestR_BITS_191_TO_128__q1[62:52] != 11'd2047 ||
		requestR_BITS_191_TO_128__q1[51:0] == 52'd0) &&
	       (requestR_BITS_191_TO_128__q1[62:52] != 11'd2047 ||
		requestR_BITS_191_TO_128__q1[51:0] != 52'd0) &&
	       (requestR_BITS_191_TO_128__q1[62:52] != 11'd0 ||
		requestR_BITS_191_TO_128__q1[51:0] != 52'd0) &&
	       IF_NEG_SEXT_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d2812 } ;
  assign x__h83895 = { {32{x__h83898[31]}}, x__h83898 } ;
  assign x__h83898 =
	     (requestR_BITS_191_TO_128__q1[62:52] == 11'd2047 &&
	      requestR_BITS_191_TO_128__q1[51:0] != 52'd0 ||
	      !requestR_BITS_191_TO_128__q1[63] &&
	      requestR_BITS_191_TO_128__q1[62:52] == 11'd2047 &&
	      requestR_BITS_191_TO_128__q1[51:0] == 52'd0) ?
	       32'hFFFFFFFF :
	       (requestR_BITS_191_TO_128__q1[63] ?
		  32'd0 :
		  ((requestR_BITS_191_TO_128__q1[62:52] == 11'd2047 &&
		    requestR_BITS_191_TO_128__q1[51:0] == 52'd0) ?
		     32'hFFFFFFFF :
		     IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2851)) ;
  assign x__h84319 =
	     { requestR_BITS_191_TO_128__q1[62:52] != 11'd0,
	       requestR_BITS_191_TO_128__q1[51:0],
	       33'd0 } >>
	     NEG_SEXT_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d2822 ;
  assign x__h84397 =
	     { requestR_BITS_191_TO_128__q1[63] ?
		 IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d2872 :
		 IF_requestR_3_BIT_214_4_THEN_requestR_3_BITS_1_ETC___d2861,
	       3'd0,
	       (requestR_BITS_191_TO_128__q1[62:52] != 11'd2047 ||
		requestR_BITS_191_TO_128__q1[51:0] == 52'd0) &&
	       (requestR_BITS_191_TO_128__q1[62:52] != 11'd2047 ||
		requestR_BITS_191_TO_128__q1[51:0] != 52'd0) &&
	       NOT_IF_requestR_3_BIT_214_4_THEN_requestR_3_BI_ETC___d2866 } ;
  assign x__h84681 =
	     { requestR[191:128] != 64'd0 &&
	       (NOT_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_ETC___d2887 ?
		  requestR_BITS_191_TO_128__q1[63] :
		  IF_64_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_2_ETC___d2937),
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2996,
	       (requestR[191:128] == 64'd0 ||
		NOT_IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_ETC___d2887) ?
		 52'd0 :
		 _theResult___snd_fst_sfd__h97197 } ;
  assign x__h96466 =
	     _64_MINUS_0_CONCAT_IF_IF_IF_requestR_3_BIT_214__ETC___d2882 +
	     12'd1023 ;
  assign x__h97358 =
	     { 2'd0,
	       requestR[191:128] != 64'd0 &&
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d3045,
	       requestR[191:128] != 64'd0 &&
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d3048,
	       requestR[191:128] != 64'd0 &&
	       IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d3057 } ;
  assign x__h97683 =
	     { 1'd0,
	       (requestR[191:128] == 64'd0) ?
		 11'd0 :
		 _theResult___snd_fst_exp__h109725,
	       (requestR[191:128] == 64'd0 ||
		NOT_IF_requestR_3_BIT_214_4_THEN_requestR_3_BI_ETC___d3156) ?
		 52'd0 :
		 _theResult___snd_fst_sfd__h109720 } ;
  always@(requestR or requestR_BITS_191_TO_128__q1)
  begin
    case (requestR[194:192])
      3'h1: CASE_requestR_BITS_194_TO_192_0x1_254_0x2_IF_r_ETC__q4 = 8'd254;
      3'h2:
	  CASE_requestR_BITS_194_TO_192_0x1_254_0x2_IF_r_ETC__q4 =
	      requestR_BITS_191_TO_128__q1[63] ? 8'd255 : 8'd254;
      3'h3:
	  CASE_requestR_BITS_194_TO_192_0x1_254_0x2_IF_r_ETC__q4 =
	      requestR_BITS_191_TO_128__q1[63] ? 8'd254 : 8'd255;
      default: CASE_requestR_BITS_194_TO_192_0x1_254_0x2_IF_r_ETC__q4 = 8'd0;
    endcase
  end
  always@(requestR or requestR_BITS_191_TO_128__q1)
  begin
    case (requestR[194:192])
      3'h1:
	  CASE_requestR_BITS_194_TO_192_0x1_8388607_0x2__ETC__q5 =
	      23'd8388607;
      3'h2:
	  CASE_requestR_BITS_194_TO_192_0x1_8388607_0x2__ETC__q5 =
	      requestR_BITS_191_TO_128__q1[63] ? 23'd0 : 23'd8388607;
      3'h3:
	  CASE_requestR_BITS_194_TO_192_0x1_8388607_0x2__ETC__q5 =
	      requestR_BITS_191_TO_128__q1[63] ? 23'd8388607 : 23'd0;
      default: CASE_requestR_BITS_194_TO_192_0x1_8388607_0x2__ETC__q5 = 23'd0;
    endcase
  end
  always@(requestR or requestR_BITS_191_TO_128__q1)
  begin
    case (requestR[194:192])
      3'h1: CASE_requestR_BITS_194_TO_192_0x1_2046_0x2_IF__ETC__q6 = 11'd2046;
      3'h2:
	  CASE_requestR_BITS_194_TO_192_0x1_2046_0x2_IF__ETC__q6 =
	      (requestR_BITS_191_TO_128__q1[63:32] == 32'hFFFFFFFF &&
	       requestR_BITS_191_TO_128__q1[31]) ?
		11'd2047 :
		11'd2046;
      3'h3:
	  CASE_requestR_BITS_194_TO_192_0x1_2046_0x2_IF__ETC__q6 =
	      (requestR_BITS_191_TO_128__q1[63:32] == 32'hFFFFFFFF &&
	       requestR_BITS_191_TO_128__q1[31]) ?
		11'd2046 :
		11'd2047;
      default: CASE_requestR_BITS_194_TO_192_0x1_2046_0x2_IF__ETC__q6 = 11'd0;
    endcase
  end
  always@(requestR or requestR_BITS_191_TO_128__q1)
  begin
    case (requestR[194:192])
      3'h1:
	  CASE_requestR_BITS_194_TO_192_0x1_450359962737_ETC__q7 =
	      52'hFFFFFFFFFFFFF;
      3'h2:
	  CASE_requestR_BITS_194_TO_192_0x1_450359962737_ETC__q7 =
	      (requestR_BITS_191_TO_128__q1[63:32] == 32'hFFFFFFFF &&
	       requestR_BITS_191_TO_128__q1[31]) ?
		52'd0 :
		52'hFFFFFFFFFFFFF;
      3'h3:
	  CASE_requestR_BITS_194_TO_192_0x1_450359962737_ETC__q7 =
	      (requestR_BITS_191_TO_128__q1[63:32] == 32'hFFFFFFFF &&
	       requestR_BITS_191_TO_128__q1[31]) ?
		52'hFFFFFFFFFFFFF :
		52'd0;
      default: CASE_requestR_BITS_194_TO_192_0x1_450359962737_ETC__q7 = 52'd0;
    endcase
  end
  always@(requestR)
  begin
    case (requestR[194:192])
      3'h0:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d61 =
	      requestR[194:192];
      3'h1: IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d61 = 3'd4;
      3'h2: IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d61 = 3'd3;
      3'h3: IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d61 = 3'd2;
      3'h4: IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d61 = 3'd1;
      default: IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d61 =
		   3'd0;
    endcase
  end
  always@(guard__h15015 or requestR_BITS_191_TO_128__q1)
  begin
    case (guard__h15015)
      2'b0, 2'b01, 2'b10:
	  CASE_guard5015_0b0_requestR_BITS_191_TO_128_BI_ETC__q13 =
	      requestR_BITS_191_TO_128__q1[63];
      2'd3:
	  CASE_guard5015_0b0_requestR_BITS_191_TO_128_BI_ETC__q13 =
	      guard__h15015 == 2'b11 && requestR_BITS_191_TO_128__q1[63];
    endcase
  end
  always@(requestR or requestR_BITS_191_TO_128__q1 or guard__h15015)
  begin
    case (requestR[194:192])
      3'h2, 3'h3:
	  CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q14 =
	      requestR_BITS_191_TO_128__q1[63];
      3'h4:
	  CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q14 =
	      (guard__h15015 == 2'b0) ?
		requestR_BITS_191_TO_128__q1[63] :
		(guard__h15015 == 2'b01 || guard__h15015 == 2'b10 ||
		 guard__h15015 == 2'b11) &&
		requestR_BITS_191_TO_128__q1[63];
      default: CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q14 =
		   requestR[194:192] == 3'h1 &&
		   requestR_BITS_191_TO_128__q1[63];
    endcase
  end
  always@(guard__h15545 or requestR_BITS_191_TO_128__q1)
  begin
    case (guard__h15545)
      2'b0, 2'b01, 2'b10:
	  CASE_guard5545_0b0_requestR_BITS_191_TO_128_BI_ETC__q15 =
	      requestR_BITS_191_TO_128__q1[63];
      2'd3:
	  CASE_guard5545_0b0_requestR_BITS_191_TO_128_BI_ETC__q15 =
	      guard__h15545 == 2'b11 && requestR_BITS_191_TO_128__q1[63];
    endcase
  end
  always@(requestR or requestR_BITS_191_TO_128__q1 or guard__h15545)
  begin
    case (requestR[194:192])
      3'h2, 3'h3:
	  CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q16 =
	      requestR_BITS_191_TO_128__q1[63];
      3'h4:
	  CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q16 =
	      (guard__h15545 == 2'b0) ?
		requestR_BITS_191_TO_128__q1[63] :
		(guard__h15545 == 2'b01 || guard__h15545 == 2'b10 ||
		 guard__h15545 == 2'b11) &&
		requestR_BITS_191_TO_128__q1[63];
      default: CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q16 =
		   requestR[194:192] == 3'h1 &&
		   requestR_BITS_191_TO_128__q1[63];
    endcase
  end
  always@(guard__h15015 or _theResult___exp__h15431)
  begin
    case (guard__h15015)
      2'b0: CASE_guard5015_0b0_0_0b1_theResult___exp5431_0_ETC__q17 = 8'd0;
      2'b01, 2'b10, 2'b11:
	  CASE_guard5015_0b0_0_0b1_theResult___exp5431_0_ETC__q17 =
	      _theResult___exp__h15431;
    endcase
  end
  always@(requestR or
	  IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d533 or
	  guard__h15015 or
	  requestR_BITS_191_TO_128__q1 or
	  _theResult___exp__h15431 or
	  CASE_guard5015_0b0_0_0b1_theResult___exp5431_0_ETC__q17)
  begin
    case (requestR[194:192])
      3'h2:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d536 =
	      IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d533;
      3'h3:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d536 =
	      (guard__h15015 == 2'b0 || requestR_BITS_191_TO_128__q1[63]) ?
		8'd0 :
		_theResult___exp__h15431;
      3'h4:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d536 =
	      CASE_guard5015_0b0_0_0b1_theResult___exp5431_0_ETC__q17;
      default: IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d536 =
		   8'd0;
    endcase
  end
  always@(guard__h15015 or out_exp__h15434 or _theResult___exp__h15431)
  begin
    case (guard__h15015)
      2'b0, 2'b01:
	  CASE_guard5015_0b0_0_0b1_0_0b10_out_exp5434_0b_ETC__q18 = 8'd0;
      2'b10:
	  CASE_guard5015_0b0_0_0b1_0_0b10_out_exp5434_0b_ETC__q18 =
	      out_exp__h15434;
      2'b11:
	  CASE_guard5015_0b0_0_0b1_0_0b10_out_exp5434_0b_ETC__q18 =
	      _theResult___exp__h15431;
    endcase
  end
  always@(guard__h15545 or x__h15560 or _theResult___exp__h15984)
  begin
    case (guard__h15545)
      2'b0:
	  CASE_guard5545_0b0_x5560_BITS_7_TO_0_0b1_theRe_ETC__q19 =
	      x__h15560[7:0];
      2'b01, 2'b10, 2'b11:
	  CASE_guard5545_0b0_x5560_BITS_7_TO_0_0b1_theRe_ETC__q19 =
	      _theResult___exp__h15984;
    endcase
  end
  always@(requestR or
	  x__h15560 or
	  IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d561 or
	  IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d559 or
	  CASE_guard5545_0b0_x5560_BITS_7_TO_0_0b1_theRe_ETC__q19)
  begin
    case (requestR[194:192])
      3'h1:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d565 =
	      x__h15560[7:0];
      3'h2:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d565 =
	      IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d561;
      3'h3:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d565 =
	      IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d559;
      3'h4:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d565 =
	      CASE_guard5545_0b0_x5560_BITS_7_TO_0_0b1_theRe_ETC__q19;
      default: IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d565 =
		   8'd0;
    endcase
  end
  always@(guard__h15545 or
	  x__h15560 or out_exp__h15987 or _theResult___exp__h15984)
  begin
    case (guard__h15545)
      2'b0, 2'b01:
	  CASE_guard5545_0b0_x5560_BITS_7_TO_0_0b1_x5560_ETC__q20 =
	      x__h15560[7:0];
      2'b10:
	  CASE_guard5545_0b0_x5560_BITS_7_TO_0_0b1_x5560_ETC__q20 =
	      out_exp__h15987;
      2'b11:
	  CASE_guard5545_0b0_x5560_BITS_7_TO_0_0b1_x5560_ETC__q20 =
	      _theResult___exp__h15984;
    endcase
  end
  always@(guard__h15015 or sfd___3__h15005 or _theResult___sfd__h15432)
  begin
    case (guard__h15015)
      2'b0:
	  CASE_guard5015_0b0_sfd___35005_BITS_63_TO_41_0_ETC__q21 =
	      sfd___3__h15005[63:41];
      2'b01, 2'b10, 2'b11:
	  CASE_guard5015_0b0_sfd___35005_BITS_63_TO_41_0_ETC__q21 =
	      _theResult___sfd__h15432;
    endcase
  end
  always@(requestR or
	  sfd___3__h15005 or
	  IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d584 or
	  IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d582 or
	  CASE_guard5015_0b0_sfd___35005_BITS_63_TO_41_0_ETC__q21)
  begin
    case (requestR[194:192])
      3'h1:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d588 =
	      sfd___3__h15005[63:41];
      3'h2:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d588 =
	      IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d584;
      3'h3:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d588 =
	      IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d582;
      3'h4:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d588 =
	      CASE_guard5015_0b0_sfd___35005_BITS_63_TO_41_0_ETC__q21;
      default: IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d588 =
		   23'd0;
    endcase
  end
  always@(guard__h15015 or
	  sfd___3__h15005 or out_sfd__h15435 or _theResult___sfd__h15432)
  begin
    case (guard__h15015)
      2'b0, 2'b01:
	  CASE_guard5015_0b0_sfd___35005_BITS_63_TO_41_0_ETC__q22 =
	      sfd___3__h15005[63:41];
      2'b10:
	  CASE_guard5015_0b0_sfd___35005_BITS_63_TO_41_0_ETC__q22 =
	      out_sfd__h15435;
      2'b11:
	  CASE_guard5015_0b0_sfd___35005_BITS_63_TO_41_0_ETC__q22 =
	      _theResult___sfd__h15432;
    endcase
  end
  always@(guard__h15545 or sfd___3__h15005 or _theResult___sfd__h15985)
  begin
    case (guard__h15545)
      2'b0:
	  CASE_guard5545_0b0_sfd___35005_BITS_62_TO_40_0_ETC__q23 =
	      sfd___3__h15005[62:40];
      2'b01, 2'b10, 2'b11:
	  CASE_guard5545_0b0_sfd___35005_BITS_62_TO_40_0_ETC__q23 =
	      _theResult___sfd__h15985;
    endcase
  end
  always@(requestR or
	  sfd___3__h15005 or
	  IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d602 or
	  IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d600 or
	  CASE_guard5545_0b0_sfd___35005_BITS_62_TO_40_0_ETC__q23)
  begin
    case (requestR[194:192])
      3'h1:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d606 =
	      sfd___3__h15005[62:40];
      3'h2:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d606 =
	      IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d602;
      3'h3:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d606 =
	      IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d600;
      3'h4:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d606 =
	      CASE_guard5545_0b0_sfd___35005_BITS_62_TO_40_0_ETC__q23;
      default: IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d606 =
		   23'd0;
    endcase
  end
  always@(guard__h15545 or
	  sfd___3__h15005 or out_sfd__h15988 or _theResult___sfd__h15985)
  begin
    case (guard__h15545)
      2'b0, 2'b01:
	  CASE_guard5545_0b0_sfd___35005_BITS_62_TO_40_0_ETC__q24 =
	      sfd___3__h15005[62:40];
      2'b10:
	  CASE_guard5545_0b0_sfd___35005_BITS_62_TO_40_0_ETC__q24 =
	      out_sfd__h15988;
      2'b11:
	  CASE_guard5545_0b0_sfd___35005_BITS_62_TO_40_0_ETC__q24 =
	      _theResult___sfd__h15985;
    endcase
  end
  always@(guard__h27296 or out_exp__h27712 or _theResult___exp__h27709)
  begin
    case (guard__h27296)
      2'b0, 2'b01:
	  CASE_guard7296_0b0_0_0b1_0_0b10_out_exp7712_0b_ETC__q29 = 8'd0;
      2'b10:
	  CASE_guard7296_0b0_0_0b1_0_0b10_out_exp7712_0b_ETC__q29 =
	      out_exp__h27712;
      2'b11:
	  CASE_guard7296_0b0_0_0b1_0_0b10_out_exp7712_0b_ETC__q29 =
	      _theResult___exp__h27709;
    endcase
  end
  always@(guard__h27296 or _theResult___exp__h27709)
  begin
    case (guard__h27296)
      2'b0: CASE_guard7296_0b0_0_0b1_theResult___exp7709_0_ETC__q30 = 8'd0;
      2'b01, 2'b10, 2'b11:
	  CASE_guard7296_0b0_0_0b1_theResult___exp7709_0_ETC__q30 =
	      _theResult___exp__h27709;
    endcase
  end
  always@(requestR or
	  guard__h27296 or
	  _theResult___exp__h27709 or
	  CASE_guard7296_0b0_0_0b1_theResult___exp7709_0_ETC__q30)
  begin
    case (requestR[194:192])
      3'h3:
	  CASE_requestR_BITS_194_TO_192_0x3_IF_guard7296_ETC__q31 =
	      (guard__h27296 == 2'b0) ? 8'd0 : _theResult___exp__h27709;
      3'h4:
	  CASE_requestR_BITS_194_TO_192_0x3_IF_guard7296_ETC__q31 =
	      CASE_guard7296_0b0_0_0b1_theResult___exp7709_0_ETC__q30;
      default: CASE_requestR_BITS_194_TO_192_0x3_IF_guard7296_ETC__q31 = 8'd0;
    endcase
  end
  always@(guard__h108246 or out_exp__h108865 or _theResult___exp__h108862)
  begin
    case (guard__h108246)
      2'b0, 2'b01:
	  CASE_guard08246_0b0_0_0b1_0_0b10_out_exp08865__ETC__q32 = 11'd0;
      2'b10:
	  CASE_guard08246_0b0_0_0b1_0_0b10_out_exp08865__ETC__q32 =
	      out_exp__h108865;
      2'b11:
	  CASE_guard08246_0b0_0_0b1_0_0b10_out_exp08865__ETC__q32 =
	      _theResult___exp__h108862;
    endcase
  end
  always@(guard__h108246 or _theResult___exp__h108862)
  begin
    case (guard__h108246)
      2'b0: CASE_guard08246_0b0_0_0b1_theResult___exp08862_ETC__q33 = 11'd0;
      2'b01, 2'b10, 2'b11:
	  CASE_guard08246_0b0_0_0b1_theResult___exp08862_ETC__q33 =
	      _theResult___exp__h108862;
    endcase
  end
  always@(requestR or
	  guard__h108246 or
	  _theResult___exp__h108862 or
	  CASE_guard08246_0b0_0_0b1_theResult___exp08862_ETC__q33)
  begin
    case (requestR[194:192])
      3'h3:
	  CASE_requestR_BITS_194_TO_192_0x3_IF_guard0824_ETC__q34 =
	      (guard__h108246 == 2'b0) ? 11'd0 : _theResult___exp__h108862;
      3'h4:
	  CASE_requestR_BITS_194_TO_192_0x3_IF_guard0824_ETC__q34 =
	      CASE_guard08246_0b0_0_0b1_theResult___exp08862_ETC__q33;
      default: CASE_requestR_BITS_194_TO_192_0x3_IF_guard0824_ETC__q34 =
		   11'd0;
    endcase
  end
  always@(guard__h27822 or x__h27837 or _theResult___exp__h28261)
  begin
    case (guard__h27822)
      2'b0:
	  CASE_guard7822_0b0_x7837_BITS_7_TO_0_0b1_theRe_ETC__q35 =
	      x__h27837[7:0];
      2'b01, 2'b10, 2'b11:
	  CASE_guard7822_0b0_x7837_BITS_7_TO_0_0b1_theRe_ETC__q35 =
	      _theResult___exp__h28261;
    endcase
  end
  always@(requestR or
	  x__h27837 or
	  guard__h27822 or
	  _theResult___exp__h28261 or
	  CASE_guard7822_0b0_x7837_BITS_7_TO_0_0b1_theRe_ETC__q35)
  begin
    case (requestR[194:192])
      3'h1, 3'h2:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1050 =
	      x__h27837[7:0];
      3'h3:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1050 =
	      (guard__h27822 == 2'b0) ?
		x__h27837[7:0] :
		_theResult___exp__h28261;
      3'h4:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1050 =
	      CASE_guard7822_0b0_x7837_BITS_7_TO_0_0b1_theRe_ETC__q35;
      default: IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1050 =
		   8'd0;
    endcase
  end
  always@(guard__h27822 or
	  x__h27837 or out_exp__h28264 or _theResult___exp__h28261)
  begin
    case (guard__h27822)
      2'b0, 2'b01:
	  CASE_guard7822_0b0_x7837_BITS_7_TO_0_0b1_x7837_ETC__q36 =
	      x__h27837[7:0];
      2'b10:
	  CASE_guard7822_0b0_x7837_BITS_7_TO_0_0b1_x7837_ETC__q36 =
	      out_exp__h28264;
      2'b11:
	  CASE_guard7822_0b0_x7837_BITS_7_TO_0_0b1_x7837_ETC__q36 =
	      _theResult___exp__h28261;
    endcase
  end
  always@(guard__h27822 or sfd___3__h27286 or _theResult___sfd__h28262)
  begin
    case (guard__h27822)
      2'b0:
	  CASE_guard7822_0b0_sfd___37286_BITS_62_TO_40_0_ETC__q37 =
	      sfd___3__h27286[62:40];
      2'b01, 2'b10, 2'b11:
	  CASE_guard7822_0b0_sfd___37286_BITS_62_TO_40_0_ETC__q37 =
	      _theResult___sfd__h28262;
    endcase
  end
  always@(requestR or
	  sfd___3__h27286 or
	  guard__h27822 or
	  _theResult___sfd__h28262 or
	  CASE_guard7822_0b0_sfd___37286_BITS_62_TO_40_0_ETC__q37)
  begin
    case (requestR[194:192])
      3'h1, 3'h2:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1088 =
	      sfd___3__h27286[62:40];
      3'h3:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1088 =
	      (guard__h27822 == 2'b0) ?
		sfd___3__h27286[62:40] :
		_theResult___sfd__h28262;
      3'h4:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1088 =
	      CASE_guard7822_0b0_sfd___37286_BITS_62_TO_40_0_ETC__q37;
      default: IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1088 =
		   23'd0;
    endcase
  end
  always@(guard__h27822 or
	  sfd___3__h27286 or out_sfd__h28265 or _theResult___sfd__h28262)
  begin
    case (guard__h27822)
      2'b0, 2'b01:
	  CASE_guard7822_0b0_sfd___37286_BITS_62_TO_40_0_ETC__q38 =
	      sfd___3__h27286[62:40];
      2'b10:
	  CASE_guard7822_0b0_sfd___37286_BITS_62_TO_40_0_ETC__q38 =
	      out_sfd__h28265;
      2'b11:
	  CASE_guard7822_0b0_sfd___37286_BITS_62_TO_40_0_ETC__q38 =
	      _theResult___sfd__h28262;
    endcase
  end
  always@(guard__h27296 or sfd___3__h27286 or _theResult___sfd__h27710)
  begin
    case (guard__h27296)
      2'b0:
	  CASE_guard7296_0b0_sfd___37286_BITS_63_TO_41_0_ETC__q39 =
	      sfd___3__h27286[63:41];
      2'b01, 2'b10, 2'b11:
	  CASE_guard7296_0b0_sfd___37286_BITS_63_TO_41_0_ETC__q39 =
	      _theResult___sfd__h27710;
    endcase
  end
  always@(requestR or
	  sfd___3__h27286 or
	  guard__h27296 or
	  _theResult___sfd__h27710 or
	  CASE_guard7296_0b0_sfd___37286_BITS_63_TO_41_0_ETC__q39)
  begin
    case (requestR[194:192])
      3'h1, 3'h2:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1073 =
	      sfd___3__h27286[63:41];
      3'h3:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1073 =
	      (guard__h27296 == 2'b0) ?
		sfd___3__h27286[63:41] :
		_theResult___sfd__h27710;
      3'h4:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1073 =
	      CASE_guard7296_0b0_sfd___37286_BITS_63_TO_41_0_ETC__q39;
      default: IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1073 =
		   23'd0;
    endcase
  end
  always@(guard__h27296 or
	  sfd___3__h27286 or out_sfd__h27713 or _theResult___sfd__h27710)
  begin
    case (guard__h27296)
      2'b0, 2'b01:
	  CASE_guard7296_0b0_sfd___37286_BITS_63_TO_41_0_ETC__q40 =
	      sfd___3__h27286[63:41];
      2'b10:
	  CASE_guard7296_0b0_sfd___37286_BITS_63_TO_41_0_ETC__q40 =
	      out_sfd__h27713;
      2'b11:
	  CASE_guard7296_0b0_sfd___37286_BITS_63_TO_41_0_ETC__q40 =
	      _theResult___sfd__h27710;
    endcase
  end
  always@(guard__h34468 or _theResult___exp__h34881)
  begin
    case (guard__h34468)
      2'b0: CASE_guard4468_0b0_0_0b1_theResult___exp4881_0_ETC__q43 = 8'd0;
      2'b01, 2'b10, 2'b11:
	  CASE_guard4468_0b0_0_0b1_theResult___exp4881_0_ETC__q43 =
	      _theResult___exp__h34881;
    endcase
  end
  always@(requestR or
	  IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d1401 or
	  guard__h34468 or
	  requestR_BITS_191_TO_128__q1 or
	  _theResult___exp__h34881 or
	  CASE_guard4468_0b0_0_0b1_theResult___exp4881_0_ETC__q43)
  begin
    case (requestR[194:192])
      3'h2:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1404 =
	      IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d1401;
      3'h3:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1404 =
	      (guard__h34468 == 2'b0 || requestR_BITS_191_TO_128__q1[31]) ?
		8'd0 :
		_theResult___exp__h34881;
      3'h4:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1404 =
	      CASE_guard4468_0b0_0_0b1_theResult___exp4881_0_ETC__q43;
      default: IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1404 =
		   8'd0;
    endcase
  end
  always@(guard__h34468 or out_exp__h34884 or _theResult___exp__h34881)
  begin
    case (guard__h34468)
      2'b0, 2'b01:
	  CASE_guard4468_0b0_0_0b1_0_0b10_out_exp4884_0b_ETC__q44 = 8'd0;
      2'b10:
	  CASE_guard4468_0b0_0_0b1_0_0b10_out_exp4884_0b_ETC__q44 =
	      out_exp__h34884;
      2'b11:
	  CASE_guard4468_0b0_0_0b1_0_0b10_out_exp4884_0b_ETC__q44 =
	      _theResult___exp__h34881;
    endcase
  end
  always@(guard__h34468 or requestR_BITS_191_TO_128__q1)
  begin
    case (guard__h34468)
      2'b0, 2'b01, 2'b10:
	  CASE_guard4468_0b0_requestR_BITS_191_TO_128_BI_ETC__q45 =
	      requestR_BITS_191_TO_128__q1[31];
      2'd3:
	  CASE_guard4468_0b0_requestR_BITS_191_TO_128_BI_ETC__q45 =
	      guard__h34468 == 2'b11 && requestR_BITS_191_TO_128__q1[31];
    endcase
  end
  always@(requestR or requestR_BITS_191_TO_128__q1 or guard__h34468)
  begin
    case (requestR[194:192])
      3'h2, 3'h3:
	  CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q46 =
	      requestR_BITS_191_TO_128__q1[31];
      3'h4:
	  CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q46 =
	      (guard__h34468 == 2'b0) ?
		requestR_BITS_191_TO_128__q1[31] :
		(guard__h34468 == 2'b01 || guard__h34468 == 2'b10 ||
		 guard__h34468 == 2'b11) &&
		requestR_BITS_191_TO_128__q1[31];
      default: CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q46 =
		   requestR[194:192] == 3'h1 &&
		   requestR_BITS_191_TO_128__q1[31];
    endcase
  end
  always@(guard__h34995 or requestR_BITS_191_TO_128__q1)
  begin
    case (guard__h34995)
      2'b0, 2'b01, 2'b10:
	  CASE_guard4995_0b0_requestR_BITS_191_TO_128_BI_ETC__q47 =
	      requestR_BITS_191_TO_128__q1[31];
      2'd3:
	  CASE_guard4995_0b0_requestR_BITS_191_TO_128_BI_ETC__q47 =
	      guard__h34995 == 2'b11 && requestR_BITS_191_TO_128__q1[31];
    endcase
  end
  always@(requestR or requestR_BITS_191_TO_128__q1 or guard__h34995)
  begin
    case (requestR[194:192])
      3'h2, 3'h3:
	  CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q48 =
	      requestR_BITS_191_TO_128__q1[31];
      3'h4:
	  CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q48 =
	      (guard__h34995 == 2'b0) ?
		requestR_BITS_191_TO_128__q1[31] :
		(guard__h34995 == 2'b01 || guard__h34995 == 2'b10 ||
		 guard__h34995 == 2'b11) &&
		requestR_BITS_191_TO_128__q1[31];
      default: CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q48 =
		   requestR[194:192] == 3'h1 &&
		   requestR_BITS_191_TO_128__q1[31];
    endcase
  end
  always@(guard__h34995 or x__h35010 or _theResult___exp__h35434)
  begin
    case (guard__h34995)
      2'b0:
	  CASE_guard4995_0b0_x5010_BITS_7_TO_0_0b1_theRe_ETC__q49 =
	      x__h35010[7:0];
      2'b01, 2'b10, 2'b11:
	  CASE_guard4995_0b0_x5010_BITS_7_TO_0_0b1_theRe_ETC__q49 =
	      _theResult___exp__h35434;
    endcase
  end
  always@(requestR or
	  x__h35010 or
	  IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d1429 or
	  IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d1427 or
	  CASE_guard4995_0b0_x5010_BITS_7_TO_0_0b1_theRe_ETC__q49)
  begin
    case (requestR[194:192])
      3'h1:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1433 =
	      x__h35010[7:0];
      3'h2:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1433 =
	      IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d1429;
      3'h3:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1433 =
	      IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d1427;
      3'h4:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1433 =
	      CASE_guard4995_0b0_x5010_BITS_7_TO_0_0b1_theRe_ETC__q49;
      default: IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1433 =
		   8'd0;
    endcase
  end
  always@(guard__h34995 or
	  x__h35010 or out_exp__h35437 or _theResult___exp__h35434)
  begin
    case (guard__h34995)
      2'b0, 2'b01:
	  CASE_guard4995_0b0_x5010_BITS_7_TO_0_0b1_x5010_ETC__q50 =
	      x__h35010[7:0];
      2'b10:
	  CASE_guard4995_0b0_x5010_BITS_7_TO_0_0b1_x5010_ETC__q50 =
	      out_exp__h35437;
      2'b11:
	  CASE_guard4995_0b0_x5010_BITS_7_TO_0_0b1_x5010_ETC__q50 =
	      _theResult___exp__h35434;
    endcase
  end
  always@(guard__h34468 or sfd___3__h34458 or _theResult___sfd__h34882)
  begin
    case (guard__h34468)
      2'b0:
	  CASE_guard4468_0b0_sfd___34458_BITS_31_TO_9_0b_ETC__q51 =
	      sfd___3__h34458[31:9];
      2'b01, 2'b10, 2'b11:
	  CASE_guard4468_0b0_sfd___34458_BITS_31_TO_9_0b_ETC__q51 =
	      _theResult___sfd__h34882;
    endcase
  end
  always@(requestR or
	  sfd___3__h34458 or
	  IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d1452 or
	  IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d1450 or
	  CASE_guard4468_0b0_sfd___34458_BITS_31_TO_9_0b_ETC__q51)
  begin
    case (requestR[194:192])
      3'h1:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1456 =
	      sfd___3__h34458[31:9];
      3'h2:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1456 =
	      IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d1452;
      3'h3:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1456 =
	      IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d1450;
      3'h4:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1456 =
	      CASE_guard4468_0b0_sfd___34458_BITS_31_TO_9_0b_ETC__q51;
      default: IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1456 =
		   23'd0;
    endcase
  end
  always@(guard__h34468 or
	  sfd___3__h34458 or out_sfd__h34885 or _theResult___sfd__h34882)
  begin
    case (guard__h34468)
      2'b0, 2'b01:
	  CASE_guard4468_0b0_sfd___34458_BITS_31_TO_9_0b_ETC__q52 =
	      sfd___3__h34458[31:9];
      2'b10:
	  CASE_guard4468_0b0_sfd___34458_BITS_31_TO_9_0b_ETC__q52 =
	      out_sfd__h34885;
      2'b11:
	  CASE_guard4468_0b0_sfd___34458_BITS_31_TO_9_0b_ETC__q52 =
	      _theResult___sfd__h34882;
    endcase
  end
  always@(guard__h34995 or sfd___3__h34458 or _theResult___sfd__h35435)
  begin
    case (guard__h34995)
      2'b0:
	  CASE_guard4995_0b0_sfd___34458_BITS_30_TO_8_0b_ETC__q53 =
	      sfd___3__h34458[30:8];
      2'b01, 2'b10, 2'b11:
	  CASE_guard4995_0b0_sfd___34458_BITS_30_TO_8_0b_ETC__q53 =
	      _theResult___sfd__h35435;
    endcase
  end
  always@(requestR or
	  sfd___3__h34458 or
	  IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d1470 or
	  IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d1468 or
	  CASE_guard4995_0b0_sfd___34458_BITS_30_TO_8_0b_ETC__q53)
  begin
    case (requestR[194:192])
      3'h1:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1474 =
	      sfd___3__h34458[30:8];
      3'h2:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1474 =
	      IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d1470;
      3'h3:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1474 =
	      IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d1468;
      3'h4:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1474 =
	      CASE_guard4995_0b0_sfd___34458_BITS_30_TO_8_0b_ETC__q53;
      default: IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1474 =
		   23'd0;
    endcase
  end
  always@(guard__h34995 or
	  sfd___3__h34458 or out_sfd__h35438 or _theResult___sfd__h35435)
  begin
    case (guard__h34995)
      2'b0, 2'b01:
	  CASE_guard4995_0b0_sfd___34458_BITS_30_TO_8_0b_ETC__q54 =
	      sfd___3__h34458[30:8];
      2'b10:
	  CASE_guard4995_0b0_sfd___34458_BITS_30_TO_8_0b_ETC__q54 =
	      out_sfd__h35438;
      2'b11:
	  CASE_guard4995_0b0_sfd___34458_BITS_30_TO_8_0b_ETC__q54 =
	      _theResult___sfd__h35435;
    endcase
  end
  always@(guard__h41384 or out_exp__h41800 or _theResult___exp__h41797)
  begin
    case (guard__h41384)
      2'b0, 2'b01:
	  CASE_guard1384_0b0_0_0b1_0_0b10_out_exp1800_0b_ETC__q57 = 8'd0;
      2'b10:
	  CASE_guard1384_0b0_0_0b1_0_0b10_out_exp1800_0b_ETC__q57 =
	      out_exp__h41800;
      2'b11:
	  CASE_guard1384_0b0_0_0b1_0_0b10_out_exp1800_0b_ETC__q57 =
	      _theResult___exp__h41797;
    endcase
  end
  always@(guard__h41384 or _theResult___exp__h41797)
  begin
    case (guard__h41384)
      2'b0: CASE_guard1384_0b0_0_0b1_theResult___exp1797_0_ETC__q58 = 8'd0;
      2'b01, 2'b10, 2'b11:
	  CASE_guard1384_0b0_0_0b1_theResult___exp1797_0_ETC__q58 =
	      _theResult___exp__h41797;
    endcase
  end
  always@(requestR or
	  guard__h41384 or
	  _theResult___exp__h41797 or
	  CASE_guard1384_0b0_0_0b1_theResult___exp1797_0_ETC__q58)
  begin
    case (requestR[194:192])
      3'h3:
	  CASE_requestR_BITS_194_TO_192_0x3_IF_guard1384_ETC__q59 =
	      (guard__h41384 == 2'b0) ? 8'd0 : _theResult___exp__h41797;
      3'h4:
	  CASE_requestR_BITS_194_TO_192_0x3_IF_guard1384_ETC__q59 =
	      CASE_guard1384_0b0_0_0b1_theResult___exp1797_0_ETC__q58;
      default: CASE_requestR_BITS_194_TO_192_0x3_IF_guard1384_ETC__q59 = 8'd0;
    endcase
  end
  always@(guard__h41910 or x__h41925 or _theResult___exp__h42349)
  begin
    case (guard__h41910)
      2'b0:
	  CASE_guard1910_0b0_x1925_BITS_7_TO_0_0b1_theRe_ETC__q60 =
	      x__h41925[7:0];
      2'b01, 2'b10, 2'b11:
	  CASE_guard1910_0b0_x1925_BITS_7_TO_0_0b1_theRe_ETC__q60 =
	      _theResult___exp__h42349;
    endcase
  end
  always@(requestR or
	  x__h41925 or
	  guard__h41910 or
	  _theResult___exp__h42349 or
	  CASE_guard1910_0b0_x1925_BITS_7_TO_0_0b1_theRe_ETC__q60)
  begin
    case (requestR[194:192])
      3'h1, 3'h2:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1657 =
	      x__h41925[7:0];
      3'h3:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1657 =
	      (guard__h41910 == 2'b0) ?
		x__h41925[7:0] :
		_theResult___exp__h42349;
      3'h4:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1657 =
	      CASE_guard1910_0b0_x1925_BITS_7_TO_0_0b1_theRe_ETC__q60;
      default: IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1657 =
		   8'd0;
    endcase
  end
  always@(guard__h41910 or
	  x__h41925 or out_exp__h42352 or _theResult___exp__h42349)
  begin
    case (guard__h41910)
      2'b0, 2'b01:
	  CASE_guard1910_0b0_x1925_BITS_7_TO_0_0b1_x1925_ETC__q61 =
	      x__h41925[7:0];
      2'b10:
	  CASE_guard1910_0b0_x1925_BITS_7_TO_0_0b1_x1925_ETC__q61 =
	      out_exp__h42352;
      2'b11:
	  CASE_guard1910_0b0_x1925_BITS_7_TO_0_0b1_x1925_ETC__q61 =
	      _theResult___exp__h42349;
    endcase
  end
  always@(guard__h41910 or sfd___3__h41374 or _theResult___sfd__h42350)
  begin
    case (guard__h41910)
      2'b0:
	  CASE_guard1910_0b0_sfd___31374_BITS_30_TO_8_0b_ETC__q62 =
	      sfd___3__h41374[30:8];
      2'b01, 2'b10, 2'b11:
	  CASE_guard1910_0b0_sfd___31374_BITS_30_TO_8_0b_ETC__q62 =
	      _theResult___sfd__h42350;
    endcase
  end
  always@(requestR or
	  sfd___3__h41374 or
	  guard__h41910 or
	  _theResult___sfd__h42350 or
	  CASE_guard1910_0b0_sfd___31374_BITS_30_TO_8_0b_ETC__q62)
  begin
    case (requestR[194:192])
      3'h1, 3'h2:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1695 =
	      sfd___3__h41374[30:8];
      3'h3:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1695 =
	      (guard__h41910 == 2'b0) ?
		sfd___3__h41374[30:8] :
		_theResult___sfd__h42350;
      3'h4:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1695 =
	      CASE_guard1910_0b0_sfd___31374_BITS_30_TO_8_0b_ETC__q62;
      default: IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1695 =
		   23'd0;
    endcase
  end
  always@(guard__h41910 or
	  sfd___3__h41374 or out_sfd__h42353 or _theResult___sfd__h42350)
  begin
    case (guard__h41910)
      2'b0, 2'b01:
	  CASE_guard1910_0b0_sfd___31374_BITS_30_TO_8_0b_ETC__q63 =
	      sfd___3__h41374[30:8];
      2'b10:
	  CASE_guard1910_0b0_sfd___31374_BITS_30_TO_8_0b_ETC__q63 =
	      out_sfd__h42353;
      2'b11:
	  CASE_guard1910_0b0_sfd___31374_BITS_30_TO_8_0b_ETC__q63 =
	      _theResult___sfd__h42350;
    endcase
  end
  always@(guard__h41384 or sfd___3__h41374 or _theResult___sfd__h41798)
  begin
    case (guard__h41384)
      2'b0:
	  CASE_guard1384_0b0_sfd___31374_BITS_31_TO_9_0b_ETC__q64 =
	      sfd___3__h41374[31:9];
      2'b01, 2'b10, 2'b11:
	  CASE_guard1384_0b0_sfd___31374_BITS_31_TO_9_0b_ETC__q64 =
	      _theResult___sfd__h41798;
    endcase
  end
  always@(requestR or
	  sfd___3__h41374 or
	  guard__h41384 or
	  _theResult___sfd__h41798 or
	  CASE_guard1384_0b0_sfd___31374_BITS_31_TO_9_0b_ETC__q64)
  begin
    case (requestR[194:192])
      3'h1, 3'h2:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1680 =
	      sfd___3__h41374[31:9];
      3'h3:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1680 =
	      (guard__h41384 == 2'b0) ?
		sfd___3__h41374[31:9] :
		_theResult___sfd__h41798;
      3'h4:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1680 =
	      CASE_guard1384_0b0_sfd___31374_BITS_31_TO_9_0b_ETC__q64;
      default: IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d1680 =
		   23'd0;
    endcase
  end
  always@(guard__h41384 or
	  sfd___3__h41374 or out_sfd__h41801 or _theResult___sfd__h41798)
  begin
    case (guard__h41384)
      2'b0, 2'b01:
	  CASE_guard1384_0b0_sfd___31374_BITS_31_TO_9_0b_ETC__q65 =
	      sfd___3__h41374[31:9];
      2'b10:
	  CASE_guard1384_0b0_sfd___31374_BITS_31_TO_9_0b_ETC__q65 =
	      out_sfd__h41801;
      2'b11:
	  CASE_guard1384_0b0_sfd___31374_BITS_31_TO_9_0b_ETC__q65 =
	      _theResult___sfd__h41798;
    endcase
  end
  always@(guard__h69399 or requestR_BITS_191_TO_128__q1)
  begin
    case (guard__h69399)
      2'b0, 2'b01, 2'b10:
	  CASE_guard9399_0b0_requestR_BITS_191_TO_128_BI_ETC__q72 =
	      requestR_BITS_191_TO_128__q1[31];
      2'd3:
	  CASE_guard9399_0b0_requestR_BITS_191_TO_128_BI_ETC__q72 =
	      guard__h69399 == 2'b11 && requestR_BITS_191_TO_128__q1[31];
    endcase
  end
  always@(requestR or requestR_BITS_191_TO_128__q1 or guard__h69399)
  begin
    case (requestR[194:192])
      3'h2, 3'h3:
	  CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q73 =
	      requestR_BITS_191_TO_128__q1[31];
      3'h4:
	  CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q73 =
	      (guard__h69399 == 2'b0) ?
		requestR_BITS_191_TO_128__q1[31] :
		(guard__h69399 == 2'b01 || guard__h69399 == 2'b10 ||
		 guard__h69399 == 2'b11) &&
		requestR_BITS_191_TO_128__q1[31];
      default: CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q73 =
		   requestR[194:192] == 3'h1 &&
		   requestR_BITS_191_TO_128__q1[31];
    endcase
  end
  always@(guard__h70129 or requestR_BITS_191_TO_128__q1)
  begin
    case (guard__h70129)
      2'b0, 2'b01, 2'b10:
	  CASE_guard0129_0b0_requestR_BITS_191_TO_128_BI_ETC__q74 =
	      requestR_BITS_191_TO_128__q1[31];
      2'd3:
	  CASE_guard0129_0b0_requestR_BITS_191_TO_128_BI_ETC__q74 =
	      guard__h70129 == 2'b11 && requestR_BITS_191_TO_128__q1[31];
    endcase
  end
  always@(requestR or requestR_BITS_191_TO_128__q1 or guard__h70129)
  begin
    case (requestR[194:192])
      3'h2, 3'h3:
	  CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q75 =
	      requestR_BITS_191_TO_128__q1[31];
      3'h4:
	  CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q75 =
	      (guard__h70129 == 2'b0) ?
		requestR_BITS_191_TO_128__q1[31] :
		(guard__h70129 == 2'b01 || guard__h70129 == 2'b10 ||
		 guard__h70129 == 2'b11) &&
		requestR_BITS_191_TO_128__q1[31];
      default: CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q75 =
		   requestR[194:192] == 3'h1 &&
		   requestR_BITS_191_TO_128__q1[31];
    endcase
  end
  always@(guard__h70129 or x__h70144 or _theResult___exp__h70771)
  begin
    case (guard__h70129)
      2'b0:
	  CASE_guard0129_0b0_x0144_BITS_10_TO_0_0b1_theR_ETC__q76 =
	      x__h70144[10:0];
      2'b01, 2'b10, 2'b11:
	  CASE_guard0129_0b0_x0144_BITS_10_TO_0_0b1_theR_ETC__q76 =
	      _theResult___exp__h70771;
    endcase
  end
  always@(requestR or
	  x__h70144 or
	  IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d2447 or
	  IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d2445 or
	  CASE_guard0129_0b0_x0144_BITS_10_TO_0_0b1_theR_ETC__q76)
  begin
    case (requestR[194:192])
      3'h1:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2451 =
	      x__h70144[10:0];
      3'h2:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2451 =
	      IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d2447;
      3'h3:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2451 =
	      IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d2445;
      3'h4:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2451 =
	      CASE_guard0129_0b0_x0144_BITS_10_TO_0_0b1_theR_ETC__q76;
      default: IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2451 =
		   11'd0;
    endcase
  end
  always@(guard__h70129 or
	  x__h70144 or out_exp__h70774 or _theResult___exp__h70771)
  begin
    case (guard__h70129)
      2'b0, 2'b01:
	  CASE_guard0129_0b0_x0144_BITS_10_TO_0_0b1_x014_ETC__q77 =
	      x__h70144[10:0];
      2'b10:
	  CASE_guard0129_0b0_x0144_BITS_10_TO_0_0b1_x014_ETC__q77 =
	      out_exp__h70774;
      2'b11:
	  CASE_guard0129_0b0_x0144_BITS_10_TO_0_0b1_x014_ETC__q77 =
	      _theResult___exp__h70771;
    endcase
  end
  always@(guard__h70129 or sfd___3__h69389 or _theResult___sfd__h70772)
  begin
    case (guard__h70129)
      2'b0:
	  CASE_guard0129_0b0_sfd___39389_BITS_53_TO_2_0b_ETC__q78 =
	      sfd___3__h69389[53:2];
      2'b01, 2'b10, 2'b11:
	  CASE_guard0129_0b0_sfd___39389_BITS_53_TO_2_0b_ETC__q78 =
	      _theResult___sfd__h70772;
    endcase
  end
  always@(requestR or
	  sfd___3__h69389 or
	  IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d2488 or
	  IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d2486 or
	  CASE_guard0129_0b0_sfd___39389_BITS_53_TO_2_0b_ETC__q78)
  begin
    case (requestR[194:192])
      3'h1:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2492 =
	      sfd___3__h69389[53:2];
      3'h2:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2492 =
	      IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d2488;
      3'h3:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2492 =
	      IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d2486;
      3'h4:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2492 =
	      CASE_guard0129_0b0_sfd___39389_BITS_53_TO_2_0b_ETC__q78;
      default: IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2492 =
		   52'd0;
    endcase
  end
  always@(guard__h70129 or
	  sfd___3__h69389 or out_sfd__h70775 or _theResult___sfd__h70772)
  begin
    case (guard__h70129)
      2'b0, 2'b01:
	  CASE_guard0129_0b0_sfd___39389_BITS_53_TO_2_0b_ETC__q79 =
	      sfd___3__h69389[53:2];
      2'b10:
	  CASE_guard0129_0b0_sfd___39389_BITS_53_TO_2_0b_ETC__q79 =
	      out_sfd__h70775;
      2'b11:
	  CASE_guard0129_0b0_sfd___39389_BITS_53_TO_2_0b_ETC__q79 =
	      _theResult___sfd__h70772;
    endcase
  end
  always@(guard__h69399 or _theResult___exp__h70015)
  begin
    case (guard__h69399)
      2'b0: CASE_guard9399_0b0_0_0b1_theResult___exp0015_0_ETC__q80 = 11'd0;
      2'b01, 2'b10, 2'b11:
	  CASE_guard9399_0b0_0_0b1_theResult___exp0015_0_ETC__q80 =
	      _theResult___exp__h70015;
    endcase
  end
  always@(requestR or
	  IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d2419 or
	  guard__h69399 or
	  requestR_BITS_191_TO_128__q1 or
	  _theResult___exp__h70015 or
	  CASE_guard9399_0b0_0_0b1_theResult___exp0015_0_ETC__q80)
  begin
    case (requestR[194:192])
      3'h2:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2422 =
	      IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d2419;
      3'h3:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2422 =
	      (guard__h69399 == 2'b0 || requestR_BITS_191_TO_128__q1[31]) ?
		11'd0 :
		_theResult___exp__h70015;
      3'h4:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2422 =
	      CASE_guard9399_0b0_0_0b1_theResult___exp0015_0_ETC__q80;
      default: IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2422 =
		   11'd0;
    endcase
  end
  always@(guard__h69399 or out_exp__h70018 or _theResult___exp__h70015)
  begin
    case (guard__h69399)
      2'b0, 2'b01:
	  CASE_guard9399_0b0_0_0b1_0_0b10_out_exp0018_0b_ETC__q81 = 11'd0;
      2'b10:
	  CASE_guard9399_0b0_0_0b1_0_0b10_out_exp0018_0b_ETC__q81 =
	      out_exp__h70018;
      2'b11:
	  CASE_guard9399_0b0_0_0b1_0_0b10_out_exp0018_0b_ETC__q81 =
	      _theResult___exp__h70015;
    endcase
  end
  always@(guard__h69399 or sfd___3__h69389 or _theResult___sfd__h70016)
  begin
    case (guard__h69399)
      2'b0:
	  CASE_guard9399_0b0_sfd___39389_BITS_54_TO_3_0b_ETC__q82 =
	      sfd___3__h69389[54:3];
      2'b01, 2'b10, 2'b11:
	  CASE_guard9399_0b0_sfd___39389_BITS_54_TO_3_0b_ETC__q82 =
	      _theResult___sfd__h70016;
    endcase
  end
  always@(requestR or
	  sfd___3__h69389 or
	  IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d2470 or
	  IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d2468 or
	  CASE_guard9399_0b0_sfd___39389_BITS_54_TO_3_0b_ETC__q82)
  begin
    case (requestR[194:192])
      3'h1:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2474 =
	      sfd___3__h69389[54:3];
      3'h2:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2474 =
	      IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d2470;
      3'h3:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2474 =
	      IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d2468;
      3'h4:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2474 =
	      CASE_guard9399_0b0_sfd___39389_BITS_54_TO_3_0b_ETC__q82;
      default: IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2474 =
		   52'd0;
    endcase
  end
  always@(guard__h69399 or
	  sfd___3__h69389 or out_sfd__h70019 or _theResult___sfd__h70016)
  begin
    case (guard__h69399)
      2'b0, 2'b01:
	  CASE_guard9399_0b0_sfd___39389_BITS_54_TO_3_0b_ETC__q83 =
	      sfd___3__h69389[54:3];
      2'b10:
	  CASE_guard9399_0b0_sfd___39389_BITS_54_TO_3_0b_ETC__q83 =
	      out_sfd__h70019;
      2'b11:
	  CASE_guard9399_0b0_sfd___39389_BITS_54_TO_3_0b_ETC__q83 =
	      _theResult___sfd__h70016;
    endcase
  end
  always@(guard__h80346 or out_exp__h80965 or _theResult___exp__h80962)
  begin
    case (guard__h80346)
      2'b0, 2'b01:
	  CASE_guard0346_0b0_0_0b1_0_0b10_out_exp0965_0b_ETC__q86 = 11'd0;
      2'b10:
	  CASE_guard0346_0b0_0_0b1_0_0b10_out_exp0965_0b_ETC__q86 =
	      out_exp__h80965;
      2'b11:
	  CASE_guard0346_0b0_0_0b1_0_0b10_out_exp0965_0b_ETC__q86 =
	      _theResult___exp__h80962;
    endcase
  end
  always@(guard__h80346 or _theResult___exp__h80962)
  begin
    case (guard__h80346)
      2'b0: CASE_guard0346_0b0_0_0b1_theResult___exp0962_0_ETC__q87 = 11'd0;
      2'b01, 2'b10, 2'b11:
	  CASE_guard0346_0b0_0_0b1_theResult___exp0962_0_ETC__q87 =
	      _theResult___exp__h80962;
    endcase
  end
  always@(requestR or
	  guard__h80346 or
	  _theResult___exp__h80962 or
	  CASE_guard0346_0b0_0_0b1_theResult___exp0962_0_ETC__q87)
  begin
    case (requestR[194:192])
      3'h3:
	  CASE_requestR_BITS_194_TO_192_0x3_IF_guard0346_ETC__q88 =
	      (guard__h80346 == 2'b0) ? 11'd0 : _theResult___exp__h80962;
      3'h4:
	  CASE_requestR_BITS_194_TO_192_0x3_IF_guard0346_ETC__q88 =
	      CASE_guard0346_0b0_0_0b1_theResult___exp0962_0_ETC__q87;
      default: CASE_requestR_BITS_194_TO_192_0x3_IF_guard0346_ETC__q88 =
		   11'd0;
    endcase
  end
  always@(guard__h81075 or x__h81090 or _theResult___exp__h81717)
  begin
    case (guard__h81075)
      2'b0:
	  CASE_guard1075_0b0_x1090_BITS_10_TO_0_0b1_theR_ETC__q89 =
	      x__h81090[10:0];
      2'b01, 2'b10, 2'b11:
	  CASE_guard1075_0b0_x1090_BITS_10_TO_0_0b1_theR_ETC__q89 =
	      _theResult___exp__h81717;
    endcase
  end
  always@(requestR or
	  x__h81090 or
	  guard__h81075 or
	  _theResult___exp__h81717 or
	  CASE_guard1075_0b0_x1090_BITS_10_TO_0_0b1_theR_ETC__q89)
  begin
    case (requestR[194:192])
      3'h1, 3'h2:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2639 =
	      x__h81090[10:0];
      3'h3:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2639 =
	      (guard__h81075 == 2'b0) ?
		x__h81090[10:0] :
		_theResult___exp__h81717;
      3'h4:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2639 =
	      CASE_guard1075_0b0_x1090_BITS_10_TO_0_0b1_theR_ETC__q89;
      default: IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2639 =
		   11'd0;
    endcase
  end
  always@(guard__h81075 or
	  x__h81090 or out_exp__h81720 or _theResult___exp__h81717)
  begin
    case (guard__h81075)
      2'b0, 2'b01:
	  CASE_guard1075_0b0_x1090_BITS_10_TO_0_0b1_x109_ETC__q90 =
	      x__h81090[10:0];
      2'b10:
	  CASE_guard1075_0b0_x1090_BITS_10_TO_0_0b1_x109_ETC__q90 =
	      out_exp__h81720;
      2'b11:
	  CASE_guard1075_0b0_x1090_BITS_10_TO_0_0b1_x109_ETC__q90 =
	      _theResult___exp__h81717;
    endcase
  end
  always@(guard__h81075 or sfd___3__h80336 or _theResult___sfd__h81718)
  begin
    case (guard__h81075)
      2'b0:
	  CASE_guard1075_0b0_sfd___30336_BITS_53_TO_2_0b_ETC__q91 =
	      sfd___3__h80336[53:2];
      2'b01, 2'b10, 2'b11:
	  CASE_guard1075_0b0_sfd___30336_BITS_53_TO_2_0b_ETC__q91 =
	      _theResult___sfd__h81718;
    endcase
  end
  always@(requestR or
	  sfd___3__h80336 or
	  guard__h81075 or
	  _theResult___sfd__h81718 or
	  CASE_guard1075_0b0_sfd___30336_BITS_53_TO_2_0b_ETC__q91)
  begin
    case (requestR[194:192])
      3'h1, 3'h2:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2676 =
	      sfd___3__h80336[53:2];
      3'h3:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2676 =
	      (guard__h81075 == 2'b0) ?
		sfd___3__h80336[53:2] :
		_theResult___sfd__h81718;
      3'h4:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2676 =
	      CASE_guard1075_0b0_sfd___30336_BITS_53_TO_2_0b_ETC__q91;
      default: IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2676 =
		   52'd0;
    endcase
  end
  always@(guard__h81075 or
	  sfd___3__h80336 or out_sfd__h81721 or _theResult___sfd__h81718)
  begin
    case (guard__h81075)
      2'b0, 2'b01:
	  CASE_guard1075_0b0_sfd___30336_BITS_53_TO_2_0b_ETC__q92 =
	      sfd___3__h80336[53:2];
      2'b10:
	  CASE_guard1075_0b0_sfd___30336_BITS_53_TO_2_0b_ETC__q92 =
	      out_sfd__h81721;
      2'b11:
	  CASE_guard1075_0b0_sfd___30336_BITS_53_TO_2_0b_ETC__q92 =
	      _theResult___sfd__h81718;
    endcase
  end
  always@(guard__h80346 or sfd___3__h80336 or _theResult___sfd__h80963)
  begin
    case (guard__h80346)
      2'b0:
	  CASE_guard0346_0b0_sfd___30336_BITS_54_TO_3_0b_ETC__q93 =
	      sfd___3__h80336[54:3];
      2'b01, 2'b10, 2'b11:
	  CASE_guard0346_0b0_sfd___30336_BITS_54_TO_3_0b_ETC__q93 =
	      _theResult___sfd__h80963;
    endcase
  end
  always@(requestR or
	  sfd___3__h80336 or
	  guard__h80346 or
	  _theResult___sfd__h80963 or
	  CASE_guard0346_0b0_sfd___30336_BITS_54_TO_3_0b_ETC__q93)
  begin
    case (requestR[194:192])
      3'h1, 3'h2:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2661 =
	      sfd___3__h80336[54:3];
      3'h3:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2661 =
	      (guard__h80346 == 2'b0) ?
		sfd___3__h80336[54:3] :
		_theResult___sfd__h80963;
      3'h4:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2661 =
	      CASE_guard0346_0b0_sfd___30336_BITS_54_TO_3_0b_ETC__q93;
      default: IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2661 =
		   52'd0;
    endcase
  end
  always@(guard__h80346 or
	  sfd___3__h80336 or out_sfd__h80966 or _theResult___sfd__h80963)
  begin
    case (guard__h80346)
      2'b0, 2'b01:
	  CASE_guard0346_0b0_sfd___30336_BITS_54_TO_3_0b_ETC__q94 =
	      sfd___3__h80336[54:3];
      2'b10:
	  CASE_guard0346_0b0_sfd___30336_BITS_54_TO_3_0b_ETC__q94 =
	      out_sfd__h80966;
      2'b11:
	  CASE_guard0346_0b0_sfd___30336_BITS_54_TO_3_0b_ETC__q94 =
	      _theResult___sfd__h80963;
    endcase
  end
  always@(guard__h95721 or requestR_BITS_191_TO_128__q1)
  begin
    case (guard__h95721)
      2'b0, 2'b01, 2'b10:
	  CASE_guard5721_0b0_requestR_BITS_191_TO_128_BI_ETC__q97 =
	      requestR_BITS_191_TO_128__q1[63];
      2'd3:
	  CASE_guard5721_0b0_requestR_BITS_191_TO_128_BI_ETC__q97 =
	      guard__h95721 == 2'b11 && requestR_BITS_191_TO_128__q1[63];
    endcase
  end
  always@(requestR or requestR_BITS_191_TO_128__q1 or guard__h95721)
  begin
    case (requestR[194:192])
      3'h2, 3'h3:
	  CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q98 =
	      requestR_BITS_191_TO_128__q1[63];
      3'h4:
	  CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q98 =
	      (guard__h95721 == 2'b0) ?
		requestR_BITS_191_TO_128__q1[63] :
		(guard__h95721 == 2'b01 || guard__h95721 == 2'b10 ||
		 guard__h95721 == 2'b11) &&
		requestR_BITS_191_TO_128__q1[63];
      default: CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q98 =
		   requestR[194:192] == 3'h1 &&
		   requestR_BITS_191_TO_128__q1[63];
    endcase
  end
  always@(guard__h96451 or requestR_BITS_191_TO_128__q1)
  begin
    case (guard__h96451)
      2'b0, 2'b01, 2'b10:
	  CASE_guard6451_0b0_requestR_BITS_191_TO_128_BI_ETC__q99 =
	      requestR_BITS_191_TO_128__q1[63];
      2'd3:
	  CASE_guard6451_0b0_requestR_BITS_191_TO_128_BI_ETC__q99 =
	      guard__h96451 == 2'b11 && requestR_BITS_191_TO_128__q1[63];
    endcase
  end
  always@(requestR or requestR_BITS_191_TO_128__q1 or guard__h96451)
  begin
    case (requestR[194:192])
      3'h2, 3'h3:
	  CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q100 =
	      requestR_BITS_191_TO_128__q1[63];
      3'h4:
	  CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q100 =
	      (guard__h96451 == 2'b0) ?
		requestR_BITS_191_TO_128__q1[63] :
		(guard__h96451 == 2'b01 || guard__h96451 == 2'b10 ||
		 guard__h96451 == 2'b11) &&
		requestR_BITS_191_TO_128__q1[63];
      default: CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q100 =
		   requestR[194:192] == 3'h1 &&
		   requestR_BITS_191_TO_128__q1[63];
    endcase
  end
  always@(guard__h96451 or x__h96466 or _theResult___exp__h97093)
  begin
    case (guard__h96451)
      2'b0:
	  CASE_guard6451_0b0_x6466_BITS_10_TO_0_0b1_theR_ETC__q101 =
	      x__h96466[10:0];
      2'b01, 2'b10, 2'b11:
	  CASE_guard6451_0b0_x6466_BITS_10_TO_0_0b1_theR_ETC__q101 =
	      _theResult___exp__h97093;
    endcase
  end
  always@(requestR or
	  x__h96466 or
	  IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d2986 or
	  IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d2984 or
	  CASE_guard6451_0b0_x6466_BITS_10_TO_0_0b1_theR_ETC__q101)
  begin
    case (requestR[194:192])
      3'h1:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2990 =
	      x__h96466[10:0];
      3'h2:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2990 =
	      IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d2986;
      3'h3:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2990 =
	      IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d2984;
      3'h4:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2990 =
	      CASE_guard6451_0b0_x6466_BITS_10_TO_0_0b1_theR_ETC__q101;
      default: IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2990 =
		   11'd0;
    endcase
  end
  always@(guard__h96451 or
	  x__h96466 or out_exp__h97096 or _theResult___exp__h97093)
  begin
    case (guard__h96451)
      2'b0, 2'b01:
	  CASE_guard6451_0b0_x6466_BITS_10_TO_0_0b1_x646_ETC__q102 =
	      x__h96466[10:0];
      2'b10:
	  CASE_guard6451_0b0_x6466_BITS_10_TO_0_0b1_x646_ETC__q102 =
	      out_exp__h97096;
      2'b11:
	  CASE_guard6451_0b0_x6466_BITS_10_TO_0_0b1_x646_ETC__q102 =
	      _theResult___exp__h97093;
    endcase
  end
  always@(guard__h96451 or sfd___3__h15005 or _theResult___sfd__h97094)
  begin
    case (guard__h96451)
      2'b0:
	  CASE_guard6451_0b0_sfd___35005_BITS_62_TO_11_0_ETC__q103 =
	      sfd___3__h15005[62:11];
      2'b01, 2'b10, 2'b11:
	  CASE_guard6451_0b0_sfd___35005_BITS_62_TO_11_0_ETC__q103 =
	      _theResult___sfd__h97094;
    endcase
  end
  always@(requestR or
	  sfd___3__h15005 or
	  IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d3027 or
	  IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d3025 or
	  CASE_guard6451_0b0_sfd___35005_BITS_62_TO_11_0_ETC__q103)
  begin
    case (requestR[194:192])
      3'h1:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d3031 =
	      sfd___3__h15005[62:11];
      3'h2:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d3031 =
	      IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d3027;
      3'h3:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d3031 =
	      IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d3025;
      3'h4:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d3031 =
	      CASE_guard6451_0b0_sfd___35005_BITS_62_TO_11_0_ETC__q103;
      default: IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d3031 =
		   52'd0;
    endcase
  end
  always@(guard__h96451 or
	  sfd___3__h15005 or out_sfd__h97097 or _theResult___sfd__h97094)
  begin
    case (guard__h96451)
      2'b0, 2'b01:
	  CASE_guard6451_0b0_sfd___35005_BITS_62_TO_11_0_ETC__q104 =
	      sfd___3__h15005[62:11];
      2'b10:
	  CASE_guard6451_0b0_sfd___35005_BITS_62_TO_11_0_ETC__q104 =
	      out_sfd__h97097;
      2'b11:
	  CASE_guard6451_0b0_sfd___35005_BITS_62_TO_11_0_ETC__q104 =
	      _theResult___sfd__h97094;
    endcase
  end
  always@(guard__h95721 or _theResult___exp__h96337)
  begin
    case (guard__h95721)
      2'b0: CASE_guard5721_0b0_0_0b1_theResult___exp6337_0_ETC__q105 = 11'd0;
      2'b01, 2'b10, 2'b11:
	  CASE_guard5721_0b0_0_0b1_theResult___exp6337_0_ETC__q105 =
	      _theResult___exp__h96337;
    endcase
  end
  always@(requestR or
	  IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d2958 or
	  guard__h95721 or
	  requestR_BITS_191_TO_128__q1 or
	  _theResult___exp__h96337 or
	  CASE_guard5721_0b0_0_0b1_theResult___exp6337_0_ETC__q105)
  begin
    case (requestR[194:192])
      3'h2:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2961 =
	      IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d2958;
      3'h3:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2961 =
	      (guard__h95721 == 2'b0 || requestR_BITS_191_TO_128__q1[63]) ?
		11'd0 :
		_theResult___exp__h96337;
      3'h4:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2961 =
	      CASE_guard5721_0b0_0_0b1_theResult___exp6337_0_ETC__q105;
      default: IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d2961 =
		   11'd0;
    endcase
  end
  always@(guard__h95721 or out_exp__h96340 or _theResult___exp__h96337)
  begin
    case (guard__h95721)
      2'b0, 2'b01:
	  CASE_guard5721_0b0_0_0b1_0_0b10_out_exp6340_0b_ETC__q106 = 11'd0;
      2'b10:
	  CASE_guard5721_0b0_0_0b1_0_0b10_out_exp6340_0b_ETC__q106 =
	      out_exp__h96340;
      2'b11:
	  CASE_guard5721_0b0_0_0b1_0_0b10_out_exp6340_0b_ETC__q106 =
	      _theResult___exp__h96337;
    endcase
  end
  always@(guard__h95721 or sfd___3__h15005 or _theResult___sfd__h96338)
  begin
    case (guard__h95721)
      2'b0:
	  CASE_guard5721_0b0_sfd___35005_BITS_63_TO_12_0_ETC__q107 =
	      sfd___3__h15005[63:12];
      2'b01, 2'b10, 2'b11:
	  CASE_guard5721_0b0_sfd___35005_BITS_63_TO_12_0_ETC__q107 =
	      _theResult___sfd__h96338;
    endcase
  end
  always@(requestR or
	  sfd___3__h15005 or
	  IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d3009 or
	  IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d3007 or
	  CASE_guard5721_0b0_sfd___35005_BITS_63_TO_12_0_ETC__q107)
  begin
    case (requestR[194:192])
      3'h1:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d3013 =
	      sfd___3__h15005[63:12];
      3'h2:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d3013 =
	      IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d3009;
      3'h3:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d3013 =
	      IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d3007;
      3'h4:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d3013 =
	      CASE_guard5721_0b0_sfd___35005_BITS_63_TO_12_0_ETC__q107;
      default: IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d3013 =
		   52'd0;
    endcase
  end
  always@(guard__h95721 or
	  sfd___3__h15005 or out_sfd__h96341 or _theResult___sfd__h96338)
  begin
    case (guard__h95721)
      2'b0, 2'b01:
	  CASE_guard5721_0b0_sfd___35005_BITS_63_TO_12_0_ETC__q108 =
	      sfd___3__h15005[63:12];
      2'b10:
	  CASE_guard5721_0b0_sfd___35005_BITS_63_TO_12_0_ETC__q108 =
	      out_sfd__h96341;
      2'b11:
	  CASE_guard5721_0b0_sfd___35005_BITS_63_TO_12_0_ETC__q108 =
	      _theResult___sfd__h96338;
    endcase
  end
  always@(guard__h108975 or x__h108990 or _theResult___exp__h109617)
  begin
    case (guard__h108975)
      2'b0:
	  CASE_guard08975_0b0_x08990_BITS_10_TO_0_0b1_th_ETC__q109 =
	      x__h108990[10:0];
      2'b01, 2'b10, 2'b11:
	  CASE_guard08975_0b0_x08990_BITS_10_TO_0_0b1_th_ETC__q109 =
	      _theResult___exp__h109617;
    endcase
  end
  always@(requestR or
	  x__h108990 or
	  guard__h108975 or
	  _theResult___exp__h109617 or
	  CASE_guard08975_0b0_x08990_BITS_10_TO_0_0b1_th_ETC__q109)
  begin
    case (requestR[194:192])
      3'h1, 3'h2:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d3147 =
	      x__h108990[10:0];
      3'h3:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d3147 =
	      (guard__h108975 == 2'b0) ?
		x__h108990[10:0] :
		_theResult___exp__h109617;
      3'h4:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d3147 =
	      CASE_guard08975_0b0_x08990_BITS_10_TO_0_0b1_th_ETC__q109;
      default: IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d3147 =
		   11'd0;
    endcase
  end
  always@(guard__h108975 or
	  x__h108990 or out_exp__h109620 or _theResult___exp__h109617)
  begin
    case (guard__h108975)
      2'b0, 2'b01:
	  CASE_guard08975_0b0_x08990_BITS_10_TO_0_0b1_x0_ETC__q110 =
	      x__h108990[10:0];
      2'b10:
	  CASE_guard08975_0b0_x08990_BITS_10_TO_0_0b1_x0_ETC__q110 =
	      out_exp__h109620;
      2'b11:
	  CASE_guard08975_0b0_x08990_BITS_10_TO_0_0b1_x0_ETC__q110 =
	      _theResult___exp__h109617;
    endcase
  end
  always@(guard__h108975 or sfd___3__h27286 or _theResult___sfd__h109618)
  begin
    case (guard__h108975)
      2'b0:
	  CASE_guard08975_0b0_sfd___37286_BITS_62_TO_11__ETC__q111 =
	      sfd___3__h27286[62:11];
      2'b01, 2'b10, 2'b11:
	  CASE_guard08975_0b0_sfd___37286_BITS_62_TO_11__ETC__q111 =
	      _theResult___sfd__h109618;
    endcase
  end
  always@(requestR or
	  sfd___3__h27286 or
	  guard__h108975 or
	  _theResult___sfd__h109618 or
	  CASE_guard08975_0b0_sfd___37286_BITS_62_TO_11__ETC__q111)
  begin
    case (requestR[194:192])
      3'h1, 3'h2:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d3185 =
	      sfd___3__h27286[62:11];
      3'h3:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d3185 =
	      (guard__h108975 == 2'b0) ?
		sfd___3__h27286[62:11] :
		_theResult___sfd__h109618;
      3'h4:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d3185 =
	      CASE_guard08975_0b0_sfd___37286_BITS_62_TO_11__ETC__q111;
      default: IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d3185 =
		   52'd0;
    endcase
  end
  always@(guard__h108975 or
	  sfd___3__h27286 or out_sfd__h109621 or _theResult___sfd__h109618)
  begin
    case (guard__h108975)
      2'b0, 2'b01:
	  CASE_guard08975_0b0_sfd___37286_BITS_62_TO_11__ETC__q112 =
	      sfd___3__h27286[62:11];
      2'b10:
	  CASE_guard08975_0b0_sfd___37286_BITS_62_TO_11__ETC__q112 =
	      out_sfd__h109621;
      2'b11:
	  CASE_guard08975_0b0_sfd___37286_BITS_62_TO_11__ETC__q112 =
	      _theResult___sfd__h109618;
    endcase
  end
  always@(guard__h108246 or sfd___3__h27286 or _theResult___sfd__h108863)
  begin
    case (guard__h108246)
      2'b0:
	  CASE_guard08246_0b0_sfd___37286_BITS_63_TO_12__ETC__q113 =
	      sfd___3__h27286[63:12];
      2'b01, 2'b10, 2'b11:
	  CASE_guard08246_0b0_sfd___37286_BITS_63_TO_12__ETC__q113 =
	      _theResult___sfd__h108863;
    endcase
  end
  always@(requestR or
	  sfd___3__h27286 or
	  guard__h108246 or
	  _theResult___sfd__h108863 or
	  CASE_guard08246_0b0_sfd___37286_BITS_63_TO_12__ETC__q113)
  begin
    case (requestR[194:192])
      3'h1, 3'h2:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d3170 =
	      sfd___3__h27286[63:12];
      3'h3:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d3170 =
	      (guard__h108246 == 2'b0) ?
		sfd___3__h27286[63:12] :
		_theResult___sfd__h108863;
      3'h4:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d3170 =
	      CASE_guard08246_0b0_sfd___37286_BITS_63_TO_12__ETC__q113;
      default: IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d3170 =
		   52'd0;
    endcase
  end
  always@(guard__h108246 or
	  sfd___3__h27286 or out_sfd__h108866 or _theResult___sfd__h108863)
  begin
    case (guard__h108246)
      2'b0, 2'b01:
	  CASE_guard08246_0b0_sfd___37286_BITS_63_TO_12__ETC__q114 =
	      sfd___3__h27286[63:12];
      2'b10:
	  CASE_guard08246_0b0_sfd___37286_BITS_63_TO_12__ETC__q114 =
	      out_sfd__h108866;
      2'b11:
	  CASE_guard08246_0b0_sfd___37286_BITS_63_TO_12__ETC__q114 =
	      _theResult___sfd__h108863;
    endcase
  end
  always@(guard__h126038 or
	  _theResult___fst_exp__h135390 or _theResult___exp__h135916)
  begin
    case (guard__h126038)
      2'b0:
	  CASE_guard26038_0b0_theResult___fst_exp35390_0_ETC__q127 =
	      _theResult___fst_exp__h135390;
      2'b01, 2'b10, 2'b11:
	  CASE_guard26038_0b0_theResult___fst_exp35390_0_ETC__q127 =
	      _theResult___exp__h135916;
    endcase
  end
  always@(requestR or
	  _theResult___fst_exp__h135390 or
	  IF_IF_IF_IF_0b0_CONCAT_NOT_IF_requestR_3_BIT_2_ETC___d3715 or
	  IF_IF_IF_IF_0b0_CONCAT_NOT_IF_requestR_3_BIT_2_ETC___d3713 or
	  CASE_guard26038_0b0_theResult___fst_exp35390_0_ETC__q127)
  begin
    case (requestR[194:192])
      3'h1:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d3719 =
	      _theResult___fst_exp__h135390;
      3'h2:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d3719 =
	      IF_IF_IF_IF_0b0_CONCAT_NOT_IF_requestR_3_BIT_2_ETC___d3715;
      3'h3:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d3719 =
	      IF_IF_IF_IF_0b0_CONCAT_NOT_IF_requestR_3_BIT_2_ETC___d3713;
      3'h4:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d3719 =
	      CASE_guard26038_0b0_theResult___fst_exp35390_0_ETC__q127;
      default: IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d3719 =
		   8'd0;
    endcase
  end
  always@(guard__h126038 or
	  _theResult___fst_exp__h135390 or
	  out_exp__h135919 or _theResult___exp__h135916)
  begin
    case (guard__h126038)
      2'b0, 2'b01:
	  CASE_guard26038_0b0_theResult___fst_exp35390_0_ETC__q128 =
	      _theResult___fst_exp__h135390;
      2'b10:
	  CASE_guard26038_0b0_theResult___fst_exp35390_0_ETC__q128 =
	      out_exp__h135919;
      2'b11:
	  CASE_guard26038_0b0_theResult___fst_exp35390_0_ETC__q128 =
	      _theResult___exp__h135916;
    endcase
  end
  always@(guard__h136028 or
	  _theResult___fst_exp__h145309 or _theResult___exp__h145761)
  begin
    case (guard__h136028)
      2'b0:
	  CASE_guard36028_0b0_theResult___fst_exp45309_0_ETC__q129 =
	      _theResult___fst_exp__h145309;
      2'b01, 2'b10, 2'b11:
	  CASE_guard36028_0b0_theResult___fst_exp45309_0_ETC__q129 =
	      _theResult___exp__h145761;
    endcase
  end
  always@(requestR or
	  _theResult___fst_exp__h145309 or
	  IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d3832 or
	  IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d3830 or
	  CASE_guard36028_0b0_theResult___fst_exp45309_0_ETC__q129)
  begin
    case (requestR[194:192])
      3'h1:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d3836 =
	      _theResult___fst_exp__h145309;
      3'h2:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d3836 =
	      IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d3832;
      3'h3:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d3836 =
	      IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d3830;
      3'h4:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d3836 =
	      CASE_guard36028_0b0_theResult___fst_exp45309_0_ETC__q129;
      default: IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d3836 =
		   8'd0;
    endcase
  end
  always@(guard__h136028 or
	  _theResult___fst_exp__h145309 or
	  out_exp__h145764 or _theResult___exp__h145761)
  begin
    case (guard__h136028)
      2'b0, 2'b01:
	  CASE_guard36028_0b0_theResult___fst_exp45309_0_ETC__q130 =
	      _theResult___fst_exp__h145309;
      2'b10:
	  CASE_guard36028_0b0_theResult___fst_exp45309_0_ETC__q130 =
	      out_exp__h145764;
      2'b11:
	  CASE_guard36028_0b0_theResult___fst_exp45309_0_ETC__q130 =
	      _theResult___exp__h145761;
    endcase
  end
  always@(guard__h146250 or
	  _theResult___fst_exp__h155731 or _theResult___exp__h156257)
  begin
    case (guard__h146250)
      2'b0:
	  CASE_guard46250_0b0_theResult___fst_exp55731_0_ETC__q131 =
	      _theResult___fst_exp__h155731;
      2'b01, 2'b10, 2'b11:
	  CASE_guard46250_0b0_theResult___fst_exp55731_0_ETC__q131 =
	      _theResult___exp__h156257;
    endcase
  end
  always@(requestR or
	  _theResult___fst_exp__h155731 or
	  IF_IF_IF_IF_3970_MINUS_SEXT_IF_requestR_3_BIT__ETC___d4159 or
	  IF_IF_IF_IF_3970_MINUS_SEXT_IF_requestR_3_BIT__ETC___d4157 or
	  CASE_guard46250_0b0_theResult___fst_exp55731_0_ETC__q131)
  begin
    case (requestR[194:192])
      3'h1:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d4163 =
	      _theResult___fst_exp__h155731;
      3'h2:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d4163 =
	      IF_IF_IF_IF_3970_MINUS_SEXT_IF_requestR_3_BIT__ETC___d4159;
      3'h3:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d4163 =
	      IF_IF_IF_IF_3970_MINUS_SEXT_IF_requestR_3_BIT__ETC___d4157;
      3'h4:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d4163 =
	      CASE_guard46250_0b0_theResult___fst_exp55731_0_ETC__q131;
      default: IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d4163 =
		   8'd0;
    endcase
  end
  always@(guard__h146250 or
	  _theResult___fst_exp__h155731 or
	  out_exp__h156260 or _theResult___exp__h156257)
  begin
    case (guard__h146250)
      2'b0, 2'b01:
	  CASE_guard46250_0b0_theResult___fst_exp55731_0_ETC__q132 =
	      _theResult___fst_exp__h155731;
      2'b10:
	  CASE_guard46250_0b0_theResult___fst_exp55731_0_ETC__q132 =
	      out_exp__h156260;
      2'b11:
	  CASE_guard46250_0b0_theResult___fst_exp55731_0_ETC__q132 =
	      _theResult___exp__h156257;
    endcase
  end
  always@(guard__h156369 or
	  _theResult___fst_exp__h165679 or _theResult___exp__h166156)
  begin
    case (guard__h156369)
      2'b0:
	  CASE_guard56369_0b0_theResult___fst_exp65679_0_ETC__q133 =
	      _theResult___fst_exp__h165679;
      2'b01, 2'b10, 2'b11:
	  CASE_guard56369_0b0_theResult___fst_exp65679_0_ETC__q133 =
	      _theResult___exp__h166156;
    endcase
  end
  always@(requestR or
	  _theResult___fst_exp__h165679 or
	  IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d4228 or
	  IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d4226 or
	  CASE_guard56369_0b0_theResult___fst_exp65679_0_ETC__q133)
  begin
    case (requestR[194:192])
      3'h1:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d4232 =
	      _theResult___fst_exp__h165679;
      3'h2:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d4232 =
	      IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d4228;
      3'h3:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d4232 =
	      IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d4226;
      3'h4:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d4232 =
	      CASE_guard56369_0b0_theResult___fst_exp65679_0_ETC__q133;
      default: IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d4232 =
		   8'd0;
    endcase
  end
  always@(guard__h156369 or
	  _theResult___fst_exp__h165679 or
	  out_exp__h166159 or _theResult___exp__h166156)
  begin
    case (guard__h156369)
      2'b0, 2'b01:
	  CASE_guard56369_0b0_theResult___fst_exp65679_0_ETC__q134 =
	      _theResult___fst_exp__h165679;
      2'b10:
	  CASE_guard56369_0b0_theResult___fst_exp65679_0_ETC__q134 =
	      out_exp__h166159;
      2'b11:
	  CASE_guard56369_0b0_theResult___fst_exp65679_0_ETC__q134 =
	      _theResult___exp__h166156;
    endcase
  end
  always@(guard__h126038 or sfdin__h135384 or _theResult___sfd__h135917)
  begin
    case (guard__h126038)
      2'b0:
	  CASE_guard26038_0b0_sfdin35384_BITS_56_TO_34_0_ETC__q135 =
	      sfdin__h135384[56:34];
      2'b01, 2'b10, 2'b11:
	  CASE_guard26038_0b0_sfdin35384_BITS_56_TO_34_0_ETC__q135 =
	      _theResult___sfd__h135917;
    endcase
  end
  always@(requestR or
	  sfdin__h135384 or
	  IF_IF_IF_IF_0b0_CONCAT_NOT_IF_requestR_3_BIT_2_ETC___d4262 or
	  IF_IF_IF_IF_0b0_CONCAT_NOT_IF_requestR_3_BIT_2_ETC___d4260 or
	  CASE_guard26038_0b0_sfdin35384_BITS_56_TO_34_0_ETC__q135)
  begin
    case (requestR[194:192])
      3'h1:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d4266 =
	      sfdin__h135384[56:34];
      3'h2:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d4266 =
	      IF_IF_IF_IF_0b0_CONCAT_NOT_IF_requestR_3_BIT_2_ETC___d4262;
      3'h3:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d4266 =
	      IF_IF_IF_IF_0b0_CONCAT_NOT_IF_requestR_3_BIT_2_ETC___d4260;
      3'h4:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d4266 =
	      CASE_guard26038_0b0_sfdin35384_BITS_56_TO_34_0_ETC__q135;
      default: IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d4266 =
		   23'd0;
    endcase
  end
  always@(guard__h126038 or
	  sfdin__h135384 or out_sfd__h135920 or _theResult___sfd__h135917)
  begin
    case (guard__h126038)
      2'b0, 2'b01:
	  CASE_guard26038_0b0_sfdin35384_BITS_56_TO_34_0_ETC__q136 =
	      sfdin__h135384[56:34];
      2'b10:
	  CASE_guard26038_0b0_sfdin35384_BITS_56_TO_34_0_ETC__q136 =
	      out_sfd__h135920;
      2'b11:
	  CASE_guard26038_0b0_sfdin35384_BITS_56_TO_34_0_ETC__q136 =
	      _theResult___sfd__h135917;
    endcase
  end
  always@(guard__h136028 or
	  _theResult___snd__h145260 or _theResult___sfd__h145762)
  begin
    case (guard__h136028)
      2'b0:
	  CASE_guard36028_0b0_theResult___snd45260_BITS__ETC__q137 =
	      _theResult___snd__h145260[56:34];
      2'b01, 2'b10, 2'b11:
	  CASE_guard36028_0b0_theResult___snd45260_BITS__ETC__q137 =
	      _theResult___sfd__h145762;
    endcase
  end
  always@(requestR or
	  _theResult___snd__h145260 or
	  IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d4281 or
	  IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d4279 or
	  CASE_guard36028_0b0_theResult___snd45260_BITS__ETC__q137)
  begin
    case (requestR[194:192])
      3'h1:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d4285 =
	      _theResult___snd__h145260[56:34];
      3'h2:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d4285 =
	      IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d4281;
      3'h3:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d4285 =
	      IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d4279;
      3'h4:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d4285 =
	      CASE_guard36028_0b0_theResult___snd45260_BITS__ETC__q137;
      default: IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d4285 =
		   23'd0;
    endcase
  end
  always@(guard__h136028 or
	  _theResult___snd__h145260 or
	  out_sfd__h145765 or _theResult___sfd__h145762)
  begin
    case (guard__h136028)
      2'b0, 2'b01:
	  CASE_guard36028_0b0_theResult___snd45260_BITS__ETC__q138 =
	      _theResult___snd__h145260[56:34];
      2'b10:
	  CASE_guard36028_0b0_theResult___snd45260_BITS__ETC__q138 =
	      out_sfd__h145765;
      2'b11:
	  CASE_guard36028_0b0_theResult___snd45260_BITS__ETC__q138 =
	      _theResult___sfd__h145762;
    endcase
  end
  always@(guard__h146250 or sfdin__h155725 or _theResult___sfd__h156258)
  begin
    case (guard__h146250)
      2'b0:
	  CASE_guard46250_0b0_sfdin55725_BITS_56_TO_34_0_ETC__q139 =
	      sfdin__h155725[56:34];
      2'b01, 2'b10, 2'b11:
	  CASE_guard46250_0b0_sfdin55725_BITS_56_TO_34_0_ETC__q139 =
	      _theResult___sfd__h156258;
    endcase
  end
  always@(requestR or
	  sfdin__h155725 or
	  IF_IF_IF_IF_3970_MINUS_SEXT_IF_requestR_3_BIT__ETC___d4308 or
	  IF_IF_IF_IF_3970_MINUS_SEXT_IF_requestR_3_BIT__ETC___d4306 or
	  CASE_guard46250_0b0_sfdin55725_BITS_56_TO_34_0_ETC__q139)
  begin
    case (requestR[194:192])
      3'h1:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d4312 =
	      sfdin__h155725[56:34];
      3'h2:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d4312 =
	      IF_IF_IF_IF_3970_MINUS_SEXT_IF_requestR_3_BIT__ETC___d4308;
      3'h3:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d4312 =
	      IF_IF_IF_IF_3970_MINUS_SEXT_IF_requestR_3_BIT__ETC___d4306;
      3'h4:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d4312 =
	      CASE_guard46250_0b0_sfdin55725_BITS_56_TO_34_0_ETC__q139;
      default: IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d4312 =
		   23'd0;
    endcase
  end
  always@(guard__h146250 or
	  sfdin__h155725 or out_sfd__h156261 or _theResult___sfd__h156258)
  begin
    case (guard__h146250)
      2'b0, 2'b01:
	  CASE_guard46250_0b0_sfdin55725_BITS_56_TO_34_0_ETC__q140 =
	      sfdin__h155725[56:34];
      2'b10:
	  CASE_guard46250_0b0_sfdin55725_BITS_56_TO_34_0_ETC__q140 =
	      out_sfd__h156261;
      2'b11:
	  CASE_guard46250_0b0_sfdin55725_BITS_56_TO_34_0_ETC__q140 =
	      _theResult___sfd__h156258;
    endcase
  end
  always@(guard__h156369 or
	  _theResult___snd__h165625 or _theResult___sfd__h166157)
  begin
    case (guard__h156369)
      2'b0:
	  CASE_guard56369_0b0_theResult___snd65625_BITS__ETC__q141 =
	      _theResult___snd__h165625[56:34];
      2'b01, 2'b10, 2'b11:
	  CASE_guard56369_0b0_theResult___snd65625_BITS__ETC__q141 =
	      _theResult___sfd__h166157;
    endcase
  end
  always@(requestR or
	  _theResult___snd__h165625 or
	  IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d4327 or
	  IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d4325 or
	  CASE_guard56369_0b0_theResult___snd65625_BITS__ETC__q141)
  begin
    case (requestR[194:192])
      3'h1:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d4331 =
	      _theResult___snd__h165625[56:34];
      3'h2:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d4331 =
	      IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d4327;
      3'h3:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d4331 =
	      IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_requestR_ETC___d4325;
      3'h4:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d4331 =
	      CASE_guard56369_0b0_theResult___snd65625_BITS__ETC__q141;
      default: IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d4331 =
		   23'd0;
    endcase
  end
  always@(guard__h156369 or
	  _theResult___snd__h165625 or
	  out_sfd__h166160 or _theResult___sfd__h166157)
  begin
    case (guard__h156369)
      2'b0, 2'b01:
	  CASE_guard56369_0b0_theResult___snd65625_BITS__ETC__q142 =
	      _theResult___snd__h165625[56:34];
      2'b10:
	  CASE_guard56369_0b0_theResult___snd65625_BITS__ETC__q142 =
	      out_sfd__h166160;
      2'b11:
	  CASE_guard56369_0b0_theResult___snd65625_BITS__ETC__q142 =
	      _theResult___sfd__h166157;
    endcase
  end
  always@(guard__h126038 or requestR_BITS_191_TO_128__q1)
  begin
    case (guard__h126038)
      2'b0, 2'b01, 2'b10:
	  CASE_guard26038_0b0_requestR_BITS_191_TO_128_B_ETC__q143 =
	      requestR_BITS_191_TO_128__q1[63];
      2'd3:
	  CASE_guard26038_0b0_requestR_BITS_191_TO_128_B_ETC__q143 =
	      guard__h126038 == 2'b11 && requestR_BITS_191_TO_128__q1[63];
    endcase
  end
  always@(requestR or requestR_BITS_191_TO_128__q1 or guard__h126038)
  begin
    case (requestR[194:192])
      3'h2, 3'h3:
	  CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q144 =
	      requestR_BITS_191_TO_128__q1[63];
      3'h4:
	  CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q144 =
	      (guard__h126038 == 2'b0) ?
		requestR_BITS_191_TO_128__q1[63] :
		(guard__h126038 == 2'b01 || guard__h126038 == 2'b10 ||
		 guard__h126038 == 2'b11) &&
		requestR_BITS_191_TO_128__q1[63];
      default: CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q144 =
		   requestR[194:192] == 3'h1 &&
		   requestR_BITS_191_TO_128__q1[63];
    endcase
  end
  always@(guard__h136028 or requestR_BITS_191_TO_128__q1)
  begin
    case (guard__h136028)
      2'b0, 2'b01, 2'b10:
	  CASE_guard36028_0b0_requestR_BITS_191_TO_128_B_ETC__q145 =
	      requestR_BITS_191_TO_128__q1[63];
      2'd3:
	  CASE_guard36028_0b0_requestR_BITS_191_TO_128_B_ETC__q145 =
	      guard__h136028 == 2'b11 && requestR_BITS_191_TO_128__q1[63];
    endcase
  end
  always@(requestR or requestR_BITS_191_TO_128__q1 or guard__h136028)
  begin
    case (requestR[194:192])
      3'h2, 3'h3:
	  CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q146 =
	      requestR_BITS_191_TO_128__q1[63];
      3'h4:
	  CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q146 =
	      (guard__h136028 == 2'b0) ?
		requestR_BITS_191_TO_128__q1[63] :
		(guard__h136028 == 2'b01 || guard__h136028 == 2'b10 ||
		 guard__h136028 == 2'b11) &&
		requestR_BITS_191_TO_128__q1[63];
      default: CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q146 =
		   requestR[194:192] == 3'h1 &&
		   requestR_BITS_191_TO_128__q1[63];
    endcase
  end
  always@(guard__h146250 or requestR_BITS_191_TO_128__q1)
  begin
    case (guard__h146250)
      2'b0, 2'b01, 2'b10:
	  CASE_guard46250_0b0_requestR_BITS_191_TO_128_B_ETC__q147 =
	      requestR_BITS_191_TO_128__q1[63];
      2'd3:
	  CASE_guard46250_0b0_requestR_BITS_191_TO_128_B_ETC__q147 =
	      guard__h146250 == 2'b11 && requestR_BITS_191_TO_128__q1[63];
    endcase
  end
  always@(requestR or requestR_BITS_191_TO_128__q1 or guard__h146250)
  begin
    case (requestR[194:192])
      3'h2, 3'h3:
	  CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q148 =
	      requestR_BITS_191_TO_128__q1[63];
      3'h4:
	  CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q148 =
	      (guard__h146250 == 2'b0) ?
		requestR_BITS_191_TO_128__q1[63] :
		(guard__h146250 == 2'b01 || guard__h146250 == 2'b10 ||
		 guard__h146250 == 2'b11) &&
		requestR_BITS_191_TO_128__q1[63];
      default: CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q148 =
		   requestR[194:192] == 3'h1 &&
		   requestR_BITS_191_TO_128__q1[63];
    endcase
  end
  always@(guard__h156369 or requestR_BITS_191_TO_128__q1)
  begin
    case (guard__h156369)
      2'b0, 2'b01, 2'b10:
	  CASE_guard56369_0b0_requestR_BITS_191_TO_128_B_ETC__q149 =
	      requestR_BITS_191_TO_128__q1[63];
      2'd3:
	  CASE_guard56369_0b0_requestR_BITS_191_TO_128_B_ETC__q149 =
	      guard__h156369 == 2'b11 && requestR_BITS_191_TO_128__q1[63];
    endcase
  end
  always@(requestR or requestR_BITS_191_TO_128__q1 or guard__h156369)
  begin
    case (requestR[194:192])
      3'h2, 3'h3:
	  CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q150 =
	      requestR_BITS_191_TO_128__q1[63];
      3'h4:
	  CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q150 =
	      (guard__h156369 == 2'b0) ?
		requestR_BITS_191_TO_128__q1[63] :
		(guard__h156369 == 2'b01 || guard__h156369 == 2'b10 ||
		 guard__h156369 == 2'b11) &&
		requestR_BITS_191_TO_128__q1[63];
      default: CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q150 =
		   requestR[194:192] == 3'h1 &&
		   requestR_BITS_191_TO_128__q1[63];
    endcase
  end
  always@(guard__h181312 or
	  _theResult___fst_exp__h190506 or _theResult___exp__h191161)
  begin
    case (guard__h181312)
      2'b0:
	  CASE_guard81312_0b0_theResult___fst_exp90506_0_ETC__q159 =
	      _theResult___fst_exp__h190506;
      2'b01, 2'b10, 2'b11:
	  CASE_guard81312_0b0_theResult___fst_exp90506_0_ETC__q159 =
	      _theResult___exp__h191161;
    endcase
  end
  always@(requestR or
	  _theResult___fst_exp__h190506 or
	  IF_IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d4669 or
	  IF_IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d4667 or
	  CASE_guard81312_0b0_theResult___fst_exp90506_0_ETC__q159)
  begin
    case (requestR[194:192])
      3'h1:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d4673 =
	      _theResult___fst_exp__h190506;
      3'h2:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d4673 =
	      IF_IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d4669;
      3'h3:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d4673 =
	      IF_IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d4667;
      3'h4:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d4673 =
	      CASE_guard81312_0b0_theResult___fst_exp90506_0_ETC__q159;
      default: IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d4673 =
		   11'd0;
    endcase
  end
  always@(guard__h181312 or
	  _theResult___fst_exp__h190506 or
	  out_exp__h191164 or _theResult___exp__h191161)
  begin
    case (guard__h181312)
      2'b0, 2'b01:
	  CASE_guard81312_0b0_theResult___fst_exp90506_0_ETC__q160 =
	      _theResult___fst_exp__h190506;
      2'b10:
	  CASE_guard81312_0b0_theResult___fst_exp90506_0_ETC__q160 =
	      out_exp__h191164;
      2'b11:
	  CASE_guard81312_0b0_theResult___fst_exp90506_0_ETC__q160 =
	      _theResult___exp__h191161;
    endcase
  end
  always@(guard__h191853 or
	  _theResult___fst_exp__h201334 or _theResult___exp__h202063)
  begin
    case (guard__h191853)
      2'b0:
	  CASE_guard91853_0b0_theResult___fst_exp01334_0_ETC__q161 =
	      _theResult___fst_exp__h201334;
      2'b01, 2'b10, 2'b11:
	  CASE_guard91853_0b0_theResult___fst_exp01334_0_ETC__q161 =
	      _theResult___exp__h202063;
    endcase
  end
  always@(requestR or
	  _theResult___fst_exp__h201334 or
	  IF_IF_IF_IF_3074_MINUS_SEXT_IF_IF_requestR_3_B_ETC___d4994 or
	  IF_IF_IF_IF_3074_MINUS_SEXT_IF_IF_requestR_3_B_ETC___d4992 or
	  CASE_guard91853_0b0_theResult___fst_exp01334_0_ETC__q161)
  begin
    case (requestR[194:192])
      3'h1:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d4998 =
	      _theResult___fst_exp__h201334;
      3'h2:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d4998 =
	      IF_IF_IF_IF_3074_MINUS_SEXT_IF_IF_requestR_3_B_ETC___d4994;
      3'h3:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d4998 =
	      IF_IF_IF_IF_3074_MINUS_SEXT_IF_IF_requestR_3_B_ETC___d4992;
      3'h4:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d4998 =
	      CASE_guard91853_0b0_theResult___fst_exp01334_0_ETC__q161;
      default: IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d4998 =
		   11'd0;
    endcase
  end
  always@(guard__h191853 or
	  _theResult___fst_exp__h201334 or
	  out_exp__h202066 or _theResult___exp__h202063)
  begin
    case (guard__h191853)
      2'b0, 2'b01:
	  CASE_guard91853_0b0_theResult___fst_exp01334_0_ETC__q162 =
	      _theResult___fst_exp__h201334;
      2'b10:
	  CASE_guard91853_0b0_theResult___fst_exp01334_0_ETC__q162 =
	      out_exp__h202066;
      2'b11:
	  CASE_guard91853_0b0_theResult___fst_exp01334_0_ETC__q162 =
	      _theResult___exp__h202063;
    endcase
  end
  always@(guard__h202175 or
	  _theResult___fst_exp__h211398 or _theResult___exp__h212078)
  begin
    case (guard__h202175)
      2'b0:
	  CASE_guard02175_0b0_theResult___fst_exp11398_0_ETC__q163 =
	      _theResult___fst_exp__h211398;
      2'b01, 2'b10, 2'b11:
	  CASE_guard02175_0b0_theResult___fst_exp11398_0_ETC__q163 =
	      _theResult___exp__h212078;
    endcase
  end
  always@(requestR or
	  _theResult___fst_exp__h211398 or
	  IF_IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d5063 or
	  IF_IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d5061 or
	  CASE_guard02175_0b0_theResult___fst_exp11398_0_ETC__q163)
  begin
    case (requestR[194:192])
      3'h1:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d5067 =
	      _theResult___fst_exp__h211398;
      3'h2:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d5067 =
	      IF_IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d5063;
      3'h3:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d5067 =
	      IF_IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d5061;
      3'h4:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d5067 =
	      CASE_guard02175_0b0_theResult___fst_exp11398_0_ETC__q163;
      default: IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d5067 =
		   11'd0;
    endcase
  end
  always@(guard__h202175 or
	  _theResult___fst_exp__h211398 or
	  out_exp__h212081 or _theResult___exp__h212078)
  begin
    case (guard__h202175)
      2'b0, 2'b01:
	  CASE_guard02175_0b0_theResult___fst_exp11398_0_ETC__q164 =
	      _theResult___fst_exp__h211398;
      2'b10:
	  CASE_guard02175_0b0_theResult___fst_exp11398_0_ETC__q164 =
	      out_exp__h212081;
      2'b11:
	  CASE_guard02175_0b0_theResult___fst_exp11398_0_ETC__q164 =
	      _theResult___exp__h212078;
    endcase
  end
  always@(guard__h181312 or requestR_BITS_191_TO_128__q1)
  begin
    case (guard__h181312)
      2'b0, 2'b01, 2'b10:
	  CASE_guard81312_0b0_requestR_BITS_191_TO_128_B_ETC__q165 =
	      requestR_BITS_191_TO_128__q1[63:32] == 32'hFFFFFFFF &&
	      requestR_BITS_191_TO_128__q1[31];
      2'd3:
	  CASE_guard81312_0b0_requestR_BITS_191_TO_128_B_ETC__q165 =
	      guard__h181312 == 2'b11 &&
	      requestR_BITS_191_TO_128__q1[63:32] == 32'hFFFFFFFF &&
	      requestR_BITS_191_TO_128__q1[31];
    endcase
  end
  always@(requestR or requestR_BITS_191_TO_128__q1 or guard__h181312)
  begin
    case (requestR[194:192])
      3'h2, 3'h3:
	  CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q166 =
	      requestR_BITS_191_TO_128__q1[63:32] == 32'hFFFFFFFF &&
	      requestR_BITS_191_TO_128__q1[31];
      3'h4:
	  CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q166 =
	      (guard__h181312 == 2'b0) ?
		requestR_BITS_191_TO_128__q1[63:32] == 32'hFFFFFFFF &&
		requestR_BITS_191_TO_128__q1[31] :
		(guard__h181312 == 2'b01 || guard__h181312 == 2'b10 ||
		 guard__h181312 == 2'b11) &&
		requestR_BITS_191_TO_128__q1[63:32] == 32'hFFFFFFFF &&
		requestR_BITS_191_TO_128__q1[31];
      default: CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q166 =
		   requestR[194:192] == 3'h1 &&
		   requestR_BITS_191_TO_128__q1[63:32] == 32'hFFFFFFFF &&
		   requestR_BITS_191_TO_128__q1[31];
    endcase
  end
  always@(guard__h191853 or requestR_BITS_191_TO_128__q1)
  begin
    case (guard__h191853)
      2'b0, 2'b01, 2'b10:
	  CASE_guard91853_0b0_requestR_BITS_191_TO_128_B_ETC__q167 =
	      requestR_BITS_191_TO_128__q1[63:32] == 32'hFFFFFFFF &&
	      requestR_BITS_191_TO_128__q1[31];
      2'd3:
	  CASE_guard91853_0b0_requestR_BITS_191_TO_128_B_ETC__q167 =
	      guard__h191853 == 2'b11 &&
	      requestR_BITS_191_TO_128__q1[63:32] == 32'hFFFFFFFF &&
	      requestR_BITS_191_TO_128__q1[31];
    endcase
  end
  always@(requestR or requestR_BITS_191_TO_128__q1 or guard__h191853)
  begin
    case (requestR[194:192])
      3'h2, 3'h3:
	  CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q168 =
	      requestR_BITS_191_TO_128__q1[63:32] == 32'hFFFFFFFF &&
	      requestR_BITS_191_TO_128__q1[31];
      3'h4:
	  CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q168 =
	      (guard__h191853 == 2'b0) ?
		requestR_BITS_191_TO_128__q1[63:32] == 32'hFFFFFFFF &&
		requestR_BITS_191_TO_128__q1[31] :
		(guard__h191853 == 2'b01 || guard__h191853 == 2'b10 ||
		 guard__h191853 == 2'b11) &&
		requestR_BITS_191_TO_128__q1[63:32] == 32'hFFFFFFFF &&
		requestR_BITS_191_TO_128__q1[31];
      default: CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q168 =
		   requestR[194:192] == 3'h1 &&
		   requestR_BITS_191_TO_128__q1[63:32] == 32'hFFFFFFFF &&
		   requestR_BITS_191_TO_128__q1[31];
    endcase
  end
  always@(guard__h202175 or requestR_BITS_191_TO_128__q1)
  begin
    case (guard__h202175)
      2'b0, 2'b01, 2'b10:
	  CASE_guard02175_0b0_requestR_BITS_191_TO_128_B_ETC__q169 =
	      requestR_BITS_191_TO_128__q1[63:32] == 32'hFFFFFFFF &&
	      requestR_BITS_191_TO_128__q1[31];
      2'd3:
	  CASE_guard02175_0b0_requestR_BITS_191_TO_128_B_ETC__q169 =
	      guard__h202175 == 2'b11 &&
	      requestR_BITS_191_TO_128__q1[63:32] == 32'hFFFFFFFF &&
	      requestR_BITS_191_TO_128__q1[31];
    endcase
  end
  always@(requestR or requestR_BITS_191_TO_128__q1 or guard__h202175)
  begin
    case (requestR[194:192])
      3'h2, 3'h3:
	  CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q170 =
	      requestR_BITS_191_TO_128__q1[63:32] == 32'hFFFFFFFF &&
	      requestR_BITS_191_TO_128__q1[31];
      3'h4:
	  CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q170 =
	      (guard__h202175 == 2'b0) ?
		requestR_BITS_191_TO_128__q1[63:32] == 32'hFFFFFFFF &&
		requestR_BITS_191_TO_128__q1[31] :
		(guard__h202175 == 2'b01 || guard__h202175 == 2'b10 ||
		 guard__h202175 == 2'b11) &&
		requestR_BITS_191_TO_128__q1[63:32] == 32'hFFFFFFFF &&
		requestR_BITS_191_TO_128__q1[31];
      default: CASE_requestR_BITS_194_TO_192_0x2_requestR_BIT_ETC__q170 =
		   requestR[194:192] == 3'h1 &&
		   requestR_BITS_191_TO_128__q1[63:32] == 32'hFFFFFFFF &&
		   requestR_BITS_191_TO_128__q1[31];
    endcase
  end
  always@(guard__h181312 or
	  _theResult___snd__h190457 or _theResult___sfd__h191162)
  begin
    case (guard__h181312)
      2'b0:
	  CASE_guard81312_0b0_theResult___snd90457_BITS__ETC__q171 =
	      _theResult___snd__h190457[56:5];
      2'b01, 2'b10, 2'b11:
	  CASE_guard81312_0b0_theResult___snd90457_BITS__ETC__q171 =
	      _theResult___sfd__h191162;
    endcase
  end
  always@(requestR or
	  _theResult___snd__h190457 or
	  IF_IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d5096 or
	  IF_IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d5094 or
	  CASE_guard81312_0b0_theResult___snd90457_BITS__ETC__q171)
  begin
    case (requestR[194:192])
      3'h1:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d5100 =
	      _theResult___snd__h190457[56:5];
      3'h2:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d5100 =
	      IF_IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d5096;
      3'h3:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d5100 =
	      IF_IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d5094;
      3'h4:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d5100 =
	      CASE_guard81312_0b0_theResult___snd90457_BITS__ETC__q171;
      default: IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d5100 =
		   52'd0;
    endcase
  end
  always@(guard__h181312 or
	  _theResult___snd__h190457 or
	  out_sfd__h191165 or _theResult___sfd__h191162)
  begin
    case (guard__h181312)
      2'b0, 2'b01:
	  CASE_guard81312_0b0_theResult___snd90457_BITS__ETC__q172 =
	      _theResult___snd__h190457[56:5];
      2'b10:
	  CASE_guard81312_0b0_theResult___snd90457_BITS__ETC__q172 =
	      out_sfd__h191165;
      2'b11:
	  CASE_guard81312_0b0_theResult___snd90457_BITS__ETC__q172 =
	      _theResult___sfd__h191162;
    endcase
  end
  always@(guard__h191853 or sfdin__h201328 or _theResult___sfd__h202064)
  begin
    case (guard__h191853)
      2'b0:
	  CASE_guard91853_0b0_sfdin01328_BITS_56_TO_5_0b_ETC__q173 =
	      sfdin__h201328[56:5];
      2'b01, 2'b10, 2'b11:
	  CASE_guard91853_0b0_sfdin01328_BITS_56_TO_5_0b_ETC__q173 =
	      _theResult___sfd__h202064;
    endcase
  end
  always@(requestR or
	  sfdin__h201328 or
	  IF_IF_IF_IF_3074_MINUS_SEXT_IF_IF_requestR_3_B_ETC___d5123 or
	  IF_IF_IF_IF_3074_MINUS_SEXT_IF_IF_requestR_3_B_ETC___d5121 or
	  CASE_guard91853_0b0_sfdin01328_BITS_56_TO_5_0b_ETC__q173)
  begin
    case (requestR[194:192])
      3'h1:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d5127 =
	      sfdin__h201328[56:5];
      3'h2:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d5127 =
	      IF_IF_IF_IF_3074_MINUS_SEXT_IF_IF_requestR_3_B_ETC___d5123;
      3'h3:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d5127 =
	      IF_IF_IF_IF_3074_MINUS_SEXT_IF_IF_requestR_3_B_ETC___d5121;
      3'h4:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d5127 =
	      CASE_guard91853_0b0_sfdin01328_BITS_56_TO_5_0b_ETC__q173;
      default: IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d5127 =
		   52'd0;
    endcase
  end
  always@(guard__h191853 or
	  sfdin__h201328 or out_sfd__h202067 or _theResult___sfd__h202064)
  begin
    case (guard__h191853)
      2'b0, 2'b01:
	  CASE_guard91853_0b0_sfdin01328_BITS_56_TO_5_0b_ETC__q174 =
	      sfdin__h201328[56:5];
      2'b10:
	  CASE_guard91853_0b0_sfdin01328_BITS_56_TO_5_0b_ETC__q174 =
	      out_sfd__h202067;
      2'b11:
	  CASE_guard91853_0b0_sfdin01328_BITS_56_TO_5_0b_ETC__q174 =
	      _theResult___sfd__h202064;
    endcase
  end
  always@(guard__h202175 or
	  _theResult___snd__h211344 or _theResult___sfd__h212079)
  begin
    case (guard__h202175)
      2'b0:
	  CASE_guard02175_0b0_theResult___snd11344_BITS__ETC__q175 =
	      _theResult___snd__h211344[56:5];
      2'b01, 2'b10, 2'b11:
	  CASE_guard02175_0b0_theResult___snd11344_BITS__ETC__q175 =
	      _theResult___sfd__h212079;
    endcase
  end
  always@(requestR or
	  _theResult___snd__h211344 or
	  IF_IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d5142 or
	  IF_IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d5140 or
	  CASE_guard02175_0b0_theResult___snd11344_BITS__ETC__q175)
  begin
    case (requestR[194:192])
      3'h1:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d5146 =
	      _theResult___snd__h211344[56:5];
      3'h2:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d5146 =
	      IF_IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d5142;
      3'h3:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d5146 =
	      IF_IF_IF_IF_IF_requestR_3_BIT_214_4_THEN_reque_ETC___d5140;
      3'h4:
	  IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d5146 =
	      CASE_guard02175_0b0_theResult___snd11344_BITS__ETC__q175;
      default: IF_IF_requestR_3_BIT_214_4_THEN_requestR_3_BIT_ETC___d5146 =
		   52'd0;
    endcase
  end
  always@(guard__h202175 or
	  _theResult___snd__h211344 or
	  out_sfd__h212082 or _theResult___sfd__h212079)
  begin
    case (guard__h202175)
      2'b0, 2'b01:
	  CASE_guard02175_0b0_theResult___snd11344_BITS__ETC__q176 =
	      _theResult___snd__h211344[56:5];
      2'b10:
	  CASE_guard02175_0b0_theResult___snd11344_BITS__ETC__q176 =
	      out_sfd__h212082;
      2'b11:
	  CASE_guard02175_0b0_theResult___snd11344_BITS__ETC__q176 =
	      _theResult___sfd__h212079;
    endcase
  end
  // handling of inlined registers
  always@(posedge CLK)
  begin
    if (RST_N == `BSV_RESET_VALUE)
      begin
        stateR <= `BSV_ASSIGNMENT_DELAY 2'd0;
      end
    else
      begin
        if (stateR$EN) stateR <= `BSV_ASSIGNMENT_DELAY stateR$D_IN;
      end
    if (requestR$EN) requestR <= `BSV_ASSIGNMENT_DELAY requestR$D_IN;
    if (resultR$EN) resultR <= `BSV_ASSIGNMENT_DELAY resultR$D_IN;
  end
  // synopsys translate_off
  `ifdef BSV_NO_INITIAL_BLOCKS
  `else // not BSV_NO_INITIAL_BLOCKS
  initial
  begin
    requestR = 215'h2AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
    resultR = 70'h2AAAAAAAAAAAAAAAAA;
    stateR = 2'h2;
  end
  `endif // BSV_NO_INITIAL_BLOCKS
  // synopsys translate_on
  // handling of system tasks
  // synopsys translate_off
  always@(negedge CLK)
  begin
    #0;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFADD_S && NOT_verbosity_ULE_1_6___d27)
	begin
	  v__h1224 = $stime;
	  #0;
	end
    v__h1218 = v__h1224 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFADD_S && NOT_verbosity_ULE_1_6___d27)
	$display("%0d: FBox_Core.doFADD: ", v__h1218);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFSUB_S && NOT_verbosity_ULE_1_6___d27)
	begin
	  v__h1777 = $stime;
	  #0;
	end
    v__h1771 = v__h1777 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFSUB_S && NOT_verbosity_ULE_1_6___d27)
	$display("%0d: FBox_Core.doFSUB: ", v__h1771);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFMUL_S && NOT_verbosity_ULE_1_6___d27)
	begin
	  v__h1966 = $stime;
	  #0;
	end
    v__h1960 = v__h1966 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFMUL_S && NOT_verbosity_ULE_1_6___d27)
	$display("%0d: FBox_Core.doFMUL: ", v__h1960);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFMADD_S && NOT_verbosity_ULE_1_6___d27)
	begin
	  v__h2168 = $stime;
	  #0;
	end
    v__h2162 = v__h2168 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFMADD_S && NOT_verbosity_ULE_1_6___d27)
	$display("%0d: FBox_Core.doFMADD_S ", v__h2162);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFMSUB_S && NOT_verbosity_ULE_1_6___d27)
	begin
	  v__h2418 = $stime;
	  #0;
	end
    v__h2412 = v__h2418 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFMSUB_S && NOT_verbosity_ULE_1_6___d27)
	$display("%0d: FBox_Core.doFMSUB_S ", v__h2412);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFNMADD_S && NOT_verbosity_ULE_1_6___d27)
	begin
	  v__h2593 = $stime;
	  #0;
	end
    v__h2587 = v__h2593 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFNMADD_S && NOT_verbosity_ULE_1_6___d27)
	$display("%0d: FBox_Core.doFNMADD_S ", v__h2587);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFNMSUB_S && NOT_verbosity_ULE_1_6___d27)
	begin
	  v__h2768 = $stime;
	  #0;
	end
    v__h2762 = v__h2768 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFNMSUB_S && NOT_verbosity_ULE_1_6___d27)
	$display("%0d: FBox_Core.doFNMSUB_S ", v__h2762);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFDIV_S && NOT_verbosity_ULE_1_6___d27)
	begin
	  v__h2950 = $stime;
	  #0;
	end
    v__h2944 = v__h2950 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFDIV_S && NOT_verbosity_ULE_1_6___d27)
	$display("%0d: FBox_Core.doFDIV_S ", v__h2944);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFSQRT_S && NOT_verbosity_ULE_1_6___d27)
	begin
	  v__h3139 = $stime;
	  #0;
	end
    v__h3133 = v__h3139 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFSQRT_S && NOT_verbosity_ULE_1_6___d27)
	$display("%0d: FBox_Core.doFSQRT_S ", v__h3133);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFSGNJ_S && NOT_verbosity_ULE_1_6___d27)
	begin
	  v__h3337 = $stime;
	  #0;
	end
    v__h3331 = v__h3337 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFSGNJ_S && NOT_verbosity_ULE_1_6___d27)
	$display("%0d: FBox_Core.doFSGNJ_S ", v__h3331);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFSGNJN_S && NOT_verbosity_ULE_1_6___d27)
	begin
	  v__h3520 = $stime;
	  #0;
	end
    v__h3514 = v__h3520 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFSGNJN_S && NOT_verbosity_ULE_1_6___d27)
	$display("%0d: FBox_Core.doFSGNJN_S ", v__h3514);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFSGNJX_S && NOT_verbosity_ULE_1_6___d27)
	begin
	  v__h3693 = $stime;
	  #0;
	end
    v__h3687 = v__h3693 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFSGNJX_S && NOT_verbosity_ULE_1_6___d27)
	$display("%0d: FBox_Core.doFSGNJX_S ", v__h3687);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFCVT_S_L && NOT_verbosity_ULE_1_6___d27)
	begin
	  v__h3882 = $stime;
	  #0;
	end
    v__h3876 = v__h3882 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFCVT_S_L && NOT_verbosity_ULE_1_6___d27)
	$display("%0d: FBox_Core.doFCVT_S_L ", v__h3876);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFCVT_S_L && NOT_verbosity_ULE_2_01___d702)
	$write("v1 = %08x, rmd = ", requestR[191:128]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFCVT_S_L && NOT_verbosity_ULE_2_01___d702 &&
	  (requestR[194:192] == 3'h0 ||
	   requestR[194:192] != 3'h1 && requestR[194:192] != 3'h2 &&
	   requestR[194:192] != 3'h3 &&
	   requestR[194:192] != 3'h4))
	$write("<Round Mode: Nearest Even>");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFCVT_S_L && NOT_verbosity_ULE_2_01___d702 &&
	  requestR[194:192] == 3'h4)
	$write("<Round Mode: Nearest Away From Zero>");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFCVT_S_L && NOT_verbosity_ULE_2_01___d702 &&
	  requestR[194:192] == 3'h3)
	$write("<Round Mode: +Infinity>");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFCVT_S_L && NOT_verbosity_ULE_2_01___d702 &&
	  requestR[194:192] == 3'h2)
	$write("<Round Mode: -Infinity>");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFCVT_S_L && NOT_verbosity_ULE_2_01___d702 &&
	  requestR[194:192] == 3'h1)
	$write("<Round Mode: Zero>");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFCVT_S_L && NOT_verbosity_ULE_2_01___d702)
	$write("\n");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFCVT_S_L && NOT_verbosity_ULE_2_01___d702)
	$display("    Result: (%08x, %05b)", res__h3932, fcsr__h3933);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFCVT_S_LU && NOT_verbosity_ULE_1_6___d27)
	begin
	  v__h16640 = $stime;
	  #0;
	end
    v__h16634 = v__h16640 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFCVT_S_LU && NOT_verbosity_ULE_1_6___d27)
	$display("%0d: FBox_Core.doFCVT_S_LU ", v__h16634);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFCVT_S_W && NOT_verbosity_ULE_1_6___d27)
	begin
	  v__h28741 = $stime;
	  #0;
	end
    v__h28735 = v__h28741 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFCVT_S_W && NOT_verbosity_ULE_1_6___d27)
	$display("%0d: FBox_Core.doFCVT_S_W ", v__h28735);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFCVT_S_WU && NOT_verbosity_ULE_1_6___d27)
	begin
	  v__h35941 = $stime;
	  #0;
	end
    v__h35935 = v__h35941 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFCVT_S_WU && NOT_verbosity_ULE_1_6___d27)
	$display("%0d: FBox_Core.doFCVT_S_WU ", v__h35935);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFCVT_L_S && NOT_verbosity_ULE_1_6___d27)
	begin
	  v__h42829 = $stime;
	  #0;
	end
    v__h42823 = v__h42829 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFCVT_L_S && NOT_verbosity_ULE_1_6___d27)
	$display("%0d: FBox_Core.doFCVT_L_S ", v__h42823);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFCVT_LU_S && NOT_verbosity_ULE_1_6___d27)
	begin
	  v__h44905 = $stime;
	  #0;
	end
    v__h44899 = v__h44905 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFCVT_LU_S && NOT_verbosity_ULE_1_6___d27)
	$display("%0d: FBox_Core.doFCVT_LU_S ", v__h44899);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFCVT_W_S && NOT_verbosity_ULE_1_6___d27)
	begin
	  v__h45689 = $stime;
	  #0;
	end
    v__h45683 = v__h45689 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFCVT_W_S && NOT_verbosity_ULE_1_6___d27)
	$display("%0d: FBox_Core.doFCVT_W_S ", v__h45683);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFCVT_WU_S && NOT_verbosity_ULE_1_6___d27)
	begin
	  v__h47303 = $stime;
	  #0;
	end
    v__h47297 = v__h47303 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFCVT_WU_S && NOT_verbosity_ULE_1_6___d27)
	$display("%0d: FBox_Core.doFCVT_WU_S ", v__h47297);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFMIN_S && NOT_verbosity_ULE_1_6___d27)
	begin
	  v__h48090 = $stime;
	  #0;
	end
    v__h48084 = v__h48090 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFMIN_S && NOT_verbosity_ULE_1_6___d27)
	$display("%0d: FBox_Core.doFMIN_S ", v__h48084);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFMAX_S && NOT_verbosity_ULE_1_6___d27)
	begin
	  v__h50764 = $stime;
	  #0;
	end
    v__h50758 = v__h50764 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFMAX_S && NOT_verbosity_ULE_1_6___d27)
	$display("%0d: FBox_Core.doFMAX_S ", v__h50758);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFMV_W_X && NOT_verbosity_ULE_1_6___d27)
	begin
	  v__h53335 = $stime;
	  #0;
	end
    v__h53329 = v__h53335 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFMV_W_X && NOT_verbosity_ULE_1_6___d27)
	$display("%0d: FBox_Core.doFMV_W_X ", v__h53329);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFMV_X_W && NOT_verbosity_ULE_1_6___d27)
	begin
	  v__h53495 = $stime;
	  #0;
	end
    v__h53489 = v__h53495 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFMV_X_W && NOT_verbosity_ULE_1_6___d27)
	$display("%0d: FBox_Core.doFMV_X_W ", v__h53489);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFEQ_S && NOT_verbosity_ULE_1_6___d27)
	begin
	  v__h53671 = $stime;
	  #0;
	end
    v__h53665 = v__h53671 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFEQ_S && NOT_verbosity_ULE_1_6___d27)
	$display("%0d: FBox_Core.doFEQ_S ", v__h53665);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFLT_S && NOT_verbosity_ULE_1_6___d27)
	begin
	  v__h55194 = $stime;
	  #0;
	end
    v__h55188 = v__h55194 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFLT_S && NOT_verbosity_ULE_1_6___d27)
	$display("%0d: FBox_Core.doFLT_S ", v__h55188);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFLE_S && NOT_verbosity_ULE_1_6___d27)
	begin
	  v__h56303 = $stime;
	  #0;
	end
    v__h56297 = v__h56303 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFLE_S && NOT_verbosity_ULE_1_6___d27)
	$display("%0d: FBox_Core.doFLE_S ", v__h56297);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFCLASS_S && NOT_verbosity_ULE_1_6___d27)
	begin
	  v__h57430 = $stime;
	  #0;
	end
    v__h57424 = v__h57430 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFCLASS_S && NOT_verbosity_ULE_1_6___d27)
	$display("%0d: FBox_Core.doFCLASS_S ", v__h57424);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFADD_D && NOT_verbosity_ULE_1_6___d27)
	begin
	  v__h57911 = $stime;
	  #0;
	end
    v__h57905 = v__h57911 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFADD_D && NOT_verbosity_ULE_1_6___d27)
	$display("%0d: FBox_Core.doFADD_D ", v__h57905);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFSUB_D && NOT_verbosity_ULE_1_6___d27)
	begin
	  v__h58124 = $stime;
	  #0;
	end
    v__h58118 = v__h58124 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFSUB_D && NOT_verbosity_ULE_1_6___d27)
	$display("%0d: FBox_Core.doFSUB_D ", v__h58118);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFMUL_D && NOT_verbosity_ULE_1_6___d27)
	begin
	  v__h58311 = $stime;
	  #0;
	end
    v__h58305 = v__h58311 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFMUL_D && NOT_verbosity_ULE_1_6___d27)
	$display("%0d: FBox_Core.doFMUL_D ", v__h58305);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFMADD_D && NOT_verbosity_ULE_1_6___d27)
	begin
	  v__h58491 = $stime;
	  #0;
	end
    v__h58485 = v__h58491 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFMADD_D && NOT_verbosity_ULE_1_6___d27)
	$display("%0d: FBox_Core.doFMADD_D ", v__h58485);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFMSUB_D && NOT_verbosity_ULE_1_6___d27)
	begin
	  v__h58676 = $stime;
	  #0;
	end
    v__h58670 = v__h58676 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFMSUB_D && NOT_verbosity_ULE_1_6___d27)
	$display("%0d: FBox_Core.doFMSUB_D ", v__h58670);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFNMADD_D && NOT_verbosity_ULE_1_6___d27)
	begin
	  v__h58848 = $stime;
	  #0;
	end
    v__h58842 = v__h58848 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFNMADD_D && NOT_verbosity_ULE_1_6___d27)
	$display("%0d: FBox_Core.doFNMADD_D ", v__h58842);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFNMSUB_D && NOT_verbosity_ULE_1_6___d27)
	begin
	  v__h59020 = $stime;
	  #0;
	end
    v__h59014 = v__h59020 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFNMSUB_D && NOT_verbosity_ULE_1_6___d27)
	$display("%0d: FBox_Core.doFNMSUB_D ", v__h59014);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFDIV_D && NOT_verbosity_ULE_1_6___d27)
	begin
	  v__h59199 = $stime;
	  #0;
	end
    v__h59193 = v__h59199 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFDIV_D && NOT_verbosity_ULE_1_6___d27)
	$display("%0d: FBox_Core.doFDIV_D ", v__h59193);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFSQRT_D && NOT_verbosity_ULE_1_6___d27)
	begin
	  v__h59386 = $stime;
	  #0;
	end
    v__h59380 = v__h59386 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFSQRT_D && NOT_verbosity_ULE_1_6___d27)
	$display("%0d: FBox_Core.doFSQRT_D ", v__h59380);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFSGNJ_D && NOT_verbosity_ULE_1_6___d27)
	begin
	  v__h59583 = $stime;
	  #0;
	end
    v__h59577 = v__h59583 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFSGNJ_D && NOT_verbosity_ULE_1_6___d27)
	$display("%0d: FBox_Core.doFSGNJ_D ", v__h59577);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFSGNJN_D && NOT_verbosity_ULE_1_6___d27)
	begin
	  v__h59744 = $stime;
	  #0;
	end
    v__h59738 = v__h59744 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFSGNJN_D && NOT_verbosity_ULE_1_6___d27)
	$display("%0d: FBox_Core.doFSGNJN_D ", v__h59738);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFSGNJX_D && NOT_verbosity_ULE_1_6___d27)
	begin
	  v__h59907 = $stime;
	  #0;
	end
    v__h59901 = v__h59907 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFSGNJX_D && NOT_verbosity_ULE_1_6___d27)
	$display("%0d: FBox_Core.doFSGNJX_D ", v__h59901);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFCVT_D_W && NOT_verbosity_ULE_1_6___d27)
	begin
	  v__h60075 = $stime;
	  #0;
	end
    v__h60069 = v__h60075 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFCVT_D_W && NOT_verbosity_ULE_1_6___d27)
	$display("%0d: FBox_Core.doFCVT_D_W ", v__h60069);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFCVT_D_WU && NOT_verbosity_ULE_1_6___d27)
	begin
	  v__h71274 = $stime;
	  #0;
	end
    v__h71268 = v__h71274 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFCVT_D_WU && NOT_verbosity_ULE_1_6___d27)
	$display("%0d: FBox_Core.doFCVT_D_WU ", v__h71268);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFCVT_W_D && NOT_verbosity_ULE_1_6___d27)
	begin
	  v__h82193 = $stime;
	  #0;
	end
    v__h82187 = v__h82193 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFCVT_W_D && NOT_verbosity_ULE_1_6___d27)
	$display("%0d: FBox_Core.doFCVT_W_D ", v__h82187);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFCVT_WU_D && NOT_verbosity_ULE_1_6___d27)
	begin
	  v__h83807 = $stime;
	  #0;
	end
    v__h83801 = v__h83807 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFCVT_WU_D && NOT_verbosity_ULE_1_6___d27)
	$display("%0d: FBox_Core.doFCVT_WU_D ", v__h83801);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFCVT_D_L && NOT_verbosity_ULE_1_6___d27)
	begin
	  v__h84594 = $stime;
	  #0;
	end
    v__h84588 = v__h84594 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFCVT_D_L && NOT_verbosity_ULE_1_6___d27)
	$display("%0d: FBox_Core.doFCVT_D_L ", v__h84588);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFCVT_D_LU && NOT_verbosity_ULE_1_6___d27)
	begin
	  v__h97596 = $stime;
	  #0;
	end
    v__h97590 = v__h97596 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFCVT_D_LU && NOT_verbosity_ULE_1_6___d27)
	$display("%0d: FBox_Core.doFCVT_D_LU ", v__h97590);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFCVT_L_D && NOT_verbosity_ULE_1_6___d27)
	begin
	  v__h110093 = $stime;
	  #0;
	end
    v__h110087 = v__h110093 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFCVT_L_D && NOT_verbosity_ULE_1_6___d27)
	$display("%0d: FBox_Core.doFCVT_L_D ", v__h110087);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFCVT_LU_D && NOT_verbosity_ULE_1_6___d27)
	begin
	  v__h112152 = $stime;
	  #0;
	end
    v__h112146 = v__h112152 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFCVT_LU_D && NOT_verbosity_ULE_1_6___d27)
	$display("%0d: FBox_Core.doFCVT_LU_D ", v__h112146);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFCVT_S_D && NOT_verbosity_ULE_1_6___d27)
	begin
	  v__h112936 = $stime;
	  #0;
	end
    v__h112930 = v__h112936 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFCVT_S_D && NOT_verbosity_ULE_1_6___d27)
	$display("%0d: FBox_Core.doFCVT_S_D ", v__h112930);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFCVT_D_S && NOT_verbosity_ULE_1_6___d27)
	begin
	  v__h167802 = $stime;
	  #0;
	end
    v__h167796 = v__h167802 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFCVT_D_S && NOT_verbosity_ULE_1_6___d27)
	$display("%0d: FBox_Core.doFCVT_D_S ", v__h167796);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFMIN_D && NOT_verbosity_ULE_1_6___d27)
	begin
	  v__h213792 = $stime;
	  #0;
	end
    v__h213786 = v__h213792 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFMIN_D && NOT_verbosity_ULE_1_6___d27)
	$display("%0d: FBox_Core.doFMIN_D ", v__h213786);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFMAX_D && NOT_verbosity_ULE_1_6___d27)
	begin
	  v__h218378 = $stime;
	  #0;
	end
    v__h218372 = v__h218378 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFMAX_D && NOT_verbosity_ULE_1_6___d27)
	$display("%0d: FBox_Core.doFMAX_D ", v__h218372);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFEQ_D && NOT_verbosity_ULE_1_6___d27)
	begin
	  v__h222864 = $stime;
	  #0;
	end
    v__h222858 = v__h222864 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFEQ_D && NOT_verbosity_ULE_1_6___d27)
	$display("%0d: FBox_Core.doFEQ_D ", v__h222858);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFLT_D && NOT_verbosity_ULE_1_6___d27)
	begin
	  v__h225599 = $stime;
	  #0;
	end
    v__h225593 = v__h225599 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFLT_D && NOT_verbosity_ULE_1_6___d27)
	$display("%0d: FBox_Core.doFLT_D ", v__h225593);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFLE_D && NOT_verbosity_ULE_1_6___d27)
	begin
	  v__h227516 = $stime;
	  #0;
	end
    v__h227510 = v__h227516 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFLE_D && NOT_verbosity_ULE_1_6___d27)
	$display("%0d: FBox_Core.doFLE_D ", v__h227510);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFMV_D_X && NOT_verbosity_ULE_1_6___d27)
	begin
	  v__h229453 = $stime;
	  #0;
	end
    v__h229447 = v__h229453 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFMV_D_X && NOT_verbosity_ULE_1_6___d27)
	$display("%0d: FBox_Core.doFMV_D_X ", v__h229447);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFMV_X_D && NOT_verbosity_ULE_1_6___d27)
	begin
	  v__h229605 = $stime;
	  #0;
	end
    v__h229599 = v__h229605 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFMV_X_D && NOT_verbosity_ULE_1_6___d27)
	$display("%0d: FBox_Core.doFMV_X_D ", v__h229599);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFCLASS_D && NOT_verbosity_ULE_1_6___d27)
	begin
	  v__h229762 = $stime;
	  #0;
	end
    v__h229756 = v__h229762 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_doFCLASS_D && NOT_verbosity_ULE_1_6___d27)
	$display("%0d: FBox_Core.doFCLASS_D ", v__h229756);
  end
  // synopsys translate_on
endmodule