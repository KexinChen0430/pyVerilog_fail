module outputs
  wire [63 : 0] axi4_slave_rdata;
  wire [3 : 0] axi4_slave_bid, axi4_slave_rid;
  wire [1 : 0] axi4_slave_bresp, axi4_slave_rresp;
  wire RDY_server_reset_request_put,
       RDY_server_reset_response_get,
       RDY_set_addr_map,
       RDY_set_verbosity,
       RDY_show_PLIC_state,
       axi4_slave_arready,
       axi4_slave_awready,
       axi4_slave_bvalid,
       axi4_slave_rlast,
       axi4_slave_rvalid,
       axi4_slave_wready,
       v_targets_0_m_eip,
       v_targets_1_m_eip;
  // register m_cfg_verbosity
  reg [3 : 0] m_cfg_verbosity;
  wire [3 : 0] m_cfg_verbosity$D_IN;
  wire m_cfg_verbosity$EN;
  // register m_rg_addr_base
  reg [63 : 0] m_rg_addr_base;
  wire [63 : 0] m_rg_addr_base$D_IN;
  wire m_rg_addr_base$EN;
  // register m_rg_addr_lim
  reg [63 : 0] m_rg_addr_lim;
  wire [63 : 0] m_rg_addr_lim$D_IN;
  wire m_rg_addr_lim$EN;
  // register m_vrg_source_busy_0
  reg m_vrg_source_busy_0;
  reg m_vrg_source_busy_0$D_IN;
  wire m_vrg_source_busy_0$EN;
  // register m_vrg_source_busy_1
  reg m_vrg_source_busy_1;
  reg m_vrg_source_busy_1$D_IN;
  wire m_vrg_source_busy_1$EN;
  // register m_vrg_source_busy_10
  reg m_vrg_source_busy_10;
  reg m_vrg_source_busy_10$D_IN;
  wire m_vrg_source_busy_10$EN;
  // register m_vrg_source_busy_11
  reg m_vrg_source_busy_11;
  reg m_vrg_source_busy_11$D_IN;
  wire m_vrg_source_busy_11$EN;
  // register m_vrg_source_busy_12
  reg m_vrg_source_busy_12;
  reg m_vrg_source_busy_12$D_IN;
  wire m_vrg_source_busy_12$EN;
  // register m_vrg_source_busy_13
  reg m_vrg_source_busy_13;
  reg m_vrg_source_busy_13$D_IN;
  wire m_vrg_source_busy_13$EN;
  // register m_vrg_source_busy_14
  reg m_vrg_source_busy_14;
  reg m_vrg_source_busy_14$D_IN;
  wire m_vrg_source_busy_14$EN;
  // register m_vrg_source_busy_15
  reg m_vrg_source_busy_15;
  reg m_vrg_source_busy_15$D_IN;
  wire m_vrg_source_busy_15$EN;
  // register m_vrg_source_busy_16
  reg m_vrg_source_busy_16;
  reg m_vrg_source_busy_16$D_IN;
  wire m_vrg_source_busy_16$EN;
  // register m_vrg_source_busy_2
  reg m_vrg_source_busy_2;
  reg m_vrg_source_busy_2$D_IN;
  wire m_vrg_source_busy_2$EN;
  // register m_vrg_source_busy_3
  reg m_vrg_source_busy_3;
  reg m_vrg_source_busy_3$D_IN;
  wire m_vrg_source_busy_3$EN;
  // register m_vrg_source_busy_4
  reg m_vrg_source_busy_4;
  reg m_vrg_source_busy_4$D_IN;
  wire m_vrg_source_busy_4$EN;
  // register m_vrg_source_busy_5
  reg m_vrg_source_busy_5;
  reg m_vrg_source_busy_5$D_IN;
  wire m_vrg_source_busy_5$EN;
  // register m_vrg_source_busy_6
  reg m_vrg_source_busy_6;
  reg m_vrg_source_busy_6$D_IN;
  wire m_vrg_source_busy_6$EN;
  // register m_vrg_source_busy_7
  reg m_vrg_source_busy_7;
  reg m_vrg_source_busy_7$D_IN;
  wire m_vrg_source_busy_7$EN;
  // register m_vrg_source_busy_8
  reg m_vrg_source_busy_8;
  reg m_vrg_source_busy_8$D_IN;
  wire m_vrg_source_busy_8$EN;
  // register m_vrg_source_busy_9
  reg m_vrg_source_busy_9;
  reg m_vrg_source_busy_9$D_IN;
  wire m_vrg_source_busy_9$EN;
  // register m_vrg_source_ip_0
  reg m_vrg_source_ip_0;
  wire m_vrg_source_ip_0$D_IN, m_vrg_source_ip_0$EN;
  // register m_vrg_source_ip_1
  reg m_vrg_source_ip_1;
  wire m_vrg_source_ip_1$D_IN, m_vrg_source_ip_1$EN;
  // register m_vrg_source_ip_10
  reg m_vrg_source_ip_10;
  wire m_vrg_source_ip_10$D_IN, m_vrg_source_ip_10$EN;
  // register m_vrg_source_ip_11
  reg m_vrg_source_ip_11;
  wire m_vrg_source_ip_11$D_IN, m_vrg_source_ip_11$EN;
  // register m_vrg_source_ip_12
  reg m_vrg_source_ip_12;
  wire m_vrg_source_ip_12$D_IN, m_vrg_source_ip_12$EN;
  // register m_vrg_source_ip_13
  reg m_vrg_source_ip_13;
  wire m_vrg_source_ip_13$D_IN, m_vrg_source_ip_13$EN;
  // register m_vrg_source_ip_14
  reg m_vrg_source_ip_14;
  wire m_vrg_source_ip_14$D_IN, m_vrg_source_ip_14$EN;
  // register m_vrg_source_ip_15
  reg m_vrg_source_ip_15;
  wire m_vrg_source_ip_15$D_IN, m_vrg_source_ip_15$EN;
  // register m_vrg_source_ip_16
  reg m_vrg_source_ip_16;
  wire m_vrg_source_ip_16$D_IN, m_vrg_source_ip_16$EN;
  // register m_vrg_source_ip_2
  reg m_vrg_source_ip_2;
  wire m_vrg_source_ip_2$D_IN, m_vrg_source_ip_2$EN;
  // register m_vrg_source_ip_3
  reg m_vrg_source_ip_3;
  wire m_vrg_source_ip_3$D_IN, m_vrg_source_ip_3$EN;
  // register m_vrg_source_ip_4
  reg m_vrg_source_ip_4;
  wire m_vrg_source_ip_4$D_IN, m_vrg_source_ip_4$EN;
  // register m_vrg_source_ip_5
  reg m_vrg_source_ip_5;
  wire m_vrg_source_ip_5$D_IN, m_vrg_source_ip_5$EN;
  // register m_vrg_source_ip_6
  reg m_vrg_source_ip_6;
  wire m_vrg_source_ip_6$D_IN, m_vrg_source_ip_6$EN;
  // register m_vrg_source_ip_7
  reg m_vrg_source_ip_7;
  wire m_vrg_source_ip_7$D_IN, m_vrg_source_ip_7$EN;
  // register m_vrg_source_ip_8
  reg m_vrg_source_ip_8;
  wire m_vrg_source_ip_8$D_IN, m_vrg_source_ip_8$EN;
  // register m_vrg_source_ip_9
  reg m_vrg_source_ip_9;
  wire m_vrg_source_ip_9$D_IN, m_vrg_source_ip_9$EN;
  // register m_vrg_source_prio_0
  reg [2 : 0] m_vrg_source_prio_0;
  wire [2 : 0] m_vrg_source_prio_0$D_IN;
  wire m_vrg_source_prio_0$EN;
  // register m_vrg_source_prio_1
  reg [2 : 0] m_vrg_source_prio_1;
  wire [2 : 0] m_vrg_source_prio_1$D_IN;
  wire m_vrg_source_prio_1$EN;
  // register m_vrg_source_prio_10
  reg [2 : 0] m_vrg_source_prio_10;
  wire [2 : 0] m_vrg_source_prio_10$D_IN;
  wire m_vrg_source_prio_10$EN;
  // register m_vrg_source_prio_11
  reg [2 : 0] m_vrg_source_prio_11;
  wire [2 : 0] m_vrg_source_prio_11$D_IN;
  wire m_vrg_source_prio_11$EN;
  // register m_vrg_source_prio_12
  reg [2 : 0] m_vrg_source_prio_12;
  wire [2 : 0] m_vrg_source_prio_12$D_IN;
  wire m_vrg_source_prio_12$EN;
  // register m_vrg_source_prio_13
  reg [2 : 0] m_vrg_source_prio_13;
  wire [2 : 0] m_vrg_source_prio_13$D_IN;
  wire m_vrg_source_prio_13$EN;
  // register m_vrg_source_prio_14
  reg [2 : 0] m_vrg_source_prio_14;
  wire [2 : 0] m_vrg_source_prio_14$D_IN;
  wire m_vrg_source_prio_14$EN;
  // register m_vrg_source_prio_15
  reg [2 : 0] m_vrg_source_prio_15;
  wire [2 : 0] m_vrg_source_prio_15$D_IN;
  wire m_vrg_source_prio_15$EN;
  // register m_vrg_source_prio_16
  reg [2 : 0] m_vrg_source_prio_16;
  wire [2 : 0] m_vrg_source_prio_16$D_IN;
  wire m_vrg_source_prio_16$EN;
  // register m_vrg_source_prio_2
  reg [2 : 0] m_vrg_source_prio_2;
  wire [2 : 0] m_vrg_source_prio_2$D_IN;
  wire m_vrg_source_prio_2$EN;
  // register m_vrg_source_prio_3
  reg [2 : 0] m_vrg_source_prio_3;
  wire [2 : 0] m_vrg_source_prio_3$D_IN;
  wire m_vrg_source_prio_3$EN;
  // register m_vrg_source_prio_4
  reg [2 : 0] m_vrg_source_prio_4;
  wire [2 : 0] m_vrg_source_prio_4$D_IN;
  wire m_vrg_source_prio_4$EN;
  // register m_vrg_source_prio_5
  reg [2 : 0] m_vrg_source_prio_5;
  wire [2 : 0] m_vrg_source_prio_5$D_IN;
  wire m_vrg_source_prio_5$EN;
  // register m_vrg_source_prio_6
  reg [2 : 0] m_vrg_source_prio_6;
  wire [2 : 0] m_vrg_source_prio_6$D_IN;
  wire m_vrg_source_prio_6$EN;
  // register m_vrg_source_prio_7
  reg [2 : 0] m_vrg_source_prio_7;
  wire [2 : 0] m_vrg_source_prio_7$D_IN;
  wire m_vrg_source_prio_7$EN;
  // register m_vrg_source_prio_8
  reg [2 : 0] m_vrg_source_prio_8;
  wire [2 : 0] m_vrg_source_prio_8$D_IN;
  wire m_vrg_source_prio_8$EN;
  // register m_vrg_source_prio_9
  reg [2 : 0] m_vrg_source_prio_9;
  wire [2 : 0] m_vrg_source_prio_9$D_IN;
  wire m_vrg_source_prio_9$EN;
  // register m_vrg_target_threshold_0
  reg [2 : 0] m_vrg_target_threshold_0;
  wire [2 : 0] m_vrg_target_threshold_0$D_IN;
  wire m_vrg_target_threshold_0$EN;
  // register m_vrg_target_threshold_1
  reg [2 : 0] m_vrg_target_threshold_1;
  wire [2 : 0] m_vrg_target_threshold_1$D_IN;
  wire m_vrg_target_threshold_1$EN;
  // register m_vvrg_ie_0_0
  reg m_vvrg_ie_0_0;
  wire m_vvrg_ie_0_0$D_IN, m_vvrg_ie_0_0$EN;
  // register m_vvrg_ie_0_1
  reg m_vvrg_ie_0_1;
  wire m_vvrg_ie_0_1$D_IN, m_vvrg_ie_0_1$EN;
  // register m_vvrg_ie_0_10
  reg m_vvrg_ie_0_10;
  wire m_vvrg_ie_0_10$D_IN, m_vvrg_ie_0_10$EN;
  // register m_vvrg_ie_0_11
  reg m_vvrg_ie_0_11;
  wire m_vvrg_ie_0_11$D_IN, m_vvrg_ie_0_11$EN;
  // register m_vvrg_ie_0_12
  reg m_vvrg_ie_0_12;
  wire m_vvrg_ie_0_12$D_IN, m_vvrg_ie_0_12$EN;
  // register m_vvrg_ie_0_13
  reg m_vvrg_ie_0_13;
  wire m_vvrg_ie_0_13$D_IN, m_vvrg_ie_0_13$EN;
  // register m_vvrg_ie_0_14
  reg m_vvrg_ie_0_14;
  wire m_vvrg_ie_0_14$D_IN, m_vvrg_ie_0_14$EN;
  // register m_vvrg_ie_0_15
  reg m_vvrg_ie_0_15;
  wire m_vvrg_ie_0_15$D_IN, m_vvrg_ie_0_15$EN;
  // register m_vvrg_ie_0_16
  reg m_vvrg_ie_0_16;
  wire m_vvrg_ie_0_16$D_IN, m_vvrg_ie_0_16$EN;
  // register m_vvrg_ie_0_2
  reg m_vvrg_ie_0_2;
  wire m_vvrg_ie_0_2$D_IN, m_vvrg_ie_0_2$EN;
  // register m_vvrg_ie_0_3
  reg m_vvrg_ie_0_3;
  wire m_vvrg_ie_0_3$D_IN, m_vvrg_ie_0_3$EN;
  // register m_vvrg_ie_0_4
  reg m_vvrg_ie_0_4;
  wire m_vvrg_ie_0_4$D_IN, m_vvrg_ie_0_4$EN;
  // register m_vvrg_ie_0_5
  reg m_vvrg_ie_0_5;
  wire m_vvrg_ie_0_5$D_IN, m_vvrg_ie_0_5$EN;
  // register m_vvrg_ie_0_6
  reg m_vvrg_ie_0_6;
  wire m_vvrg_ie_0_6$D_IN, m_vvrg_ie_0_6$EN;
  // register m_vvrg_ie_0_7
  reg m_vvrg_ie_0_7;
  wire m_vvrg_ie_0_7$D_IN, m_vvrg_ie_0_7$EN;
  // register m_vvrg_ie_0_8
  reg m_vvrg_ie_0_8;
  wire m_vvrg_ie_0_8$D_IN, m_vvrg_ie_0_8$EN;
  // register m_vvrg_ie_0_9
  reg m_vvrg_ie_0_9;
  wire m_vvrg_ie_0_9$D_IN, m_vvrg_ie_0_9$EN;
  // register m_vvrg_ie_1_0
  reg m_vvrg_ie_1_0;
  wire m_vvrg_ie_1_0$D_IN, m_vvrg_ie_1_0$EN;
  // register m_vvrg_ie_1_1
  reg m_vvrg_ie_1_1;
  wire m_vvrg_ie_1_1$D_IN, m_vvrg_ie_1_1$EN;
  // register m_vvrg_ie_1_10
  reg m_vvrg_ie_1_10;
  wire m_vvrg_ie_1_10$D_IN, m_vvrg_ie_1_10$EN;
  // register m_vvrg_ie_1_11
  reg m_vvrg_ie_1_11;
  wire m_vvrg_ie_1_11$D_IN, m_vvrg_ie_1_11$EN;
  // register m_vvrg_ie_1_12
  reg m_vvrg_ie_1_12;
  wire m_vvrg_ie_1_12$D_IN, m_vvrg_ie_1_12$EN;
  // register m_vvrg_ie_1_13
  reg m_vvrg_ie_1_13;
  wire m_vvrg_ie_1_13$D_IN, m_vvrg_ie_1_13$EN;
  // register m_vvrg_ie_1_14
  reg m_vvrg_ie_1_14;
  wire m_vvrg_ie_1_14$D_IN, m_vvrg_ie_1_14$EN;
  // register m_vvrg_ie_1_15
  reg m_vvrg_ie_1_15;
  wire m_vvrg_ie_1_15$D_IN, m_vvrg_ie_1_15$EN;
  // register m_vvrg_ie_1_16
  reg m_vvrg_ie_1_16;
  wire m_vvrg_ie_1_16$D_IN, m_vvrg_ie_1_16$EN;
  // register m_vvrg_ie_1_2
  reg m_vvrg_ie_1_2;
  wire m_vvrg_ie_1_2$D_IN, m_vvrg_ie_1_2$EN;
  // register m_vvrg_ie_1_3
  reg m_vvrg_ie_1_3;
  wire m_vvrg_ie_1_3$D_IN, m_vvrg_ie_1_3$EN;
  // register m_vvrg_ie_1_4
  reg m_vvrg_ie_1_4;
  wire m_vvrg_ie_1_4$D_IN, m_vvrg_ie_1_4$EN;
  // register m_vvrg_ie_1_5
  reg m_vvrg_ie_1_5;
  wire m_vvrg_ie_1_5$D_IN, m_vvrg_ie_1_5$EN;
  // register m_vvrg_ie_1_6
  reg m_vvrg_ie_1_6;
  wire m_vvrg_ie_1_6$D_IN, m_vvrg_ie_1_6$EN;
  // register m_vvrg_ie_1_7
  reg m_vvrg_ie_1_7;
  wire m_vvrg_ie_1_7$D_IN, m_vvrg_ie_1_7$EN;
  // register m_vvrg_ie_1_8
  reg m_vvrg_ie_1_8;
  wire m_vvrg_ie_1_8$D_IN, m_vvrg_ie_1_8$EN;
  // register m_vvrg_ie_1_9
  reg m_vvrg_ie_1_9;
  wire m_vvrg_ie_1_9$D_IN, m_vvrg_ie_1_9$EN;
  // ports of submodule m_f_reset_reqs
  wire m_f_reset_reqs$CLR,
       m_f_reset_reqs$DEQ,
       m_f_reset_reqs$EMPTY_N,
       m_f_reset_reqs$ENQ,
       m_f_reset_reqs$FULL_N;
  // ports of submodule m_f_reset_rsps
  wire m_f_reset_rsps$CLR,
       m_f_reset_rsps$DEQ,
       m_f_reset_rsps$EMPTY_N,
       m_f_reset_rsps$ENQ,
       m_f_reset_rsps$FULL_N;
  // ports of submodule m_slave_xactor_f_rd_addr
  wire [96 : 0] m_slave_xactor_f_rd_addr$D_IN, m_slave_xactor_f_rd_addr$D_OUT;
  wire m_slave_xactor_f_rd_addr$CLR,
       m_slave_xactor_f_rd_addr$DEQ,
       m_slave_xactor_f_rd_addr$EMPTY_N,
       m_slave_xactor_f_rd_addr$ENQ,
       m_slave_xactor_f_rd_addr$FULL_N;
  // ports of submodule m_slave_xactor_f_rd_data
  wire [70 : 0] m_slave_xactor_f_rd_data$D_IN, m_slave_xactor_f_rd_data$D_OUT;
  wire m_slave_xactor_f_rd_data$CLR,
       m_slave_xactor_f_rd_data$DEQ,
       m_slave_xactor_f_rd_data$EMPTY_N,
       m_slave_xactor_f_rd_data$ENQ,
       m_slave_xactor_f_rd_data$FULL_N;
  // ports of submodule m_slave_xactor_f_wr_addr
  wire [96 : 0] m_slave_xactor_f_wr_addr$D_IN, m_slave_xactor_f_wr_addr$D_OUT;
  wire m_slave_xactor_f_wr_addr$CLR,
       m_slave_xactor_f_wr_addr$DEQ,
       m_slave_xactor_f_wr_addr$EMPTY_N,
       m_slave_xactor_f_wr_addr$ENQ,
       m_slave_xactor_f_wr_addr$FULL_N;
  // ports of submodule m_slave_xactor_f_wr_data
  wire [72 : 0] m_slave_xactor_f_wr_data$D_IN, m_slave_xactor_f_wr_data$D_OUT;
  wire m_slave_xactor_f_wr_data$CLR,
       m_slave_xactor_f_wr_data$DEQ,
       m_slave_xactor_f_wr_data$EMPTY_N,
       m_slave_xactor_f_wr_data$ENQ,
       m_slave_xactor_f_wr_data$FULL_N;
  // ports of submodule m_slave_xactor_f_wr_resp
  wire [5 : 0] m_slave_xactor_f_wr_resp$D_IN, m_slave_xactor_f_wr_resp$D_OUT;
  wire m_slave_xactor_f_wr_resp$CLR,
       m_slave_xactor_f_wr_resp$DEQ,
       m_slave_xactor_f_wr_resp$EMPTY_N,
       m_slave_xactor_f_wr_resp$ENQ,
       m_slave_xactor_f_wr_resp$FULL_N;
  // rule scheduling signals
  wire CAN_FIRE_RL_m_rl_process_rd_req,
       CAN_FIRE_RL_m_rl_process_wr_req,
       CAN_FIRE_RL_m_rl_reset,
       CAN_FIRE_axi4_slave_m_arvalid,
       CAN_FIRE_axi4_slave_m_awvalid,
       CAN_FIRE_axi4_slave_m_bready,
       CAN_FIRE_axi4_slave_m_rready,
       CAN_FIRE_axi4_slave_m_wvalid,
       CAN_FIRE_server_reset_request_put,
       CAN_FIRE_server_reset_response_get,
       CAN_FIRE_set_addr_map,
       CAN_FIRE_set_verbosity,
       CAN_FIRE_show_PLIC_state,
       CAN_FIRE_v_sources_0_m_interrupt_req,
       CAN_FIRE_v_sources_10_m_interrupt_req,
       CAN_FIRE_v_sources_11_m_interrupt_req,
       CAN_FIRE_v_sources_12_m_interrupt_req,
       CAN_FIRE_v_sources_13_m_interrupt_req,
       CAN_FIRE_v_sources_14_m_interrupt_req,
       CAN_FIRE_v_sources_15_m_interrupt_req,
       CAN_FIRE_v_sources_1_m_interrupt_req,
       CAN_FIRE_v_sources_2_m_interrupt_req,
       CAN_FIRE_v_sources_3_m_interrupt_req,
       CAN_FIRE_v_sources_4_m_interrupt_req,
       CAN_FIRE_v_sources_5_m_interrupt_req,
       CAN_FIRE_v_sources_6_m_interrupt_req,
       CAN_FIRE_v_sources_7_m_interrupt_req,
       CAN_FIRE_v_sources_8_m_interrupt_req,
       CAN_FIRE_v_sources_9_m_interrupt_req,
       WILL_FIRE_RL_m_rl_process_rd_req,
       WILL_FIRE_RL_m_rl_process_wr_req,
       WILL_FIRE_RL_m_rl_reset,
       WILL_FIRE_axi4_slave_m_arvalid,
       WILL_FIRE_axi4_slave_m_awvalid,
       WILL_FIRE_axi4_slave_m_bready,
       WILL_FIRE_axi4_slave_m_rready,
       WILL_FIRE_axi4_slave_m_wvalid,
       WILL_FIRE_server_reset_request_put,
       WILL_FIRE_server_reset_response_get,
       WILL_FIRE_set_addr_map,
       WILL_FIRE_set_verbosity,
       WILL_FIRE_show_PLIC_state,
       WILL_FIRE_v_sources_0_m_interrupt_req,
       WILL_FIRE_v_sources_10_m_interrupt_req,
       WILL_FIRE_v_sources_11_m_interrupt_req,
       WILL_FIRE_v_sources_12_m_interrupt_req,
       WILL_FIRE_v_sources_13_m_interrupt_req,
       WILL_FIRE_v_sources_14_m_interrupt_req,
       WILL_FIRE_v_sources_15_m_interrupt_req,
       WILL_FIRE_v_sources_1_m_interrupt_req,
       WILL_FIRE_v_sources_2_m_interrupt_req,
       WILL_FIRE_v_sources_3_m_interrupt_req,
       WILL_FIRE_v_sources_4_m_interrupt_req,
       WILL_FIRE_v_sources_5_m_interrupt_req,
       WILL_FIRE_v_sources_6_m_interrupt_req,
       WILL_FIRE_v_sources_7_m_interrupt_req,
       WILL_FIRE_v_sources_8_m_interrupt_req,
       WILL_FIRE_v_sources_9_m_interrupt_req;
  // inputs to muxes for submodule ports
  wire MUX_m_vrg_source_busy_0$write_1__SEL_1,
       MUX_m_vrg_source_busy_0$write_1__SEL_2,
       MUX_m_vrg_source_busy_1$write_1__SEL_1,
       MUX_m_vrg_source_busy_1$write_1__SEL_2,
       MUX_m_vrg_source_busy_10$write_1__SEL_1,
       MUX_m_vrg_source_busy_10$write_1__SEL_2,
       MUX_m_vrg_source_busy_11$write_1__SEL_1,
       MUX_m_vrg_source_busy_11$write_1__SEL_2,
       MUX_m_vrg_source_busy_12$write_1__SEL_1,
       MUX_m_vrg_source_busy_12$write_1__SEL_2,
       MUX_m_vrg_source_busy_13$write_1__SEL_1,
       MUX_m_vrg_source_busy_13$write_1__SEL_2,
       MUX_m_vrg_source_busy_14$write_1__SEL_1,
       MUX_m_vrg_source_busy_14$write_1__SEL_2,
       MUX_m_vrg_source_busy_15$write_1__SEL_1,
       MUX_m_vrg_source_busy_15$write_1__SEL_2,
       MUX_m_vrg_source_busy_16$write_1__SEL_1,
       MUX_m_vrg_source_busy_16$write_1__SEL_2,
       MUX_m_vrg_source_busy_2$write_1__SEL_1,
       MUX_m_vrg_source_busy_2$write_1__SEL_2,
       MUX_m_vrg_source_busy_3$write_1__SEL_1,
       MUX_m_vrg_source_busy_3$write_1__SEL_2,
       MUX_m_vrg_source_busy_4$write_1__SEL_1,
       MUX_m_vrg_source_busy_4$write_1__SEL_2,
       MUX_m_vrg_source_busy_5$write_1__SEL_1,
       MUX_m_vrg_source_busy_5$write_1__SEL_2,
       MUX_m_vrg_source_busy_6$write_1__SEL_1,
       MUX_m_vrg_source_busy_6$write_1__SEL_2,
       MUX_m_vrg_source_busy_7$write_1__SEL_1,
       MUX_m_vrg_source_busy_7$write_1__SEL_2,
       MUX_m_vrg_source_busy_8$write_1__SEL_1,
       MUX_m_vrg_source_busy_8$write_1__SEL_2,
       MUX_m_vrg_source_busy_9$write_1__SEL_1,
       MUX_m_vrg_source_busy_9$write_1__SEL_2,
       MUX_m_vrg_source_prio_0$write_1__SEL_1,
       MUX_m_vrg_source_prio_1$write_1__SEL_1,
       MUX_m_vrg_source_prio_10$write_1__SEL_1,
       MUX_m_vrg_source_prio_11$write_1__SEL_1,
       MUX_m_vrg_source_prio_12$write_1__SEL_1,
       MUX_m_vrg_source_prio_13$write_1__SEL_1,
       MUX_m_vrg_source_prio_14$write_1__SEL_1,
       MUX_m_vrg_source_prio_15$write_1__SEL_1,
       MUX_m_vrg_source_prio_16$write_1__SEL_1,
       MUX_m_vrg_source_prio_2$write_1__SEL_1,
       MUX_m_vrg_source_prio_3$write_1__SEL_1,
       MUX_m_vrg_source_prio_4$write_1__SEL_1,
       MUX_m_vrg_source_prio_5$write_1__SEL_1,
       MUX_m_vrg_source_prio_6$write_1__SEL_1,
       MUX_m_vrg_source_prio_7$write_1__SEL_1,
       MUX_m_vrg_source_prio_8$write_1__SEL_1,
       MUX_m_vrg_source_prio_9$write_1__SEL_1,
       MUX_m_vrg_target_threshold_0$write_1__SEL_1,
       MUX_m_vrg_target_threshold_1$write_1__SEL_1,
       MUX_m_vvrg_ie_0_0$write_1__SEL_1,
       MUX_m_vvrg_ie_0_0$write_1__VAL_1,
       MUX_m_vvrg_ie_0_1$write_1__SEL_1,
       MUX_m_vvrg_ie_0_1$write_1__VAL_1,
       MUX_m_vvrg_ie_0_10$write_1__SEL_1,
       MUX_m_vvrg_ie_0_10$write_1__VAL_1,
       MUX_m_vvrg_ie_0_11$write_1__SEL_1,
       MUX_m_vvrg_ie_0_11$write_1__VAL_1,
       MUX_m_vvrg_ie_0_12$write_1__SEL_1,
       MUX_m_vvrg_ie_0_12$write_1__VAL_1,
       MUX_m_vvrg_ie_0_13$write_1__SEL_1,
       MUX_m_vvrg_ie_0_13$write_1__VAL_1,
       MUX_m_vvrg_ie_0_14$write_1__SEL_1,
       MUX_m_vvrg_ie_0_14$write_1__VAL_1,
       MUX_m_vvrg_ie_0_15$write_1__SEL_1,
       MUX_m_vvrg_ie_0_15$write_1__VAL_1,
       MUX_m_vvrg_ie_0_16$write_1__SEL_1,
       MUX_m_vvrg_ie_0_16$write_1__VAL_1,
       MUX_m_vvrg_ie_0_2$write_1__SEL_1,
       MUX_m_vvrg_ie_0_2$write_1__VAL_1,
       MUX_m_vvrg_ie_0_3$write_1__SEL_1,
       MUX_m_vvrg_ie_0_3$write_1__VAL_1,
       MUX_m_vvrg_ie_0_4$write_1__SEL_1,
       MUX_m_vvrg_ie_0_4$write_1__VAL_1,
       MUX_m_vvrg_ie_0_5$write_1__SEL_1,
       MUX_m_vvrg_ie_0_5$write_1__VAL_1,
       MUX_m_vvrg_ie_0_6$write_1__SEL_1,
       MUX_m_vvrg_ie_0_6$write_1__VAL_1,
       MUX_m_vvrg_ie_0_7$write_1__SEL_1,
       MUX_m_vvrg_ie_0_7$write_1__VAL_1,
       MUX_m_vvrg_ie_0_8$write_1__SEL_1,
       MUX_m_vvrg_ie_0_8$write_1__VAL_1,
       MUX_m_vvrg_ie_0_9$write_1__SEL_1,
       MUX_m_vvrg_ie_0_9$write_1__VAL_1,
       MUX_m_vvrg_ie_1_0$write_1__SEL_1,
       MUX_m_vvrg_ie_1_0$write_1__VAL_1,
       MUX_m_vvrg_ie_1_1$write_1__SEL_1,
       MUX_m_vvrg_ie_1_1$write_1__VAL_1,
       MUX_m_vvrg_ie_1_10$write_1__SEL_1,
       MUX_m_vvrg_ie_1_10$write_1__VAL_1,
       MUX_m_vvrg_ie_1_11$write_1__SEL_1,
       MUX_m_vvrg_ie_1_11$write_1__VAL_1,
       MUX_m_vvrg_ie_1_12$write_1__SEL_1,
       MUX_m_vvrg_ie_1_12$write_1__VAL_1,
       MUX_m_vvrg_ie_1_13$write_1__SEL_1,
       MUX_m_vvrg_ie_1_13$write_1__VAL_1,
       MUX_m_vvrg_ie_1_14$write_1__SEL_1,
       MUX_m_vvrg_ie_1_14$write_1__VAL_1,
       MUX_m_vvrg_ie_1_15$write_1__SEL_1,
       MUX_m_vvrg_ie_1_15$write_1__VAL_1,
       MUX_m_vvrg_ie_1_16$write_1__SEL_1,
       MUX_m_vvrg_ie_1_16$write_1__VAL_1,
       MUX_m_vvrg_ie_1_2$write_1__SEL_1,
       MUX_m_vvrg_ie_1_2$write_1__VAL_1,
       MUX_m_vvrg_ie_1_3$write_1__SEL_1,
       MUX_m_vvrg_ie_1_3$write_1__VAL_1,
       MUX_m_vvrg_ie_1_4$write_1__SEL_1,
       MUX_m_vvrg_ie_1_4$write_1__VAL_1,
       MUX_m_vvrg_ie_1_5$write_1__SEL_1,
       MUX_m_vvrg_ie_1_5$write_1__VAL_1,
       MUX_m_vvrg_ie_1_6$write_1__SEL_1,
       MUX_m_vvrg_ie_1_6$write_1__VAL_1,
       MUX_m_vvrg_ie_1_7$write_1__SEL_1,
       MUX_m_vvrg_ie_1_7$write_1__VAL_1,
       MUX_m_vvrg_ie_1_8$write_1__SEL_1,
       MUX_m_vvrg_ie_1_8$write_1__VAL_1,
       MUX_m_vvrg_ie_1_9$write_1__SEL_1,
       MUX_m_vvrg_ie_1_9$write_1__VAL_1;
  // declarations used by system tasks
  // synopsys translate_off
  reg [31 : 0] v__h86248;
  reg [31 : 0] v__h86443;
  reg [31 : 0] v__h86638;
  reg [31 : 0] v__h86833;
  reg [31 : 0] v__h87028;
  reg [31 : 0] v__h87223;
  reg [31 : 0] v__h87418;
  reg [31 : 0] v__h87613;
  reg [31 : 0] v__h87808;
  reg [31 : 0] v__h88003;
  reg [31 : 0] v__h88198;
  reg [31 : 0] v__h88393;
  reg [31 : 0] v__h88588;
  reg [31 : 0] v__h88783;
  reg [31 : 0] v__h88978;
  reg [31 : 0] v__h89173;
  reg [31 : 0] v__h5962;
  reg [31 : 0] v__h13331;
  reg [31 : 0] v__h13514;
  reg [31 : 0] v__h13730;
  reg [31 : 0] v__h13976;
  reg [31 : 0] v__h18445;
  reg [31 : 0] v__h24057;
  reg [31 : 0] v__h26355;
  reg [31 : 0] v__h26568;
  reg [31 : 0] v__h26773;
  reg [31 : 0] v__h27053;
  reg [31 : 0] v__h27284;
  reg [31 : 0] v__h28359;
  reg [31 : 0] v__h28531;
  reg [31 : 0] v__h76647;
  reg [31 : 0] v__h76947;
  reg [31 : 0] v__h77579;
  reg [31 : 0] v__h77673;
  reg [31 : 0] v__h77844;
  reg [31 : 0] v__h78064;
  reg [31 : 0] v__h85245;
  reg [31 : 0] v__h85351;
  reg [31 : 0] v__h85478;
  reg [31 : 0] v__h5956;
  reg [31 : 0] v__h13325;
  reg [31 : 0] v__h13508;
  reg [31 : 0] v__h13724;
  reg [31 : 0] v__h13970;
  reg [31 : 0] v__h18439;
  reg [31 : 0] v__h24051;
  reg [31 : 0] v__h26349;
  reg [31 : 0] v__h26562;
  reg [31 : 0] v__h26767;
  reg [31 : 0] v__h27047;
  reg [31 : 0] v__h27278;
  reg [31 : 0] v__h28353;
  reg [31 : 0] v__h28525;
  reg [31 : 0] v__h76641;
  reg [31 : 0] v__h76941;
  reg [31 : 0] v__h77573;
  reg [31 : 0] v__h77667;
  reg [31 : 0] v__h77838;
  reg [31 : 0] v__h78058;
  reg [31 : 0] v__h85239;
  reg [31 : 0] v__h85345;
  reg [31 : 0] v__h85472;
  reg [31 : 0] v__h86242;
  reg [31 : 0] v__h86437;
  reg [31 : 0] v__h86632;
  reg [31 : 0] v__h86827;
  reg [31 : 0] v__h87022;
  reg [31 : 0] v__h87217;
  reg [31 : 0] v__h87412;
  reg [31 : 0] v__h87607;
  reg [31 : 0] v__h87802;
  reg [31 : 0] v__h87997;
  reg [31 : 0] v__h88192;
  reg [31 : 0] v__h88387;
  reg [31 : 0] v__h88582;
  reg [31 : 0] v__h88777;
  reg [31 : 0] v__h88972;
  reg [31 : 0] v__h89167;
  // synopsys translate_on
  // remaining internal signals
  reg [63 : 0] y_avValue_fst__h26466;
  reg [2 : 0] x__h13769, x__h24096;
  reg [1 : 0] v__h76713, y_avValue_snd__h26467;
  reg CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q1,
      CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q10,
      CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q11,
      CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q12,
      CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q13,
      CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q14,
      CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q15,
      CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q16,
      CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q17,
      CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q18,
      CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q19,
      CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q2,
      CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q20,
      CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q21,
      CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q22,
      CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q23,
      CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q24,
      CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q25,
      CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q26,
      CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q27,
      CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q28,
      CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q29,
      CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q3,
      CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q30,
      CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q31,
      CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q32,
      CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q4,
      CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q5,
      CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q6,
      CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q7,
      CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q8,
      CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q9,
      CASE_addr_offset3465_BITS_16_TO_12_0_m_vvrg_ie_ETC__q33,
      CASE_addr_offset3465_BITS_16_TO_12_0_m_vvrg_ie_ETC__q34,
      CASE_addr_offset3465_BITS_16_TO_12_0_m_vvrg_ie_ETC__q35,
      CASE_addr_offset3465_BITS_16_TO_12_0_m_vvrg_ie_ETC__q36,
      CASE_addr_offset3465_BITS_16_TO_12_0_m_vvrg_ie_ETC__q37,
      CASE_addr_offset3465_BITS_16_TO_12_0_m_vvrg_ie_ETC__q38,
      CASE_addr_offset3465_BITS_16_TO_12_0_m_vvrg_ie_ETC__q39,
      CASE_addr_offset3465_BITS_16_TO_12_0_m_vvrg_ie_ETC__q40,
      CASE_addr_offset3465_BITS_16_TO_12_0_m_vvrg_ie_ETC__q41,
      CASE_addr_offset3465_BITS_16_TO_12_0_m_vvrg_ie_ETC__q42,
      CASE_addr_offset3465_BITS_16_TO_12_0_m_vvrg_ie_ETC__q43,
      CASE_addr_offset3465_BITS_16_TO_12_0_m_vvrg_ie_ETC__q44,
      CASE_addr_offset3465_BITS_16_TO_12_0_m_vvrg_ie_ETC__q45,
      CASE_addr_offset3465_BITS_16_TO_12_0_m_vvrg_ie_ETC__q46,
      CASE_addr_offset3465_BITS_16_TO_12_0_m_vvrg_ie_ETC__q47,
      CASE_addr_offset3465_BITS_16_TO_12_0_m_vvrg_ie_ETC__q48,
      SEL_ARR_SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_ETC___d2878,
      SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d102,
      SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d107,
      SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d111,
      SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d116,
      SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d120,
      SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d125,
      SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d129,
      SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d134,
      SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d138,
      SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d143,
      SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d147,
      SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d152,
      SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d156,
      SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d161,
      SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d165,
      SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d170,
      SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d174,
      SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d179,
      SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d183,
      SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d188,
      SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d192,
      SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d197,
      SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d201,
      SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d206,
      SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d210,
      SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d215,
      SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d219,
      SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d224,
      SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d228,
      SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d233,
      SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d235,
      SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d98,
      SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d271,
      SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d2875,
      SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d296,
      SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d304,
      SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d311,
      SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d319,
      SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d326,
      SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d334,
      SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d341,
      SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d349,
      SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d356,
      SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d364,
      SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d371,
      SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d379,
      SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d386,
      SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d394,
      SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d401,
      SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d409,
      SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d416,
      SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d424,
      SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d431,
      SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d439,
      SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d446,
      SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d454,
      SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d461,
      SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d469,
      SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d476,
      SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d484,
      SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d491,
      SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d499,
      SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d506,
      SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d514,
      SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d519,
      SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d2876,
      SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d290,
      SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d297,
      SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d305,
      SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d312,
      SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d320,
      SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d327,
      SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d335,
      SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d342,
      SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d350,
      SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d357,
      SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d365,
      SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d372,
      SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d380,
      SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d387,
      SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d395,
      SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d402,
      SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d410,
      SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d417,
      SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d425,
      SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d432,
      SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d440,
      SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d447,
      SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d455,
      SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d462,
      SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d470,
      SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d477,
      SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d485,
      SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d492,
      SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d500,
      SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d507,
      SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d515,
      SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d520;
  wire [63 : 0] addr_offset__h13465,
		addr_offset__h27245,
		rdata___1__h26714,
		rdata__h26520,
		v__h13689,
		v__h13934,
		v__h18403,
		v__h24016,
		v__h24251,
		v__h25556,
		x__h26677,
		y_avValue_fst__h26433,
		y_avValue_fst__h26445,
		y_avValue_fst__h26461,
		y_avValue_fst__h26477,
		y_avValue_fst__h26482,
		y_avValue_fst__h26493,
		y_avValue_fst__h26498,
		y_avValue_fst__h26512;
  wire [31 : 0] v_ie__h18406,
		v_ip__h13937,
		wdata32__h27246,
		x__h23928,
		x__h76716;
  wire [9 : 0] source_id__h15937,
	       source_id__h16044,
	       source_id__h16117,
	       source_id__h16190,
	       source_id__h16263,
	       source_id__h16336,
	       source_id__h16409,
	       source_id__h16482,
	       source_id__h16555,
	       source_id__h16628,
	       source_id__h16701,
	       source_id__h16774,
	       source_id__h16847,
	       source_id__h16920,
	       source_id__h16993,
	       source_id__h17066,
	       source_id__h17139,
	       source_id__h17212,
	       source_id__h17285,
	       source_id__h17358,
	       source_id__h17431,
	       source_id__h17504,
	       source_id__h17577,
	       source_id__h17650,
	       source_id__h17723,
	       source_id__h17796,
	       source_id__h17869,
	       source_id__h17942,
	       source_id__h18015,
	       source_id__h18088,
	       source_id__h18161,
	       source_id__h20405,
	       source_id__h20581,
	       source_id__h20689,
	       source_id__h20797,
	       source_id__h20905,
	       source_id__h21013,
	       source_id__h21121,
	       source_id__h21229,
	       source_id__h21337,
	       source_id__h21445,
	       source_id__h21553,
	       source_id__h21661,
	       source_id__h21769,
	       source_id__h21877,
	       source_id__h21985,
	       source_id__h22093,
	       source_id__h22201,
	       source_id__h22309,
	       source_id__h22417,
	       source_id__h22525,
	       source_id__h22633,
	       source_id__h22741,
	       source_id__h22849,
	       source_id__h22957,
	       source_id__h23065,
	       source_id__h23173,
	       source_id__h23281,
	       source_id__h23389,
	       source_id__h23497,
	       source_id__h23605,
	       source_id__h23713,
	       source_id__h30233,
	       source_id__h31729,
	       source_id__h33225,
	       source_id__h34721,
	       source_id__h36217,
	       source_id__h37713,
	       source_id__h39209,
	       source_id__h40705,
	       source_id__h42201,
	       source_id__h43697,
	       source_id__h45193,
	       source_id__h46689,
	       source_id__h48185,
	       source_id__h49681,
	       source_id__h51177,
	       source_id__h52673,
	       source_id__h54169,
	       source_id__h55665,
	       source_id__h57161,
	       source_id__h58657,
	       source_id__h60153,
	       source_id__h61649,
	       source_id__h63145,
	       source_id__h64641,
	       source_id__h66137,
	       source_id__h67633,
	       source_id__h69129,
	       source_id__h70625,
	       source_id__h72121,
	       source_id__h73617,
	       source_id__h75113,
	       source_id_base__h13893,
	       source_id_base__h28620;
  wire [4 : 0] IF_m_vrg_source_ip_11_read__1_AND_NOT_m_vrg_so_ETC___d3078,
	       IF_m_vrg_source_ip_11_read__1_AND_NOT_m_vrg_so_ETC___d3172,
	       IF_m_vrg_source_ip_11_read__1_AND_NOT_m_vrg_so_ETC___d667,
	       IF_m_vrg_source_ip_13_read__3_AND_NOT_m_vrg_so_ETC___d3080,
	       IF_m_vrg_source_ip_13_read__3_AND_NOT_m_vrg_so_ETC___d3174,
	       IF_m_vrg_source_ip_13_read__3_AND_NOT_m_vrg_so_ETC___d669,
	       IF_m_vrg_source_ip_15_read__5_AND_NOT_m_vrg_so_ETC___d3082,
	       IF_m_vrg_source_ip_15_read__5_AND_NOT_m_vrg_so_ETC___d3176,
	       IF_m_vrg_source_ip_15_read__5_AND_NOT_m_vrg_so_ETC___d671,
	       IF_m_vrg_source_ip_3_read__3_AND_NOT_m_vrg_sou_ETC___d3070,
	       IF_m_vrg_source_ip_3_read__3_AND_NOT_m_vrg_sou_ETC___d3164,
	       IF_m_vrg_source_ip_3_read__3_AND_NOT_m_vrg_sou_ETC___d659,
	       IF_m_vrg_source_ip_5_read__5_AND_NOT_m_vrg_sou_ETC___d3072,
	       IF_m_vrg_source_ip_5_read__5_AND_NOT_m_vrg_sou_ETC___d3166,
	       IF_m_vrg_source_ip_5_read__5_AND_NOT_m_vrg_sou_ETC___d661,
	       IF_m_vrg_source_ip_7_read__7_AND_NOT_m_vrg_sou_ETC___d3074,
	       IF_m_vrg_source_ip_7_read__7_AND_NOT_m_vrg_sou_ETC___d3168,
	       IF_m_vrg_source_ip_7_read__7_AND_NOT_m_vrg_sou_ETC___d663,
	       IF_m_vrg_source_ip_9_read__9_AND_NOT_m_vrg_sou_ETC___d3076,
	       IF_m_vrg_source_ip_9_read__9_AND_NOT_m_vrg_sou_ETC___d3170,
	       IF_m_vrg_source_ip_9_read__9_AND_NOT_m_vrg_sou_ETC___d665,
	       b__h81741,
	       b__h83895,
	       max_id__h24210;
  wire [2 : 0] IF_m_vrg_source_ip_10_read__0_AND_NOT_m_vrg_so_ETC___d3037,
	       IF_m_vrg_source_ip_10_read__0_AND_NOT_m_vrg_so_ETC___d3131,
	       IF_m_vrg_source_ip_10_read__0_AND_NOT_m_vrg_so_ETC___d615,
	       IF_m_vrg_source_ip_11_read__1_AND_NOT_m_vrg_so_ETC___d3042,
	       IF_m_vrg_source_ip_11_read__1_AND_NOT_m_vrg_so_ETC___d3136,
	       IF_m_vrg_source_ip_11_read__1_AND_NOT_m_vrg_so_ETC___d622,
	       IF_m_vrg_source_ip_12_read__2_AND_NOT_m_vrg_so_ETC___d3047,
	       IF_m_vrg_source_ip_12_read__2_AND_NOT_m_vrg_so_ETC___d3141,
	       IF_m_vrg_source_ip_12_read__2_AND_NOT_m_vrg_so_ETC___d629,
	       IF_m_vrg_source_ip_13_read__3_AND_NOT_m_vrg_so_ETC___d3052,
	       IF_m_vrg_source_ip_13_read__3_AND_NOT_m_vrg_so_ETC___d3146,
	       IF_m_vrg_source_ip_13_read__3_AND_NOT_m_vrg_so_ETC___d636,
	       IF_m_vrg_source_ip_14_read__4_AND_NOT_m_vrg_so_ETC___d3057,
	       IF_m_vrg_source_ip_14_read__4_AND_NOT_m_vrg_so_ETC___d3151,
	       IF_m_vrg_source_ip_14_read__4_AND_NOT_m_vrg_so_ETC___d643,
	       IF_m_vrg_source_ip_15_read__5_AND_NOT_m_vrg_so_ETC___d3062,
	       IF_m_vrg_source_ip_15_read__5_AND_NOT_m_vrg_so_ETC___d3156,
	       IF_m_vrg_source_ip_1_read__1_AND_NOT_m_vrg_sou_ETC___d2992,
	       IF_m_vrg_source_ip_1_read__1_AND_NOT_m_vrg_sou_ETC___d3086,
	       IF_m_vrg_source_ip_1_read__1_AND_NOT_m_vrg_sou_ETC___d552,
	       IF_m_vrg_source_ip_2_read__2_AND_NOT_m_vrg_sou_ETC___d2997,
	       IF_m_vrg_source_ip_2_read__2_AND_NOT_m_vrg_sou_ETC___d3091,
	       IF_m_vrg_source_ip_2_read__2_AND_NOT_m_vrg_sou_ETC___d559,
	       IF_m_vrg_source_ip_3_read__3_AND_NOT_m_vrg_sou_ETC___d3002,
	       IF_m_vrg_source_ip_3_read__3_AND_NOT_m_vrg_sou_ETC___d3096,
	       IF_m_vrg_source_ip_3_read__3_AND_NOT_m_vrg_sou_ETC___d566,
	       IF_m_vrg_source_ip_4_read__4_AND_NOT_m_vrg_sou_ETC___d3007,
	       IF_m_vrg_source_ip_4_read__4_AND_NOT_m_vrg_sou_ETC___d3101,
	       IF_m_vrg_source_ip_4_read__4_AND_NOT_m_vrg_sou_ETC___d573,
	       IF_m_vrg_source_ip_5_read__5_AND_NOT_m_vrg_sou_ETC___d3012,
	       IF_m_vrg_source_ip_5_read__5_AND_NOT_m_vrg_sou_ETC___d3106,
	       IF_m_vrg_source_ip_5_read__5_AND_NOT_m_vrg_sou_ETC___d580,
	       IF_m_vrg_source_ip_6_read__6_AND_NOT_m_vrg_sou_ETC___d3017,
	       IF_m_vrg_source_ip_6_read__6_AND_NOT_m_vrg_sou_ETC___d3111,
	       IF_m_vrg_source_ip_6_read__6_AND_NOT_m_vrg_sou_ETC___d587,
	       IF_m_vrg_source_ip_7_read__7_AND_NOT_m_vrg_sou_ETC___d3022,
	       IF_m_vrg_source_ip_7_read__7_AND_NOT_m_vrg_sou_ETC___d3116,
	       IF_m_vrg_source_ip_7_read__7_AND_NOT_m_vrg_sou_ETC___d594,
	       IF_m_vrg_source_ip_8_read__8_AND_NOT_m_vrg_sou_ETC___d3027,
	       IF_m_vrg_source_ip_8_read__8_AND_NOT_m_vrg_sou_ETC___d3121,
	       IF_m_vrg_source_ip_8_read__8_AND_NOT_m_vrg_sou_ETC___d601,
	       IF_m_vrg_source_ip_9_read__9_AND_NOT_m_vrg_sou_ETC___d3032,
	       IF_m_vrg_source_ip_9_read__9_AND_NOT_m_vrg_sou_ETC___d3126,
	       IF_m_vrg_source_ip_9_read__9_AND_NOT_m_vrg_sou_ETC___d608,
	       a__h81740,
	       a__h83894;
  wire [1 : 0] rresp__h26521,
	       v__h27250,
	       v__h27435,
	       v__h27448,
	       v__h28425,
	       v__h28444,
	       v__h28597,
	       v__h28616,
	       v__h76750,
	       y_avValue_snd__h26446,
	       y_avValue_snd__h26462,
	       y_avValue_snd__h26478,
	       y_avValue_snd__h26483,
	       y_avValue_snd__h26494,
	       y_avValue_snd__h26499,
	       y_avValue_snd__h26513;
  wire IF_m_slave_xactor_f_rd_addr_first__9_BITS_92_T_ETC___d748,
       IF_m_slave_xactor_f_rd_addr_first__9_BITS_92_T_ETC___d750,
       IF_m_slave_xactor_f_wr_addr_first__94_BITS_92__ETC___d2874,
       IF_m_slave_xactor_f_wr_addr_first__94_BITS_92__ETC___d2950,
       IF_m_slave_xactor_f_wr_addr_first__94_BITS_92__ETC___d2952,
       NOT_m_cfg_verbosity_read_ULE_1_5___d16,
       NOT_m_slave_xactor_f_rd_addr_first__9_BITS_92__ETC___d248,
       NOT_m_slave_xactor_f_rd_addr_first__9_BITS_92__ETC___d538,
       NOT_m_slave_xactor_f_rd_addr_first__9_BITS_92__ETC___d695,
       NOT_m_slave_xactor_f_rd_addr_first__9_BITS_92__ETC___d733,
       NOT_m_slave_xactor_f_rd_addr_first__9_BITS_92__ETC___d74,
       NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1017,
       NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1078,
       NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1139,
       NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1200,
       NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1261,
       NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1322,
       NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1383,
       NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1444,
       NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1505,
       NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1566,
       NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1627,
       NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1688,
       NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1749,
       NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1810,
       NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1871,
       NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1932,
       NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1993,
       NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2054,
       NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2115,
       NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2176,
       NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2237,
       NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2298,
       NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2359,
       NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2420,
       NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2481,
       NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2542,
       NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2603,
       NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2664,
       NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2725,
       NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2786,
       NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2844,
       NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2857,
       NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2868,
       NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2884,
       NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2923,
       NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2935,
       NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d826,
       NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d880,
       NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d892,
       NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d956,
       NOT_m_vrg_source_busy_10_983_284_AND_NOT_m_cfg_ETC___d3288,
       NOT_m_vrg_source_busy_11_984_292_AND_NOT_m_cfg_ETC___d3296,
       NOT_m_vrg_source_busy_12_985_300_AND_NOT_m_cfg_ETC___d3304,
       NOT_m_vrg_source_busy_13_986_308_AND_NOT_m_cfg_ETC___d3312,
       NOT_m_vrg_source_busy_14_987_316_AND_NOT_m_cfg_ETC___d3320,
       NOT_m_vrg_source_busy_15_988_324_AND_NOT_m_cfg_ETC___d3328,
       NOT_m_vrg_source_busy_16_989_332_AND_NOT_m_cfg_ETC___d3336,
       NOT_m_vrg_source_busy_1_974_213_AND_NOT_m_cfg__ETC___d3217,
       NOT_m_vrg_source_busy_2_975_220_AND_NOT_m_cfg__ETC___d3224,
       NOT_m_vrg_source_busy_3_976_228_AND_NOT_m_cfg__ETC___d3232,
       NOT_m_vrg_source_busy_4_977_236_AND_NOT_m_cfg__ETC___d3240,
       NOT_m_vrg_source_busy_5_978_244_AND_NOT_m_cfg__ETC___d3248,
       NOT_m_vrg_source_busy_6_979_252_AND_NOT_m_cfg__ETC___d3256,
       NOT_m_vrg_source_busy_7_980_260_AND_NOT_m_cfg__ETC___d3264,
       NOT_m_vrg_source_busy_8_981_268_AND_NOT_m_cfg__ETC___d3272,
       NOT_m_vrg_source_busy_9_982_276_AND_NOT_m_cfg__ETC___d3280,
       _dfoo1,
       _dfoo10,
       _dfoo100,
       _dfoo1000,
       _dfoo1001,
       _dfoo1002,
       _dfoo1003,
       _dfoo1004,
       _dfoo1005,
       _dfoo1006,
       _dfoo1007,
       _dfoo1008,
       _dfoo1009,
       _dfoo1010,
       _dfoo1011,
       _dfoo1012,
       _dfoo1013,
       _dfoo1014,
       _dfoo1015,
       _dfoo1016,
       _dfoo1017,
       _dfoo1018,
       _dfoo1019,
       _dfoo102,
       _dfoo1020,
       _dfoo1022,
       _dfoo1024,
       _dfoo1026,
       _dfoo1028,
       _dfoo1030,
       _dfoo1032,
       _dfoo1034,
       _dfoo1036,
       _dfoo1038,
       _dfoo104,
       _dfoo1040,
       _dfoo1042,
       _dfoo1044,
       _dfoo1046,
       _dfoo1048,
       _dfoo1050,
       _dfoo1052,
       _dfoo1054,
       _dfoo1056,
       _dfoo1058,
       _dfoo106,
       _dfoo1060,
       _dfoo1062,
       _dfoo1064,
       _dfoo1066,
       _dfoo1068,
       _dfoo1070,
       _dfoo1072,
       _dfoo1074,
       _dfoo1076,
       _dfoo1078,
       _dfoo108,
       _dfoo1080,
       _dfoo1082,
       _dfoo1084,
       _dfoo1086,
       _dfoo1088,
       _dfoo1089,
       _dfoo1090,
       _dfoo1091,
       _dfoo1092,
       _dfoo1093,
       _dfoo1094,
       _dfoo1095,
       _dfoo1096,
       _dfoo1097,
       _dfoo1098,
       _dfoo1099,
       _dfoo11,
       _dfoo110,
       _dfoo1100,
       _dfoo1101,
       _dfoo1102,
       _dfoo1103,
       _dfoo1104,
       _dfoo1105,
       _dfoo1106,
       _dfoo1107,
       _dfoo1108,
       _dfoo1109,
       _dfoo1110,
       _dfoo1111,
       _dfoo1112,
       _dfoo1113,
       _dfoo1114,
       _dfoo1115,
       _dfoo1116,
       _dfoo1117,
       _dfoo1118,
       _dfoo1119,
       _dfoo112,
       _dfoo1120,
       _dfoo1121,
       _dfoo1122,
       _dfoo1123,
       _dfoo1124,
       _dfoo1125,
       _dfoo1126,
       _dfoo1127,
       _dfoo1128,
       _dfoo1129,
       _dfoo1130,
       _dfoo1131,
       _dfoo1132,
       _dfoo1133,
       _dfoo1134,
       _dfoo1135,
       _dfoo1136,
       _dfoo1137,
       _dfoo1138,
       _dfoo1139,
       _dfoo114,
       _dfoo1140,
       _dfoo1141,
       _dfoo1142,
       _dfoo1143,
       _dfoo1144,
       _dfoo1145,
       _dfoo1146,
       _dfoo1147,
       _dfoo1148,
       _dfoo1149,
       _dfoo1150,
       _dfoo1151,
       _dfoo1152,
       _dfoo1153,
       _dfoo1154,
       _dfoo1155,
       _dfoo1156,
       _dfoo1158,
       _dfoo116,
       _dfoo1160,
       _dfoo1162,
       _dfoo1164,
       _dfoo1166,
       _dfoo1168,
       _dfoo1170,
       _dfoo1172,
       _dfoo1174,
       _dfoo1176,
       _dfoo1178,
       _dfoo118,
       _dfoo1180,
       _dfoo1182,
       _dfoo1184,
       _dfoo1186,
       _dfoo1188,
       _dfoo1190,
       _dfoo1192,
       _dfoo1194,
       _dfoo1196,
       _dfoo1198,
       _dfoo12,
       _dfoo120,
       _dfoo1200,
       _dfoo1202,
       _dfoo1204,
       _dfoo1206,
       _dfoo1208,
       _dfoo1210,
       _dfoo1212,
       _dfoo1214,
       _dfoo1216,
       _dfoo1218,
       _dfoo122,
       _dfoo1220,
       _dfoo1222,
       _dfoo1224,
       _dfoo1225,
       _dfoo1226,
       _dfoo1227,
       _dfoo1228,
       _dfoo1229,
       _dfoo1230,
       _dfoo1231,
       _dfoo1232,
       _dfoo1233,
       _dfoo1234,
       _dfoo1235,
       _dfoo1236,
       _dfoo1237,
       _dfoo1238,
       _dfoo1239,
       _dfoo124,
       _dfoo1240,
       _dfoo1241,
       _dfoo1242,
       _dfoo1243,
       _dfoo1244,
       _dfoo1245,
       _dfoo1246,
       _dfoo1247,
       _dfoo1248,
       _dfoo1249,
       _dfoo1250,
       _dfoo1251,
       _dfoo1252,
       _dfoo1253,
       _dfoo1254,
       _dfoo1255,
       _dfoo1256,
       _dfoo1257,
       _dfoo1258,
       _dfoo1259,
       _dfoo126,
       _dfoo1260,
       _dfoo1261,
       _dfoo1262,
       _dfoo1263,
       _dfoo1264,
       _dfoo1265,
       _dfoo1266,
       _dfoo1267,
       _dfoo1268,
       _dfoo1269,
       _dfoo1270,
       _dfoo1271,
       _dfoo1272,
       _dfoo1273,
       _dfoo1274,
       _dfoo1275,
       _dfoo1276,
       _dfoo1277,
       _dfoo1278,
       _dfoo1279,
       _dfoo128,
       _dfoo1280,
       _dfoo1281,
       _dfoo1282,
       _dfoo1283,
       _dfoo1284,
       _dfoo1285,
       _dfoo1286,
       _dfoo1287,
       _dfoo1288,
       _dfoo1289,
       _dfoo1290,
       _dfoo1291,
       _dfoo1292,
       _dfoo1294,
       _dfoo1296,
       _dfoo1298,
       _dfoo13,
       _dfoo130,
       _dfoo1300,
       _dfoo1302,
       _dfoo1304,
       _dfoo1306,
       _dfoo1308,
       _dfoo1310,
       _dfoo1312,
       _dfoo1314,
       _dfoo1316,
       _dfoo1318,
       _dfoo132,
       _dfoo1320,
       _dfoo1322,
       _dfoo1324,
       _dfoo1326,
       _dfoo1328,
       _dfoo1330,
       _dfoo1332,
       _dfoo1334,
       _dfoo1336,
       _dfoo1338,
       _dfoo134,
       _dfoo1340,
       _dfoo1342,
       _dfoo1344,
       _dfoo1346,
       _dfoo1348,
       _dfoo1350,
       _dfoo1352,
       _dfoo1354,
       _dfoo1356,
       _dfoo1358,
       _dfoo136,
       _dfoo1360,
       _dfoo1361,
       _dfoo1362,
       _dfoo1363,
       _dfoo1364,
       _dfoo1365,
       _dfoo1366,
       _dfoo1367,
       _dfoo1368,
       _dfoo1369,
       _dfoo137,
       _dfoo1370,
       _dfoo1371,
       _dfoo1372,
       _dfoo1373,
       _dfoo1374,
       _dfoo1375,
       _dfoo1376,
       _dfoo1377,
       _dfoo1378,
       _dfoo1379,
       _dfoo138,
       _dfoo1380,
       _dfoo1381,
       _dfoo1382,
       _dfoo1383,
       _dfoo1384,
       _dfoo1385,
       _dfoo1386,
       _dfoo1387,
       _dfoo1388,
       _dfoo1389,
       _dfoo139,
       _dfoo1390,
       _dfoo1391,
       _dfoo1392,
       _dfoo1393,
       _dfoo1394,
       _dfoo1395,
       _dfoo1396,
       _dfoo1397,
       _dfoo1398,
       _dfoo1399,
       _dfoo14,
       _dfoo140,
       _dfoo1400,
       _dfoo1401,
       _dfoo1402,
       _dfoo1403,
       _dfoo1404,
       _dfoo1405,
       _dfoo1406,
       _dfoo1407,
       _dfoo1408,
       _dfoo1409,
       _dfoo141,
       _dfoo1410,
       _dfoo1411,
       _dfoo1412,
       _dfoo1413,
       _dfoo1414,
       _dfoo1415,
       _dfoo1416,
       _dfoo1417,
       _dfoo1418,
       _dfoo1419,
       _dfoo142,
       _dfoo1420,
       _dfoo1421,
       _dfoo1422,
       _dfoo1423,
       _dfoo1424,
       _dfoo1425,
       _dfoo1426,
       _dfoo1427,
       _dfoo1428,
       _dfoo143,
       _dfoo1430,
       _dfoo1432,
       _dfoo1434,
       _dfoo1436,
       _dfoo1438,
       _dfoo144,
       _dfoo1440,
       _dfoo1442,
       _dfoo1444,
       _dfoo1446,
       _dfoo1448,
       _dfoo145,
       _dfoo1450,
       _dfoo1452,
       _dfoo1454,
       _dfoo1456,
       _dfoo1458,
       _dfoo146,
       _dfoo1460,
       _dfoo1462,
       _dfoo1464,
       _dfoo1466,
       _dfoo1468,
       _dfoo147,
       _dfoo1470,
       _dfoo1472,
       _dfoo1474,
       _dfoo1476,
       _dfoo1478,
       _dfoo148,
       _dfoo1480,
       _dfoo1482,
       _dfoo1484,
       _dfoo1486,
       _dfoo1488,
       _dfoo149,
       _dfoo1490,
       _dfoo1492,
       _dfoo1494,
       _dfoo1496,
       _dfoo1497,
       _dfoo1498,
       _dfoo1499,
       _dfoo15,
       _dfoo150,
       _dfoo1500,
       _dfoo1501,
       _dfoo1502,
       _dfoo1503,
       _dfoo1504,
       _dfoo1505,
       _dfoo1506,
       _dfoo1507,
       _dfoo1508,
       _dfoo1509,
       _dfoo151,
       _dfoo1510,
       _dfoo1511,
       _dfoo1512,
       _dfoo1513,
       _dfoo1514,
       _dfoo1515,
       _dfoo1516,
       _dfoo1517,
       _dfoo1518,
       _dfoo1519,
       _dfoo152,
       _dfoo1520,
       _dfoo1521,
       _dfoo1522,
       _dfoo1523,
       _dfoo1524,
       _dfoo1525,
       _dfoo1526,
       _dfoo1527,
       _dfoo1528,
       _dfoo1529,
       _dfoo153,
       _dfoo1530,
       _dfoo1531,
       _dfoo1532,
       _dfoo1533,
       _dfoo1534,
       _dfoo1535,
       _dfoo1536,
       _dfoo1537,
       _dfoo1538,
       _dfoo1539,
       _dfoo154,
       _dfoo1540,
       _dfoo1541,
       _dfoo1542,
       _dfoo1543,
       _dfoo1544,
       _dfoo1545,
       _dfoo1546,
       _dfoo1547,
       _dfoo1548,
       _dfoo1549,
       _dfoo155,
       _dfoo1550,
       _dfoo1551,
       _dfoo1552,
       _dfoo1553,
       _dfoo1554,
       _dfoo1555,
       _dfoo1556,
       _dfoo1557,
       _dfoo1558,
       _dfoo1559,
       _dfoo156,
       _dfoo1560,
       _dfoo1561,
       _dfoo1562,
       _dfoo1563,
       _dfoo1564,
       _dfoo1566,
       _dfoo1568,
       _dfoo157,
       _dfoo1570,
       _dfoo1572,
       _dfoo1574,
       _dfoo1576,
       _dfoo1578,
       _dfoo158,
       _dfoo1580,
       _dfoo1582,
       _dfoo1584,
       _dfoo1586,
       _dfoo1588,
       _dfoo159,
       _dfoo1590,
       _dfoo1592,
       _dfoo1594,
       _dfoo1596,
       _dfoo1598,
       _dfoo16,
       _dfoo160,
       _dfoo1600,
       _dfoo1602,
       _dfoo1604,
       _dfoo1606,
       _dfoo1608,
       _dfoo161,
       _dfoo1610,
       _dfoo1612,
       _dfoo1614,
       _dfoo1616,
       _dfoo1618,
       _dfoo162,
       _dfoo1620,
       _dfoo1622,
       _dfoo1624,
       _dfoo1626,
       _dfoo1628,
       _dfoo163,
       _dfoo1630,
       _dfoo1632,
       _dfoo1633,
       _dfoo1634,
       _dfoo1635,
       _dfoo1636,
       _dfoo1637,
       _dfoo1638,
       _dfoo1639,
       _dfoo164,
       _dfoo1640,
       _dfoo1641,
       _dfoo1642,
       _dfoo1643,
       _dfoo1644,
       _dfoo1645,
       _dfoo1646,
       _dfoo1647,
       _dfoo1648,
       _dfoo1649,
       _dfoo165,
       _dfoo1650,
       _dfoo1651,
       _dfoo1652,
       _dfoo1653,
       _dfoo1654,
       _dfoo1655,
       _dfoo1656,
       _dfoo1657,
       _dfoo1658,
       _dfoo1659,
       _dfoo166,
       _dfoo1660,
       _dfoo1661,
       _dfoo1662,
       _dfoo1663,
       _dfoo1664,
       _dfoo1665,
       _dfoo1666,
       _dfoo1667,
       _dfoo1668,
       _dfoo1669,
       _dfoo167,
       _dfoo1670,
       _dfoo1671,
       _dfoo1672,
       _dfoo1673,
       _dfoo1674,
       _dfoo1675,
       _dfoo1676,
       _dfoo1677,
       _dfoo1678,
       _dfoo1679,
       _dfoo168,
       _dfoo1680,
       _dfoo1681,
       _dfoo1682,
       _dfoo1683,
       _dfoo1684,
       _dfoo1685,
       _dfoo1686,
       _dfoo1687,
       _dfoo1688,
       _dfoo1689,
       _dfoo169,
       _dfoo1690,
       _dfoo1691,
       _dfoo1692,
       _dfoo1693,
       _dfoo1694,
       _dfoo1695,
       _dfoo1696,
       _dfoo1697,
       _dfoo1698,
       _dfoo1699,
       _dfoo17,
       _dfoo170,
       _dfoo1700,
       _dfoo1702,
       _dfoo1704,
       _dfoo1706,
       _dfoo1708,
       _dfoo171,
       _dfoo1710,
       _dfoo1712,
       _dfoo1714,
       _dfoo1716,
       _dfoo1718,
       _dfoo172,
       _dfoo1720,
       _dfoo1722,
       _dfoo1724,
       _dfoo1726,
       _dfoo1728,
       _dfoo173,
       _dfoo1730,
       _dfoo1732,
       _dfoo1734,
       _dfoo1736,
       _dfoo1738,
       _dfoo174,
       _dfoo1740,
       _dfoo1742,
       _dfoo1744,
       _dfoo1746,
       _dfoo1748,
       _dfoo175,
       _dfoo1750,
       _dfoo1752,
       _dfoo1754,
       _dfoo1756,
       _dfoo1758,
       _dfoo176,
       _dfoo1760,
       _dfoo1762,
       _dfoo1764,
       _dfoo1766,
       _dfoo1768,
       _dfoo1769,
       _dfoo177,
       _dfoo1770,
       _dfoo1771,
       _dfoo1772,
       _dfoo1773,
       _dfoo1774,
       _dfoo1775,
       _dfoo1776,
       _dfoo1777,
       _dfoo1778,
       _dfoo1779,
       _dfoo178,
       _dfoo1780,
       _dfoo1781,
       _dfoo1782,
       _dfoo1783,
       _dfoo1784,
       _dfoo1785,
       _dfoo1786,
       _dfoo1787,
       _dfoo1788,
       _dfoo1789,
       _dfoo179,
       _dfoo1790,
       _dfoo1791,
       _dfoo1792,
       _dfoo1793,
       _dfoo1794,
       _dfoo1795,
       _dfoo1796,
       _dfoo1797,
       _dfoo1798,
       _dfoo1799,
       _dfoo18,
       _dfoo180,
       _dfoo1800,
       _dfoo1801,
       _dfoo1802,
       _dfoo1803,
       _dfoo1804,
       _dfoo1805,
       _dfoo1806,
       _dfoo1807,
       _dfoo1808,
       _dfoo1809,
       _dfoo181,
       _dfoo1810,
       _dfoo1811,
       _dfoo1812,
       _dfoo1813,
       _dfoo1814,
       _dfoo1815,
       _dfoo1816,
       _dfoo1817,
       _dfoo1818,
       _dfoo1819,
       _dfoo182,
       _dfoo1820,
       _dfoo1821,
       _dfoo1822,
       _dfoo1823,
       _dfoo1824,
       _dfoo1825,
       _dfoo1826,
       _dfoo1827,
       _dfoo1828,
       _dfoo1829,
       _dfoo183,
       _dfoo1830,
       _dfoo1831,
       _dfoo1832,
       _dfoo1833,
       _dfoo1834,
       _dfoo1835,
       _dfoo1836,
       _dfoo1838,
       _dfoo184,
       _dfoo1840,
       _dfoo1842,
       _dfoo1844,
       _dfoo1846,
       _dfoo1848,
       _dfoo185,
       _dfoo1850,
       _dfoo1852,
       _dfoo1854,
       _dfoo1856,
       _dfoo1858,
       _dfoo186,
       _dfoo1860,
       _dfoo1862,
       _dfoo1864,
       _dfoo1866,
       _dfoo1868,
       _dfoo187,
       _dfoo1870,
       _dfoo1872,
       _dfoo1874,
       _dfoo1876,
       _dfoo1878,
       _dfoo188,
       _dfoo1880,
       _dfoo1882,
       _dfoo1884,
       _dfoo1886,
       _dfoo1888,
       _dfoo189,
       _dfoo1890,
       _dfoo1892,
       _dfoo1894,
       _dfoo1896,
       _dfoo1898,
       _dfoo19,
       _dfoo190,
       _dfoo1900,
       _dfoo1902,
       _dfoo1904,
       _dfoo1905,
       _dfoo1906,
       _dfoo1907,
       _dfoo1908,
       _dfoo1909,
       _dfoo191,
       _dfoo1910,
       _dfoo1911,
       _dfoo1912,
       _dfoo1913,
       _dfoo1914,
       _dfoo1915,
       _dfoo1916,
       _dfoo1917,
       _dfoo1918,
       _dfoo1919,
       _dfoo192,
       _dfoo1920,
       _dfoo1921,
       _dfoo1922,
       _dfoo1923,
       _dfoo1924,
       _dfoo1925,
       _dfoo1926,
       _dfoo1927,
       _dfoo1928,
       _dfoo1929,
       _dfoo193,
       _dfoo1930,
       _dfoo1931,
       _dfoo1932,
       _dfoo1933,
       _dfoo1934,
       _dfoo1935,
       _dfoo1936,
       _dfoo1937,
       _dfoo1938,
       _dfoo1939,
       _dfoo194,
       _dfoo1940,
       _dfoo1941,
       _dfoo1942,
       _dfoo1943,
       _dfoo1944,
       _dfoo1945,
       _dfoo1946,
       _dfoo1947,
       _dfoo1948,
       _dfoo1949,
       _dfoo195,
       _dfoo1950,
       _dfoo1951,
       _dfoo1952,
       _dfoo1953,
       _dfoo1954,
       _dfoo1955,
       _dfoo1956,
       _dfoo1957,
       _dfoo1958,
       _dfoo1959,
       _dfoo196,
       _dfoo1960,
       _dfoo1961,
       _dfoo1962,
       _dfoo1963,
       _dfoo1964,
       _dfoo1965,
       _dfoo1966,
       _dfoo1967,
       _dfoo1968,
       _dfoo1969,
       _dfoo197,
       _dfoo1970,
       _dfoo1971,
       _dfoo1972,
       _dfoo1974,
       _dfoo1976,
       _dfoo1978,
       _dfoo198,
       _dfoo1980,
       _dfoo1982,
       _dfoo1984,
       _dfoo1986,
       _dfoo1988,
       _dfoo199,
       _dfoo1990,
       _dfoo1992,
       _dfoo1994,
       _dfoo1996,
       _dfoo1998,
       _dfoo2,
       _dfoo20,
       _dfoo200,
       _dfoo2000,
       _dfoo2002,
       _dfoo2004,
       _dfoo2006,
       _dfoo2008,
       _dfoo201,
       _dfoo2010,
       _dfoo2012,
       _dfoo2014,
       _dfoo2016,
       _dfoo2018,
       _dfoo202,
       _dfoo2020,
       _dfoo2022,
       _dfoo2024,
       _dfoo2026,
       _dfoo2028,
       _dfoo203,
       _dfoo2030,
       _dfoo2032,
       _dfoo2034,
       _dfoo2036,
       _dfoo2038,
       _dfoo204,
       _dfoo2040,
       _dfoo2041,
       _dfoo2043,
       _dfoo2045,
       _dfoo2047,
       _dfoo2049,
       _dfoo2051,
       _dfoo2053,
       _dfoo2055,
       _dfoo2057,
       _dfoo2059,
       _dfoo206,
       _dfoo2061,
       _dfoo2063,
       _dfoo2065,
       _dfoo2067,
       _dfoo2069,
       _dfoo2071,
       _dfoo2073,
       _dfoo2075,
       _dfoo2077,
       _dfoo2079,
       _dfoo208,
       _dfoo2081,
       _dfoo2083,
       _dfoo2085,
       _dfoo2087,
       _dfoo2089,
       _dfoo2091,
       _dfoo2093,
       _dfoo2095,
       _dfoo2097,
       _dfoo2099,
       _dfoo21,
       _dfoo210,
       _dfoo2101,
       _dfoo2103,
       _dfoo2105,
       _dfoo2107,
       _dfoo212,
       _dfoo214,
       _dfoo216,
       _dfoo218,
       _dfoo22,
       _dfoo220,
       _dfoo222,
       _dfoo224,
       _dfoo226,
       _dfoo228,
       _dfoo23,
       _dfoo230,
       _dfoo232,
       _dfoo234,
       _dfoo236,
       _dfoo238,
       _dfoo24,
       _dfoo240,
       _dfoo242,
       _dfoo244,
       _dfoo246,
       _dfoo248,
       _dfoo25,
       _dfoo250,
       _dfoo252,
       _dfoo254,
       _dfoo256,
       _dfoo258,
       _dfoo26,
       _dfoo260,
       _dfoo262,
       _dfoo264,
       _dfoo266,
       _dfoo268,
       _dfoo27,
       _dfoo270,
       _dfoo272,
       _dfoo273,
       _dfoo274,
       _dfoo275,
       _dfoo276,
       _dfoo277,
       _dfoo278,
       _dfoo279,
       _dfoo28,
       _dfoo280,
       _dfoo281,
       _dfoo282,
       _dfoo283,
       _dfoo284,
       _dfoo285,
       _dfoo286,
       _dfoo287,
       _dfoo288,
       _dfoo289,
       _dfoo29,
       _dfoo290,
       _dfoo291,
       _dfoo292,
       _dfoo293,
       _dfoo294,
       _dfoo295,
       _dfoo296,
       _dfoo297,
       _dfoo298,
       _dfoo299,
       _dfoo3,
       _dfoo30,
       _dfoo300,
       _dfoo301,
       _dfoo302,
       _dfoo303,
       _dfoo304,
       _dfoo305,
       _dfoo306,
       _dfoo307,
       _dfoo308,
       _dfoo309,
       _dfoo31,
       _dfoo310,
       _dfoo311,
       _dfoo312,
       _dfoo313,
       _dfoo314,
       _dfoo315,
       _dfoo316,
       _dfoo317,
       _dfoo318,
       _dfoo319,
       _dfoo32,
       _dfoo320,
       _dfoo321,
       _dfoo322,
       _dfoo323,
       _dfoo324,
       _dfoo325,
       _dfoo326,
       _dfoo327,
       _dfoo328,
       _dfoo329,
       _dfoo33,
       _dfoo330,
       _dfoo331,
       _dfoo332,
       _dfoo333,
       _dfoo334,
       _dfoo335,
       _dfoo336,
       _dfoo337,
       _dfoo338,
       _dfoo339,
       _dfoo34,
       _dfoo340,
       _dfoo342,
       _dfoo344,
       _dfoo346,
       _dfoo348,
       _dfoo35,
       _dfoo350,
       _dfoo352,
       _dfoo354,
       _dfoo356,
       _dfoo358,
       _dfoo36,
       _dfoo360,
       _dfoo362,
       _dfoo364,
       _dfoo366,
       _dfoo368,
       _dfoo37,
       _dfoo370,
       _dfoo372,
       _dfoo374,
       _dfoo376,
       _dfoo378,
       _dfoo38,
       _dfoo380,
       _dfoo382,
       _dfoo384,
       _dfoo386,
       _dfoo388,
       _dfoo39,
       _dfoo390,
       _dfoo392,
       _dfoo394,
       _dfoo396,
       _dfoo398,
       _dfoo4,
       _dfoo40,
       _dfoo400,
       _dfoo402,
       _dfoo404,
       _dfoo406,
       _dfoo408,
       _dfoo409,
       _dfoo41,
       _dfoo410,
       _dfoo411,
       _dfoo412,
       _dfoo413,
       _dfoo414,
       _dfoo415,
       _dfoo416,
       _dfoo417,
       _dfoo418,
       _dfoo419,
       _dfoo42,
       _dfoo420,
       _dfoo421,
       _dfoo422,
       _dfoo423,
       _dfoo424,
       _dfoo425,
       _dfoo426,
       _dfoo427,
       _dfoo428,
       _dfoo429,
       _dfoo43,
       _dfoo430,
       _dfoo431,
       _dfoo432,
       _dfoo433,
       _dfoo434,
       _dfoo435,
       _dfoo436,
       _dfoo437,
       _dfoo438,
       _dfoo439,
       _dfoo44,
       _dfoo440,
       _dfoo441,
       _dfoo442,
       _dfoo443,
       _dfoo444,
       _dfoo445,
       _dfoo446,
       _dfoo447,
       _dfoo448,
       _dfoo449,
       _dfoo45,
       _dfoo450,
       _dfoo451,
       _dfoo452,
       _dfoo453,
       _dfoo454,
       _dfoo455,
       _dfoo456,
       _dfoo457,
       _dfoo458,
       _dfoo459,
       _dfoo46,
       _dfoo460,
       _dfoo461,
       _dfoo462,
       _dfoo463,
       _dfoo464,
       _dfoo465,
       _dfoo466,
       _dfoo467,
       _dfoo468,
       _dfoo469,
       _dfoo47,
       _dfoo470,
       _dfoo471,
       _dfoo472,
       _dfoo473,
       _dfoo474,
       _dfoo475,
       _dfoo476,
       _dfoo478,
       _dfoo48,
       _dfoo480,
       _dfoo482,
       _dfoo484,
       _dfoo486,
       _dfoo488,
       _dfoo49,
       _dfoo490,
       _dfoo492,
       _dfoo494,
       _dfoo496,
       _dfoo498,
       _dfoo5,
       _dfoo50,
       _dfoo500,
       _dfoo502,
       _dfoo504,
       _dfoo506,
       _dfoo508,
       _dfoo51,
       _dfoo510,
       _dfoo512,
       _dfoo514,
       _dfoo516,
       _dfoo518,
       _dfoo52,
       _dfoo520,
       _dfoo522,
       _dfoo524,
       _dfoo526,
       _dfoo528,
       _dfoo53,
       _dfoo530,
       _dfoo532,
       _dfoo534,
       _dfoo536,
       _dfoo538,
       _dfoo54,
       _dfoo540,
       _dfoo542,
       _dfoo544,
       _dfoo545,
       _dfoo546,
       _dfoo547,
       _dfoo548,
       _dfoo549,
       _dfoo55,
       _dfoo550,
       _dfoo551,
       _dfoo552,
       _dfoo553,
       _dfoo554,
       _dfoo555,
       _dfoo556,
       _dfoo557,
       _dfoo558,
       _dfoo559,
       _dfoo56,
       _dfoo560,
       _dfoo561,
       _dfoo562,
       _dfoo563,
       _dfoo564,
       _dfoo565,
       _dfoo566,
       _dfoo567,
       _dfoo568,
       _dfoo569,
       _dfoo57,
       _dfoo570,
       _dfoo571,
       _dfoo572,
       _dfoo573,
       _dfoo574,
       _dfoo575,
       _dfoo576,
       _dfoo577,
       _dfoo578,
       _dfoo579,
       _dfoo58,
       _dfoo580,
       _dfoo581,
       _dfoo582,
       _dfoo583,
       _dfoo584,
       _dfoo585,
       _dfoo586,
       _dfoo587,
       _dfoo588,
       _dfoo589,
       _dfoo59,
       _dfoo590,
       _dfoo591,
       _dfoo592,
       _dfoo593,
       _dfoo594,
       _dfoo595,
       _dfoo596,
       _dfoo597,
       _dfoo598,
       _dfoo599,
       _dfoo6,
       _dfoo60,
       _dfoo600,
       _dfoo601,
       _dfoo602,
       _dfoo603,
       _dfoo604,
       _dfoo605,
       _dfoo606,
       _dfoo607,
       _dfoo608,
       _dfoo609,
       _dfoo61,
       _dfoo610,
       _dfoo611,
       _dfoo612,
       _dfoo614,
       _dfoo616,
       _dfoo618,
       _dfoo62,
       _dfoo620,
       _dfoo622,
       _dfoo624,
       _dfoo626,
       _dfoo628,
       _dfoo63,
       _dfoo630,
       _dfoo632,
       _dfoo634,
       _dfoo636,
       _dfoo638,
       _dfoo64,
       _dfoo640,
       _dfoo642,
       _dfoo644,
       _dfoo646,
       _dfoo648,
       _dfoo65,
       _dfoo650,
       _dfoo652,
       _dfoo654,
       _dfoo656,
       _dfoo658,
       _dfoo66,
       _dfoo660,
       _dfoo662,
       _dfoo664,
       _dfoo666,
       _dfoo668,
       _dfoo67,
       _dfoo670,
       _dfoo672,
       _dfoo674,
       _dfoo676,
       _dfoo678,
       _dfoo68,
       _dfoo680,
       _dfoo681,
       _dfoo682,
       _dfoo683,
       _dfoo684,
       _dfoo685,
       _dfoo686,
       _dfoo687,
       _dfoo688,
       _dfoo689,
       _dfoo690,
       _dfoo691,
       _dfoo692,
       _dfoo693,
       _dfoo694,
       _dfoo695,
       _dfoo696,
       _dfoo697,
       _dfoo698,
       _dfoo699,
       _dfoo7,
       _dfoo70,
       _dfoo700,
       _dfoo701,
       _dfoo702,
       _dfoo703,
       _dfoo704,
       _dfoo705,
       _dfoo706,
       _dfoo707,
       _dfoo708,
       _dfoo709,
       _dfoo710,
       _dfoo711,
       _dfoo712,
       _dfoo713,
       _dfoo714,
       _dfoo715,
       _dfoo716,
       _dfoo717,
       _dfoo718,
       _dfoo719,
       _dfoo72,
       _dfoo720,
       _dfoo721,
       _dfoo722,
       _dfoo723,
       _dfoo724,
       _dfoo725,
       _dfoo726,
       _dfoo727,
       _dfoo728,
       _dfoo729,
       _dfoo730,
       _dfoo731,
       _dfoo732,
       _dfoo733,
       _dfoo734,
       _dfoo735,
       _dfoo736,
       _dfoo737,
       _dfoo738,
       _dfoo739,
       _dfoo74,
       _dfoo740,
       _dfoo741,
       _dfoo742,
       _dfoo743,
       _dfoo744,
       _dfoo745,
       _dfoo746,
       _dfoo747,
       _dfoo748,
       _dfoo750,
       _dfoo752,
       _dfoo754,
       _dfoo756,
       _dfoo758,
       _dfoo76,
       _dfoo760,
       _dfoo762,
       _dfoo764,
       _dfoo766,
       _dfoo768,
       _dfoo770,
       _dfoo772,
       _dfoo774,
       _dfoo776,
       _dfoo778,
       _dfoo78,
       _dfoo780,
       _dfoo782,
       _dfoo784,
       _dfoo786,
       _dfoo788,
       _dfoo790,
       _dfoo792,
       _dfoo794,
       _dfoo796,
       _dfoo798,
       _dfoo8,
       _dfoo80,
       _dfoo800,
       _dfoo802,
       _dfoo804,
       _dfoo806,
       _dfoo808,
       _dfoo810,
       _dfoo812,
       _dfoo814,
       _dfoo816,
       _dfoo817,
       _dfoo818,
       _dfoo819,
       _dfoo82,
       _dfoo820,
       _dfoo821,
       _dfoo822,
       _dfoo823,
       _dfoo824,
       _dfoo825,
       _dfoo826,
       _dfoo827,
       _dfoo828,
       _dfoo829,
       _dfoo830,
       _dfoo831,
       _dfoo832,
       _dfoo833,
       _dfoo834,
       _dfoo835,
       _dfoo836,
       _dfoo837,
       _dfoo838,
       _dfoo839,
       _dfoo84,
       _dfoo840,
       _dfoo841,
       _dfoo842,
       _dfoo843,
       _dfoo844,
       _dfoo845,
       _dfoo846,
       _dfoo847,
       _dfoo848,
       _dfoo849,
       _dfoo850,
       _dfoo851,
       _dfoo852,
       _dfoo853,
       _dfoo854,
       _dfoo855,
       _dfoo856,
       _dfoo857,
       _dfoo858,
       _dfoo859,
       _dfoo86,
       _dfoo860,
       _dfoo861,
       _dfoo862,
       _dfoo863,
       _dfoo864,
       _dfoo865,
       _dfoo866,
       _dfoo867,
       _dfoo868,
       _dfoo869,
       _dfoo870,
       _dfoo871,
       _dfoo872,
       _dfoo873,
       _dfoo874,
       _dfoo875,
       _dfoo876,
       _dfoo877,
       _dfoo878,
       _dfoo879,
       _dfoo88,
       _dfoo880,
       _dfoo881,
       _dfoo882,
       _dfoo883,
       _dfoo884,
       _dfoo886,
       _dfoo888,
       _dfoo890,
       _dfoo892,
       _dfoo894,
       _dfoo896,
       _dfoo898,
       _dfoo9,
       _dfoo90,
       _dfoo900,
       _dfoo902,
       _dfoo904,
       _dfoo906,
       _dfoo908,
       _dfoo910,
       _dfoo912,
       _dfoo914,
       _dfoo916,
       _dfoo918,
       _dfoo92,
       _dfoo920,
       _dfoo922,
       _dfoo924,
       _dfoo926,
       _dfoo928,
       _dfoo930,
       _dfoo932,
       _dfoo934,
       _dfoo936,
       _dfoo938,
       _dfoo94,
       _dfoo940,
       _dfoo942,
       _dfoo944,
       _dfoo946,
       _dfoo948,
       _dfoo950,
       _dfoo952,
       _dfoo953,
       _dfoo954,
       _dfoo955,
       _dfoo956,
       _dfoo957,
       _dfoo958,
       _dfoo959,
       _dfoo96,
       _dfoo960,
       _dfoo961,
       _dfoo962,
       _dfoo963,
       _dfoo964,
       _dfoo965,
       _dfoo966,
       _dfoo967,
       _dfoo968,
       _dfoo969,
       _dfoo970,
       _dfoo971,
       _dfoo972,
       _dfoo973,
       _dfoo974,
       _dfoo975,
       _dfoo976,
       _dfoo977,
       _dfoo978,
       _dfoo979,
       _dfoo98,
       _dfoo980,
       _dfoo981,
       _dfoo982,
       _dfoo983,
       _dfoo984,
       _dfoo985,
       _dfoo986,
       _dfoo987,
       _dfoo988,
       _dfoo989,
       _dfoo990,
       _dfoo991,
       _dfoo992,
       _dfoo993,
       _dfoo994,
       _dfoo995,
       _dfoo996,
       _dfoo997,
       _dfoo998,
       _dfoo999,
       m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d240,
       m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d242,
       m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d31,
       m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d36,
       m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d40,
       m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d43,
       m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d532,
       m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d68,
       m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d71,
       m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d2854,
       m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d2860,
       m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d2862,
       m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812,
       m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d821,
       m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d823,
       m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d837,
       m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d839,
       m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d841,
       m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d843,
       m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d845,
       m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d847,
       m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d849,
       m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d851,
       m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d853,
       m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d855,
       m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d857,
       m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d859,
       m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d861,
       m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d863,
       m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d865,
       m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d867,
       m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d869,
       m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d874,
       m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d877,
       m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d888,
       m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d889,
       m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d895,
       m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d931,
       m_vrg_source_ip_10_read__0_AND_NOT_m_vrg_sourc_ETC___d3036,
       m_vrg_source_ip_10_read__0_AND_NOT_m_vrg_sourc_ETC___d3130,
       m_vrg_source_ip_10_read__0_AND_NOT_m_vrg_sourc_ETC___d614,
       m_vrg_source_ip_11_read__1_AND_NOT_m_vrg_sourc_ETC___d3041,
       m_vrg_source_ip_11_read__1_AND_NOT_m_vrg_sourc_ETC___d3135,
       m_vrg_source_ip_11_read__1_AND_NOT_m_vrg_sourc_ETC___d621,
       m_vrg_source_ip_12_read__2_AND_NOT_m_vrg_sourc_ETC___d3046,
       m_vrg_source_ip_12_read__2_AND_NOT_m_vrg_sourc_ETC___d3140,
       m_vrg_source_ip_12_read__2_AND_NOT_m_vrg_sourc_ETC___d628,
       m_vrg_source_ip_13_read__3_AND_NOT_m_vrg_sourc_ETC___d3051,
       m_vrg_source_ip_13_read__3_AND_NOT_m_vrg_sourc_ETC___d3145,
       m_vrg_source_ip_13_read__3_AND_NOT_m_vrg_sourc_ETC___d635,
       m_vrg_source_ip_13_read__3_AND_NOT_m_vrg_sourc_ETC___d686,
       m_vrg_source_ip_14_read__4_AND_NOT_m_vrg_sourc_ETC___d3056,
       m_vrg_source_ip_14_read__4_AND_NOT_m_vrg_sourc_ETC___d3150,
       m_vrg_source_ip_14_read__4_AND_NOT_m_vrg_sourc_ETC___d642,
       m_vrg_source_ip_15_read__5_AND_NOT_m_vrg_sourc_ETC___d3061,
       m_vrg_source_ip_15_read__5_AND_NOT_m_vrg_sourc_ETC___d3155,
       m_vrg_source_ip_15_read__5_AND_NOT_m_vrg_sourc_ETC___d649,
       m_vrg_source_ip_16_read__6_AND_NOT_m_vrg_sourc_ETC___d3066,
       m_vrg_source_ip_16_read__6_AND_NOT_m_vrg_sourc_ETC___d3160,
       m_vrg_source_ip_16_read__6_AND_NOT_m_vrg_sourc_ETC___d656,
       m_vrg_source_ip_16_read__6_AND_NOT_m_vrg_sourc_ETC___d689,
       m_vrg_source_ip_1_read__1_AND_NOT_m_vrg_source_ETC___d551,
       m_vrg_source_ip_2_read__2_AND_NOT_m_vrg_source_ETC___d2996,
       m_vrg_source_ip_2_read__2_AND_NOT_m_vrg_source_ETC___d3090,
       m_vrg_source_ip_2_read__2_AND_NOT_m_vrg_source_ETC___d558,
       m_vrg_source_ip_3_read__3_AND_NOT_m_vrg_source_ETC___d3001,
       m_vrg_source_ip_3_read__3_AND_NOT_m_vrg_source_ETC___d3095,
       m_vrg_source_ip_3_read__3_AND_NOT_m_vrg_source_ETC___d565,
       m_vrg_source_ip_4_read__4_AND_NOT_m_vrg_source_ETC___d3006,
       m_vrg_source_ip_4_read__4_AND_NOT_m_vrg_source_ETC___d3100,
       m_vrg_source_ip_4_read__4_AND_NOT_m_vrg_source_ETC___d572,
       m_vrg_source_ip_5_read__5_AND_NOT_m_vrg_source_ETC___d3011,
       m_vrg_source_ip_5_read__5_AND_NOT_m_vrg_source_ETC___d3105,
       m_vrg_source_ip_5_read__5_AND_NOT_m_vrg_source_ETC___d579,
       m_vrg_source_ip_6_read__6_AND_NOT_m_vrg_source_ETC___d3016,
       m_vrg_source_ip_6_read__6_AND_NOT_m_vrg_source_ETC___d3110,
       m_vrg_source_ip_6_read__6_AND_NOT_m_vrg_source_ETC___d586,
       m_vrg_source_ip_7_read__7_AND_NOT_m_vrg_source_ETC___d3021,
       m_vrg_source_ip_7_read__7_AND_NOT_m_vrg_source_ETC___d3115,
       m_vrg_source_ip_7_read__7_AND_NOT_m_vrg_source_ETC___d593,
       m_vrg_source_ip_7_read__7_AND_NOT_m_vrg_source_ETC___d680,
       m_vrg_source_ip_8_read__8_AND_NOT_m_vrg_source_ETC___d3026,
       m_vrg_source_ip_8_read__8_AND_NOT_m_vrg_source_ETC___d3120,
       m_vrg_source_ip_8_read__8_AND_NOT_m_vrg_source_ETC___d600,
       m_vrg_source_ip_9_read__9_AND_NOT_m_vrg_source_ETC___d3031,
       m_vrg_source_ip_9_read__9_AND_NOT_m_vrg_source_ETC___d3125,
       m_vrg_source_ip_9_read__9_AND_NOT_m_vrg_source_ETC___d607,
       m_vrg_source_prio_16_3_ULE_IF_m_vrg_source_ip__ETC___d651;
  // action method set_verbosity
  assign RDY_set_verbosity = 1'd1 ;
  assign CAN_FIRE_set_verbosity = 1'd1 ;
  assign WILL_FIRE_set_verbosity = EN_set_verbosity ;
  // action method show_PLIC_state
  assign RDY_show_PLIC_state = 1'd1 ;
  assign CAN_FIRE_show_PLIC_state = 1'd1 ;
  assign WILL_FIRE_show_PLIC_state = EN_show_PLIC_state ;
  // action method server_reset_request_put
  assign RDY_server_reset_request_put = m_f_reset_reqs$FULL_N ;
  assign CAN_FIRE_server_reset_request_put = m_f_reset_reqs$FULL_N ;
  assign WILL_FIRE_server_reset_request_put = EN_server_reset_request_put ;
  // action method server_reset_response_get
  assign RDY_server_reset_response_get = m_f_reset_rsps$EMPTY_N ;
  assign CAN_FIRE_server_reset_response_get = m_f_reset_rsps$EMPTY_N ;
  assign WILL_FIRE_server_reset_response_get = EN_server_reset_response_get ;
  // action method set_addr_map
  assign RDY_set_addr_map = 1'd1 ;
  assign CAN_FIRE_set_addr_map = 1'd1 ;
  assign WILL_FIRE_set_addr_map = EN_set_addr_map ;
  // action method axi4_slave_m_awvalid
  assign CAN_FIRE_axi4_slave_m_awvalid = 1'd1 ;
  assign WILL_FIRE_axi4_slave_m_awvalid = 1'd1 ;
  // value method axi4_slave_m_awready
  assign axi4_slave_awready = m_slave_xactor_f_wr_addr$FULL_N ;
  // action method axi4_slave_m_wvalid
  assign CAN_FIRE_axi4_slave_m_wvalid = 1'd1 ;
  assign WILL_FIRE_axi4_slave_m_wvalid = 1'd1 ;
  // value method axi4_slave_m_wready
  assign axi4_slave_wready = m_slave_xactor_f_wr_data$FULL_N ;
  // value method axi4_slave_m_bvalid
  assign axi4_slave_bvalid = m_slave_xactor_f_wr_resp$EMPTY_N ;
  // value method axi4_slave_m_bid
  assign axi4_slave_bid = m_slave_xactor_f_wr_resp$D_OUT[5:2] ;
  // value method axi4_slave_m_bresp
  assign axi4_slave_bresp = m_slave_xactor_f_wr_resp$D_OUT[1:0] ;
  // action method axi4_slave_m_bready
  assign CAN_FIRE_axi4_slave_m_bready = 1'd1 ;
  assign WILL_FIRE_axi4_slave_m_bready = 1'd1 ;
  // action method axi4_slave_m_arvalid
  assign CAN_FIRE_axi4_slave_m_arvalid = 1'd1 ;
  assign WILL_FIRE_axi4_slave_m_arvalid = 1'd1 ;
  // value method axi4_slave_m_arready
  assign axi4_slave_arready = m_slave_xactor_f_rd_addr$FULL_N ;
  // value method axi4_slave_m_rvalid
  assign axi4_slave_rvalid = m_slave_xactor_f_rd_data$EMPTY_N ;
  // value method axi4_slave_m_rid
  assign axi4_slave_rid = m_slave_xactor_f_rd_data$D_OUT[70:67] ;
  // value method axi4_slave_m_rdata
  assign axi4_slave_rdata = m_slave_xactor_f_rd_data$D_OUT[66:3] ;
  // value method axi4_slave_m_rresp
  assign axi4_slave_rresp = m_slave_xactor_f_rd_data$D_OUT[2:1] ;
  // value method axi4_slave_m_rlast
  assign axi4_slave_rlast = m_slave_xactor_f_rd_data$D_OUT[0] ;
  // action method axi4_slave_m_rready
  assign CAN_FIRE_axi4_slave_m_rready = 1'd1 ;
  assign WILL_FIRE_axi4_slave_m_rready = 1'd1 ;
  // action method v_sources_0_m_interrupt_req
  assign CAN_FIRE_v_sources_0_m_interrupt_req = 1'd1 ;
  assign WILL_FIRE_v_sources_0_m_interrupt_req = 1'd1 ;
  // action method v_sources_1_m_interrupt_req
  assign CAN_FIRE_v_sources_1_m_interrupt_req = 1'd1 ;
  assign WILL_FIRE_v_sources_1_m_interrupt_req = 1'd1 ;
  // action method v_sources_2_m_interrupt_req
  assign CAN_FIRE_v_sources_2_m_interrupt_req = 1'd1 ;
  assign WILL_FIRE_v_sources_2_m_interrupt_req = 1'd1 ;
  // action method v_sources_3_m_interrupt_req
  assign CAN_FIRE_v_sources_3_m_interrupt_req = 1'd1 ;
  assign WILL_FIRE_v_sources_3_m_interrupt_req = 1'd1 ;
  // action method v_sources_4_m_interrupt_req
  assign CAN_FIRE_v_sources_4_m_interrupt_req = 1'd1 ;
  assign WILL_FIRE_v_sources_4_m_interrupt_req = 1'd1 ;
  // action method v_sources_5_m_interrupt_req
  assign CAN_FIRE_v_sources_5_m_interrupt_req = 1'd1 ;
  assign WILL_FIRE_v_sources_5_m_interrupt_req = 1'd1 ;
  // action method v_sources_6_m_interrupt_req
  assign CAN_FIRE_v_sources_6_m_interrupt_req = 1'd1 ;
  assign WILL_FIRE_v_sources_6_m_interrupt_req = 1'd1 ;
  // action method v_sources_7_m_interrupt_req
  assign CAN_FIRE_v_sources_7_m_interrupt_req = 1'd1 ;
  assign WILL_FIRE_v_sources_7_m_interrupt_req = 1'd1 ;
  // action method v_sources_8_m_interrupt_req
  assign CAN_FIRE_v_sources_8_m_interrupt_req = 1'd1 ;
  assign WILL_FIRE_v_sources_8_m_interrupt_req = 1'd1 ;
  // action method v_sources_9_m_interrupt_req
  assign CAN_FIRE_v_sources_9_m_interrupt_req = 1'd1 ;
  assign WILL_FIRE_v_sources_9_m_interrupt_req = 1'd1 ;
  // action method v_sources_10_m_interrupt_req
  assign CAN_FIRE_v_sources_10_m_interrupt_req = 1'd1 ;
  assign WILL_FIRE_v_sources_10_m_interrupt_req = 1'd1 ;
  // action method v_sources_11_m_interrupt_req
  assign CAN_FIRE_v_sources_11_m_interrupt_req = 1'd1 ;
  assign WILL_FIRE_v_sources_11_m_interrupt_req = 1'd1 ;
  // action method v_sources_12_m_interrupt_req
  assign CAN_FIRE_v_sources_12_m_interrupt_req = 1'd1 ;
  assign WILL_FIRE_v_sources_12_m_interrupt_req = 1'd1 ;
  // action method v_sources_13_m_interrupt_req
  assign CAN_FIRE_v_sources_13_m_interrupt_req = 1'd1 ;
  assign WILL_FIRE_v_sources_13_m_interrupt_req = 1'd1 ;
  // action method v_sources_14_m_interrupt_req
  assign CAN_FIRE_v_sources_14_m_interrupt_req = 1'd1 ;
  assign WILL_FIRE_v_sources_14_m_interrupt_req = 1'd1 ;
  // action method v_sources_15_m_interrupt_req
  assign CAN_FIRE_v_sources_15_m_interrupt_req = 1'd1 ;
  assign WILL_FIRE_v_sources_15_m_interrupt_req = 1'd1 ;
  // value method v_targets_0_m_eip
  assign v_targets_0_m_eip = a__h81740 > m_vrg_target_threshold_0 ;
  // value method v_targets_1_m_eip
  assign v_targets_1_m_eip = a__h83894 > m_vrg_target_threshold_1 ;
  // submodule m_f_reset_reqs
  FIFO20 #(.guarded(1'd1)) m_f_reset_reqs(.RST(RST_N),
					  .CLK(CLK),
					  .ENQ(m_f_reset_reqs$ENQ),
					  .DEQ(m_f_reset_reqs$DEQ),
					  .CLR(m_f_reset_reqs$CLR),
					  .FULL_N(m_f_reset_reqs$FULL_N),
					  .EMPTY_N(m_f_reset_reqs$EMPTY_N));
  // submodule m_f_reset_rsps
  FIFO20 #(.guarded(1'd1)) m_f_reset_rsps(.RST(RST_N),
					  .CLK(CLK),
					  .ENQ(m_f_reset_rsps$ENQ),
					  .DEQ(m_f_reset_rsps$DEQ),
					  .CLR(m_f_reset_rsps$CLR),
					  .FULL_N(m_f_reset_rsps$FULL_N),
					  .EMPTY_N(m_f_reset_rsps$EMPTY_N));
  // submodule m_slave_xactor_f_rd_addr
  FIFO2 #(.width(32'd97),
	  .guarded(1'd1)) m_slave_xactor_f_rd_addr(.RST(RST_N),
						   .CLK(CLK),
						   .D_IN(m_slave_xactor_f_rd_addr$D_IN),
						   .ENQ(m_slave_xactor_f_rd_addr$ENQ),
						   .DEQ(m_slave_xactor_f_rd_addr$DEQ),
						   .CLR(m_slave_xactor_f_rd_addr$CLR),
						   .D_OUT(m_slave_xactor_f_rd_addr$D_OUT),
						   .FULL_N(m_slave_xactor_f_rd_addr$FULL_N),
						   .EMPTY_N(m_slave_xactor_f_rd_addr$EMPTY_N));
  // submodule m_slave_xactor_f_rd_data
  FIFO2 #(.width(32'd71),
	  .guarded(1'd1)) m_slave_xactor_f_rd_data(.RST(RST_N),
						   .CLK(CLK),
						   .D_IN(m_slave_xactor_f_rd_data$D_IN),
						   .ENQ(m_slave_xactor_f_rd_data$ENQ),
						   .DEQ(m_slave_xactor_f_rd_data$DEQ),
						   .CLR(m_slave_xactor_f_rd_data$CLR),
						   .D_OUT(m_slave_xactor_f_rd_data$D_OUT),
						   .FULL_N(m_slave_xactor_f_rd_data$FULL_N),
						   .EMPTY_N(m_slave_xactor_f_rd_data$EMPTY_N));
  // submodule m_slave_xactor_f_wr_addr
  FIFO2 #(.width(32'd97),
	  .guarded(1'd1)) m_slave_xactor_f_wr_addr(.RST(RST_N),
						   .CLK(CLK),
						   .D_IN(m_slave_xactor_f_wr_addr$D_IN),
						   .ENQ(m_slave_xactor_f_wr_addr$ENQ),
						   .DEQ(m_slave_xactor_f_wr_addr$DEQ),
						   .CLR(m_slave_xactor_f_wr_addr$CLR),
						   .D_OUT(m_slave_xactor_f_wr_addr$D_OUT),
						   .FULL_N(m_slave_xactor_f_wr_addr$FULL_N),
						   .EMPTY_N(m_slave_xactor_f_wr_addr$EMPTY_N));
  // submodule m_slave_xactor_f_wr_data
  FIFO2 #(.width(32'd73),
	  .guarded(1'd1)) m_slave_xactor_f_wr_data(.RST(RST_N),
						   .CLK(CLK),
						   .D_IN(m_slave_xactor_f_wr_data$D_IN),
						   .ENQ(m_slave_xactor_f_wr_data$ENQ),
						   .DEQ(m_slave_xactor_f_wr_data$DEQ),
						   .CLR(m_slave_xactor_f_wr_data$CLR),
						   .D_OUT(m_slave_xactor_f_wr_data$D_OUT),
						   .FULL_N(m_slave_xactor_f_wr_data$FULL_N),
						   .EMPTY_N(m_slave_xactor_f_wr_data$EMPTY_N));
  // submodule m_slave_xactor_f_wr_resp
  FIFO2 #(.width(32'd6), .guarded(1'd1)) m_slave_xactor_f_wr_resp(.RST(RST_N),
								  .CLK(CLK),
								  .D_IN(m_slave_xactor_f_wr_resp$D_IN),
								  .ENQ(m_slave_xactor_f_wr_resp$ENQ),
								  .DEQ(m_slave_xactor_f_wr_resp$DEQ),
								  .CLR(m_slave_xactor_f_wr_resp$CLR),
								  .D_OUT(m_slave_xactor_f_wr_resp$D_OUT),
								  .FULL_N(m_slave_xactor_f_wr_resp$FULL_N),
								  .EMPTY_N(m_slave_xactor_f_wr_resp$EMPTY_N));
  // rule RL_m_rl_reset
  assign CAN_FIRE_RL_m_rl_reset =
	     m_f_reset_reqs$EMPTY_N && m_f_reset_rsps$FULL_N ;
  assign WILL_FIRE_RL_m_rl_reset = CAN_FIRE_RL_m_rl_reset ;
  // rule RL_m_rl_process_rd_req
  assign CAN_FIRE_RL_m_rl_process_rd_req =
	     m_slave_xactor_f_rd_addr$EMPTY_N &&
	     m_slave_xactor_f_rd_data$FULL_N &&
	     !m_f_reset_reqs$EMPTY_N ;
  assign WILL_FIRE_RL_m_rl_process_rd_req = CAN_FIRE_RL_m_rl_process_rd_req ;
  // rule RL_m_rl_process_wr_req
  assign CAN_FIRE_RL_m_rl_process_wr_req =
	     m_slave_xactor_f_wr_addr$EMPTY_N &&
	     m_slave_xactor_f_wr_data$EMPTY_N &&
	     m_slave_xactor_f_wr_resp$FULL_N &&
	     !m_f_reset_reqs$EMPTY_N ;
  assign WILL_FIRE_RL_m_rl_process_wr_req = CAN_FIRE_RL_m_rl_process_wr_req ;
  // inputs to muxes for submodule ports
  assign MUX_m_vrg_source_busy_0$write_1__SEL_1 =
	     WILL_FIRE_RL_m_rl_process_wr_req &&
	     wdata32__h27246[9:0] == 10'd0 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2884 ;
  assign MUX_m_vrg_source_busy_0$write_1__SEL_2 =
	     WILL_FIRE_RL_m_rl_process_rd_req && max_id__h24210 == 5'd0 &&
	     NOT_m_slave_xactor_f_rd_addr_first__9_BITS_92__ETC___d695 ;
  assign MUX_m_vrg_source_busy_1$write_1__SEL_1 =
	     WILL_FIRE_RL_m_rl_process_wr_req &&
	     wdata32__h27246[9:0] == 10'd1 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2884 ;
  assign MUX_m_vrg_source_busy_1$write_1__SEL_2 =
	     WILL_FIRE_RL_m_rl_process_rd_req && max_id__h24210 == 5'd1 &&
	     NOT_m_slave_xactor_f_rd_addr_first__9_BITS_92__ETC___d695 ;
  assign MUX_m_vrg_source_busy_10$write_1__SEL_1 =
	     WILL_FIRE_RL_m_rl_process_wr_req &&
	     wdata32__h27246[9:0] == 10'd10 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2884 ;
  assign MUX_m_vrg_source_busy_10$write_1__SEL_2 =
	     WILL_FIRE_RL_m_rl_process_rd_req && max_id__h24210 == 5'd10 &&
	     NOT_m_slave_xactor_f_rd_addr_first__9_BITS_92__ETC___d695 ;
  assign MUX_m_vrg_source_busy_11$write_1__SEL_1 =
	     WILL_FIRE_RL_m_rl_process_wr_req &&
	     wdata32__h27246[9:0] == 10'd11 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2884 ;
  assign MUX_m_vrg_source_busy_11$write_1__SEL_2 =
	     WILL_FIRE_RL_m_rl_process_rd_req && max_id__h24210 == 5'd11 &&
	     NOT_m_slave_xactor_f_rd_addr_first__9_BITS_92__ETC___d695 ;
  assign MUX_m_vrg_source_busy_12$write_1__SEL_1 =
	     WILL_FIRE_RL_m_rl_process_wr_req &&
	     wdata32__h27246[9:0] == 10'd12 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2884 ;
  assign MUX_m_vrg_source_busy_12$write_1__SEL_2 =
	     WILL_FIRE_RL_m_rl_process_rd_req && max_id__h24210 == 5'd12 &&
	     NOT_m_slave_xactor_f_rd_addr_first__9_BITS_92__ETC___d695 ;
  assign MUX_m_vrg_source_busy_13$write_1__SEL_1 =
	     WILL_FIRE_RL_m_rl_process_wr_req &&
	     wdata32__h27246[9:0] == 10'd13 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2884 ;
  assign MUX_m_vrg_source_busy_13$write_1__SEL_2 =
	     WILL_FIRE_RL_m_rl_process_rd_req && max_id__h24210 == 5'd13 &&
	     NOT_m_slave_xactor_f_rd_addr_first__9_BITS_92__ETC___d695 ;
  assign MUX_m_vrg_source_busy_14$write_1__SEL_1 =
	     WILL_FIRE_RL_m_rl_process_wr_req &&
	     wdata32__h27246[9:0] == 10'd14 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2884 ;
  assign MUX_m_vrg_source_busy_14$write_1__SEL_2 =
	     WILL_FIRE_RL_m_rl_process_rd_req && max_id__h24210 == 5'd14 &&
	     NOT_m_slave_xactor_f_rd_addr_first__9_BITS_92__ETC___d695 ;
  assign MUX_m_vrg_source_busy_15$write_1__SEL_1 =
	     WILL_FIRE_RL_m_rl_process_wr_req &&
	     wdata32__h27246[9:0] == 10'd15 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2884 ;
  assign MUX_m_vrg_source_busy_15$write_1__SEL_2 =
	     WILL_FIRE_RL_m_rl_process_rd_req && max_id__h24210 == 5'd15 &&
	     NOT_m_slave_xactor_f_rd_addr_first__9_BITS_92__ETC___d695 ;
  assign MUX_m_vrg_source_busy_16$write_1__SEL_1 =
	     WILL_FIRE_RL_m_rl_process_wr_req &&
	     wdata32__h27246[9:0] == 10'd16 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2884 ;
  assign MUX_m_vrg_source_busy_16$write_1__SEL_2 =
	     WILL_FIRE_RL_m_rl_process_rd_req && max_id__h24210 == 5'd16 &&
	     NOT_m_slave_xactor_f_rd_addr_first__9_BITS_92__ETC___d695 ;
  assign MUX_m_vrg_source_busy_2$write_1__SEL_1 =
	     WILL_FIRE_RL_m_rl_process_wr_req &&
	     wdata32__h27246[9:0] == 10'd2 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2884 ;
  assign MUX_m_vrg_source_busy_2$write_1__SEL_2 =
	     WILL_FIRE_RL_m_rl_process_rd_req && max_id__h24210 == 5'd2 &&
	     NOT_m_slave_xactor_f_rd_addr_first__9_BITS_92__ETC___d695 ;
  assign MUX_m_vrg_source_busy_3$write_1__SEL_1 =
	     WILL_FIRE_RL_m_rl_process_wr_req &&
	     wdata32__h27246[9:0] == 10'd3 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2884 ;
  assign MUX_m_vrg_source_busy_3$write_1__SEL_2 =
	     WILL_FIRE_RL_m_rl_process_rd_req && max_id__h24210 == 5'd3 &&
	     NOT_m_slave_xactor_f_rd_addr_first__9_BITS_92__ETC___d695 ;
  assign MUX_m_vrg_source_busy_4$write_1__SEL_1 =
	     WILL_FIRE_RL_m_rl_process_wr_req &&
	     wdata32__h27246[9:0] == 10'd4 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2884 ;
  assign MUX_m_vrg_source_busy_4$write_1__SEL_2 =
	     WILL_FIRE_RL_m_rl_process_rd_req && max_id__h24210 == 5'd4 &&
	     NOT_m_slave_xactor_f_rd_addr_first__9_BITS_92__ETC___d695 ;
  assign MUX_m_vrg_source_busy_5$write_1__SEL_1 =
	     WILL_FIRE_RL_m_rl_process_wr_req &&
	     wdata32__h27246[9:0] == 10'd5 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2884 ;
  assign MUX_m_vrg_source_busy_5$write_1__SEL_2 =
	     WILL_FIRE_RL_m_rl_process_rd_req && max_id__h24210 == 5'd5 &&
	     NOT_m_slave_xactor_f_rd_addr_first__9_BITS_92__ETC___d695 ;
  assign MUX_m_vrg_source_busy_6$write_1__SEL_1 =
	     WILL_FIRE_RL_m_rl_process_wr_req &&
	     wdata32__h27246[9:0] == 10'd6 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2884 ;
  assign MUX_m_vrg_source_busy_6$write_1__SEL_2 =
	     WILL_FIRE_RL_m_rl_process_rd_req && max_id__h24210 == 5'd6 &&
	     NOT_m_slave_xactor_f_rd_addr_first__9_BITS_92__ETC___d695 ;
  assign MUX_m_vrg_source_busy_7$write_1__SEL_1 =
	     WILL_FIRE_RL_m_rl_process_wr_req &&
	     wdata32__h27246[9:0] == 10'd7 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2884 ;
  assign MUX_m_vrg_source_busy_7$write_1__SEL_2 =
	     WILL_FIRE_RL_m_rl_process_rd_req && max_id__h24210 == 5'd7 &&
	     NOT_m_slave_xactor_f_rd_addr_first__9_BITS_92__ETC___d695 ;
  assign MUX_m_vrg_source_busy_8$write_1__SEL_1 =
	     WILL_FIRE_RL_m_rl_process_wr_req &&
	     wdata32__h27246[9:0] == 10'd8 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2884 ;
  assign MUX_m_vrg_source_busy_8$write_1__SEL_2 =
	     WILL_FIRE_RL_m_rl_process_rd_req && max_id__h24210 == 5'd8 &&
	     NOT_m_slave_xactor_f_rd_addr_first__9_BITS_92__ETC___d695 ;
  assign MUX_m_vrg_source_busy_9$write_1__SEL_1 =
	     WILL_FIRE_RL_m_rl_process_wr_req &&
	     wdata32__h27246[9:0] == 10'd9 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2884 ;
  assign MUX_m_vrg_source_busy_9$write_1__SEL_2 =
	     WILL_FIRE_RL_m_rl_process_rd_req && max_id__h24210 == 5'd9 &&
	     NOT_m_slave_xactor_f_rd_addr_first__9_BITS_92__ETC___d695 ;
  assign MUX_m_vrg_source_prio_0$write_1__SEL_1 =
	     WILL_FIRE_RL_m_rl_process_wr_req &&
	     addr_offset__h27245[11:2] == 10'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d826 ;
  assign MUX_m_vrg_source_prio_1$write_1__SEL_1 =
	     WILL_FIRE_RL_m_rl_process_wr_req &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d837 ;
  assign MUX_m_vrg_source_prio_10$write_1__SEL_1 =
	     WILL_FIRE_RL_m_rl_process_wr_req &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d855 ;
  assign MUX_m_vrg_source_prio_11$write_1__SEL_1 =
	     WILL_FIRE_RL_m_rl_process_wr_req &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d857 ;
  assign MUX_m_vrg_source_prio_12$write_1__SEL_1 =
	     WILL_FIRE_RL_m_rl_process_wr_req &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d859 ;
  assign MUX_m_vrg_source_prio_13$write_1__SEL_1 =
	     WILL_FIRE_RL_m_rl_process_wr_req &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d861 ;
  assign MUX_m_vrg_source_prio_14$write_1__SEL_1 =
	     WILL_FIRE_RL_m_rl_process_wr_req &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d863 ;
  assign MUX_m_vrg_source_prio_15$write_1__SEL_1 =
	     WILL_FIRE_RL_m_rl_process_wr_req &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d865 ;
  assign MUX_m_vrg_source_prio_16$write_1__SEL_1 =
	     WILL_FIRE_RL_m_rl_process_wr_req &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d867 ;
  assign MUX_m_vrg_source_prio_2$write_1__SEL_1 =
	     WILL_FIRE_RL_m_rl_process_wr_req &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d839 ;
  assign MUX_m_vrg_source_prio_3$write_1__SEL_1 =
	     WILL_FIRE_RL_m_rl_process_wr_req &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d841 ;
  assign MUX_m_vrg_source_prio_4$write_1__SEL_1 =
	     WILL_FIRE_RL_m_rl_process_wr_req &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d843 ;
  assign MUX_m_vrg_source_prio_5$write_1__SEL_1 =
	     WILL_FIRE_RL_m_rl_process_wr_req &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d845 ;
  assign MUX_m_vrg_source_prio_6$write_1__SEL_1 =
	     WILL_FIRE_RL_m_rl_process_wr_req &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d847 ;
  assign MUX_m_vrg_source_prio_7$write_1__SEL_1 =
	     WILL_FIRE_RL_m_rl_process_wr_req &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d849 ;
  assign MUX_m_vrg_source_prio_8$write_1__SEL_1 =
	     WILL_FIRE_RL_m_rl_process_wr_req &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d851 ;
  assign MUX_m_vrg_source_prio_9$write_1__SEL_1 =
	     WILL_FIRE_RL_m_rl_process_wr_req &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d853 ;
  assign MUX_m_vrg_target_threshold_0$write_1__SEL_1 =
	     WILL_FIRE_RL_m_rl_process_wr_req &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d2860 ;
  assign MUX_m_vrg_target_threshold_1$write_1__SEL_1 =
	     WILL_FIRE_RL_m_rl_process_wr_req &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d2862 ;
  assign MUX_m_vvrg_ie_0_0$write_1__SEL_1 =
	     WILL_FIRE_RL_m_rl_process_wr_req && _dfoo2107 ;
  assign MUX_m_vvrg_ie_0_1$write_1__SEL_1 =
	     WILL_FIRE_RL_m_rl_process_wr_req && _dfoo2105 ;
  assign MUX_m_vvrg_ie_0_10$write_1__SEL_1 =
	     WILL_FIRE_RL_m_rl_process_wr_req && _dfoo2087 ;
  assign MUX_m_vvrg_ie_0_11$write_1__SEL_1 =
	     WILL_FIRE_RL_m_rl_process_wr_req && _dfoo2085 ;
  assign MUX_m_vvrg_ie_0_12$write_1__SEL_1 =
	     WILL_FIRE_RL_m_rl_process_wr_req && _dfoo2083 ;
  assign MUX_m_vvrg_ie_0_13$write_1__SEL_1 =
	     WILL_FIRE_RL_m_rl_process_wr_req && _dfoo2081 ;
  assign MUX_m_vvrg_ie_0_14$write_1__SEL_1 =
	     WILL_FIRE_RL_m_rl_process_wr_req && _dfoo2079 ;
  assign MUX_m_vvrg_ie_0_15$write_1__SEL_1 =
	     WILL_FIRE_RL_m_rl_process_wr_req && _dfoo2077 ;
  assign MUX_m_vvrg_ie_0_16$write_1__SEL_1 =
	     WILL_FIRE_RL_m_rl_process_wr_req && _dfoo2075 ;
  assign MUX_m_vvrg_ie_0_2$write_1__SEL_1 =
	     WILL_FIRE_RL_m_rl_process_wr_req && _dfoo2103 ;
  assign MUX_m_vvrg_ie_0_3$write_1__SEL_1 =
	     WILL_FIRE_RL_m_rl_process_wr_req && _dfoo2101 ;
  assign MUX_m_vvrg_ie_0_4$write_1__SEL_1 =
	     WILL_FIRE_RL_m_rl_process_wr_req && _dfoo2099 ;
  assign MUX_m_vvrg_ie_0_5$write_1__SEL_1 =
	     WILL_FIRE_RL_m_rl_process_wr_req && _dfoo2097 ;
  assign MUX_m_vvrg_ie_0_6$write_1__SEL_1 =
	     WILL_FIRE_RL_m_rl_process_wr_req && _dfoo2095 ;
  assign MUX_m_vvrg_ie_0_7$write_1__SEL_1 =
	     WILL_FIRE_RL_m_rl_process_wr_req && _dfoo2093 ;
  assign MUX_m_vvrg_ie_0_8$write_1__SEL_1 =
	     WILL_FIRE_RL_m_rl_process_wr_req && _dfoo2091 ;
  assign MUX_m_vvrg_ie_0_9$write_1__SEL_1 =
	     WILL_FIRE_RL_m_rl_process_wr_req && _dfoo2089 ;
  assign MUX_m_vvrg_ie_1_0$write_1__SEL_1 =
	     WILL_FIRE_RL_m_rl_process_wr_req && _dfoo2073 ;
  assign MUX_m_vvrg_ie_1_1$write_1__SEL_1 =
	     WILL_FIRE_RL_m_rl_process_wr_req && _dfoo2071 ;
  assign MUX_m_vvrg_ie_1_10$write_1__SEL_1 =
	     WILL_FIRE_RL_m_rl_process_wr_req && _dfoo2053 ;
  assign MUX_m_vvrg_ie_1_11$write_1__SEL_1 =
	     WILL_FIRE_RL_m_rl_process_wr_req && _dfoo2051 ;
  assign MUX_m_vvrg_ie_1_12$write_1__SEL_1 =
	     WILL_FIRE_RL_m_rl_process_wr_req && _dfoo2049 ;
  assign MUX_m_vvrg_ie_1_13$write_1__SEL_1 =
	     WILL_FIRE_RL_m_rl_process_wr_req && _dfoo2047 ;
  assign MUX_m_vvrg_ie_1_14$write_1__SEL_1 =
	     WILL_FIRE_RL_m_rl_process_wr_req && _dfoo2045 ;
  assign MUX_m_vvrg_ie_1_15$write_1__SEL_1 =
	     WILL_FIRE_RL_m_rl_process_wr_req && _dfoo2043 ;
  assign MUX_m_vvrg_ie_1_16$write_1__SEL_1 =
	     WILL_FIRE_RL_m_rl_process_wr_req && _dfoo2041 ;
  assign MUX_m_vvrg_ie_1_2$write_1__SEL_1 =
	     WILL_FIRE_RL_m_rl_process_wr_req && _dfoo2069 ;
  assign MUX_m_vvrg_ie_1_3$write_1__SEL_1 =
	     WILL_FIRE_RL_m_rl_process_wr_req && _dfoo2067 ;
  assign MUX_m_vvrg_ie_1_4$write_1__SEL_1 =
	     WILL_FIRE_RL_m_rl_process_wr_req && _dfoo2065 ;
  assign MUX_m_vvrg_ie_1_5$write_1__SEL_1 =
	     WILL_FIRE_RL_m_rl_process_wr_req && _dfoo2063 ;
  assign MUX_m_vvrg_ie_1_6$write_1__SEL_1 =
	     WILL_FIRE_RL_m_rl_process_wr_req && _dfoo2061 ;
  assign MUX_m_vvrg_ie_1_7$write_1__SEL_1 =
	     WILL_FIRE_RL_m_rl_process_wr_req && _dfoo2059 ;
  assign MUX_m_vvrg_ie_1_8$write_1__SEL_1 =
	     WILL_FIRE_RL_m_rl_process_wr_req && _dfoo2057 ;
  assign MUX_m_vvrg_ie_1_9$write_1__SEL_1 =
	     WILL_FIRE_RL_m_rl_process_wr_req && _dfoo2055 ;
  assign MUX_m_vvrg_ie_0_0$write_1__VAL_1 =
	     (source_id_base__h28620 == 10'd0 &&
	      m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d895) ?
	       wdata32__h27246[0] :
	       _dfoo2040 ;
  assign MUX_m_vvrg_ie_0_1$write_1__VAL_1 =
	     (source_id_base__h28620 == 10'd1 &&
	      m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d895) ?
	       wdata32__h27246[0] :
	       _dfoo2038 ;
  assign MUX_m_vvrg_ie_0_10$write_1__VAL_1 =
	     (source_id_base__h28620 == 10'd10 &&
	      m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d895) ?
	       wdata32__h27246[0] :
	       _dfoo2020 ;
  assign MUX_m_vvrg_ie_0_11$write_1__VAL_1 =
	     (source_id_base__h28620 == 10'd11 &&
	      m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d895) ?
	       wdata32__h27246[0] :
	       _dfoo2018 ;
  assign MUX_m_vvrg_ie_0_12$write_1__VAL_1 =
	     (source_id_base__h28620 == 10'd12 &&
	      m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d895) ?
	       wdata32__h27246[0] :
	       _dfoo2016 ;
  assign MUX_m_vvrg_ie_0_13$write_1__VAL_1 =
	     (source_id_base__h28620 == 10'd13 &&
	      m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d895) ?
	       wdata32__h27246[0] :
	       _dfoo2014 ;
  assign MUX_m_vvrg_ie_0_14$write_1__VAL_1 =
	     (source_id_base__h28620 == 10'd14 &&
	      m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d895) ?
	       wdata32__h27246[0] :
	       _dfoo2012 ;
  assign MUX_m_vvrg_ie_0_15$write_1__VAL_1 =
	     (source_id_base__h28620 == 10'd15 &&
	      m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d895) ?
	       wdata32__h27246[0] :
	       _dfoo2010 ;
  assign MUX_m_vvrg_ie_0_16$write_1__VAL_1 =
	     (source_id_base__h28620 == 10'd16 &&
	      m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d895) ?
	       wdata32__h27246[0] :
	       _dfoo2008 ;
  assign MUX_m_vvrg_ie_0_2$write_1__VAL_1 =
	     (source_id_base__h28620 == 10'd2 &&
	      m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d895) ?
	       wdata32__h27246[0] :
	       _dfoo2036 ;
  assign MUX_m_vvrg_ie_0_3$write_1__VAL_1 =
	     (source_id_base__h28620 == 10'd3 &&
	      m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d895) ?
	       wdata32__h27246[0] :
	       _dfoo2034 ;
  assign MUX_m_vvrg_ie_0_4$write_1__VAL_1 =
	     (source_id_base__h28620 == 10'd4 &&
	      m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d895) ?
	       wdata32__h27246[0] :
	       _dfoo2032 ;
  assign MUX_m_vvrg_ie_0_5$write_1__VAL_1 =
	     (source_id_base__h28620 == 10'd5 &&
	      m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d895) ?
	       wdata32__h27246[0] :
	       _dfoo2030 ;
  assign MUX_m_vvrg_ie_0_6$write_1__VAL_1 =
	     (source_id_base__h28620 == 10'd6 &&
	      m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d895) ?
	       wdata32__h27246[0] :
	       _dfoo2028 ;
  assign MUX_m_vvrg_ie_0_7$write_1__VAL_1 =
	     (source_id_base__h28620 == 10'd7 &&
	      m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d895) ?
	       wdata32__h27246[0] :
	       _dfoo2026 ;
  assign MUX_m_vvrg_ie_0_8$write_1__VAL_1 =
	     (source_id_base__h28620 == 10'd8 &&
	      m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d895) ?
	       wdata32__h27246[0] :
	       _dfoo2024 ;
  assign MUX_m_vvrg_ie_0_9$write_1__VAL_1 =
	     (source_id_base__h28620 == 10'd9 &&
	      m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d895) ?
	       wdata32__h27246[0] :
	       _dfoo2022 ;
  assign MUX_m_vvrg_ie_1_0$write_1__VAL_1 =
	     (source_id_base__h28620 == 10'd0 &&
	      m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d931) ?
	       wdata32__h27246[0] :
	       _dfoo2006 ;
  assign MUX_m_vvrg_ie_1_1$write_1__VAL_1 =
	     (source_id_base__h28620 == 10'd1 &&
	      m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d931) ?
	       wdata32__h27246[0] :
	       _dfoo2004 ;
  assign MUX_m_vvrg_ie_1_10$write_1__VAL_1 =
	     (source_id_base__h28620 == 10'd10 &&
	      m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d931) ?
	       wdata32__h27246[0] :
	       _dfoo1986 ;
  assign MUX_m_vvrg_ie_1_11$write_1__VAL_1 =
	     (source_id_base__h28620 == 10'd11 &&
	      m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d931) ?
	       wdata32__h27246[0] :
	       _dfoo1984 ;
  assign MUX_m_vvrg_ie_1_12$write_1__VAL_1 =
	     (source_id_base__h28620 == 10'd12 &&
	      m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d931) ?
	       wdata32__h27246[0] :
	       _dfoo1982 ;
  assign MUX_m_vvrg_ie_1_13$write_1__VAL_1 =
	     (source_id_base__h28620 == 10'd13 &&
	      m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d931) ?
	       wdata32__h27246[0] :
	       _dfoo1980 ;
  assign MUX_m_vvrg_ie_1_14$write_1__VAL_1 =
	     (source_id_base__h28620 == 10'd14 &&
	      m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d931) ?
	       wdata32__h27246[0] :
	       _dfoo1978 ;
  assign MUX_m_vvrg_ie_1_15$write_1__VAL_1 =
	     (source_id_base__h28620 == 10'd15 &&
	      m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d931) ?
	       wdata32__h27246[0] :
	       _dfoo1976 ;
  assign MUX_m_vvrg_ie_1_16$write_1__VAL_1 =
	     (source_id_base__h28620 == 10'd16 &&
	      m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d931) ?
	       wdata32__h27246[0] :
	       _dfoo1974 ;
  assign MUX_m_vvrg_ie_1_2$write_1__VAL_1 =
	     (source_id_base__h28620 == 10'd2 &&
	      m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d931) ?
	       wdata32__h27246[0] :
	       _dfoo2002 ;
  assign MUX_m_vvrg_ie_1_3$write_1__VAL_1 =
	     (source_id_base__h28620 == 10'd3 &&
	      m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d931) ?
	       wdata32__h27246[0] :
	       _dfoo2000 ;
  assign MUX_m_vvrg_ie_1_4$write_1__VAL_1 =
	     (source_id_base__h28620 == 10'd4 &&
	      m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d931) ?
	       wdata32__h27246[0] :
	       _dfoo1998 ;
  assign MUX_m_vvrg_ie_1_5$write_1__VAL_1 =
	     (source_id_base__h28620 == 10'd5 &&
	      m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d931) ?
	       wdata32__h27246[0] :
	       _dfoo1996 ;
  assign MUX_m_vvrg_ie_1_6$write_1__VAL_1 =
	     (source_id_base__h28620 == 10'd6 &&
	      m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d931) ?
	       wdata32__h27246[0] :
	       _dfoo1994 ;
  assign MUX_m_vvrg_ie_1_7$write_1__VAL_1 =
	     (source_id_base__h28620 == 10'd7 &&
	      m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d931) ?
	       wdata32__h27246[0] :
	       _dfoo1992 ;
  assign MUX_m_vvrg_ie_1_8$write_1__VAL_1 =
	     (source_id_base__h28620 == 10'd8 &&
	      m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d931) ?
	       wdata32__h27246[0] :
	       _dfoo1990 ;
  assign MUX_m_vvrg_ie_1_9$write_1__VAL_1 =
	     (source_id_base__h28620 == 10'd9 &&
	      m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d931) ?
	       wdata32__h27246[0] :
	       _dfoo1988 ;
  // register m_cfg_verbosity
  assign m_cfg_verbosity$D_IN = set_verbosity_verbosity ;
  assign m_cfg_verbosity$EN = EN_set_verbosity ;
  // register m_rg_addr_base
  assign m_rg_addr_base$D_IN = set_addr_map_addr_base ;
  assign m_rg_addr_base$EN = EN_set_addr_map ;
  // register m_rg_addr_lim
  assign m_rg_addr_lim$D_IN = set_addr_map_addr_lim ;
  assign m_rg_addr_lim$EN = EN_set_addr_map ;
  // register m_vrg_source_busy_0
  always@(MUX_m_vrg_source_busy_0$write_1__SEL_1 or
	  MUX_m_vrg_source_busy_0$write_1__SEL_2 or WILL_FIRE_RL_m_rl_reset)
  case (1'b1)
    MUX_m_vrg_source_busy_0$write_1__SEL_1: m_vrg_source_busy_0$D_IN = 1'd0;
    MUX_m_vrg_source_busy_0$write_1__SEL_2: m_vrg_source_busy_0$D_IN = 1'd1;
    WILL_FIRE_RL_m_rl_reset: m_vrg_source_busy_0$D_IN = 1'd0;
    default: m_vrg_source_busy_0$D_IN = 1'b0 /* unspecified value */ ;
  endcase
  assign m_vrg_source_busy_0$EN =
	     WILL_FIRE_RL_m_rl_process_rd_req && max_id__h24210 == 5'd0 &&
	     NOT_m_slave_xactor_f_rd_addr_first__9_BITS_92__ETC___d695 ||
	     WILL_FIRE_RL_m_rl_process_wr_req &&
	     wdata32__h27246[9:0] == 10'd0 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2884 ||
	     WILL_FIRE_RL_m_rl_reset ;
  // register m_vrg_source_busy_1
  always@(MUX_m_vrg_source_busy_1$write_1__SEL_1 or
	  MUX_m_vrg_source_busy_1$write_1__SEL_2 or WILL_FIRE_RL_m_rl_reset)
  case (1'b1)
    MUX_m_vrg_source_busy_1$write_1__SEL_1: m_vrg_source_busy_1$D_IN = 1'd0;
    MUX_m_vrg_source_busy_1$write_1__SEL_2: m_vrg_source_busy_1$D_IN = 1'd1;
    WILL_FIRE_RL_m_rl_reset: m_vrg_source_busy_1$D_IN = 1'd0;
    default: m_vrg_source_busy_1$D_IN = 1'b0 /* unspecified value */ ;
  endcase
  assign m_vrg_source_busy_1$EN =
	     WILL_FIRE_RL_m_rl_process_rd_req && max_id__h24210 == 5'd1 &&
	     NOT_m_slave_xactor_f_rd_addr_first__9_BITS_92__ETC___d695 ||
	     WILL_FIRE_RL_m_rl_process_wr_req &&
	     wdata32__h27246[9:0] == 10'd1 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2884 ||
	     WILL_FIRE_RL_m_rl_reset ;
  // register m_vrg_source_busy_10
  always@(MUX_m_vrg_source_busy_10$write_1__SEL_1 or
	  MUX_m_vrg_source_busy_10$write_1__SEL_2 or WILL_FIRE_RL_m_rl_reset)
  case (1'b1)
    MUX_m_vrg_source_busy_10$write_1__SEL_1: m_vrg_source_busy_10$D_IN = 1'd0;
    MUX_m_vrg_source_busy_10$write_1__SEL_2: m_vrg_source_busy_10$D_IN = 1'd1;
    WILL_FIRE_RL_m_rl_reset: m_vrg_source_busy_10$D_IN = 1'd0;
    default: m_vrg_source_busy_10$D_IN = 1'b0 /* unspecified value */ ;
  endcase
  assign m_vrg_source_busy_10$EN =
	     WILL_FIRE_RL_m_rl_process_rd_req && max_id__h24210 == 5'd10 &&
	     NOT_m_slave_xactor_f_rd_addr_first__9_BITS_92__ETC___d695 ||
	     WILL_FIRE_RL_m_rl_process_wr_req &&
	     wdata32__h27246[9:0] == 10'd10 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2884 ||
	     WILL_FIRE_RL_m_rl_reset ;
  // register m_vrg_source_busy_11
  always@(MUX_m_vrg_source_busy_11$write_1__SEL_1 or
	  MUX_m_vrg_source_busy_11$write_1__SEL_2 or WILL_FIRE_RL_m_rl_reset)
  case (1'b1)
    MUX_m_vrg_source_busy_11$write_1__SEL_1: m_vrg_source_busy_11$D_IN = 1'd0;
    MUX_m_vrg_source_busy_11$write_1__SEL_2: m_vrg_source_busy_11$D_IN = 1'd1;
    WILL_FIRE_RL_m_rl_reset: m_vrg_source_busy_11$D_IN = 1'd0;
    default: m_vrg_source_busy_11$D_IN = 1'b0 /* unspecified value */ ;
  endcase
  assign m_vrg_source_busy_11$EN =
	     WILL_FIRE_RL_m_rl_process_rd_req && max_id__h24210 == 5'd11 &&
	     NOT_m_slave_xactor_f_rd_addr_first__9_BITS_92__ETC___d695 ||
	     WILL_FIRE_RL_m_rl_process_wr_req &&
	     wdata32__h27246[9:0] == 10'd11 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2884 ||
	     WILL_FIRE_RL_m_rl_reset ;
  // register m_vrg_source_busy_12
  always@(MUX_m_vrg_source_busy_12$write_1__SEL_1 or
	  MUX_m_vrg_source_busy_12$write_1__SEL_2 or WILL_FIRE_RL_m_rl_reset)
  case (1'b1)
    MUX_m_vrg_source_busy_12$write_1__SEL_1: m_vrg_source_busy_12$D_IN = 1'd0;
    MUX_m_vrg_source_busy_12$write_1__SEL_2: m_vrg_source_busy_12$D_IN = 1'd1;
    WILL_FIRE_RL_m_rl_reset: m_vrg_source_busy_12$D_IN = 1'd0;
    default: m_vrg_source_busy_12$D_IN = 1'b0 /* unspecified value */ ;
  endcase
  assign m_vrg_source_busy_12$EN =
	     WILL_FIRE_RL_m_rl_process_rd_req && max_id__h24210 == 5'd12 &&
	     NOT_m_slave_xactor_f_rd_addr_first__9_BITS_92__ETC___d695 ||
	     WILL_FIRE_RL_m_rl_process_wr_req &&
	     wdata32__h27246[9:0] == 10'd12 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2884 ||
	     WILL_FIRE_RL_m_rl_reset ;
  // register m_vrg_source_busy_13
  always@(MUX_m_vrg_source_busy_13$write_1__SEL_1 or
	  MUX_m_vrg_source_busy_13$write_1__SEL_2 or WILL_FIRE_RL_m_rl_reset)
  case (1'b1)
    MUX_m_vrg_source_busy_13$write_1__SEL_1: m_vrg_source_busy_13$D_IN = 1'd0;
    MUX_m_vrg_source_busy_13$write_1__SEL_2: m_vrg_source_busy_13$D_IN = 1'd1;
    WILL_FIRE_RL_m_rl_reset: m_vrg_source_busy_13$D_IN = 1'd0;
    default: m_vrg_source_busy_13$D_IN = 1'b0 /* unspecified value */ ;
  endcase
  assign m_vrg_source_busy_13$EN =
	     WILL_FIRE_RL_m_rl_process_rd_req && max_id__h24210 == 5'd13 &&
	     NOT_m_slave_xactor_f_rd_addr_first__9_BITS_92__ETC___d695 ||
	     WILL_FIRE_RL_m_rl_process_wr_req &&
	     wdata32__h27246[9:0] == 10'd13 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2884 ||
	     WILL_FIRE_RL_m_rl_reset ;
  // register m_vrg_source_busy_14
  always@(MUX_m_vrg_source_busy_14$write_1__SEL_1 or
	  MUX_m_vrg_source_busy_14$write_1__SEL_2 or WILL_FIRE_RL_m_rl_reset)
  case (1'b1)
    MUX_m_vrg_source_busy_14$write_1__SEL_1: m_vrg_source_busy_14$D_IN = 1'd0;
    MUX_m_vrg_source_busy_14$write_1__SEL_2: m_vrg_source_busy_14$D_IN = 1'd1;
    WILL_FIRE_RL_m_rl_reset: m_vrg_source_busy_14$D_IN = 1'd0;
    default: m_vrg_source_busy_14$D_IN = 1'b0 /* unspecified value */ ;
  endcase
  assign m_vrg_source_busy_14$EN =
	     WILL_FIRE_RL_m_rl_process_rd_req && max_id__h24210 == 5'd14 &&
	     NOT_m_slave_xactor_f_rd_addr_first__9_BITS_92__ETC___d695 ||
	     WILL_FIRE_RL_m_rl_process_wr_req &&
	     wdata32__h27246[9:0] == 10'd14 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2884 ||
	     WILL_FIRE_RL_m_rl_reset ;
  // register m_vrg_source_busy_15
  always@(MUX_m_vrg_source_busy_15$write_1__SEL_1 or
	  MUX_m_vrg_source_busy_15$write_1__SEL_2 or WILL_FIRE_RL_m_rl_reset)
  case (1'b1)
    MUX_m_vrg_source_busy_15$write_1__SEL_1: m_vrg_source_busy_15$D_IN = 1'd0;
    MUX_m_vrg_source_busy_15$write_1__SEL_2: m_vrg_source_busy_15$D_IN = 1'd1;
    WILL_FIRE_RL_m_rl_reset: m_vrg_source_busy_15$D_IN = 1'd0;
    default: m_vrg_source_busy_15$D_IN = 1'b0 /* unspecified value */ ;
  endcase
  assign m_vrg_source_busy_15$EN =
	     WILL_FIRE_RL_m_rl_process_rd_req && max_id__h24210 == 5'd15 &&
	     NOT_m_slave_xactor_f_rd_addr_first__9_BITS_92__ETC___d695 ||
	     WILL_FIRE_RL_m_rl_process_wr_req &&
	     wdata32__h27246[9:0] == 10'd15 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2884 ||
	     WILL_FIRE_RL_m_rl_reset ;
  // register m_vrg_source_busy_16
  always@(MUX_m_vrg_source_busy_16$write_1__SEL_1 or
	  MUX_m_vrg_source_busy_16$write_1__SEL_2 or WILL_FIRE_RL_m_rl_reset)
  case (1'b1)
    MUX_m_vrg_source_busy_16$write_1__SEL_1: m_vrg_source_busy_16$D_IN = 1'd0;
    MUX_m_vrg_source_busy_16$write_1__SEL_2: m_vrg_source_busy_16$D_IN = 1'd1;
    WILL_FIRE_RL_m_rl_reset: m_vrg_source_busy_16$D_IN = 1'd0;
    default: m_vrg_source_busy_16$D_IN = 1'b0 /* unspecified value */ ;
  endcase
  assign m_vrg_source_busy_16$EN =
	     WILL_FIRE_RL_m_rl_process_rd_req && max_id__h24210 == 5'd16 &&
	     NOT_m_slave_xactor_f_rd_addr_first__9_BITS_92__ETC___d695 ||
	     WILL_FIRE_RL_m_rl_process_wr_req &&
	     wdata32__h27246[9:0] == 10'd16 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2884 ||
	     WILL_FIRE_RL_m_rl_reset ;
  // register m_vrg_source_busy_2
  always@(MUX_m_vrg_source_busy_2$write_1__SEL_1 or
	  MUX_m_vrg_source_busy_2$write_1__SEL_2 or WILL_FIRE_RL_m_rl_reset)
  case (1'b1)
    MUX_m_vrg_source_busy_2$write_1__SEL_1: m_vrg_source_busy_2$D_IN = 1'd0;
    MUX_m_vrg_source_busy_2$write_1__SEL_2: m_vrg_source_busy_2$D_IN = 1'd1;
    WILL_FIRE_RL_m_rl_reset: m_vrg_source_busy_2$D_IN = 1'd0;
    default: m_vrg_source_busy_2$D_IN = 1'b0 /* unspecified value */ ;
  endcase
  assign m_vrg_source_busy_2$EN =
	     WILL_FIRE_RL_m_rl_process_rd_req && max_id__h24210 == 5'd2 &&
	     NOT_m_slave_xactor_f_rd_addr_first__9_BITS_92__ETC___d695 ||
	     WILL_FIRE_RL_m_rl_process_wr_req &&
	     wdata32__h27246[9:0] == 10'd2 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2884 ||
	     WILL_FIRE_RL_m_rl_reset ;
  // register m_vrg_source_busy_3
  always@(MUX_m_vrg_source_busy_3$write_1__SEL_1 or
	  MUX_m_vrg_source_busy_3$write_1__SEL_2 or WILL_FIRE_RL_m_rl_reset)
  case (1'b1)
    MUX_m_vrg_source_busy_3$write_1__SEL_1: m_vrg_source_busy_3$D_IN = 1'd0;
    MUX_m_vrg_source_busy_3$write_1__SEL_2: m_vrg_source_busy_3$D_IN = 1'd1;
    WILL_FIRE_RL_m_rl_reset: m_vrg_source_busy_3$D_IN = 1'd0;
    default: m_vrg_source_busy_3$D_IN = 1'b0 /* unspecified value */ ;
  endcase
  assign m_vrg_source_busy_3$EN =
	     WILL_FIRE_RL_m_rl_process_rd_req && max_id__h24210 == 5'd3 &&
	     NOT_m_slave_xactor_f_rd_addr_first__9_BITS_92__ETC___d695 ||
	     WILL_FIRE_RL_m_rl_process_wr_req &&
	     wdata32__h27246[9:0] == 10'd3 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2884 ||
	     WILL_FIRE_RL_m_rl_reset ;
  // register m_vrg_source_busy_4
  always@(MUX_m_vrg_source_busy_4$write_1__SEL_1 or
	  MUX_m_vrg_source_busy_4$write_1__SEL_2 or WILL_FIRE_RL_m_rl_reset)
  case (1'b1)
    MUX_m_vrg_source_busy_4$write_1__SEL_1: m_vrg_source_busy_4$D_IN = 1'd0;
    MUX_m_vrg_source_busy_4$write_1__SEL_2: m_vrg_source_busy_4$D_IN = 1'd1;
    WILL_FIRE_RL_m_rl_reset: m_vrg_source_busy_4$D_IN = 1'd0;
    default: m_vrg_source_busy_4$D_IN = 1'b0 /* unspecified value */ ;
  endcase
  assign m_vrg_source_busy_4$EN =
	     WILL_FIRE_RL_m_rl_process_rd_req && max_id__h24210 == 5'd4 &&
	     NOT_m_slave_xactor_f_rd_addr_first__9_BITS_92__ETC___d695 ||
	     WILL_FIRE_RL_m_rl_process_wr_req &&
	     wdata32__h27246[9:0] == 10'd4 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2884 ||
	     WILL_FIRE_RL_m_rl_reset ;
  // register m_vrg_source_busy_5
  always@(MUX_m_vrg_source_busy_5$write_1__SEL_1 or
	  MUX_m_vrg_source_busy_5$write_1__SEL_2 or WILL_FIRE_RL_m_rl_reset)
  case (1'b1)
    MUX_m_vrg_source_busy_5$write_1__SEL_1: m_vrg_source_busy_5$D_IN = 1'd0;
    MUX_m_vrg_source_busy_5$write_1__SEL_2: m_vrg_source_busy_5$D_IN = 1'd1;
    WILL_FIRE_RL_m_rl_reset: m_vrg_source_busy_5$D_IN = 1'd0;
    default: m_vrg_source_busy_5$D_IN = 1'b0 /* unspecified value */ ;
  endcase
  assign m_vrg_source_busy_5$EN =
	     WILL_FIRE_RL_m_rl_process_rd_req && max_id__h24210 == 5'd5 &&
	     NOT_m_slave_xactor_f_rd_addr_first__9_BITS_92__ETC___d695 ||
	     WILL_FIRE_RL_m_rl_process_wr_req &&
	     wdata32__h27246[9:0] == 10'd5 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2884 ||
	     WILL_FIRE_RL_m_rl_reset ;
  // register m_vrg_source_busy_6
  always@(MUX_m_vrg_source_busy_6$write_1__SEL_1 or
	  MUX_m_vrg_source_busy_6$write_1__SEL_2 or WILL_FIRE_RL_m_rl_reset)
  case (1'b1)
    MUX_m_vrg_source_busy_6$write_1__SEL_1: m_vrg_source_busy_6$D_IN = 1'd0;
    MUX_m_vrg_source_busy_6$write_1__SEL_2: m_vrg_source_busy_6$D_IN = 1'd1;
    WILL_FIRE_RL_m_rl_reset: m_vrg_source_busy_6$D_IN = 1'd0;
    default: m_vrg_source_busy_6$D_IN = 1'b0 /* unspecified value */ ;
  endcase
  assign m_vrg_source_busy_6$EN =
	     WILL_FIRE_RL_m_rl_process_rd_req && max_id__h24210 == 5'd6 &&
	     NOT_m_slave_xactor_f_rd_addr_first__9_BITS_92__ETC___d695 ||
	     WILL_FIRE_RL_m_rl_process_wr_req &&
	     wdata32__h27246[9:0] == 10'd6 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2884 ||
	     WILL_FIRE_RL_m_rl_reset ;
  // register m_vrg_source_busy_7
  always@(MUX_m_vrg_source_busy_7$write_1__SEL_1 or
	  MUX_m_vrg_source_busy_7$write_1__SEL_2 or WILL_FIRE_RL_m_rl_reset)
  case (1'b1)
    MUX_m_vrg_source_busy_7$write_1__SEL_1: m_vrg_source_busy_7$D_IN = 1'd0;
    MUX_m_vrg_source_busy_7$write_1__SEL_2: m_vrg_source_busy_7$D_IN = 1'd1;
    WILL_FIRE_RL_m_rl_reset: m_vrg_source_busy_7$D_IN = 1'd0;
    default: m_vrg_source_busy_7$D_IN = 1'b0 /* unspecified value */ ;
  endcase
  assign m_vrg_source_busy_7$EN =
	     WILL_FIRE_RL_m_rl_process_rd_req && max_id__h24210 == 5'd7 &&
	     NOT_m_slave_xactor_f_rd_addr_first__9_BITS_92__ETC___d695 ||
	     WILL_FIRE_RL_m_rl_process_wr_req &&
	     wdata32__h27246[9:0] == 10'd7 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2884 ||
	     WILL_FIRE_RL_m_rl_reset ;
  // register m_vrg_source_busy_8
  always@(MUX_m_vrg_source_busy_8$write_1__SEL_1 or
	  MUX_m_vrg_source_busy_8$write_1__SEL_2 or WILL_FIRE_RL_m_rl_reset)
  case (1'b1)
    MUX_m_vrg_source_busy_8$write_1__SEL_1: m_vrg_source_busy_8$D_IN = 1'd0;
    MUX_m_vrg_source_busy_8$write_1__SEL_2: m_vrg_source_busy_8$D_IN = 1'd1;
    WILL_FIRE_RL_m_rl_reset: m_vrg_source_busy_8$D_IN = 1'd0;
    default: m_vrg_source_busy_8$D_IN = 1'b0 /* unspecified value */ ;
  endcase
  assign m_vrg_source_busy_8$EN =
	     WILL_FIRE_RL_m_rl_process_rd_req && max_id__h24210 == 5'd8 &&
	     NOT_m_slave_xactor_f_rd_addr_first__9_BITS_92__ETC___d695 ||
	     WILL_FIRE_RL_m_rl_process_wr_req &&
	     wdata32__h27246[9:0] == 10'd8 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2884 ||
	     WILL_FIRE_RL_m_rl_reset ;
  // register m_vrg_source_busy_9
  always@(MUX_m_vrg_source_busy_9$write_1__SEL_1 or
	  MUX_m_vrg_source_busy_9$write_1__SEL_2 or WILL_FIRE_RL_m_rl_reset)
  case (1'b1)
    MUX_m_vrg_source_busy_9$write_1__SEL_1: m_vrg_source_busy_9$D_IN = 1'd0;
    MUX_m_vrg_source_busy_9$write_1__SEL_2: m_vrg_source_busy_9$D_IN = 1'd1;
    WILL_FIRE_RL_m_rl_reset: m_vrg_source_busy_9$D_IN = 1'd0;
    default: m_vrg_source_busy_9$D_IN = 1'b0 /* unspecified value */ ;
  endcase
  assign m_vrg_source_busy_9$EN =
	     WILL_FIRE_RL_m_rl_process_rd_req && max_id__h24210 == 5'd9 &&
	     NOT_m_slave_xactor_f_rd_addr_first__9_BITS_92__ETC___d695 ||
	     WILL_FIRE_RL_m_rl_process_wr_req &&
	     wdata32__h27246[9:0] == 10'd9 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2884 ||
	     WILL_FIRE_RL_m_rl_reset ;
  // register m_vrg_source_ip_0
  assign m_vrg_source_ip_0$D_IN = 1'd0 ;
  assign m_vrg_source_ip_0$EN =
	     WILL_FIRE_RL_m_rl_process_rd_req && max_id__h24210 == 5'd0 &&
	     NOT_m_slave_xactor_f_rd_addr_first__9_BITS_92__ETC___d695 ||
	     WILL_FIRE_RL_m_rl_reset ;
  // register m_vrg_source_ip_1
  assign m_vrg_source_ip_1$D_IN =
	     !MUX_m_vrg_source_busy_1$write_1__SEL_2 &&
	     !WILL_FIRE_RL_m_rl_reset &&
	     v_sources_0_m_interrupt_req_set_not_clear ;
  assign m_vrg_source_ip_1$EN =
	     !m_vrg_source_busy_1 ||
	     WILL_FIRE_RL_m_rl_process_rd_req && max_id__h24210 == 5'd1 &&
	     NOT_m_slave_xactor_f_rd_addr_first__9_BITS_92__ETC___d695 ||
	     WILL_FIRE_RL_m_rl_reset ;
  // register m_vrg_source_ip_10
  assign m_vrg_source_ip_10$D_IN =
	     !MUX_m_vrg_source_busy_10$write_1__SEL_2 &&
	     !WILL_FIRE_RL_m_rl_reset &&
	     v_sources_9_m_interrupt_req_set_not_clear ;
  assign m_vrg_source_ip_10$EN =
	     !m_vrg_source_busy_10 ||
	     WILL_FIRE_RL_m_rl_process_rd_req && max_id__h24210 == 5'd10 &&
	     NOT_m_slave_xactor_f_rd_addr_first__9_BITS_92__ETC___d695 ||
	     WILL_FIRE_RL_m_rl_reset ;
  // register m_vrg_source_ip_11
  assign m_vrg_source_ip_11$D_IN =
	     !MUX_m_vrg_source_busy_11$write_1__SEL_2 &&
	     !WILL_FIRE_RL_m_rl_reset &&
	     v_sources_10_m_interrupt_req_set_not_clear ;
  assign m_vrg_source_ip_11$EN =
	     !m_vrg_source_busy_11 ||
	     WILL_FIRE_RL_m_rl_process_rd_req && max_id__h24210 == 5'd11 &&
	     NOT_m_slave_xactor_f_rd_addr_first__9_BITS_92__ETC___d695 ||
	     WILL_FIRE_RL_m_rl_reset ;
  // register m_vrg_source_ip_12
  assign m_vrg_source_ip_12$D_IN =
	     !MUX_m_vrg_source_busy_12$write_1__SEL_2 &&
	     !WILL_FIRE_RL_m_rl_reset &&
	     v_sources_11_m_interrupt_req_set_not_clear ;
  assign m_vrg_source_ip_12$EN =
	     !m_vrg_source_busy_12 ||
	     WILL_FIRE_RL_m_rl_process_rd_req && max_id__h24210 == 5'd12 &&
	     NOT_m_slave_xactor_f_rd_addr_first__9_BITS_92__ETC___d695 ||
	     WILL_FIRE_RL_m_rl_reset ;
  // register m_vrg_source_ip_13
  assign m_vrg_source_ip_13$D_IN =
	     !MUX_m_vrg_source_busy_13$write_1__SEL_2 &&
	     !WILL_FIRE_RL_m_rl_reset &&
	     v_sources_12_m_interrupt_req_set_not_clear ;
  assign m_vrg_source_ip_13$EN =
	     !m_vrg_source_busy_13 ||
	     WILL_FIRE_RL_m_rl_process_rd_req && max_id__h24210 == 5'd13 &&
	     NOT_m_slave_xactor_f_rd_addr_first__9_BITS_92__ETC___d695 ||
	     WILL_FIRE_RL_m_rl_reset ;
  // register m_vrg_source_ip_14
  assign m_vrg_source_ip_14$D_IN =
	     !MUX_m_vrg_source_busy_14$write_1__SEL_2 &&
	     !WILL_FIRE_RL_m_rl_reset &&
	     v_sources_13_m_interrupt_req_set_not_clear ;
  assign m_vrg_source_ip_14$EN =
	     !m_vrg_source_busy_14 ||
	     WILL_FIRE_RL_m_rl_process_rd_req && max_id__h24210 == 5'd14 &&
	     NOT_m_slave_xactor_f_rd_addr_first__9_BITS_92__ETC___d695 ||
	     WILL_FIRE_RL_m_rl_reset ;
  // register m_vrg_source_ip_15
  assign m_vrg_source_ip_15$D_IN =
	     !MUX_m_vrg_source_busy_15$write_1__SEL_2 &&
	     !WILL_FIRE_RL_m_rl_reset &&
	     v_sources_14_m_interrupt_req_set_not_clear ;
  assign m_vrg_source_ip_15$EN =
	     !m_vrg_source_busy_15 ||
	     WILL_FIRE_RL_m_rl_process_rd_req && max_id__h24210 == 5'd15 &&
	     NOT_m_slave_xactor_f_rd_addr_first__9_BITS_92__ETC___d695 ||
	     WILL_FIRE_RL_m_rl_reset ;
  // register m_vrg_source_ip_16
  assign m_vrg_source_ip_16$D_IN =
	     !MUX_m_vrg_source_busy_16$write_1__SEL_2 &&
	     !WILL_FIRE_RL_m_rl_reset &&
	     v_sources_15_m_interrupt_req_set_not_clear ;
  assign m_vrg_source_ip_16$EN =
	     !m_vrg_source_busy_16 ||
	     WILL_FIRE_RL_m_rl_process_rd_req && max_id__h24210 == 5'd16 &&
	     NOT_m_slave_xactor_f_rd_addr_first__9_BITS_92__ETC___d695 ||
	     WILL_FIRE_RL_m_rl_reset ;
  // register m_vrg_source_ip_2
  assign m_vrg_source_ip_2$D_IN =
	     !MUX_m_vrg_source_busy_2$write_1__SEL_2 &&
	     !WILL_FIRE_RL_m_rl_reset &&
	     v_sources_1_m_interrupt_req_set_not_clear ;
  assign m_vrg_source_ip_2$EN =
	     !m_vrg_source_busy_2 ||
	     WILL_FIRE_RL_m_rl_process_rd_req && max_id__h24210 == 5'd2 &&
	     NOT_m_slave_xactor_f_rd_addr_first__9_BITS_92__ETC___d695 ||
	     WILL_FIRE_RL_m_rl_reset ;
  // register m_vrg_source_ip_3
  assign m_vrg_source_ip_3$D_IN =
	     !MUX_m_vrg_source_busy_3$write_1__SEL_2 &&
	     !WILL_FIRE_RL_m_rl_reset &&
	     v_sources_2_m_interrupt_req_set_not_clear ;
  assign m_vrg_source_ip_3$EN =
	     !m_vrg_source_busy_3 ||
	     WILL_FIRE_RL_m_rl_process_rd_req && max_id__h24210 == 5'd3 &&
	     NOT_m_slave_xactor_f_rd_addr_first__9_BITS_92__ETC___d695 ||
	     WILL_FIRE_RL_m_rl_reset ;
  // register m_vrg_source_ip_4
  assign m_vrg_source_ip_4$D_IN =
	     !MUX_m_vrg_source_busy_4$write_1__SEL_2 &&
	     !WILL_FIRE_RL_m_rl_reset &&
	     v_sources_3_m_interrupt_req_set_not_clear ;
  assign m_vrg_source_ip_4$EN =
	     !m_vrg_source_busy_4 ||
	     WILL_FIRE_RL_m_rl_process_rd_req && max_id__h24210 == 5'd4 &&
	     NOT_m_slave_xactor_f_rd_addr_first__9_BITS_92__ETC___d695 ||
	     WILL_FIRE_RL_m_rl_reset ;
  // register m_vrg_source_ip_5
  assign m_vrg_source_ip_5$D_IN =
	     !MUX_m_vrg_source_busy_5$write_1__SEL_2 &&
	     !WILL_FIRE_RL_m_rl_reset &&
	     v_sources_4_m_interrupt_req_set_not_clear ;
  assign m_vrg_source_ip_5$EN =
	     !m_vrg_source_busy_5 ||
	     WILL_FIRE_RL_m_rl_process_rd_req && max_id__h24210 == 5'd5 &&
	     NOT_m_slave_xactor_f_rd_addr_first__9_BITS_92__ETC___d695 ||
	     WILL_FIRE_RL_m_rl_reset ;
  // register m_vrg_source_ip_6
  assign m_vrg_source_ip_6$D_IN =
	     !MUX_m_vrg_source_busy_6$write_1__SEL_2 &&
	     !WILL_FIRE_RL_m_rl_reset &&
	     v_sources_5_m_interrupt_req_set_not_clear ;
  assign m_vrg_source_ip_6$EN =
	     !m_vrg_source_busy_6 ||
	     WILL_FIRE_RL_m_rl_process_rd_req && max_id__h24210 == 5'd6 &&
	     NOT_m_slave_xactor_f_rd_addr_first__9_BITS_92__ETC___d695 ||
	     WILL_FIRE_RL_m_rl_reset ;
  // register m_vrg_source_ip_7
  assign m_vrg_source_ip_7$D_IN =
	     !MUX_m_vrg_source_busy_7$write_1__SEL_2 &&
	     !WILL_FIRE_RL_m_rl_reset &&
	     v_sources_6_m_interrupt_req_set_not_clear ;
  assign m_vrg_source_ip_7$EN =
	     !m_vrg_source_busy_7 ||
	     WILL_FIRE_RL_m_rl_process_rd_req && max_id__h24210 == 5'd7 &&
	     NOT_m_slave_xactor_f_rd_addr_first__9_BITS_92__ETC___d695 ||
	     WILL_FIRE_RL_m_rl_reset ;
  // register m_vrg_source_ip_8
  assign m_vrg_source_ip_8$D_IN =
	     !MUX_m_vrg_source_busy_8$write_1__SEL_2 &&
	     !WILL_FIRE_RL_m_rl_reset &&
	     v_sources_7_m_interrupt_req_set_not_clear ;
  assign m_vrg_source_ip_8$EN =
	     !m_vrg_source_busy_8 ||
	     WILL_FIRE_RL_m_rl_process_rd_req && max_id__h24210 == 5'd8 &&
	     NOT_m_slave_xactor_f_rd_addr_first__9_BITS_92__ETC___d695 ||
	     WILL_FIRE_RL_m_rl_reset ;
  // register m_vrg_source_ip_9
  assign m_vrg_source_ip_9$D_IN =
	     !MUX_m_vrg_source_busy_9$write_1__SEL_2 &&
	     !WILL_FIRE_RL_m_rl_reset &&
	     v_sources_8_m_interrupt_req_set_not_clear ;
  assign m_vrg_source_ip_9$EN =
	     !m_vrg_source_busy_9 ||
	     WILL_FIRE_RL_m_rl_process_rd_req && max_id__h24210 == 5'd9 &&
	     NOT_m_slave_xactor_f_rd_addr_first__9_BITS_92__ETC___d695 ||
	     WILL_FIRE_RL_m_rl_reset ;
  // register m_vrg_source_prio_0
  assign m_vrg_source_prio_0$D_IN =
	     MUX_m_vrg_source_prio_0$write_1__SEL_1 ?
	       wdata32__h27246[2:0] :
	       3'd0 ;
  assign m_vrg_source_prio_0$EN =
	     WILL_FIRE_RL_m_rl_process_wr_req &&
	     addr_offset__h27245[11:2] == 10'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d826 ||
	     WILL_FIRE_RL_m_rl_reset ;
  // register m_vrg_source_prio_1
  assign m_vrg_source_prio_1$D_IN =
	     MUX_m_vrg_source_prio_1$write_1__SEL_1 ?
	       wdata32__h27246[2:0] :
	       3'd0 ;
  assign m_vrg_source_prio_1$EN =
	     WILL_FIRE_RL_m_rl_process_wr_req &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d837 ||
	     WILL_FIRE_RL_m_rl_reset ;
  // register m_vrg_source_prio_10
  assign m_vrg_source_prio_10$D_IN =
	     MUX_m_vrg_source_prio_10$write_1__SEL_1 ?
	       wdata32__h27246[2:0] :
	       3'd0 ;
  assign m_vrg_source_prio_10$EN =
	     WILL_FIRE_RL_m_rl_process_wr_req &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d855 ||
	     WILL_FIRE_RL_m_rl_reset ;
  // register m_vrg_source_prio_11
  assign m_vrg_source_prio_11$D_IN =
	     MUX_m_vrg_source_prio_11$write_1__SEL_1 ?
	       wdata32__h27246[2:0] :
	       3'd0 ;
  assign m_vrg_source_prio_11$EN =
	     WILL_FIRE_RL_m_rl_process_wr_req &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d857 ||
	     WILL_FIRE_RL_m_rl_reset ;
  // register m_vrg_source_prio_12
  assign m_vrg_source_prio_12$D_IN =
	     MUX_m_vrg_source_prio_12$write_1__SEL_1 ?
	       wdata32__h27246[2:0] :
	       3'd0 ;
  assign m_vrg_source_prio_12$EN =
	     WILL_FIRE_RL_m_rl_process_wr_req &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d859 ||
	     WILL_FIRE_RL_m_rl_reset ;
  // register m_vrg_source_prio_13
  assign m_vrg_source_prio_13$D_IN =
	     MUX_m_vrg_source_prio_13$write_1__SEL_1 ?
	       wdata32__h27246[2:0] :
	       3'd0 ;
  assign m_vrg_source_prio_13$EN =
	     WILL_FIRE_RL_m_rl_process_wr_req &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d861 ||
	     WILL_FIRE_RL_m_rl_reset ;
  // register m_vrg_source_prio_14
  assign m_vrg_source_prio_14$D_IN =
	     MUX_m_vrg_source_prio_14$write_1__SEL_1 ?
	       wdata32__h27246[2:0] :
	       3'd0 ;
  assign m_vrg_source_prio_14$EN =
	     WILL_FIRE_RL_m_rl_process_wr_req &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d863 ||
	     WILL_FIRE_RL_m_rl_reset ;
  // register m_vrg_source_prio_15
  assign m_vrg_source_prio_15$D_IN =
	     MUX_m_vrg_source_prio_15$write_1__SEL_1 ?
	       wdata32__h27246[2:0] :
	       3'd0 ;
  assign m_vrg_source_prio_15$EN =
	     WILL_FIRE_RL_m_rl_process_wr_req &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d865 ||
	     WILL_FIRE_RL_m_rl_reset ;
  // register m_vrg_source_prio_16
  assign m_vrg_source_prio_16$D_IN =
	     MUX_m_vrg_source_prio_16$write_1__SEL_1 ?
	       wdata32__h27246[2:0] :
	       3'd0 ;
  assign m_vrg_source_prio_16$EN =
	     WILL_FIRE_RL_m_rl_process_wr_req &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d867 ||
	     WILL_FIRE_RL_m_rl_reset ;
  // register m_vrg_source_prio_2
  assign m_vrg_source_prio_2$D_IN =
	     MUX_m_vrg_source_prio_2$write_1__SEL_1 ?
	       wdata32__h27246[2:0] :
	       3'd0 ;
  assign m_vrg_source_prio_2$EN =
	     WILL_FIRE_RL_m_rl_process_wr_req &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d839 ||
	     WILL_FIRE_RL_m_rl_reset ;
  // register m_vrg_source_prio_3
  assign m_vrg_source_prio_3$D_IN =
	     MUX_m_vrg_source_prio_3$write_1__SEL_1 ?
	       wdata32__h27246[2:0] :
	       3'd0 ;
  assign m_vrg_source_prio_3$EN =
	     WILL_FIRE_RL_m_rl_process_wr_req &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d841 ||
	     WILL_FIRE_RL_m_rl_reset ;
  // register m_vrg_source_prio_4
  assign m_vrg_source_prio_4$D_IN =
	     MUX_m_vrg_source_prio_4$write_1__SEL_1 ?
	       wdata32__h27246[2:0] :
	       3'd0 ;
  assign m_vrg_source_prio_4$EN =
	     WILL_FIRE_RL_m_rl_process_wr_req &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d843 ||
	     WILL_FIRE_RL_m_rl_reset ;
  // register m_vrg_source_prio_5
  assign m_vrg_source_prio_5$D_IN =
	     MUX_m_vrg_source_prio_5$write_1__SEL_1 ?
	       wdata32__h27246[2:0] :
	       3'd0 ;
  assign m_vrg_source_prio_5$EN =
	     WILL_FIRE_RL_m_rl_process_wr_req &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d845 ||
	     WILL_FIRE_RL_m_rl_reset ;
  // register m_vrg_source_prio_6
  assign m_vrg_source_prio_6$D_IN =
	     MUX_m_vrg_source_prio_6$write_1__SEL_1 ?
	       wdata32__h27246[2:0] :
	       3'd0 ;
  assign m_vrg_source_prio_6$EN =
	     WILL_FIRE_RL_m_rl_process_wr_req &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d847 ||
	     WILL_FIRE_RL_m_rl_reset ;
  // register m_vrg_source_prio_7
  assign m_vrg_source_prio_7$D_IN =
	     MUX_m_vrg_source_prio_7$write_1__SEL_1 ?
	       wdata32__h27246[2:0] :
	       3'd0 ;
  assign m_vrg_source_prio_7$EN =
	     WILL_FIRE_RL_m_rl_process_wr_req &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d849 ||
	     WILL_FIRE_RL_m_rl_reset ;
  // register m_vrg_source_prio_8
  assign m_vrg_source_prio_8$D_IN =
	     MUX_m_vrg_source_prio_8$write_1__SEL_1 ?
	       wdata32__h27246[2:0] :
	       3'd0 ;
  assign m_vrg_source_prio_8$EN =
	     WILL_FIRE_RL_m_rl_process_wr_req &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d851 ||
	     WILL_FIRE_RL_m_rl_reset ;
  // register m_vrg_source_prio_9
  assign m_vrg_source_prio_9$D_IN =
	     MUX_m_vrg_source_prio_9$write_1__SEL_1 ?
	       wdata32__h27246[2:0] :
	       3'd0 ;
  assign m_vrg_source_prio_9$EN =
	     WILL_FIRE_RL_m_rl_process_wr_req &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d853 ||
	     WILL_FIRE_RL_m_rl_reset ;
  // register m_vrg_target_threshold_0
  assign m_vrg_target_threshold_0$D_IN =
	     MUX_m_vrg_target_threshold_0$write_1__SEL_1 ?
	       wdata32__h27246[2:0] :
	       3'd7 ;
  assign m_vrg_target_threshold_0$EN =
	     WILL_FIRE_RL_m_rl_process_wr_req &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d2860 ||
	     WILL_FIRE_RL_m_rl_reset ;
  // register m_vrg_target_threshold_1
  assign m_vrg_target_threshold_1$D_IN =
	     MUX_m_vrg_target_threshold_1$write_1__SEL_1 ?
	       wdata32__h27246[2:0] :
	       3'd7 ;
  assign m_vrg_target_threshold_1$EN =
	     WILL_FIRE_RL_m_rl_process_wr_req &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d2862 ||
	     WILL_FIRE_RL_m_rl_reset ;
  // register m_vvrg_ie_0_0
  assign m_vvrg_ie_0_0$D_IN =
	     MUX_m_vvrg_ie_0_0$write_1__SEL_1 &&
	     MUX_m_vvrg_ie_0_0$write_1__VAL_1 ;
  assign m_vvrg_ie_0_0$EN =
	     WILL_FIRE_RL_m_rl_process_wr_req && _dfoo2107 ||
	     WILL_FIRE_RL_m_rl_reset ;
  // register m_vvrg_ie_0_1
  assign m_vvrg_ie_0_1$D_IN =
	     MUX_m_vvrg_ie_0_1$write_1__SEL_1 &&
	     MUX_m_vvrg_ie_0_1$write_1__VAL_1 ;
  assign m_vvrg_ie_0_1$EN =
	     WILL_FIRE_RL_m_rl_process_wr_req && _dfoo2105 ||
	     WILL_FIRE_RL_m_rl_reset ;
  // register m_vvrg_ie_0_10
  assign m_vvrg_ie_0_10$D_IN =
	     MUX_m_vvrg_ie_0_10$write_1__SEL_1 &&
	     MUX_m_vvrg_ie_0_10$write_1__VAL_1 ;
  assign m_vvrg_ie_0_10$EN =
	     WILL_FIRE_RL_m_rl_process_wr_req && _dfoo2087 ||
	     WILL_FIRE_RL_m_rl_reset ;
  // register m_vvrg_ie_0_11
  assign m_vvrg_ie_0_11$D_IN =
	     MUX_m_vvrg_ie_0_11$write_1__SEL_1 &&
	     MUX_m_vvrg_ie_0_11$write_1__VAL_1 ;
  assign m_vvrg_ie_0_11$EN =
	     WILL_FIRE_RL_m_rl_process_wr_req && _dfoo2085 ||
	     WILL_FIRE_RL_m_rl_reset ;
  // register m_vvrg_ie_0_12
  assign m_vvrg_ie_0_12$D_IN =
	     MUX_m_vvrg_ie_0_12$write_1__SEL_1 &&
	     MUX_m_vvrg_ie_0_12$write_1__VAL_1 ;
  assign m_vvrg_ie_0_12$EN =
	     WILL_FIRE_RL_m_rl_process_wr_req && _dfoo2083 ||
	     WILL_FIRE_RL_m_rl_reset ;
  // register m_vvrg_ie_0_13
  assign m_vvrg_ie_0_13$D_IN =
	     MUX_m_vvrg_ie_0_13$write_1__SEL_1 &&
	     MUX_m_vvrg_ie_0_13$write_1__VAL_1 ;
  assign m_vvrg_ie_0_13$EN =
	     WILL_FIRE_RL_m_rl_process_wr_req && _dfoo2081 ||
	     WILL_FIRE_RL_m_rl_reset ;
  // register m_vvrg_ie_0_14
  assign m_vvrg_ie_0_14$D_IN =
	     MUX_m_vvrg_ie_0_14$write_1__SEL_1 &&
	     MUX_m_vvrg_ie_0_14$write_1__VAL_1 ;
  assign m_vvrg_ie_0_14$EN =
	     WILL_FIRE_RL_m_rl_process_wr_req && _dfoo2079 ||
	     WILL_FIRE_RL_m_rl_reset ;
  // register m_vvrg_ie_0_15
  assign m_vvrg_ie_0_15$D_IN =
	     MUX_m_vvrg_ie_0_15$write_1__SEL_1 &&
	     MUX_m_vvrg_ie_0_15$write_1__VAL_1 ;
  assign m_vvrg_ie_0_15$EN =
	     WILL_FIRE_RL_m_rl_process_wr_req && _dfoo2077 ||
	     WILL_FIRE_RL_m_rl_reset ;
  // register m_vvrg_ie_0_16
  assign m_vvrg_ie_0_16$D_IN =
	     MUX_m_vvrg_ie_0_16$write_1__SEL_1 &&
	     MUX_m_vvrg_ie_0_16$write_1__VAL_1 ;
  assign m_vvrg_ie_0_16$EN =
	     WILL_FIRE_RL_m_rl_process_wr_req && _dfoo2075 ||
	     WILL_FIRE_RL_m_rl_reset ;
  // register m_vvrg_ie_0_2
  assign m_vvrg_ie_0_2$D_IN =
	     MUX_m_vvrg_ie_0_2$write_1__SEL_1 &&
	     MUX_m_vvrg_ie_0_2$write_1__VAL_1 ;
  assign m_vvrg_ie_0_2$EN =
	     WILL_FIRE_RL_m_rl_process_wr_req && _dfoo2103 ||
	     WILL_FIRE_RL_m_rl_reset ;
  // register m_vvrg_ie_0_3
  assign m_vvrg_ie_0_3$D_IN =
	     MUX_m_vvrg_ie_0_3$write_1__SEL_1 &&
	     MUX_m_vvrg_ie_0_3$write_1__VAL_1 ;
  assign m_vvrg_ie_0_3$EN =
	     WILL_FIRE_RL_m_rl_process_wr_req && _dfoo2101 ||
	     WILL_FIRE_RL_m_rl_reset ;
  // register m_vvrg_ie_0_4
  assign m_vvrg_ie_0_4$D_IN =
	     MUX_m_vvrg_ie_0_4$write_1__SEL_1 &&
	     MUX_m_vvrg_ie_0_4$write_1__VAL_1 ;
  assign m_vvrg_ie_0_4$EN =
	     WILL_FIRE_RL_m_rl_process_wr_req && _dfoo2099 ||
	     WILL_FIRE_RL_m_rl_reset ;
  // register m_vvrg_ie_0_5
  assign m_vvrg_ie_0_5$D_IN =
	     MUX_m_vvrg_ie_0_5$write_1__SEL_1 &&
	     MUX_m_vvrg_ie_0_5$write_1__VAL_1 ;
  assign m_vvrg_ie_0_5$EN =
	     WILL_FIRE_RL_m_rl_process_wr_req && _dfoo2097 ||
	     WILL_FIRE_RL_m_rl_reset ;
  // register m_vvrg_ie_0_6
  assign m_vvrg_ie_0_6$D_IN =
	     MUX_m_vvrg_ie_0_6$write_1__SEL_1 &&
	     MUX_m_vvrg_ie_0_6$write_1__VAL_1 ;
  assign m_vvrg_ie_0_6$EN =
	     WILL_FIRE_RL_m_rl_process_wr_req && _dfoo2095 ||
	     WILL_FIRE_RL_m_rl_reset ;
  // register m_vvrg_ie_0_7
  assign m_vvrg_ie_0_7$D_IN =
	     MUX_m_vvrg_ie_0_7$write_1__SEL_1 &&
	     MUX_m_vvrg_ie_0_7$write_1__VAL_1 ;
  assign m_vvrg_ie_0_7$EN =
	     WILL_FIRE_RL_m_rl_process_wr_req && _dfoo2093 ||
	     WILL_FIRE_RL_m_rl_reset ;
  // register m_vvrg_ie_0_8
  assign m_vvrg_ie_0_8$D_IN =
	     MUX_m_vvrg_ie_0_8$write_1__SEL_1 &&
	     MUX_m_vvrg_ie_0_8$write_1__VAL_1 ;
  assign m_vvrg_ie_0_8$EN =
	     WILL_FIRE_RL_m_rl_process_wr_req && _dfoo2091 ||
	     WILL_FIRE_RL_m_rl_reset ;
  // register m_vvrg_ie_0_9
  assign m_vvrg_ie_0_9$D_IN =
	     MUX_m_vvrg_ie_0_9$write_1__SEL_1 &&
	     MUX_m_vvrg_ie_0_9$write_1__VAL_1 ;
  assign m_vvrg_ie_0_9$EN =
	     WILL_FIRE_RL_m_rl_process_wr_req && _dfoo2089 ||
	     WILL_FIRE_RL_m_rl_reset ;
  // register m_vvrg_ie_1_0
  assign m_vvrg_ie_1_0$D_IN =
	     MUX_m_vvrg_ie_1_0$write_1__SEL_1 &&
	     MUX_m_vvrg_ie_1_0$write_1__VAL_1 ;
  assign m_vvrg_ie_1_0$EN =
	     WILL_FIRE_RL_m_rl_process_wr_req && _dfoo2073 ||
	     WILL_FIRE_RL_m_rl_reset ;
  // register m_vvrg_ie_1_1
  assign m_vvrg_ie_1_1$D_IN =
	     MUX_m_vvrg_ie_1_1$write_1__SEL_1 &&
	     MUX_m_vvrg_ie_1_1$write_1__VAL_1 ;
  assign m_vvrg_ie_1_1$EN =
	     WILL_FIRE_RL_m_rl_process_wr_req && _dfoo2071 ||
	     WILL_FIRE_RL_m_rl_reset ;
  // register m_vvrg_ie_1_10
  assign m_vvrg_ie_1_10$D_IN =
	     MUX_m_vvrg_ie_1_10$write_1__SEL_1 &&
	     MUX_m_vvrg_ie_1_10$write_1__VAL_1 ;
  assign m_vvrg_ie_1_10$EN =
	     WILL_FIRE_RL_m_rl_process_wr_req && _dfoo2053 ||
	     WILL_FIRE_RL_m_rl_reset ;
  // register m_vvrg_ie_1_11
  assign m_vvrg_ie_1_11$D_IN =
	     MUX_m_vvrg_ie_1_11$write_1__SEL_1 &&
	     MUX_m_vvrg_ie_1_11$write_1__VAL_1 ;
  assign m_vvrg_ie_1_11$EN =
	     WILL_FIRE_RL_m_rl_process_wr_req && _dfoo2051 ||
	     WILL_FIRE_RL_m_rl_reset ;
  // register m_vvrg_ie_1_12
  assign m_vvrg_ie_1_12$D_IN =
	     MUX_m_vvrg_ie_1_12$write_1__SEL_1 &&
	     MUX_m_vvrg_ie_1_12$write_1__VAL_1 ;
  assign m_vvrg_ie_1_12$EN =
	     WILL_FIRE_RL_m_rl_process_wr_req && _dfoo2049 ||
	     WILL_FIRE_RL_m_rl_reset ;
  // register m_vvrg_ie_1_13
  assign m_vvrg_ie_1_13$D_IN =
	     MUX_m_vvrg_ie_1_13$write_1__SEL_1 &&
	     MUX_m_vvrg_ie_1_13$write_1__VAL_1 ;
  assign m_vvrg_ie_1_13$EN =
	     WILL_FIRE_RL_m_rl_process_wr_req && _dfoo2047 ||
	     WILL_FIRE_RL_m_rl_reset ;
  // register m_vvrg_ie_1_14
  assign m_vvrg_ie_1_14$D_IN =
	     MUX_m_vvrg_ie_1_14$write_1__SEL_1 &&
	     MUX_m_vvrg_ie_1_14$write_1__VAL_1 ;
  assign m_vvrg_ie_1_14$EN =
	     WILL_FIRE_RL_m_rl_process_wr_req && _dfoo2045 ||
	     WILL_FIRE_RL_m_rl_reset ;
  // register m_vvrg_ie_1_15
  assign m_vvrg_ie_1_15$D_IN =
	     MUX_m_vvrg_ie_1_15$write_1__SEL_1 &&
	     MUX_m_vvrg_ie_1_15$write_1__VAL_1 ;
  assign m_vvrg_ie_1_15$EN =
	     WILL_FIRE_RL_m_rl_process_wr_req && _dfoo2043 ||
	     WILL_FIRE_RL_m_rl_reset ;
  // register m_vvrg_ie_1_16
  assign m_vvrg_ie_1_16$D_IN =
	     MUX_m_vvrg_ie_1_16$write_1__SEL_1 &&
	     MUX_m_vvrg_ie_1_16$write_1__VAL_1 ;
  assign m_vvrg_ie_1_16$EN =
	     WILL_FIRE_RL_m_rl_process_wr_req && _dfoo2041 ||
	     WILL_FIRE_RL_m_rl_reset ;
  // register m_vvrg_ie_1_2
  assign m_vvrg_ie_1_2$D_IN =
	     MUX_m_vvrg_ie_1_2$write_1__SEL_1 &&
	     MUX_m_vvrg_ie_1_2$write_1__VAL_1 ;
  assign m_vvrg_ie_1_2$EN =
	     WILL_FIRE_RL_m_rl_process_wr_req && _dfoo2069 ||
	     WILL_FIRE_RL_m_rl_reset ;
  // register m_vvrg_ie_1_3
  assign m_vvrg_ie_1_3$D_IN =
	     MUX_m_vvrg_ie_1_3$write_1__SEL_1 &&
	     MUX_m_vvrg_ie_1_3$write_1__VAL_1 ;
  assign m_vvrg_ie_1_3$EN =
	     WILL_FIRE_RL_m_rl_process_wr_req && _dfoo2067 ||
	     WILL_FIRE_RL_m_rl_reset ;
  // register m_vvrg_ie_1_4
  assign m_vvrg_ie_1_4$D_IN =
	     MUX_m_vvrg_ie_1_4$write_1__SEL_1 &&
	     MUX_m_vvrg_ie_1_4$write_1__VAL_1 ;
  assign m_vvrg_ie_1_4$EN =
	     WILL_FIRE_RL_m_rl_process_wr_req && _dfoo2065 ||
	     WILL_FIRE_RL_m_rl_reset ;
  // register m_vvrg_ie_1_5
  assign m_vvrg_ie_1_5$D_IN =
	     MUX_m_vvrg_ie_1_5$write_1__SEL_1 &&
	     MUX_m_vvrg_ie_1_5$write_1__VAL_1 ;
  assign m_vvrg_ie_1_5$EN =
	     WILL_FIRE_RL_m_rl_process_wr_req && _dfoo2063 ||
	     WILL_FIRE_RL_m_rl_reset ;
  // register m_vvrg_ie_1_6
  assign m_vvrg_ie_1_6$D_IN =
	     MUX_m_vvrg_ie_1_6$write_1__SEL_1 &&
	     MUX_m_vvrg_ie_1_6$write_1__VAL_1 ;
  assign m_vvrg_ie_1_6$EN =
	     WILL_FIRE_RL_m_rl_process_wr_req && _dfoo2061 ||
	     WILL_FIRE_RL_m_rl_reset ;
  // register m_vvrg_ie_1_7
  assign m_vvrg_ie_1_7$D_IN =
	     MUX_m_vvrg_ie_1_7$write_1__SEL_1 &&
	     MUX_m_vvrg_ie_1_7$write_1__VAL_1 ;
  assign m_vvrg_ie_1_7$EN =
	     WILL_FIRE_RL_m_rl_process_wr_req && _dfoo2059 ||
	     WILL_FIRE_RL_m_rl_reset ;
  // register m_vvrg_ie_1_8
  assign m_vvrg_ie_1_8$D_IN =
	     MUX_m_vvrg_ie_1_8$write_1__SEL_1 &&
	     MUX_m_vvrg_ie_1_8$write_1__VAL_1 ;
  assign m_vvrg_ie_1_8$EN =
	     WILL_FIRE_RL_m_rl_process_wr_req && _dfoo2057 ||
	     WILL_FIRE_RL_m_rl_reset ;
  // register m_vvrg_ie_1_9
  assign m_vvrg_ie_1_9$D_IN =
	     MUX_m_vvrg_ie_1_9$write_1__SEL_1 &&
	     MUX_m_vvrg_ie_1_9$write_1__VAL_1 ;
  assign m_vvrg_ie_1_9$EN =
	     WILL_FIRE_RL_m_rl_process_wr_req && _dfoo2055 ||
	     WILL_FIRE_RL_m_rl_reset ;
  // submodule m_f_reset_reqs
  assign m_f_reset_reqs$ENQ = EN_server_reset_request_put ;
  assign m_f_reset_reqs$DEQ = CAN_FIRE_RL_m_rl_reset ;
  assign m_f_reset_reqs$CLR = 1'b0 ;
  // submodule m_f_reset_rsps
  assign m_f_reset_rsps$ENQ = CAN_FIRE_RL_m_rl_reset ;
  assign m_f_reset_rsps$DEQ = EN_server_reset_response_get ;
  assign m_f_reset_rsps$CLR = 1'b0 ;
  // submodule m_slave_xactor_f_rd_addr
  assign m_slave_xactor_f_rd_addr$D_IN =
	     { axi4_slave_arid,
	       axi4_slave_araddr,
	       axi4_slave_arlen,
	       axi4_slave_arsize,
	       axi4_slave_arburst,
	       axi4_slave_arlock,
	       axi4_slave_arcache,
	       axi4_slave_arprot,
	       axi4_slave_arqos,
	       axi4_slave_arregion } ;
  assign m_slave_xactor_f_rd_addr$ENQ =
	     axi4_slave_arvalid && m_slave_xactor_f_rd_addr$FULL_N ;
  assign m_slave_xactor_f_rd_addr$DEQ = CAN_FIRE_RL_m_rl_process_rd_req ;
  assign m_slave_xactor_f_rd_addr$CLR = CAN_FIRE_RL_m_rl_reset ;
  // submodule m_slave_xactor_f_rd_data
  assign m_slave_xactor_f_rd_data$D_IN =
	     { m_slave_xactor_f_rd_addr$D_OUT[96:93],
	       x__h26677,
	       rresp__h26521,
	       1'd1 } ;
  assign m_slave_xactor_f_rd_data$ENQ = CAN_FIRE_RL_m_rl_process_rd_req ;
  assign m_slave_xactor_f_rd_data$DEQ =
	     axi4_slave_rready && m_slave_xactor_f_rd_data$EMPTY_N ;
  assign m_slave_xactor_f_rd_data$CLR = CAN_FIRE_RL_m_rl_reset ;
  // submodule m_slave_xactor_f_wr_addr
  assign m_slave_xactor_f_wr_addr$D_IN =
	     { axi4_slave_awid,
	       axi4_slave_awaddr,
	       axi4_slave_awlen,
	       axi4_slave_awsize,
	       axi4_slave_awburst,
	       axi4_slave_awlock,
	       axi4_slave_awcache,
	       axi4_slave_awprot,
	       axi4_slave_awqos,
	       axi4_slave_awregion } ;
  assign m_slave_xactor_f_wr_addr$ENQ =
	     axi4_slave_awvalid && m_slave_xactor_f_wr_addr$FULL_N ;
  assign m_slave_xactor_f_wr_addr$DEQ = CAN_FIRE_RL_m_rl_process_wr_req ;
  assign m_slave_xactor_f_wr_addr$CLR = CAN_FIRE_RL_m_rl_reset ;
  // submodule m_slave_xactor_f_wr_data
  assign m_slave_xactor_f_wr_data$D_IN =
	     { axi4_slave_wdata, axi4_slave_wstrb, axi4_slave_wlast } ;
  assign m_slave_xactor_f_wr_data$ENQ =
	     axi4_slave_wvalid && m_slave_xactor_f_wr_data$FULL_N ;
  assign m_slave_xactor_f_wr_data$DEQ = CAN_FIRE_RL_m_rl_process_wr_req ;
  assign m_slave_xactor_f_wr_data$CLR = CAN_FIRE_RL_m_rl_reset ;
  // submodule m_slave_xactor_f_wr_resp
  assign m_slave_xactor_f_wr_resp$D_IN =
	     { m_slave_xactor_f_wr_addr$D_OUT[96:93], v__h27250 } ;
  assign m_slave_xactor_f_wr_resp$ENQ = CAN_FIRE_RL_m_rl_process_wr_req ;
  assign m_slave_xactor_f_wr_resp$DEQ =
	     axi4_slave_bready && m_slave_xactor_f_wr_resp$EMPTY_N ;
  assign m_slave_xactor_f_wr_resp$CLR = CAN_FIRE_RL_m_rl_reset ;
  // remaining internal signals
  assign IF_m_slave_xactor_f_rd_addr_first__9_BITS_92_T_ETC___d748 =
	     m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d240 ?
	       !m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d71 ||
	       !m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d242 :
	       x__h23928 != 32'h00200000 && x__h23928 != 32'h00200004 ||
	       !m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d532 ;
  assign IF_m_slave_xactor_f_rd_addr_first__9_BITS_92_T_ETC___d750 =
	     m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d36 ?
	       addr_offset__h13465[11:2] == 10'd0 ||
	       !m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d40 :
	       (m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d68 ?
		  !m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d71 :
		  IF_m_slave_xactor_f_rd_addr_first__9_BITS_92_T_ETC___d748) ;
  assign IF_m_slave_xactor_f_wr_addr_first__94_BITS_92__ETC___d2874 =
	     wdata32__h27246[9:0] <= 10'd17 ;
  assign IF_m_slave_xactor_f_wr_addr_first__94_BITS_92__ETC___d2950 =
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d888 ?
	       !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d877 ||
	       !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d889 :
	       x__h76716 != 32'h00200000 && x__h76716 != 32'h00200004 ||
	       !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d2854 ;
  assign IF_m_slave_xactor_f_wr_addr_first__94_BITS_92__ETC___d2952 =
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d821 ?
	       addr_offset__h27245[11:2] == 10'd0 ||
	       !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d823 :
	       (m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d874 ?
		  !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d877 :
		  IF_m_slave_xactor_f_wr_addr_first__94_BITS_92__ETC___d2950) ;
  assign IF_m_vrg_source_ip_10_read__0_AND_NOT_m_vrg_so_ETC___d3037 =
	     m_vrg_source_ip_10_read__0_AND_NOT_m_vrg_sourc_ETC___d3036 ?
	       m_vrg_source_prio_10 :
	       IF_m_vrg_source_ip_9_read__9_AND_NOT_m_vrg_sou_ETC___d3032 ;
  assign IF_m_vrg_source_ip_10_read__0_AND_NOT_m_vrg_so_ETC___d3131 =
	     m_vrg_source_ip_10_read__0_AND_NOT_m_vrg_sourc_ETC___d3130 ?
	       m_vrg_source_prio_10 :
	       IF_m_vrg_source_ip_9_read__9_AND_NOT_m_vrg_sou_ETC___d3126 ;
  assign IF_m_vrg_source_ip_10_read__0_AND_NOT_m_vrg_so_ETC___d615 =
	     m_vrg_source_ip_10_read__0_AND_NOT_m_vrg_sourc_ETC___d614 ?
	       m_vrg_source_prio_10 :
	       IF_m_vrg_source_ip_9_read__9_AND_NOT_m_vrg_sou_ETC___d608 ;
  assign IF_m_vrg_source_ip_11_read__1_AND_NOT_m_vrg_so_ETC___d3042 =
	     m_vrg_source_ip_11_read__1_AND_NOT_m_vrg_sourc_ETC___d3041 ?
	       m_vrg_source_prio_11 :
	       IF_m_vrg_source_ip_10_read__0_AND_NOT_m_vrg_so_ETC___d3037 ;
  assign IF_m_vrg_source_ip_11_read__1_AND_NOT_m_vrg_so_ETC___d3078 =
	     m_vrg_source_ip_11_read__1_AND_NOT_m_vrg_sourc_ETC___d3041 ?
	       5'd11 :
	       (m_vrg_source_ip_10_read__0_AND_NOT_m_vrg_sourc_ETC___d3036 ?
		  5'd10 :
		  IF_m_vrg_source_ip_9_read__9_AND_NOT_m_vrg_sou_ETC___d3076) ;
  assign IF_m_vrg_source_ip_11_read__1_AND_NOT_m_vrg_so_ETC___d3136 =
	     m_vrg_source_ip_11_read__1_AND_NOT_m_vrg_sourc_ETC___d3135 ?
	       m_vrg_source_prio_11 :
	       IF_m_vrg_source_ip_10_read__0_AND_NOT_m_vrg_so_ETC___d3131 ;
  assign IF_m_vrg_source_ip_11_read__1_AND_NOT_m_vrg_so_ETC___d3172 =
	     m_vrg_source_ip_11_read__1_AND_NOT_m_vrg_sourc_ETC___d3135 ?
	       5'd11 :
	       (m_vrg_source_ip_10_read__0_AND_NOT_m_vrg_sourc_ETC___d3130 ?
		  5'd10 :
		  IF_m_vrg_source_ip_9_read__9_AND_NOT_m_vrg_sou_ETC___d3170) ;
  assign IF_m_vrg_source_ip_11_read__1_AND_NOT_m_vrg_so_ETC___d622 =
	     m_vrg_source_ip_11_read__1_AND_NOT_m_vrg_sourc_ETC___d621 ?
	       m_vrg_source_prio_11 :
	       IF_m_vrg_source_ip_10_read__0_AND_NOT_m_vrg_so_ETC___d615 ;
  assign IF_m_vrg_source_ip_11_read__1_AND_NOT_m_vrg_so_ETC___d667 =
	     m_vrg_source_ip_11_read__1_AND_NOT_m_vrg_sourc_ETC___d621 ?
	       5'd11 :
	       (m_vrg_source_ip_10_read__0_AND_NOT_m_vrg_sourc_ETC___d614 ?
		  5'd10 :
		  IF_m_vrg_source_ip_9_read__9_AND_NOT_m_vrg_sou_ETC___d665) ;
  assign IF_m_vrg_source_ip_12_read__2_AND_NOT_m_vrg_so_ETC___d3047 =
	     m_vrg_source_ip_12_read__2_AND_NOT_m_vrg_sourc_ETC___d3046 ?
	       m_vrg_source_prio_12 :
	       IF_m_vrg_source_ip_11_read__1_AND_NOT_m_vrg_so_ETC___d3042 ;
  assign IF_m_vrg_source_ip_12_read__2_AND_NOT_m_vrg_so_ETC___d3141 =
	     m_vrg_source_ip_12_read__2_AND_NOT_m_vrg_sourc_ETC___d3140 ?
	       m_vrg_source_prio_12 :
	       IF_m_vrg_source_ip_11_read__1_AND_NOT_m_vrg_so_ETC___d3136 ;
  assign IF_m_vrg_source_ip_12_read__2_AND_NOT_m_vrg_so_ETC___d629 =
	     m_vrg_source_ip_12_read__2_AND_NOT_m_vrg_sourc_ETC___d628 ?
	       m_vrg_source_prio_12 :
	       IF_m_vrg_source_ip_11_read__1_AND_NOT_m_vrg_so_ETC___d622 ;
  assign IF_m_vrg_source_ip_13_read__3_AND_NOT_m_vrg_so_ETC___d3052 =
	     m_vrg_source_ip_13_read__3_AND_NOT_m_vrg_sourc_ETC___d3051 ?
	       m_vrg_source_prio_13 :
	       IF_m_vrg_source_ip_12_read__2_AND_NOT_m_vrg_so_ETC___d3047 ;
  assign IF_m_vrg_source_ip_13_read__3_AND_NOT_m_vrg_so_ETC___d3080 =
	     m_vrg_source_ip_13_read__3_AND_NOT_m_vrg_sourc_ETC___d3051 ?
	       5'd13 :
	       (m_vrg_source_ip_12_read__2_AND_NOT_m_vrg_sourc_ETC___d3046 ?
		  5'd12 :
		  IF_m_vrg_source_ip_11_read__1_AND_NOT_m_vrg_so_ETC___d3078) ;
  assign IF_m_vrg_source_ip_13_read__3_AND_NOT_m_vrg_so_ETC___d3146 =
	     m_vrg_source_ip_13_read__3_AND_NOT_m_vrg_sourc_ETC___d3145 ?
	       m_vrg_source_prio_13 :
	       IF_m_vrg_source_ip_12_read__2_AND_NOT_m_vrg_so_ETC___d3141 ;
  assign IF_m_vrg_source_ip_13_read__3_AND_NOT_m_vrg_so_ETC___d3174 =
	     m_vrg_source_ip_13_read__3_AND_NOT_m_vrg_sourc_ETC___d3145 ?
	       5'd13 :
	       (m_vrg_source_ip_12_read__2_AND_NOT_m_vrg_sourc_ETC___d3140 ?
		  5'd12 :
		  IF_m_vrg_source_ip_11_read__1_AND_NOT_m_vrg_so_ETC___d3172) ;
  assign IF_m_vrg_source_ip_13_read__3_AND_NOT_m_vrg_so_ETC___d636 =
	     m_vrg_source_ip_13_read__3_AND_NOT_m_vrg_sourc_ETC___d635 ?
	       m_vrg_source_prio_13 :
	       IF_m_vrg_source_ip_12_read__2_AND_NOT_m_vrg_so_ETC___d629 ;
  assign IF_m_vrg_source_ip_13_read__3_AND_NOT_m_vrg_so_ETC___d669 =
	     m_vrg_source_ip_13_read__3_AND_NOT_m_vrg_sourc_ETC___d635 ?
	       5'd13 :
	       (m_vrg_source_ip_12_read__2_AND_NOT_m_vrg_sourc_ETC___d628 ?
		  5'd12 :
		  IF_m_vrg_source_ip_11_read__1_AND_NOT_m_vrg_so_ETC___d667) ;
  assign IF_m_vrg_source_ip_14_read__4_AND_NOT_m_vrg_so_ETC___d3057 =
	     m_vrg_source_ip_14_read__4_AND_NOT_m_vrg_sourc_ETC___d3056 ?
	       m_vrg_source_prio_14 :
	       IF_m_vrg_source_ip_13_read__3_AND_NOT_m_vrg_so_ETC___d3052 ;
  assign IF_m_vrg_source_ip_14_read__4_AND_NOT_m_vrg_so_ETC___d3151 =
	     m_vrg_source_ip_14_read__4_AND_NOT_m_vrg_sourc_ETC___d3150 ?
	       m_vrg_source_prio_14 :
	       IF_m_vrg_source_ip_13_read__3_AND_NOT_m_vrg_so_ETC___d3146 ;
  assign IF_m_vrg_source_ip_14_read__4_AND_NOT_m_vrg_so_ETC___d643 =
	     m_vrg_source_ip_14_read__4_AND_NOT_m_vrg_sourc_ETC___d642 ?
	       m_vrg_source_prio_14 :
	       IF_m_vrg_source_ip_13_read__3_AND_NOT_m_vrg_so_ETC___d636 ;
  assign IF_m_vrg_source_ip_15_read__5_AND_NOT_m_vrg_so_ETC___d3062 =
	     m_vrg_source_ip_15_read__5_AND_NOT_m_vrg_sourc_ETC___d3061 ?
	       m_vrg_source_prio_15 :
	       IF_m_vrg_source_ip_14_read__4_AND_NOT_m_vrg_so_ETC___d3057 ;
  assign IF_m_vrg_source_ip_15_read__5_AND_NOT_m_vrg_so_ETC___d3082 =
	     m_vrg_source_ip_15_read__5_AND_NOT_m_vrg_sourc_ETC___d3061 ?
	       5'd15 :
	       (m_vrg_source_ip_14_read__4_AND_NOT_m_vrg_sourc_ETC___d3056 ?
		  5'd14 :
		  IF_m_vrg_source_ip_13_read__3_AND_NOT_m_vrg_so_ETC___d3080) ;
  assign IF_m_vrg_source_ip_15_read__5_AND_NOT_m_vrg_so_ETC___d3156 =
	     m_vrg_source_ip_15_read__5_AND_NOT_m_vrg_sourc_ETC___d3155 ?
	       m_vrg_source_prio_15 :
	       IF_m_vrg_source_ip_14_read__4_AND_NOT_m_vrg_so_ETC___d3151 ;
  assign IF_m_vrg_source_ip_15_read__5_AND_NOT_m_vrg_so_ETC___d3176 =
	     m_vrg_source_ip_15_read__5_AND_NOT_m_vrg_sourc_ETC___d3155 ?
	       5'd15 :
	       (m_vrg_source_ip_14_read__4_AND_NOT_m_vrg_sourc_ETC___d3150 ?
		  5'd14 :
		  IF_m_vrg_source_ip_13_read__3_AND_NOT_m_vrg_so_ETC___d3174) ;
  assign IF_m_vrg_source_ip_15_read__5_AND_NOT_m_vrg_so_ETC___d671 =
	     m_vrg_source_ip_15_read__5_AND_NOT_m_vrg_sourc_ETC___d649 ?
	       5'd15 :
	       (m_vrg_source_ip_14_read__4_AND_NOT_m_vrg_sourc_ETC___d642 ?
		  5'd14 :
		  IF_m_vrg_source_ip_13_read__3_AND_NOT_m_vrg_so_ETC___d669) ;
  assign IF_m_vrg_source_ip_1_read__1_AND_NOT_m_vrg_sou_ETC___d2992 =
	     (m_vrg_source_ip_1 && m_vrg_source_prio_1 != 3'd0 &&
	      m_vvrg_ie_0_1) ?
	       m_vrg_source_prio_1 :
	       3'd0 ;
  assign IF_m_vrg_source_ip_1_read__1_AND_NOT_m_vrg_sou_ETC___d3086 =
	     (m_vrg_source_ip_1 && m_vrg_source_prio_1 != 3'd0 &&
	      m_vvrg_ie_1_1) ?
	       m_vrg_source_prio_1 :
	       3'd0 ;
  assign IF_m_vrg_source_ip_1_read__1_AND_NOT_m_vrg_sou_ETC___d552 =
	     m_vrg_source_ip_1_read__1_AND_NOT_m_vrg_source_ETC___d551 ?
	       m_vrg_source_prio_1 :
	       3'd0 ;
  assign IF_m_vrg_source_ip_2_read__2_AND_NOT_m_vrg_sou_ETC___d2997 =
	     m_vrg_source_ip_2_read__2_AND_NOT_m_vrg_source_ETC___d2996 ?
	       m_vrg_source_prio_2 :
	       IF_m_vrg_source_ip_1_read__1_AND_NOT_m_vrg_sou_ETC___d2992 ;
  assign IF_m_vrg_source_ip_2_read__2_AND_NOT_m_vrg_sou_ETC___d3091 =
	     m_vrg_source_ip_2_read__2_AND_NOT_m_vrg_source_ETC___d3090 ?
	       m_vrg_source_prio_2 :
	       IF_m_vrg_source_ip_1_read__1_AND_NOT_m_vrg_sou_ETC___d3086 ;
  assign IF_m_vrg_source_ip_2_read__2_AND_NOT_m_vrg_sou_ETC___d559 =
	     m_vrg_source_ip_2_read__2_AND_NOT_m_vrg_source_ETC___d558 ?
	       m_vrg_source_prio_2 :
	       IF_m_vrg_source_ip_1_read__1_AND_NOT_m_vrg_sou_ETC___d552 ;
  assign IF_m_vrg_source_ip_3_read__3_AND_NOT_m_vrg_sou_ETC___d3002 =
	     m_vrg_source_ip_3_read__3_AND_NOT_m_vrg_source_ETC___d3001 ?
	       m_vrg_source_prio_3 :
	       IF_m_vrg_source_ip_2_read__2_AND_NOT_m_vrg_sou_ETC___d2997 ;
  assign IF_m_vrg_source_ip_3_read__3_AND_NOT_m_vrg_sou_ETC___d3070 =
	     m_vrg_source_ip_3_read__3_AND_NOT_m_vrg_source_ETC___d3001 ?
	       5'd3 :
	       (m_vrg_source_ip_2_read__2_AND_NOT_m_vrg_source_ETC___d2996 ?
		  5'd2 :
		  ((m_vrg_source_ip_1 && m_vrg_source_prio_1 != 3'd0 &&
		    m_vvrg_ie_0_1) ?
		     5'd1 :
		     5'd0)) ;
  assign IF_m_vrg_source_ip_3_read__3_AND_NOT_m_vrg_sou_ETC___d3096 =
	     m_vrg_source_ip_3_read__3_AND_NOT_m_vrg_source_ETC___d3095 ?
	       m_vrg_source_prio_3 :
	       IF_m_vrg_source_ip_2_read__2_AND_NOT_m_vrg_sou_ETC___d3091 ;
  assign IF_m_vrg_source_ip_3_read__3_AND_NOT_m_vrg_sou_ETC___d3164 =
	     m_vrg_source_ip_3_read__3_AND_NOT_m_vrg_source_ETC___d3095 ?
	       5'd3 :
	       (m_vrg_source_ip_2_read__2_AND_NOT_m_vrg_source_ETC___d3090 ?
		  5'd2 :
		  ((m_vrg_source_ip_1 && m_vrg_source_prio_1 != 3'd0 &&
		    m_vvrg_ie_1_1) ?
		     5'd1 :
		     5'd0)) ;
  assign IF_m_vrg_source_ip_3_read__3_AND_NOT_m_vrg_sou_ETC___d566 =
	     m_vrg_source_ip_3_read__3_AND_NOT_m_vrg_source_ETC___d565 ?
	       m_vrg_source_prio_3 :
	       IF_m_vrg_source_ip_2_read__2_AND_NOT_m_vrg_sou_ETC___d559 ;
  assign IF_m_vrg_source_ip_3_read__3_AND_NOT_m_vrg_sou_ETC___d659 =
	     m_vrg_source_ip_3_read__3_AND_NOT_m_vrg_source_ETC___d565 ?
	       5'd3 :
	       (m_vrg_source_ip_2_read__2_AND_NOT_m_vrg_source_ETC___d558 ?
		  5'd2 :
		  (m_vrg_source_ip_1_read__1_AND_NOT_m_vrg_source_ETC___d551 ?
		     5'd1 :
		     5'd0)) ;
  assign IF_m_vrg_source_ip_4_read__4_AND_NOT_m_vrg_sou_ETC___d3007 =
	     m_vrg_source_ip_4_read__4_AND_NOT_m_vrg_source_ETC___d3006 ?
	       m_vrg_source_prio_4 :
	       IF_m_vrg_source_ip_3_read__3_AND_NOT_m_vrg_sou_ETC___d3002 ;
  assign IF_m_vrg_source_ip_4_read__4_AND_NOT_m_vrg_sou_ETC___d3101 =
	     m_vrg_source_ip_4_read__4_AND_NOT_m_vrg_source_ETC___d3100 ?
	       m_vrg_source_prio_4 :
	       IF_m_vrg_source_ip_3_read__3_AND_NOT_m_vrg_sou_ETC___d3096 ;
  assign IF_m_vrg_source_ip_4_read__4_AND_NOT_m_vrg_sou_ETC___d573 =
	     m_vrg_source_ip_4_read__4_AND_NOT_m_vrg_source_ETC___d572 ?
	       m_vrg_source_prio_4 :
	       IF_m_vrg_source_ip_3_read__3_AND_NOT_m_vrg_sou_ETC___d566 ;
  assign IF_m_vrg_source_ip_5_read__5_AND_NOT_m_vrg_sou_ETC___d3012 =
	     m_vrg_source_ip_5_read__5_AND_NOT_m_vrg_source_ETC___d3011 ?
	       m_vrg_source_prio_5 :
	       IF_m_vrg_source_ip_4_read__4_AND_NOT_m_vrg_sou_ETC___d3007 ;
  assign IF_m_vrg_source_ip_5_read__5_AND_NOT_m_vrg_sou_ETC___d3072 =
	     m_vrg_source_ip_5_read__5_AND_NOT_m_vrg_source_ETC___d3011 ?
	       5'd5 :
	       (m_vrg_source_ip_4_read__4_AND_NOT_m_vrg_source_ETC___d3006 ?
		  5'd4 :
		  IF_m_vrg_source_ip_3_read__3_AND_NOT_m_vrg_sou_ETC___d3070) ;
  assign IF_m_vrg_source_ip_5_read__5_AND_NOT_m_vrg_sou_ETC___d3106 =
	     m_vrg_source_ip_5_read__5_AND_NOT_m_vrg_source_ETC___d3105 ?
	       m_vrg_source_prio_5 :
	       IF_m_vrg_source_ip_4_read__4_AND_NOT_m_vrg_sou_ETC___d3101 ;
  assign IF_m_vrg_source_ip_5_read__5_AND_NOT_m_vrg_sou_ETC___d3166 =
	     m_vrg_source_ip_5_read__5_AND_NOT_m_vrg_source_ETC___d3105 ?
	       5'd5 :
	       (m_vrg_source_ip_4_read__4_AND_NOT_m_vrg_source_ETC___d3100 ?
		  5'd4 :
		  IF_m_vrg_source_ip_3_read__3_AND_NOT_m_vrg_sou_ETC___d3164) ;
  assign IF_m_vrg_source_ip_5_read__5_AND_NOT_m_vrg_sou_ETC___d580 =
	     m_vrg_source_ip_5_read__5_AND_NOT_m_vrg_source_ETC___d579 ?
	       m_vrg_source_prio_5 :
	       IF_m_vrg_source_ip_4_read__4_AND_NOT_m_vrg_sou_ETC___d573 ;
  assign IF_m_vrg_source_ip_5_read__5_AND_NOT_m_vrg_sou_ETC___d661 =
	     m_vrg_source_ip_5_read__5_AND_NOT_m_vrg_source_ETC___d579 ?
	       5'd5 :
	       (m_vrg_source_ip_4_read__4_AND_NOT_m_vrg_source_ETC___d572 ?
		  5'd4 :
		  IF_m_vrg_source_ip_3_read__3_AND_NOT_m_vrg_sou_ETC___d659) ;
  assign IF_m_vrg_source_ip_6_read__6_AND_NOT_m_vrg_sou_ETC___d3017 =
	     m_vrg_source_ip_6_read__6_AND_NOT_m_vrg_source_ETC___d3016 ?
	       m_vrg_source_prio_6 :
	       IF_m_vrg_source_ip_5_read__5_AND_NOT_m_vrg_sou_ETC___d3012 ;
  assign IF_m_vrg_source_ip_6_read__6_AND_NOT_m_vrg_sou_ETC___d3111 =
	     m_vrg_source_ip_6_read__6_AND_NOT_m_vrg_source_ETC___d3110 ?
	       m_vrg_source_prio_6 :
	       IF_m_vrg_source_ip_5_read__5_AND_NOT_m_vrg_sou_ETC___d3106 ;
  assign IF_m_vrg_source_ip_6_read__6_AND_NOT_m_vrg_sou_ETC___d587 =
	     m_vrg_source_ip_6_read__6_AND_NOT_m_vrg_source_ETC___d586 ?
	       m_vrg_source_prio_6 :
	       IF_m_vrg_source_ip_5_read__5_AND_NOT_m_vrg_sou_ETC___d580 ;
  assign IF_m_vrg_source_ip_7_read__7_AND_NOT_m_vrg_sou_ETC___d3022 =
	     m_vrg_source_ip_7_read__7_AND_NOT_m_vrg_source_ETC___d3021 ?
	       m_vrg_source_prio_7 :
	       IF_m_vrg_source_ip_6_read__6_AND_NOT_m_vrg_sou_ETC___d3017 ;
  assign IF_m_vrg_source_ip_7_read__7_AND_NOT_m_vrg_sou_ETC___d3074 =
	     m_vrg_source_ip_7_read__7_AND_NOT_m_vrg_source_ETC___d3021 ?
	       5'd7 :
	       (m_vrg_source_ip_6_read__6_AND_NOT_m_vrg_source_ETC___d3016 ?
		  5'd6 :
		  IF_m_vrg_source_ip_5_read__5_AND_NOT_m_vrg_sou_ETC___d3072) ;
  assign IF_m_vrg_source_ip_7_read__7_AND_NOT_m_vrg_sou_ETC___d3116 =
	     m_vrg_source_ip_7_read__7_AND_NOT_m_vrg_source_ETC___d3115 ?
	       m_vrg_source_prio_7 :
	       IF_m_vrg_source_ip_6_read__6_AND_NOT_m_vrg_sou_ETC___d3111 ;
  assign IF_m_vrg_source_ip_7_read__7_AND_NOT_m_vrg_sou_ETC___d3168 =
	     m_vrg_source_ip_7_read__7_AND_NOT_m_vrg_source_ETC___d3115 ?
	       5'd7 :
	       (m_vrg_source_ip_6_read__6_AND_NOT_m_vrg_source_ETC___d3110 ?
		  5'd6 :
		  IF_m_vrg_source_ip_5_read__5_AND_NOT_m_vrg_sou_ETC___d3166) ;
  assign IF_m_vrg_source_ip_7_read__7_AND_NOT_m_vrg_sou_ETC___d594 =
	     m_vrg_source_ip_7_read__7_AND_NOT_m_vrg_source_ETC___d593 ?
	       m_vrg_source_prio_7 :
	       IF_m_vrg_source_ip_6_read__6_AND_NOT_m_vrg_sou_ETC___d587 ;
  assign IF_m_vrg_source_ip_7_read__7_AND_NOT_m_vrg_sou_ETC___d663 =
	     m_vrg_source_ip_7_read__7_AND_NOT_m_vrg_source_ETC___d593 ?
	       5'd7 :
	       (m_vrg_source_ip_6_read__6_AND_NOT_m_vrg_source_ETC___d586 ?
		  5'd6 :
		  IF_m_vrg_source_ip_5_read__5_AND_NOT_m_vrg_sou_ETC___d661) ;
  assign IF_m_vrg_source_ip_8_read__8_AND_NOT_m_vrg_sou_ETC___d3027 =
	     m_vrg_source_ip_8_read__8_AND_NOT_m_vrg_source_ETC___d3026 ?
	       m_vrg_source_prio_8 :
	       IF_m_vrg_source_ip_7_read__7_AND_NOT_m_vrg_sou_ETC___d3022 ;
  assign IF_m_vrg_source_ip_8_read__8_AND_NOT_m_vrg_sou_ETC___d3121 =
	     m_vrg_source_ip_8_read__8_AND_NOT_m_vrg_source_ETC___d3120 ?
	       m_vrg_source_prio_8 :
	       IF_m_vrg_source_ip_7_read__7_AND_NOT_m_vrg_sou_ETC___d3116 ;
  assign IF_m_vrg_source_ip_8_read__8_AND_NOT_m_vrg_sou_ETC___d601 =
	     m_vrg_source_ip_8_read__8_AND_NOT_m_vrg_source_ETC___d600 ?
	       m_vrg_source_prio_8 :
	       IF_m_vrg_source_ip_7_read__7_AND_NOT_m_vrg_sou_ETC___d594 ;
  assign IF_m_vrg_source_ip_9_read__9_AND_NOT_m_vrg_sou_ETC___d3032 =
	     m_vrg_source_ip_9_read__9_AND_NOT_m_vrg_source_ETC___d3031 ?
	       m_vrg_source_prio_9 :
	       IF_m_vrg_source_ip_8_read__8_AND_NOT_m_vrg_sou_ETC___d3027 ;
  assign IF_m_vrg_source_ip_9_read__9_AND_NOT_m_vrg_sou_ETC___d3076 =
	     m_vrg_source_ip_9_read__9_AND_NOT_m_vrg_source_ETC___d3031 ?
	       5'd9 :
	       (m_vrg_source_ip_8_read__8_AND_NOT_m_vrg_source_ETC___d3026 ?
		  5'd8 :
		  IF_m_vrg_source_ip_7_read__7_AND_NOT_m_vrg_sou_ETC___d3074) ;
  assign IF_m_vrg_source_ip_9_read__9_AND_NOT_m_vrg_sou_ETC___d3126 =
	     m_vrg_source_ip_9_read__9_AND_NOT_m_vrg_source_ETC___d3125 ?
	       m_vrg_source_prio_9 :
	       IF_m_vrg_source_ip_8_read__8_AND_NOT_m_vrg_sou_ETC___d3121 ;
  assign IF_m_vrg_source_ip_9_read__9_AND_NOT_m_vrg_sou_ETC___d3170 =
	     m_vrg_source_ip_9_read__9_AND_NOT_m_vrg_source_ETC___d3125 ?
	       5'd9 :
	       (m_vrg_source_ip_8_read__8_AND_NOT_m_vrg_source_ETC___d3120 ?
		  5'd8 :
		  IF_m_vrg_source_ip_7_read__7_AND_NOT_m_vrg_sou_ETC___d3168) ;
  assign IF_m_vrg_source_ip_9_read__9_AND_NOT_m_vrg_sou_ETC___d608 =
	     m_vrg_source_ip_9_read__9_AND_NOT_m_vrg_source_ETC___d607 ?
	       m_vrg_source_prio_9 :
	       IF_m_vrg_source_ip_8_read__8_AND_NOT_m_vrg_sou_ETC___d601 ;
  assign IF_m_vrg_source_ip_9_read__9_AND_NOT_m_vrg_sou_ETC___d665 =
	     m_vrg_source_ip_9_read__9_AND_NOT_m_vrg_source_ETC___d607 ?
	       5'd9 :
	       (m_vrg_source_ip_8_read__8_AND_NOT_m_vrg_source_ETC___d600 ?
		  5'd8 :
		  IF_m_vrg_source_ip_7_read__7_AND_NOT_m_vrg_sou_ETC___d663) ;
  assign NOT_m_cfg_verbosity_read_ULE_1_5___d16 = m_cfg_verbosity > 4'd1 ;
  assign NOT_m_slave_xactor_f_rd_addr_first__9_BITS_92__ETC___d248 =
	     !m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d31 &&
	     !m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d36 &&
	     !m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d68 &&
	     m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d240 &&
	     m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d71 &&
	     m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d242 &&
	     m_cfg_verbosity != 4'd0 ;
  assign NOT_m_slave_xactor_f_rd_addr_first__9_BITS_92__ETC___d538 =
	     !m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d31 &&
	     !m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d36 &&
	     !m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d68 &&
	     !m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d240 &&
	     x__h23928 == 32'h00200000 &&
	     m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d532 &&
	     m_cfg_verbosity != 4'd0 ;
  assign NOT_m_slave_xactor_f_rd_addr_first__9_BITS_92__ETC___d695 =
	     !m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d31 &&
	     !m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d36 &&
	     !m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d68 &&
	     !m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d240 &&
	     x__h23928 == 32'h00200004 &&
	     m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d532 &&
	     m_vrg_source_ip_16_read__6_AND_NOT_m_vrg_sourc_ETC___d689 ;
  assign NOT_m_slave_xactor_f_rd_addr_first__9_BITS_92__ETC___d733 =
	     !m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d31 &&
	     !m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d36 &&
	     !m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d68 &&
	     !m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d240 &&
	     x__h23928 == 32'h00200004 &&
	     m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d532 &&
	     m_cfg_verbosity != 4'd0 ;
  assign NOT_m_slave_xactor_f_rd_addr_first__9_BITS_92__ETC___d74 =
	     !m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d36 &&
	     m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d68 &&
	     m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d71 &&
	     m_cfg_verbosity != 4'd0 ;
  assign NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1017 =
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d821 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d874 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d888 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d877 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d889 &&
	     source_id__h31729 <= 10'd16 ;
  assign NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1078 =
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d821 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d874 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d888 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d877 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d889 &&
	     source_id__h33225 <= 10'd16 ;
  assign NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1139 =
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d821 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d874 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d888 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d877 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d889 &&
	     source_id__h34721 <= 10'd16 ;
  assign NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1200 =
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d821 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d874 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d888 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d877 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d889 &&
	     source_id__h36217 <= 10'd16 ;
  assign NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1261 =
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d821 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d874 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d888 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d877 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d889 &&
	     source_id__h37713 <= 10'd16 ;
  assign NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1322 =
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d821 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d874 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d888 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d877 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d889 &&
	     source_id__h39209 <= 10'd16 ;
  assign NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1383 =
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d821 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d874 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d888 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d877 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d889 &&
	     source_id__h40705 <= 10'd16 ;
  assign NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1444 =
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d821 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d874 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d888 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d877 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d889 &&
	     source_id__h42201 <= 10'd16 ;
  assign NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1505 =
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d821 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d874 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d888 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d877 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d889 &&
	     source_id__h43697 <= 10'd16 ;
  assign NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1566 =
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d821 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d874 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d888 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d877 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d889 &&
	     source_id__h45193 <= 10'd16 ;
  assign NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1627 =
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d821 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d874 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d888 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d877 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d889 &&
	     source_id__h46689 <= 10'd16 ;
  assign NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1688 =
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d821 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d874 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d888 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d877 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d889 &&
	     source_id__h48185 <= 10'd16 ;
  assign NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1749 =
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d821 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d874 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d888 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d877 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d889 &&
	     source_id__h49681 <= 10'd16 ;
  assign NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1810 =
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d821 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d874 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d888 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d877 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d889 &&
	     source_id__h51177 <= 10'd16 ;
  assign NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1871 =
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d821 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d874 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d888 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d877 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d889 &&
	     source_id__h52673 <= 10'd16 ;
  assign NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1932 =
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d821 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d874 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d888 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d877 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d889 &&
	     source_id__h54169 <= 10'd16 ;
  assign NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1993 =
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d821 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d874 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d888 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d877 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d889 &&
	     source_id__h55665 <= 10'd16 ;
  assign NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2054 =
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d821 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d874 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d888 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d877 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d889 &&
	     source_id__h57161 <= 10'd16 ;
  assign NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2115 =
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d821 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d874 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d888 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d877 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d889 &&
	     source_id__h58657 <= 10'd16 ;
  assign NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2176 =
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d821 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d874 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d888 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d877 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d889 &&
	     source_id__h60153 <= 10'd16 ;
  assign NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2237 =
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d821 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d874 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d888 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d877 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d889 &&
	     source_id__h61649 <= 10'd16 ;
  assign NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2298 =
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d821 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d874 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d888 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d877 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d889 &&
	     source_id__h63145 <= 10'd16 ;
  assign NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2359 =
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d821 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d874 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d888 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d877 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d889 &&
	     source_id__h64641 <= 10'd16 ;
  assign NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2420 =
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d821 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d874 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d888 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d877 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d889 &&
	     source_id__h66137 <= 10'd16 ;
  assign NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2481 =
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d821 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d874 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d888 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d877 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d889 &&
	     source_id__h67633 <= 10'd16 ;
  assign NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2542 =
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d821 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d874 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d888 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d877 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d889 &&
	     source_id__h69129 <= 10'd16 ;
  assign NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2603 =
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d821 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d874 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d888 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d877 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d889 &&
	     source_id__h70625 <= 10'd16 ;
  assign NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2664 =
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d821 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d874 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d888 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d877 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d889 &&
	     source_id__h72121 <= 10'd16 ;
  assign NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2725 =
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d821 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d874 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d888 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d877 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d889 &&
	     source_id__h73617 <= 10'd16 ;
  assign NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2786 =
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d821 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d874 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d888 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d877 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d889 &&
	     source_id__h75113 <= 10'd16 ;
  assign NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2844 =
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d821 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d874 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d888 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d877 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d889 &&
	     m_cfg_verbosity != 4'd0 ;
  assign NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2857 =
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d874 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d888 &&
	     x__h76716 == 32'h00200000 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d2854 ;
  assign NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2868 =
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d821 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d874 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d888 &&
	     x__h76716 == 32'h00200000 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d2854 &&
	     m_cfg_verbosity != 4'd0 ;
  assign NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2884 =
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d821 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d874 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d888 &&
	     x__h76716 == 32'h00200004 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d2854 &&
	     IF_m_slave_xactor_f_wr_addr_first__94_BITS_92__ETC___d2874 &&
	     SEL_ARR_SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_ETC___d2878 ;
  assign NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2923 =
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d874 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d888 &&
	     x__h76716 == 32'h00200004 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d2854 &&
	     IF_m_slave_xactor_f_wr_addr_first__94_BITS_92__ETC___d2874 &&
	     SEL_ARR_SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_ETC___d2878 &&
	     m_cfg_verbosity != 4'd0 ;
  assign NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2935 =
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d874 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d888 &&
	     x__h76716 == 32'h00200004 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d2854 &&
	     (!IF_m_slave_xactor_f_wr_addr_first__94_BITS_92__ETC___d2874 ||
	      !SEL_ARR_SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_ETC___d2878) &&
	     m_cfg_verbosity != 4'd0 ;
  assign NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d826 =
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d821 &&
	     addr_offset__h27245[11:2] != 10'd0 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d823 ;
  assign NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d880 =
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d821 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d874 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d877 &&
	     m_cfg_verbosity != 4'd0 ;
  assign NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d892 =
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d874 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d888 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d877 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d889 ;
  assign NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d956 =
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d821 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d874 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d888 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d877 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d889 &&
	     source_id__h30233 <= 10'd16 ;
  assign NOT_m_vrg_source_busy_10_983_284_AND_NOT_m_cfg_ETC___d3288 =
	     !m_vrg_source_busy_10 && m_cfg_verbosity != 4'd0 &&
	     m_vrg_source_ip_10 != v_sources_9_m_interrupt_req_set_not_clear ;
  assign NOT_m_vrg_source_busy_11_984_292_AND_NOT_m_cfg_ETC___d3296 =
	     !m_vrg_source_busy_11 && m_cfg_verbosity != 4'd0 &&
	     m_vrg_source_ip_11 !=
	     v_sources_10_m_interrupt_req_set_not_clear ;
  assign NOT_m_vrg_source_busy_12_985_300_AND_NOT_m_cfg_ETC___d3304 =
	     !m_vrg_source_busy_12 && m_cfg_verbosity != 4'd0 &&
	     m_vrg_source_ip_12 !=
	     v_sources_11_m_interrupt_req_set_not_clear ;
  assign NOT_m_vrg_source_busy_13_986_308_AND_NOT_m_cfg_ETC___d3312 =
	     !m_vrg_source_busy_13 && m_cfg_verbosity != 4'd0 &&
	     m_vrg_source_ip_13 !=
	     v_sources_12_m_interrupt_req_set_not_clear ;
  assign NOT_m_vrg_source_busy_14_987_316_AND_NOT_m_cfg_ETC___d3320 =
	     !m_vrg_source_busy_14 && m_cfg_verbosity != 4'd0 &&
	     m_vrg_source_ip_14 !=
	     v_sources_13_m_interrupt_req_set_not_clear ;
  assign NOT_m_vrg_source_busy_15_988_324_AND_NOT_m_cfg_ETC___d3328 =
	     !m_vrg_source_busy_15 && m_cfg_verbosity != 4'd0 &&
	     m_vrg_source_ip_15 !=
	     v_sources_14_m_interrupt_req_set_not_clear ;
  assign NOT_m_vrg_source_busy_16_989_332_AND_NOT_m_cfg_ETC___d3336 =
	     !m_vrg_source_busy_16 && m_cfg_verbosity != 4'd0 &&
	     m_vrg_source_ip_16 !=
	     v_sources_15_m_interrupt_req_set_not_clear ;
  assign NOT_m_vrg_source_busy_1_974_213_AND_NOT_m_cfg__ETC___d3217 =
	     !m_vrg_source_busy_1 && m_cfg_verbosity != 4'd0 &&
	     m_vrg_source_ip_1 != v_sources_0_m_interrupt_req_set_not_clear ;
  assign NOT_m_vrg_source_busy_2_975_220_AND_NOT_m_cfg__ETC___d3224 =
	     !m_vrg_source_busy_2 && m_cfg_verbosity != 4'd0 &&
	     m_vrg_source_ip_2 != v_sources_1_m_interrupt_req_set_not_clear ;
  assign NOT_m_vrg_source_busy_3_976_228_AND_NOT_m_cfg__ETC___d3232 =
	     !m_vrg_source_busy_3 && m_cfg_verbosity != 4'd0 &&
	     m_vrg_source_ip_3 != v_sources_2_m_interrupt_req_set_not_clear ;
  assign NOT_m_vrg_source_busy_4_977_236_AND_NOT_m_cfg__ETC___d3240 =
	     !m_vrg_source_busy_4 && m_cfg_verbosity != 4'd0 &&
	     m_vrg_source_ip_4 != v_sources_3_m_interrupt_req_set_not_clear ;
  assign NOT_m_vrg_source_busy_5_978_244_AND_NOT_m_cfg__ETC___d3248 =
	     !m_vrg_source_busy_5 && m_cfg_verbosity != 4'd0 &&
	     m_vrg_source_ip_5 != v_sources_4_m_interrupt_req_set_not_clear ;
  assign NOT_m_vrg_source_busy_6_979_252_AND_NOT_m_cfg__ETC___d3256 =
	     !m_vrg_source_busy_6 && m_cfg_verbosity != 4'd0 &&
	     m_vrg_source_ip_6 != v_sources_5_m_interrupt_req_set_not_clear ;
  assign NOT_m_vrg_source_busy_7_980_260_AND_NOT_m_cfg__ETC___d3264 =
	     !m_vrg_source_busy_7 && m_cfg_verbosity != 4'd0 &&
	     m_vrg_source_ip_7 != v_sources_6_m_interrupt_req_set_not_clear ;
  assign NOT_m_vrg_source_busy_8_981_268_AND_NOT_m_cfg__ETC___d3272 =
	     !m_vrg_source_busy_8 && m_cfg_verbosity != 4'd0 &&
	     m_vrg_source_ip_8 != v_sources_7_m_interrupt_req_set_not_clear ;
  assign NOT_m_vrg_source_busy_9_982_276_AND_NOT_m_cfg__ETC___d3280 =
	     !m_vrg_source_busy_9 && m_cfg_verbosity != 4'd0 &&
	     m_vrg_source_ip_9 != v_sources_8_m_interrupt_req_set_not_clear ;
  assign _dfoo1 =
	     source_id__h73617 == 10'd16 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2725 ||
	     source_id__h75113 == 10'd16 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2786 ;
  assign _dfoo10 =
	     (source_id__h73617 == 10'd12 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2725) ?
	       wdata32__h27246[30] :
	       wdata32__h27246[31] ;
  assign _dfoo100 =
	     (source_id__h72121 == 10'd1 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2664) ?
	       wdata32__h27246[29] :
	       _dfoo32 ;
  assign _dfoo1000 =
	     (source_id__h52673 == 10'd10 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1871) ?
	       wdata32__h27246[16] :
	       _dfoo932 ;
  assign _dfoo1001 =
	     source_id__h52673 == 10'd9 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1871 ||
	     source_id__h54169 == 10'd9 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1932 ||
	     _dfoo865 ;
  assign _dfoo1002 =
	     (source_id__h52673 == 10'd9 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1871) ?
	       wdata32__h27246[16] :
	       _dfoo934 ;
  assign _dfoo1003 =
	     source_id__h52673 == 10'd8 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1871 ||
	     source_id__h54169 == 10'd8 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1932 ||
	     _dfoo867 ;
  assign _dfoo1004 =
	     (source_id__h52673 == 10'd8 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1871) ?
	       wdata32__h27246[16] :
	       _dfoo936 ;
  assign _dfoo1005 =
	     source_id__h52673 == 10'd7 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1871 ||
	     source_id__h54169 == 10'd7 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1932 ||
	     _dfoo869 ;
  assign _dfoo1006 =
	     (source_id__h52673 == 10'd7 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1871) ?
	       wdata32__h27246[16] :
	       _dfoo938 ;
  assign _dfoo1007 =
	     source_id__h52673 == 10'd6 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1871 ||
	     source_id__h54169 == 10'd6 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1932 ||
	     _dfoo871 ;
  assign _dfoo1008 =
	     (source_id__h52673 == 10'd6 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1871) ?
	       wdata32__h27246[16] :
	       _dfoo940 ;
  assign _dfoo1009 =
	     source_id__h52673 == 10'd5 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1871 ||
	     source_id__h54169 == 10'd5 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1932 ||
	     _dfoo873 ;
  assign _dfoo1010 =
	     (source_id__h52673 == 10'd5 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1871) ?
	       wdata32__h27246[16] :
	       _dfoo942 ;
  assign _dfoo1011 =
	     source_id__h52673 == 10'd4 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1871 ||
	     source_id__h54169 == 10'd4 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1932 ||
	     _dfoo875 ;
  assign _dfoo1012 =
	     (source_id__h52673 == 10'd4 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1871) ?
	       wdata32__h27246[16] :
	       _dfoo944 ;
  assign _dfoo1013 =
	     source_id__h52673 == 10'd3 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1871 ||
	     source_id__h54169 == 10'd3 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1932 ||
	     _dfoo877 ;
  assign _dfoo1014 =
	     (source_id__h52673 == 10'd3 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1871) ?
	       wdata32__h27246[16] :
	       _dfoo946 ;
  assign _dfoo1015 =
	     source_id__h52673 == 10'd2 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1871 ||
	     source_id__h54169 == 10'd2 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1932 ||
	     _dfoo879 ;
  assign _dfoo1016 =
	     (source_id__h52673 == 10'd2 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1871) ?
	       wdata32__h27246[16] :
	       _dfoo948 ;
  assign _dfoo1017 =
	     source_id__h52673 == 10'd1 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1871 ||
	     source_id__h54169 == 10'd1 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1932 ||
	     _dfoo881 ;
  assign _dfoo1018 =
	     (source_id__h52673 == 10'd1 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1871) ?
	       wdata32__h27246[16] :
	       _dfoo950 ;
  assign _dfoo1019 =
	     source_id__h52673 == 10'd0 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1871 ||
	     source_id__h54169 == 10'd0 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1932 ||
	     _dfoo883 ;
  assign _dfoo102 =
	     (source_id__h72121 == 10'd0 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2664) ?
	       wdata32__h27246[29] :
	       _dfoo34 ;
  assign _dfoo1020 =
	     (source_id__h52673 == 10'd0 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1871) ?
	       wdata32__h27246[16] :
	       _dfoo952 ;
  assign _dfoo1022 =
	     (source_id__h51177 == 10'd16 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1810) ?
	       wdata32__h27246[15] :
	       _dfoo954 ;
  assign _dfoo1024 =
	     (source_id__h51177 == 10'd15 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1810) ?
	       wdata32__h27246[15] :
	       _dfoo956 ;
  assign _dfoo1026 =
	     (source_id__h51177 == 10'd14 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1810) ?
	       wdata32__h27246[15] :
	       _dfoo958 ;
  assign _dfoo1028 =
	     (source_id__h51177 == 10'd13 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1810) ?
	       wdata32__h27246[15] :
	       _dfoo960 ;
  assign _dfoo1030 =
	     (source_id__h51177 == 10'd12 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1810) ?
	       wdata32__h27246[15] :
	       _dfoo962 ;
  assign _dfoo1032 =
	     (source_id__h51177 == 10'd11 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1810) ?
	       wdata32__h27246[15] :
	       _dfoo964 ;
  assign _dfoo1034 =
	     (source_id__h51177 == 10'd10 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1810) ?
	       wdata32__h27246[15] :
	       _dfoo966 ;
  assign _dfoo1036 =
	     (source_id__h51177 == 10'd9 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1810) ?
	       wdata32__h27246[15] :
	       _dfoo968 ;
  assign _dfoo1038 =
	     (source_id__h51177 == 10'd8 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1810) ?
	       wdata32__h27246[15] :
	       _dfoo970 ;
  assign _dfoo104 =
	     (source_id__h72121 == 10'd16 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2664) ?
	       wdata32__h27246[29] :
	       _dfoo36 ;
  assign _dfoo1040 =
	     (source_id__h51177 == 10'd7 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1810) ?
	       wdata32__h27246[15] :
	       _dfoo972 ;
  assign _dfoo1042 =
	     (source_id__h51177 == 10'd6 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1810) ?
	       wdata32__h27246[15] :
	       _dfoo974 ;
  assign _dfoo1044 =
	     (source_id__h51177 == 10'd5 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1810) ?
	       wdata32__h27246[15] :
	       _dfoo976 ;
  assign _dfoo1046 =
	     (source_id__h51177 == 10'd4 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1810) ?
	       wdata32__h27246[15] :
	       _dfoo978 ;
  assign _dfoo1048 =
	     (source_id__h51177 == 10'd3 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1810) ?
	       wdata32__h27246[15] :
	       _dfoo980 ;
  assign _dfoo1050 =
	     (source_id__h51177 == 10'd2 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1810) ?
	       wdata32__h27246[15] :
	       _dfoo982 ;
  assign _dfoo1052 =
	     (source_id__h51177 == 10'd1 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1810) ?
	       wdata32__h27246[15] :
	       _dfoo984 ;
  assign _dfoo1054 =
	     (source_id__h51177 == 10'd0 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1810) ?
	       wdata32__h27246[15] :
	       _dfoo986 ;
  assign _dfoo1056 =
	     (source_id__h51177 == 10'd16 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1810) ?
	       wdata32__h27246[15] :
	       _dfoo988 ;
  assign _dfoo1058 =
	     (source_id__h51177 == 10'd15 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1810) ?
	       wdata32__h27246[15] :
	       _dfoo990 ;
  assign _dfoo106 =
	     (source_id__h72121 == 10'd15 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2664) ?
	       wdata32__h27246[29] :
	       _dfoo38 ;
  assign _dfoo1060 =
	     (source_id__h51177 == 10'd14 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1810) ?
	       wdata32__h27246[15] :
	       _dfoo992 ;
  assign _dfoo1062 =
	     (source_id__h51177 == 10'd13 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1810) ?
	       wdata32__h27246[15] :
	       _dfoo994 ;
  assign _dfoo1064 =
	     (source_id__h51177 == 10'd12 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1810) ?
	       wdata32__h27246[15] :
	       _dfoo996 ;
  assign _dfoo1066 =
	     (source_id__h51177 == 10'd11 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1810) ?
	       wdata32__h27246[15] :
	       _dfoo998 ;
  assign _dfoo1068 =
	     (source_id__h51177 == 10'd10 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1810) ?
	       wdata32__h27246[15] :
	       _dfoo1000 ;
  assign _dfoo1070 =
	     (source_id__h51177 == 10'd9 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1810) ?
	       wdata32__h27246[15] :
	       _dfoo1002 ;
  assign _dfoo1072 =
	     (source_id__h51177 == 10'd8 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1810) ?
	       wdata32__h27246[15] :
	       _dfoo1004 ;
  assign _dfoo1074 =
	     (source_id__h51177 == 10'd7 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1810) ?
	       wdata32__h27246[15] :
	       _dfoo1006 ;
  assign _dfoo1076 =
	     (source_id__h51177 == 10'd6 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1810) ?
	       wdata32__h27246[15] :
	       _dfoo1008 ;
  assign _dfoo1078 =
	     (source_id__h51177 == 10'd5 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1810) ?
	       wdata32__h27246[15] :
	       _dfoo1010 ;
  assign _dfoo108 =
	     (source_id__h72121 == 10'd14 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2664) ?
	       wdata32__h27246[29] :
	       _dfoo40 ;
  assign _dfoo1080 =
	     (source_id__h51177 == 10'd4 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1810) ?
	       wdata32__h27246[15] :
	       _dfoo1012 ;
  assign _dfoo1082 =
	     (source_id__h51177 == 10'd3 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1810) ?
	       wdata32__h27246[15] :
	       _dfoo1014 ;
  assign _dfoo1084 =
	     (source_id__h51177 == 10'd2 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1810) ?
	       wdata32__h27246[15] :
	       _dfoo1016 ;
  assign _dfoo1086 =
	     (source_id__h51177 == 10'd1 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1810) ?
	       wdata32__h27246[15] :
	       _dfoo1018 ;
  assign _dfoo1088 =
	     (source_id__h51177 == 10'd0 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1810) ?
	       wdata32__h27246[15] :
	       _dfoo1020 ;
  assign _dfoo1089 =
	     source_id__h49681 == 10'd16 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1749 ||
	     source_id__h51177 == 10'd16 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1810 ||
	     _dfoo953 ;
  assign _dfoo1090 =
	     (source_id__h49681 == 10'd16 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1749) ?
	       wdata32__h27246[14] :
	       _dfoo1022 ;
  assign _dfoo1091 =
	     source_id__h49681 == 10'd15 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1749 ||
	     source_id__h51177 == 10'd15 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1810 ||
	     _dfoo955 ;
  assign _dfoo1092 =
	     (source_id__h49681 == 10'd15 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1749) ?
	       wdata32__h27246[14] :
	       _dfoo1024 ;
  assign _dfoo1093 =
	     source_id__h49681 == 10'd14 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1749 ||
	     source_id__h51177 == 10'd14 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1810 ||
	     _dfoo957 ;
  assign _dfoo1094 =
	     (source_id__h49681 == 10'd14 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1749) ?
	       wdata32__h27246[14] :
	       _dfoo1026 ;
  assign _dfoo1095 =
	     source_id__h49681 == 10'd13 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1749 ||
	     source_id__h51177 == 10'd13 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1810 ||
	     _dfoo959 ;
  assign _dfoo1096 =
	     (source_id__h49681 == 10'd13 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1749) ?
	       wdata32__h27246[14] :
	       _dfoo1028 ;
  assign _dfoo1097 =
	     source_id__h49681 == 10'd12 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1749 ||
	     source_id__h51177 == 10'd12 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1810 ||
	     _dfoo961 ;
  assign _dfoo1098 =
	     (source_id__h49681 == 10'd12 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1749) ?
	       wdata32__h27246[14] :
	       _dfoo1030 ;
  assign _dfoo1099 =
	     source_id__h49681 == 10'd11 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1749 ||
	     source_id__h51177 == 10'd11 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1810 ||
	     _dfoo963 ;
  assign _dfoo11 =
	     source_id__h73617 == 10'd11 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2725 ||
	     source_id__h75113 == 10'd11 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2786 ;
  assign _dfoo110 =
	     (source_id__h72121 == 10'd13 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2664) ?
	       wdata32__h27246[29] :
	       _dfoo42 ;
  assign _dfoo1100 =
	     (source_id__h49681 == 10'd11 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1749) ?
	       wdata32__h27246[14] :
	       _dfoo1032 ;
  assign _dfoo1101 =
	     source_id__h49681 == 10'd10 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1749 ||
	     source_id__h51177 == 10'd10 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1810 ||
	     _dfoo965 ;
  assign _dfoo1102 =
	     (source_id__h49681 == 10'd10 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1749) ?
	       wdata32__h27246[14] :
	       _dfoo1034 ;
  assign _dfoo1103 =
	     source_id__h49681 == 10'd9 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1749 ||
	     source_id__h51177 == 10'd9 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1810 ||
	     _dfoo967 ;
  assign _dfoo1104 =
	     (source_id__h49681 == 10'd9 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1749) ?
	       wdata32__h27246[14] :
	       _dfoo1036 ;
  assign _dfoo1105 =
	     source_id__h49681 == 10'd8 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1749 ||
	     source_id__h51177 == 10'd8 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1810 ||
	     _dfoo969 ;
  assign _dfoo1106 =
	     (source_id__h49681 == 10'd8 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1749) ?
	       wdata32__h27246[14] :
	       _dfoo1038 ;
  assign _dfoo1107 =
	     source_id__h49681 == 10'd7 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1749 ||
	     source_id__h51177 == 10'd7 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1810 ||
	     _dfoo971 ;
  assign _dfoo1108 =
	     (source_id__h49681 == 10'd7 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1749) ?
	       wdata32__h27246[14] :
	       _dfoo1040 ;
  assign _dfoo1109 =
	     source_id__h49681 == 10'd6 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1749 ||
	     source_id__h51177 == 10'd6 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1810 ||
	     _dfoo973 ;
  assign _dfoo1110 =
	     (source_id__h49681 == 10'd6 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1749) ?
	       wdata32__h27246[14] :
	       _dfoo1042 ;
  assign _dfoo1111 =
	     source_id__h49681 == 10'd5 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1749 ||
	     source_id__h51177 == 10'd5 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1810 ||
	     _dfoo975 ;
  assign _dfoo1112 =
	     (source_id__h49681 == 10'd5 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1749) ?
	       wdata32__h27246[14] :
	       _dfoo1044 ;
  assign _dfoo1113 =
	     source_id__h49681 == 10'd4 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1749 ||
	     source_id__h51177 == 10'd4 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1810 ||
	     _dfoo977 ;
  assign _dfoo1114 =
	     (source_id__h49681 == 10'd4 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1749) ?
	       wdata32__h27246[14] :
	       _dfoo1046 ;
  assign _dfoo1115 =
	     source_id__h49681 == 10'd3 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1749 ||
	     source_id__h51177 == 10'd3 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1810 ||
	     _dfoo979 ;
  assign _dfoo1116 =
	     (source_id__h49681 == 10'd3 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1749) ?
	       wdata32__h27246[14] :
	       _dfoo1048 ;
  assign _dfoo1117 =
	     source_id__h49681 == 10'd2 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1749 ||
	     source_id__h51177 == 10'd2 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1810 ||
	     _dfoo981 ;
  assign _dfoo1118 =
	     (source_id__h49681 == 10'd2 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1749) ?
	       wdata32__h27246[14] :
	       _dfoo1050 ;
  assign _dfoo1119 =
	     source_id__h49681 == 10'd1 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1749 ||
	     source_id__h51177 == 10'd1 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1810 ||
	     _dfoo983 ;
  assign _dfoo112 =
	     (source_id__h72121 == 10'd12 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2664) ?
	       wdata32__h27246[29] :
	       _dfoo44 ;
  assign _dfoo1120 =
	     (source_id__h49681 == 10'd1 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1749) ?
	       wdata32__h27246[14] :
	       _dfoo1052 ;
  assign _dfoo1121 =
	     source_id__h49681 == 10'd0 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1749 ||
	     source_id__h51177 == 10'd0 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1810 ||
	     _dfoo985 ;
  assign _dfoo1122 =
	     (source_id__h49681 == 10'd0 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1749) ?
	       wdata32__h27246[14] :
	       _dfoo1054 ;
  assign _dfoo1123 =
	     source_id__h49681 == 10'd16 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1749 ||
	     source_id__h51177 == 10'd16 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1810 ||
	     _dfoo987 ;
  assign _dfoo1124 =
	     (source_id__h49681 == 10'd16 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1749) ?
	       wdata32__h27246[14] :
	       _dfoo1056 ;
  assign _dfoo1125 =
	     source_id__h49681 == 10'd15 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1749 ||
	     source_id__h51177 == 10'd15 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1810 ||
	     _dfoo989 ;
  assign _dfoo1126 =
	     (source_id__h49681 == 10'd15 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1749) ?
	       wdata32__h27246[14] :
	       _dfoo1058 ;
  assign _dfoo1127 =
	     source_id__h49681 == 10'd14 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1749 ||
	     source_id__h51177 == 10'd14 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1810 ||
	     _dfoo991 ;
  assign _dfoo1128 =
	     (source_id__h49681 == 10'd14 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1749) ?
	       wdata32__h27246[14] :
	       _dfoo1060 ;
  assign _dfoo1129 =
	     source_id__h49681 == 10'd13 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1749 ||
	     source_id__h51177 == 10'd13 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1810 ||
	     _dfoo993 ;
  assign _dfoo1130 =
	     (source_id__h49681 == 10'd13 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1749) ?
	       wdata32__h27246[14] :
	       _dfoo1062 ;
  assign _dfoo1131 =
	     source_id__h49681 == 10'd12 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1749 ||
	     source_id__h51177 == 10'd12 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1810 ||
	     _dfoo995 ;
  assign _dfoo1132 =
	     (source_id__h49681 == 10'd12 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1749) ?
	       wdata32__h27246[14] :
	       _dfoo1064 ;
  assign _dfoo1133 =
	     source_id__h49681 == 10'd11 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1749 ||
	     source_id__h51177 == 10'd11 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1810 ||
	     _dfoo997 ;
  assign _dfoo1134 =
	     (source_id__h49681 == 10'd11 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1749) ?
	       wdata32__h27246[14] :
	       _dfoo1066 ;
  assign _dfoo1135 =
	     source_id__h49681 == 10'd10 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1749 ||
	     source_id__h51177 == 10'd10 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1810 ||
	     _dfoo999 ;
  assign _dfoo1136 =
	     (source_id__h49681 == 10'd10 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1749) ?
	       wdata32__h27246[14] :
	       _dfoo1068 ;
  assign _dfoo1137 =
	     source_id__h49681 == 10'd9 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1749 ||
	     source_id__h51177 == 10'd9 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1810 ||
	     _dfoo1001 ;
  assign _dfoo1138 =
	     (source_id__h49681 == 10'd9 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1749) ?
	       wdata32__h27246[14] :
	       _dfoo1070 ;
  assign _dfoo1139 =
	     source_id__h49681 == 10'd8 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1749 ||
	     source_id__h51177 == 10'd8 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1810 ||
	     _dfoo1003 ;
  assign _dfoo114 =
	     (source_id__h72121 == 10'd11 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2664) ?
	       wdata32__h27246[29] :
	       _dfoo46 ;
  assign _dfoo1140 =
	     (source_id__h49681 == 10'd8 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1749) ?
	       wdata32__h27246[14] :
	       _dfoo1072 ;
  assign _dfoo1141 =
	     source_id__h49681 == 10'd7 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1749 ||
	     source_id__h51177 == 10'd7 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1810 ||
	     _dfoo1005 ;
  assign _dfoo1142 =
	     (source_id__h49681 == 10'd7 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1749) ?
	       wdata32__h27246[14] :
	       _dfoo1074 ;
  assign _dfoo1143 =
	     source_id__h49681 == 10'd6 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1749 ||
	     source_id__h51177 == 10'd6 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1810 ||
	     _dfoo1007 ;
  assign _dfoo1144 =
	     (source_id__h49681 == 10'd6 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1749) ?
	       wdata32__h27246[14] :
	       _dfoo1076 ;
  assign _dfoo1145 =
	     source_id__h49681 == 10'd5 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1749 ||
	     source_id__h51177 == 10'd5 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1810 ||
	     _dfoo1009 ;
  assign _dfoo1146 =
	     (source_id__h49681 == 10'd5 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1749) ?
	       wdata32__h27246[14] :
	       _dfoo1078 ;
  assign _dfoo1147 =
	     source_id__h49681 == 10'd4 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1749 ||
	     source_id__h51177 == 10'd4 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1810 ||
	     _dfoo1011 ;
  assign _dfoo1148 =
	     (source_id__h49681 == 10'd4 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1749) ?
	       wdata32__h27246[14] :
	       _dfoo1080 ;
  assign _dfoo1149 =
	     source_id__h49681 == 10'd3 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1749 ||
	     source_id__h51177 == 10'd3 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1810 ||
	     _dfoo1013 ;
  assign _dfoo1150 =
	     (source_id__h49681 == 10'd3 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1749) ?
	       wdata32__h27246[14] :
	       _dfoo1082 ;
  assign _dfoo1151 =
	     source_id__h49681 == 10'd2 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1749 ||
	     source_id__h51177 == 10'd2 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1810 ||
	     _dfoo1015 ;
  assign _dfoo1152 =
	     (source_id__h49681 == 10'd2 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1749) ?
	       wdata32__h27246[14] :
	       _dfoo1084 ;
  assign _dfoo1153 =
	     source_id__h49681 == 10'd1 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1749 ||
	     source_id__h51177 == 10'd1 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1810 ||
	     _dfoo1017 ;
  assign _dfoo1154 =
	     (source_id__h49681 == 10'd1 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1749) ?
	       wdata32__h27246[14] :
	       _dfoo1086 ;
  assign _dfoo1155 =
	     source_id__h49681 == 10'd0 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1749 ||
	     source_id__h51177 == 10'd0 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1810 ||
	     _dfoo1019 ;
  assign _dfoo1156 =
	     (source_id__h49681 == 10'd0 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1749) ?
	       wdata32__h27246[14] :
	       _dfoo1088 ;
  assign _dfoo1158 =
	     (source_id__h48185 == 10'd16 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1688) ?
	       wdata32__h27246[13] :
	       _dfoo1090 ;
  assign _dfoo116 =
	     (source_id__h72121 == 10'd10 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2664) ?
	       wdata32__h27246[29] :
	       _dfoo48 ;
  assign _dfoo1160 =
	     (source_id__h48185 == 10'd15 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1688) ?
	       wdata32__h27246[13] :
	       _dfoo1092 ;
  assign _dfoo1162 =
	     (source_id__h48185 == 10'd14 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1688) ?
	       wdata32__h27246[13] :
	       _dfoo1094 ;
  assign _dfoo1164 =
	     (source_id__h48185 == 10'd13 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1688) ?
	       wdata32__h27246[13] :
	       _dfoo1096 ;
  assign _dfoo1166 =
	     (source_id__h48185 == 10'd12 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1688) ?
	       wdata32__h27246[13] :
	       _dfoo1098 ;
  assign _dfoo1168 =
	     (source_id__h48185 == 10'd11 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1688) ?
	       wdata32__h27246[13] :
	       _dfoo1100 ;
  assign _dfoo1170 =
	     (source_id__h48185 == 10'd10 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1688) ?
	       wdata32__h27246[13] :
	       _dfoo1102 ;
  assign _dfoo1172 =
	     (source_id__h48185 == 10'd9 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1688) ?
	       wdata32__h27246[13] :
	       _dfoo1104 ;
  assign _dfoo1174 =
	     (source_id__h48185 == 10'd8 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1688) ?
	       wdata32__h27246[13] :
	       _dfoo1106 ;
  assign _dfoo1176 =
	     (source_id__h48185 == 10'd7 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1688) ?
	       wdata32__h27246[13] :
	       _dfoo1108 ;
  assign _dfoo1178 =
	     (source_id__h48185 == 10'd6 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1688) ?
	       wdata32__h27246[13] :
	       _dfoo1110 ;
  assign _dfoo118 =
	     (source_id__h72121 == 10'd9 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2664) ?
	       wdata32__h27246[29] :
	       _dfoo50 ;
  assign _dfoo1180 =
	     (source_id__h48185 == 10'd5 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1688) ?
	       wdata32__h27246[13] :
	       _dfoo1112 ;
  assign _dfoo1182 =
	     (source_id__h48185 == 10'd4 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1688) ?
	       wdata32__h27246[13] :
	       _dfoo1114 ;
  assign _dfoo1184 =
	     (source_id__h48185 == 10'd3 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1688) ?
	       wdata32__h27246[13] :
	       _dfoo1116 ;
  assign _dfoo1186 =
	     (source_id__h48185 == 10'd2 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1688) ?
	       wdata32__h27246[13] :
	       _dfoo1118 ;
  assign _dfoo1188 =
	     (source_id__h48185 == 10'd1 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1688) ?
	       wdata32__h27246[13] :
	       _dfoo1120 ;
  assign _dfoo1190 =
	     (source_id__h48185 == 10'd0 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1688) ?
	       wdata32__h27246[13] :
	       _dfoo1122 ;
  assign _dfoo1192 =
	     (source_id__h48185 == 10'd16 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1688) ?
	       wdata32__h27246[13] :
	       _dfoo1124 ;
  assign _dfoo1194 =
	     (source_id__h48185 == 10'd15 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1688) ?
	       wdata32__h27246[13] :
	       _dfoo1126 ;
  assign _dfoo1196 =
	     (source_id__h48185 == 10'd14 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1688) ?
	       wdata32__h27246[13] :
	       _dfoo1128 ;
  assign _dfoo1198 =
	     (source_id__h48185 == 10'd13 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1688) ?
	       wdata32__h27246[13] :
	       _dfoo1130 ;
  assign _dfoo12 =
	     (source_id__h73617 == 10'd11 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2725) ?
	       wdata32__h27246[30] :
	       wdata32__h27246[31] ;
  assign _dfoo120 =
	     (source_id__h72121 == 10'd8 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2664) ?
	       wdata32__h27246[29] :
	       _dfoo52 ;
  assign _dfoo1200 =
	     (source_id__h48185 == 10'd12 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1688) ?
	       wdata32__h27246[13] :
	       _dfoo1132 ;
  assign _dfoo1202 =
	     (source_id__h48185 == 10'd11 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1688) ?
	       wdata32__h27246[13] :
	       _dfoo1134 ;
  assign _dfoo1204 =
	     (source_id__h48185 == 10'd10 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1688) ?
	       wdata32__h27246[13] :
	       _dfoo1136 ;
  assign _dfoo1206 =
	     (source_id__h48185 == 10'd9 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1688) ?
	       wdata32__h27246[13] :
	       _dfoo1138 ;
  assign _dfoo1208 =
	     (source_id__h48185 == 10'd8 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1688) ?
	       wdata32__h27246[13] :
	       _dfoo1140 ;
  assign _dfoo1210 =
	     (source_id__h48185 == 10'd7 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1688) ?
	       wdata32__h27246[13] :
	       _dfoo1142 ;
  assign _dfoo1212 =
	     (source_id__h48185 == 10'd6 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1688) ?
	       wdata32__h27246[13] :
	       _dfoo1144 ;
  assign _dfoo1214 =
	     (source_id__h48185 == 10'd5 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1688) ?
	       wdata32__h27246[13] :
	       _dfoo1146 ;
  assign _dfoo1216 =
	     (source_id__h48185 == 10'd4 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1688) ?
	       wdata32__h27246[13] :
	       _dfoo1148 ;
  assign _dfoo1218 =
	     (source_id__h48185 == 10'd3 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1688) ?
	       wdata32__h27246[13] :
	       _dfoo1150 ;
  assign _dfoo122 =
	     (source_id__h72121 == 10'd7 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2664) ?
	       wdata32__h27246[29] :
	       _dfoo54 ;
  assign _dfoo1220 =
	     (source_id__h48185 == 10'd2 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1688) ?
	       wdata32__h27246[13] :
	       _dfoo1152 ;
  assign _dfoo1222 =
	     (source_id__h48185 == 10'd1 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1688) ?
	       wdata32__h27246[13] :
	       _dfoo1154 ;
  assign _dfoo1224 =
	     (source_id__h48185 == 10'd0 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1688) ?
	       wdata32__h27246[13] :
	       _dfoo1156 ;
  assign _dfoo1225 =
	     source_id__h46689 == 10'd16 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1627 ||
	     source_id__h48185 == 10'd16 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1688 ||
	     _dfoo1089 ;
  assign _dfoo1226 =
	     (source_id__h46689 == 10'd16 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1627) ?
	       wdata32__h27246[12] :
	       _dfoo1158 ;
  assign _dfoo1227 =
	     source_id__h46689 == 10'd15 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1627 ||
	     source_id__h48185 == 10'd15 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1688 ||
	     _dfoo1091 ;
  assign _dfoo1228 =
	     (source_id__h46689 == 10'd15 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1627) ?
	       wdata32__h27246[12] :
	       _dfoo1160 ;
  assign _dfoo1229 =
	     source_id__h46689 == 10'd14 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1627 ||
	     source_id__h48185 == 10'd14 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1688 ||
	     _dfoo1093 ;
  assign _dfoo1230 =
	     (source_id__h46689 == 10'd14 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1627) ?
	       wdata32__h27246[12] :
	       _dfoo1162 ;
  assign _dfoo1231 =
	     source_id__h46689 == 10'd13 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1627 ||
	     source_id__h48185 == 10'd13 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1688 ||
	     _dfoo1095 ;
  assign _dfoo1232 =
	     (source_id__h46689 == 10'd13 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1627) ?
	       wdata32__h27246[12] :
	       _dfoo1164 ;
  assign _dfoo1233 =
	     source_id__h46689 == 10'd12 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1627 ||
	     source_id__h48185 == 10'd12 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1688 ||
	     _dfoo1097 ;
  assign _dfoo1234 =
	     (source_id__h46689 == 10'd12 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1627) ?
	       wdata32__h27246[12] :
	       _dfoo1166 ;
  assign _dfoo1235 =
	     source_id__h46689 == 10'd11 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1627 ||
	     source_id__h48185 == 10'd11 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1688 ||
	     _dfoo1099 ;
  assign _dfoo1236 =
	     (source_id__h46689 == 10'd11 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1627) ?
	       wdata32__h27246[12] :
	       _dfoo1168 ;
  assign _dfoo1237 =
	     source_id__h46689 == 10'd10 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1627 ||
	     source_id__h48185 == 10'd10 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1688 ||
	     _dfoo1101 ;
  assign _dfoo1238 =
	     (source_id__h46689 == 10'd10 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1627) ?
	       wdata32__h27246[12] :
	       _dfoo1170 ;
  assign _dfoo1239 =
	     source_id__h46689 == 10'd9 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1627 ||
	     source_id__h48185 == 10'd9 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1688 ||
	     _dfoo1103 ;
  assign _dfoo124 =
	     (source_id__h72121 == 10'd6 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2664) ?
	       wdata32__h27246[29] :
	       _dfoo56 ;
  assign _dfoo1240 =
	     (source_id__h46689 == 10'd9 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1627) ?
	       wdata32__h27246[12] :
	       _dfoo1172 ;
  assign _dfoo1241 =
	     source_id__h46689 == 10'd8 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1627 ||
	     source_id__h48185 == 10'd8 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1688 ||
	     _dfoo1105 ;
  assign _dfoo1242 =
	     (source_id__h46689 == 10'd8 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1627) ?
	       wdata32__h27246[12] :
	       _dfoo1174 ;
  assign _dfoo1243 =
	     source_id__h46689 == 10'd7 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1627 ||
	     source_id__h48185 == 10'd7 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1688 ||
	     _dfoo1107 ;
  assign _dfoo1244 =
	     (source_id__h46689 == 10'd7 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1627) ?
	       wdata32__h27246[12] :
	       _dfoo1176 ;
  assign _dfoo1245 =
	     source_id__h46689 == 10'd6 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1627 ||
	     source_id__h48185 == 10'd6 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1688 ||
	     _dfoo1109 ;
  assign _dfoo1246 =
	     (source_id__h46689 == 10'd6 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1627) ?
	       wdata32__h27246[12] :
	       _dfoo1178 ;
  assign _dfoo1247 =
	     source_id__h46689 == 10'd5 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1627 ||
	     source_id__h48185 == 10'd5 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1688 ||
	     _dfoo1111 ;
  assign _dfoo1248 =
	     (source_id__h46689 == 10'd5 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1627) ?
	       wdata32__h27246[12] :
	       _dfoo1180 ;
  assign _dfoo1249 =
	     source_id__h46689 == 10'd4 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1627 ||
	     source_id__h48185 == 10'd4 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1688 ||
	     _dfoo1113 ;
  assign _dfoo1250 =
	     (source_id__h46689 == 10'd4 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1627) ?
	       wdata32__h27246[12] :
	       _dfoo1182 ;
  assign _dfoo1251 =
	     source_id__h46689 == 10'd3 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1627 ||
	     source_id__h48185 == 10'd3 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1688 ||
	     _dfoo1115 ;
  assign _dfoo1252 =
	     (source_id__h46689 == 10'd3 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1627) ?
	       wdata32__h27246[12] :
	       _dfoo1184 ;
  assign _dfoo1253 =
	     source_id__h46689 == 10'd2 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1627 ||
	     source_id__h48185 == 10'd2 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1688 ||
	     _dfoo1117 ;
  assign _dfoo1254 =
	     (source_id__h46689 == 10'd2 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1627) ?
	       wdata32__h27246[12] :
	       _dfoo1186 ;
  assign _dfoo1255 =
	     source_id__h46689 == 10'd1 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1627 ||
	     source_id__h48185 == 10'd1 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1688 ||
	     _dfoo1119 ;
  assign _dfoo1256 =
	     (source_id__h46689 == 10'd1 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1627) ?
	       wdata32__h27246[12] :
	       _dfoo1188 ;
  assign _dfoo1257 =
	     source_id__h46689 == 10'd0 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1627 ||
	     source_id__h48185 == 10'd0 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1688 ||
	     _dfoo1121 ;
  assign _dfoo1258 =
	     (source_id__h46689 == 10'd0 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1627) ?
	       wdata32__h27246[12] :
	       _dfoo1190 ;
  assign _dfoo1259 =
	     source_id__h46689 == 10'd16 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1627 ||
	     source_id__h48185 == 10'd16 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1688 ||
	     _dfoo1123 ;
  assign _dfoo126 =
	     (source_id__h72121 == 10'd5 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2664) ?
	       wdata32__h27246[29] :
	       _dfoo58 ;
  assign _dfoo1260 =
	     (source_id__h46689 == 10'd16 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1627) ?
	       wdata32__h27246[12] :
	       _dfoo1192 ;
  assign _dfoo1261 =
	     source_id__h46689 == 10'd15 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1627 ||
	     source_id__h48185 == 10'd15 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1688 ||
	     _dfoo1125 ;
  assign _dfoo1262 =
	     (source_id__h46689 == 10'd15 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1627) ?
	       wdata32__h27246[12] :
	       _dfoo1194 ;
  assign _dfoo1263 =
	     source_id__h46689 == 10'd14 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1627 ||
	     source_id__h48185 == 10'd14 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1688 ||
	     _dfoo1127 ;
  assign _dfoo1264 =
	     (source_id__h46689 == 10'd14 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1627) ?
	       wdata32__h27246[12] :
	       _dfoo1196 ;
  assign _dfoo1265 =
	     source_id__h46689 == 10'd13 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1627 ||
	     source_id__h48185 == 10'd13 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1688 ||
	     _dfoo1129 ;
  assign _dfoo1266 =
	     (source_id__h46689 == 10'd13 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1627) ?
	       wdata32__h27246[12] :
	       _dfoo1198 ;
  assign _dfoo1267 =
	     source_id__h46689 == 10'd12 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1627 ||
	     source_id__h48185 == 10'd12 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1688 ||
	     _dfoo1131 ;
  assign _dfoo1268 =
	     (source_id__h46689 == 10'd12 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1627) ?
	       wdata32__h27246[12] :
	       _dfoo1200 ;
  assign _dfoo1269 =
	     source_id__h46689 == 10'd11 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1627 ||
	     source_id__h48185 == 10'd11 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1688 ||
	     _dfoo1133 ;
  assign _dfoo1270 =
	     (source_id__h46689 == 10'd11 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1627) ?
	       wdata32__h27246[12] :
	       _dfoo1202 ;
  assign _dfoo1271 =
	     source_id__h46689 == 10'd10 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1627 ||
	     source_id__h48185 == 10'd10 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1688 ||
	     _dfoo1135 ;
  assign _dfoo1272 =
	     (source_id__h46689 == 10'd10 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1627) ?
	       wdata32__h27246[12] :
	       _dfoo1204 ;
  assign _dfoo1273 =
	     source_id__h46689 == 10'd9 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1627 ||
	     source_id__h48185 == 10'd9 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1688 ||
	     _dfoo1137 ;
  assign _dfoo1274 =
	     (source_id__h46689 == 10'd9 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1627) ?
	       wdata32__h27246[12] :
	       _dfoo1206 ;
  assign _dfoo1275 =
	     source_id__h46689 == 10'd8 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1627 ||
	     source_id__h48185 == 10'd8 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1688 ||
	     _dfoo1139 ;
  assign _dfoo1276 =
	     (source_id__h46689 == 10'd8 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1627) ?
	       wdata32__h27246[12] :
	       _dfoo1208 ;
  assign _dfoo1277 =
	     source_id__h46689 == 10'd7 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1627 ||
	     source_id__h48185 == 10'd7 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1688 ||
	     _dfoo1141 ;
  assign _dfoo1278 =
	     (source_id__h46689 == 10'd7 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1627) ?
	       wdata32__h27246[12] :
	       _dfoo1210 ;
  assign _dfoo1279 =
	     source_id__h46689 == 10'd6 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1627 ||
	     source_id__h48185 == 10'd6 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1688 ||
	     _dfoo1143 ;
  assign _dfoo128 =
	     (source_id__h72121 == 10'd4 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2664) ?
	       wdata32__h27246[29] :
	       _dfoo60 ;
  assign _dfoo1280 =
	     (source_id__h46689 == 10'd6 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1627) ?
	       wdata32__h27246[12] :
	       _dfoo1212 ;
  assign _dfoo1281 =
	     source_id__h46689 == 10'd5 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1627 ||
	     source_id__h48185 == 10'd5 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1688 ||
	     _dfoo1145 ;
  assign _dfoo1282 =
	     (source_id__h46689 == 10'd5 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1627) ?
	       wdata32__h27246[12] :
	       _dfoo1214 ;
  assign _dfoo1283 =
	     source_id__h46689 == 10'd4 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1627 ||
	     source_id__h48185 == 10'd4 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1688 ||
	     _dfoo1147 ;
  assign _dfoo1284 =
	     (source_id__h46689 == 10'd4 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1627) ?
	       wdata32__h27246[12] :
	       _dfoo1216 ;
  assign _dfoo1285 =
	     source_id__h46689 == 10'd3 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1627 ||
	     source_id__h48185 == 10'd3 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1688 ||
	     _dfoo1149 ;
  assign _dfoo1286 =
	     (source_id__h46689 == 10'd3 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1627) ?
	       wdata32__h27246[12] :
	       _dfoo1218 ;
  assign _dfoo1287 =
	     source_id__h46689 == 10'd2 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1627 ||
	     source_id__h48185 == 10'd2 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1688 ||
	     _dfoo1151 ;
  assign _dfoo1288 =
	     (source_id__h46689 == 10'd2 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1627) ?
	       wdata32__h27246[12] :
	       _dfoo1220 ;
  assign _dfoo1289 =
	     source_id__h46689 == 10'd1 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1627 ||
	     source_id__h48185 == 10'd1 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1688 ||
	     _dfoo1153 ;
  assign _dfoo1290 =
	     (source_id__h46689 == 10'd1 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1627) ?
	       wdata32__h27246[12] :
	       _dfoo1222 ;
  assign _dfoo1291 =
	     source_id__h46689 == 10'd0 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1627 ||
	     source_id__h48185 == 10'd0 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1688 ||
	     _dfoo1155 ;
  assign _dfoo1292 =
	     (source_id__h46689 == 10'd0 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1627) ?
	       wdata32__h27246[12] :
	       _dfoo1224 ;
  assign _dfoo1294 =
	     (source_id__h45193 == 10'd16 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1566) ?
	       wdata32__h27246[11] :
	       _dfoo1226 ;
  assign _dfoo1296 =
	     (source_id__h45193 == 10'd15 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1566) ?
	       wdata32__h27246[11] :
	       _dfoo1228 ;
  assign _dfoo1298 =
	     (source_id__h45193 == 10'd14 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1566) ?
	       wdata32__h27246[11] :
	       _dfoo1230 ;
  assign _dfoo13 =
	     source_id__h73617 == 10'd10 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2725 ||
	     source_id__h75113 == 10'd10 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2786 ;
  assign _dfoo130 =
	     (source_id__h72121 == 10'd3 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2664) ?
	       wdata32__h27246[29] :
	       _dfoo62 ;
  assign _dfoo1300 =
	     (source_id__h45193 == 10'd13 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1566) ?
	       wdata32__h27246[11] :
	       _dfoo1232 ;
  assign _dfoo1302 =
	     (source_id__h45193 == 10'd12 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1566) ?
	       wdata32__h27246[11] :
	       _dfoo1234 ;
  assign _dfoo1304 =
	     (source_id__h45193 == 10'd11 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1566) ?
	       wdata32__h27246[11] :
	       _dfoo1236 ;
  assign _dfoo1306 =
	     (source_id__h45193 == 10'd10 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1566) ?
	       wdata32__h27246[11] :
	       _dfoo1238 ;
  assign _dfoo1308 =
	     (source_id__h45193 == 10'd9 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1566) ?
	       wdata32__h27246[11] :
	       _dfoo1240 ;
  assign _dfoo1310 =
	     (source_id__h45193 == 10'd8 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1566) ?
	       wdata32__h27246[11] :
	       _dfoo1242 ;
  assign _dfoo1312 =
	     (source_id__h45193 == 10'd7 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1566) ?
	       wdata32__h27246[11] :
	       _dfoo1244 ;
  assign _dfoo1314 =
	     (source_id__h45193 == 10'd6 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1566) ?
	       wdata32__h27246[11] :
	       _dfoo1246 ;
  assign _dfoo1316 =
	     (source_id__h45193 == 10'd5 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1566) ?
	       wdata32__h27246[11] :
	       _dfoo1248 ;
  assign _dfoo1318 =
	     (source_id__h45193 == 10'd4 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1566) ?
	       wdata32__h27246[11] :
	       _dfoo1250 ;
  assign _dfoo132 =
	     (source_id__h72121 == 10'd2 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2664) ?
	       wdata32__h27246[29] :
	       _dfoo64 ;
  assign _dfoo1320 =
	     (source_id__h45193 == 10'd3 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1566) ?
	       wdata32__h27246[11] :
	       _dfoo1252 ;
  assign _dfoo1322 =
	     (source_id__h45193 == 10'd2 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1566) ?
	       wdata32__h27246[11] :
	       _dfoo1254 ;
  assign _dfoo1324 =
	     (source_id__h45193 == 10'd1 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1566) ?
	       wdata32__h27246[11] :
	       _dfoo1256 ;
  assign _dfoo1326 =
	     (source_id__h45193 == 10'd0 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1566) ?
	       wdata32__h27246[11] :
	       _dfoo1258 ;
  assign _dfoo1328 =
	     (source_id__h45193 == 10'd16 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1566) ?
	       wdata32__h27246[11] :
	       _dfoo1260 ;
  assign _dfoo1330 =
	     (source_id__h45193 == 10'd15 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1566) ?
	       wdata32__h27246[11] :
	       _dfoo1262 ;
  assign _dfoo1332 =
	     (source_id__h45193 == 10'd14 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1566) ?
	       wdata32__h27246[11] :
	       _dfoo1264 ;
  assign _dfoo1334 =
	     (source_id__h45193 == 10'd13 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1566) ?
	       wdata32__h27246[11] :
	       _dfoo1266 ;
  assign _dfoo1336 =
	     (source_id__h45193 == 10'd12 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1566) ?
	       wdata32__h27246[11] :
	       _dfoo1268 ;
  assign _dfoo1338 =
	     (source_id__h45193 == 10'd11 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1566) ?
	       wdata32__h27246[11] :
	       _dfoo1270 ;
  assign _dfoo134 =
	     (source_id__h72121 == 10'd1 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2664) ?
	       wdata32__h27246[29] :
	       _dfoo66 ;
  assign _dfoo1340 =
	     (source_id__h45193 == 10'd10 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1566) ?
	       wdata32__h27246[11] :
	       _dfoo1272 ;
  assign _dfoo1342 =
	     (source_id__h45193 == 10'd9 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1566) ?
	       wdata32__h27246[11] :
	       _dfoo1274 ;
  assign _dfoo1344 =
	     (source_id__h45193 == 10'd8 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1566) ?
	       wdata32__h27246[11] :
	       _dfoo1276 ;
  assign _dfoo1346 =
	     (source_id__h45193 == 10'd7 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1566) ?
	       wdata32__h27246[11] :
	       _dfoo1278 ;
  assign _dfoo1348 =
	     (source_id__h45193 == 10'd6 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1566) ?
	       wdata32__h27246[11] :
	       _dfoo1280 ;
  assign _dfoo1350 =
	     (source_id__h45193 == 10'd5 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1566) ?
	       wdata32__h27246[11] :
	       _dfoo1282 ;
  assign _dfoo1352 =
	     (source_id__h45193 == 10'd4 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1566) ?
	       wdata32__h27246[11] :
	       _dfoo1284 ;
  assign _dfoo1354 =
	     (source_id__h45193 == 10'd3 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1566) ?
	       wdata32__h27246[11] :
	       _dfoo1286 ;
  assign _dfoo1356 =
	     (source_id__h45193 == 10'd2 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1566) ?
	       wdata32__h27246[11] :
	       _dfoo1288 ;
  assign _dfoo1358 =
	     (source_id__h45193 == 10'd1 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1566) ?
	       wdata32__h27246[11] :
	       _dfoo1290 ;
  assign _dfoo136 =
	     (source_id__h72121 == 10'd0 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2664) ?
	       wdata32__h27246[29] :
	       _dfoo68 ;
  assign _dfoo1360 =
	     (source_id__h45193 == 10'd0 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1566) ?
	       wdata32__h27246[11] :
	       _dfoo1292 ;
  assign _dfoo1361 =
	     source_id__h43697 == 10'd16 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1505 ||
	     source_id__h45193 == 10'd16 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1566 ||
	     _dfoo1225 ;
  assign _dfoo1362 =
	     (source_id__h43697 == 10'd16 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1505) ?
	       wdata32__h27246[10] :
	       _dfoo1294 ;
  assign _dfoo1363 =
	     source_id__h43697 == 10'd15 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1505 ||
	     source_id__h45193 == 10'd15 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1566 ||
	     _dfoo1227 ;
  assign _dfoo1364 =
	     (source_id__h43697 == 10'd15 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1505) ?
	       wdata32__h27246[10] :
	       _dfoo1296 ;
  assign _dfoo1365 =
	     source_id__h43697 == 10'd14 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1505 ||
	     source_id__h45193 == 10'd14 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1566 ||
	     _dfoo1229 ;
  assign _dfoo1366 =
	     (source_id__h43697 == 10'd14 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1505) ?
	       wdata32__h27246[10] :
	       _dfoo1298 ;
  assign _dfoo1367 =
	     source_id__h43697 == 10'd13 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1505 ||
	     source_id__h45193 == 10'd13 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1566 ||
	     _dfoo1231 ;
  assign _dfoo1368 =
	     (source_id__h43697 == 10'd13 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1505) ?
	       wdata32__h27246[10] :
	       _dfoo1300 ;
  assign _dfoo1369 =
	     source_id__h43697 == 10'd12 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1505 ||
	     source_id__h45193 == 10'd12 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1566 ||
	     _dfoo1233 ;
  assign _dfoo137 =
	     source_id__h70625 == 10'd16 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2603 ||
	     source_id__h72121 == 10'd16 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2664 ||
	     _dfoo1 ;
  assign _dfoo1370 =
	     (source_id__h43697 == 10'd12 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1505) ?
	       wdata32__h27246[10] :
	       _dfoo1302 ;
  assign _dfoo1371 =
	     source_id__h43697 == 10'd11 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1505 ||
	     source_id__h45193 == 10'd11 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1566 ||
	     _dfoo1235 ;
  assign _dfoo1372 =
	     (source_id__h43697 == 10'd11 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1505) ?
	       wdata32__h27246[10] :
	       _dfoo1304 ;
  assign _dfoo1373 =
	     source_id__h43697 == 10'd10 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1505 ||
	     source_id__h45193 == 10'd10 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1566 ||
	     _dfoo1237 ;
  assign _dfoo1374 =
	     (source_id__h43697 == 10'd10 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1505) ?
	       wdata32__h27246[10] :
	       _dfoo1306 ;
  assign _dfoo1375 =
	     source_id__h43697 == 10'd9 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1505 ||
	     source_id__h45193 == 10'd9 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1566 ||
	     _dfoo1239 ;
  assign _dfoo1376 =
	     (source_id__h43697 == 10'd9 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1505) ?
	       wdata32__h27246[10] :
	       _dfoo1308 ;
  assign _dfoo1377 =
	     source_id__h43697 == 10'd8 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1505 ||
	     source_id__h45193 == 10'd8 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1566 ||
	     _dfoo1241 ;
  assign _dfoo1378 =
	     (source_id__h43697 == 10'd8 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1505) ?
	       wdata32__h27246[10] :
	       _dfoo1310 ;
  assign _dfoo1379 =
	     source_id__h43697 == 10'd7 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1505 ||
	     source_id__h45193 == 10'd7 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1566 ||
	     _dfoo1243 ;
  assign _dfoo138 =
	     (source_id__h70625 == 10'd16 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2603) ?
	       wdata32__h27246[28] :
	       _dfoo70 ;
  assign _dfoo1380 =
	     (source_id__h43697 == 10'd7 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1505) ?
	       wdata32__h27246[10] :
	       _dfoo1312 ;
  assign _dfoo1381 =
	     source_id__h43697 == 10'd6 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1505 ||
	     source_id__h45193 == 10'd6 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1566 ||
	     _dfoo1245 ;
  assign _dfoo1382 =
	     (source_id__h43697 == 10'd6 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1505) ?
	       wdata32__h27246[10] :
	       _dfoo1314 ;
  assign _dfoo1383 =
	     source_id__h43697 == 10'd5 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1505 ||
	     source_id__h45193 == 10'd5 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1566 ||
	     _dfoo1247 ;
  assign _dfoo1384 =
	     (source_id__h43697 == 10'd5 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1505) ?
	       wdata32__h27246[10] :
	       _dfoo1316 ;
  assign _dfoo1385 =
	     source_id__h43697 == 10'd4 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1505 ||
	     source_id__h45193 == 10'd4 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1566 ||
	     _dfoo1249 ;
  assign _dfoo1386 =
	     (source_id__h43697 == 10'd4 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1505) ?
	       wdata32__h27246[10] :
	       _dfoo1318 ;
  assign _dfoo1387 =
	     source_id__h43697 == 10'd3 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1505 ||
	     source_id__h45193 == 10'd3 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1566 ||
	     _dfoo1251 ;
  assign _dfoo1388 =
	     (source_id__h43697 == 10'd3 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1505) ?
	       wdata32__h27246[10] :
	       _dfoo1320 ;
  assign _dfoo1389 =
	     source_id__h43697 == 10'd2 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1505 ||
	     source_id__h45193 == 10'd2 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1566 ||
	     _dfoo1253 ;
  assign _dfoo139 =
	     source_id__h70625 == 10'd15 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2603 ||
	     source_id__h72121 == 10'd15 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2664 ||
	     _dfoo3 ;
  assign _dfoo1390 =
	     (source_id__h43697 == 10'd2 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1505) ?
	       wdata32__h27246[10] :
	       _dfoo1322 ;
  assign _dfoo1391 =
	     source_id__h43697 == 10'd1 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1505 ||
	     source_id__h45193 == 10'd1 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1566 ||
	     _dfoo1255 ;
  assign _dfoo1392 =
	     (source_id__h43697 == 10'd1 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1505) ?
	       wdata32__h27246[10] :
	       _dfoo1324 ;
  assign _dfoo1393 =
	     source_id__h43697 == 10'd0 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1505 ||
	     source_id__h45193 == 10'd0 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1566 ||
	     _dfoo1257 ;
  assign _dfoo1394 =
	     (source_id__h43697 == 10'd0 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1505) ?
	       wdata32__h27246[10] :
	       _dfoo1326 ;
  assign _dfoo1395 =
	     source_id__h43697 == 10'd16 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1505 ||
	     source_id__h45193 == 10'd16 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1566 ||
	     _dfoo1259 ;
  assign _dfoo1396 =
	     (source_id__h43697 == 10'd16 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1505) ?
	       wdata32__h27246[10] :
	       _dfoo1328 ;
  assign _dfoo1397 =
	     source_id__h43697 == 10'd15 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1505 ||
	     source_id__h45193 == 10'd15 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1566 ||
	     _dfoo1261 ;
  assign _dfoo1398 =
	     (source_id__h43697 == 10'd15 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1505) ?
	       wdata32__h27246[10] :
	       _dfoo1330 ;
  assign _dfoo1399 =
	     source_id__h43697 == 10'd14 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1505 ||
	     source_id__h45193 == 10'd14 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1566 ||
	     _dfoo1263 ;
  assign _dfoo14 =
	     (source_id__h73617 == 10'd10 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2725) ?
	       wdata32__h27246[30] :
	       wdata32__h27246[31] ;
  assign _dfoo140 =
	     (source_id__h70625 == 10'd15 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2603) ?
	       wdata32__h27246[28] :
	       _dfoo72 ;
  assign _dfoo1400 =
	     (source_id__h43697 == 10'd14 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1505) ?
	       wdata32__h27246[10] :
	       _dfoo1332 ;
  assign _dfoo1401 =
	     source_id__h43697 == 10'd13 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1505 ||
	     source_id__h45193 == 10'd13 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1566 ||
	     _dfoo1265 ;
  assign _dfoo1402 =
	     (source_id__h43697 == 10'd13 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1505) ?
	       wdata32__h27246[10] :
	       _dfoo1334 ;
  assign _dfoo1403 =
	     source_id__h43697 == 10'd12 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1505 ||
	     source_id__h45193 == 10'd12 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1566 ||
	     _dfoo1267 ;
  assign _dfoo1404 =
	     (source_id__h43697 == 10'd12 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1505) ?
	       wdata32__h27246[10] :
	       _dfoo1336 ;
  assign _dfoo1405 =
	     source_id__h43697 == 10'd11 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1505 ||
	     source_id__h45193 == 10'd11 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1566 ||
	     _dfoo1269 ;
  assign _dfoo1406 =
	     (source_id__h43697 == 10'd11 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1505) ?
	       wdata32__h27246[10] :
	       _dfoo1338 ;
  assign _dfoo1407 =
	     source_id__h43697 == 10'd10 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1505 ||
	     source_id__h45193 == 10'd10 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1566 ||
	     _dfoo1271 ;
  assign _dfoo1408 =
	     (source_id__h43697 == 10'd10 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1505) ?
	       wdata32__h27246[10] :
	       _dfoo1340 ;
  assign _dfoo1409 =
	     source_id__h43697 == 10'd9 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1505 ||
	     source_id__h45193 == 10'd9 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1566 ||
	     _dfoo1273 ;
  assign _dfoo141 =
	     source_id__h70625 == 10'd14 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2603 ||
	     source_id__h72121 == 10'd14 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2664 ||
	     _dfoo5 ;
  assign _dfoo1410 =
	     (source_id__h43697 == 10'd9 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1505) ?
	       wdata32__h27246[10] :
	       _dfoo1342 ;
  assign _dfoo1411 =
	     source_id__h43697 == 10'd8 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1505 ||
	     source_id__h45193 == 10'd8 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1566 ||
	     _dfoo1275 ;
  assign _dfoo1412 =
	     (source_id__h43697 == 10'd8 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1505) ?
	       wdata32__h27246[10] :
	       _dfoo1344 ;
  assign _dfoo1413 =
	     source_id__h43697 == 10'd7 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1505 ||
	     source_id__h45193 == 10'd7 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1566 ||
	     _dfoo1277 ;
  assign _dfoo1414 =
	     (source_id__h43697 == 10'd7 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1505) ?
	       wdata32__h27246[10] :
	       _dfoo1346 ;
  assign _dfoo1415 =
	     source_id__h43697 == 10'd6 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1505 ||
	     source_id__h45193 == 10'd6 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1566 ||
	     _dfoo1279 ;
  assign _dfoo1416 =
	     (source_id__h43697 == 10'd6 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1505) ?
	       wdata32__h27246[10] :
	       _dfoo1348 ;
  assign _dfoo1417 =
	     source_id__h43697 == 10'd5 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1505 ||
	     source_id__h45193 == 10'd5 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1566 ||
	     _dfoo1281 ;
  assign _dfoo1418 =
	     (source_id__h43697 == 10'd5 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1505) ?
	       wdata32__h27246[10] :
	       _dfoo1350 ;
  assign _dfoo1419 =
	     source_id__h43697 == 10'd4 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1505 ||
	     source_id__h45193 == 10'd4 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1566 ||
	     _dfoo1283 ;
  assign _dfoo142 =
	     (source_id__h70625 == 10'd14 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2603) ?
	       wdata32__h27246[28] :
	       _dfoo74 ;
  assign _dfoo1420 =
	     (source_id__h43697 == 10'd4 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1505) ?
	       wdata32__h27246[10] :
	       _dfoo1352 ;
  assign _dfoo1421 =
	     source_id__h43697 == 10'd3 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1505 ||
	     source_id__h45193 == 10'd3 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1566 ||
	     _dfoo1285 ;
  assign _dfoo1422 =
	     (source_id__h43697 == 10'd3 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1505) ?
	       wdata32__h27246[10] :
	       _dfoo1354 ;
  assign _dfoo1423 =
	     source_id__h43697 == 10'd2 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1505 ||
	     source_id__h45193 == 10'd2 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1566 ||
	     _dfoo1287 ;
  assign _dfoo1424 =
	     (source_id__h43697 == 10'd2 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1505) ?
	       wdata32__h27246[10] :
	       _dfoo1356 ;
  assign _dfoo1425 =
	     source_id__h43697 == 10'd1 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1505 ||
	     source_id__h45193 == 10'd1 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1566 ||
	     _dfoo1289 ;
  assign _dfoo1426 =
	     (source_id__h43697 == 10'd1 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1505) ?
	       wdata32__h27246[10] :
	       _dfoo1358 ;
  assign _dfoo1427 =
	     source_id__h43697 == 10'd0 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1505 ||
	     source_id__h45193 == 10'd0 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1566 ||
	     _dfoo1291 ;
  assign _dfoo1428 =
	     (source_id__h43697 == 10'd0 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1505) ?
	       wdata32__h27246[10] :
	       _dfoo1360 ;
  assign _dfoo143 =
	     source_id__h70625 == 10'd13 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2603 ||
	     source_id__h72121 == 10'd13 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2664 ||
	     _dfoo7 ;
  assign _dfoo1430 =
	     (source_id__h42201 == 10'd16 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1444) ?
	       wdata32__h27246[9] :
	       _dfoo1362 ;
  assign _dfoo1432 =
	     (source_id__h42201 == 10'd15 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1444) ?
	       wdata32__h27246[9] :
	       _dfoo1364 ;
  assign _dfoo1434 =
	     (source_id__h42201 == 10'd14 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1444) ?
	       wdata32__h27246[9] :
	       _dfoo1366 ;
  assign _dfoo1436 =
	     (source_id__h42201 == 10'd13 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1444) ?
	       wdata32__h27246[9] :
	       _dfoo1368 ;
  assign _dfoo1438 =
	     (source_id__h42201 == 10'd12 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1444) ?
	       wdata32__h27246[9] :
	       _dfoo1370 ;
  assign _dfoo144 =
	     (source_id__h70625 == 10'd13 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2603) ?
	       wdata32__h27246[28] :
	       _dfoo76 ;
  assign _dfoo1440 =
	     (source_id__h42201 == 10'd11 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1444) ?
	       wdata32__h27246[9] :
	       _dfoo1372 ;
  assign _dfoo1442 =
	     (source_id__h42201 == 10'd10 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1444) ?
	       wdata32__h27246[9] :
	       _dfoo1374 ;
  assign _dfoo1444 =
	     (source_id__h42201 == 10'd9 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1444) ?
	       wdata32__h27246[9] :
	       _dfoo1376 ;
  assign _dfoo1446 =
	     (source_id__h42201 == 10'd8 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1444) ?
	       wdata32__h27246[9] :
	       _dfoo1378 ;
  assign _dfoo1448 =
	     (source_id__h42201 == 10'd7 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1444) ?
	       wdata32__h27246[9] :
	       _dfoo1380 ;
  assign _dfoo145 =
	     source_id__h70625 == 10'd12 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2603 ||
	     source_id__h72121 == 10'd12 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2664 ||
	     _dfoo9 ;
  assign _dfoo1450 =
	     (source_id__h42201 == 10'd6 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1444) ?
	       wdata32__h27246[9] :
	       _dfoo1382 ;
  assign _dfoo1452 =
	     (source_id__h42201 == 10'd5 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1444) ?
	       wdata32__h27246[9] :
	       _dfoo1384 ;
  assign _dfoo1454 =
	     (source_id__h42201 == 10'd4 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1444) ?
	       wdata32__h27246[9] :
	       _dfoo1386 ;
  assign _dfoo1456 =
	     (source_id__h42201 == 10'd3 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1444) ?
	       wdata32__h27246[9] :
	       _dfoo1388 ;
  assign _dfoo1458 =
	     (source_id__h42201 == 10'd2 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1444) ?
	       wdata32__h27246[9] :
	       _dfoo1390 ;
  assign _dfoo146 =
	     (source_id__h70625 == 10'd12 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2603) ?
	       wdata32__h27246[28] :
	       _dfoo78 ;
  assign _dfoo1460 =
	     (source_id__h42201 == 10'd1 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1444) ?
	       wdata32__h27246[9] :
	       _dfoo1392 ;
  assign _dfoo1462 =
	     (source_id__h42201 == 10'd0 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1444) ?
	       wdata32__h27246[9] :
	       _dfoo1394 ;
  assign _dfoo1464 =
	     (source_id__h42201 == 10'd16 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1444) ?
	       wdata32__h27246[9] :
	       _dfoo1396 ;
  assign _dfoo1466 =
	     (source_id__h42201 == 10'd15 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1444) ?
	       wdata32__h27246[9] :
	       _dfoo1398 ;
  assign _dfoo1468 =
	     (source_id__h42201 == 10'd14 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1444) ?
	       wdata32__h27246[9] :
	       _dfoo1400 ;
  assign _dfoo147 =
	     source_id__h70625 == 10'd11 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2603 ||
	     source_id__h72121 == 10'd11 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2664 ||
	     _dfoo11 ;
  assign _dfoo1470 =
	     (source_id__h42201 == 10'd13 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1444) ?
	       wdata32__h27246[9] :
	       _dfoo1402 ;
  assign _dfoo1472 =
	     (source_id__h42201 == 10'd12 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1444) ?
	       wdata32__h27246[9] :
	       _dfoo1404 ;
  assign _dfoo1474 =
	     (source_id__h42201 == 10'd11 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1444) ?
	       wdata32__h27246[9] :
	       _dfoo1406 ;
  assign _dfoo1476 =
	     (source_id__h42201 == 10'd10 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1444) ?
	       wdata32__h27246[9] :
	       _dfoo1408 ;
  assign _dfoo1478 =
	     (source_id__h42201 == 10'd9 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1444) ?
	       wdata32__h27246[9] :
	       _dfoo1410 ;
  assign _dfoo148 =
	     (source_id__h70625 == 10'd11 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2603) ?
	       wdata32__h27246[28] :
	       _dfoo80 ;
  assign _dfoo1480 =
	     (source_id__h42201 == 10'd8 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1444) ?
	       wdata32__h27246[9] :
	       _dfoo1412 ;
  assign _dfoo1482 =
	     (source_id__h42201 == 10'd7 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1444) ?
	       wdata32__h27246[9] :
	       _dfoo1414 ;
  assign _dfoo1484 =
	     (source_id__h42201 == 10'd6 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1444) ?
	       wdata32__h27246[9] :
	       _dfoo1416 ;
  assign _dfoo1486 =
	     (source_id__h42201 == 10'd5 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1444) ?
	       wdata32__h27246[9] :
	       _dfoo1418 ;
  assign _dfoo1488 =
	     (source_id__h42201 == 10'd4 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1444) ?
	       wdata32__h27246[9] :
	       _dfoo1420 ;
  assign _dfoo149 =
	     source_id__h70625 == 10'd10 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2603 ||
	     source_id__h72121 == 10'd10 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2664 ||
	     _dfoo13 ;
  assign _dfoo1490 =
	     (source_id__h42201 == 10'd3 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1444) ?
	       wdata32__h27246[9] :
	       _dfoo1422 ;
  assign _dfoo1492 =
	     (source_id__h42201 == 10'd2 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1444) ?
	       wdata32__h27246[9] :
	       _dfoo1424 ;
  assign _dfoo1494 =
	     (source_id__h42201 == 10'd1 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1444) ?
	       wdata32__h27246[9] :
	       _dfoo1426 ;
  assign _dfoo1496 =
	     (source_id__h42201 == 10'd0 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1444) ?
	       wdata32__h27246[9] :
	       _dfoo1428 ;
  assign _dfoo1497 =
	     source_id__h40705 == 10'd16 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1383 ||
	     source_id__h42201 == 10'd16 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1444 ||
	     _dfoo1361 ;
  assign _dfoo1498 =
	     (source_id__h40705 == 10'd16 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1383) ?
	       wdata32__h27246[8] :
	       _dfoo1430 ;
  assign _dfoo1499 =
	     source_id__h40705 == 10'd15 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1383 ||
	     source_id__h42201 == 10'd15 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1444 ||
	     _dfoo1363 ;
  assign _dfoo15 =
	     source_id__h73617 == 10'd9 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2725 ||
	     source_id__h75113 == 10'd9 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2786 ;
  assign _dfoo150 =
	     (source_id__h70625 == 10'd10 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2603) ?
	       wdata32__h27246[28] :
	       _dfoo82 ;
  assign _dfoo1500 =
	     (source_id__h40705 == 10'd15 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1383) ?
	       wdata32__h27246[8] :
	       _dfoo1432 ;
  assign _dfoo1501 =
	     source_id__h40705 == 10'd14 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1383 ||
	     source_id__h42201 == 10'd14 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1444 ||
	     _dfoo1365 ;
  assign _dfoo1502 =
	     (source_id__h40705 == 10'd14 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1383) ?
	       wdata32__h27246[8] :
	       _dfoo1434 ;
  assign _dfoo1503 =
	     source_id__h40705 == 10'd13 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1383 ||
	     source_id__h42201 == 10'd13 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1444 ||
	     _dfoo1367 ;
  assign _dfoo1504 =
	     (source_id__h40705 == 10'd13 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1383) ?
	       wdata32__h27246[8] :
	       _dfoo1436 ;
  assign _dfoo1505 =
	     source_id__h40705 == 10'd12 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1383 ||
	     source_id__h42201 == 10'd12 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1444 ||
	     _dfoo1369 ;
  assign _dfoo1506 =
	     (source_id__h40705 == 10'd12 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1383) ?
	       wdata32__h27246[8] :
	       _dfoo1438 ;
  assign _dfoo1507 =
	     source_id__h40705 == 10'd11 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1383 ||
	     source_id__h42201 == 10'd11 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1444 ||
	     _dfoo1371 ;
  assign _dfoo1508 =
	     (source_id__h40705 == 10'd11 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1383) ?
	       wdata32__h27246[8] :
	       _dfoo1440 ;
  assign _dfoo1509 =
	     source_id__h40705 == 10'd10 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1383 ||
	     source_id__h42201 == 10'd10 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1444 ||
	     _dfoo1373 ;
  assign _dfoo151 =
	     source_id__h70625 == 10'd9 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2603 ||
	     source_id__h72121 == 10'd9 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2664 ||
	     _dfoo15 ;
  assign _dfoo1510 =
	     (source_id__h40705 == 10'd10 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1383) ?
	       wdata32__h27246[8] :
	       _dfoo1442 ;
  assign _dfoo1511 =
	     source_id__h40705 == 10'd9 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1383 ||
	     source_id__h42201 == 10'd9 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1444 ||
	     _dfoo1375 ;
  assign _dfoo1512 =
	     (source_id__h40705 == 10'd9 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1383) ?
	       wdata32__h27246[8] :
	       _dfoo1444 ;
  assign _dfoo1513 =
	     source_id__h40705 == 10'd8 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1383 ||
	     source_id__h42201 == 10'd8 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1444 ||
	     _dfoo1377 ;
  assign _dfoo1514 =
	     (source_id__h40705 == 10'd8 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1383) ?
	       wdata32__h27246[8] :
	       _dfoo1446 ;
  assign _dfoo1515 =
	     source_id__h40705 == 10'd7 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1383 ||
	     source_id__h42201 == 10'd7 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1444 ||
	     _dfoo1379 ;
  assign _dfoo1516 =
	     (source_id__h40705 == 10'd7 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1383) ?
	       wdata32__h27246[8] :
	       _dfoo1448 ;
  assign _dfoo1517 =
	     source_id__h40705 == 10'd6 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1383 ||
	     source_id__h42201 == 10'd6 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1444 ||
	     _dfoo1381 ;
  assign _dfoo1518 =
	     (source_id__h40705 == 10'd6 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1383) ?
	       wdata32__h27246[8] :
	       _dfoo1450 ;
  assign _dfoo1519 =
	     source_id__h40705 == 10'd5 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1383 ||
	     source_id__h42201 == 10'd5 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1444 ||
	     _dfoo1383 ;
  assign _dfoo152 =
	     (source_id__h70625 == 10'd9 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2603) ?
	       wdata32__h27246[28] :
	       _dfoo84 ;
  assign _dfoo1520 =
	     (source_id__h40705 == 10'd5 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1383) ?
	       wdata32__h27246[8] :
	       _dfoo1452 ;
  assign _dfoo1521 =
	     source_id__h40705 == 10'd4 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1383 ||
	     source_id__h42201 == 10'd4 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1444 ||
	     _dfoo1385 ;
  assign _dfoo1522 =
	     (source_id__h40705 == 10'd4 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1383) ?
	       wdata32__h27246[8] :
	       _dfoo1454 ;
  assign _dfoo1523 =
	     source_id__h40705 == 10'd3 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1383 ||
	     source_id__h42201 == 10'd3 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1444 ||
	     _dfoo1387 ;
  assign _dfoo1524 =
	     (source_id__h40705 == 10'd3 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1383) ?
	       wdata32__h27246[8] :
	       _dfoo1456 ;
  assign _dfoo1525 =
	     source_id__h40705 == 10'd2 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1383 ||
	     source_id__h42201 == 10'd2 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1444 ||
	     _dfoo1389 ;
  assign _dfoo1526 =
	     (source_id__h40705 == 10'd2 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1383) ?
	       wdata32__h27246[8] :
	       _dfoo1458 ;
  assign _dfoo1527 =
	     source_id__h40705 == 10'd1 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1383 ||
	     source_id__h42201 == 10'd1 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1444 ||
	     _dfoo1391 ;
  assign _dfoo1528 =
	     (source_id__h40705 == 10'd1 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1383) ?
	       wdata32__h27246[8] :
	       _dfoo1460 ;
  assign _dfoo1529 =
	     source_id__h40705 == 10'd0 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1383 ||
	     source_id__h42201 == 10'd0 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1444 ||
	     _dfoo1393 ;
  assign _dfoo153 =
	     source_id__h70625 == 10'd8 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2603 ||
	     source_id__h72121 == 10'd8 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2664 ||
	     _dfoo17 ;
  assign _dfoo1530 =
	     (source_id__h40705 == 10'd0 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1383) ?
	       wdata32__h27246[8] :
	       _dfoo1462 ;
  assign _dfoo1531 =
	     source_id__h40705 == 10'd16 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1383 ||
	     source_id__h42201 == 10'd16 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1444 ||
	     _dfoo1395 ;
  assign _dfoo1532 =
	     (source_id__h40705 == 10'd16 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1383) ?
	       wdata32__h27246[8] :
	       _dfoo1464 ;
  assign _dfoo1533 =
	     source_id__h40705 == 10'd15 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1383 ||
	     source_id__h42201 == 10'd15 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1444 ||
	     _dfoo1397 ;
  assign _dfoo1534 =
	     (source_id__h40705 == 10'd15 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1383) ?
	       wdata32__h27246[8] :
	       _dfoo1466 ;
  assign _dfoo1535 =
	     source_id__h40705 == 10'd14 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1383 ||
	     source_id__h42201 == 10'd14 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1444 ||
	     _dfoo1399 ;
  assign _dfoo1536 =
	     (source_id__h40705 == 10'd14 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1383) ?
	       wdata32__h27246[8] :
	       _dfoo1468 ;
  assign _dfoo1537 =
	     source_id__h40705 == 10'd13 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1383 ||
	     source_id__h42201 == 10'd13 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1444 ||
	     _dfoo1401 ;
  assign _dfoo1538 =
	     (source_id__h40705 == 10'd13 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1383) ?
	       wdata32__h27246[8] :
	       _dfoo1470 ;
  assign _dfoo1539 =
	     source_id__h40705 == 10'd12 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1383 ||
	     source_id__h42201 == 10'd12 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1444 ||
	     _dfoo1403 ;
  assign _dfoo154 =
	     (source_id__h70625 == 10'd8 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2603) ?
	       wdata32__h27246[28] :
	       _dfoo86 ;
  assign _dfoo1540 =
	     (source_id__h40705 == 10'd12 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1383) ?
	       wdata32__h27246[8] :
	       _dfoo1472 ;
  assign _dfoo1541 =
	     source_id__h40705 == 10'd11 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1383 ||
	     source_id__h42201 == 10'd11 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1444 ||
	     _dfoo1405 ;
  assign _dfoo1542 =
	     (source_id__h40705 == 10'd11 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1383) ?
	       wdata32__h27246[8] :
	       _dfoo1474 ;
  assign _dfoo1543 =
	     source_id__h40705 == 10'd10 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1383 ||
	     source_id__h42201 == 10'd10 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1444 ||
	     _dfoo1407 ;
  assign _dfoo1544 =
	     (source_id__h40705 == 10'd10 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1383) ?
	       wdata32__h27246[8] :
	       _dfoo1476 ;
  assign _dfoo1545 =
	     source_id__h40705 == 10'd9 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1383 ||
	     source_id__h42201 == 10'd9 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1444 ||
	     _dfoo1409 ;
  assign _dfoo1546 =
	     (source_id__h40705 == 10'd9 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1383) ?
	       wdata32__h27246[8] :
	       _dfoo1478 ;
  assign _dfoo1547 =
	     source_id__h40705 == 10'd8 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1383 ||
	     source_id__h42201 == 10'd8 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1444 ||
	     _dfoo1411 ;
  assign _dfoo1548 =
	     (source_id__h40705 == 10'd8 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1383) ?
	       wdata32__h27246[8] :
	       _dfoo1480 ;
  assign _dfoo1549 =
	     source_id__h40705 == 10'd7 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1383 ||
	     source_id__h42201 == 10'd7 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1444 ||
	     _dfoo1413 ;
  assign _dfoo155 =
	     source_id__h70625 == 10'd7 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2603 ||
	     source_id__h72121 == 10'd7 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2664 ||
	     _dfoo19 ;
  assign _dfoo1550 =
	     (source_id__h40705 == 10'd7 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1383) ?
	       wdata32__h27246[8] :
	       _dfoo1482 ;
  assign _dfoo1551 =
	     source_id__h40705 == 10'd6 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1383 ||
	     source_id__h42201 == 10'd6 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1444 ||
	     _dfoo1415 ;
  assign _dfoo1552 =
	     (source_id__h40705 == 10'd6 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1383) ?
	       wdata32__h27246[8] :
	       _dfoo1484 ;
  assign _dfoo1553 =
	     source_id__h40705 == 10'd5 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1383 ||
	     source_id__h42201 == 10'd5 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1444 ||
	     _dfoo1417 ;
  assign _dfoo1554 =
	     (source_id__h40705 == 10'd5 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1383) ?
	       wdata32__h27246[8] :
	       _dfoo1486 ;
  assign _dfoo1555 =
	     source_id__h40705 == 10'd4 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1383 ||
	     source_id__h42201 == 10'd4 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1444 ||
	     _dfoo1419 ;
  assign _dfoo1556 =
	     (source_id__h40705 == 10'd4 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1383) ?
	       wdata32__h27246[8] :
	       _dfoo1488 ;
  assign _dfoo1557 =
	     source_id__h40705 == 10'd3 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1383 ||
	     source_id__h42201 == 10'd3 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1444 ||
	     _dfoo1421 ;
  assign _dfoo1558 =
	     (source_id__h40705 == 10'd3 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1383) ?
	       wdata32__h27246[8] :
	       _dfoo1490 ;
  assign _dfoo1559 =
	     source_id__h40705 == 10'd2 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1383 ||
	     source_id__h42201 == 10'd2 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1444 ||
	     _dfoo1423 ;
  assign _dfoo156 =
	     (source_id__h70625 == 10'd7 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2603) ?
	       wdata32__h27246[28] :
	       _dfoo88 ;
  assign _dfoo1560 =
	     (source_id__h40705 == 10'd2 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1383) ?
	       wdata32__h27246[8] :
	       _dfoo1492 ;
  assign _dfoo1561 =
	     source_id__h40705 == 10'd1 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1383 ||
	     source_id__h42201 == 10'd1 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1444 ||
	     _dfoo1425 ;
  assign _dfoo1562 =
	     (source_id__h40705 == 10'd1 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1383) ?
	       wdata32__h27246[8] :
	       _dfoo1494 ;
  assign _dfoo1563 =
	     source_id__h40705 == 10'd0 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1383 ||
	     source_id__h42201 == 10'd0 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1444 ||
	     _dfoo1427 ;
  assign _dfoo1564 =
	     (source_id__h40705 == 10'd0 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1383) ?
	       wdata32__h27246[8] :
	       _dfoo1496 ;
  assign _dfoo1566 =
	     (source_id__h39209 == 10'd16 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1322) ?
	       wdata32__h27246[7] :
	       _dfoo1498 ;
  assign _dfoo1568 =
	     (source_id__h39209 == 10'd15 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1322) ?
	       wdata32__h27246[7] :
	       _dfoo1500 ;
  assign _dfoo157 =
	     source_id__h70625 == 10'd6 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2603 ||
	     source_id__h72121 == 10'd6 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2664 ||
	     _dfoo21 ;
  assign _dfoo1570 =
	     (source_id__h39209 == 10'd14 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1322) ?
	       wdata32__h27246[7] :
	       _dfoo1502 ;
  assign _dfoo1572 =
	     (source_id__h39209 == 10'd13 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1322) ?
	       wdata32__h27246[7] :
	       _dfoo1504 ;
  assign _dfoo1574 =
	     (source_id__h39209 == 10'd12 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1322) ?
	       wdata32__h27246[7] :
	       _dfoo1506 ;
  assign _dfoo1576 =
	     (source_id__h39209 == 10'd11 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1322) ?
	       wdata32__h27246[7] :
	       _dfoo1508 ;
  assign _dfoo1578 =
	     (source_id__h39209 == 10'd10 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1322) ?
	       wdata32__h27246[7] :
	       _dfoo1510 ;
  assign _dfoo158 =
	     (source_id__h70625 == 10'd6 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2603) ?
	       wdata32__h27246[28] :
	       _dfoo90 ;
  assign _dfoo1580 =
	     (source_id__h39209 == 10'd9 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1322) ?
	       wdata32__h27246[7] :
	       _dfoo1512 ;
  assign _dfoo1582 =
	     (source_id__h39209 == 10'd8 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1322) ?
	       wdata32__h27246[7] :
	       _dfoo1514 ;
  assign _dfoo1584 =
	     (source_id__h39209 == 10'd7 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1322) ?
	       wdata32__h27246[7] :
	       _dfoo1516 ;
  assign _dfoo1586 =
	     (source_id__h39209 == 10'd6 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1322) ?
	       wdata32__h27246[7] :
	       _dfoo1518 ;
  assign _dfoo1588 =
	     (source_id__h39209 == 10'd5 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1322) ?
	       wdata32__h27246[7] :
	       _dfoo1520 ;
  assign _dfoo159 =
	     source_id__h70625 == 10'd5 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2603 ||
	     source_id__h72121 == 10'd5 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2664 ||
	     _dfoo23 ;
  assign _dfoo1590 =
	     (source_id__h39209 == 10'd4 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1322) ?
	       wdata32__h27246[7] :
	       _dfoo1522 ;
  assign _dfoo1592 =
	     (source_id__h39209 == 10'd3 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1322) ?
	       wdata32__h27246[7] :
	       _dfoo1524 ;
  assign _dfoo1594 =
	     (source_id__h39209 == 10'd2 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1322) ?
	       wdata32__h27246[7] :
	       _dfoo1526 ;
  assign _dfoo1596 =
	     (source_id__h39209 == 10'd1 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1322) ?
	       wdata32__h27246[7] :
	       _dfoo1528 ;
  assign _dfoo1598 =
	     (source_id__h39209 == 10'd0 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1322) ?
	       wdata32__h27246[7] :
	       _dfoo1530 ;
  assign _dfoo16 =
	     (source_id__h73617 == 10'd9 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2725) ?
	       wdata32__h27246[30] :
	       wdata32__h27246[31] ;
  assign _dfoo160 =
	     (source_id__h70625 == 10'd5 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2603) ?
	       wdata32__h27246[28] :
	       _dfoo92 ;
  assign _dfoo1600 =
	     (source_id__h39209 == 10'd16 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1322) ?
	       wdata32__h27246[7] :
	       _dfoo1532 ;
  assign _dfoo1602 =
	     (source_id__h39209 == 10'd15 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1322) ?
	       wdata32__h27246[7] :
	       _dfoo1534 ;
  assign _dfoo1604 =
	     (source_id__h39209 == 10'd14 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1322) ?
	       wdata32__h27246[7] :
	       _dfoo1536 ;
  assign _dfoo1606 =
	     (source_id__h39209 == 10'd13 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1322) ?
	       wdata32__h27246[7] :
	       _dfoo1538 ;
  assign _dfoo1608 =
	     (source_id__h39209 == 10'd12 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1322) ?
	       wdata32__h27246[7] :
	       _dfoo1540 ;
  assign _dfoo161 =
	     source_id__h70625 == 10'd4 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2603 ||
	     source_id__h72121 == 10'd4 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2664 ||
	     _dfoo25 ;
  assign _dfoo1610 =
	     (source_id__h39209 == 10'd11 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1322) ?
	       wdata32__h27246[7] :
	       _dfoo1542 ;
  assign _dfoo1612 =
	     (source_id__h39209 == 10'd10 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1322) ?
	       wdata32__h27246[7] :
	       _dfoo1544 ;
  assign _dfoo1614 =
	     (source_id__h39209 == 10'd9 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1322) ?
	       wdata32__h27246[7] :
	       _dfoo1546 ;
  assign _dfoo1616 =
	     (source_id__h39209 == 10'd8 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1322) ?
	       wdata32__h27246[7] :
	       _dfoo1548 ;
  assign _dfoo1618 =
	     (source_id__h39209 == 10'd7 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1322) ?
	       wdata32__h27246[7] :
	       _dfoo1550 ;
  assign _dfoo162 =
	     (source_id__h70625 == 10'd4 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2603) ?
	       wdata32__h27246[28] :
	       _dfoo94 ;
  assign _dfoo1620 =
	     (source_id__h39209 == 10'd6 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1322) ?
	       wdata32__h27246[7] :
	       _dfoo1552 ;
  assign _dfoo1622 =
	     (source_id__h39209 == 10'd5 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1322) ?
	       wdata32__h27246[7] :
	       _dfoo1554 ;
  assign _dfoo1624 =
	     (source_id__h39209 == 10'd4 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1322) ?
	       wdata32__h27246[7] :
	       _dfoo1556 ;
  assign _dfoo1626 =
	     (source_id__h39209 == 10'd3 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1322) ?
	       wdata32__h27246[7] :
	       _dfoo1558 ;
  assign _dfoo1628 =
	     (source_id__h39209 == 10'd2 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1322) ?
	       wdata32__h27246[7] :
	       _dfoo1560 ;
  assign _dfoo163 =
	     source_id__h70625 == 10'd3 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2603 ||
	     source_id__h72121 == 10'd3 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2664 ||
	     _dfoo27 ;
  assign _dfoo1630 =
	     (source_id__h39209 == 10'd1 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1322) ?
	       wdata32__h27246[7] :
	       _dfoo1562 ;
  assign _dfoo1632 =
	     (source_id__h39209 == 10'd0 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1322) ?
	       wdata32__h27246[7] :
	       _dfoo1564 ;
  assign _dfoo1633 =
	     source_id__h37713 == 10'd16 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1261 ||
	     source_id__h39209 == 10'd16 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1322 ||
	     _dfoo1497 ;
  assign _dfoo1634 =
	     (source_id__h37713 == 10'd16 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1261) ?
	       wdata32__h27246[6] :
	       _dfoo1566 ;
  assign _dfoo1635 =
	     source_id__h37713 == 10'd15 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1261 ||
	     source_id__h39209 == 10'd15 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1322 ||
	     _dfoo1499 ;
  assign _dfoo1636 =
	     (source_id__h37713 == 10'd15 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1261) ?
	       wdata32__h27246[6] :
	       _dfoo1568 ;
  assign _dfoo1637 =
	     source_id__h37713 == 10'd14 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1261 ||
	     source_id__h39209 == 10'd14 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1322 ||
	     _dfoo1501 ;
  assign _dfoo1638 =
	     (source_id__h37713 == 10'd14 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1261) ?
	       wdata32__h27246[6] :
	       _dfoo1570 ;
  assign _dfoo1639 =
	     source_id__h37713 == 10'd13 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1261 ||
	     source_id__h39209 == 10'd13 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1322 ||
	     _dfoo1503 ;
  assign _dfoo164 =
	     (source_id__h70625 == 10'd3 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2603) ?
	       wdata32__h27246[28] :
	       _dfoo96 ;
  assign _dfoo1640 =
	     (source_id__h37713 == 10'd13 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1261) ?
	       wdata32__h27246[6] :
	       _dfoo1572 ;
  assign _dfoo1641 =
	     source_id__h37713 == 10'd12 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1261 ||
	     source_id__h39209 == 10'd12 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1322 ||
	     _dfoo1505 ;
  assign _dfoo1642 =
	     (source_id__h37713 == 10'd12 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1261) ?
	       wdata32__h27246[6] :
	       _dfoo1574 ;
  assign _dfoo1643 =
	     source_id__h37713 == 10'd11 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1261 ||
	     source_id__h39209 == 10'd11 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1322 ||
	     _dfoo1507 ;
  assign _dfoo1644 =
	     (source_id__h37713 == 10'd11 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1261) ?
	       wdata32__h27246[6] :
	       _dfoo1576 ;
  assign _dfoo1645 =
	     source_id__h37713 == 10'd10 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1261 ||
	     source_id__h39209 == 10'd10 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1322 ||
	     _dfoo1509 ;
  assign _dfoo1646 =
	     (source_id__h37713 == 10'd10 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1261) ?
	       wdata32__h27246[6] :
	       _dfoo1578 ;
  assign _dfoo1647 =
	     source_id__h37713 == 10'd9 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1261 ||
	     source_id__h39209 == 10'd9 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1322 ||
	     _dfoo1511 ;
  assign _dfoo1648 =
	     (source_id__h37713 == 10'd9 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1261) ?
	       wdata32__h27246[6] :
	       _dfoo1580 ;
  assign _dfoo1649 =
	     source_id__h37713 == 10'd8 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1261 ||
	     source_id__h39209 == 10'd8 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1322 ||
	     _dfoo1513 ;
  assign _dfoo165 =
	     source_id__h70625 == 10'd2 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2603 ||
	     source_id__h72121 == 10'd2 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2664 ||
	     _dfoo29 ;
  assign _dfoo1650 =
	     (source_id__h37713 == 10'd8 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1261) ?
	       wdata32__h27246[6] :
	       _dfoo1582 ;
  assign _dfoo1651 =
	     source_id__h37713 == 10'd7 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1261 ||
	     source_id__h39209 == 10'd7 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1322 ||
	     _dfoo1515 ;
  assign _dfoo1652 =
	     (source_id__h37713 == 10'd7 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1261) ?
	       wdata32__h27246[6] :
	       _dfoo1584 ;
  assign _dfoo1653 =
	     source_id__h37713 == 10'd6 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1261 ||
	     source_id__h39209 == 10'd6 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1322 ||
	     _dfoo1517 ;
  assign _dfoo1654 =
	     (source_id__h37713 == 10'd6 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1261) ?
	       wdata32__h27246[6] :
	       _dfoo1586 ;
  assign _dfoo1655 =
	     source_id__h37713 == 10'd5 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1261 ||
	     source_id__h39209 == 10'd5 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1322 ||
	     _dfoo1519 ;
  assign _dfoo1656 =
	     (source_id__h37713 == 10'd5 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1261) ?
	       wdata32__h27246[6] :
	       _dfoo1588 ;
  assign _dfoo1657 =
	     source_id__h37713 == 10'd4 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1261 ||
	     source_id__h39209 == 10'd4 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1322 ||
	     _dfoo1521 ;
  assign _dfoo1658 =
	     (source_id__h37713 == 10'd4 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1261) ?
	       wdata32__h27246[6] :
	       _dfoo1590 ;
  assign _dfoo1659 =
	     source_id__h37713 == 10'd3 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1261 ||
	     source_id__h39209 == 10'd3 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1322 ||
	     _dfoo1523 ;
  assign _dfoo166 =
	     (source_id__h70625 == 10'd2 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2603) ?
	       wdata32__h27246[28] :
	       _dfoo98 ;
  assign _dfoo1660 =
	     (source_id__h37713 == 10'd3 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1261) ?
	       wdata32__h27246[6] :
	       _dfoo1592 ;
  assign _dfoo1661 =
	     source_id__h37713 == 10'd2 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1261 ||
	     source_id__h39209 == 10'd2 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1322 ||
	     _dfoo1525 ;
  assign _dfoo1662 =
	     (source_id__h37713 == 10'd2 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1261) ?
	       wdata32__h27246[6] :
	       _dfoo1594 ;
  assign _dfoo1663 =
	     source_id__h37713 == 10'd1 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1261 ||
	     source_id__h39209 == 10'd1 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1322 ||
	     _dfoo1527 ;
  assign _dfoo1664 =
	     (source_id__h37713 == 10'd1 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1261) ?
	       wdata32__h27246[6] :
	       _dfoo1596 ;
  assign _dfoo1665 =
	     source_id__h37713 == 10'd0 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1261 ||
	     source_id__h39209 == 10'd0 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1322 ||
	     _dfoo1529 ;
  assign _dfoo1666 =
	     (source_id__h37713 == 10'd0 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1261) ?
	       wdata32__h27246[6] :
	       _dfoo1598 ;
  assign _dfoo1667 =
	     source_id__h37713 == 10'd16 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1261 ||
	     source_id__h39209 == 10'd16 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1322 ||
	     _dfoo1531 ;
  assign _dfoo1668 =
	     (source_id__h37713 == 10'd16 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1261) ?
	       wdata32__h27246[6] :
	       _dfoo1600 ;
  assign _dfoo1669 =
	     source_id__h37713 == 10'd15 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1261 ||
	     source_id__h39209 == 10'd15 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1322 ||
	     _dfoo1533 ;
  assign _dfoo167 =
	     source_id__h70625 == 10'd1 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2603 ||
	     source_id__h72121 == 10'd1 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2664 ||
	     _dfoo31 ;
  assign _dfoo1670 =
	     (source_id__h37713 == 10'd15 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1261) ?
	       wdata32__h27246[6] :
	       _dfoo1602 ;
  assign _dfoo1671 =
	     source_id__h37713 == 10'd14 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1261 ||
	     source_id__h39209 == 10'd14 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1322 ||
	     _dfoo1535 ;
  assign _dfoo1672 =
	     (source_id__h37713 == 10'd14 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1261) ?
	       wdata32__h27246[6] :
	       _dfoo1604 ;
  assign _dfoo1673 =
	     source_id__h37713 == 10'd13 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1261 ||
	     source_id__h39209 == 10'd13 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1322 ||
	     _dfoo1537 ;
  assign _dfoo1674 =
	     (source_id__h37713 == 10'd13 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1261) ?
	       wdata32__h27246[6] :
	       _dfoo1606 ;
  assign _dfoo1675 =
	     source_id__h37713 == 10'd12 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1261 ||
	     source_id__h39209 == 10'd12 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1322 ||
	     _dfoo1539 ;
  assign _dfoo1676 =
	     (source_id__h37713 == 10'd12 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1261) ?
	       wdata32__h27246[6] :
	       _dfoo1608 ;
  assign _dfoo1677 =
	     source_id__h37713 == 10'd11 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1261 ||
	     source_id__h39209 == 10'd11 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1322 ||
	     _dfoo1541 ;
  assign _dfoo1678 =
	     (source_id__h37713 == 10'd11 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1261) ?
	       wdata32__h27246[6] :
	       _dfoo1610 ;
  assign _dfoo1679 =
	     source_id__h37713 == 10'd10 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1261 ||
	     source_id__h39209 == 10'd10 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1322 ||
	     _dfoo1543 ;
  assign _dfoo168 =
	     (source_id__h70625 == 10'd1 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2603) ?
	       wdata32__h27246[28] :
	       _dfoo100 ;
  assign _dfoo1680 =
	     (source_id__h37713 == 10'd10 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1261) ?
	       wdata32__h27246[6] :
	       _dfoo1612 ;
  assign _dfoo1681 =
	     source_id__h37713 == 10'd9 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1261 ||
	     source_id__h39209 == 10'd9 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1322 ||
	     _dfoo1545 ;
  assign _dfoo1682 =
	     (source_id__h37713 == 10'd9 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1261) ?
	       wdata32__h27246[6] :
	       _dfoo1614 ;
  assign _dfoo1683 =
	     source_id__h37713 == 10'd8 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1261 ||
	     source_id__h39209 == 10'd8 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1322 ||
	     _dfoo1547 ;
  assign _dfoo1684 =
	     (source_id__h37713 == 10'd8 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1261) ?
	       wdata32__h27246[6] :
	       _dfoo1616 ;
  assign _dfoo1685 =
	     source_id__h37713 == 10'd7 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1261 ||
	     source_id__h39209 == 10'd7 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1322 ||
	     _dfoo1549 ;
  assign _dfoo1686 =
	     (source_id__h37713 == 10'd7 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1261) ?
	       wdata32__h27246[6] :
	       _dfoo1618 ;
  assign _dfoo1687 =
	     source_id__h37713 == 10'd6 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1261 ||
	     source_id__h39209 == 10'd6 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1322 ||
	     _dfoo1551 ;
  assign _dfoo1688 =
	     (source_id__h37713 == 10'd6 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1261) ?
	       wdata32__h27246[6] :
	       _dfoo1620 ;
  assign _dfoo1689 =
	     source_id__h37713 == 10'd5 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1261 ||
	     source_id__h39209 == 10'd5 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1322 ||
	     _dfoo1553 ;
  assign _dfoo169 =
	     source_id__h70625 == 10'd0 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2603 ||
	     source_id__h72121 == 10'd0 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2664 ||
	     _dfoo33 ;
  assign _dfoo1690 =
	     (source_id__h37713 == 10'd5 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1261) ?
	       wdata32__h27246[6] :
	       _dfoo1622 ;
  assign _dfoo1691 =
	     source_id__h37713 == 10'd4 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1261 ||
	     source_id__h39209 == 10'd4 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1322 ||
	     _dfoo1555 ;
  assign _dfoo1692 =
	     (source_id__h37713 == 10'd4 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1261) ?
	       wdata32__h27246[6] :
	       _dfoo1624 ;
  assign _dfoo1693 =
	     source_id__h37713 == 10'd3 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1261 ||
	     source_id__h39209 == 10'd3 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1322 ||
	     _dfoo1557 ;
  assign _dfoo1694 =
	     (source_id__h37713 == 10'd3 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1261) ?
	       wdata32__h27246[6] :
	       _dfoo1626 ;
  assign _dfoo1695 =
	     source_id__h37713 == 10'd2 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1261 ||
	     source_id__h39209 == 10'd2 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1322 ||
	     _dfoo1559 ;
  assign _dfoo1696 =
	     (source_id__h37713 == 10'd2 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1261) ?
	       wdata32__h27246[6] :
	       _dfoo1628 ;
  assign _dfoo1697 =
	     source_id__h37713 == 10'd1 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1261 ||
	     source_id__h39209 == 10'd1 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1322 ||
	     _dfoo1561 ;
  assign _dfoo1698 =
	     (source_id__h37713 == 10'd1 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1261) ?
	       wdata32__h27246[6] :
	       _dfoo1630 ;
  assign _dfoo1699 =
	     source_id__h37713 == 10'd0 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1261 ||
	     source_id__h39209 == 10'd0 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1322 ||
	     _dfoo1563 ;
  assign _dfoo17 =
	     source_id__h73617 == 10'd8 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2725 ||
	     source_id__h75113 == 10'd8 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2786 ;
  assign _dfoo170 =
	     (source_id__h70625 == 10'd0 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2603) ?
	       wdata32__h27246[28] :
	       _dfoo102 ;
  assign _dfoo1700 =
	     (source_id__h37713 == 10'd0 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1261) ?
	       wdata32__h27246[6] :
	       _dfoo1632 ;
  assign _dfoo1702 =
	     (source_id__h36217 == 10'd16 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1200) ?
	       wdata32__h27246[5] :
	       _dfoo1634 ;
  assign _dfoo1704 =
	     (source_id__h36217 == 10'd15 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1200) ?
	       wdata32__h27246[5] :
	       _dfoo1636 ;
  assign _dfoo1706 =
	     (source_id__h36217 == 10'd14 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1200) ?
	       wdata32__h27246[5] :
	       _dfoo1638 ;
  assign _dfoo1708 =
	     (source_id__h36217 == 10'd13 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1200) ?
	       wdata32__h27246[5] :
	       _dfoo1640 ;
  assign _dfoo171 =
	     source_id__h70625 == 10'd16 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2603 ||
	     source_id__h72121 == 10'd16 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2664 ||
	     _dfoo35 ;
  assign _dfoo1710 =
	     (source_id__h36217 == 10'd12 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1200) ?
	       wdata32__h27246[5] :
	       _dfoo1642 ;
  assign _dfoo1712 =
	     (source_id__h36217 == 10'd11 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1200) ?
	       wdata32__h27246[5] :
	       _dfoo1644 ;
  assign _dfoo1714 =
	     (source_id__h36217 == 10'd10 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1200) ?
	       wdata32__h27246[5] :
	       _dfoo1646 ;
  assign _dfoo1716 =
	     (source_id__h36217 == 10'd9 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1200) ?
	       wdata32__h27246[5] :
	       _dfoo1648 ;
  assign _dfoo1718 =
	     (source_id__h36217 == 10'd8 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1200) ?
	       wdata32__h27246[5] :
	       _dfoo1650 ;
  assign _dfoo172 =
	     (source_id__h70625 == 10'd16 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2603) ?
	       wdata32__h27246[28] :
	       _dfoo104 ;
  assign _dfoo1720 =
	     (source_id__h36217 == 10'd7 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1200) ?
	       wdata32__h27246[5] :
	       _dfoo1652 ;
  assign _dfoo1722 =
	     (source_id__h36217 == 10'd6 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1200) ?
	       wdata32__h27246[5] :
	       _dfoo1654 ;
  assign _dfoo1724 =
	     (source_id__h36217 == 10'd5 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1200) ?
	       wdata32__h27246[5] :
	       _dfoo1656 ;
  assign _dfoo1726 =
	     (source_id__h36217 == 10'd4 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1200) ?
	       wdata32__h27246[5] :
	       _dfoo1658 ;
  assign _dfoo1728 =
	     (source_id__h36217 == 10'd3 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1200) ?
	       wdata32__h27246[5] :
	       _dfoo1660 ;
  assign _dfoo173 =
	     source_id__h70625 == 10'd15 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2603 ||
	     source_id__h72121 == 10'd15 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2664 ||
	     _dfoo37 ;
  assign _dfoo1730 =
	     (source_id__h36217 == 10'd2 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1200) ?
	       wdata32__h27246[5] :
	       _dfoo1662 ;
  assign _dfoo1732 =
	     (source_id__h36217 == 10'd1 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1200) ?
	       wdata32__h27246[5] :
	       _dfoo1664 ;
  assign _dfoo1734 =
	     (source_id__h36217 == 10'd0 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1200) ?
	       wdata32__h27246[5] :
	       _dfoo1666 ;
  assign _dfoo1736 =
	     (source_id__h36217 == 10'd16 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1200) ?
	       wdata32__h27246[5] :
	       _dfoo1668 ;
  assign _dfoo1738 =
	     (source_id__h36217 == 10'd15 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1200) ?
	       wdata32__h27246[5] :
	       _dfoo1670 ;
  assign _dfoo174 =
	     (source_id__h70625 == 10'd15 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2603) ?
	       wdata32__h27246[28] :
	       _dfoo106 ;
  assign _dfoo1740 =
	     (source_id__h36217 == 10'd14 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1200) ?
	       wdata32__h27246[5] :
	       _dfoo1672 ;
  assign _dfoo1742 =
	     (source_id__h36217 == 10'd13 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1200) ?
	       wdata32__h27246[5] :
	       _dfoo1674 ;
  assign _dfoo1744 =
	     (source_id__h36217 == 10'd12 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1200) ?
	       wdata32__h27246[5] :
	       _dfoo1676 ;
  assign _dfoo1746 =
	     (source_id__h36217 == 10'd11 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1200) ?
	       wdata32__h27246[5] :
	       _dfoo1678 ;
  assign _dfoo1748 =
	     (source_id__h36217 == 10'd10 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1200) ?
	       wdata32__h27246[5] :
	       _dfoo1680 ;
  assign _dfoo175 =
	     source_id__h70625 == 10'd14 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2603 ||
	     source_id__h72121 == 10'd14 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2664 ||
	     _dfoo39 ;
  assign _dfoo1750 =
	     (source_id__h36217 == 10'd9 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1200) ?
	       wdata32__h27246[5] :
	       _dfoo1682 ;
  assign _dfoo1752 =
	     (source_id__h36217 == 10'd8 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1200) ?
	       wdata32__h27246[5] :
	       _dfoo1684 ;
  assign _dfoo1754 =
	     (source_id__h36217 == 10'd7 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1200) ?
	       wdata32__h27246[5] :
	       _dfoo1686 ;
  assign _dfoo1756 =
	     (source_id__h36217 == 10'd6 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1200) ?
	       wdata32__h27246[5] :
	       _dfoo1688 ;
  assign _dfoo1758 =
	     (source_id__h36217 == 10'd5 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1200) ?
	       wdata32__h27246[5] :
	       _dfoo1690 ;
  assign _dfoo176 =
	     (source_id__h70625 == 10'd14 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2603) ?
	       wdata32__h27246[28] :
	       _dfoo108 ;
  assign _dfoo1760 =
	     (source_id__h36217 == 10'd4 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1200) ?
	       wdata32__h27246[5] :
	       _dfoo1692 ;
  assign _dfoo1762 =
	     (source_id__h36217 == 10'd3 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1200) ?
	       wdata32__h27246[5] :
	       _dfoo1694 ;
  assign _dfoo1764 =
	     (source_id__h36217 == 10'd2 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1200) ?
	       wdata32__h27246[5] :
	       _dfoo1696 ;
  assign _dfoo1766 =
	     (source_id__h36217 == 10'd1 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1200) ?
	       wdata32__h27246[5] :
	       _dfoo1698 ;
  assign _dfoo1768 =
	     (source_id__h36217 == 10'd0 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1200) ?
	       wdata32__h27246[5] :
	       _dfoo1700 ;
  assign _dfoo1769 =
	     source_id__h34721 == 10'd16 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1139 ||
	     source_id__h36217 == 10'd16 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1200 ||
	     _dfoo1633 ;
  assign _dfoo177 =
	     source_id__h70625 == 10'd13 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2603 ||
	     source_id__h72121 == 10'd13 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2664 ||
	     _dfoo41 ;
  assign _dfoo1770 =
	     (source_id__h34721 == 10'd16 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1139) ?
	       wdata32__h27246[4] :
	       _dfoo1702 ;
  assign _dfoo1771 =
	     source_id__h34721 == 10'd15 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1139 ||
	     source_id__h36217 == 10'd15 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1200 ||
	     _dfoo1635 ;
  assign _dfoo1772 =
	     (source_id__h34721 == 10'd15 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1139) ?
	       wdata32__h27246[4] :
	       _dfoo1704 ;
  assign _dfoo1773 =
	     source_id__h34721 == 10'd14 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1139 ||
	     source_id__h36217 == 10'd14 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1200 ||
	     _dfoo1637 ;
  assign _dfoo1774 =
	     (source_id__h34721 == 10'd14 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1139) ?
	       wdata32__h27246[4] :
	       _dfoo1706 ;
  assign _dfoo1775 =
	     source_id__h34721 == 10'd13 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1139 ||
	     source_id__h36217 == 10'd13 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1200 ||
	     _dfoo1639 ;
  assign _dfoo1776 =
	     (source_id__h34721 == 10'd13 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1139) ?
	       wdata32__h27246[4] :
	       _dfoo1708 ;
  assign _dfoo1777 =
	     source_id__h34721 == 10'd12 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1139 ||
	     source_id__h36217 == 10'd12 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1200 ||
	     _dfoo1641 ;
  assign _dfoo1778 =
	     (source_id__h34721 == 10'd12 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1139) ?
	       wdata32__h27246[4] :
	       _dfoo1710 ;
  assign _dfoo1779 =
	     source_id__h34721 == 10'd11 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1139 ||
	     source_id__h36217 == 10'd11 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1200 ||
	     _dfoo1643 ;
  assign _dfoo178 =
	     (source_id__h70625 == 10'd13 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2603) ?
	       wdata32__h27246[28] :
	       _dfoo110 ;
  assign _dfoo1780 =
	     (source_id__h34721 == 10'd11 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1139) ?
	       wdata32__h27246[4] :
	       _dfoo1712 ;
  assign _dfoo1781 =
	     source_id__h34721 == 10'd10 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1139 ||
	     source_id__h36217 == 10'd10 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1200 ||
	     _dfoo1645 ;
  assign _dfoo1782 =
	     (source_id__h34721 == 10'd10 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1139) ?
	       wdata32__h27246[4] :
	       _dfoo1714 ;
  assign _dfoo1783 =
	     source_id__h34721 == 10'd9 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1139 ||
	     source_id__h36217 == 10'd9 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1200 ||
	     _dfoo1647 ;
  assign _dfoo1784 =
	     (source_id__h34721 == 10'd9 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1139) ?
	       wdata32__h27246[4] :
	       _dfoo1716 ;
  assign _dfoo1785 =
	     source_id__h34721 == 10'd8 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1139 ||
	     source_id__h36217 == 10'd8 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1200 ||
	     _dfoo1649 ;
  assign _dfoo1786 =
	     (source_id__h34721 == 10'd8 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1139) ?
	       wdata32__h27246[4] :
	       _dfoo1718 ;
  assign _dfoo1787 =
	     source_id__h34721 == 10'd7 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1139 ||
	     source_id__h36217 == 10'd7 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1200 ||
	     _dfoo1651 ;
  assign _dfoo1788 =
	     (source_id__h34721 == 10'd7 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1139) ?
	       wdata32__h27246[4] :
	       _dfoo1720 ;
  assign _dfoo1789 =
	     source_id__h34721 == 10'd6 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1139 ||
	     source_id__h36217 == 10'd6 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1200 ||
	     _dfoo1653 ;
  assign _dfoo179 =
	     source_id__h70625 == 10'd12 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2603 ||
	     source_id__h72121 == 10'd12 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2664 ||
	     _dfoo43 ;
  assign _dfoo1790 =
	     (source_id__h34721 == 10'd6 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1139) ?
	       wdata32__h27246[4] :
	       _dfoo1722 ;
  assign _dfoo1791 =
	     source_id__h34721 == 10'd5 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1139 ||
	     source_id__h36217 == 10'd5 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1200 ||
	     _dfoo1655 ;
  assign _dfoo1792 =
	     (source_id__h34721 == 10'd5 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1139) ?
	       wdata32__h27246[4] :
	       _dfoo1724 ;
  assign _dfoo1793 =
	     source_id__h34721 == 10'd4 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1139 ||
	     source_id__h36217 == 10'd4 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1200 ||
	     _dfoo1657 ;
  assign _dfoo1794 =
	     (source_id__h34721 == 10'd4 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1139) ?
	       wdata32__h27246[4] :
	       _dfoo1726 ;
  assign _dfoo1795 =
	     source_id__h34721 == 10'd3 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1139 ||
	     source_id__h36217 == 10'd3 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1200 ||
	     _dfoo1659 ;
  assign _dfoo1796 =
	     (source_id__h34721 == 10'd3 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1139) ?
	       wdata32__h27246[4] :
	       _dfoo1728 ;
  assign _dfoo1797 =
	     source_id__h34721 == 10'd2 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1139 ||
	     source_id__h36217 == 10'd2 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1200 ||
	     _dfoo1661 ;
  assign _dfoo1798 =
	     (source_id__h34721 == 10'd2 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1139) ?
	       wdata32__h27246[4] :
	       _dfoo1730 ;
  assign _dfoo1799 =
	     source_id__h34721 == 10'd1 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1139 ||
	     source_id__h36217 == 10'd1 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1200 ||
	     _dfoo1663 ;
  assign _dfoo18 =
	     (source_id__h73617 == 10'd8 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2725) ?
	       wdata32__h27246[30] :
	       wdata32__h27246[31] ;
  assign _dfoo180 =
	     (source_id__h70625 == 10'd12 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2603) ?
	       wdata32__h27246[28] :
	       _dfoo112 ;
  assign _dfoo1800 =
	     (source_id__h34721 == 10'd1 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1139) ?
	       wdata32__h27246[4] :
	       _dfoo1732 ;
  assign _dfoo1801 =
	     source_id__h34721 == 10'd0 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1139 ||
	     source_id__h36217 == 10'd0 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1200 ||
	     _dfoo1665 ;
  assign _dfoo1802 =
	     (source_id__h34721 == 10'd0 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1139) ?
	       wdata32__h27246[4] :
	       _dfoo1734 ;
  assign _dfoo1803 =
	     source_id__h34721 == 10'd16 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1139 ||
	     source_id__h36217 == 10'd16 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1200 ||
	     _dfoo1667 ;
  assign _dfoo1804 =
	     (source_id__h34721 == 10'd16 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1139) ?
	       wdata32__h27246[4] :
	       _dfoo1736 ;
  assign _dfoo1805 =
	     source_id__h34721 == 10'd15 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1139 ||
	     source_id__h36217 == 10'd15 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1200 ||
	     _dfoo1669 ;
  assign _dfoo1806 =
	     (source_id__h34721 == 10'd15 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1139) ?
	       wdata32__h27246[4] :
	       _dfoo1738 ;
  assign _dfoo1807 =
	     source_id__h34721 == 10'd14 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1139 ||
	     source_id__h36217 == 10'd14 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1200 ||
	     _dfoo1671 ;
  assign _dfoo1808 =
	     (source_id__h34721 == 10'd14 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1139) ?
	       wdata32__h27246[4] :
	       _dfoo1740 ;
  assign _dfoo1809 =
	     source_id__h34721 == 10'd13 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1139 ||
	     source_id__h36217 == 10'd13 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1200 ||
	     _dfoo1673 ;
  assign _dfoo181 =
	     source_id__h70625 == 10'd11 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2603 ||
	     source_id__h72121 == 10'd11 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2664 ||
	     _dfoo45 ;
  assign _dfoo1810 =
	     (source_id__h34721 == 10'd13 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1139) ?
	       wdata32__h27246[4] :
	       _dfoo1742 ;
  assign _dfoo1811 =
	     source_id__h34721 == 10'd12 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1139 ||
	     source_id__h36217 == 10'd12 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1200 ||
	     _dfoo1675 ;
  assign _dfoo1812 =
	     (source_id__h34721 == 10'd12 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1139) ?
	       wdata32__h27246[4] :
	       _dfoo1744 ;
  assign _dfoo1813 =
	     source_id__h34721 == 10'd11 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1139 ||
	     source_id__h36217 == 10'd11 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1200 ||
	     _dfoo1677 ;
  assign _dfoo1814 =
	     (source_id__h34721 == 10'd11 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1139) ?
	       wdata32__h27246[4] :
	       _dfoo1746 ;
  assign _dfoo1815 =
	     source_id__h34721 == 10'd10 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1139 ||
	     source_id__h36217 == 10'd10 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1200 ||
	     _dfoo1679 ;
  assign _dfoo1816 =
	     (source_id__h34721 == 10'd10 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1139) ?
	       wdata32__h27246[4] :
	       _dfoo1748 ;
  assign _dfoo1817 =
	     source_id__h34721 == 10'd9 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1139 ||
	     source_id__h36217 == 10'd9 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1200 ||
	     _dfoo1681 ;
  assign _dfoo1818 =
	     (source_id__h34721 == 10'd9 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1139) ?
	       wdata32__h27246[4] :
	       _dfoo1750 ;
  assign _dfoo1819 =
	     source_id__h34721 == 10'd8 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1139 ||
	     source_id__h36217 == 10'd8 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1200 ||
	     _dfoo1683 ;
  assign _dfoo182 =
	     (source_id__h70625 == 10'd11 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2603) ?
	       wdata32__h27246[28] :
	       _dfoo114 ;
  assign _dfoo1820 =
	     (source_id__h34721 == 10'd8 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1139) ?
	       wdata32__h27246[4] :
	       _dfoo1752 ;
  assign _dfoo1821 =
	     source_id__h34721 == 10'd7 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1139 ||
	     source_id__h36217 == 10'd7 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1200 ||
	     _dfoo1685 ;
  assign _dfoo1822 =
	     (source_id__h34721 == 10'd7 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1139) ?
	       wdata32__h27246[4] :
	       _dfoo1754 ;
  assign _dfoo1823 =
	     source_id__h34721 == 10'd6 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1139 ||
	     source_id__h36217 == 10'd6 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1200 ||
	     _dfoo1687 ;
  assign _dfoo1824 =
	     (source_id__h34721 == 10'd6 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1139) ?
	       wdata32__h27246[4] :
	       _dfoo1756 ;
  assign _dfoo1825 =
	     source_id__h34721 == 10'd5 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1139 ||
	     source_id__h36217 == 10'd5 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1200 ||
	     _dfoo1689 ;
  assign _dfoo1826 =
	     (source_id__h34721 == 10'd5 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1139) ?
	       wdata32__h27246[4] :
	       _dfoo1758 ;
  assign _dfoo1827 =
	     source_id__h34721 == 10'd4 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1139 ||
	     source_id__h36217 == 10'd4 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1200 ||
	     _dfoo1691 ;
  assign _dfoo1828 =
	     (source_id__h34721 == 10'd4 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1139) ?
	       wdata32__h27246[4] :
	       _dfoo1760 ;
  assign _dfoo1829 =
	     source_id__h34721 == 10'd3 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1139 ||
	     source_id__h36217 == 10'd3 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1200 ||
	     _dfoo1693 ;
  assign _dfoo183 =
	     source_id__h70625 == 10'd10 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2603 ||
	     source_id__h72121 == 10'd10 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2664 ||
	     _dfoo47 ;
  assign _dfoo1830 =
	     (source_id__h34721 == 10'd3 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1139) ?
	       wdata32__h27246[4] :
	       _dfoo1762 ;
  assign _dfoo1831 =
	     source_id__h34721 == 10'd2 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1139 ||
	     source_id__h36217 == 10'd2 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1200 ||
	     _dfoo1695 ;
  assign _dfoo1832 =
	     (source_id__h34721 == 10'd2 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1139) ?
	       wdata32__h27246[4] :
	       _dfoo1764 ;
  assign _dfoo1833 =
	     source_id__h34721 == 10'd1 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1139 ||
	     source_id__h36217 == 10'd1 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1200 ||
	     _dfoo1697 ;
  assign _dfoo1834 =
	     (source_id__h34721 == 10'd1 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1139) ?
	       wdata32__h27246[4] :
	       _dfoo1766 ;
  assign _dfoo1835 =
	     source_id__h34721 == 10'd0 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1139 ||
	     source_id__h36217 == 10'd0 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1200 ||
	     _dfoo1699 ;
  assign _dfoo1836 =
	     (source_id__h34721 == 10'd0 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1139) ?
	       wdata32__h27246[4] :
	       _dfoo1768 ;
  assign _dfoo1838 =
	     (source_id__h33225 == 10'd16 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1078) ?
	       wdata32__h27246[3] :
	       _dfoo1770 ;
  assign _dfoo184 =
	     (source_id__h70625 == 10'd10 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2603) ?
	       wdata32__h27246[28] :
	       _dfoo116 ;
  assign _dfoo1840 =
	     (source_id__h33225 == 10'd15 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1078) ?
	       wdata32__h27246[3] :
	       _dfoo1772 ;
  assign _dfoo1842 =
	     (source_id__h33225 == 10'd14 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1078) ?
	       wdata32__h27246[3] :
	       _dfoo1774 ;
  assign _dfoo1844 =
	     (source_id__h33225 == 10'd13 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1078) ?
	       wdata32__h27246[3] :
	       _dfoo1776 ;
  assign _dfoo1846 =
	     (source_id__h33225 == 10'd12 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1078) ?
	       wdata32__h27246[3] :
	       _dfoo1778 ;
  assign _dfoo1848 =
	     (source_id__h33225 == 10'd11 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1078) ?
	       wdata32__h27246[3] :
	       _dfoo1780 ;
  assign _dfoo185 =
	     source_id__h70625 == 10'd9 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2603 ||
	     source_id__h72121 == 10'd9 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2664 ||
	     _dfoo49 ;
  assign _dfoo1850 =
	     (source_id__h33225 == 10'd10 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1078) ?
	       wdata32__h27246[3] :
	       _dfoo1782 ;
  assign _dfoo1852 =
	     (source_id__h33225 == 10'd9 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1078) ?
	       wdata32__h27246[3] :
	       _dfoo1784 ;
  assign _dfoo1854 =
	     (source_id__h33225 == 10'd8 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1078) ?
	       wdata32__h27246[3] :
	       _dfoo1786 ;
  assign _dfoo1856 =
	     (source_id__h33225 == 10'd7 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1078) ?
	       wdata32__h27246[3] :
	       _dfoo1788 ;
  assign _dfoo1858 =
	     (source_id__h33225 == 10'd6 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1078) ?
	       wdata32__h27246[3] :
	       _dfoo1790 ;
  assign _dfoo186 =
	     (source_id__h70625 == 10'd9 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2603) ?
	       wdata32__h27246[28] :
	       _dfoo118 ;
  assign _dfoo1860 =
	     (source_id__h33225 == 10'd5 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1078) ?
	       wdata32__h27246[3] :
	       _dfoo1792 ;
  assign _dfoo1862 =
	     (source_id__h33225 == 10'd4 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1078) ?
	       wdata32__h27246[3] :
	       _dfoo1794 ;
  assign _dfoo1864 =
	     (source_id__h33225 == 10'd3 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1078) ?
	       wdata32__h27246[3] :
	       _dfoo1796 ;
  assign _dfoo1866 =
	     (source_id__h33225 == 10'd2 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1078) ?
	       wdata32__h27246[3] :
	       _dfoo1798 ;
  assign _dfoo1868 =
	     (source_id__h33225 == 10'd1 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1078) ?
	       wdata32__h27246[3] :
	       _dfoo1800 ;
  assign _dfoo187 =
	     source_id__h70625 == 10'd8 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2603 ||
	     source_id__h72121 == 10'd8 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2664 ||
	     _dfoo51 ;
  assign _dfoo1870 =
	     (source_id__h33225 == 10'd0 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1078) ?
	       wdata32__h27246[3] :
	       _dfoo1802 ;
  assign _dfoo1872 =
	     (source_id__h33225 == 10'd16 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1078) ?
	       wdata32__h27246[3] :
	       _dfoo1804 ;
  assign _dfoo1874 =
	     (source_id__h33225 == 10'd15 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1078) ?
	       wdata32__h27246[3] :
	       _dfoo1806 ;
  assign _dfoo1876 =
	     (source_id__h33225 == 10'd14 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1078) ?
	       wdata32__h27246[3] :
	       _dfoo1808 ;
  assign _dfoo1878 =
	     (source_id__h33225 == 10'd13 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1078) ?
	       wdata32__h27246[3] :
	       _dfoo1810 ;
  assign _dfoo188 =
	     (source_id__h70625 == 10'd8 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2603) ?
	       wdata32__h27246[28] :
	       _dfoo120 ;
  assign _dfoo1880 =
	     (source_id__h33225 == 10'd12 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1078) ?
	       wdata32__h27246[3] :
	       _dfoo1812 ;
  assign _dfoo1882 =
	     (source_id__h33225 == 10'd11 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1078) ?
	       wdata32__h27246[3] :
	       _dfoo1814 ;
  assign _dfoo1884 =
	     (source_id__h33225 == 10'd10 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1078) ?
	       wdata32__h27246[3] :
	       _dfoo1816 ;
  assign _dfoo1886 =
	     (source_id__h33225 == 10'd9 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1078) ?
	       wdata32__h27246[3] :
	       _dfoo1818 ;
  assign _dfoo1888 =
	     (source_id__h33225 == 10'd8 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1078) ?
	       wdata32__h27246[3] :
	       _dfoo1820 ;
  assign _dfoo189 =
	     source_id__h70625 == 10'd7 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2603 ||
	     source_id__h72121 == 10'd7 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2664 ||
	     _dfoo53 ;
  assign _dfoo1890 =
	     (source_id__h33225 == 10'd7 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1078) ?
	       wdata32__h27246[3] :
	       _dfoo1822 ;
  assign _dfoo1892 =
	     (source_id__h33225 == 10'd6 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1078) ?
	       wdata32__h27246[3] :
	       _dfoo1824 ;
  assign _dfoo1894 =
	     (source_id__h33225 == 10'd5 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1078) ?
	       wdata32__h27246[3] :
	       _dfoo1826 ;
  assign _dfoo1896 =
	     (source_id__h33225 == 10'd4 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1078) ?
	       wdata32__h27246[3] :
	       _dfoo1828 ;
  assign _dfoo1898 =
	     (source_id__h33225 == 10'd3 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1078) ?
	       wdata32__h27246[3] :
	       _dfoo1830 ;
  assign _dfoo19 =
	     source_id__h73617 == 10'd7 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2725 ||
	     source_id__h75113 == 10'd7 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2786 ;
  assign _dfoo190 =
	     (source_id__h70625 == 10'd7 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2603) ?
	       wdata32__h27246[28] :
	       _dfoo122 ;
  assign _dfoo1900 =
	     (source_id__h33225 == 10'd2 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1078) ?
	       wdata32__h27246[3] :
	       _dfoo1832 ;
  assign _dfoo1902 =
	     (source_id__h33225 == 10'd1 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1078) ?
	       wdata32__h27246[3] :
	       _dfoo1834 ;
  assign _dfoo1904 =
	     (source_id__h33225 == 10'd0 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1078) ?
	       wdata32__h27246[3] :
	       _dfoo1836 ;
  assign _dfoo1905 =
	     source_id__h31729 == 10'd16 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1017 ||
	     source_id__h33225 == 10'd16 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1078 ||
	     _dfoo1769 ;
  assign _dfoo1906 =
	     (source_id__h31729 == 10'd16 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1017) ?
	       wdata32__h27246[2] :
	       _dfoo1838 ;
  assign _dfoo1907 =
	     source_id__h31729 == 10'd15 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1017 ||
	     source_id__h33225 == 10'd15 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1078 ||
	     _dfoo1771 ;
  assign _dfoo1908 =
	     (source_id__h31729 == 10'd15 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1017) ?
	       wdata32__h27246[2] :
	       _dfoo1840 ;
  assign _dfoo1909 =
	     source_id__h31729 == 10'd14 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1017 ||
	     source_id__h33225 == 10'd14 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1078 ||
	     _dfoo1773 ;
  assign _dfoo191 =
	     source_id__h70625 == 10'd6 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2603 ||
	     source_id__h72121 == 10'd6 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2664 ||
	     _dfoo55 ;
  assign _dfoo1910 =
	     (source_id__h31729 == 10'd14 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1017) ?
	       wdata32__h27246[2] :
	       _dfoo1842 ;
  assign _dfoo1911 =
	     source_id__h31729 == 10'd13 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1017 ||
	     source_id__h33225 == 10'd13 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1078 ||
	     _dfoo1775 ;
  assign _dfoo1912 =
	     (source_id__h31729 == 10'd13 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1017) ?
	       wdata32__h27246[2] :
	       _dfoo1844 ;
  assign _dfoo1913 =
	     source_id__h31729 == 10'd12 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1017 ||
	     source_id__h33225 == 10'd12 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1078 ||
	     _dfoo1777 ;
  assign _dfoo1914 =
	     (source_id__h31729 == 10'd12 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1017) ?
	       wdata32__h27246[2] :
	       _dfoo1846 ;
  assign _dfoo1915 =
	     source_id__h31729 == 10'd11 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1017 ||
	     source_id__h33225 == 10'd11 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1078 ||
	     _dfoo1779 ;
  assign _dfoo1916 =
	     (source_id__h31729 == 10'd11 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1017) ?
	       wdata32__h27246[2] :
	       _dfoo1848 ;
  assign _dfoo1917 =
	     source_id__h31729 == 10'd10 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1017 ||
	     source_id__h33225 == 10'd10 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1078 ||
	     _dfoo1781 ;
  assign _dfoo1918 =
	     (source_id__h31729 == 10'd10 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1017) ?
	       wdata32__h27246[2] :
	       _dfoo1850 ;
  assign _dfoo1919 =
	     source_id__h31729 == 10'd9 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1017 ||
	     source_id__h33225 == 10'd9 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1078 ||
	     _dfoo1783 ;
  assign _dfoo192 =
	     (source_id__h70625 == 10'd6 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2603) ?
	       wdata32__h27246[28] :
	       _dfoo124 ;
  assign _dfoo1920 =
	     (source_id__h31729 == 10'd9 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1017) ?
	       wdata32__h27246[2] :
	       _dfoo1852 ;
  assign _dfoo1921 =
	     source_id__h31729 == 10'd8 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1017 ||
	     source_id__h33225 == 10'd8 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1078 ||
	     _dfoo1785 ;
  assign _dfoo1922 =
	     (source_id__h31729 == 10'd8 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1017) ?
	       wdata32__h27246[2] :
	       _dfoo1854 ;
  assign _dfoo1923 =
	     source_id__h31729 == 10'd7 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1017 ||
	     source_id__h33225 == 10'd7 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1078 ||
	     _dfoo1787 ;
  assign _dfoo1924 =
	     (source_id__h31729 == 10'd7 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1017) ?
	       wdata32__h27246[2] :
	       _dfoo1856 ;
  assign _dfoo1925 =
	     source_id__h31729 == 10'd6 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1017 ||
	     source_id__h33225 == 10'd6 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1078 ||
	     _dfoo1789 ;
  assign _dfoo1926 =
	     (source_id__h31729 == 10'd6 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1017) ?
	       wdata32__h27246[2] :
	       _dfoo1858 ;
  assign _dfoo1927 =
	     source_id__h31729 == 10'd5 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1017 ||
	     source_id__h33225 == 10'd5 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1078 ||
	     _dfoo1791 ;
  assign _dfoo1928 =
	     (source_id__h31729 == 10'd5 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1017) ?
	       wdata32__h27246[2] :
	       _dfoo1860 ;
  assign _dfoo1929 =
	     source_id__h31729 == 10'd4 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1017 ||
	     source_id__h33225 == 10'd4 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1078 ||
	     _dfoo1793 ;
  assign _dfoo193 =
	     source_id__h70625 == 10'd5 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2603 ||
	     source_id__h72121 == 10'd5 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2664 ||
	     _dfoo57 ;
  assign _dfoo1930 =
	     (source_id__h31729 == 10'd4 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1017) ?
	       wdata32__h27246[2] :
	       _dfoo1862 ;
  assign _dfoo1931 =
	     source_id__h31729 == 10'd3 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1017 ||
	     source_id__h33225 == 10'd3 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1078 ||
	     _dfoo1795 ;
  assign _dfoo1932 =
	     (source_id__h31729 == 10'd3 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1017) ?
	       wdata32__h27246[2] :
	       _dfoo1864 ;
  assign _dfoo1933 =
	     source_id__h31729 == 10'd2 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1017 ||
	     source_id__h33225 == 10'd2 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1078 ||
	     _dfoo1797 ;
  assign _dfoo1934 =
	     (source_id__h31729 == 10'd2 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1017) ?
	       wdata32__h27246[2] :
	       _dfoo1866 ;
  assign _dfoo1935 =
	     source_id__h31729 == 10'd1 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1017 ||
	     source_id__h33225 == 10'd1 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1078 ||
	     _dfoo1799 ;
  assign _dfoo1936 =
	     (source_id__h31729 == 10'd1 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1017) ?
	       wdata32__h27246[2] :
	       _dfoo1868 ;
  assign _dfoo1937 =
	     source_id__h31729 == 10'd0 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1017 ||
	     source_id__h33225 == 10'd0 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1078 ||
	     _dfoo1801 ;
  assign _dfoo1938 =
	     (source_id__h31729 == 10'd0 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1017) ?
	       wdata32__h27246[2] :
	       _dfoo1870 ;
  assign _dfoo1939 =
	     source_id__h31729 == 10'd16 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1017 ||
	     source_id__h33225 == 10'd16 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1078 ||
	     _dfoo1803 ;
  assign _dfoo194 =
	     (source_id__h70625 == 10'd5 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2603) ?
	       wdata32__h27246[28] :
	       _dfoo126 ;
  assign _dfoo1940 =
	     (source_id__h31729 == 10'd16 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1017) ?
	       wdata32__h27246[2] :
	       _dfoo1872 ;
  assign _dfoo1941 =
	     source_id__h31729 == 10'd15 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1017 ||
	     source_id__h33225 == 10'd15 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1078 ||
	     _dfoo1805 ;
  assign _dfoo1942 =
	     (source_id__h31729 == 10'd15 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1017) ?
	       wdata32__h27246[2] :
	       _dfoo1874 ;
  assign _dfoo1943 =
	     source_id__h31729 == 10'd14 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1017 ||
	     source_id__h33225 == 10'd14 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1078 ||
	     _dfoo1807 ;
  assign _dfoo1944 =
	     (source_id__h31729 == 10'd14 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1017) ?
	       wdata32__h27246[2] :
	       _dfoo1876 ;
  assign _dfoo1945 =
	     source_id__h31729 == 10'd13 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1017 ||
	     source_id__h33225 == 10'd13 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1078 ||
	     _dfoo1809 ;
  assign _dfoo1946 =
	     (source_id__h31729 == 10'd13 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1017) ?
	       wdata32__h27246[2] :
	       _dfoo1878 ;
  assign _dfoo1947 =
	     source_id__h31729 == 10'd12 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1017 ||
	     source_id__h33225 == 10'd12 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1078 ||
	     _dfoo1811 ;
  assign _dfoo1948 =
	     (source_id__h31729 == 10'd12 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1017) ?
	       wdata32__h27246[2] :
	       _dfoo1880 ;
  assign _dfoo1949 =
	     source_id__h31729 == 10'd11 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1017 ||
	     source_id__h33225 == 10'd11 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1078 ||
	     _dfoo1813 ;
  assign _dfoo195 =
	     source_id__h70625 == 10'd4 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2603 ||
	     source_id__h72121 == 10'd4 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2664 ||
	     _dfoo59 ;
  assign _dfoo1950 =
	     (source_id__h31729 == 10'd11 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1017) ?
	       wdata32__h27246[2] :
	       _dfoo1882 ;
  assign _dfoo1951 =
	     source_id__h31729 == 10'd10 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1017 ||
	     source_id__h33225 == 10'd10 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1078 ||
	     _dfoo1815 ;
  assign _dfoo1952 =
	     (source_id__h31729 == 10'd10 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1017) ?
	       wdata32__h27246[2] :
	       _dfoo1884 ;
  assign _dfoo1953 =
	     source_id__h31729 == 10'd9 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1017 ||
	     source_id__h33225 == 10'd9 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1078 ||
	     _dfoo1817 ;
  assign _dfoo1954 =
	     (source_id__h31729 == 10'd9 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1017) ?
	       wdata32__h27246[2] :
	       _dfoo1886 ;
  assign _dfoo1955 =
	     source_id__h31729 == 10'd8 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1017 ||
	     source_id__h33225 == 10'd8 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1078 ||
	     _dfoo1819 ;
  assign _dfoo1956 =
	     (source_id__h31729 == 10'd8 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1017) ?
	       wdata32__h27246[2] :
	       _dfoo1888 ;
  assign _dfoo1957 =
	     source_id__h31729 == 10'd7 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1017 ||
	     source_id__h33225 == 10'd7 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1078 ||
	     _dfoo1821 ;
  assign _dfoo1958 =
	     (source_id__h31729 == 10'd7 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1017) ?
	       wdata32__h27246[2] :
	       _dfoo1890 ;
  assign _dfoo1959 =
	     source_id__h31729 == 10'd6 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1017 ||
	     source_id__h33225 == 10'd6 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1078 ||
	     _dfoo1823 ;
  assign _dfoo196 =
	     (source_id__h70625 == 10'd4 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2603) ?
	       wdata32__h27246[28] :
	       _dfoo128 ;
  assign _dfoo1960 =
	     (source_id__h31729 == 10'd6 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1017) ?
	       wdata32__h27246[2] :
	       _dfoo1892 ;
  assign _dfoo1961 =
	     source_id__h31729 == 10'd5 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1017 ||
	     source_id__h33225 == 10'd5 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1078 ||
	     _dfoo1825 ;
  assign _dfoo1962 =
	     (source_id__h31729 == 10'd5 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1017) ?
	       wdata32__h27246[2] :
	       _dfoo1894 ;
  assign _dfoo1963 =
	     source_id__h31729 == 10'd4 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1017 ||
	     source_id__h33225 == 10'd4 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1078 ||
	     _dfoo1827 ;
  assign _dfoo1964 =
	     (source_id__h31729 == 10'd4 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1017) ?
	       wdata32__h27246[2] :
	       _dfoo1896 ;
  assign _dfoo1965 =
	     source_id__h31729 == 10'd3 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1017 ||
	     source_id__h33225 == 10'd3 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1078 ||
	     _dfoo1829 ;
  assign _dfoo1966 =
	     (source_id__h31729 == 10'd3 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1017) ?
	       wdata32__h27246[2] :
	       _dfoo1898 ;
  assign _dfoo1967 =
	     source_id__h31729 == 10'd2 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1017 ||
	     source_id__h33225 == 10'd2 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1078 ||
	     _dfoo1831 ;
  assign _dfoo1968 =
	     (source_id__h31729 == 10'd2 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1017) ?
	       wdata32__h27246[2] :
	       _dfoo1900 ;
  assign _dfoo1969 =
	     source_id__h31729 == 10'd1 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1017 ||
	     source_id__h33225 == 10'd1 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1078 ||
	     _dfoo1833 ;
  assign _dfoo197 =
	     source_id__h70625 == 10'd3 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2603 ||
	     source_id__h72121 == 10'd3 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2664 ||
	     _dfoo61 ;
  assign _dfoo1970 =
	     (source_id__h31729 == 10'd1 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1017) ?
	       wdata32__h27246[2] :
	       _dfoo1902 ;
  assign _dfoo1971 =
	     source_id__h31729 == 10'd0 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1017 ||
	     source_id__h33225 == 10'd0 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1078 ||
	     _dfoo1835 ;
  assign _dfoo1972 =
	     (source_id__h31729 == 10'd0 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1017) ?
	       wdata32__h27246[2] :
	       _dfoo1904 ;
  assign _dfoo1974 =
	     (source_id__h30233 == 10'd16 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d956) ?
	       wdata32__h27246[1] :
	       _dfoo1906 ;
  assign _dfoo1976 =
	     (source_id__h30233 == 10'd15 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d956) ?
	       wdata32__h27246[1] :
	       _dfoo1908 ;
  assign _dfoo1978 =
	     (source_id__h30233 == 10'd14 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d956) ?
	       wdata32__h27246[1] :
	       _dfoo1910 ;
  assign _dfoo198 =
	     (source_id__h70625 == 10'd3 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2603) ?
	       wdata32__h27246[28] :
	       _dfoo130 ;
  assign _dfoo1980 =
	     (source_id__h30233 == 10'd13 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d956) ?
	       wdata32__h27246[1] :
	       _dfoo1912 ;
  assign _dfoo1982 =
	     (source_id__h30233 == 10'd12 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d956) ?
	       wdata32__h27246[1] :
	       _dfoo1914 ;
  assign _dfoo1984 =
	     (source_id__h30233 == 10'd11 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d956) ?
	       wdata32__h27246[1] :
	       _dfoo1916 ;
  assign _dfoo1986 =
	     (source_id__h30233 == 10'd10 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d956) ?
	       wdata32__h27246[1] :
	       _dfoo1918 ;
  assign _dfoo1988 =
	     (source_id__h30233 == 10'd9 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d956) ?
	       wdata32__h27246[1] :
	       _dfoo1920 ;
  assign _dfoo199 =
	     source_id__h70625 == 10'd2 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2603 ||
	     source_id__h72121 == 10'd2 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2664 ||
	     _dfoo63 ;
  assign _dfoo1990 =
	     (source_id__h30233 == 10'd8 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d956) ?
	       wdata32__h27246[1] :
	       _dfoo1922 ;
  assign _dfoo1992 =
	     (source_id__h30233 == 10'd7 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d956) ?
	       wdata32__h27246[1] :
	       _dfoo1924 ;
  assign _dfoo1994 =
	     (source_id__h30233 == 10'd6 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d956) ?
	       wdata32__h27246[1] :
	       _dfoo1926 ;
  assign _dfoo1996 =
	     (source_id__h30233 == 10'd5 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d956) ?
	       wdata32__h27246[1] :
	       _dfoo1928 ;
  assign _dfoo1998 =
	     (source_id__h30233 == 10'd4 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d956) ?
	       wdata32__h27246[1] :
	       _dfoo1930 ;
  assign _dfoo2 =
	     (source_id__h73617 == 10'd16 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2725) ?
	       wdata32__h27246[30] :
	       wdata32__h27246[31] ;
  assign _dfoo20 =
	     (source_id__h73617 == 10'd7 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2725) ?
	       wdata32__h27246[30] :
	       wdata32__h27246[31] ;
  assign _dfoo200 =
	     (source_id__h70625 == 10'd2 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2603) ?
	       wdata32__h27246[28] :
	       _dfoo132 ;
  assign _dfoo2000 =
	     (source_id__h30233 == 10'd3 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d956) ?
	       wdata32__h27246[1] :
	       _dfoo1932 ;
  assign _dfoo2002 =
	     (source_id__h30233 == 10'd2 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d956) ?
	       wdata32__h27246[1] :
	       _dfoo1934 ;
  assign _dfoo2004 =
	     (source_id__h30233 == 10'd1 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d956) ?
	       wdata32__h27246[1] :
	       _dfoo1936 ;
  assign _dfoo2006 =
	     (source_id__h30233 == 10'd0 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d956) ?
	       wdata32__h27246[1] :
	       _dfoo1938 ;
  assign _dfoo2008 =
	     (source_id__h30233 == 10'd16 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d956) ?
	       wdata32__h27246[1] :
	       _dfoo1940 ;
  assign _dfoo201 =
	     source_id__h70625 == 10'd1 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2603 ||
	     source_id__h72121 == 10'd1 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2664 ||
	     _dfoo65 ;
  assign _dfoo2010 =
	     (source_id__h30233 == 10'd15 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d956) ?
	       wdata32__h27246[1] :
	       _dfoo1942 ;
  assign _dfoo2012 =
	     (source_id__h30233 == 10'd14 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d956) ?
	       wdata32__h27246[1] :
	       _dfoo1944 ;
  assign _dfoo2014 =
	     (source_id__h30233 == 10'd13 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d956) ?
	       wdata32__h27246[1] :
	       _dfoo1946 ;
  assign _dfoo2016 =
	     (source_id__h30233 == 10'd12 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d956) ?
	       wdata32__h27246[1] :
	       _dfoo1948 ;
  assign _dfoo2018 =
	     (source_id__h30233 == 10'd11 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d956) ?
	       wdata32__h27246[1] :
	       _dfoo1950 ;
  assign _dfoo202 =
	     (source_id__h70625 == 10'd1 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2603) ?
	       wdata32__h27246[28] :
	       _dfoo134 ;
  assign _dfoo2020 =
	     (source_id__h30233 == 10'd10 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d956) ?
	       wdata32__h27246[1] :
	       _dfoo1952 ;
  assign _dfoo2022 =
	     (source_id__h30233 == 10'd9 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d956) ?
	       wdata32__h27246[1] :
	       _dfoo1954 ;
  assign _dfoo2024 =
	     (source_id__h30233 == 10'd8 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d956) ?
	       wdata32__h27246[1] :
	       _dfoo1956 ;
  assign _dfoo2026 =
	     (source_id__h30233 == 10'd7 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d956) ?
	       wdata32__h27246[1] :
	       _dfoo1958 ;
  assign _dfoo2028 =
	     (source_id__h30233 == 10'd6 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d956) ?
	       wdata32__h27246[1] :
	       _dfoo1960 ;
  assign _dfoo203 =
	     source_id__h70625 == 10'd0 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2603 ||
	     source_id__h72121 == 10'd0 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2664 ||
	     _dfoo67 ;
  assign _dfoo2030 =
	     (source_id__h30233 == 10'd5 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d956) ?
	       wdata32__h27246[1] :
	       _dfoo1962 ;
  assign _dfoo2032 =
	     (source_id__h30233 == 10'd4 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d956) ?
	       wdata32__h27246[1] :
	       _dfoo1964 ;
  assign _dfoo2034 =
	     (source_id__h30233 == 10'd3 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d956) ?
	       wdata32__h27246[1] :
	       _dfoo1966 ;
  assign _dfoo2036 =
	     (source_id__h30233 == 10'd2 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d956) ?
	       wdata32__h27246[1] :
	       _dfoo1968 ;
  assign _dfoo2038 =
	     (source_id__h30233 == 10'd1 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d956) ?
	       wdata32__h27246[1] :
	       _dfoo1970 ;
  assign _dfoo204 =
	     (source_id__h70625 == 10'd0 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2603) ?
	       wdata32__h27246[28] :
	       _dfoo136 ;
  assign _dfoo2040 =
	     (source_id__h30233 == 10'd0 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d956) ?
	       wdata32__h27246[1] :
	       _dfoo1972 ;
  assign _dfoo2041 =
	     source_id_base__h28620 == 10'd16 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d931 ||
	     source_id__h30233 == 10'd16 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d956 ||
	     _dfoo1905 ;
  assign _dfoo2043 =
	     source_id_base__h28620 == 10'd15 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d931 ||
	     source_id__h30233 == 10'd15 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d956 ||
	     _dfoo1907 ;
  assign _dfoo2045 =
	     source_id_base__h28620 == 10'd14 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d931 ||
	     source_id__h30233 == 10'd14 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d956 ||
	     _dfoo1909 ;
  assign _dfoo2047 =
	     source_id_base__h28620 == 10'd13 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d931 ||
	     source_id__h30233 == 10'd13 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d956 ||
	     _dfoo1911 ;
  assign _dfoo2049 =
	     source_id_base__h28620 == 10'd12 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d931 ||
	     source_id__h30233 == 10'd12 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d956 ||
	     _dfoo1913 ;
  assign _dfoo2051 =
	     source_id_base__h28620 == 10'd11 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d931 ||
	     source_id__h30233 == 10'd11 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d956 ||
	     _dfoo1915 ;
  assign _dfoo2053 =
	     source_id_base__h28620 == 10'd10 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d931 ||
	     source_id__h30233 == 10'd10 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d956 ||
	     _dfoo1917 ;
  assign _dfoo2055 =
	     source_id_base__h28620 == 10'd9 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d931 ||
	     source_id__h30233 == 10'd9 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d956 ||
	     _dfoo1919 ;
  assign _dfoo2057 =
	     source_id_base__h28620 == 10'd8 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d931 ||
	     source_id__h30233 == 10'd8 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d956 ||
	     _dfoo1921 ;
  assign _dfoo2059 =
	     source_id_base__h28620 == 10'd7 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d931 ||
	     source_id__h30233 == 10'd7 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d956 ||
	     _dfoo1923 ;
  assign _dfoo206 =
	     (source_id__h69129 == 10'd16 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2542) ?
	       wdata32__h27246[27] :
	       _dfoo138 ;
  assign _dfoo2061 =
	     source_id_base__h28620 == 10'd6 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d931 ||
	     source_id__h30233 == 10'd6 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d956 ||
	     _dfoo1925 ;
  assign _dfoo2063 =
	     source_id_base__h28620 == 10'd5 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d931 ||
	     source_id__h30233 == 10'd5 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d956 ||
	     _dfoo1927 ;
  assign _dfoo2065 =
	     source_id_base__h28620 == 10'd4 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d931 ||
	     source_id__h30233 == 10'd4 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d956 ||
	     _dfoo1929 ;
  assign _dfoo2067 =
	     source_id_base__h28620 == 10'd3 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d931 ||
	     source_id__h30233 == 10'd3 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d956 ||
	     _dfoo1931 ;
  assign _dfoo2069 =
	     source_id_base__h28620 == 10'd2 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d931 ||
	     source_id__h30233 == 10'd2 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d956 ||
	     _dfoo1933 ;
  assign _dfoo2071 =
	     source_id_base__h28620 == 10'd1 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d931 ||
	     source_id__h30233 == 10'd1 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d956 ||
	     _dfoo1935 ;
  assign _dfoo2073 =
	     source_id_base__h28620 == 10'd0 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d931 ||
	     source_id__h30233 == 10'd0 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d956 ||
	     _dfoo1937 ;
  assign _dfoo2075 =
	     source_id_base__h28620 == 10'd16 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d895 ||
	     source_id__h30233 == 10'd16 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d956 ||
	     _dfoo1939 ;
  assign _dfoo2077 =
	     source_id_base__h28620 == 10'd15 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d895 ||
	     source_id__h30233 == 10'd15 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d956 ||
	     _dfoo1941 ;
  assign _dfoo2079 =
	     source_id_base__h28620 == 10'd14 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d895 ||
	     source_id__h30233 == 10'd14 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d956 ||
	     _dfoo1943 ;
  assign _dfoo208 =
	     (source_id__h69129 == 10'd15 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2542) ?
	       wdata32__h27246[27] :
	       _dfoo140 ;
  assign _dfoo2081 =
	     source_id_base__h28620 == 10'd13 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d895 ||
	     source_id__h30233 == 10'd13 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d956 ||
	     _dfoo1945 ;
  assign _dfoo2083 =
	     source_id_base__h28620 == 10'd12 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d895 ||
	     source_id__h30233 == 10'd12 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d956 ||
	     _dfoo1947 ;
  assign _dfoo2085 =
	     source_id_base__h28620 == 10'd11 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d895 ||
	     source_id__h30233 == 10'd11 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d956 ||
	     _dfoo1949 ;
  assign _dfoo2087 =
	     source_id_base__h28620 == 10'd10 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d895 ||
	     source_id__h30233 == 10'd10 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d956 ||
	     _dfoo1951 ;
  assign _dfoo2089 =
	     source_id_base__h28620 == 10'd9 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d895 ||
	     source_id__h30233 == 10'd9 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d956 ||
	     _dfoo1953 ;
  assign _dfoo2091 =
	     source_id_base__h28620 == 10'd8 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d895 ||
	     source_id__h30233 == 10'd8 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d956 ||
	     _dfoo1955 ;
  assign _dfoo2093 =
	     source_id_base__h28620 == 10'd7 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d895 ||
	     source_id__h30233 == 10'd7 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d956 ||
	     _dfoo1957 ;
  assign _dfoo2095 =
	     source_id_base__h28620 == 10'd6 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d895 ||
	     source_id__h30233 == 10'd6 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d956 ||
	     _dfoo1959 ;
  assign _dfoo2097 =
	     source_id_base__h28620 == 10'd5 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d895 ||
	     source_id__h30233 == 10'd5 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d956 ||
	     _dfoo1961 ;
  assign _dfoo2099 =
	     source_id_base__h28620 == 10'd4 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d895 ||
	     source_id__h30233 == 10'd4 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d956 ||
	     _dfoo1963 ;
  assign _dfoo21 =
	     source_id__h73617 == 10'd6 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2725 ||
	     source_id__h75113 == 10'd6 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2786 ;
  assign _dfoo210 =
	     (source_id__h69129 == 10'd14 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2542) ?
	       wdata32__h27246[27] :
	       _dfoo142 ;
  assign _dfoo2101 =
	     source_id_base__h28620 == 10'd3 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d895 ||
	     source_id__h30233 == 10'd3 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d956 ||
	     _dfoo1965 ;
  assign _dfoo2103 =
	     source_id_base__h28620 == 10'd2 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d895 ||
	     source_id__h30233 == 10'd2 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d956 ||
	     _dfoo1967 ;
  assign _dfoo2105 =
	     source_id_base__h28620 == 10'd1 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d895 ||
	     source_id__h30233 == 10'd1 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d956 ||
	     _dfoo1969 ;
  assign _dfoo2107 =
	     source_id_base__h28620 == 10'd0 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d895 ||
	     source_id__h30233 == 10'd0 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d956 ||
	     _dfoo1971 ;
  assign _dfoo212 =
	     (source_id__h69129 == 10'd13 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2542) ?
	       wdata32__h27246[27] :
	       _dfoo144 ;
  assign _dfoo214 =
	     (source_id__h69129 == 10'd12 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2542) ?
	       wdata32__h27246[27] :
	       _dfoo146 ;
  assign _dfoo216 =
	     (source_id__h69129 == 10'd11 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2542) ?
	       wdata32__h27246[27] :
	       _dfoo148 ;
  assign _dfoo218 =
	     (source_id__h69129 == 10'd10 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2542) ?
	       wdata32__h27246[27] :
	       _dfoo150 ;
  assign _dfoo22 =
	     (source_id__h73617 == 10'd6 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2725) ?
	       wdata32__h27246[30] :
	       wdata32__h27246[31] ;
  assign _dfoo220 =
	     (source_id__h69129 == 10'd9 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2542) ?
	       wdata32__h27246[27] :
	       _dfoo152 ;
  assign _dfoo222 =
	     (source_id__h69129 == 10'd8 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2542) ?
	       wdata32__h27246[27] :
	       _dfoo154 ;
  assign _dfoo224 =
	     (source_id__h69129 == 10'd7 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2542) ?
	       wdata32__h27246[27] :
	       _dfoo156 ;
  assign _dfoo226 =
	     (source_id__h69129 == 10'd6 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2542) ?
	       wdata32__h27246[27] :
	       _dfoo158 ;
  assign _dfoo228 =
	     (source_id__h69129 == 10'd5 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2542) ?
	       wdata32__h27246[27] :
	       _dfoo160 ;
  assign _dfoo23 =
	     source_id__h73617 == 10'd5 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2725 ||
	     source_id__h75113 == 10'd5 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2786 ;
  assign _dfoo230 =
	     (source_id__h69129 == 10'd4 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2542) ?
	       wdata32__h27246[27] :
	       _dfoo162 ;
  assign _dfoo232 =
	     (source_id__h69129 == 10'd3 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2542) ?
	       wdata32__h27246[27] :
	       _dfoo164 ;
  assign _dfoo234 =
	     (source_id__h69129 == 10'd2 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2542) ?
	       wdata32__h27246[27] :
	       _dfoo166 ;
  assign _dfoo236 =
	     (source_id__h69129 == 10'd1 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2542) ?
	       wdata32__h27246[27] :
	       _dfoo168 ;
  assign _dfoo238 =
	     (source_id__h69129 == 10'd0 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2542) ?
	       wdata32__h27246[27] :
	       _dfoo170 ;
  assign _dfoo24 =
	     (source_id__h73617 == 10'd5 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2725) ?
	       wdata32__h27246[30] :
	       wdata32__h27246[31] ;
  assign _dfoo240 =
	     (source_id__h69129 == 10'd16 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2542) ?
	       wdata32__h27246[27] :
	       _dfoo172 ;
  assign _dfoo242 =
	     (source_id__h69129 == 10'd15 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2542) ?
	       wdata32__h27246[27] :
	       _dfoo174 ;
  assign _dfoo244 =
	     (source_id__h69129 == 10'd14 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2542) ?
	       wdata32__h27246[27] :
	       _dfoo176 ;
  assign _dfoo246 =
	     (source_id__h69129 == 10'd13 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2542) ?
	       wdata32__h27246[27] :
	       _dfoo178 ;
  assign _dfoo248 =
	     (source_id__h69129 == 10'd12 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2542) ?
	       wdata32__h27246[27] :
	       _dfoo180 ;
  assign _dfoo25 =
	     source_id__h73617 == 10'd4 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2725 ||
	     source_id__h75113 == 10'd4 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2786 ;
  assign _dfoo250 =
	     (source_id__h69129 == 10'd11 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2542) ?
	       wdata32__h27246[27] :
	       _dfoo182 ;
  assign _dfoo252 =
	     (source_id__h69129 == 10'd10 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2542) ?
	       wdata32__h27246[27] :
	       _dfoo184 ;
  assign _dfoo254 =
	     (source_id__h69129 == 10'd9 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2542) ?
	       wdata32__h27246[27] :
	       _dfoo186 ;
  assign _dfoo256 =
	     (source_id__h69129 == 10'd8 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2542) ?
	       wdata32__h27246[27] :
	       _dfoo188 ;
  assign _dfoo258 =
	     (source_id__h69129 == 10'd7 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2542) ?
	       wdata32__h27246[27] :
	       _dfoo190 ;
  assign _dfoo26 =
	     (source_id__h73617 == 10'd4 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2725) ?
	       wdata32__h27246[30] :
	       wdata32__h27246[31] ;
  assign _dfoo260 =
	     (source_id__h69129 == 10'd6 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2542) ?
	       wdata32__h27246[27] :
	       _dfoo192 ;
  assign _dfoo262 =
	     (source_id__h69129 == 10'd5 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2542) ?
	       wdata32__h27246[27] :
	       _dfoo194 ;
  assign _dfoo264 =
	     (source_id__h69129 == 10'd4 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2542) ?
	       wdata32__h27246[27] :
	       _dfoo196 ;
  assign _dfoo266 =
	     (source_id__h69129 == 10'd3 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2542) ?
	       wdata32__h27246[27] :
	       _dfoo198 ;
  assign _dfoo268 =
	     (source_id__h69129 == 10'd2 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2542) ?
	       wdata32__h27246[27] :
	       _dfoo200 ;
  assign _dfoo27 =
	     source_id__h73617 == 10'd3 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2725 ||
	     source_id__h75113 == 10'd3 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2786 ;
  assign _dfoo270 =
	     (source_id__h69129 == 10'd1 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2542) ?
	       wdata32__h27246[27] :
	       _dfoo202 ;
  assign _dfoo272 =
	     (source_id__h69129 == 10'd0 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2542) ?
	       wdata32__h27246[27] :
	       _dfoo204 ;
  assign _dfoo273 =
	     source_id__h67633 == 10'd16 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2481 ||
	     source_id__h69129 == 10'd16 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2542 ||
	     _dfoo137 ;
  assign _dfoo274 =
	     (source_id__h67633 == 10'd16 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2481) ?
	       wdata32__h27246[26] :
	       _dfoo206 ;
  assign _dfoo275 =
	     source_id__h67633 == 10'd15 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2481 ||
	     source_id__h69129 == 10'd15 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2542 ||
	     _dfoo139 ;
  assign _dfoo276 =
	     (source_id__h67633 == 10'd15 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2481) ?
	       wdata32__h27246[26] :
	       _dfoo208 ;
  assign _dfoo277 =
	     source_id__h67633 == 10'd14 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2481 ||
	     source_id__h69129 == 10'd14 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2542 ||
	     _dfoo141 ;
  assign _dfoo278 =
	     (source_id__h67633 == 10'd14 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2481) ?
	       wdata32__h27246[26] :
	       _dfoo210 ;
  assign _dfoo279 =
	     source_id__h67633 == 10'd13 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2481 ||
	     source_id__h69129 == 10'd13 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2542 ||
	     _dfoo143 ;
  assign _dfoo28 =
	     (source_id__h73617 == 10'd3 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2725) ?
	       wdata32__h27246[30] :
	       wdata32__h27246[31] ;
  assign _dfoo280 =
	     (source_id__h67633 == 10'd13 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2481) ?
	       wdata32__h27246[26] :
	       _dfoo212 ;
  assign _dfoo281 =
	     source_id__h67633 == 10'd12 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2481 ||
	     source_id__h69129 == 10'd12 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2542 ||
	     _dfoo145 ;
  assign _dfoo282 =
	     (source_id__h67633 == 10'd12 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2481) ?
	       wdata32__h27246[26] :
	       _dfoo214 ;
  assign _dfoo283 =
	     source_id__h67633 == 10'd11 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2481 ||
	     source_id__h69129 == 10'd11 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2542 ||
	     _dfoo147 ;
  assign _dfoo284 =
	     (source_id__h67633 == 10'd11 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2481) ?
	       wdata32__h27246[26] :
	       _dfoo216 ;
  assign _dfoo285 =
	     source_id__h67633 == 10'd10 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2481 ||
	     source_id__h69129 == 10'd10 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2542 ||
	     _dfoo149 ;
  assign _dfoo286 =
	     (source_id__h67633 == 10'd10 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2481) ?
	       wdata32__h27246[26] :
	       _dfoo218 ;
  assign _dfoo287 =
	     source_id__h67633 == 10'd9 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2481 ||
	     source_id__h69129 == 10'd9 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2542 ||
	     _dfoo151 ;
  assign _dfoo288 =
	     (source_id__h67633 == 10'd9 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2481) ?
	       wdata32__h27246[26] :
	       _dfoo220 ;
  assign _dfoo289 =
	     source_id__h67633 == 10'd8 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2481 ||
	     source_id__h69129 == 10'd8 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2542 ||
	     _dfoo153 ;
  assign _dfoo29 =
	     source_id__h73617 == 10'd2 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2725 ||
	     source_id__h75113 == 10'd2 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2786 ;
  assign _dfoo290 =
	     (source_id__h67633 == 10'd8 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2481) ?
	       wdata32__h27246[26] :
	       _dfoo222 ;
  assign _dfoo291 =
	     source_id__h67633 == 10'd7 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2481 ||
	     source_id__h69129 == 10'd7 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2542 ||
	     _dfoo155 ;
  assign _dfoo292 =
	     (source_id__h67633 == 10'd7 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2481) ?
	       wdata32__h27246[26] :
	       _dfoo224 ;
  assign _dfoo293 =
	     source_id__h67633 == 10'd6 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2481 ||
	     source_id__h69129 == 10'd6 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2542 ||
	     _dfoo157 ;
  assign _dfoo294 =
	     (source_id__h67633 == 10'd6 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2481) ?
	       wdata32__h27246[26] :
	       _dfoo226 ;
  assign _dfoo295 =
	     source_id__h67633 == 10'd5 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2481 ||
	     source_id__h69129 == 10'd5 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2542 ||
	     _dfoo159 ;
  assign _dfoo296 =
	     (source_id__h67633 == 10'd5 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2481) ?
	       wdata32__h27246[26] :
	       _dfoo228 ;
  assign _dfoo297 =
	     source_id__h67633 == 10'd4 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2481 ||
	     source_id__h69129 == 10'd4 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2542 ||
	     _dfoo161 ;
  assign _dfoo298 =
	     (source_id__h67633 == 10'd4 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2481) ?
	       wdata32__h27246[26] :
	       _dfoo230 ;
  assign _dfoo299 =
	     source_id__h67633 == 10'd3 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2481 ||
	     source_id__h69129 == 10'd3 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2542 ||
	     _dfoo163 ;
  assign _dfoo3 =
	     source_id__h73617 == 10'd15 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2725 ||
	     source_id__h75113 == 10'd15 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2786 ;
  assign _dfoo30 =
	     (source_id__h73617 == 10'd2 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2725) ?
	       wdata32__h27246[30] :
	       wdata32__h27246[31] ;
  assign _dfoo300 =
	     (source_id__h67633 == 10'd3 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2481) ?
	       wdata32__h27246[26] :
	       _dfoo232 ;
  assign _dfoo301 =
	     source_id__h67633 == 10'd2 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2481 ||
	     source_id__h69129 == 10'd2 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2542 ||
	     _dfoo165 ;
  assign _dfoo302 =
	     (source_id__h67633 == 10'd2 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2481) ?
	       wdata32__h27246[26] :
	       _dfoo234 ;
  assign _dfoo303 =
	     source_id__h67633 == 10'd1 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2481 ||
	     source_id__h69129 == 10'd1 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2542 ||
	     _dfoo167 ;
  assign _dfoo304 =
	     (source_id__h67633 == 10'd1 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2481) ?
	       wdata32__h27246[26] :
	       _dfoo236 ;
  assign _dfoo305 =
	     source_id__h67633 == 10'd0 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2481 ||
	     source_id__h69129 == 10'd0 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2542 ||
	     _dfoo169 ;
  assign _dfoo306 =
	     (source_id__h67633 == 10'd0 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2481) ?
	       wdata32__h27246[26] :
	       _dfoo238 ;
  assign _dfoo307 =
	     source_id__h67633 == 10'd16 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2481 ||
	     source_id__h69129 == 10'd16 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2542 ||
	     _dfoo171 ;
  assign _dfoo308 =
	     (source_id__h67633 == 10'd16 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2481) ?
	       wdata32__h27246[26] :
	       _dfoo240 ;
  assign _dfoo309 =
	     source_id__h67633 == 10'd15 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2481 ||
	     source_id__h69129 == 10'd15 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2542 ||
	     _dfoo173 ;
  assign _dfoo31 =
	     source_id__h73617 == 10'd1 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2725 ||
	     source_id__h75113 == 10'd1 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2786 ;
  assign _dfoo310 =
	     (source_id__h67633 == 10'd15 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2481) ?
	       wdata32__h27246[26] :
	       _dfoo242 ;
  assign _dfoo311 =
	     source_id__h67633 == 10'd14 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2481 ||
	     source_id__h69129 == 10'd14 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2542 ||
	     _dfoo175 ;
  assign _dfoo312 =
	     (source_id__h67633 == 10'd14 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2481) ?
	       wdata32__h27246[26] :
	       _dfoo244 ;
  assign _dfoo313 =
	     source_id__h67633 == 10'd13 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2481 ||
	     source_id__h69129 == 10'd13 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2542 ||
	     _dfoo177 ;
  assign _dfoo314 =
	     (source_id__h67633 == 10'd13 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2481) ?
	       wdata32__h27246[26] :
	       _dfoo246 ;
  assign _dfoo315 =
	     source_id__h67633 == 10'd12 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2481 ||
	     source_id__h69129 == 10'd12 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2542 ||
	     _dfoo179 ;
  assign _dfoo316 =
	     (source_id__h67633 == 10'd12 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2481) ?
	       wdata32__h27246[26] :
	       _dfoo248 ;
  assign _dfoo317 =
	     source_id__h67633 == 10'd11 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2481 ||
	     source_id__h69129 == 10'd11 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2542 ||
	     _dfoo181 ;
  assign _dfoo318 =
	     (source_id__h67633 == 10'd11 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2481) ?
	       wdata32__h27246[26] :
	       _dfoo250 ;
  assign _dfoo319 =
	     source_id__h67633 == 10'd10 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2481 ||
	     source_id__h69129 == 10'd10 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2542 ||
	     _dfoo183 ;
  assign _dfoo32 =
	     (source_id__h73617 == 10'd1 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2725) ?
	       wdata32__h27246[30] :
	       wdata32__h27246[31] ;
  assign _dfoo320 =
	     (source_id__h67633 == 10'd10 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2481) ?
	       wdata32__h27246[26] :
	       _dfoo252 ;
  assign _dfoo321 =
	     source_id__h67633 == 10'd9 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2481 ||
	     source_id__h69129 == 10'd9 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2542 ||
	     _dfoo185 ;
  assign _dfoo322 =
	     (source_id__h67633 == 10'd9 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2481) ?
	       wdata32__h27246[26] :
	       _dfoo254 ;
  assign _dfoo323 =
	     source_id__h67633 == 10'd8 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2481 ||
	     source_id__h69129 == 10'd8 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2542 ||
	     _dfoo187 ;
  assign _dfoo324 =
	     (source_id__h67633 == 10'd8 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2481) ?
	       wdata32__h27246[26] :
	       _dfoo256 ;
  assign _dfoo325 =
	     source_id__h67633 == 10'd7 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2481 ||
	     source_id__h69129 == 10'd7 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2542 ||
	     _dfoo189 ;
  assign _dfoo326 =
	     (source_id__h67633 == 10'd7 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2481) ?
	       wdata32__h27246[26] :
	       _dfoo258 ;
  assign _dfoo327 =
	     source_id__h67633 == 10'd6 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2481 ||
	     source_id__h69129 == 10'd6 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2542 ||
	     _dfoo191 ;
  assign _dfoo328 =
	     (source_id__h67633 == 10'd6 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2481) ?
	       wdata32__h27246[26] :
	       _dfoo260 ;
  assign _dfoo329 =
	     source_id__h67633 == 10'd5 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2481 ||
	     source_id__h69129 == 10'd5 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2542 ||
	     _dfoo193 ;
  assign _dfoo33 =
	     source_id__h73617 == 10'd0 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2725 ||
	     source_id__h75113 == 10'd0 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2786 ;
  assign _dfoo330 =
	     (source_id__h67633 == 10'd5 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2481) ?
	       wdata32__h27246[26] :
	       _dfoo262 ;
  assign _dfoo331 =
	     source_id__h67633 == 10'd4 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2481 ||
	     source_id__h69129 == 10'd4 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2542 ||
	     _dfoo195 ;
  assign _dfoo332 =
	     (source_id__h67633 == 10'd4 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2481) ?
	       wdata32__h27246[26] :
	       _dfoo264 ;
  assign _dfoo333 =
	     source_id__h67633 == 10'd3 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2481 ||
	     source_id__h69129 == 10'd3 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2542 ||
	     _dfoo197 ;
  assign _dfoo334 =
	     (source_id__h67633 == 10'd3 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2481) ?
	       wdata32__h27246[26] :
	       _dfoo266 ;
  assign _dfoo335 =
	     source_id__h67633 == 10'd2 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2481 ||
	     source_id__h69129 == 10'd2 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2542 ||
	     _dfoo199 ;
  assign _dfoo336 =
	     (source_id__h67633 == 10'd2 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2481) ?
	       wdata32__h27246[26] :
	       _dfoo268 ;
  assign _dfoo337 =
	     source_id__h67633 == 10'd1 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2481 ||
	     source_id__h69129 == 10'd1 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2542 ||
	     _dfoo201 ;
  assign _dfoo338 =
	     (source_id__h67633 == 10'd1 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2481) ?
	       wdata32__h27246[26] :
	       _dfoo270 ;
  assign _dfoo339 =
	     source_id__h67633 == 10'd0 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2481 ||
	     source_id__h69129 == 10'd0 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2542 ||
	     _dfoo203 ;
  assign _dfoo34 =
	     (source_id__h73617 == 10'd0 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2725) ?
	       wdata32__h27246[30] :
	       wdata32__h27246[31] ;
  assign _dfoo340 =
	     (source_id__h67633 == 10'd0 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2481) ?
	       wdata32__h27246[26] :
	       _dfoo272 ;
  assign _dfoo342 =
	     (source_id__h66137 == 10'd16 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2420) ?
	       wdata32__h27246[25] :
	       _dfoo274 ;
  assign _dfoo344 =
	     (source_id__h66137 == 10'd15 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2420) ?
	       wdata32__h27246[25] :
	       _dfoo276 ;
  assign _dfoo346 =
	     (source_id__h66137 == 10'd14 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2420) ?
	       wdata32__h27246[25] :
	       _dfoo278 ;
  assign _dfoo348 =
	     (source_id__h66137 == 10'd13 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2420) ?
	       wdata32__h27246[25] :
	       _dfoo280 ;
  assign _dfoo35 =
	     source_id__h73617 == 10'd16 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2725 ||
	     source_id__h75113 == 10'd16 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2786 ;
  assign _dfoo350 =
	     (source_id__h66137 == 10'd12 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2420) ?
	       wdata32__h27246[25] :
	       _dfoo282 ;
  assign _dfoo352 =
	     (source_id__h66137 == 10'd11 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2420) ?
	       wdata32__h27246[25] :
	       _dfoo284 ;
  assign _dfoo354 =
	     (source_id__h66137 == 10'd10 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2420) ?
	       wdata32__h27246[25] :
	       _dfoo286 ;
  assign _dfoo356 =
	     (source_id__h66137 == 10'd9 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2420) ?
	       wdata32__h27246[25] :
	       _dfoo288 ;
  assign _dfoo358 =
	     (source_id__h66137 == 10'd8 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2420) ?
	       wdata32__h27246[25] :
	       _dfoo290 ;
  assign _dfoo36 =
	     (source_id__h73617 == 10'd16 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2725) ?
	       wdata32__h27246[30] :
	       wdata32__h27246[31] ;
  assign _dfoo360 =
	     (source_id__h66137 == 10'd7 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2420) ?
	       wdata32__h27246[25] :
	       _dfoo292 ;
  assign _dfoo362 =
	     (source_id__h66137 == 10'd6 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2420) ?
	       wdata32__h27246[25] :
	       _dfoo294 ;
  assign _dfoo364 =
	     (source_id__h66137 == 10'd5 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2420) ?
	       wdata32__h27246[25] :
	       _dfoo296 ;
  assign _dfoo366 =
	     (source_id__h66137 == 10'd4 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2420) ?
	       wdata32__h27246[25] :
	       _dfoo298 ;
  assign _dfoo368 =
	     (source_id__h66137 == 10'd3 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2420) ?
	       wdata32__h27246[25] :
	       _dfoo300 ;
  assign _dfoo37 =
	     source_id__h73617 == 10'd15 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2725 ||
	     source_id__h75113 == 10'd15 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2786 ;
  assign _dfoo370 =
	     (source_id__h66137 == 10'd2 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2420) ?
	       wdata32__h27246[25] :
	       _dfoo302 ;
  assign _dfoo372 =
	     (source_id__h66137 == 10'd1 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2420) ?
	       wdata32__h27246[25] :
	       _dfoo304 ;
  assign _dfoo374 =
	     (source_id__h66137 == 10'd0 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2420) ?
	       wdata32__h27246[25] :
	       _dfoo306 ;
  assign _dfoo376 =
	     (source_id__h66137 == 10'd16 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2420) ?
	       wdata32__h27246[25] :
	       _dfoo308 ;
  assign _dfoo378 =
	     (source_id__h66137 == 10'd15 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2420) ?
	       wdata32__h27246[25] :
	       _dfoo310 ;
  assign _dfoo38 =
	     (source_id__h73617 == 10'd15 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2725) ?
	       wdata32__h27246[30] :
	       wdata32__h27246[31] ;
  assign _dfoo380 =
	     (source_id__h66137 == 10'd14 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2420) ?
	       wdata32__h27246[25] :
	       _dfoo312 ;
  assign _dfoo382 =
	     (source_id__h66137 == 10'd13 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2420) ?
	       wdata32__h27246[25] :
	       _dfoo314 ;
  assign _dfoo384 =
	     (source_id__h66137 == 10'd12 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2420) ?
	       wdata32__h27246[25] :
	       _dfoo316 ;
  assign _dfoo386 =
	     (source_id__h66137 == 10'd11 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2420) ?
	       wdata32__h27246[25] :
	       _dfoo318 ;
  assign _dfoo388 =
	     (source_id__h66137 == 10'd10 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2420) ?
	       wdata32__h27246[25] :
	       _dfoo320 ;
  assign _dfoo39 =
	     source_id__h73617 == 10'd14 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2725 ||
	     source_id__h75113 == 10'd14 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2786 ;
  assign _dfoo390 =
	     (source_id__h66137 == 10'd9 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2420) ?
	       wdata32__h27246[25] :
	       _dfoo322 ;
  assign _dfoo392 =
	     (source_id__h66137 == 10'd8 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2420) ?
	       wdata32__h27246[25] :
	       _dfoo324 ;
  assign _dfoo394 =
	     (source_id__h66137 == 10'd7 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2420) ?
	       wdata32__h27246[25] :
	       _dfoo326 ;
  assign _dfoo396 =
	     (source_id__h66137 == 10'd6 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2420) ?
	       wdata32__h27246[25] :
	       _dfoo328 ;
  assign _dfoo398 =
	     (source_id__h66137 == 10'd5 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2420) ?
	       wdata32__h27246[25] :
	       _dfoo330 ;
  assign _dfoo4 =
	     (source_id__h73617 == 10'd15 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2725) ?
	       wdata32__h27246[30] :
	       wdata32__h27246[31] ;
  assign _dfoo40 =
	     (source_id__h73617 == 10'd14 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2725) ?
	       wdata32__h27246[30] :
	       wdata32__h27246[31] ;
  assign _dfoo400 =
	     (source_id__h66137 == 10'd4 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2420) ?
	       wdata32__h27246[25] :
	       _dfoo332 ;
  assign _dfoo402 =
	     (source_id__h66137 == 10'd3 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2420) ?
	       wdata32__h27246[25] :
	       _dfoo334 ;
  assign _dfoo404 =
	     (source_id__h66137 == 10'd2 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2420) ?
	       wdata32__h27246[25] :
	       _dfoo336 ;
  assign _dfoo406 =
	     (source_id__h66137 == 10'd1 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2420) ?
	       wdata32__h27246[25] :
	       _dfoo338 ;
  assign _dfoo408 =
	     (source_id__h66137 == 10'd0 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2420) ?
	       wdata32__h27246[25] :
	       _dfoo340 ;
  assign _dfoo409 =
	     source_id__h64641 == 10'd16 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2359 ||
	     source_id__h66137 == 10'd16 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2420 ||
	     _dfoo273 ;
  assign _dfoo41 =
	     source_id__h73617 == 10'd13 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2725 ||
	     source_id__h75113 == 10'd13 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2786 ;
  assign _dfoo410 =
	     (source_id__h64641 == 10'd16 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2359) ?
	       wdata32__h27246[24] :
	       _dfoo342 ;
  assign _dfoo411 =
	     source_id__h64641 == 10'd15 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2359 ||
	     source_id__h66137 == 10'd15 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2420 ||
	     _dfoo275 ;
  assign _dfoo412 =
	     (source_id__h64641 == 10'd15 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2359) ?
	       wdata32__h27246[24] :
	       _dfoo344 ;
  assign _dfoo413 =
	     source_id__h64641 == 10'd14 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2359 ||
	     source_id__h66137 == 10'd14 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2420 ||
	     _dfoo277 ;
  assign _dfoo414 =
	     (source_id__h64641 == 10'd14 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2359) ?
	       wdata32__h27246[24] :
	       _dfoo346 ;
  assign _dfoo415 =
	     source_id__h64641 == 10'd13 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2359 ||
	     source_id__h66137 == 10'd13 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2420 ||
	     _dfoo279 ;
  assign _dfoo416 =
	     (source_id__h64641 == 10'd13 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2359) ?
	       wdata32__h27246[24] :
	       _dfoo348 ;
  assign _dfoo417 =
	     source_id__h64641 == 10'd12 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2359 ||
	     source_id__h66137 == 10'd12 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2420 ||
	     _dfoo281 ;
  assign _dfoo418 =
	     (source_id__h64641 == 10'd12 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2359) ?
	       wdata32__h27246[24] :
	       _dfoo350 ;
  assign _dfoo419 =
	     source_id__h64641 == 10'd11 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2359 ||
	     source_id__h66137 == 10'd11 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2420 ||
	     _dfoo283 ;
  assign _dfoo42 =
	     (source_id__h73617 == 10'd13 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2725) ?
	       wdata32__h27246[30] :
	       wdata32__h27246[31] ;
  assign _dfoo420 =
	     (source_id__h64641 == 10'd11 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2359) ?
	       wdata32__h27246[24] :
	       _dfoo352 ;
  assign _dfoo421 =
	     source_id__h64641 == 10'd10 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2359 ||
	     source_id__h66137 == 10'd10 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2420 ||
	     _dfoo285 ;
  assign _dfoo422 =
	     (source_id__h64641 == 10'd10 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2359) ?
	       wdata32__h27246[24] :
	       _dfoo354 ;
  assign _dfoo423 =
	     source_id__h64641 == 10'd9 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2359 ||
	     source_id__h66137 == 10'd9 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2420 ||
	     _dfoo287 ;
  assign _dfoo424 =
	     (source_id__h64641 == 10'd9 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2359) ?
	       wdata32__h27246[24] :
	       _dfoo356 ;
  assign _dfoo425 =
	     source_id__h64641 == 10'd8 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2359 ||
	     source_id__h66137 == 10'd8 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2420 ||
	     _dfoo289 ;
  assign _dfoo426 =
	     (source_id__h64641 == 10'd8 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2359) ?
	       wdata32__h27246[24] :
	       _dfoo358 ;
  assign _dfoo427 =
	     source_id__h64641 == 10'd7 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2359 ||
	     source_id__h66137 == 10'd7 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2420 ||
	     _dfoo291 ;
  assign _dfoo428 =
	     (source_id__h64641 == 10'd7 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2359) ?
	       wdata32__h27246[24] :
	       _dfoo360 ;
  assign _dfoo429 =
	     source_id__h64641 == 10'd6 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2359 ||
	     source_id__h66137 == 10'd6 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2420 ||
	     _dfoo293 ;
  assign _dfoo43 =
	     source_id__h73617 == 10'd12 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2725 ||
	     source_id__h75113 == 10'd12 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2786 ;
  assign _dfoo430 =
	     (source_id__h64641 == 10'd6 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2359) ?
	       wdata32__h27246[24] :
	       _dfoo362 ;
  assign _dfoo431 =
	     source_id__h64641 == 10'd5 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2359 ||
	     source_id__h66137 == 10'd5 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2420 ||
	     _dfoo295 ;
  assign _dfoo432 =
	     (source_id__h64641 == 10'd5 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2359) ?
	       wdata32__h27246[24] :
	       _dfoo364 ;
  assign _dfoo433 =
	     source_id__h64641 == 10'd4 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2359 ||
	     source_id__h66137 == 10'd4 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2420 ||
	     _dfoo297 ;
  assign _dfoo434 =
	     (source_id__h64641 == 10'd4 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2359) ?
	       wdata32__h27246[24] :
	       _dfoo366 ;
  assign _dfoo435 =
	     source_id__h64641 == 10'd3 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2359 ||
	     source_id__h66137 == 10'd3 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2420 ||
	     _dfoo299 ;
  assign _dfoo436 =
	     (source_id__h64641 == 10'd3 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2359) ?
	       wdata32__h27246[24] :
	       _dfoo368 ;
  assign _dfoo437 =
	     source_id__h64641 == 10'd2 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2359 ||
	     source_id__h66137 == 10'd2 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2420 ||
	     _dfoo301 ;
  assign _dfoo438 =
	     (source_id__h64641 == 10'd2 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2359) ?
	       wdata32__h27246[24] :
	       _dfoo370 ;
  assign _dfoo439 =
	     source_id__h64641 == 10'd1 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2359 ||
	     source_id__h66137 == 10'd1 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2420 ||
	     _dfoo303 ;
  assign _dfoo44 =
	     (source_id__h73617 == 10'd12 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2725) ?
	       wdata32__h27246[30] :
	       wdata32__h27246[31] ;
  assign _dfoo440 =
	     (source_id__h64641 == 10'd1 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2359) ?
	       wdata32__h27246[24] :
	       _dfoo372 ;
  assign _dfoo441 =
	     source_id__h64641 == 10'd0 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2359 ||
	     source_id__h66137 == 10'd0 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2420 ||
	     _dfoo305 ;
  assign _dfoo442 =
	     (source_id__h64641 == 10'd0 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2359) ?
	       wdata32__h27246[24] :
	       _dfoo374 ;
  assign _dfoo443 =
	     source_id__h64641 == 10'd16 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2359 ||
	     source_id__h66137 == 10'd16 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2420 ||
	     _dfoo307 ;
  assign _dfoo444 =
	     (source_id__h64641 == 10'd16 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2359) ?
	       wdata32__h27246[24] :
	       _dfoo376 ;
  assign _dfoo445 =
	     source_id__h64641 == 10'd15 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2359 ||
	     source_id__h66137 == 10'd15 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2420 ||
	     _dfoo309 ;
  assign _dfoo446 =
	     (source_id__h64641 == 10'd15 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2359) ?
	       wdata32__h27246[24] :
	       _dfoo378 ;
  assign _dfoo447 =
	     source_id__h64641 == 10'd14 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2359 ||
	     source_id__h66137 == 10'd14 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2420 ||
	     _dfoo311 ;
  assign _dfoo448 =
	     (source_id__h64641 == 10'd14 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2359) ?
	       wdata32__h27246[24] :
	       _dfoo380 ;
  assign _dfoo449 =
	     source_id__h64641 == 10'd13 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2359 ||
	     source_id__h66137 == 10'd13 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2420 ||
	     _dfoo313 ;
  assign _dfoo45 =
	     source_id__h73617 == 10'd11 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2725 ||
	     source_id__h75113 == 10'd11 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2786 ;
  assign _dfoo450 =
	     (source_id__h64641 == 10'd13 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2359) ?
	       wdata32__h27246[24] :
	       _dfoo382 ;
  assign _dfoo451 =
	     source_id__h64641 == 10'd12 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2359 ||
	     source_id__h66137 == 10'd12 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2420 ||
	     _dfoo315 ;
  assign _dfoo452 =
	     (source_id__h64641 == 10'd12 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2359) ?
	       wdata32__h27246[24] :
	       _dfoo384 ;
  assign _dfoo453 =
	     source_id__h64641 == 10'd11 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2359 ||
	     source_id__h66137 == 10'd11 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2420 ||
	     _dfoo317 ;
  assign _dfoo454 =
	     (source_id__h64641 == 10'd11 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2359) ?
	       wdata32__h27246[24] :
	       _dfoo386 ;
  assign _dfoo455 =
	     source_id__h64641 == 10'd10 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2359 ||
	     source_id__h66137 == 10'd10 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2420 ||
	     _dfoo319 ;
  assign _dfoo456 =
	     (source_id__h64641 == 10'd10 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2359) ?
	       wdata32__h27246[24] :
	       _dfoo388 ;
  assign _dfoo457 =
	     source_id__h64641 == 10'd9 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2359 ||
	     source_id__h66137 == 10'd9 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2420 ||
	     _dfoo321 ;
  assign _dfoo458 =
	     (source_id__h64641 == 10'd9 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2359) ?
	       wdata32__h27246[24] :
	       _dfoo390 ;
  assign _dfoo459 =
	     source_id__h64641 == 10'd8 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2359 ||
	     source_id__h66137 == 10'd8 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2420 ||
	     _dfoo323 ;
  assign _dfoo46 =
	     (source_id__h73617 == 10'd11 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2725) ?
	       wdata32__h27246[30] :
	       wdata32__h27246[31] ;
  assign _dfoo460 =
	     (source_id__h64641 == 10'd8 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2359) ?
	       wdata32__h27246[24] :
	       _dfoo392 ;
  assign _dfoo461 =
	     source_id__h64641 == 10'd7 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2359 ||
	     source_id__h66137 == 10'd7 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2420 ||
	     _dfoo325 ;
  assign _dfoo462 =
	     (source_id__h64641 == 10'd7 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2359) ?
	       wdata32__h27246[24] :
	       _dfoo394 ;
  assign _dfoo463 =
	     source_id__h64641 == 10'd6 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2359 ||
	     source_id__h66137 == 10'd6 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2420 ||
	     _dfoo327 ;
  assign _dfoo464 =
	     (source_id__h64641 == 10'd6 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2359) ?
	       wdata32__h27246[24] :
	       _dfoo396 ;
  assign _dfoo465 =
	     source_id__h64641 == 10'd5 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2359 ||
	     source_id__h66137 == 10'd5 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2420 ||
	     _dfoo329 ;
  assign _dfoo466 =
	     (source_id__h64641 == 10'd5 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2359) ?
	       wdata32__h27246[24] :
	       _dfoo398 ;
  assign _dfoo467 =
	     source_id__h64641 == 10'd4 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2359 ||
	     source_id__h66137 == 10'd4 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2420 ||
	     _dfoo331 ;
  assign _dfoo468 =
	     (source_id__h64641 == 10'd4 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2359) ?
	       wdata32__h27246[24] :
	       _dfoo400 ;
  assign _dfoo469 =
	     source_id__h64641 == 10'd3 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2359 ||
	     source_id__h66137 == 10'd3 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2420 ||
	     _dfoo333 ;
  assign _dfoo47 =
	     source_id__h73617 == 10'd10 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2725 ||
	     source_id__h75113 == 10'd10 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2786 ;
  assign _dfoo470 =
	     (source_id__h64641 == 10'd3 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2359) ?
	       wdata32__h27246[24] :
	       _dfoo402 ;
  assign _dfoo471 =
	     source_id__h64641 == 10'd2 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2359 ||
	     source_id__h66137 == 10'd2 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2420 ||
	     _dfoo335 ;
  assign _dfoo472 =
	     (source_id__h64641 == 10'd2 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2359) ?
	       wdata32__h27246[24] :
	       _dfoo404 ;
  assign _dfoo473 =
	     source_id__h64641 == 10'd1 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2359 ||
	     source_id__h66137 == 10'd1 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2420 ||
	     _dfoo337 ;
  assign _dfoo474 =
	     (source_id__h64641 == 10'd1 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2359) ?
	       wdata32__h27246[24] :
	       _dfoo406 ;
  assign _dfoo475 =
	     source_id__h64641 == 10'd0 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2359 ||
	     source_id__h66137 == 10'd0 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2420 ||
	     _dfoo339 ;
  assign _dfoo476 =
	     (source_id__h64641 == 10'd0 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2359) ?
	       wdata32__h27246[24] :
	       _dfoo408 ;
  assign _dfoo478 =
	     (source_id__h63145 == 10'd16 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2298) ?
	       wdata32__h27246[23] :
	       _dfoo410 ;
  assign _dfoo48 =
	     (source_id__h73617 == 10'd10 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2725) ?
	       wdata32__h27246[30] :
	       wdata32__h27246[31] ;
  assign _dfoo480 =
	     (source_id__h63145 == 10'd15 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2298) ?
	       wdata32__h27246[23] :
	       _dfoo412 ;
  assign _dfoo482 =
	     (source_id__h63145 == 10'd14 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2298) ?
	       wdata32__h27246[23] :
	       _dfoo414 ;
  assign _dfoo484 =
	     (source_id__h63145 == 10'd13 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2298) ?
	       wdata32__h27246[23] :
	       _dfoo416 ;
  assign _dfoo486 =
	     (source_id__h63145 == 10'd12 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2298) ?
	       wdata32__h27246[23] :
	       _dfoo418 ;
  assign _dfoo488 =
	     (source_id__h63145 == 10'd11 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2298) ?
	       wdata32__h27246[23] :
	       _dfoo420 ;
  assign _dfoo49 =
	     source_id__h73617 == 10'd9 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2725 ||
	     source_id__h75113 == 10'd9 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2786 ;
  assign _dfoo490 =
	     (source_id__h63145 == 10'd10 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2298) ?
	       wdata32__h27246[23] :
	       _dfoo422 ;
  assign _dfoo492 =
	     (source_id__h63145 == 10'd9 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2298) ?
	       wdata32__h27246[23] :
	       _dfoo424 ;
  assign _dfoo494 =
	     (source_id__h63145 == 10'd8 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2298) ?
	       wdata32__h27246[23] :
	       _dfoo426 ;
  assign _dfoo496 =
	     (source_id__h63145 == 10'd7 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2298) ?
	       wdata32__h27246[23] :
	       _dfoo428 ;
  assign _dfoo498 =
	     (source_id__h63145 == 10'd6 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2298) ?
	       wdata32__h27246[23] :
	       _dfoo430 ;
  assign _dfoo5 =
	     source_id__h73617 == 10'd14 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2725 ||
	     source_id__h75113 == 10'd14 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2786 ;
  assign _dfoo50 =
	     (source_id__h73617 == 10'd9 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2725) ?
	       wdata32__h27246[30] :
	       wdata32__h27246[31] ;
  assign _dfoo500 =
	     (source_id__h63145 == 10'd5 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2298) ?
	       wdata32__h27246[23] :
	       _dfoo432 ;
  assign _dfoo502 =
	     (source_id__h63145 == 10'd4 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2298) ?
	       wdata32__h27246[23] :
	       _dfoo434 ;
  assign _dfoo504 =
	     (source_id__h63145 == 10'd3 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2298) ?
	       wdata32__h27246[23] :
	       _dfoo436 ;
  assign _dfoo506 =
	     (source_id__h63145 == 10'd2 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2298) ?
	       wdata32__h27246[23] :
	       _dfoo438 ;
  assign _dfoo508 =
	     (source_id__h63145 == 10'd1 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2298) ?
	       wdata32__h27246[23] :
	       _dfoo440 ;
  assign _dfoo51 =
	     source_id__h73617 == 10'd8 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2725 ||
	     source_id__h75113 == 10'd8 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2786 ;
  assign _dfoo510 =
	     (source_id__h63145 == 10'd0 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2298) ?
	       wdata32__h27246[23] :
	       _dfoo442 ;
  assign _dfoo512 =
	     (source_id__h63145 == 10'd16 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2298) ?
	       wdata32__h27246[23] :
	       _dfoo444 ;
  assign _dfoo514 =
	     (source_id__h63145 == 10'd15 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2298) ?
	       wdata32__h27246[23] :
	       _dfoo446 ;
  assign _dfoo516 =
	     (source_id__h63145 == 10'd14 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2298) ?
	       wdata32__h27246[23] :
	       _dfoo448 ;
  assign _dfoo518 =
	     (source_id__h63145 == 10'd13 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2298) ?
	       wdata32__h27246[23] :
	       _dfoo450 ;
  assign _dfoo52 =
	     (source_id__h73617 == 10'd8 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2725) ?
	       wdata32__h27246[30] :
	       wdata32__h27246[31] ;
  assign _dfoo520 =
	     (source_id__h63145 == 10'd12 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2298) ?
	       wdata32__h27246[23] :
	       _dfoo452 ;
  assign _dfoo522 =
	     (source_id__h63145 == 10'd11 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2298) ?
	       wdata32__h27246[23] :
	       _dfoo454 ;
  assign _dfoo524 =
	     (source_id__h63145 == 10'd10 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2298) ?
	       wdata32__h27246[23] :
	       _dfoo456 ;
  assign _dfoo526 =
	     (source_id__h63145 == 10'd9 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2298) ?
	       wdata32__h27246[23] :
	       _dfoo458 ;
  assign _dfoo528 =
	     (source_id__h63145 == 10'd8 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2298) ?
	       wdata32__h27246[23] :
	       _dfoo460 ;
  assign _dfoo53 =
	     source_id__h73617 == 10'd7 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2725 ||
	     source_id__h75113 == 10'd7 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2786 ;
  assign _dfoo530 =
	     (source_id__h63145 == 10'd7 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2298) ?
	       wdata32__h27246[23] :
	       _dfoo462 ;
  assign _dfoo532 =
	     (source_id__h63145 == 10'd6 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2298) ?
	       wdata32__h27246[23] :
	       _dfoo464 ;
  assign _dfoo534 =
	     (source_id__h63145 == 10'd5 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2298) ?
	       wdata32__h27246[23] :
	       _dfoo466 ;
  assign _dfoo536 =
	     (source_id__h63145 == 10'd4 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2298) ?
	       wdata32__h27246[23] :
	       _dfoo468 ;
  assign _dfoo538 =
	     (source_id__h63145 == 10'd3 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2298) ?
	       wdata32__h27246[23] :
	       _dfoo470 ;
  assign _dfoo54 =
	     (source_id__h73617 == 10'd7 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2725) ?
	       wdata32__h27246[30] :
	       wdata32__h27246[31] ;
  assign _dfoo540 =
	     (source_id__h63145 == 10'd2 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2298) ?
	       wdata32__h27246[23] :
	       _dfoo472 ;
  assign _dfoo542 =
	     (source_id__h63145 == 10'd1 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2298) ?
	       wdata32__h27246[23] :
	       _dfoo474 ;
  assign _dfoo544 =
	     (source_id__h63145 == 10'd0 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2298) ?
	       wdata32__h27246[23] :
	       _dfoo476 ;
  assign _dfoo545 =
	     source_id__h61649 == 10'd16 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2237 ||
	     source_id__h63145 == 10'd16 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2298 ||
	     _dfoo409 ;
  assign _dfoo546 =
	     (source_id__h61649 == 10'd16 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2237) ?
	       wdata32__h27246[22] :
	       _dfoo478 ;
  assign _dfoo547 =
	     source_id__h61649 == 10'd15 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2237 ||
	     source_id__h63145 == 10'd15 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2298 ||
	     _dfoo411 ;
  assign _dfoo548 =
	     (source_id__h61649 == 10'd15 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2237) ?
	       wdata32__h27246[22] :
	       _dfoo480 ;
  assign _dfoo549 =
	     source_id__h61649 == 10'd14 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2237 ||
	     source_id__h63145 == 10'd14 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2298 ||
	     _dfoo413 ;
  assign _dfoo55 =
	     source_id__h73617 == 10'd6 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2725 ||
	     source_id__h75113 == 10'd6 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2786 ;
  assign _dfoo550 =
	     (source_id__h61649 == 10'd14 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2237) ?
	       wdata32__h27246[22] :
	       _dfoo482 ;
  assign _dfoo551 =
	     source_id__h61649 == 10'd13 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2237 ||
	     source_id__h63145 == 10'd13 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2298 ||
	     _dfoo415 ;
  assign _dfoo552 =
	     (source_id__h61649 == 10'd13 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2237) ?
	       wdata32__h27246[22] :
	       _dfoo484 ;
  assign _dfoo553 =
	     source_id__h61649 == 10'd12 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2237 ||
	     source_id__h63145 == 10'd12 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2298 ||
	     _dfoo417 ;
  assign _dfoo554 =
	     (source_id__h61649 == 10'd12 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2237) ?
	       wdata32__h27246[22] :
	       _dfoo486 ;
  assign _dfoo555 =
	     source_id__h61649 == 10'd11 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2237 ||
	     source_id__h63145 == 10'd11 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2298 ||
	     _dfoo419 ;
  assign _dfoo556 =
	     (source_id__h61649 == 10'd11 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2237) ?
	       wdata32__h27246[22] :
	       _dfoo488 ;
  assign _dfoo557 =
	     source_id__h61649 == 10'd10 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2237 ||
	     source_id__h63145 == 10'd10 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2298 ||
	     _dfoo421 ;
  assign _dfoo558 =
	     (source_id__h61649 == 10'd10 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2237) ?
	       wdata32__h27246[22] :
	       _dfoo490 ;
  assign _dfoo559 =
	     source_id__h61649 == 10'd9 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2237 ||
	     source_id__h63145 == 10'd9 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2298 ||
	     _dfoo423 ;
  assign _dfoo56 =
	     (source_id__h73617 == 10'd6 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2725) ?
	       wdata32__h27246[30] :
	       wdata32__h27246[31] ;
  assign _dfoo560 =
	     (source_id__h61649 == 10'd9 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2237) ?
	       wdata32__h27246[22] :
	       _dfoo492 ;
  assign _dfoo561 =
	     source_id__h61649 == 10'd8 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2237 ||
	     source_id__h63145 == 10'd8 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2298 ||
	     _dfoo425 ;
  assign _dfoo562 =
	     (source_id__h61649 == 10'd8 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2237) ?
	       wdata32__h27246[22] :
	       _dfoo494 ;
  assign _dfoo563 =
	     source_id__h61649 == 10'd7 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2237 ||
	     source_id__h63145 == 10'd7 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2298 ||
	     _dfoo427 ;
  assign _dfoo564 =
	     (source_id__h61649 == 10'd7 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2237) ?
	       wdata32__h27246[22] :
	       _dfoo496 ;
  assign _dfoo565 =
	     source_id__h61649 == 10'd6 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2237 ||
	     source_id__h63145 == 10'd6 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2298 ||
	     _dfoo429 ;
  assign _dfoo566 =
	     (source_id__h61649 == 10'd6 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2237) ?
	       wdata32__h27246[22] :
	       _dfoo498 ;
  assign _dfoo567 =
	     source_id__h61649 == 10'd5 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2237 ||
	     source_id__h63145 == 10'd5 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2298 ||
	     _dfoo431 ;
  assign _dfoo568 =
	     (source_id__h61649 == 10'd5 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2237) ?
	       wdata32__h27246[22] :
	       _dfoo500 ;
  assign _dfoo569 =
	     source_id__h61649 == 10'd4 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2237 ||
	     source_id__h63145 == 10'd4 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2298 ||
	     _dfoo433 ;
  assign _dfoo57 =
	     source_id__h73617 == 10'd5 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2725 ||
	     source_id__h75113 == 10'd5 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2786 ;
  assign _dfoo570 =
	     (source_id__h61649 == 10'd4 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2237) ?
	       wdata32__h27246[22] :
	       _dfoo502 ;
  assign _dfoo571 =
	     source_id__h61649 == 10'd3 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2237 ||
	     source_id__h63145 == 10'd3 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2298 ||
	     _dfoo435 ;
  assign _dfoo572 =
	     (source_id__h61649 == 10'd3 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2237) ?
	       wdata32__h27246[22] :
	       _dfoo504 ;
  assign _dfoo573 =
	     source_id__h61649 == 10'd2 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2237 ||
	     source_id__h63145 == 10'd2 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2298 ||
	     _dfoo437 ;
  assign _dfoo574 =
	     (source_id__h61649 == 10'd2 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2237) ?
	       wdata32__h27246[22] :
	       _dfoo506 ;
  assign _dfoo575 =
	     source_id__h61649 == 10'd1 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2237 ||
	     source_id__h63145 == 10'd1 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2298 ||
	     _dfoo439 ;
  assign _dfoo576 =
	     (source_id__h61649 == 10'd1 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2237) ?
	       wdata32__h27246[22] :
	       _dfoo508 ;
  assign _dfoo577 =
	     source_id__h61649 == 10'd0 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2237 ||
	     source_id__h63145 == 10'd0 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2298 ||
	     _dfoo441 ;
  assign _dfoo578 =
	     (source_id__h61649 == 10'd0 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2237) ?
	       wdata32__h27246[22] :
	       _dfoo510 ;
  assign _dfoo579 =
	     source_id__h61649 == 10'd16 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2237 ||
	     source_id__h63145 == 10'd16 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2298 ||
	     _dfoo443 ;
  assign _dfoo58 =
	     (source_id__h73617 == 10'd5 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2725) ?
	       wdata32__h27246[30] :
	       wdata32__h27246[31] ;
  assign _dfoo580 =
	     (source_id__h61649 == 10'd16 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2237) ?
	       wdata32__h27246[22] :
	       _dfoo512 ;
  assign _dfoo581 =
	     source_id__h61649 == 10'd15 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2237 ||
	     source_id__h63145 == 10'd15 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2298 ||
	     _dfoo445 ;
  assign _dfoo582 =
	     (source_id__h61649 == 10'd15 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2237) ?
	       wdata32__h27246[22] :
	       _dfoo514 ;
  assign _dfoo583 =
	     source_id__h61649 == 10'd14 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2237 ||
	     source_id__h63145 == 10'd14 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2298 ||
	     _dfoo447 ;
  assign _dfoo584 =
	     (source_id__h61649 == 10'd14 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2237) ?
	       wdata32__h27246[22] :
	       _dfoo516 ;
  assign _dfoo585 =
	     source_id__h61649 == 10'd13 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2237 ||
	     source_id__h63145 == 10'd13 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2298 ||
	     _dfoo449 ;
  assign _dfoo586 =
	     (source_id__h61649 == 10'd13 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2237) ?
	       wdata32__h27246[22] :
	       _dfoo518 ;
  assign _dfoo587 =
	     source_id__h61649 == 10'd12 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2237 ||
	     source_id__h63145 == 10'd12 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2298 ||
	     _dfoo451 ;
  assign _dfoo588 =
	     (source_id__h61649 == 10'd12 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2237) ?
	       wdata32__h27246[22] :
	       _dfoo520 ;
  assign _dfoo589 =
	     source_id__h61649 == 10'd11 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2237 ||
	     source_id__h63145 == 10'd11 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2298 ||
	     _dfoo453 ;
  assign _dfoo59 =
	     source_id__h73617 == 10'd4 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2725 ||
	     source_id__h75113 == 10'd4 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2786 ;
  assign _dfoo590 =
	     (source_id__h61649 == 10'd11 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2237) ?
	       wdata32__h27246[22] :
	       _dfoo522 ;
  assign _dfoo591 =
	     source_id__h61649 == 10'd10 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2237 ||
	     source_id__h63145 == 10'd10 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2298 ||
	     _dfoo455 ;
  assign _dfoo592 =
	     (source_id__h61649 == 10'd10 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2237) ?
	       wdata32__h27246[22] :
	       _dfoo524 ;
  assign _dfoo593 =
	     source_id__h61649 == 10'd9 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2237 ||
	     source_id__h63145 == 10'd9 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2298 ||
	     _dfoo457 ;
  assign _dfoo594 =
	     (source_id__h61649 == 10'd9 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2237) ?
	       wdata32__h27246[22] :
	       _dfoo526 ;
  assign _dfoo595 =
	     source_id__h61649 == 10'd8 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2237 ||
	     source_id__h63145 == 10'd8 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2298 ||
	     _dfoo459 ;
  assign _dfoo596 =
	     (source_id__h61649 == 10'd8 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2237) ?
	       wdata32__h27246[22] :
	       _dfoo528 ;
  assign _dfoo597 =
	     source_id__h61649 == 10'd7 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2237 ||
	     source_id__h63145 == 10'd7 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2298 ||
	     _dfoo461 ;
  assign _dfoo598 =
	     (source_id__h61649 == 10'd7 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2237) ?
	       wdata32__h27246[22] :
	       _dfoo530 ;
  assign _dfoo599 =
	     source_id__h61649 == 10'd6 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2237 ||
	     source_id__h63145 == 10'd6 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2298 ||
	     _dfoo463 ;
  assign _dfoo6 =
	     (source_id__h73617 == 10'd14 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2725) ?
	       wdata32__h27246[30] :
	       wdata32__h27246[31] ;
  assign _dfoo60 =
	     (source_id__h73617 == 10'd4 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2725) ?
	       wdata32__h27246[30] :
	       wdata32__h27246[31] ;
  assign _dfoo600 =
	     (source_id__h61649 == 10'd6 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2237) ?
	       wdata32__h27246[22] :
	       _dfoo532 ;
  assign _dfoo601 =
	     source_id__h61649 == 10'd5 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2237 ||
	     source_id__h63145 == 10'd5 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2298 ||
	     _dfoo465 ;
  assign _dfoo602 =
	     (source_id__h61649 == 10'd5 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2237) ?
	       wdata32__h27246[22] :
	       _dfoo534 ;
  assign _dfoo603 =
	     source_id__h61649 == 10'd4 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2237 ||
	     source_id__h63145 == 10'd4 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2298 ||
	     _dfoo467 ;
  assign _dfoo604 =
	     (source_id__h61649 == 10'd4 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2237) ?
	       wdata32__h27246[22] :
	       _dfoo536 ;
  assign _dfoo605 =
	     source_id__h61649 == 10'd3 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2237 ||
	     source_id__h63145 == 10'd3 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2298 ||
	     _dfoo469 ;
  assign _dfoo606 =
	     (source_id__h61649 == 10'd3 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2237) ?
	       wdata32__h27246[22] :
	       _dfoo538 ;
  assign _dfoo607 =
	     source_id__h61649 == 10'd2 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2237 ||
	     source_id__h63145 == 10'd2 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2298 ||
	     _dfoo471 ;
  assign _dfoo608 =
	     (source_id__h61649 == 10'd2 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2237) ?
	       wdata32__h27246[22] :
	       _dfoo540 ;
  assign _dfoo609 =
	     source_id__h61649 == 10'd1 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2237 ||
	     source_id__h63145 == 10'd1 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2298 ||
	     _dfoo473 ;
  assign _dfoo61 =
	     source_id__h73617 == 10'd3 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2725 ||
	     source_id__h75113 == 10'd3 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2786 ;
  assign _dfoo610 =
	     (source_id__h61649 == 10'd1 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2237) ?
	       wdata32__h27246[22] :
	       _dfoo542 ;
  assign _dfoo611 =
	     source_id__h61649 == 10'd0 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2237 ||
	     source_id__h63145 == 10'd0 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2298 ||
	     _dfoo475 ;
  assign _dfoo612 =
	     (source_id__h61649 == 10'd0 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2237) ?
	       wdata32__h27246[22] :
	       _dfoo544 ;
  assign _dfoo614 =
	     (source_id__h60153 == 10'd16 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2176) ?
	       wdata32__h27246[21] :
	       _dfoo546 ;
  assign _dfoo616 =
	     (source_id__h60153 == 10'd15 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2176) ?
	       wdata32__h27246[21] :
	       _dfoo548 ;
  assign _dfoo618 =
	     (source_id__h60153 == 10'd14 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2176) ?
	       wdata32__h27246[21] :
	       _dfoo550 ;
  assign _dfoo62 =
	     (source_id__h73617 == 10'd3 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2725) ?
	       wdata32__h27246[30] :
	       wdata32__h27246[31] ;
  assign _dfoo620 =
	     (source_id__h60153 == 10'd13 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2176) ?
	       wdata32__h27246[21] :
	       _dfoo552 ;
  assign _dfoo622 =
	     (source_id__h60153 == 10'd12 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2176) ?
	       wdata32__h27246[21] :
	       _dfoo554 ;
  assign _dfoo624 =
	     (source_id__h60153 == 10'd11 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2176) ?
	       wdata32__h27246[21] :
	       _dfoo556 ;
  assign _dfoo626 =
	     (source_id__h60153 == 10'd10 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2176) ?
	       wdata32__h27246[21] :
	       _dfoo558 ;
  assign _dfoo628 =
	     (source_id__h60153 == 10'd9 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2176) ?
	       wdata32__h27246[21] :
	       _dfoo560 ;
  assign _dfoo63 =
	     source_id__h73617 == 10'd2 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2725 ||
	     source_id__h75113 == 10'd2 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2786 ;
  assign _dfoo630 =
	     (source_id__h60153 == 10'd8 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2176) ?
	       wdata32__h27246[21] :
	       _dfoo562 ;
  assign _dfoo632 =
	     (source_id__h60153 == 10'd7 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2176) ?
	       wdata32__h27246[21] :
	       _dfoo564 ;
  assign _dfoo634 =
	     (source_id__h60153 == 10'd6 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2176) ?
	       wdata32__h27246[21] :
	       _dfoo566 ;
  assign _dfoo636 =
	     (source_id__h60153 == 10'd5 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2176) ?
	       wdata32__h27246[21] :
	       _dfoo568 ;
  assign _dfoo638 =
	     (source_id__h60153 == 10'd4 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2176) ?
	       wdata32__h27246[21] :
	       _dfoo570 ;
  assign _dfoo64 =
	     (source_id__h73617 == 10'd2 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2725) ?
	       wdata32__h27246[30] :
	       wdata32__h27246[31] ;
  assign _dfoo640 =
	     (source_id__h60153 == 10'd3 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2176) ?
	       wdata32__h27246[21] :
	       _dfoo572 ;
  assign _dfoo642 =
	     (source_id__h60153 == 10'd2 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2176) ?
	       wdata32__h27246[21] :
	       _dfoo574 ;
  assign _dfoo644 =
	     (source_id__h60153 == 10'd1 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2176) ?
	       wdata32__h27246[21] :
	       _dfoo576 ;
  assign _dfoo646 =
	     (source_id__h60153 == 10'd0 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2176) ?
	       wdata32__h27246[21] :
	       _dfoo578 ;
  assign _dfoo648 =
	     (source_id__h60153 == 10'd16 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2176) ?
	       wdata32__h27246[21] :
	       _dfoo580 ;
  assign _dfoo65 =
	     source_id__h73617 == 10'd1 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2725 ||
	     source_id__h75113 == 10'd1 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2786 ;
  assign _dfoo650 =
	     (source_id__h60153 == 10'd15 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2176) ?
	       wdata32__h27246[21] :
	       _dfoo582 ;
  assign _dfoo652 =
	     (source_id__h60153 == 10'd14 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2176) ?
	       wdata32__h27246[21] :
	       _dfoo584 ;
  assign _dfoo654 =
	     (source_id__h60153 == 10'd13 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2176) ?
	       wdata32__h27246[21] :
	       _dfoo586 ;
  assign _dfoo656 =
	     (source_id__h60153 == 10'd12 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2176) ?
	       wdata32__h27246[21] :
	       _dfoo588 ;
  assign _dfoo658 =
	     (source_id__h60153 == 10'd11 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2176) ?
	       wdata32__h27246[21] :
	       _dfoo590 ;
  assign _dfoo66 =
	     (source_id__h73617 == 10'd1 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2725) ?
	       wdata32__h27246[30] :
	       wdata32__h27246[31] ;
  assign _dfoo660 =
	     (source_id__h60153 == 10'd10 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2176) ?
	       wdata32__h27246[21] :
	       _dfoo592 ;
  assign _dfoo662 =
	     (source_id__h60153 == 10'd9 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2176) ?
	       wdata32__h27246[21] :
	       _dfoo594 ;
  assign _dfoo664 =
	     (source_id__h60153 == 10'd8 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2176) ?
	       wdata32__h27246[21] :
	       _dfoo596 ;
  assign _dfoo666 =
	     (source_id__h60153 == 10'd7 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2176) ?
	       wdata32__h27246[21] :
	       _dfoo598 ;
  assign _dfoo668 =
	     (source_id__h60153 == 10'd6 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2176) ?
	       wdata32__h27246[21] :
	       _dfoo600 ;
  assign _dfoo67 =
	     source_id__h73617 == 10'd0 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2725 ||
	     source_id__h75113 == 10'd0 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2786 ;
  assign _dfoo670 =
	     (source_id__h60153 == 10'd5 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2176) ?
	       wdata32__h27246[21] :
	       _dfoo602 ;
  assign _dfoo672 =
	     (source_id__h60153 == 10'd4 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2176) ?
	       wdata32__h27246[21] :
	       _dfoo604 ;
  assign _dfoo674 =
	     (source_id__h60153 == 10'd3 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2176) ?
	       wdata32__h27246[21] :
	       _dfoo606 ;
  assign _dfoo676 =
	     (source_id__h60153 == 10'd2 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2176) ?
	       wdata32__h27246[21] :
	       _dfoo608 ;
  assign _dfoo678 =
	     (source_id__h60153 == 10'd1 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2176) ?
	       wdata32__h27246[21] :
	       _dfoo610 ;
  assign _dfoo68 =
	     (source_id__h73617 == 10'd0 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2725) ?
	       wdata32__h27246[30] :
	       wdata32__h27246[31] ;
  assign _dfoo680 =
	     (source_id__h60153 == 10'd0 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2176) ?
	       wdata32__h27246[21] :
	       _dfoo612 ;
  assign _dfoo681 =
	     source_id__h58657 == 10'd16 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2115 ||
	     source_id__h60153 == 10'd16 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2176 ||
	     _dfoo545 ;
  assign _dfoo682 =
	     (source_id__h58657 == 10'd16 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2115) ?
	       wdata32__h27246[20] :
	       _dfoo614 ;
  assign _dfoo683 =
	     source_id__h58657 == 10'd15 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2115 ||
	     source_id__h60153 == 10'd15 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2176 ||
	     _dfoo547 ;
  assign _dfoo684 =
	     (source_id__h58657 == 10'd15 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2115) ?
	       wdata32__h27246[20] :
	       _dfoo616 ;
  assign _dfoo685 =
	     source_id__h58657 == 10'd14 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2115 ||
	     source_id__h60153 == 10'd14 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2176 ||
	     _dfoo549 ;
  assign _dfoo686 =
	     (source_id__h58657 == 10'd14 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2115) ?
	       wdata32__h27246[20] :
	       _dfoo618 ;
  assign _dfoo687 =
	     source_id__h58657 == 10'd13 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2115 ||
	     source_id__h60153 == 10'd13 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2176 ||
	     _dfoo551 ;
  assign _dfoo688 =
	     (source_id__h58657 == 10'd13 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2115) ?
	       wdata32__h27246[20] :
	       _dfoo620 ;
  assign _dfoo689 =
	     source_id__h58657 == 10'd12 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2115 ||
	     source_id__h60153 == 10'd12 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2176 ||
	     _dfoo553 ;
  assign _dfoo690 =
	     (source_id__h58657 == 10'd12 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2115) ?
	       wdata32__h27246[20] :
	       _dfoo622 ;
  assign _dfoo691 =
	     source_id__h58657 == 10'd11 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2115 ||
	     source_id__h60153 == 10'd11 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2176 ||
	     _dfoo555 ;
  assign _dfoo692 =
	     (source_id__h58657 == 10'd11 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2115) ?
	       wdata32__h27246[20] :
	       _dfoo624 ;
  assign _dfoo693 =
	     source_id__h58657 == 10'd10 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2115 ||
	     source_id__h60153 == 10'd10 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2176 ||
	     _dfoo557 ;
  assign _dfoo694 =
	     (source_id__h58657 == 10'd10 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2115) ?
	       wdata32__h27246[20] :
	       _dfoo626 ;
  assign _dfoo695 =
	     source_id__h58657 == 10'd9 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2115 ||
	     source_id__h60153 == 10'd9 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2176 ||
	     _dfoo559 ;
  assign _dfoo696 =
	     (source_id__h58657 == 10'd9 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2115) ?
	       wdata32__h27246[20] :
	       _dfoo628 ;
  assign _dfoo697 =
	     source_id__h58657 == 10'd8 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2115 ||
	     source_id__h60153 == 10'd8 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2176 ||
	     _dfoo561 ;
  assign _dfoo698 =
	     (source_id__h58657 == 10'd8 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2115) ?
	       wdata32__h27246[20] :
	       _dfoo630 ;
  assign _dfoo699 =
	     source_id__h58657 == 10'd7 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2115 ||
	     source_id__h60153 == 10'd7 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2176 ||
	     _dfoo563 ;
  assign _dfoo7 =
	     source_id__h73617 == 10'd13 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2725 ||
	     source_id__h75113 == 10'd13 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2786 ;
  assign _dfoo70 =
	     (source_id__h72121 == 10'd16 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2664) ?
	       wdata32__h27246[29] :
	       _dfoo2 ;
  assign _dfoo700 =
	     (source_id__h58657 == 10'd7 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2115) ?
	       wdata32__h27246[20] :
	       _dfoo632 ;
  assign _dfoo701 =
	     source_id__h58657 == 10'd6 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2115 ||
	     source_id__h60153 == 10'd6 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2176 ||
	     _dfoo565 ;
  assign _dfoo702 =
	     (source_id__h58657 == 10'd6 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2115) ?
	       wdata32__h27246[20] :
	       _dfoo634 ;
  assign _dfoo703 =
	     source_id__h58657 == 10'd5 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2115 ||
	     source_id__h60153 == 10'd5 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2176 ||
	     _dfoo567 ;
  assign _dfoo704 =
	     (source_id__h58657 == 10'd5 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2115) ?
	       wdata32__h27246[20] :
	       _dfoo636 ;
  assign _dfoo705 =
	     source_id__h58657 == 10'd4 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2115 ||
	     source_id__h60153 == 10'd4 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2176 ||
	     _dfoo569 ;
  assign _dfoo706 =
	     (source_id__h58657 == 10'd4 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2115) ?
	       wdata32__h27246[20] :
	       _dfoo638 ;
  assign _dfoo707 =
	     source_id__h58657 == 10'd3 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2115 ||
	     source_id__h60153 == 10'd3 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2176 ||
	     _dfoo571 ;
  assign _dfoo708 =
	     (source_id__h58657 == 10'd3 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2115) ?
	       wdata32__h27246[20] :
	       _dfoo640 ;
  assign _dfoo709 =
	     source_id__h58657 == 10'd2 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2115 ||
	     source_id__h60153 == 10'd2 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2176 ||
	     _dfoo573 ;
  assign _dfoo710 =
	     (source_id__h58657 == 10'd2 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2115) ?
	       wdata32__h27246[20] :
	       _dfoo642 ;
  assign _dfoo711 =
	     source_id__h58657 == 10'd1 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2115 ||
	     source_id__h60153 == 10'd1 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2176 ||
	     _dfoo575 ;
  assign _dfoo712 =
	     (source_id__h58657 == 10'd1 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2115) ?
	       wdata32__h27246[20] :
	       _dfoo644 ;
  assign _dfoo713 =
	     source_id__h58657 == 10'd0 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2115 ||
	     source_id__h60153 == 10'd0 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2176 ||
	     _dfoo577 ;
  assign _dfoo714 =
	     (source_id__h58657 == 10'd0 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2115) ?
	       wdata32__h27246[20] :
	       _dfoo646 ;
  assign _dfoo715 =
	     source_id__h58657 == 10'd16 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2115 ||
	     source_id__h60153 == 10'd16 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2176 ||
	     _dfoo579 ;
  assign _dfoo716 =
	     (source_id__h58657 == 10'd16 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2115) ?
	       wdata32__h27246[20] :
	       _dfoo648 ;
  assign _dfoo717 =
	     source_id__h58657 == 10'd15 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2115 ||
	     source_id__h60153 == 10'd15 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2176 ||
	     _dfoo581 ;
  assign _dfoo718 =
	     (source_id__h58657 == 10'd15 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2115) ?
	       wdata32__h27246[20] :
	       _dfoo650 ;
  assign _dfoo719 =
	     source_id__h58657 == 10'd14 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2115 ||
	     source_id__h60153 == 10'd14 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2176 ||
	     _dfoo583 ;
  assign _dfoo72 =
	     (source_id__h72121 == 10'd15 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2664) ?
	       wdata32__h27246[29] :
	       _dfoo4 ;
  assign _dfoo720 =
	     (source_id__h58657 == 10'd14 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2115) ?
	       wdata32__h27246[20] :
	       _dfoo652 ;
  assign _dfoo721 =
	     source_id__h58657 == 10'd13 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2115 ||
	     source_id__h60153 == 10'd13 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2176 ||
	     _dfoo585 ;
  assign _dfoo722 =
	     (source_id__h58657 == 10'd13 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2115) ?
	       wdata32__h27246[20] :
	       _dfoo654 ;
  assign _dfoo723 =
	     source_id__h58657 == 10'd12 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2115 ||
	     source_id__h60153 == 10'd12 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2176 ||
	     _dfoo587 ;
  assign _dfoo724 =
	     (source_id__h58657 == 10'd12 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2115) ?
	       wdata32__h27246[20] :
	       _dfoo656 ;
  assign _dfoo725 =
	     source_id__h58657 == 10'd11 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2115 ||
	     source_id__h60153 == 10'd11 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2176 ||
	     _dfoo589 ;
  assign _dfoo726 =
	     (source_id__h58657 == 10'd11 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2115) ?
	       wdata32__h27246[20] :
	       _dfoo658 ;
  assign _dfoo727 =
	     source_id__h58657 == 10'd10 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2115 ||
	     source_id__h60153 == 10'd10 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2176 ||
	     _dfoo591 ;
  assign _dfoo728 =
	     (source_id__h58657 == 10'd10 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2115) ?
	       wdata32__h27246[20] :
	       _dfoo660 ;
  assign _dfoo729 =
	     source_id__h58657 == 10'd9 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2115 ||
	     source_id__h60153 == 10'd9 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2176 ||
	     _dfoo593 ;
  assign _dfoo730 =
	     (source_id__h58657 == 10'd9 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2115) ?
	       wdata32__h27246[20] :
	       _dfoo662 ;
  assign _dfoo731 =
	     source_id__h58657 == 10'd8 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2115 ||
	     source_id__h60153 == 10'd8 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2176 ||
	     _dfoo595 ;
  assign _dfoo732 =
	     (source_id__h58657 == 10'd8 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2115) ?
	       wdata32__h27246[20] :
	       _dfoo664 ;
  assign _dfoo733 =
	     source_id__h58657 == 10'd7 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2115 ||
	     source_id__h60153 == 10'd7 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2176 ||
	     _dfoo597 ;
  assign _dfoo734 =
	     (source_id__h58657 == 10'd7 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2115) ?
	       wdata32__h27246[20] :
	       _dfoo666 ;
  assign _dfoo735 =
	     source_id__h58657 == 10'd6 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2115 ||
	     source_id__h60153 == 10'd6 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2176 ||
	     _dfoo599 ;
  assign _dfoo736 =
	     (source_id__h58657 == 10'd6 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2115) ?
	       wdata32__h27246[20] :
	       _dfoo668 ;
  assign _dfoo737 =
	     source_id__h58657 == 10'd5 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2115 ||
	     source_id__h60153 == 10'd5 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2176 ||
	     _dfoo601 ;
  assign _dfoo738 =
	     (source_id__h58657 == 10'd5 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2115) ?
	       wdata32__h27246[20] :
	       _dfoo670 ;
  assign _dfoo739 =
	     source_id__h58657 == 10'd4 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2115 ||
	     source_id__h60153 == 10'd4 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2176 ||
	     _dfoo603 ;
  assign _dfoo74 =
	     (source_id__h72121 == 10'd14 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2664) ?
	       wdata32__h27246[29] :
	       _dfoo6 ;
  assign _dfoo740 =
	     (source_id__h58657 == 10'd4 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2115) ?
	       wdata32__h27246[20] :
	       _dfoo672 ;
  assign _dfoo741 =
	     source_id__h58657 == 10'd3 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2115 ||
	     source_id__h60153 == 10'd3 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2176 ||
	     _dfoo605 ;
  assign _dfoo742 =
	     (source_id__h58657 == 10'd3 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2115) ?
	       wdata32__h27246[20] :
	       _dfoo674 ;
  assign _dfoo743 =
	     source_id__h58657 == 10'd2 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2115 ||
	     source_id__h60153 == 10'd2 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2176 ||
	     _dfoo607 ;
  assign _dfoo744 =
	     (source_id__h58657 == 10'd2 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2115) ?
	       wdata32__h27246[20] :
	       _dfoo676 ;
  assign _dfoo745 =
	     source_id__h58657 == 10'd1 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2115 ||
	     source_id__h60153 == 10'd1 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2176 ||
	     _dfoo609 ;
  assign _dfoo746 =
	     (source_id__h58657 == 10'd1 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2115) ?
	       wdata32__h27246[20] :
	       _dfoo678 ;
  assign _dfoo747 =
	     source_id__h58657 == 10'd0 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2115 ||
	     source_id__h60153 == 10'd0 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2176 ||
	     _dfoo611 ;
  assign _dfoo748 =
	     (source_id__h58657 == 10'd0 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2115) ?
	       wdata32__h27246[20] :
	       _dfoo680 ;
  assign _dfoo750 =
	     (source_id__h57161 == 10'd16 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2054) ?
	       wdata32__h27246[19] :
	       _dfoo682 ;
  assign _dfoo752 =
	     (source_id__h57161 == 10'd15 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2054) ?
	       wdata32__h27246[19] :
	       _dfoo684 ;
  assign _dfoo754 =
	     (source_id__h57161 == 10'd14 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2054) ?
	       wdata32__h27246[19] :
	       _dfoo686 ;
  assign _dfoo756 =
	     (source_id__h57161 == 10'd13 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2054) ?
	       wdata32__h27246[19] :
	       _dfoo688 ;
  assign _dfoo758 =
	     (source_id__h57161 == 10'd12 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2054) ?
	       wdata32__h27246[19] :
	       _dfoo690 ;
  assign _dfoo76 =
	     (source_id__h72121 == 10'd13 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2664) ?
	       wdata32__h27246[29] :
	       _dfoo8 ;
  assign _dfoo760 =
	     (source_id__h57161 == 10'd11 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2054) ?
	       wdata32__h27246[19] :
	       _dfoo692 ;
  assign _dfoo762 =
	     (source_id__h57161 == 10'd10 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2054) ?
	       wdata32__h27246[19] :
	       _dfoo694 ;
  assign _dfoo764 =
	     (source_id__h57161 == 10'd9 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2054) ?
	       wdata32__h27246[19] :
	       _dfoo696 ;
  assign _dfoo766 =
	     (source_id__h57161 == 10'd8 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2054) ?
	       wdata32__h27246[19] :
	       _dfoo698 ;
  assign _dfoo768 =
	     (source_id__h57161 == 10'd7 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2054) ?
	       wdata32__h27246[19] :
	       _dfoo700 ;
  assign _dfoo770 =
	     (source_id__h57161 == 10'd6 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2054) ?
	       wdata32__h27246[19] :
	       _dfoo702 ;
  assign _dfoo772 =
	     (source_id__h57161 == 10'd5 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2054) ?
	       wdata32__h27246[19] :
	       _dfoo704 ;
  assign _dfoo774 =
	     (source_id__h57161 == 10'd4 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2054) ?
	       wdata32__h27246[19] :
	       _dfoo706 ;
  assign _dfoo776 =
	     (source_id__h57161 == 10'd3 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2054) ?
	       wdata32__h27246[19] :
	       _dfoo708 ;
  assign _dfoo778 =
	     (source_id__h57161 == 10'd2 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2054) ?
	       wdata32__h27246[19] :
	       _dfoo710 ;
  assign _dfoo78 =
	     (source_id__h72121 == 10'd12 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2664) ?
	       wdata32__h27246[29] :
	       _dfoo10 ;
  assign _dfoo780 =
	     (source_id__h57161 == 10'd1 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2054) ?
	       wdata32__h27246[19] :
	       _dfoo712 ;
  assign _dfoo782 =
	     (source_id__h57161 == 10'd0 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2054) ?
	       wdata32__h27246[19] :
	       _dfoo714 ;
  assign _dfoo784 =
	     (source_id__h57161 == 10'd16 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2054) ?
	       wdata32__h27246[19] :
	       _dfoo716 ;
  assign _dfoo786 =
	     (source_id__h57161 == 10'd15 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2054) ?
	       wdata32__h27246[19] :
	       _dfoo718 ;
  assign _dfoo788 =
	     (source_id__h57161 == 10'd14 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2054) ?
	       wdata32__h27246[19] :
	       _dfoo720 ;
  assign _dfoo790 =
	     (source_id__h57161 == 10'd13 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2054) ?
	       wdata32__h27246[19] :
	       _dfoo722 ;
  assign _dfoo792 =
	     (source_id__h57161 == 10'd12 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2054) ?
	       wdata32__h27246[19] :
	       _dfoo724 ;
  assign _dfoo794 =
	     (source_id__h57161 == 10'd11 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2054) ?
	       wdata32__h27246[19] :
	       _dfoo726 ;
  assign _dfoo796 =
	     (source_id__h57161 == 10'd10 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2054) ?
	       wdata32__h27246[19] :
	       _dfoo728 ;
  assign _dfoo798 =
	     (source_id__h57161 == 10'd9 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2054) ?
	       wdata32__h27246[19] :
	       _dfoo730 ;
  assign _dfoo8 =
	     (source_id__h73617 == 10'd13 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2725) ?
	       wdata32__h27246[30] :
	       wdata32__h27246[31] ;
  assign _dfoo80 =
	     (source_id__h72121 == 10'd11 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2664) ?
	       wdata32__h27246[29] :
	       _dfoo12 ;
  assign _dfoo800 =
	     (source_id__h57161 == 10'd8 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2054) ?
	       wdata32__h27246[19] :
	       _dfoo732 ;
  assign _dfoo802 =
	     (source_id__h57161 == 10'd7 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2054) ?
	       wdata32__h27246[19] :
	       _dfoo734 ;
  assign _dfoo804 =
	     (source_id__h57161 == 10'd6 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2054) ?
	       wdata32__h27246[19] :
	       _dfoo736 ;
  assign _dfoo806 =
	     (source_id__h57161 == 10'd5 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2054) ?
	       wdata32__h27246[19] :
	       _dfoo738 ;
  assign _dfoo808 =
	     (source_id__h57161 == 10'd4 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2054) ?
	       wdata32__h27246[19] :
	       _dfoo740 ;
  assign _dfoo810 =
	     (source_id__h57161 == 10'd3 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2054) ?
	       wdata32__h27246[19] :
	       _dfoo742 ;
  assign _dfoo812 =
	     (source_id__h57161 == 10'd2 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2054) ?
	       wdata32__h27246[19] :
	       _dfoo744 ;
  assign _dfoo814 =
	     (source_id__h57161 == 10'd1 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2054) ?
	       wdata32__h27246[19] :
	       _dfoo746 ;
  assign _dfoo816 =
	     (source_id__h57161 == 10'd0 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2054) ?
	       wdata32__h27246[19] :
	       _dfoo748 ;
  assign _dfoo817 =
	     source_id__h55665 == 10'd16 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1993 ||
	     source_id__h57161 == 10'd16 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2054 ||
	     _dfoo681 ;
  assign _dfoo818 =
	     (source_id__h55665 == 10'd16 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1993) ?
	       wdata32__h27246[18] :
	       _dfoo750 ;
  assign _dfoo819 =
	     source_id__h55665 == 10'd15 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1993 ||
	     source_id__h57161 == 10'd15 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2054 ||
	     _dfoo683 ;
  assign _dfoo82 =
	     (source_id__h72121 == 10'd10 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2664) ?
	       wdata32__h27246[29] :
	       _dfoo14 ;
  assign _dfoo820 =
	     (source_id__h55665 == 10'd15 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1993) ?
	       wdata32__h27246[18] :
	       _dfoo752 ;
  assign _dfoo821 =
	     source_id__h55665 == 10'd14 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1993 ||
	     source_id__h57161 == 10'd14 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2054 ||
	     _dfoo685 ;
  assign _dfoo822 =
	     (source_id__h55665 == 10'd14 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1993) ?
	       wdata32__h27246[18] :
	       _dfoo754 ;
  assign _dfoo823 =
	     source_id__h55665 == 10'd13 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1993 ||
	     source_id__h57161 == 10'd13 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2054 ||
	     _dfoo687 ;
  assign _dfoo824 =
	     (source_id__h55665 == 10'd13 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1993) ?
	       wdata32__h27246[18] :
	       _dfoo756 ;
  assign _dfoo825 =
	     source_id__h55665 == 10'd12 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1993 ||
	     source_id__h57161 == 10'd12 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2054 ||
	     _dfoo689 ;
  assign _dfoo826 =
	     (source_id__h55665 == 10'd12 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1993) ?
	       wdata32__h27246[18] :
	       _dfoo758 ;
  assign _dfoo827 =
	     source_id__h55665 == 10'd11 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1993 ||
	     source_id__h57161 == 10'd11 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2054 ||
	     _dfoo691 ;
  assign _dfoo828 =
	     (source_id__h55665 == 10'd11 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1993) ?
	       wdata32__h27246[18] :
	       _dfoo760 ;
  assign _dfoo829 =
	     source_id__h55665 == 10'd10 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1993 ||
	     source_id__h57161 == 10'd10 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2054 ||
	     _dfoo693 ;
  assign _dfoo830 =
	     (source_id__h55665 == 10'd10 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1993) ?
	       wdata32__h27246[18] :
	       _dfoo762 ;
  assign _dfoo831 =
	     source_id__h55665 == 10'd9 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1993 ||
	     source_id__h57161 == 10'd9 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2054 ||
	     _dfoo695 ;
  assign _dfoo832 =
	     (source_id__h55665 == 10'd9 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1993) ?
	       wdata32__h27246[18] :
	       _dfoo764 ;
  assign _dfoo833 =
	     source_id__h55665 == 10'd8 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1993 ||
	     source_id__h57161 == 10'd8 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2054 ||
	     _dfoo697 ;
  assign _dfoo834 =
	     (source_id__h55665 == 10'd8 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1993) ?
	       wdata32__h27246[18] :
	       _dfoo766 ;
  assign _dfoo835 =
	     source_id__h55665 == 10'd7 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1993 ||
	     source_id__h57161 == 10'd7 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2054 ||
	     _dfoo699 ;
  assign _dfoo836 =
	     (source_id__h55665 == 10'd7 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1993) ?
	       wdata32__h27246[18] :
	       _dfoo768 ;
  assign _dfoo837 =
	     source_id__h55665 == 10'd6 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1993 ||
	     source_id__h57161 == 10'd6 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2054 ||
	     _dfoo701 ;
  assign _dfoo838 =
	     (source_id__h55665 == 10'd6 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1993) ?
	       wdata32__h27246[18] :
	       _dfoo770 ;
  assign _dfoo839 =
	     source_id__h55665 == 10'd5 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1993 ||
	     source_id__h57161 == 10'd5 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2054 ||
	     _dfoo703 ;
  assign _dfoo84 =
	     (source_id__h72121 == 10'd9 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2664) ?
	       wdata32__h27246[29] :
	       _dfoo16 ;
  assign _dfoo840 =
	     (source_id__h55665 == 10'd5 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1993) ?
	       wdata32__h27246[18] :
	       _dfoo772 ;
  assign _dfoo841 =
	     source_id__h55665 == 10'd4 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1993 ||
	     source_id__h57161 == 10'd4 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2054 ||
	     _dfoo705 ;
  assign _dfoo842 =
	     (source_id__h55665 == 10'd4 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1993) ?
	       wdata32__h27246[18] :
	       _dfoo774 ;
  assign _dfoo843 =
	     source_id__h55665 == 10'd3 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1993 ||
	     source_id__h57161 == 10'd3 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2054 ||
	     _dfoo707 ;
  assign _dfoo844 =
	     (source_id__h55665 == 10'd3 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1993) ?
	       wdata32__h27246[18] :
	       _dfoo776 ;
  assign _dfoo845 =
	     source_id__h55665 == 10'd2 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1993 ||
	     source_id__h57161 == 10'd2 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2054 ||
	     _dfoo709 ;
  assign _dfoo846 =
	     (source_id__h55665 == 10'd2 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1993) ?
	       wdata32__h27246[18] :
	       _dfoo778 ;
  assign _dfoo847 =
	     source_id__h55665 == 10'd1 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1993 ||
	     source_id__h57161 == 10'd1 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2054 ||
	     _dfoo711 ;
  assign _dfoo848 =
	     (source_id__h55665 == 10'd1 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1993) ?
	       wdata32__h27246[18] :
	       _dfoo780 ;
  assign _dfoo849 =
	     source_id__h55665 == 10'd0 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1993 ||
	     source_id__h57161 == 10'd0 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2054 ||
	     _dfoo713 ;
  assign _dfoo850 =
	     (source_id__h55665 == 10'd0 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1993) ?
	       wdata32__h27246[18] :
	       _dfoo782 ;
  assign _dfoo851 =
	     source_id__h55665 == 10'd16 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1993 ||
	     source_id__h57161 == 10'd16 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2054 ||
	     _dfoo715 ;
  assign _dfoo852 =
	     (source_id__h55665 == 10'd16 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1993) ?
	       wdata32__h27246[18] :
	       _dfoo784 ;
  assign _dfoo853 =
	     source_id__h55665 == 10'd15 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1993 ||
	     source_id__h57161 == 10'd15 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2054 ||
	     _dfoo717 ;
  assign _dfoo854 =
	     (source_id__h55665 == 10'd15 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1993) ?
	       wdata32__h27246[18] :
	       _dfoo786 ;
  assign _dfoo855 =
	     source_id__h55665 == 10'd14 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1993 ||
	     source_id__h57161 == 10'd14 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2054 ||
	     _dfoo719 ;
  assign _dfoo856 =
	     (source_id__h55665 == 10'd14 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1993) ?
	       wdata32__h27246[18] :
	       _dfoo788 ;
  assign _dfoo857 =
	     source_id__h55665 == 10'd13 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1993 ||
	     source_id__h57161 == 10'd13 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2054 ||
	     _dfoo721 ;
  assign _dfoo858 =
	     (source_id__h55665 == 10'd13 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1993) ?
	       wdata32__h27246[18] :
	       _dfoo790 ;
  assign _dfoo859 =
	     source_id__h55665 == 10'd12 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1993 ||
	     source_id__h57161 == 10'd12 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2054 ||
	     _dfoo723 ;
  assign _dfoo86 =
	     (source_id__h72121 == 10'd8 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2664) ?
	       wdata32__h27246[29] :
	       _dfoo18 ;
  assign _dfoo860 =
	     (source_id__h55665 == 10'd12 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1993) ?
	       wdata32__h27246[18] :
	       _dfoo792 ;
  assign _dfoo861 =
	     source_id__h55665 == 10'd11 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1993 ||
	     source_id__h57161 == 10'd11 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2054 ||
	     _dfoo725 ;
  assign _dfoo862 =
	     (source_id__h55665 == 10'd11 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1993) ?
	       wdata32__h27246[18] :
	       _dfoo794 ;
  assign _dfoo863 =
	     source_id__h55665 == 10'd10 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1993 ||
	     source_id__h57161 == 10'd10 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2054 ||
	     _dfoo727 ;
  assign _dfoo864 =
	     (source_id__h55665 == 10'd10 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1993) ?
	       wdata32__h27246[18] :
	       _dfoo796 ;
  assign _dfoo865 =
	     source_id__h55665 == 10'd9 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1993 ||
	     source_id__h57161 == 10'd9 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2054 ||
	     _dfoo729 ;
  assign _dfoo866 =
	     (source_id__h55665 == 10'd9 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1993) ?
	       wdata32__h27246[18] :
	       _dfoo798 ;
  assign _dfoo867 =
	     source_id__h55665 == 10'd8 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1993 ||
	     source_id__h57161 == 10'd8 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2054 ||
	     _dfoo731 ;
  assign _dfoo868 =
	     (source_id__h55665 == 10'd8 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1993) ?
	       wdata32__h27246[18] :
	       _dfoo800 ;
  assign _dfoo869 =
	     source_id__h55665 == 10'd7 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1993 ||
	     source_id__h57161 == 10'd7 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2054 ||
	     _dfoo733 ;
  assign _dfoo870 =
	     (source_id__h55665 == 10'd7 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1993) ?
	       wdata32__h27246[18] :
	       _dfoo802 ;
  assign _dfoo871 =
	     source_id__h55665 == 10'd6 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1993 ||
	     source_id__h57161 == 10'd6 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2054 ||
	     _dfoo735 ;
  assign _dfoo872 =
	     (source_id__h55665 == 10'd6 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1993) ?
	       wdata32__h27246[18] :
	       _dfoo804 ;
  assign _dfoo873 =
	     source_id__h55665 == 10'd5 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1993 ||
	     source_id__h57161 == 10'd5 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2054 ||
	     _dfoo737 ;
  assign _dfoo874 =
	     (source_id__h55665 == 10'd5 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1993) ?
	       wdata32__h27246[18] :
	       _dfoo806 ;
  assign _dfoo875 =
	     source_id__h55665 == 10'd4 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1993 ||
	     source_id__h57161 == 10'd4 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2054 ||
	     _dfoo739 ;
  assign _dfoo876 =
	     (source_id__h55665 == 10'd4 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1993) ?
	       wdata32__h27246[18] :
	       _dfoo808 ;
  assign _dfoo877 =
	     source_id__h55665 == 10'd3 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1993 ||
	     source_id__h57161 == 10'd3 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2054 ||
	     _dfoo741 ;
  assign _dfoo878 =
	     (source_id__h55665 == 10'd3 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1993) ?
	       wdata32__h27246[18] :
	       _dfoo810 ;
  assign _dfoo879 =
	     source_id__h55665 == 10'd2 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1993 ||
	     source_id__h57161 == 10'd2 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2054 ||
	     _dfoo743 ;
  assign _dfoo88 =
	     (source_id__h72121 == 10'd7 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2664) ?
	       wdata32__h27246[29] :
	       _dfoo20 ;
  assign _dfoo880 =
	     (source_id__h55665 == 10'd2 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1993) ?
	       wdata32__h27246[18] :
	       _dfoo812 ;
  assign _dfoo881 =
	     source_id__h55665 == 10'd1 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1993 ||
	     source_id__h57161 == 10'd1 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2054 ||
	     _dfoo745 ;
  assign _dfoo882 =
	     (source_id__h55665 == 10'd1 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1993) ?
	       wdata32__h27246[18] :
	       _dfoo814 ;
  assign _dfoo883 =
	     source_id__h55665 == 10'd0 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1993 ||
	     source_id__h57161 == 10'd0 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2054 ||
	     _dfoo747 ;
  assign _dfoo884 =
	     (source_id__h55665 == 10'd0 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1993) ?
	       wdata32__h27246[18] :
	       _dfoo816 ;
  assign _dfoo886 =
	     (source_id__h54169 == 10'd16 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1932) ?
	       wdata32__h27246[17] :
	       _dfoo818 ;
  assign _dfoo888 =
	     (source_id__h54169 == 10'd15 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1932) ?
	       wdata32__h27246[17] :
	       _dfoo820 ;
  assign _dfoo890 =
	     (source_id__h54169 == 10'd14 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1932) ?
	       wdata32__h27246[17] :
	       _dfoo822 ;
  assign _dfoo892 =
	     (source_id__h54169 == 10'd13 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1932) ?
	       wdata32__h27246[17] :
	       _dfoo824 ;
  assign _dfoo894 =
	     (source_id__h54169 == 10'd12 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1932) ?
	       wdata32__h27246[17] :
	       _dfoo826 ;
  assign _dfoo896 =
	     (source_id__h54169 == 10'd11 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1932) ?
	       wdata32__h27246[17] :
	       _dfoo828 ;
  assign _dfoo898 =
	     (source_id__h54169 == 10'd10 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1932) ?
	       wdata32__h27246[17] :
	       _dfoo830 ;
  assign _dfoo9 =
	     source_id__h73617 == 10'd12 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2725 ||
	     source_id__h75113 == 10'd12 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2786 ;
  assign _dfoo90 =
	     (source_id__h72121 == 10'd6 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2664) ?
	       wdata32__h27246[29] :
	       _dfoo22 ;
  assign _dfoo900 =
	     (source_id__h54169 == 10'd9 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1932) ?
	       wdata32__h27246[17] :
	       _dfoo832 ;
  assign _dfoo902 =
	     (source_id__h54169 == 10'd8 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1932) ?
	       wdata32__h27246[17] :
	       _dfoo834 ;
  assign _dfoo904 =
	     (source_id__h54169 == 10'd7 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1932) ?
	       wdata32__h27246[17] :
	       _dfoo836 ;
  assign _dfoo906 =
	     (source_id__h54169 == 10'd6 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1932) ?
	       wdata32__h27246[17] :
	       _dfoo838 ;
  assign _dfoo908 =
	     (source_id__h54169 == 10'd5 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1932) ?
	       wdata32__h27246[17] :
	       _dfoo840 ;
  assign _dfoo910 =
	     (source_id__h54169 == 10'd4 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1932) ?
	       wdata32__h27246[17] :
	       _dfoo842 ;
  assign _dfoo912 =
	     (source_id__h54169 == 10'd3 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1932) ?
	       wdata32__h27246[17] :
	       _dfoo844 ;
  assign _dfoo914 =
	     (source_id__h54169 == 10'd2 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1932) ?
	       wdata32__h27246[17] :
	       _dfoo846 ;
  assign _dfoo916 =
	     (source_id__h54169 == 10'd1 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1932) ?
	       wdata32__h27246[17] :
	       _dfoo848 ;
  assign _dfoo918 =
	     (source_id__h54169 == 10'd0 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1932) ?
	       wdata32__h27246[17] :
	       _dfoo850 ;
  assign _dfoo92 =
	     (source_id__h72121 == 10'd5 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2664) ?
	       wdata32__h27246[29] :
	       _dfoo24 ;
  assign _dfoo920 =
	     (source_id__h54169 == 10'd16 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1932) ?
	       wdata32__h27246[17] :
	       _dfoo852 ;
  assign _dfoo922 =
	     (source_id__h54169 == 10'd15 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1932) ?
	       wdata32__h27246[17] :
	       _dfoo854 ;
  assign _dfoo924 =
	     (source_id__h54169 == 10'd14 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1932) ?
	       wdata32__h27246[17] :
	       _dfoo856 ;
  assign _dfoo926 =
	     (source_id__h54169 == 10'd13 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1932) ?
	       wdata32__h27246[17] :
	       _dfoo858 ;
  assign _dfoo928 =
	     (source_id__h54169 == 10'd12 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1932) ?
	       wdata32__h27246[17] :
	       _dfoo860 ;
  assign _dfoo930 =
	     (source_id__h54169 == 10'd11 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1932) ?
	       wdata32__h27246[17] :
	       _dfoo862 ;
  assign _dfoo932 =
	     (source_id__h54169 == 10'd10 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1932) ?
	       wdata32__h27246[17] :
	       _dfoo864 ;
  assign _dfoo934 =
	     (source_id__h54169 == 10'd9 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1932) ?
	       wdata32__h27246[17] :
	       _dfoo866 ;
  assign _dfoo936 =
	     (source_id__h54169 == 10'd8 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1932) ?
	       wdata32__h27246[17] :
	       _dfoo868 ;
  assign _dfoo938 =
	     (source_id__h54169 == 10'd7 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1932) ?
	       wdata32__h27246[17] :
	       _dfoo870 ;
  assign _dfoo94 =
	     (source_id__h72121 == 10'd4 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2664) ?
	       wdata32__h27246[29] :
	       _dfoo26 ;
  assign _dfoo940 =
	     (source_id__h54169 == 10'd6 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1932) ?
	       wdata32__h27246[17] :
	       _dfoo872 ;
  assign _dfoo942 =
	     (source_id__h54169 == 10'd5 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1932) ?
	       wdata32__h27246[17] :
	       _dfoo874 ;
  assign _dfoo944 =
	     (source_id__h54169 == 10'd4 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1932) ?
	       wdata32__h27246[17] :
	       _dfoo876 ;
  assign _dfoo946 =
	     (source_id__h54169 == 10'd3 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1932) ?
	       wdata32__h27246[17] :
	       _dfoo878 ;
  assign _dfoo948 =
	     (source_id__h54169 == 10'd2 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1932) ?
	       wdata32__h27246[17] :
	       _dfoo880 ;
  assign _dfoo950 =
	     (source_id__h54169 == 10'd1 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1932) ?
	       wdata32__h27246[17] :
	       _dfoo882 ;
  assign _dfoo952 =
	     (source_id__h54169 == 10'd0 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1932) ?
	       wdata32__h27246[17] :
	       _dfoo884 ;
  assign _dfoo953 =
	     source_id__h52673 == 10'd16 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1871 ||
	     source_id__h54169 == 10'd16 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1932 ||
	     _dfoo817 ;
  assign _dfoo954 =
	     (source_id__h52673 == 10'd16 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1871) ?
	       wdata32__h27246[16] :
	       _dfoo886 ;
  assign _dfoo955 =
	     source_id__h52673 == 10'd15 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1871 ||
	     source_id__h54169 == 10'd15 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1932 ||
	     _dfoo819 ;
  assign _dfoo956 =
	     (source_id__h52673 == 10'd15 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1871) ?
	       wdata32__h27246[16] :
	       _dfoo888 ;
  assign _dfoo957 =
	     source_id__h52673 == 10'd14 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1871 ||
	     source_id__h54169 == 10'd14 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1932 ||
	     _dfoo821 ;
  assign _dfoo958 =
	     (source_id__h52673 == 10'd14 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1871) ?
	       wdata32__h27246[16] :
	       _dfoo890 ;
  assign _dfoo959 =
	     source_id__h52673 == 10'd13 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1871 ||
	     source_id__h54169 == 10'd13 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1932 ||
	     _dfoo823 ;
  assign _dfoo96 =
	     (source_id__h72121 == 10'd3 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2664) ?
	       wdata32__h27246[29] :
	       _dfoo28 ;
  assign _dfoo960 =
	     (source_id__h52673 == 10'd13 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1871) ?
	       wdata32__h27246[16] :
	       _dfoo892 ;
  assign _dfoo961 =
	     source_id__h52673 == 10'd12 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1871 ||
	     source_id__h54169 == 10'd12 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1932 ||
	     _dfoo825 ;
  assign _dfoo962 =
	     (source_id__h52673 == 10'd12 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1871) ?
	       wdata32__h27246[16] :
	       _dfoo894 ;
  assign _dfoo963 =
	     source_id__h52673 == 10'd11 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1871 ||
	     source_id__h54169 == 10'd11 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1932 ||
	     _dfoo827 ;
  assign _dfoo964 =
	     (source_id__h52673 == 10'd11 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1871) ?
	       wdata32__h27246[16] :
	       _dfoo896 ;
  assign _dfoo965 =
	     source_id__h52673 == 10'd10 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1871 ||
	     source_id__h54169 == 10'd10 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1932 ||
	     _dfoo829 ;
  assign _dfoo966 =
	     (source_id__h52673 == 10'd10 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1871) ?
	       wdata32__h27246[16] :
	       _dfoo898 ;
  assign _dfoo967 =
	     source_id__h52673 == 10'd9 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1871 ||
	     source_id__h54169 == 10'd9 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1932 ||
	     _dfoo831 ;
  assign _dfoo968 =
	     (source_id__h52673 == 10'd9 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1871) ?
	       wdata32__h27246[16] :
	       _dfoo900 ;
  assign _dfoo969 =
	     source_id__h52673 == 10'd8 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1871 ||
	     source_id__h54169 == 10'd8 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1932 ||
	     _dfoo833 ;
  assign _dfoo970 =
	     (source_id__h52673 == 10'd8 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1871) ?
	       wdata32__h27246[16] :
	       _dfoo902 ;
  assign _dfoo971 =
	     source_id__h52673 == 10'd7 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1871 ||
	     source_id__h54169 == 10'd7 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1932 ||
	     _dfoo835 ;
  assign _dfoo972 =
	     (source_id__h52673 == 10'd7 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1871) ?
	       wdata32__h27246[16] :
	       _dfoo904 ;
  assign _dfoo973 =
	     source_id__h52673 == 10'd6 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1871 ||
	     source_id__h54169 == 10'd6 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1932 ||
	     _dfoo837 ;
  assign _dfoo974 =
	     (source_id__h52673 == 10'd6 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1871) ?
	       wdata32__h27246[16] :
	       _dfoo906 ;
  assign _dfoo975 =
	     source_id__h52673 == 10'd5 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1871 ||
	     source_id__h54169 == 10'd5 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1932 ||
	     _dfoo839 ;
  assign _dfoo976 =
	     (source_id__h52673 == 10'd5 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1871) ?
	       wdata32__h27246[16] :
	       _dfoo908 ;
  assign _dfoo977 =
	     source_id__h52673 == 10'd4 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1871 ||
	     source_id__h54169 == 10'd4 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1932 ||
	     _dfoo841 ;
  assign _dfoo978 =
	     (source_id__h52673 == 10'd4 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1871) ?
	       wdata32__h27246[16] :
	       _dfoo910 ;
  assign _dfoo979 =
	     source_id__h52673 == 10'd3 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1871 ||
	     source_id__h54169 == 10'd3 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1932 ||
	     _dfoo843 ;
  assign _dfoo98 =
	     (source_id__h72121 == 10'd2 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2664) ?
	       wdata32__h27246[29] :
	       _dfoo30 ;
  assign _dfoo980 =
	     (source_id__h52673 == 10'd3 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1871) ?
	       wdata32__h27246[16] :
	       _dfoo912 ;
  assign _dfoo981 =
	     source_id__h52673 == 10'd2 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1871 ||
	     source_id__h54169 == 10'd2 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1932 ||
	     _dfoo845 ;
  assign _dfoo982 =
	     (source_id__h52673 == 10'd2 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1871) ?
	       wdata32__h27246[16] :
	       _dfoo914 ;
  assign _dfoo983 =
	     source_id__h52673 == 10'd1 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1871 ||
	     source_id__h54169 == 10'd1 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1932 ||
	     _dfoo847 ;
  assign _dfoo984 =
	     (source_id__h52673 == 10'd1 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1871) ?
	       wdata32__h27246[16] :
	       _dfoo916 ;
  assign _dfoo985 =
	     source_id__h52673 == 10'd0 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1871 ||
	     source_id__h54169 == 10'd0 &&
	     addr_offset__h27245[11:7] == 5'd1 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1932 ||
	     _dfoo849 ;
  assign _dfoo986 =
	     (source_id__h52673 == 10'd0 &&
	      addr_offset__h27245[11:7] == 5'd1 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1871) ?
	       wdata32__h27246[16] :
	       _dfoo918 ;
  assign _dfoo987 =
	     source_id__h52673 == 10'd16 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1871 ||
	     source_id__h54169 == 10'd16 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1932 ||
	     _dfoo851 ;
  assign _dfoo988 =
	     (source_id__h52673 == 10'd16 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1871) ?
	       wdata32__h27246[16] :
	       _dfoo920 ;
  assign _dfoo989 =
	     source_id__h52673 == 10'd15 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1871 ||
	     source_id__h54169 == 10'd15 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1932 ||
	     _dfoo853 ;
  assign _dfoo990 =
	     (source_id__h52673 == 10'd15 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1871) ?
	       wdata32__h27246[16] :
	       _dfoo922 ;
  assign _dfoo991 =
	     source_id__h52673 == 10'd14 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1871 ||
	     source_id__h54169 == 10'd14 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1932 ||
	     _dfoo855 ;
  assign _dfoo992 =
	     (source_id__h52673 == 10'd14 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1871) ?
	       wdata32__h27246[16] :
	       _dfoo924 ;
  assign _dfoo993 =
	     source_id__h52673 == 10'd13 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1871 ||
	     source_id__h54169 == 10'd13 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1932 ||
	     _dfoo857 ;
  assign _dfoo994 =
	     (source_id__h52673 == 10'd13 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1871) ?
	       wdata32__h27246[16] :
	       _dfoo926 ;
  assign _dfoo995 =
	     source_id__h52673 == 10'd12 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1871 ||
	     source_id__h54169 == 10'd12 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1932 ||
	     _dfoo859 ;
  assign _dfoo996 =
	     (source_id__h52673 == 10'd12 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1871) ?
	       wdata32__h27246[16] :
	       _dfoo928 ;
  assign _dfoo997 =
	     source_id__h52673 == 10'd11 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1871 ||
	     source_id__h54169 == 10'd11 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1932 ||
	     _dfoo861 ;
  assign _dfoo998 =
	     (source_id__h52673 == 10'd11 &&
	      addr_offset__h27245[11:7] == 5'd0 &&
	      NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1871) ?
	       wdata32__h27246[16] :
	       _dfoo930 ;
  assign _dfoo999 =
	     source_id__h52673 == 10'd10 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1871 ||
	     source_id__h54169 == 10'd10 &&
	     addr_offset__h27245[11:7] == 5'd0 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d1932 ||
	     _dfoo863 ;
  assign a__h81740 =
	     m_vrg_source_ip_16_read__6_AND_NOT_m_vrg_sourc_ETC___d3066 ?
	       m_vrg_source_prio_16 :
	       IF_m_vrg_source_ip_15_read__5_AND_NOT_m_vrg_so_ETC___d3062 ;
  assign a__h83894 =
	     m_vrg_source_ip_16_read__6_AND_NOT_m_vrg_sourc_ETC___d3160 ?
	       m_vrg_source_prio_16 :
	       IF_m_vrg_source_ip_15_read__5_AND_NOT_m_vrg_so_ETC___d3156 ;
  assign addr_offset__h13465 =
	     m_slave_xactor_f_rd_addr$D_OUT[92:29] - m_rg_addr_base ;
  assign addr_offset__h27245 =
	     m_slave_xactor_f_wr_addr$D_OUT[92:29] - m_rg_addr_base ;
  assign b__h81741 =
	     m_vrg_source_ip_16_read__6_AND_NOT_m_vrg_sourc_ETC___d3066 ?
	       5'd16 :
	       IF_m_vrg_source_ip_15_read__5_AND_NOT_m_vrg_so_ETC___d3082 ;
  assign b__h83895 =
	     m_vrg_source_ip_16_read__6_AND_NOT_m_vrg_sourc_ETC___d3160 ?
	       5'd16 :
	       IF_m_vrg_source_ip_15_read__5_AND_NOT_m_vrg_so_ETC___d3176 ;
  assign m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d240 =
	     addr_offset__h13465 < 64'h0000000000003000 ;
  assign m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d242 =
	     addr_offset__h13465[11:7] <= 5'd1 ;
  assign m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d31 =
	     m_slave_xactor_f_rd_addr$D_OUT[92:29] < m_rg_addr_base ;
  assign m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d36 =
	     addr_offset__h13465 < 64'h0000000000001000 ;
  assign m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d40 =
	     addr_offset__h13465[11:2] <= 10'd16 ;
  assign m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d43 =
	     m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d36 &&
	     addr_offset__h13465[11:2] != 10'd0 &&
	     m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d40 &&
	     m_cfg_verbosity != 4'd0 ;
  assign m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d532 =
	     addr_offset__h13465[16:12] <= 5'd1 ;
  assign m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d68 =
	     addr_offset__h13465 < 64'h0000000000002000 ;
  assign m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d71 =
	     source_id_base__h13893 <= 10'd16 ;
  assign m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d2854 =
	     addr_offset__h27245[16:12] <= 5'd1 ;
  assign m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d2860 =
	     addr_offset__h27245[16:12] == 5'd0 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d821 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2857 ;
  assign m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d2862 =
	     addr_offset__h27245[16:12] == 5'd1 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d821 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2857 ;
  assign m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 =
	     m_slave_xactor_f_wr_addr$D_OUT[92:29] < m_rg_addr_base ;
  assign m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d821 =
	     addr_offset__h27245 < 64'h0000000000001000 ;
  assign m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d823 =
	     addr_offset__h27245[11:2] <= 10'd16 ;
  assign m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d837 =
	     addr_offset__h27245[11:2] == 10'd1 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d821 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d823 ;
  assign m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d839 =
	     addr_offset__h27245[11:2] == 10'd2 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d821 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d823 ;
  assign m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d841 =
	     addr_offset__h27245[11:2] == 10'd3 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d821 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d823 ;
  assign m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d843 =
	     addr_offset__h27245[11:2] == 10'd4 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d821 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d823 ;
  assign m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d845 =
	     addr_offset__h27245[11:2] == 10'd5 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d821 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d823 ;
  assign m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d847 =
	     addr_offset__h27245[11:2] == 10'd6 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d821 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d823 ;
  assign m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d849 =
	     addr_offset__h27245[11:2] == 10'd7 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d821 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d823 ;
  assign m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d851 =
	     addr_offset__h27245[11:2] == 10'd8 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d821 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d823 ;
  assign m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d853 =
	     addr_offset__h27245[11:2] == 10'd9 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d821 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d823 ;
  assign m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d855 =
	     addr_offset__h27245[11:2] == 10'd10 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d821 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d823 ;
  assign m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d857 =
	     addr_offset__h27245[11:2] == 10'd11 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d821 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d823 ;
  assign m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d859 =
	     addr_offset__h27245[11:2] == 10'd12 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d821 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d823 ;
  assign m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d861 =
	     addr_offset__h27245[11:2] == 10'd13 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d821 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d823 ;
  assign m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d863 =
	     addr_offset__h27245[11:2] == 10'd14 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d821 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d823 ;
  assign m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d865 =
	     addr_offset__h27245[11:2] == 10'd15 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d821 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d823 ;
  assign m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d867 =
	     addr_offset__h27245[11:2] == 10'd16 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d821 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d823 ;
  assign m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d869 =
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d821 &&
	     addr_offset__h27245[11:2] != 10'd0 &&
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d823 &&
	     m_cfg_verbosity != 4'd0 ;
  assign m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d874 =
	     addr_offset__h27245 < 64'h0000000000002000 ;
  assign m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d877 =
	     source_id_base__h28620 <= 10'd16 ;
  assign m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d888 =
	     addr_offset__h27245 < 64'h0000000000003000 ;
  assign m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d889 =
	     addr_offset__h27245[11:7] <= 5'd1 ;
  assign m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d895 =
	     addr_offset__h27245[11:7] == 5'd0 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d821 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d892 ;
  assign m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d931 =
	     addr_offset__h27245[11:7] == 5'd1 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 &&
	     !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d821 &&
	     NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d892 ;
  assign m_vrg_source_ip_10_read__0_AND_NOT_m_vrg_sourc_ETC___d3036 =
	     m_vrg_source_ip_10 &&
	     m_vrg_source_prio_10 >
	     IF_m_vrg_source_ip_9_read__9_AND_NOT_m_vrg_sou_ETC___d3032 &&
	     m_vvrg_ie_0_10 ;
  assign m_vrg_source_ip_10_read__0_AND_NOT_m_vrg_sourc_ETC___d3130 =
	     m_vrg_source_ip_10 &&
	     m_vrg_source_prio_10 >
	     IF_m_vrg_source_ip_9_read__9_AND_NOT_m_vrg_sou_ETC___d3126 &&
	     m_vvrg_ie_1_10 ;
  assign m_vrg_source_ip_10_read__0_AND_NOT_m_vrg_sourc_ETC___d614 =
	     m_vrg_source_ip_10 &&
	     m_vrg_source_prio_10 >
	     IF_m_vrg_source_ip_9_read__9_AND_NOT_m_vrg_sou_ETC___d608 &&
	     CASE_addr_offset3465_BITS_16_TO_12_0_m_vvrg_ie_ETC__q42 ;
  assign m_vrg_source_ip_11_read__1_AND_NOT_m_vrg_sourc_ETC___d3041 =
	     m_vrg_source_ip_11 &&
	     m_vrg_source_prio_11 >
	     IF_m_vrg_source_ip_10_read__0_AND_NOT_m_vrg_so_ETC___d3037 &&
	     m_vvrg_ie_0_11 ;
  assign m_vrg_source_ip_11_read__1_AND_NOT_m_vrg_sourc_ETC___d3135 =
	     m_vrg_source_ip_11 &&
	     m_vrg_source_prio_11 >
	     IF_m_vrg_source_ip_10_read__0_AND_NOT_m_vrg_so_ETC___d3131 &&
	     m_vvrg_ie_1_11 ;
  assign m_vrg_source_ip_11_read__1_AND_NOT_m_vrg_sourc_ETC___d621 =
	     m_vrg_source_ip_11 &&
	     m_vrg_source_prio_11 >
	     IF_m_vrg_source_ip_10_read__0_AND_NOT_m_vrg_so_ETC___d615 &&
	     CASE_addr_offset3465_BITS_16_TO_12_0_m_vvrg_ie_ETC__q43 ;
  assign m_vrg_source_ip_12_read__2_AND_NOT_m_vrg_sourc_ETC___d3046 =
	     m_vrg_source_ip_12 &&
	     m_vrg_source_prio_12 >
	     IF_m_vrg_source_ip_11_read__1_AND_NOT_m_vrg_so_ETC___d3042 &&
	     m_vvrg_ie_0_12 ;
  assign m_vrg_source_ip_12_read__2_AND_NOT_m_vrg_sourc_ETC___d3140 =
	     m_vrg_source_ip_12 &&
	     m_vrg_source_prio_12 >
	     IF_m_vrg_source_ip_11_read__1_AND_NOT_m_vrg_so_ETC___d3136 &&
	     m_vvrg_ie_1_12 ;
  assign m_vrg_source_ip_12_read__2_AND_NOT_m_vrg_sourc_ETC___d628 =
	     m_vrg_source_ip_12 &&
	     m_vrg_source_prio_12 >
	     IF_m_vrg_source_ip_11_read__1_AND_NOT_m_vrg_so_ETC___d622 &&
	     CASE_addr_offset3465_BITS_16_TO_12_0_m_vvrg_ie_ETC__q44 ;
  assign m_vrg_source_ip_13_read__3_AND_NOT_m_vrg_sourc_ETC___d3051 =
	     m_vrg_source_ip_13 &&
	     m_vrg_source_prio_13 >
	     IF_m_vrg_source_ip_12_read__2_AND_NOT_m_vrg_so_ETC___d3047 &&
	     m_vvrg_ie_0_13 ;
  assign m_vrg_source_ip_13_read__3_AND_NOT_m_vrg_sourc_ETC___d3145 =
	     m_vrg_source_ip_13 &&
	     m_vrg_source_prio_13 >
	     IF_m_vrg_source_ip_12_read__2_AND_NOT_m_vrg_so_ETC___d3141 &&
	     m_vvrg_ie_1_13 ;
  assign m_vrg_source_ip_13_read__3_AND_NOT_m_vrg_sourc_ETC___d635 =
	     m_vrg_source_ip_13 &&
	     m_vrg_source_prio_13 >
	     IF_m_vrg_source_ip_12_read__2_AND_NOT_m_vrg_so_ETC___d629 &&
	     CASE_addr_offset3465_BITS_16_TO_12_0_m_vvrg_ie_ETC__q45 ;
  assign m_vrg_source_ip_13_read__3_AND_NOT_m_vrg_sourc_ETC___d686 =
	     m_vrg_source_ip_13_read__3_AND_NOT_m_vrg_sourc_ETC___d635 ||
	     m_vrg_source_ip_12_read__2_AND_NOT_m_vrg_sourc_ETC___d628 ||
	     m_vrg_source_ip_11_read__1_AND_NOT_m_vrg_sourc_ETC___d621 ||
	     m_vrg_source_ip_10_read__0_AND_NOT_m_vrg_sourc_ETC___d614 ||
	     m_vrg_source_ip_9_read__9_AND_NOT_m_vrg_source_ETC___d607 ||
	     m_vrg_source_ip_8_read__8_AND_NOT_m_vrg_source_ETC___d600 ||
	     m_vrg_source_ip_7_read__7_AND_NOT_m_vrg_source_ETC___d680 ;
  assign m_vrg_source_ip_14_read__4_AND_NOT_m_vrg_sourc_ETC___d3056 =
	     m_vrg_source_ip_14 &&
	     m_vrg_source_prio_14 >
	     IF_m_vrg_source_ip_13_read__3_AND_NOT_m_vrg_so_ETC___d3052 &&
	     m_vvrg_ie_0_14 ;
  assign m_vrg_source_ip_14_read__4_AND_NOT_m_vrg_sourc_ETC___d3150 =
	     m_vrg_source_ip_14 &&
	     m_vrg_source_prio_14 >
	     IF_m_vrg_source_ip_13_read__3_AND_NOT_m_vrg_so_ETC___d3146 &&
	     m_vvrg_ie_1_14 ;
  assign m_vrg_source_ip_14_read__4_AND_NOT_m_vrg_sourc_ETC___d642 =
	     m_vrg_source_ip_14 &&
	     m_vrg_source_prio_14 >
	     IF_m_vrg_source_ip_13_read__3_AND_NOT_m_vrg_so_ETC___d636 &&
	     CASE_addr_offset3465_BITS_16_TO_12_0_m_vvrg_ie_ETC__q46 ;
  assign m_vrg_source_ip_15_read__5_AND_NOT_m_vrg_sourc_ETC___d3061 =
	     m_vrg_source_ip_15 &&
	     m_vrg_source_prio_15 >
	     IF_m_vrg_source_ip_14_read__4_AND_NOT_m_vrg_so_ETC___d3057 &&
	     m_vvrg_ie_0_15 ;
  assign m_vrg_source_ip_15_read__5_AND_NOT_m_vrg_sourc_ETC___d3155 =
	     m_vrg_source_ip_15 &&
	     m_vrg_source_prio_15 >
	     IF_m_vrg_source_ip_14_read__4_AND_NOT_m_vrg_so_ETC___d3151 &&
	     m_vvrg_ie_1_15 ;
  assign m_vrg_source_ip_15_read__5_AND_NOT_m_vrg_sourc_ETC___d649 =
	     m_vrg_source_ip_15 &&
	     m_vrg_source_prio_15 >
	     IF_m_vrg_source_ip_14_read__4_AND_NOT_m_vrg_so_ETC___d643 &&
	     CASE_addr_offset3465_BITS_16_TO_12_0_m_vvrg_ie_ETC__q47 ;
  assign m_vrg_source_ip_16_read__6_AND_NOT_m_vrg_sourc_ETC___d3066 =
	     m_vrg_source_ip_16 &&
	     m_vrg_source_prio_16 >
	     IF_m_vrg_source_ip_15_read__5_AND_NOT_m_vrg_so_ETC___d3062 &&
	     m_vvrg_ie_0_16 ;
  assign m_vrg_source_ip_16_read__6_AND_NOT_m_vrg_sourc_ETC___d3160 =
	     m_vrg_source_ip_16 &&
	     m_vrg_source_prio_16 >
	     IF_m_vrg_source_ip_15_read__5_AND_NOT_m_vrg_so_ETC___d3156 &&
	     m_vvrg_ie_1_16 ;
  assign m_vrg_source_ip_16_read__6_AND_NOT_m_vrg_sourc_ETC___d656 =
	     m_vrg_source_ip_16 &&
	     !m_vrg_source_prio_16_3_ULE_IF_m_vrg_source_ip__ETC___d651 &&
	     CASE_addr_offset3465_BITS_16_TO_12_0_m_vvrg_ie_ETC__q48 ;
  assign m_vrg_source_ip_16_read__6_AND_NOT_m_vrg_sourc_ETC___d689 =
	     m_vrg_source_ip_16_read__6_AND_NOT_m_vrg_sourc_ETC___d656 ||
	     m_vrg_source_ip_15_read__5_AND_NOT_m_vrg_sourc_ETC___d649 ||
	     m_vrg_source_ip_14_read__4_AND_NOT_m_vrg_sourc_ETC___d642 ||
	     m_vrg_source_ip_13_read__3_AND_NOT_m_vrg_sourc_ETC___d686 ;
  assign m_vrg_source_ip_1_read__1_AND_NOT_m_vrg_source_ETC___d551 =
	     m_vrg_source_ip_1 && m_vrg_source_prio_1 != 3'd0 &&
	     CASE_addr_offset3465_BITS_16_TO_12_0_m_vvrg_ie_ETC__q33 ;
  assign m_vrg_source_ip_2_read__2_AND_NOT_m_vrg_source_ETC___d2996 =
	     m_vrg_source_ip_2 &&
	     m_vrg_source_prio_2 >
	     IF_m_vrg_source_ip_1_read__1_AND_NOT_m_vrg_sou_ETC___d2992 &&
	     m_vvrg_ie_0_2 ;
  assign m_vrg_source_ip_2_read__2_AND_NOT_m_vrg_source_ETC___d3090 =
	     m_vrg_source_ip_2 &&
	     m_vrg_source_prio_2 >
	     IF_m_vrg_source_ip_1_read__1_AND_NOT_m_vrg_sou_ETC___d3086 &&
	     m_vvrg_ie_1_2 ;
  assign m_vrg_source_ip_2_read__2_AND_NOT_m_vrg_source_ETC___d558 =
	     m_vrg_source_ip_2 &&
	     m_vrg_source_prio_2 >
	     IF_m_vrg_source_ip_1_read__1_AND_NOT_m_vrg_sou_ETC___d552 &&
	     CASE_addr_offset3465_BITS_16_TO_12_0_m_vvrg_ie_ETC__q34 ;
  assign m_vrg_source_ip_3_read__3_AND_NOT_m_vrg_source_ETC___d3001 =
	     m_vrg_source_ip_3 &&
	     m_vrg_source_prio_3 >
	     IF_m_vrg_source_ip_2_read__2_AND_NOT_m_vrg_sou_ETC___d2997 &&
	     m_vvrg_ie_0_3 ;
  assign m_vrg_source_ip_3_read__3_AND_NOT_m_vrg_source_ETC___d3095 =
	     m_vrg_source_ip_3 &&
	     m_vrg_source_prio_3 >
	     IF_m_vrg_source_ip_2_read__2_AND_NOT_m_vrg_sou_ETC___d3091 &&
	     m_vvrg_ie_1_3 ;
  assign m_vrg_source_ip_3_read__3_AND_NOT_m_vrg_source_ETC___d565 =
	     m_vrg_source_ip_3 &&
	     m_vrg_source_prio_3 >
	     IF_m_vrg_source_ip_2_read__2_AND_NOT_m_vrg_sou_ETC___d559 &&
	     CASE_addr_offset3465_BITS_16_TO_12_0_m_vvrg_ie_ETC__q35 ;
  assign m_vrg_source_ip_4_read__4_AND_NOT_m_vrg_source_ETC___d3006 =
	     m_vrg_source_ip_4 &&
	     m_vrg_source_prio_4 >
	     IF_m_vrg_source_ip_3_read__3_AND_NOT_m_vrg_sou_ETC___d3002 &&
	     m_vvrg_ie_0_4 ;
  assign m_vrg_source_ip_4_read__4_AND_NOT_m_vrg_source_ETC___d3100 =
	     m_vrg_source_ip_4 &&
	     m_vrg_source_prio_4 >
	     IF_m_vrg_source_ip_3_read__3_AND_NOT_m_vrg_sou_ETC___d3096 &&
	     m_vvrg_ie_1_4 ;
  assign m_vrg_source_ip_4_read__4_AND_NOT_m_vrg_source_ETC___d572 =
	     m_vrg_source_ip_4 &&
	     m_vrg_source_prio_4 >
	     IF_m_vrg_source_ip_3_read__3_AND_NOT_m_vrg_sou_ETC___d566 &&
	     CASE_addr_offset3465_BITS_16_TO_12_0_m_vvrg_ie_ETC__q36 ;
  assign m_vrg_source_ip_5_read__5_AND_NOT_m_vrg_source_ETC___d3011 =
	     m_vrg_source_ip_5 &&
	     m_vrg_source_prio_5 >
	     IF_m_vrg_source_ip_4_read__4_AND_NOT_m_vrg_sou_ETC___d3007 &&
	     m_vvrg_ie_0_5 ;
  assign m_vrg_source_ip_5_read__5_AND_NOT_m_vrg_source_ETC___d3105 =
	     m_vrg_source_ip_5 &&
	     m_vrg_source_prio_5 >
	     IF_m_vrg_source_ip_4_read__4_AND_NOT_m_vrg_sou_ETC___d3101 &&
	     m_vvrg_ie_1_5 ;
  assign m_vrg_source_ip_5_read__5_AND_NOT_m_vrg_source_ETC___d579 =
	     m_vrg_source_ip_5 &&
	     m_vrg_source_prio_5 >
	     IF_m_vrg_source_ip_4_read__4_AND_NOT_m_vrg_sou_ETC___d573 &&
	     CASE_addr_offset3465_BITS_16_TO_12_0_m_vvrg_ie_ETC__q37 ;
  assign m_vrg_source_ip_6_read__6_AND_NOT_m_vrg_source_ETC___d3016 =
	     m_vrg_source_ip_6 &&
	     m_vrg_source_prio_6 >
	     IF_m_vrg_source_ip_5_read__5_AND_NOT_m_vrg_sou_ETC___d3012 &&
	     m_vvrg_ie_0_6 ;
  assign m_vrg_source_ip_6_read__6_AND_NOT_m_vrg_source_ETC___d3110 =
	     m_vrg_source_ip_6 &&
	     m_vrg_source_prio_6 >
	     IF_m_vrg_source_ip_5_read__5_AND_NOT_m_vrg_sou_ETC___d3106 &&
	     m_vvrg_ie_1_6 ;
  assign m_vrg_source_ip_6_read__6_AND_NOT_m_vrg_source_ETC___d586 =
	     m_vrg_source_ip_6 &&
	     m_vrg_source_prio_6 >
	     IF_m_vrg_source_ip_5_read__5_AND_NOT_m_vrg_sou_ETC___d580 &&
	     CASE_addr_offset3465_BITS_16_TO_12_0_m_vvrg_ie_ETC__q38 ;
  assign m_vrg_source_ip_7_read__7_AND_NOT_m_vrg_source_ETC___d3021 =
	     m_vrg_source_ip_7 &&
	     m_vrg_source_prio_7 >
	     IF_m_vrg_source_ip_6_read__6_AND_NOT_m_vrg_sou_ETC___d3017 &&
	     m_vvrg_ie_0_7 ;
  assign m_vrg_source_ip_7_read__7_AND_NOT_m_vrg_source_ETC___d3115 =
	     m_vrg_source_ip_7 &&
	     m_vrg_source_prio_7 >
	     IF_m_vrg_source_ip_6_read__6_AND_NOT_m_vrg_sou_ETC___d3111 &&
	     m_vvrg_ie_1_7 ;
  assign m_vrg_source_ip_7_read__7_AND_NOT_m_vrg_source_ETC___d593 =
	     m_vrg_source_ip_7 &&
	     m_vrg_source_prio_7 >
	     IF_m_vrg_source_ip_6_read__6_AND_NOT_m_vrg_sou_ETC___d587 &&
	     CASE_addr_offset3465_BITS_16_TO_12_0_m_vvrg_ie_ETC__q39 ;
  assign m_vrg_source_ip_7_read__7_AND_NOT_m_vrg_source_ETC___d680 =
	     m_vrg_source_ip_7_read__7_AND_NOT_m_vrg_source_ETC___d593 ||
	     m_vrg_source_ip_6_read__6_AND_NOT_m_vrg_source_ETC___d586 ||
	     m_vrg_source_ip_5_read__5_AND_NOT_m_vrg_source_ETC___d579 ||
	     m_vrg_source_ip_4_read__4_AND_NOT_m_vrg_source_ETC___d572 ||
	     m_vrg_source_ip_3_read__3_AND_NOT_m_vrg_source_ETC___d565 ||
	     m_vrg_source_ip_2_read__2_AND_NOT_m_vrg_source_ETC___d558 ||
	     m_vrg_source_ip_1_read__1_AND_NOT_m_vrg_source_ETC___d551 ;
  assign m_vrg_source_ip_8_read__8_AND_NOT_m_vrg_source_ETC___d3026 =
	     m_vrg_source_ip_8 &&
	     m_vrg_source_prio_8 >
	     IF_m_vrg_source_ip_7_read__7_AND_NOT_m_vrg_sou_ETC___d3022 &&
	     m_vvrg_ie_0_8 ;
  assign m_vrg_source_ip_8_read__8_AND_NOT_m_vrg_source_ETC___d3120 =
	     m_vrg_source_ip_8 &&
	     m_vrg_source_prio_8 >
	     IF_m_vrg_source_ip_7_read__7_AND_NOT_m_vrg_sou_ETC___d3116 &&
	     m_vvrg_ie_1_8 ;
  assign m_vrg_source_ip_8_read__8_AND_NOT_m_vrg_source_ETC___d600 =
	     m_vrg_source_ip_8 &&
	     m_vrg_source_prio_8 >
	     IF_m_vrg_source_ip_7_read__7_AND_NOT_m_vrg_sou_ETC___d594 &&
	     CASE_addr_offset3465_BITS_16_TO_12_0_m_vvrg_ie_ETC__q40 ;
  assign m_vrg_source_ip_9_read__9_AND_NOT_m_vrg_source_ETC___d3031 =
	     m_vrg_source_ip_9 &&
	     m_vrg_source_prio_9 >
	     IF_m_vrg_source_ip_8_read__8_AND_NOT_m_vrg_sou_ETC___d3027 &&
	     m_vvrg_ie_0_9 ;
  assign m_vrg_source_ip_9_read__9_AND_NOT_m_vrg_source_ETC___d3125 =
	     m_vrg_source_ip_9 &&
	     m_vrg_source_prio_9 >
	     IF_m_vrg_source_ip_8_read__8_AND_NOT_m_vrg_sou_ETC___d3121 &&
	     m_vvrg_ie_1_9 ;
  assign m_vrg_source_ip_9_read__9_AND_NOT_m_vrg_source_ETC___d607 =
	     m_vrg_source_ip_9 &&
	     m_vrg_source_prio_9 >
	     IF_m_vrg_source_ip_8_read__8_AND_NOT_m_vrg_sou_ETC___d601 &&
	     CASE_addr_offset3465_BITS_16_TO_12_0_m_vvrg_ie_ETC__q41 ;
  assign m_vrg_source_prio_16_3_ULE_IF_m_vrg_source_ip__ETC___d651 =
	     m_vrg_source_prio_16 <=
	     (m_vrg_source_ip_15_read__5_AND_NOT_m_vrg_sourc_ETC___d649 ?
		m_vrg_source_prio_15 :
		IF_m_vrg_source_ip_14_read__4_AND_NOT_m_vrg_so_ETC___d643) ;
  assign max_id__h24210 =
	     m_vrg_source_ip_16_read__6_AND_NOT_m_vrg_sourc_ETC___d656 ?
	       5'd16 :
	       IF_m_vrg_source_ip_15_read__5_AND_NOT_m_vrg_so_ETC___d671 ;
  assign rdata___1__h26714 = { rdata__h26520[31:0], 32'h0 } ;
  assign rdata__h26520 =
	     m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d31 ?
	       64'd0 :
	       y_avValue_fst__h26512 ;
  assign rresp__h26521 =
	     m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d31 ?
	       2'b11 :
	       y_avValue_snd__h26513 ;
  assign source_id__h15937 = { addr_offset__h13465[4:0], 5'd31 } ;
  assign source_id__h16044 = { addr_offset__h13465[4:0], 5'd30 } ;
  assign source_id__h16117 = { addr_offset__h13465[4:0], 5'd29 } ;
  assign source_id__h16190 = { addr_offset__h13465[4:0], 5'd28 } ;
  assign source_id__h16263 = { addr_offset__h13465[4:0], 5'd27 } ;
  assign source_id__h16336 = { addr_offset__h13465[4:0], 5'd26 } ;
  assign source_id__h16409 = { addr_offset__h13465[4:0], 5'd25 } ;
  assign source_id__h16482 = { addr_offset__h13465[4:0], 5'd24 } ;
  assign source_id__h16555 = { addr_offset__h13465[4:0], 5'd23 } ;
  assign source_id__h16628 = { addr_offset__h13465[4:0], 5'd22 } ;
  assign source_id__h16701 = { addr_offset__h13465[4:0], 5'd21 } ;
  assign source_id__h16774 = { addr_offset__h13465[4:0], 5'd20 } ;
  assign source_id__h16847 = { addr_offset__h13465[4:0], 5'd19 } ;
  assign source_id__h16920 = { addr_offset__h13465[4:0], 5'd18 } ;
  assign source_id__h16993 = { addr_offset__h13465[4:0], 5'd17 } ;
  assign source_id__h17066 = { addr_offset__h13465[4:0], 5'd16 } ;
  assign source_id__h17139 = { addr_offset__h13465[4:0], 5'd15 } ;
  assign source_id__h17212 = { addr_offset__h13465[4:0], 5'd14 } ;
  assign source_id__h17285 = { addr_offset__h13465[4:0], 5'd13 } ;
  assign source_id__h17358 = { addr_offset__h13465[4:0], 5'd12 } ;
  assign source_id__h17431 = { addr_offset__h13465[4:0], 5'd11 } ;
  assign source_id__h17504 = { addr_offset__h13465[4:0], 5'd10 } ;
  assign source_id__h17577 = { addr_offset__h13465[4:0], 5'd9 } ;
  assign source_id__h17650 = { addr_offset__h13465[4:0], 5'd8 } ;
  assign source_id__h17723 = { addr_offset__h13465[4:0], 5'd7 } ;
  assign source_id__h17796 = { addr_offset__h13465[4:0], 5'd6 } ;
  assign source_id__h17869 = { addr_offset__h13465[4:0], 5'd5 } ;
  assign source_id__h17942 = { addr_offset__h13465[4:0], 5'd4 } ;
  assign source_id__h18015 = { addr_offset__h13465[4:0], 5'd3 } ;
  assign source_id__h18088 = { addr_offset__h13465[4:0], 5'd2 } ;
  assign source_id__h18161 = { addr_offset__h13465[4:0], 5'd1 } ;
  assign source_id__h20405 = 10'd31 + source_id_base__h13893 ;
  assign source_id__h20581 = 10'd30 + source_id_base__h13893 ;
  assign source_id__h20689 = 10'd29 + source_id_base__h13893 ;
  assign source_id__h20797 = 10'd28 + source_id_base__h13893 ;
  assign source_id__h20905 = 10'd27 + source_id_base__h13893 ;
  assign source_id__h21013 = 10'd26 + source_id_base__h13893 ;
  assign source_id__h21121 = 10'd25 + source_id_base__h13893 ;
  assign source_id__h21229 = 10'd24 + source_id_base__h13893 ;
  assign source_id__h21337 = 10'd23 + source_id_base__h13893 ;
  assign source_id__h21445 = 10'd22 + source_id_base__h13893 ;
  assign source_id__h21553 = 10'd21 + source_id_base__h13893 ;
  assign source_id__h21661 = 10'd20 + source_id_base__h13893 ;
  assign source_id__h21769 = 10'd19 + source_id_base__h13893 ;
  assign source_id__h21877 = 10'd18 + source_id_base__h13893 ;
  assign source_id__h21985 = 10'd17 + source_id_base__h13893 ;
  assign source_id__h22093 = 10'd16 + source_id_base__h13893 ;
  assign source_id__h22201 = 10'd15 + source_id_base__h13893 ;
  assign source_id__h22309 = 10'd14 + source_id_base__h13893 ;
  assign source_id__h22417 = 10'd13 + source_id_base__h13893 ;
  assign source_id__h22525 = 10'd12 + source_id_base__h13893 ;
  assign source_id__h22633 = 10'd11 + source_id_base__h13893 ;
  assign source_id__h22741 = 10'd10 + source_id_base__h13893 ;
  assign source_id__h22849 = 10'd9 + source_id_base__h13893 ;
  assign source_id__h22957 = 10'd8 + source_id_base__h13893 ;
  assign source_id__h23065 = 10'd7 + source_id_base__h13893 ;
  assign source_id__h23173 = 10'd6 + source_id_base__h13893 ;
  assign source_id__h23281 = 10'd5 + source_id_base__h13893 ;
  assign source_id__h23389 = 10'd4 + source_id_base__h13893 ;
  assign source_id__h23497 = 10'd3 + source_id_base__h13893 ;
  assign source_id__h23605 = 10'd2 + source_id_base__h13893 ;
  assign source_id__h23713 = 10'd1 + source_id_base__h13893 ;
  assign source_id__h30233 = { addr_offset__h27245[4:0], 5'd1 } ;
  assign source_id__h31729 = { addr_offset__h27245[4:0], 5'd2 } ;
  assign source_id__h33225 = { addr_offset__h27245[4:0], 5'd3 } ;
  assign source_id__h34721 = { addr_offset__h27245[4:0], 5'd4 } ;
  assign source_id__h36217 = { addr_offset__h27245[4:0], 5'd5 } ;
  assign source_id__h37713 = { addr_offset__h27245[4:0], 5'd6 } ;
  assign source_id__h39209 = { addr_offset__h27245[4:0], 5'd7 } ;
  assign source_id__h40705 = { addr_offset__h27245[4:0], 5'd8 } ;
  assign source_id__h42201 = { addr_offset__h27245[4:0], 5'd9 } ;
  assign source_id__h43697 = { addr_offset__h27245[4:0], 5'd10 } ;
  assign source_id__h45193 = { addr_offset__h27245[4:0], 5'd11 } ;
  assign source_id__h46689 = { addr_offset__h27245[4:0], 5'd12 } ;
  assign source_id__h48185 = { addr_offset__h27245[4:0], 5'd13 } ;
  assign source_id__h49681 = { addr_offset__h27245[4:0], 5'd14 } ;
  assign source_id__h51177 = { addr_offset__h27245[4:0], 5'd15 } ;
  assign source_id__h52673 = { addr_offset__h27245[4:0], 5'd16 } ;
  assign source_id__h54169 = { addr_offset__h27245[4:0], 5'd17 } ;
  assign source_id__h55665 = { addr_offset__h27245[4:0], 5'd18 } ;
  assign source_id__h57161 = { addr_offset__h27245[4:0], 5'd19 } ;
  assign source_id__h58657 = { addr_offset__h27245[4:0], 5'd20 } ;
  assign source_id__h60153 = { addr_offset__h27245[4:0], 5'd21 } ;
  assign source_id__h61649 = { addr_offset__h27245[4:0], 5'd22 } ;
  assign source_id__h63145 = { addr_offset__h27245[4:0], 5'd23 } ;
  assign source_id__h64641 = { addr_offset__h27245[4:0], 5'd24 } ;
  assign source_id__h66137 = { addr_offset__h27245[4:0], 5'd25 } ;
  assign source_id__h67633 = { addr_offset__h27245[4:0], 5'd26 } ;
  assign source_id__h69129 = { addr_offset__h27245[4:0], 5'd27 } ;
  assign source_id__h70625 = { addr_offset__h27245[4:0], 5'd28 } ;
  assign source_id__h72121 = { addr_offset__h27245[4:0], 5'd29 } ;
  assign source_id__h73617 = { addr_offset__h27245[4:0], 5'd30 } ;
  assign source_id__h75113 = { addr_offset__h27245[4:0], 5'd31 } ;
  assign source_id_base__h13893 = { addr_offset__h13465[4:0], 5'h0 } ;
  assign source_id_base__h28620 = { addr_offset__h27245[4:0], 5'h0 } ;
  assign v__h13689 = { 61'd0, x__h13769 } ;
  assign v__h13934 = { 32'd0, v_ip__h13937 } ;
  assign v__h18403 = { 32'd0, v_ie__h18406 } ;
  assign v__h24016 = { 61'd0, x__h24096 } ;
  assign v__h24251 =
	     m_vrg_source_ip_16_read__6_AND_NOT_m_vrg_sourc_ETC___d689 ?
	       v__h25556 :
	       64'd0 ;
  assign v__h25556 = { 59'd0, max_id__h24210 } ;
  assign v__h27250 =
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 ?
	       2'b11 :
	       v__h27435 ;
  assign v__h27435 =
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d821 ?
	       v__h27448 :
	       v__h28425 ;
  assign v__h27448 =
	     (addr_offset__h27245[11:2] != 10'd0 &&
	      m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d823) ?
	       2'b0 :
	       2'b10 ;
  assign v__h28425 =
	     (!m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d821 &&
	      m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d874) ?
	       v__h28444 :
	       v__h28597 ;
  assign v__h28444 =
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d877 ?
	       2'b0 :
	       2'b10 ;
  assign v__h28597 =
	     (!m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d874 &&
	      m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d888) ?
	       v__h28616 :
	       v__h76713 ;
  assign v__h28616 =
	     (m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d877 &&
	      m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d889) ?
	       2'b0 :
	       2'b10 ;
  assign v__h76750 =
	     m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d2854 ?
	       2'b0 :
	       2'b10 ;
  assign v_ie__h18406 =
	     { source_id__h20405 <= 10'd16 &&
	       CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q1,
	       source_id__h20581 <= 10'd16 &&
	       CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q2,
	       source_id__h20689 <= 10'd16 &&
	       CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q3,
	       source_id__h20797 <= 10'd16 &&
	       CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q4,
	       source_id__h20905 <= 10'd16 &&
	       CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q5,
	       source_id__h21013 <= 10'd16 &&
	       CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q6,
	       source_id__h21121 <= 10'd16 &&
	       CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q7,
	       source_id__h21229 <= 10'd16 &&
	       CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q8,
	       source_id__h21337 <= 10'd16 &&
	       CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q9,
	       source_id__h21445 <= 10'd16 &&
	       CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q10,
	       source_id__h21553 <= 10'd16 &&
	       CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q11,
	       source_id__h21661 <= 10'd16 &&
	       CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q12,
	       source_id__h21769 <= 10'd16 &&
	       CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q13,
	       source_id__h21877 <= 10'd16 &&
	       CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q14,
	       source_id__h21985 <= 10'd16 &&
	       CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q15,
	       source_id__h22093 <= 10'd16 &&
	       CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q16,
	       source_id__h22201 <= 10'd16 &&
	       CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q17,
	       source_id__h22309 <= 10'd16 &&
	       CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q18,
	       source_id__h22417 <= 10'd16 &&
	       CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q19,
	       source_id__h22525 <= 10'd16 &&
	       CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q20,
	       source_id__h22633 <= 10'd16 &&
	       CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q21,
	       source_id__h22741 <= 10'd16 &&
	       CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q22,
	       source_id__h22849 <= 10'd16 &&
	       CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q23,
	       source_id__h22957 <= 10'd16 &&
	       CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q24,
	       source_id__h23065 <= 10'd16 &&
	       CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q25,
	       source_id__h23173 <= 10'd16 &&
	       CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q26,
	       source_id__h23281 <= 10'd16 &&
	       CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q27,
	       source_id__h23389 <= 10'd16 &&
	       CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q28,
	       source_id__h23497 <= 10'd16 &&
	       CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q29,
	       source_id__h23605 <= 10'd16 &&
	       CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q30,
	       source_id__h23713 <= 10'd16 &&
	       CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q31,
	       m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d71 &&
	       CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q32 } ;
  assign v_ip__h13937 =
	     { source_id__h15937 <= 10'd16 &&
	       SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d98,
	       source_id__h16044 <= 10'd16 &&
	       SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d102,
	       source_id__h16117 <= 10'd16 &&
	       SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d107,
	       source_id__h16190 <= 10'd16 &&
	       SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d111,
	       source_id__h16263 <= 10'd16 &&
	       SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d116,
	       source_id__h16336 <= 10'd16 &&
	       SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d120,
	       source_id__h16409 <= 10'd16 &&
	       SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d125,
	       source_id__h16482 <= 10'd16 &&
	       SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d129,
	       source_id__h16555 <= 10'd16 &&
	       SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d134,
	       source_id__h16628 <= 10'd16 &&
	       SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d138,
	       source_id__h16701 <= 10'd16 &&
	       SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d143,
	       source_id__h16774 <= 10'd16 &&
	       SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d147,
	       source_id__h16847 <= 10'd16 &&
	       SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d152,
	       source_id__h16920 <= 10'd16 &&
	       SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d156,
	       source_id__h16993 <= 10'd16 &&
	       SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d161,
	       source_id__h17066 <= 10'd16 &&
	       SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d165,
	       source_id__h17139 <= 10'd16 &&
	       SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d170,
	       source_id__h17212 <= 10'd16 &&
	       SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d174,
	       source_id__h17285 <= 10'd16 &&
	       SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d179,
	       source_id__h17358 <= 10'd16 &&
	       SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d183,
	       source_id__h17431 <= 10'd16 &&
	       SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d188,
	       source_id__h17504 <= 10'd16 &&
	       SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d192,
	       source_id__h17577 <= 10'd16 &&
	       SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d197,
	       source_id__h17650 <= 10'd16 &&
	       SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d201,
	       source_id__h17723 <= 10'd16 &&
	       SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d206,
	       source_id__h17796 <= 10'd16 &&
	       SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d210,
	       source_id__h17869 <= 10'd16 &&
	       SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d215,
	       source_id__h17942 <= 10'd16 &&
	       SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d219,
	       source_id__h18015 <= 10'd16 &&
	       SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d224,
	       source_id__h18088 <= 10'd16 &&
	       SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d228,
	       source_id__h18161 <= 10'd16 &&
	       SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d233,
	       m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d71 &&
	       SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d235 } ;
  assign wdata32__h27246 =
	     (addr_offset__h27245[2:0] == 3'd4) ?
	       m_slave_xactor_f_wr_data$D_OUT[72:41] :
	       m_slave_xactor_f_wr_data$D_OUT[40:9] ;
  assign x__h23928 =
	     { addr_offset__h13465[31:16], 4'd0, addr_offset__h13465[11:0] } ;
  assign x__h26677 =
	     (addr_offset__h13465[2:0] == 3'd4) ?
	       rdata___1__h26714 :
	       rdata__h26520 ;
  assign x__h76716 =
	     { addr_offset__h27245[31:16], 4'd0, addr_offset__h27245[11:0] } ;
  assign y_avValue_fst__h26433 =
	     m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d532 ?
	       v__h24251 :
	       64'd0 ;
  assign y_avValue_fst__h26445 =
	     m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d532 ?
	       v__h24016 :
	       64'd0 ;
  assign y_avValue_fst__h26461 =
	     (m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d71 &&
	      m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d242) ?
	       v__h18403 :
	       64'd0 ;
  assign y_avValue_fst__h26477 =
	     m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d71 ?
	       v__h13934 :
	       64'd0 ;
  assign y_avValue_fst__h26482 =
	     (!m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d68 &&
	      m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d240) ?
	       y_avValue_fst__h26461 :
	       y_avValue_fst__h26466 ;
  assign y_avValue_fst__h26493 =
	     (addr_offset__h13465[11:2] != 10'd0 &&
	      m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d40) ?
	       v__h13689 :
	       64'd0 ;
  assign y_avValue_fst__h26498 =
	     (!m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d36 &&
	      m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d68) ?
	       y_avValue_fst__h26477 :
	       y_avValue_fst__h26482 ;
  assign y_avValue_fst__h26512 =
	     m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d36 ?
	       y_avValue_fst__h26493 :
	       y_avValue_fst__h26498 ;
  assign y_avValue_snd__h26446 =
	     m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d532 ?
	       2'b0 :
	       2'b10 ;
  assign y_avValue_snd__h26462 =
	     (m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d71 &&
	      m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d242) ?
	       2'b0 :
	       2'b10 ;
  assign y_avValue_snd__h26478 =
	     m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d71 ?
	       2'b0 :
	       2'b10 ;
  assign y_avValue_snd__h26483 =
	     (!m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d68 &&
	      m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d240) ?
	       y_avValue_snd__h26462 :
	       y_avValue_snd__h26467 ;
  assign y_avValue_snd__h26494 =
	     (addr_offset__h13465[11:2] != 10'd0 &&
	      m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d40) ?
	       2'b0 :
	       2'b10 ;
  assign y_avValue_snd__h26499 =
	     (!m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d36 &&
	      m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d68) ?
	       y_avValue_snd__h26478 :
	       y_avValue_snd__h26483 ;
  assign y_avValue_snd__h26513 =
	     m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d36 ?
	       y_avValue_snd__h26494 :
	       y_avValue_snd__h26499 ;
  always@(addr_offset__h13465 or
	  m_vrg_source_prio_0 or
	  m_vrg_source_prio_1 or
	  m_vrg_source_prio_2 or
	  m_vrg_source_prio_3 or
	  m_vrg_source_prio_4 or
	  m_vrg_source_prio_5 or
	  m_vrg_source_prio_6 or
	  m_vrg_source_prio_7 or
	  m_vrg_source_prio_8 or
	  m_vrg_source_prio_9 or
	  m_vrg_source_prio_10 or
	  m_vrg_source_prio_11 or
	  m_vrg_source_prio_12 or
	  m_vrg_source_prio_13 or
	  m_vrg_source_prio_14 or
	  m_vrg_source_prio_15 or m_vrg_source_prio_16)
  begin
    case (addr_offset__h13465[11:2])
      10'd0: x__h13769 = m_vrg_source_prio_0;
      10'd1: x__h13769 = m_vrg_source_prio_1;
      10'd2: x__h13769 = m_vrg_source_prio_2;
      10'd3: x__h13769 = m_vrg_source_prio_3;
      10'd4: x__h13769 = m_vrg_source_prio_4;
      10'd5: x__h13769 = m_vrg_source_prio_5;
      10'd6: x__h13769 = m_vrg_source_prio_6;
      10'd7: x__h13769 = m_vrg_source_prio_7;
      10'd8: x__h13769 = m_vrg_source_prio_8;
      10'd9: x__h13769 = m_vrg_source_prio_9;
      10'd10: x__h13769 = m_vrg_source_prio_10;
      10'd11: x__h13769 = m_vrg_source_prio_11;
      10'd12: x__h13769 = m_vrg_source_prio_12;
      10'd13: x__h13769 = m_vrg_source_prio_13;
      10'd14: x__h13769 = m_vrg_source_prio_14;
      10'd15: x__h13769 = m_vrg_source_prio_15;
      10'd16: x__h13769 = m_vrg_source_prio_16;
      default: x__h13769 = 3'b010 /* unspecified value */ ;
    endcase
  end
  always@(addr_offset__h13465 or
	  m_vrg_target_threshold_0 or m_vrg_target_threshold_1)
  begin
    case (addr_offset__h13465[16:12])
      5'd0: x__h24096 = m_vrg_target_threshold_0;
      5'd1: x__h24096 = m_vrg_target_threshold_1;
      default: x__h24096 = 3'b010 /* unspecified value */ ;
    endcase
  end
  always@(source_id_base__h13893 or
	  m_vrg_source_ip_0 or
	  m_vrg_source_ip_1 or
	  m_vrg_source_ip_2 or
	  m_vrg_source_ip_3 or
	  m_vrg_source_ip_4 or
	  m_vrg_source_ip_5 or
	  m_vrg_source_ip_6 or
	  m_vrg_source_ip_7 or
	  m_vrg_source_ip_8 or
	  m_vrg_source_ip_9 or
	  m_vrg_source_ip_10 or
	  m_vrg_source_ip_11 or
	  m_vrg_source_ip_12 or
	  m_vrg_source_ip_13 or
	  m_vrg_source_ip_14 or m_vrg_source_ip_15 or m_vrg_source_ip_16)
  begin
    case (source_id_base__h13893)
      10'd0:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d235 =
	      m_vrg_source_ip_0;
      10'd1:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d235 =
	      m_vrg_source_ip_1;
      10'd2:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d235 =
	      m_vrg_source_ip_2;
      10'd3:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d235 =
	      m_vrg_source_ip_3;
      10'd4:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d235 =
	      m_vrg_source_ip_4;
      10'd5:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d235 =
	      m_vrg_source_ip_5;
      10'd6:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d235 =
	      m_vrg_source_ip_6;
      10'd7:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d235 =
	      m_vrg_source_ip_7;
      10'd8:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d235 =
	      m_vrg_source_ip_8;
      10'd9:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d235 =
	      m_vrg_source_ip_9;
      10'd10:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d235 =
	      m_vrg_source_ip_10;
      10'd11:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d235 =
	      m_vrg_source_ip_11;
      10'd12:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d235 =
	      m_vrg_source_ip_12;
      10'd13:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d235 =
	      m_vrg_source_ip_13;
      10'd14:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d235 =
	      m_vrg_source_ip_14;
      10'd15:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d235 =
	      m_vrg_source_ip_15;
      10'd16:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d235 =
	      m_vrg_source_ip_16;
      default: SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d235 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(source_id__h20581 or
	  m_vvrg_ie_0_0 or
	  m_vvrg_ie_0_1 or
	  m_vvrg_ie_0_2 or
	  m_vvrg_ie_0_3 or
	  m_vvrg_ie_0_4 or
	  m_vvrg_ie_0_5 or
	  m_vvrg_ie_0_6 or
	  m_vvrg_ie_0_7 or
	  m_vvrg_ie_0_8 or
	  m_vvrg_ie_0_9 or
	  m_vvrg_ie_0_10 or
	  m_vvrg_ie_0_11 or
	  m_vvrg_ie_0_12 or
	  m_vvrg_ie_0_13 or
	  m_vvrg_ie_0_14 or m_vvrg_ie_0_15 or m_vvrg_ie_0_16)
  begin
    case (source_id__h20581)
      10'd0:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d296 =
	      m_vvrg_ie_0_0;
      10'd1:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d296 =
	      m_vvrg_ie_0_1;
      10'd2:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d296 =
	      m_vvrg_ie_0_2;
      10'd3:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d296 =
	      m_vvrg_ie_0_3;
      10'd4:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d296 =
	      m_vvrg_ie_0_4;
      10'd5:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d296 =
	      m_vvrg_ie_0_5;
      10'd6:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d296 =
	      m_vvrg_ie_0_6;
      10'd7:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d296 =
	      m_vvrg_ie_0_7;
      10'd8:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d296 =
	      m_vvrg_ie_0_8;
      10'd9:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d296 =
	      m_vvrg_ie_0_9;
      10'd10:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d296 =
	      m_vvrg_ie_0_10;
      10'd11:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d296 =
	      m_vvrg_ie_0_11;
      10'd12:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d296 =
	      m_vvrg_ie_0_12;
      10'd13:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d296 =
	      m_vvrg_ie_0_13;
      10'd14:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d296 =
	      m_vvrg_ie_0_14;
      10'd15:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d296 =
	      m_vvrg_ie_0_15;
      10'd16:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d296 =
	      m_vvrg_ie_0_16;
      default: SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d296 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(source_id__h20405 or
	  m_vvrg_ie_0_0 or
	  m_vvrg_ie_0_1 or
	  m_vvrg_ie_0_2 or
	  m_vvrg_ie_0_3 or
	  m_vvrg_ie_0_4 or
	  m_vvrg_ie_0_5 or
	  m_vvrg_ie_0_6 or
	  m_vvrg_ie_0_7 or
	  m_vvrg_ie_0_8 or
	  m_vvrg_ie_0_9 or
	  m_vvrg_ie_0_10 or
	  m_vvrg_ie_0_11 or
	  m_vvrg_ie_0_12 or
	  m_vvrg_ie_0_13 or
	  m_vvrg_ie_0_14 or m_vvrg_ie_0_15 or m_vvrg_ie_0_16)
  begin
    case (source_id__h20405)
      10'd0:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d271 =
	      m_vvrg_ie_0_0;
      10'd1:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d271 =
	      m_vvrg_ie_0_1;
      10'd2:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d271 =
	      m_vvrg_ie_0_2;
      10'd3:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d271 =
	      m_vvrg_ie_0_3;
      10'd4:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d271 =
	      m_vvrg_ie_0_4;
      10'd5:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d271 =
	      m_vvrg_ie_0_5;
      10'd6:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d271 =
	      m_vvrg_ie_0_6;
      10'd7:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d271 =
	      m_vvrg_ie_0_7;
      10'd8:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d271 =
	      m_vvrg_ie_0_8;
      10'd9:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d271 =
	      m_vvrg_ie_0_9;
      10'd10:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d271 =
	      m_vvrg_ie_0_10;
      10'd11:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d271 =
	      m_vvrg_ie_0_11;
      10'd12:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d271 =
	      m_vvrg_ie_0_12;
      10'd13:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d271 =
	      m_vvrg_ie_0_13;
      10'd14:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d271 =
	      m_vvrg_ie_0_14;
      10'd15:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d271 =
	      m_vvrg_ie_0_15;
      10'd16:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d271 =
	      m_vvrg_ie_0_16;
      default: SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d271 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(source_id__h20405 or
	  m_vvrg_ie_1_0 or
	  m_vvrg_ie_1_1 or
	  m_vvrg_ie_1_2 or
	  m_vvrg_ie_1_3 or
	  m_vvrg_ie_1_4 or
	  m_vvrg_ie_1_5 or
	  m_vvrg_ie_1_6 or
	  m_vvrg_ie_1_7 or
	  m_vvrg_ie_1_8 or
	  m_vvrg_ie_1_9 or
	  m_vvrg_ie_1_10 or
	  m_vvrg_ie_1_11 or
	  m_vvrg_ie_1_12 or
	  m_vvrg_ie_1_13 or
	  m_vvrg_ie_1_14 or m_vvrg_ie_1_15 or m_vvrg_ie_1_16)
  begin
    case (source_id__h20405)
      10'd0:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d290 =
	      m_vvrg_ie_1_0;
      10'd1:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d290 =
	      m_vvrg_ie_1_1;
      10'd2:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d290 =
	      m_vvrg_ie_1_2;
      10'd3:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d290 =
	      m_vvrg_ie_1_3;
      10'd4:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d290 =
	      m_vvrg_ie_1_4;
      10'd5:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d290 =
	      m_vvrg_ie_1_5;
      10'd6:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d290 =
	      m_vvrg_ie_1_6;
      10'd7:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d290 =
	      m_vvrg_ie_1_7;
      10'd8:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d290 =
	      m_vvrg_ie_1_8;
      10'd9:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d290 =
	      m_vvrg_ie_1_9;
      10'd10:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d290 =
	      m_vvrg_ie_1_10;
      10'd11:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d290 =
	      m_vvrg_ie_1_11;
      10'd12:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d290 =
	      m_vvrg_ie_1_12;
      10'd13:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d290 =
	      m_vvrg_ie_1_13;
      10'd14:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d290 =
	      m_vvrg_ie_1_14;
      10'd15:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d290 =
	      m_vvrg_ie_1_15;
      10'd16:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d290 =
	      m_vvrg_ie_1_16;
      default: SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d290 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(source_id__h20581 or
	  m_vvrg_ie_1_0 or
	  m_vvrg_ie_1_1 or
	  m_vvrg_ie_1_2 or
	  m_vvrg_ie_1_3 or
	  m_vvrg_ie_1_4 or
	  m_vvrg_ie_1_5 or
	  m_vvrg_ie_1_6 or
	  m_vvrg_ie_1_7 or
	  m_vvrg_ie_1_8 or
	  m_vvrg_ie_1_9 or
	  m_vvrg_ie_1_10 or
	  m_vvrg_ie_1_11 or
	  m_vvrg_ie_1_12 or
	  m_vvrg_ie_1_13 or
	  m_vvrg_ie_1_14 or m_vvrg_ie_1_15 or m_vvrg_ie_1_16)
  begin
    case (source_id__h20581)
      10'd0:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d297 =
	      m_vvrg_ie_1_0;
      10'd1:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d297 =
	      m_vvrg_ie_1_1;
      10'd2:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d297 =
	      m_vvrg_ie_1_2;
      10'd3:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d297 =
	      m_vvrg_ie_1_3;
      10'd4:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d297 =
	      m_vvrg_ie_1_4;
      10'd5:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d297 =
	      m_vvrg_ie_1_5;
      10'd6:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d297 =
	      m_vvrg_ie_1_6;
      10'd7:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d297 =
	      m_vvrg_ie_1_7;
      10'd8:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d297 =
	      m_vvrg_ie_1_8;
      10'd9:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d297 =
	      m_vvrg_ie_1_9;
      10'd10:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d297 =
	      m_vvrg_ie_1_10;
      10'd11:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d297 =
	      m_vvrg_ie_1_11;
      10'd12:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d297 =
	      m_vvrg_ie_1_12;
      10'd13:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d297 =
	      m_vvrg_ie_1_13;
      10'd14:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d297 =
	      m_vvrg_ie_1_14;
      10'd15:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d297 =
	      m_vvrg_ie_1_15;
      10'd16:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d297 =
	      m_vvrg_ie_1_16;
      default: SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d297 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(source_id__h15937 or
	  m_vrg_source_ip_0 or
	  m_vrg_source_ip_1 or
	  m_vrg_source_ip_2 or
	  m_vrg_source_ip_3 or
	  m_vrg_source_ip_4 or
	  m_vrg_source_ip_5 or
	  m_vrg_source_ip_6 or
	  m_vrg_source_ip_7 or
	  m_vrg_source_ip_8 or
	  m_vrg_source_ip_9 or
	  m_vrg_source_ip_10 or
	  m_vrg_source_ip_11 or
	  m_vrg_source_ip_12 or
	  m_vrg_source_ip_13 or
	  m_vrg_source_ip_14 or m_vrg_source_ip_15 or m_vrg_source_ip_16)
  begin
    case (source_id__h15937)
      10'd0:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d98 =
	      m_vrg_source_ip_0;
      10'd1:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d98 =
	      m_vrg_source_ip_1;
      10'd2:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d98 =
	      m_vrg_source_ip_2;
      10'd3:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d98 =
	      m_vrg_source_ip_3;
      10'd4:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d98 =
	      m_vrg_source_ip_4;
      10'd5:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d98 =
	      m_vrg_source_ip_5;
      10'd6:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d98 =
	      m_vrg_source_ip_6;
      10'd7:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d98 =
	      m_vrg_source_ip_7;
      10'd8:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d98 =
	      m_vrg_source_ip_8;
      10'd9:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d98 =
	      m_vrg_source_ip_9;
      10'd10:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d98 =
	      m_vrg_source_ip_10;
      10'd11:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d98 =
	      m_vrg_source_ip_11;
      10'd12:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d98 =
	      m_vrg_source_ip_12;
      10'd13:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d98 =
	      m_vrg_source_ip_13;
      10'd14:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d98 =
	      m_vrg_source_ip_14;
      10'd15:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d98 =
	      m_vrg_source_ip_15;
      10'd16:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d98 =
	      m_vrg_source_ip_16;
      default: SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d98 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(source_id__h20689 or
	  m_vvrg_ie_1_0 or
	  m_vvrg_ie_1_1 or
	  m_vvrg_ie_1_2 or
	  m_vvrg_ie_1_3 or
	  m_vvrg_ie_1_4 or
	  m_vvrg_ie_1_5 or
	  m_vvrg_ie_1_6 or
	  m_vvrg_ie_1_7 or
	  m_vvrg_ie_1_8 or
	  m_vvrg_ie_1_9 or
	  m_vvrg_ie_1_10 or
	  m_vvrg_ie_1_11 or
	  m_vvrg_ie_1_12 or
	  m_vvrg_ie_1_13 or
	  m_vvrg_ie_1_14 or m_vvrg_ie_1_15 or m_vvrg_ie_1_16)
  begin
    case (source_id__h20689)
      10'd0:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d305 =
	      m_vvrg_ie_1_0;
      10'd1:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d305 =
	      m_vvrg_ie_1_1;
      10'd2:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d305 =
	      m_vvrg_ie_1_2;
      10'd3:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d305 =
	      m_vvrg_ie_1_3;
      10'd4:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d305 =
	      m_vvrg_ie_1_4;
      10'd5:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d305 =
	      m_vvrg_ie_1_5;
      10'd6:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d305 =
	      m_vvrg_ie_1_6;
      10'd7:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d305 =
	      m_vvrg_ie_1_7;
      10'd8:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d305 =
	      m_vvrg_ie_1_8;
      10'd9:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d305 =
	      m_vvrg_ie_1_9;
      10'd10:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d305 =
	      m_vvrg_ie_1_10;
      10'd11:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d305 =
	      m_vvrg_ie_1_11;
      10'd12:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d305 =
	      m_vvrg_ie_1_12;
      10'd13:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d305 =
	      m_vvrg_ie_1_13;
      10'd14:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d305 =
	      m_vvrg_ie_1_14;
      10'd15:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d305 =
	      m_vvrg_ie_1_15;
      10'd16:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d305 =
	      m_vvrg_ie_1_16;
      default: SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d305 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(source_id__h20689 or
	  m_vvrg_ie_0_0 or
	  m_vvrg_ie_0_1 or
	  m_vvrg_ie_0_2 or
	  m_vvrg_ie_0_3 or
	  m_vvrg_ie_0_4 or
	  m_vvrg_ie_0_5 or
	  m_vvrg_ie_0_6 or
	  m_vvrg_ie_0_7 or
	  m_vvrg_ie_0_8 or
	  m_vvrg_ie_0_9 or
	  m_vvrg_ie_0_10 or
	  m_vvrg_ie_0_11 or
	  m_vvrg_ie_0_12 or
	  m_vvrg_ie_0_13 or
	  m_vvrg_ie_0_14 or m_vvrg_ie_0_15 or m_vvrg_ie_0_16)
  begin
    case (source_id__h20689)
      10'd0:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d304 =
	      m_vvrg_ie_0_0;
      10'd1:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d304 =
	      m_vvrg_ie_0_1;
      10'd2:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d304 =
	      m_vvrg_ie_0_2;
      10'd3:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d304 =
	      m_vvrg_ie_0_3;
      10'd4:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d304 =
	      m_vvrg_ie_0_4;
      10'd5:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d304 =
	      m_vvrg_ie_0_5;
      10'd6:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d304 =
	      m_vvrg_ie_0_6;
      10'd7:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d304 =
	      m_vvrg_ie_0_7;
      10'd8:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d304 =
	      m_vvrg_ie_0_8;
      10'd9:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d304 =
	      m_vvrg_ie_0_9;
      10'd10:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d304 =
	      m_vvrg_ie_0_10;
      10'd11:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d304 =
	      m_vvrg_ie_0_11;
      10'd12:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d304 =
	      m_vvrg_ie_0_12;
      10'd13:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d304 =
	      m_vvrg_ie_0_13;
      10'd14:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d304 =
	      m_vvrg_ie_0_14;
      10'd15:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d304 =
	      m_vvrg_ie_0_15;
      10'd16:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d304 =
	      m_vvrg_ie_0_16;
      default: SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d304 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(source_id__h20797 or
	  m_vvrg_ie_0_0 or
	  m_vvrg_ie_0_1 or
	  m_vvrg_ie_0_2 or
	  m_vvrg_ie_0_3 or
	  m_vvrg_ie_0_4 or
	  m_vvrg_ie_0_5 or
	  m_vvrg_ie_0_6 or
	  m_vvrg_ie_0_7 or
	  m_vvrg_ie_0_8 or
	  m_vvrg_ie_0_9 or
	  m_vvrg_ie_0_10 or
	  m_vvrg_ie_0_11 or
	  m_vvrg_ie_0_12 or
	  m_vvrg_ie_0_13 or
	  m_vvrg_ie_0_14 or m_vvrg_ie_0_15 or m_vvrg_ie_0_16)
  begin
    case (source_id__h20797)
      10'd0:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d311 =
	      m_vvrg_ie_0_0;
      10'd1:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d311 =
	      m_vvrg_ie_0_1;
      10'd2:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d311 =
	      m_vvrg_ie_0_2;
      10'd3:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d311 =
	      m_vvrg_ie_0_3;
      10'd4:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d311 =
	      m_vvrg_ie_0_4;
      10'd5:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d311 =
	      m_vvrg_ie_0_5;
      10'd6:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d311 =
	      m_vvrg_ie_0_6;
      10'd7:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d311 =
	      m_vvrg_ie_0_7;
      10'd8:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d311 =
	      m_vvrg_ie_0_8;
      10'd9:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d311 =
	      m_vvrg_ie_0_9;
      10'd10:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d311 =
	      m_vvrg_ie_0_10;
      10'd11:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d311 =
	      m_vvrg_ie_0_11;
      10'd12:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d311 =
	      m_vvrg_ie_0_12;
      10'd13:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d311 =
	      m_vvrg_ie_0_13;
      10'd14:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d311 =
	      m_vvrg_ie_0_14;
      10'd15:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d311 =
	      m_vvrg_ie_0_15;
      10'd16:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d311 =
	      m_vvrg_ie_0_16;
      default: SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d311 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(source_id__h16044 or
	  m_vrg_source_ip_0 or
	  m_vrg_source_ip_1 or
	  m_vrg_source_ip_2 or
	  m_vrg_source_ip_3 or
	  m_vrg_source_ip_4 or
	  m_vrg_source_ip_5 or
	  m_vrg_source_ip_6 or
	  m_vrg_source_ip_7 or
	  m_vrg_source_ip_8 or
	  m_vrg_source_ip_9 or
	  m_vrg_source_ip_10 or
	  m_vrg_source_ip_11 or
	  m_vrg_source_ip_12 or
	  m_vrg_source_ip_13 or
	  m_vrg_source_ip_14 or m_vrg_source_ip_15 or m_vrg_source_ip_16)
  begin
    case (source_id__h16044)
      10'd0:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d102 =
	      m_vrg_source_ip_0;
      10'd1:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d102 =
	      m_vrg_source_ip_1;
      10'd2:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d102 =
	      m_vrg_source_ip_2;
      10'd3:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d102 =
	      m_vrg_source_ip_3;
      10'd4:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d102 =
	      m_vrg_source_ip_4;
      10'd5:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d102 =
	      m_vrg_source_ip_5;
      10'd6:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d102 =
	      m_vrg_source_ip_6;
      10'd7:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d102 =
	      m_vrg_source_ip_7;
      10'd8:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d102 =
	      m_vrg_source_ip_8;
      10'd9:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d102 =
	      m_vrg_source_ip_9;
      10'd10:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d102 =
	      m_vrg_source_ip_10;
      10'd11:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d102 =
	      m_vrg_source_ip_11;
      10'd12:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d102 =
	      m_vrg_source_ip_12;
      10'd13:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d102 =
	      m_vrg_source_ip_13;
      10'd14:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d102 =
	      m_vrg_source_ip_14;
      10'd15:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d102 =
	      m_vrg_source_ip_15;
      10'd16:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d102 =
	      m_vrg_source_ip_16;
      default: SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d102 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(source_id__h20797 or
	  m_vvrg_ie_1_0 or
	  m_vvrg_ie_1_1 or
	  m_vvrg_ie_1_2 or
	  m_vvrg_ie_1_3 or
	  m_vvrg_ie_1_4 or
	  m_vvrg_ie_1_5 or
	  m_vvrg_ie_1_6 or
	  m_vvrg_ie_1_7 or
	  m_vvrg_ie_1_8 or
	  m_vvrg_ie_1_9 or
	  m_vvrg_ie_1_10 or
	  m_vvrg_ie_1_11 or
	  m_vvrg_ie_1_12 or
	  m_vvrg_ie_1_13 or
	  m_vvrg_ie_1_14 or m_vvrg_ie_1_15 or m_vvrg_ie_1_16)
  begin
    case (source_id__h20797)
      10'd0:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d312 =
	      m_vvrg_ie_1_0;
      10'd1:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d312 =
	      m_vvrg_ie_1_1;
      10'd2:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d312 =
	      m_vvrg_ie_1_2;
      10'd3:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d312 =
	      m_vvrg_ie_1_3;
      10'd4:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d312 =
	      m_vvrg_ie_1_4;
      10'd5:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d312 =
	      m_vvrg_ie_1_5;
      10'd6:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d312 =
	      m_vvrg_ie_1_6;
      10'd7:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d312 =
	      m_vvrg_ie_1_7;
      10'd8:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d312 =
	      m_vvrg_ie_1_8;
      10'd9:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d312 =
	      m_vvrg_ie_1_9;
      10'd10:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d312 =
	      m_vvrg_ie_1_10;
      10'd11:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d312 =
	      m_vvrg_ie_1_11;
      10'd12:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d312 =
	      m_vvrg_ie_1_12;
      10'd13:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d312 =
	      m_vvrg_ie_1_13;
      10'd14:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d312 =
	      m_vvrg_ie_1_14;
      10'd15:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d312 =
	      m_vvrg_ie_1_15;
      10'd16:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d312 =
	      m_vvrg_ie_1_16;
      default: SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d312 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(source_id__h20905 or
	  m_vvrg_ie_0_0 or
	  m_vvrg_ie_0_1 or
	  m_vvrg_ie_0_2 or
	  m_vvrg_ie_0_3 or
	  m_vvrg_ie_0_4 or
	  m_vvrg_ie_0_5 or
	  m_vvrg_ie_0_6 or
	  m_vvrg_ie_0_7 or
	  m_vvrg_ie_0_8 or
	  m_vvrg_ie_0_9 or
	  m_vvrg_ie_0_10 or
	  m_vvrg_ie_0_11 or
	  m_vvrg_ie_0_12 or
	  m_vvrg_ie_0_13 or
	  m_vvrg_ie_0_14 or m_vvrg_ie_0_15 or m_vvrg_ie_0_16)
  begin
    case (source_id__h20905)
      10'd0:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d319 =
	      m_vvrg_ie_0_0;
      10'd1:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d319 =
	      m_vvrg_ie_0_1;
      10'd2:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d319 =
	      m_vvrg_ie_0_2;
      10'd3:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d319 =
	      m_vvrg_ie_0_3;
      10'd4:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d319 =
	      m_vvrg_ie_0_4;
      10'd5:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d319 =
	      m_vvrg_ie_0_5;
      10'd6:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d319 =
	      m_vvrg_ie_0_6;
      10'd7:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d319 =
	      m_vvrg_ie_0_7;
      10'd8:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d319 =
	      m_vvrg_ie_0_8;
      10'd9:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d319 =
	      m_vvrg_ie_0_9;
      10'd10:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d319 =
	      m_vvrg_ie_0_10;
      10'd11:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d319 =
	      m_vvrg_ie_0_11;
      10'd12:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d319 =
	      m_vvrg_ie_0_12;
      10'd13:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d319 =
	      m_vvrg_ie_0_13;
      10'd14:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d319 =
	      m_vvrg_ie_0_14;
      10'd15:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d319 =
	      m_vvrg_ie_0_15;
      10'd16:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d319 =
	      m_vvrg_ie_0_16;
      default: SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d319 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(source_id__h20905 or
	  m_vvrg_ie_1_0 or
	  m_vvrg_ie_1_1 or
	  m_vvrg_ie_1_2 or
	  m_vvrg_ie_1_3 or
	  m_vvrg_ie_1_4 or
	  m_vvrg_ie_1_5 or
	  m_vvrg_ie_1_6 or
	  m_vvrg_ie_1_7 or
	  m_vvrg_ie_1_8 or
	  m_vvrg_ie_1_9 or
	  m_vvrg_ie_1_10 or
	  m_vvrg_ie_1_11 or
	  m_vvrg_ie_1_12 or
	  m_vvrg_ie_1_13 or
	  m_vvrg_ie_1_14 or m_vvrg_ie_1_15 or m_vvrg_ie_1_16)
  begin
    case (source_id__h20905)
      10'd0:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d320 =
	      m_vvrg_ie_1_0;
      10'd1:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d320 =
	      m_vvrg_ie_1_1;
      10'd2:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d320 =
	      m_vvrg_ie_1_2;
      10'd3:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d320 =
	      m_vvrg_ie_1_3;
      10'd4:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d320 =
	      m_vvrg_ie_1_4;
      10'd5:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d320 =
	      m_vvrg_ie_1_5;
      10'd6:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d320 =
	      m_vvrg_ie_1_6;
      10'd7:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d320 =
	      m_vvrg_ie_1_7;
      10'd8:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d320 =
	      m_vvrg_ie_1_8;
      10'd9:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d320 =
	      m_vvrg_ie_1_9;
      10'd10:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d320 =
	      m_vvrg_ie_1_10;
      10'd11:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d320 =
	      m_vvrg_ie_1_11;
      10'd12:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d320 =
	      m_vvrg_ie_1_12;
      10'd13:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d320 =
	      m_vvrg_ie_1_13;
      10'd14:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d320 =
	      m_vvrg_ie_1_14;
      10'd15:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d320 =
	      m_vvrg_ie_1_15;
      10'd16:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d320 =
	      m_vvrg_ie_1_16;
      default: SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d320 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(source_id__h21013 or
	  m_vvrg_ie_0_0 or
	  m_vvrg_ie_0_1 or
	  m_vvrg_ie_0_2 or
	  m_vvrg_ie_0_3 or
	  m_vvrg_ie_0_4 or
	  m_vvrg_ie_0_5 or
	  m_vvrg_ie_0_6 or
	  m_vvrg_ie_0_7 or
	  m_vvrg_ie_0_8 or
	  m_vvrg_ie_0_9 or
	  m_vvrg_ie_0_10 or
	  m_vvrg_ie_0_11 or
	  m_vvrg_ie_0_12 or
	  m_vvrg_ie_0_13 or
	  m_vvrg_ie_0_14 or m_vvrg_ie_0_15 or m_vvrg_ie_0_16)
  begin
    case (source_id__h21013)
      10'd0:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d326 =
	      m_vvrg_ie_0_0;
      10'd1:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d326 =
	      m_vvrg_ie_0_1;
      10'd2:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d326 =
	      m_vvrg_ie_0_2;
      10'd3:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d326 =
	      m_vvrg_ie_0_3;
      10'd4:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d326 =
	      m_vvrg_ie_0_4;
      10'd5:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d326 =
	      m_vvrg_ie_0_5;
      10'd6:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d326 =
	      m_vvrg_ie_0_6;
      10'd7:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d326 =
	      m_vvrg_ie_0_7;
      10'd8:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d326 =
	      m_vvrg_ie_0_8;
      10'd9:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d326 =
	      m_vvrg_ie_0_9;
      10'd10:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d326 =
	      m_vvrg_ie_0_10;
      10'd11:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d326 =
	      m_vvrg_ie_0_11;
      10'd12:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d326 =
	      m_vvrg_ie_0_12;
      10'd13:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d326 =
	      m_vvrg_ie_0_13;
      10'd14:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d326 =
	      m_vvrg_ie_0_14;
      10'd15:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d326 =
	      m_vvrg_ie_0_15;
      10'd16:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d326 =
	      m_vvrg_ie_0_16;
      default: SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d326 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(source_id__h21013 or
	  m_vvrg_ie_1_0 or
	  m_vvrg_ie_1_1 or
	  m_vvrg_ie_1_2 or
	  m_vvrg_ie_1_3 or
	  m_vvrg_ie_1_4 or
	  m_vvrg_ie_1_5 or
	  m_vvrg_ie_1_6 or
	  m_vvrg_ie_1_7 or
	  m_vvrg_ie_1_8 or
	  m_vvrg_ie_1_9 or
	  m_vvrg_ie_1_10 or
	  m_vvrg_ie_1_11 or
	  m_vvrg_ie_1_12 or
	  m_vvrg_ie_1_13 or
	  m_vvrg_ie_1_14 or m_vvrg_ie_1_15 or m_vvrg_ie_1_16)
  begin
    case (source_id__h21013)
      10'd0:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d327 =
	      m_vvrg_ie_1_0;
      10'd1:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d327 =
	      m_vvrg_ie_1_1;
      10'd2:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d327 =
	      m_vvrg_ie_1_2;
      10'd3:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d327 =
	      m_vvrg_ie_1_3;
      10'd4:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d327 =
	      m_vvrg_ie_1_4;
      10'd5:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d327 =
	      m_vvrg_ie_1_5;
      10'd6:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d327 =
	      m_vvrg_ie_1_6;
      10'd7:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d327 =
	      m_vvrg_ie_1_7;
      10'd8:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d327 =
	      m_vvrg_ie_1_8;
      10'd9:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d327 =
	      m_vvrg_ie_1_9;
      10'd10:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d327 =
	      m_vvrg_ie_1_10;
      10'd11:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d327 =
	      m_vvrg_ie_1_11;
      10'd12:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d327 =
	      m_vvrg_ie_1_12;
      10'd13:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d327 =
	      m_vvrg_ie_1_13;
      10'd14:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d327 =
	      m_vvrg_ie_1_14;
      10'd15:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d327 =
	      m_vvrg_ie_1_15;
      10'd16:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d327 =
	      m_vvrg_ie_1_16;
      default: SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d327 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(source_id__h16117 or
	  m_vrg_source_ip_0 or
	  m_vrg_source_ip_1 or
	  m_vrg_source_ip_2 or
	  m_vrg_source_ip_3 or
	  m_vrg_source_ip_4 or
	  m_vrg_source_ip_5 or
	  m_vrg_source_ip_6 or
	  m_vrg_source_ip_7 or
	  m_vrg_source_ip_8 or
	  m_vrg_source_ip_9 or
	  m_vrg_source_ip_10 or
	  m_vrg_source_ip_11 or
	  m_vrg_source_ip_12 or
	  m_vrg_source_ip_13 or
	  m_vrg_source_ip_14 or m_vrg_source_ip_15 or m_vrg_source_ip_16)
  begin
    case (source_id__h16117)
      10'd0:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d107 =
	      m_vrg_source_ip_0;
      10'd1:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d107 =
	      m_vrg_source_ip_1;
      10'd2:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d107 =
	      m_vrg_source_ip_2;
      10'd3:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d107 =
	      m_vrg_source_ip_3;
      10'd4:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d107 =
	      m_vrg_source_ip_4;
      10'd5:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d107 =
	      m_vrg_source_ip_5;
      10'd6:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d107 =
	      m_vrg_source_ip_6;
      10'd7:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d107 =
	      m_vrg_source_ip_7;
      10'd8:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d107 =
	      m_vrg_source_ip_8;
      10'd9:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d107 =
	      m_vrg_source_ip_9;
      10'd10:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d107 =
	      m_vrg_source_ip_10;
      10'd11:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d107 =
	      m_vrg_source_ip_11;
      10'd12:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d107 =
	      m_vrg_source_ip_12;
      10'd13:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d107 =
	      m_vrg_source_ip_13;
      10'd14:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d107 =
	      m_vrg_source_ip_14;
      10'd15:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d107 =
	      m_vrg_source_ip_15;
      10'd16:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d107 =
	      m_vrg_source_ip_16;
      default: SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d107 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(source_id__h16190 or
	  m_vrg_source_ip_0 or
	  m_vrg_source_ip_1 or
	  m_vrg_source_ip_2 or
	  m_vrg_source_ip_3 or
	  m_vrg_source_ip_4 or
	  m_vrg_source_ip_5 or
	  m_vrg_source_ip_6 or
	  m_vrg_source_ip_7 or
	  m_vrg_source_ip_8 or
	  m_vrg_source_ip_9 or
	  m_vrg_source_ip_10 or
	  m_vrg_source_ip_11 or
	  m_vrg_source_ip_12 or
	  m_vrg_source_ip_13 or
	  m_vrg_source_ip_14 or m_vrg_source_ip_15 or m_vrg_source_ip_16)
  begin
    case (source_id__h16190)
      10'd0:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d111 =
	      m_vrg_source_ip_0;
      10'd1:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d111 =
	      m_vrg_source_ip_1;
      10'd2:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d111 =
	      m_vrg_source_ip_2;
      10'd3:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d111 =
	      m_vrg_source_ip_3;
      10'd4:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d111 =
	      m_vrg_source_ip_4;
      10'd5:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d111 =
	      m_vrg_source_ip_5;
      10'd6:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d111 =
	      m_vrg_source_ip_6;
      10'd7:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d111 =
	      m_vrg_source_ip_7;
      10'd8:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d111 =
	      m_vrg_source_ip_8;
      10'd9:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d111 =
	      m_vrg_source_ip_9;
      10'd10:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d111 =
	      m_vrg_source_ip_10;
      10'd11:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d111 =
	      m_vrg_source_ip_11;
      10'd12:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d111 =
	      m_vrg_source_ip_12;
      10'd13:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d111 =
	      m_vrg_source_ip_13;
      10'd14:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d111 =
	      m_vrg_source_ip_14;
      10'd15:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d111 =
	      m_vrg_source_ip_15;
      10'd16:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d111 =
	      m_vrg_source_ip_16;
      default: SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d111 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(source_id__h21121 or
	  m_vvrg_ie_0_0 or
	  m_vvrg_ie_0_1 or
	  m_vvrg_ie_0_2 or
	  m_vvrg_ie_0_3 or
	  m_vvrg_ie_0_4 or
	  m_vvrg_ie_0_5 or
	  m_vvrg_ie_0_6 or
	  m_vvrg_ie_0_7 or
	  m_vvrg_ie_0_8 or
	  m_vvrg_ie_0_9 or
	  m_vvrg_ie_0_10 or
	  m_vvrg_ie_0_11 or
	  m_vvrg_ie_0_12 or
	  m_vvrg_ie_0_13 or
	  m_vvrg_ie_0_14 or m_vvrg_ie_0_15 or m_vvrg_ie_0_16)
  begin
    case (source_id__h21121)
      10'd0:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d334 =
	      m_vvrg_ie_0_0;
      10'd1:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d334 =
	      m_vvrg_ie_0_1;
      10'd2:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d334 =
	      m_vvrg_ie_0_2;
      10'd3:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d334 =
	      m_vvrg_ie_0_3;
      10'd4:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d334 =
	      m_vvrg_ie_0_4;
      10'd5:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d334 =
	      m_vvrg_ie_0_5;
      10'd6:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d334 =
	      m_vvrg_ie_0_6;
      10'd7:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d334 =
	      m_vvrg_ie_0_7;
      10'd8:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d334 =
	      m_vvrg_ie_0_8;
      10'd9:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d334 =
	      m_vvrg_ie_0_9;
      10'd10:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d334 =
	      m_vvrg_ie_0_10;
      10'd11:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d334 =
	      m_vvrg_ie_0_11;
      10'd12:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d334 =
	      m_vvrg_ie_0_12;
      10'd13:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d334 =
	      m_vvrg_ie_0_13;
      10'd14:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d334 =
	      m_vvrg_ie_0_14;
      10'd15:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d334 =
	      m_vvrg_ie_0_15;
      10'd16:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d334 =
	      m_vvrg_ie_0_16;
      default: SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d334 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(source_id__h21121 or
	  m_vvrg_ie_1_0 or
	  m_vvrg_ie_1_1 or
	  m_vvrg_ie_1_2 or
	  m_vvrg_ie_1_3 or
	  m_vvrg_ie_1_4 or
	  m_vvrg_ie_1_5 or
	  m_vvrg_ie_1_6 or
	  m_vvrg_ie_1_7 or
	  m_vvrg_ie_1_8 or
	  m_vvrg_ie_1_9 or
	  m_vvrg_ie_1_10 or
	  m_vvrg_ie_1_11 or
	  m_vvrg_ie_1_12 or
	  m_vvrg_ie_1_13 or
	  m_vvrg_ie_1_14 or m_vvrg_ie_1_15 or m_vvrg_ie_1_16)
  begin
    case (source_id__h21121)
      10'd0:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d335 =
	      m_vvrg_ie_1_0;
      10'd1:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d335 =
	      m_vvrg_ie_1_1;
      10'd2:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d335 =
	      m_vvrg_ie_1_2;
      10'd3:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d335 =
	      m_vvrg_ie_1_3;
      10'd4:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d335 =
	      m_vvrg_ie_1_4;
      10'd5:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d335 =
	      m_vvrg_ie_1_5;
      10'd6:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d335 =
	      m_vvrg_ie_1_6;
      10'd7:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d335 =
	      m_vvrg_ie_1_7;
      10'd8:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d335 =
	      m_vvrg_ie_1_8;
      10'd9:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d335 =
	      m_vvrg_ie_1_9;
      10'd10:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d335 =
	      m_vvrg_ie_1_10;
      10'd11:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d335 =
	      m_vvrg_ie_1_11;
      10'd12:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d335 =
	      m_vvrg_ie_1_12;
      10'd13:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d335 =
	      m_vvrg_ie_1_13;
      10'd14:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d335 =
	      m_vvrg_ie_1_14;
      10'd15:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d335 =
	      m_vvrg_ie_1_15;
      10'd16:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d335 =
	      m_vvrg_ie_1_16;
      default: SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d335 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(source_id__h21229 or
	  m_vvrg_ie_0_0 or
	  m_vvrg_ie_0_1 or
	  m_vvrg_ie_0_2 or
	  m_vvrg_ie_0_3 or
	  m_vvrg_ie_0_4 or
	  m_vvrg_ie_0_5 or
	  m_vvrg_ie_0_6 or
	  m_vvrg_ie_0_7 or
	  m_vvrg_ie_0_8 or
	  m_vvrg_ie_0_9 or
	  m_vvrg_ie_0_10 or
	  m_vvrg_ie_0_11 or
	  m_vvrg_ie_0_12 or
	  m_vvrg_ie_0_13 or
	  m_vvrg_ie_0_14 or m_vvrg_ie_0_15 or m_vvrg_ie_0_16)
  begin
    case (source_id__h21229)
      10'd0:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d341 =
	      m_vvrg_ie_0_0;
      10'd1:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d341 =
	      m_vvrg_ie_0_1;
      10'd2:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d341 =
	      m_vvrg_ie_0_2;
      10'd3:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d341 =
	      m_vvrg_ie_0_3;
      10'd4:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d341 =
	      m_vvrg_ie_0_4;
      10'd5:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d341 =
	      m_vvrg_ie_0_5;
      10'd6:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d341 =
	      m_vvrg_ie_0_6;
      10'd7:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d341 =
	      m_vvrg_ie_0_7;
      10'd8:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d341 =
	      m_vvrg_ie_0_8;
      10'd9:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d341 =
	      m_vvrg_ie_0_9;
      10'd10:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d341 =
	      m_vvrg_ie_0_10;
      10'd11:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d341 =
	      m_vvrg_ie_0_11;
      10'd12:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d341 =
	      m_vvrg_ie_0_12;
      10'd13:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d341 =
	      m_vvrg_ie_0_13;
      10'd14:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d341 =
	      m_vvrg_ie_0_14;
      10'd15:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d341 =
	      m_vvrg_ie_0_15;
      10'd16:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d341 =
	      m_vvrg_ie_0_16;
      default: SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d341 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(source_id__h16263 or
	  m_vrg_source_ip_0 or
	  m_vrg_source_ip_1 or
	  m_vrg_source_ip_2 or
	  m_vrg_source_ip_3 or
	  m_vrg_source_ip_4 or
	  m_vrg_source_ip_5 or
	  m_vrg_source_ip_6 or
	  m_vrg_source_ip_7 or
	  m_vrg_source_ip_8 or
	  m_vrg_source_ip_9 or
	  m_vrg_source_ip_10 or
	  m_vrg_source_ip_11 or
	  m_vrg_source_ip_12 or
	  m_vrg_source_ip_13 or
	  m_vrg_source_ip_14 or m_vrg_source_ip_15 or m_vrg_source_ip_16)
  begin
    case (source_id__h16263)
      10'd0:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d116 =
	      m_vrg_source_ip_0;
      10'd1:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d116 =
	      m_vrg_source_ip_1;
      10'd2:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d116 =
	      m_vrg_source_ip_2;
      10'd3:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d116 =
	      m_vrg_source_ip_3;
      10'd4:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d116 =
	      m_vrg_source_ip_4;
      10'd5:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d116 =
	      m_vrg_source_ip_5;
      10'd6:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d116 =
	      m_vrg_source_ip_6;
      10'd7:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d116 =
	      m_vrg_source_ip_7;
      10'd8:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d116 =
	      m_vrg_source_ip_8;
      10'd9:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d116 =
	      m_vrg_source_ip_9;
      10'd10:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d116 =
	      m_vrg_source_ip_10;
      10'd11:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d116 =
	      m_vrg_source_ip_11;
      10'd12:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d116 =
	      m_vrg_source_ip_12;
      10'd13:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d116 =
	      m_vrg_source_ip_13;
      10'd14:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d116 =
	      m_vrg_source_ip_14;
      10'd15:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d116 =
	      m_vrg_source_ip_15;
      10'd16:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d116 =
	      m_vrg_source_ip_16;
      default: SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d116 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(source_id__h21229 or
	  m_vvrg_ie_1_0 or
	  m_vvrg_ie_1_1 or
	  m_vvrg_ie_1_2 or
	  m_vvrg_ie_1_3 or
	  m_vvrg_ie_1_4 or
	  m_vvrg_ie_1_5 or
	  m_vvrg_ie_1_6 or
	  m_vvrg_ie_1_7 or
	  m_vvrg_ie_1_8 or
	  m_vvrg_ie_1_9 or
	  m_vvrg_ie_1_10 or
	  m_vvrg_ie_1_11 or
	  m_vvrg_ie_1_12 or
	  m_vvrg_ie_1_13 or
	  m_vvrg_ie_1_14 or m_vvrg_ie_1_15 or m_vvrg_ie_1_16)
  begin
    case (source_id__h21229)
      10'd0:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d342 =
	      m_vvrg_ie_1_0;
      10'd1:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d342 =
	      m_vvrg_ie_1_1;
      10'd2:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d342 =
	      m_vvrg_ie_1_2;
      10'd3:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d342 =
	      m_vvrg_ie_1_3;
      10'd4:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d342 =
	      m_vvrg_ie_1_4;
      10'd5:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d342 =
	      m_vvrg_ie_1_5;
      10'd6:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d342 =
	      m_vvrg_ie_1_6;
      10'd7:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d342 =
	      m_vvrg_ie_1_7;
      10'd8:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d342 =
	      m_vvrg_ie_1_8;
      10'd9:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d342 =
	      m_vvrg_ie_1_9;
      10'd10:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d342 =
	      m_vvrg_ie_1_10;
      10'd11:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d342 =
	      m_vvrg_ie_1_11;
      10'd12:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d342 =
	      m_vvrg_ie_1_12;
      10'd13:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d342 =
	      m_vvrg_ie_1_13;
      10'd14:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d342 =
	      m_vvrg_ie_1_14;
      10'd15:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d342 =
	      m_vvrg_ie_1_15;
      10'd16:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d342 =
	      m_vvrg_ie_1_16;
      default: SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d342 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(source_id__h16336 or
	  m_vrg_source_ip_0 or
	  m_vrg_source_ip_1 or
	  m_vrg_source_ip_2 or
	  m_vrg_source_ip_3 or
	  m_vrg_source_ip_4 or
	  m_vrg_source_ip_5 or
	  m_vrg_source_ip_6 or
	  m_vrg_source_ip_7 or
	  m_vrg_source_ip_8 or
	  m_vrg_source_ip_9 or
	  m_vrg_source_ip_10 or
	  m_vrg_source_ip_11 or
	  m_vrg_source_ip_12 or
	  m_vrg_source_ip_13 or
	  m_vrg_source_ip_14 or m_vrg_source_ip_15 or m_vrg_source_ip_16)
  begin
    case (source_id__h16336)
      10'd0:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d120 =
	      m_vrg_source_ip_0;
      10'd1:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d120 =
	      m_vrg_source_ip_1;
      10'd2:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d120 =
	      m_vrg_source_ip_2;
      10'd3:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d120 =
	      m_vrg_source_ip_3;
      10'd4:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d120 =
	      m_vrg_source_ip_4;
      10'd5:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d120 =
	      m_vrg_source_ip_5;
      10'd6:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d120 =
	      m_vrg_source_ip_6;
      10'd7:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d120 =
	      m_vrg_source_ip_7;
      10'd8:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d120 =
	      m_vrg_source_ip_8;
      10'd9:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d120 =
	      m_vrg_source_ip_9;
      10'd10:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d120 =
	      m_vrg_source_ip_10;
      10'd11:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d120 =
	      m_vrg_source_ip_11;
      10'd12:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d120 =
	      m_vrg_source_ip_12;
      10'd13:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d120 =
	      m_vrg_source_ip_13;
      10'd14:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d120 =
	      m_vrg_source_ip_14;
      10'd15:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d120 =
	      m_vrg_source_ip_15;
      10'd16:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d120 =
	      m_vrg_source_ip_16;
      default: SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d120 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(source_id__h21337 or
	  m_vvrg_ie_0_0 or
	  m_vvrg_ie_0_1 or
	  m_vvrg_ie_0_2 or
	  m_vvrg_ie_0_3 or
	  m_vvrg_ie_0_4 or
	  m_vvrg_ie_0_5 or
	  m_vvrg_ie_0_6 or
	  m_vvrg_ie_0_7 or
	  m_vvrg_ie_0_8 or
	  m_vvrg_ie_0_9 or
	  m_vvrg_ie_0_10 or
	  m_vvrg_ie_0_11 or
	  m_vvrg_ie_0_12 or
	  m_vvrg_ie_0_13 or
	  m_vvrg_ie_0_14 or m_vvrg_ie_0_15 or m_vvrg_ie_0_16)
  begin
    case (source_id__h21337)
      10'd0:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d349 =
	      m_vvrg_ie_0_0;
      10'd1:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d349 =
	      m_vvrg_ie_0_1;
      10'd2:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d349 =
	      m_vvrg_ie_0_2;
      10'd3:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d349 =
	      m_vvrg_ie_0_3;
      10'd4:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d349 =
	      m_vvrg_ie_0_4;
      10'd5:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d349 =
	      m_vvrg_ie_0_5;
      10'd6:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d349 =
	      m_vvrg_ie_0_6;
      10'd7:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d349 =
	      m_vvrg_ie_0_7;
      10'd8:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d349 =
	      m_vvrg_ie_0_8;
      10'd9:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d349 =
	      m_vvrg_ie_0_9;
      10'd10:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d349 =
	      m_vvrg_ie_0_10;
      10'd11:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d349 =
	      m_vvrg_ie_0_11;
      10'd12:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d349 =
	      m_vvrg_ie_0_12;
      10'd13:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d349 =
	      m_vvrg_ie_0_13;
      10'd14:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d349 =
	      m_vvrg_ie_0_14;
      10'd15:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d349 =
	      m_vvrg_ie_0_15;
      10'd16:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d349 =
	      m_vvrg_ie_0_16;
      default: SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d349 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(source_id__h21337 or
	  m_vvrg_ie_1_0 or
	  m_vvrg_ie_1_1 or
	  m_vvrg_ie_1_2 or
	  m_vvrg_ie_1_3 or
	  m_vvrg_ie_1_4 or
	  m_vvrg_ie_1_5 or
	  m_vvrg_ie_1_6 or
	  m_vvrg_ie_1_7 or
	  m_vvrg_ie_1_8 or
	  m_vvrg_ie_1_9 or
	  m_vvrg_ie_1_10 or
	  m_vvrg_ie_1_11 or
	  m_vvrg_ie_1_12 or
	  m_vvrg_ie_1_13 or
	  m_vvrg_ie_1_14 or m_vvrg_ie_1_15 or m_vvrg_ie_1_16)
  begin
    case (source_id__h21337)
      10'd0:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d350 =
	      m_vvrg_ie_1_0;
      10'd1:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d350 =
	      m_vvrg_ie_1_1;
      10'd2:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d350 =
	      m_vvrg_ie_1_2;
      10'd3:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d350 =
	      m_vvrg_ie_1_3;
      10'd4:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d350 =
	      m_vvrg_ie_1_4;
      10'd5:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d350 =
	      m_vvrg_ie_1_5;
      10'd6:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d350 =
	      m_vvrg_ie_1_6;
      10'd7:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d350 =
	      m_vvrg_ie_1_7;
      10'd8:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d350 =
	      m_vvrg_ie_1_8;
      10'd9:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d350 =
	      m_vvrg_ie_1_9;
      10'd10:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d350 =
	      m_vvrg_ie_1_10;
      10'd11:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d350 =
	      m_vvrg_ie_1_11;
      10'd12:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d350 =
	      m_vvrg_ie_1_12;
      10'd13:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d350 =
	      m_vvrg_ie_1_13;
      10'd14:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d350 =
	      m_vvrg_ie_1_14;
      10'd15:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d350 =
	      m_vvrg_ie_1_15;
      10'd16:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d350 =
	      m_vvrg_ie_1_16;
      default: SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d350 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(source_id__h21445 or
	  m_vvrg_ie_0_0 or
	  m_vvrg_ie_0_1 or
	  m_vvrg_ie_0_2 or
	  m_vvrg_ie_0_3 or
	  m_vvrg_ie_0_4 or
	  m_vvrg_ie_0_5 or
	  m_vvrg_ie_0_6 or
	  m_vvrg_ie_0_7 or
	  m_vvrg_ie_0_8 or
	  m_vvrg_ie_0_9 or
	  m_vvrg_ie_0_10 or
	  m_vvrg_ie_0_11 or
	  m_vvrg_ie_0_12 or
	  m_vvrg_ie_0_13 or
	  m_vvrg_ie_0_14 or m_vvrg_ie_0_15 or m_vvrg_ie_0_16)
  begin
    case (source_id__h21445)
      10'd0:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d356 =
	      m_vvrg_ie_0_0;
      10'd1:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d356 =
	      m_vvrg_ie_0_1;
      10'd2:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d356 =
	      m_vvrg_ie_0_2;
      10'd3:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d356 =
	      m_vvrg_ie_0_3;
      10'd4:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d356 =
	      m_vvrg_ie_0_4;
      10'd5:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d356 =
	      m_vvrg_ie_0_5;
      10'd6:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d356 =
	      m_vvrg_ie_0_6;
      10'd7:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d356 =
	      m_vvrg_ie_0_7;
      10'd8:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d356 =
	      m_vvrg_ie_0_8;
      10'd9:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d356 =
	      m_vvrg_ie_0_9;
      10'd10:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d356 =
	      m_vvrg_ie_0_10;
      10'd11:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d356 =
	      m_vvrg_ie_0_11;
      10'd12:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d356 =
	      m_vvrg_ie_0_12;
      10'd13:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d356 =
	      m_vvrg_ie_0_13;
      10'd14:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d356 =
	      m_vvrg_ie_0_14;
      10'd15:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d356 =
	      m_vvrg_ie_0_15;
      10'd16:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d356 =
	      m_vvrg_ie_0_16;
      default: SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d356 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(source_id__h16409 or
	  m_vrg_source_ip_0 or
	  m_vrg_source_ip_1 or
	  m_vrg_source_ip_2 or
	  m_vrg_source_ip_3 or
	  m_vrg_source_ip_4 or
	  m_vrg_source_ip_5 or
	  m_vrg_source_ip_6 or
	  m_vrg_source_ip_7 or
	  m_vrg_source_ip_8 or
	  m_vrg_source_ip_9 or
	  m_vrg_source_ip_10 or
	  m_vrg_source_ip_11 or
	  m_vrg_source_ip_12 or
	  m_vrg_source_ip_13 or
	  m_vrg_source_ip_14 or m_vrg_source_ip_15 or m_vrg_source_ip_16)
  begin
    case (source_id__h16409)
      10'd0:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d125 =
	      m_vrg_source_ip_0;
      10'd1:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d125 =
	      m_vrg_source_ip_1;
      10'd2:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d125 =
	      m_vrg_source_ip_2;
      10'd3:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d125 =
	      m_vrg_source_ip_3;
      10'd4:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d125 =
	      m_vrg_source_ip_4;
      10'd5:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d125 =
	      m_vrg_source_ip_5;
      10'd6:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d125 =
	      m_vrg_source_ip_6;
      10'd7:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d125 =
	      m_vrg_source_ip_7;
      10'd8:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d125 =
	      m_vrg_source_ip_8;
      10'd9:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d125 =
	      m_vrg_source_ip_9;
      10'd10:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d125 =
	      m_vrg_source_ip_10;
      10'd11:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d125 =
	      m_vrg_source_ip_11;
      10'd12:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d125 =
	      m_vrg_source_ip_12;
      10'd13:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d125 =
	      m_vrg_source_ip_13;
      10'd14:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d125 =
	      m_vrg_source_ip_14;
      10'd15:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d125 =
	      m_vrg_source_ip_15;
      10'd16:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d125 =
	      m_vrg_source_ip_16;
      default: SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d125 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(source_id__h21445 or
	  m_vvrg_ie_1_0 or
	  m_vvrg_ie_1_1 or
	  m_vvrg_ie_1_2 or
	  m_vvrg_ie_1_3 or
	  m_vvrg_ie_1_4 or
	  m_vvrg_ie_1_5 or
	  m_vvrg_ie_1_6 or
	  m_vvrg_ie_1_7 or
	  m_vvrg_ie_1_8 or
	  m_vvrg_ie_1_9 or
	  m_vvrg_ie_1_10 or
	  m_vvrg_ie_1_11 or
	  m_vvrg_ie_1_12 or
	  m_vvrg_ie_1_13 or
	  m_vvrg_ie_1_14 or m_vvrg_ie_1_15 or m_vvrg_ie_1_16)
  begin
    case (source_id__h21445)
      10'd0:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d357 =
	      m_vvrg_ie_1_0;
      10'd1:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d357 =
	      m_vvrg_ie_1_1;
      10'd2:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d357 =
	      m_vvrg_ie_1_2;
      10'd3:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d357 =
	      m_vvrg_ie_1_3;
      10'd4:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d357 =
	      m_vvrg_ie_1_4;
      10'd5:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d357 =
	      m_vvrg_ie_1_5;
      10'd6:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d357 =
	      m_vvrg_ie_1_6;
      10'd7:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d357 =
	      m_vvrg_ie_1_7;
      10'd8:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d357 =
	      m_vvrg_ie_1_8;
      10'd9:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d357 =
	      m_vvrg_ie_1_9;
      10'd10:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d357 =
	      m_vvrg_ie_1_10;
      10'd11:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d357 =
	      m_vvrg_ie_1_11;
      10'd12:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d357 =
	      m_vvrg_ie_1_12;
      10'd13:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d357 =
	      m_vvrg_ie_1_13;
      10'd14:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d357 =
	      m_vvrg_ie_1_14;
      10'd15:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d357 =
	      m_vvrg_ie_1_15;
      10'd16:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d357 =
	      m_vvrg_ie_1_16;
      default: SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d357 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(source_id__h16482 or
	  m_vrg_source_ip_0 or
	  m_vrg_source_ip_1 or
	  m_vrg_source_ip_2 or
	  m_vrg_source_ip_3 or
	  m_vrg_source_ip_4 or
	  m_vrg_source_ip_5 or
	  m_vrg_source_ip_6 or
	  m_vrg_source_ip_7 or
	  m_vrg_source_ip_8 or
	  m_vrg_source_ip_9 or
	  m_vrg_source_ip_10 or
	  m_vrg_source_ip_11 or
	  m_vrg_source_ip_12 or
	  m_vrg_source_ip_13 or
	  m_vrg_source_ip_14 or m_vrg_source_ip_15 or m_vrg_source_ip_16)
  begin
    case (source_id__h16482)
      10'd0:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d129 =
	      m_vrg_source_ip_0;
      10'd1:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d129 =
	      m_vrg_source_ip_1;
      10'd2:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d129 =
	      m_vrg_source_ip_2;
      10'd3:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d129 =
	      m_vrg_source_ip_3;
      10'd4:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d129 =
	      m_vrg_source_ip_4;
      10'd5:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d129 =
	      m_vrg_source_ip_5;
      10'd6:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d129 =
	      m_vrg_source_ip_6;
      10'd7:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d129 =
	      m_vrg_source_ip_7;
      10'd8:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d129 =
	      m_vrg_source_ip_8;
      10'd9:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d129 =
	      m_vrg_source_ip_9;
      10'd10:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d129 =
	      m_vrg_source_ip_10;
      10'd11:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d129 =
	      m_vrg_source_ip_11;
      10'd12:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d129 =
	      m_vrg_source_ip_12;
      10'd13:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d129 =
	      m_vrg_source_ip_13;
      10'd14:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d129 =
	      m_vrg_source_ip_14;
      10'd15:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d129 =
	      m_vrg_source_ip_15;
      10'd16:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d129 =
	      m_vrg_source_ip_16;
      default: SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d129 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(source_id__h21553 or
	  m_vvrg_ie_1_0 or
	  m_vvrg_ie_1_1 or
	  m_vvrg_ie_1_2 or
	  m_vvrg_ie_1_3 or
	  m_vvrg_ie_1_4 or
	  m_vvrg_ie_1_5 or
	  m_vvrg_ie_1_6 or
	  m_vvrg_ie_1_7 or
	  m_vvrg_ie_1_8 or
	  m_vvrg_ie_1_9 or
	  m_vvrg_ie_1_10 or
	  m_vvrg_ie_1_11 or
	  m_vvrg_ie_1_12 or
	  m_vvrg_ie_1_13 or
	  m_vvrg_ie_1_14 or m_vvrg_ie_1_15 or m_vvrg_ie_1_16)
  begin
    case (source_id__h21553)
      10'd0:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d365 =
	      m_vvrg_ie_1_0;
      10'd1:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d365 =
	      m_vvrg_ie_1_1;
      10'd2:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d365 =
	      m_vvrg_ie_1_2;
      10'd3:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d365 =
	      m_vvrg_ie_1_3;
      10'd4:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d365 =
	      m_vvrg_ie_1_4;
      10'd5:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d365 =
	      m_vvrg_ie_1_5;
      10'd6:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d365 =
	      m_vvrg_ie_1_6;
      10'd7:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d365 =
	      m_vvrg_ie_1_7;
      10'd8:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d365 =
	      m_vvrg_ie_1_8;
      10'd9:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d365 =
	      m_vvrg_ie_1_9;
      10'd10:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d365 =
	      m_vvrg_ie_1_10;
      10'd11:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d365 =
	      m_vvrg_ie_1_11;
      10'd12:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d365 =
	      m_vvrg_ie_1_12;
      10'd13:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d365 =
	      m_vvrg_ie_1_13;
      10'd14:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d365 =
	      m_vvrg_ie_1_14;
      10'd15:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d365 =
	      m_vvrg_ie_1_15;
      10'd16:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d365 =
	      m_vvrg_ie_1_16;
      default: SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d365 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(source_id__h21553 or
	  m_vvrg_ie_0_0 or
	  m_vvrg_ie_0_1 or
	  m_vvrg_ie_0_2 or
	  m_vvrg_ie_0_3 or
	  m_vvrg_ie_0_4 or
	  m_vvrg_ie_0_5 or
	  m_vvrg_ie_0_6 or
	  m_vvrg_ie_0_7 or
	  m_vvrg_ie_0_8 or
	  m_vvrg_ie_0_9 or
	  m_vvrg_ie_0_10 or
	  m_vvrg_ie_0_11 or
	  m_vvrg_ie_0_12 or
	  m_vvrg_ie_0_13 or
	  m_vvrg_ie_0_14 or m_vvrg_ie_0_15 or m_vvrg_ie_0_16)
  begin
    case (source_id__h21553)
      10'd0:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d364 =
	      m_vvrg_ie_0_0;
      10'd1:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d364 =
	      m_vvrg_ie_0_1;
      10'd2:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d364 =
	      m_vvrg_ie_0_2;
      10'd3:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d364 =
	      m_vvrg_ie_0_3;
      10'd4:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d364 =
	      m_vvrg_ie_0_4;
      10'd5:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d364 =
	      m_vvrg_ie_0_5;
      10'd6:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d364 =
	      m_vvrg_ie_0_6;
      10'd7:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d364 =
	      m_vvrg_ie_0_7;
      10'd8:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d364 =
	      m_vvrg_ie_0_8;
      10'd9:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d364 =
	      m_vvrg_ie_0_9;
      10'd10:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d364 =
	      m_vvrg_ie_0_10;
      10'd11:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d364 =
	      m_vvrg_ie_0_11;
      10'd12:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d364 =
	      m_vvrg_ie_0_12;
      10'd13:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d364 =
	      m_vvrg_ie_0_13;
      10'd14:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d364 =
	      m_vvrg_ie_0_14;
      10'd15:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d364 =
	      m_vvrg_ie_0_15;
      10'd16:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d364 =
	      m_vvrg_ie_0_16;
      default: SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d364 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(source_id__h21661 or
	  m_vvrg_ie_0_0 or
	  m_vvrg_ie_0_1 or
	  m_vvrg_ie_0_2 or
	  m_vvrg_ie_0_3 or
	  m_vvrg_ie_0_4 or
	  m_vvrg_ie_0_5 or
	  m_vvrg_ie_0_6 or
	  m_vvrg_ie_0_7 or
	  m_vvrg_ie_0_8 or
	  m_vvrg_ie_0_9 or
	  m_vvrg_ie_0_10 or
	  m_vvrg_ie_0_11 or
	  m_vvrg_ie_0_12 or
	  m_vvrg_ie_0_13 or
	  m_vvrg_ie_0_14 or m_vvrg_ie_0_15 or m_vvrg_ie_0_16)
  begin
    case (source_id__h21661)
      10'd0:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d371 =
	      m_vvrg_ie_0_0;
      10'd1:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d371 =
	      m_vvrg_ie_0_1;
      10'd2:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d371 =
	      m_vvrg_ie_0_2;
      10'd3:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d371 =
	      m_vvrg_ie_0_3;
      10'd4:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d371 =
	      m_vvrg_ie_0_4;
      10'd5:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d371 =
	      m_vvrg_ie_0_5;
      10'd6:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d371 =
	      m_vvrg_ie_0_6;
      10'd7:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d371 =
	      m_vvrg_ie_0_7;
      10'd8:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d371 =
	      m_vvrg_ie_0_8;
      10'd9:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d371 =
	      m_vvrg_ie_0_9;
      10'd10:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d371 =
	      m_vvrg_ie_0_10;
      10'd11:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d371 =
	      m_vvrg_ie_0_11;
      10'd12:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d371 =
	      m_vvrg_ie_0_12;
      10'd13:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d371 =
	      m_vvrg_ie_0_13;
      10'd14:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d371 =
	      m_vvrg_ie_0_14;
      10'd15:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d371 =
	      m_vvrg_ie_0_15;
      10'd16:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d371 =
	      m_vvrg_ie_0_16;
      default: SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d371 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(source_id__h16555 or
	  m_vrg_source_ip_0 or
	  m_vrg_source_ip_1 or
	  m_vrg_source_ip_2 or
	  m_vrg_source_ip_3 or
	  m_vrg_source_ip_4 or
	  m_vrg_source_ip_5 or
	  m_vrg_source_ip_6 or
	  m_vrg_source_ip_7 or
	  m_vrg_source_ip_8 or
	  m_vrg_source_ip_9 or
	  m_vrg_source_ip_10 or
	  m_vrg_source_ip_11 or
	  m_vrg_source_ip_12 or
	  m_vrg_source_ip_13 or
	  m_vrg_source_ip_14 or m_vrg_source_ip_15 or m_vrg_source_ip_16)
  begin
    case (source_id__h16555)
      10'd0:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d134 =
	      m_vrg_source_ip_0;
      10'd1:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d134 =
	      m_vrg_source_ip_1;
      10'd2:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d134 =
	      m_vrg_source_ip_2;
      10'd3:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d134 =
	      m_vrg_source_ip_3;
      10'd4:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d134 =
	      m_vrg_source_ip_4;
      10'd5:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d134 =
	      m_vrg_source_ip_5;
      10'd6:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d134 =
	      m_vrg_source_ip_6;
      10'd7:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d134 =
	      m_vrg_source_ip_7;
      10'd8:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d134 =
	      m_vrg_source_ip_8;
      10'd9:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d134 =
	      m_vrg_source_ip_9;
      10'd10:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d134 =
	      m_vrg_source_ip_10;
      10'd11:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d134 =
	      m_vrg_source_ip_11;
      10'd12:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d134 =
	      m_vrg_source_ip_12;
      10'd13:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d134 =
	      m_vrg_source_ip_13;
      10'd14:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d134 =
	      m_vrg_source_ip_14;
      10'd15:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d134 =
	      m_vrg_source_ip_15;
      10'd16:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d134 =
	      m_vrg_source_ip_16;
      default: SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d134 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(source_id__h21661 or
	  m_vvrg_ie_1_0 or
	  m_vvrg_ie_1_1 or
	  m_vvrg_ie_1_2 or
	  m_vvrg_ie_1_3 or
	  m_vvrg_ie_1_4 or
	  m_vvrg_ie_1_5 or
	  m_vvrg_ie_1_6 or
	  m_vvrg_ie_1_7 or
	  m_vvrg_ie_1_8 or
	  m_vvrg_ie_1_9 or
	  m_vvrg_ie_1_10 or
	  m_vvrg_ie_1_11 or
	  m_vvrg_ie_1_12 or
	  m_vvrg_ie_1_13 or
	  m_vvrg_ie_1_14 or m_vvrg_ie_1_15 or m_vvrg_ie_1_16)
  begin
    case (source_id__h21661)
      10'd0:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d372 =
	      m_vvrg_ie_1_0;
      10'd1:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d372 =
	      m_vvrg_ie_1_1;
      10'd2:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d372 =
	      m_vvrg_ie_1_2;
      10'd3:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d372 =
	      m_vvrg_ie_1_3;
      10'd4:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d372 =
	      m_vvrg_ie_1_4;
      10'd5:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d372 =
	      m_vvrg_ie_1_5;
      10'd6:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d372 =
	      m_vvrg_ie_1_6;
      10'd7:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d372 =
	      m_vvrg_ie_1_7;
      10'd8:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d372 =
	      m_vvrg_ie_1_8;
      10'd9:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d372 =
	      m_vvrg_ie_1_9;
      10'd10:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d372 =
	      m_vvrg_ie_1_10;
      10'd11:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d372 =
	      m_vvrg_ie_1_11;
      10'd12:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d372 =
	      m_vvrg_ie_1_12;
      10'd13:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d372 =
	      m_vvrg_ie_1_13;
      10'd14:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d372 =
	      m_vvrg_ie_1_14;
      10'd15:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d372 =
	      m_vvrg_ie_1_15;
      10'd16:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d372 =
	      m_vvrg_ie_1_16;
      default: SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d372 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(source_id__h16628 or
	  m_vrg_source_ip_0 or
	  m_vrg_source_ip_1 or
	  m_vrg_source_ip_2 or
	  m_vrg_source_ip_3 or
	  m_vrg_source_ip_4 or
	  m_vrg_source_ip_5 or
	  m_vrg_source_ip_6 or
	  m_vrg_source_ip_7 or
	  m_vrg_source_ip_8 or
	  m_vrg_source_ip_9 or
	  m_vrg_source_ip_10 or
	  m_vrg_source_ip_11 or
	  m_vrg_source_ip_12 or
	  m_vrg_source_ip_13 or
	  m_vrg_source_ip_14 or m_vrg_source_ip_15 or m_vrg_source_ip_16)
  begin
    case (source_id__h16628)
      10'd0:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d138 =
	      m_vrg_source_ip_0;
      10'd1:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d138 =
	      m_vrg_source_ip_1;
      10'd2:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d138 =
	      m_vrg_source_ip_2;
      10'd3:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d138 =
	      m_vrg_source_ip_3;
      10'd4:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d138 =
	      m_vrg_source_ip_4;
      10'd5:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d138 =
	      m_vrg_source_ip_5;
      10'd6:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d138 =
	      m_vrg_source_ip_6;
      10'd7:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d138 =
	      m_vrg_source_ip_7;
      10'd8:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d138 =
	      m_vrg_source_ip_8;
      10'd9:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d138 =
	      m_vrg_source_ip_9;
      10'd10:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d138 =
	      m_vrg_source_ip_10;
      10'd11:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d138 =
	      m_vrg_source_ip_11;
      10'd12:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d138 =
	      m_vrg_source_ip_12;
      10'd13:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d138 =
	      m_vrg_source_ip_13;
      10'd14:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d138 =
	      m_vrg_source_ip_14;
      10'd15:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d138 =
	      m_vrg_source_ip_15;
      10'd16:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d138 =
	      m_vrg_source_ip_16;
      default: SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d138 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(source_id__h21769 or
	  m_vvrg_ie_0_0 or
	  m_vvrg_ie_0_1 or
	  m_vvrg_ie_0_2 or
	  m_vvrg_ie_0_3 or
	  m_vvrg_ie_0_4 or
	  m_vvrg_ie_0_5 or
	  m_vvrg_ie_0_6 or
	  m_vvrg_ie_0_7 or
	  m_vvrg_ie_0_8 or
	  m_vvrg_ie_0_9 or
	  m_vvrg_ie_0_10 or
	  m_vvrg_ie_0_11 or
	  m_vvrg_ie_0_12 or
	  m_vvrg_ie_0_13 or
	  m_vvrg_ie_0_14 or m_vvrg_ie_0_15 or m_vvrg_ie_0_16)
  begin
    case (source_id__h21769)
      10'd0:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d379 =
	      m_vvrg_ie_0_0;
      10'd1:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d379 =
	      m_vvrg_ie_0_1;
      10'd2:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d379 =
	      m_vvrg_ie_0_2;
      10'd3:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d379 =
	      m_vvrg_ie_0_3;
      10'd4:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d379 =
	      m_vvrg_ie_0_4;
      10'd5:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d379 =
	      m_vvrg_ie_0_5;
      10'd6:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d379 =
	      m_vvrg_ie_0_6;
      10'd7:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d379 =
	      m_vvrg_ie_0_7;
      10'd8:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d379 =
	      m_vvrg_ie_0_8;
      10'd9:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d379 =
	      m_vvrg_ie_0_9;
      10'd10:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d379 =
	      m_vvrg_ie_0_10;
      10'd11:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d379 =
	      m_vvrg_ie_0_11;
      10'd12:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d379 =
	      m_vvrg_ie_0_12;
      10'd13:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d379 =
	      m_vvrg_ie_0_13;
      10'd14:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d379 =
	      m_vvrg_ie_0_14;
      10'd15:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d379 =
	      m_vvrg_ie_0_15;
      10'd16:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d379 =
	      m_vvrg_ie_0_16;
      default: SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d379 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(source_id__h21769 or
	  m_vvrg_ie_1_0 or
	  m_vvrg_ie_1_1 or
	  m_vvrg_ie_1_2 or
	  m_vvrg_ie_1_3 or
	  m_vvrg_ie_1_4 or
	  m_vvrg_ie_1_5 or
	  m_vvrg_ie_1_6 or
	  m_vvrg_ie_1_7 or
	  m_vvrg_ie_1_8 or
	  m_vvrg_ie_1_9 or
	  m_vvrg_ie_1_10 or
	  m_vvrg_ie_1_11 or
	  m_vvrg_ie_1_12 or
	  m_vvrg_ie_1_13 or
	  m_vvrg_ie_1_14 or m_vvrg_ie_1_15 or m_vvrg_ie_1_16)
  begin
    case (source_id__h21769)
      10'd0:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d380 =
	      m_vvrg_ie_1_0;
      10'd1:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d380 =
	      m_vvrg_ie_1_1;
      10'd2:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d380 =
	      m_vvrg_ie_1_2;
      10'd3:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d380 =
	      m_vvrg_ie_1_3;
      10'd4:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d380 =
	      m_vvrg_ie_1_4;
      10'd5:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d380 =
	      m_vvrg_ie_1_5;
      10'd6:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d380 =
	      m_vvrg_ie_1_6;
      10'd7:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d380 =
	      m_vvrg_ie_1_7;
      10'd8:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d380 =
	      m_vvrg_ie_1_8;
      10'd9:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d380 =
	      m_vvrg_ie_1_9;
      10'd10:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d380 =
	      m_vvrg_ie_1_10;
      10'd11:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d380 =
	      m_vvrg_ie_1_11;
      10'd12:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d380 =
	      m_vvrg_ie_1_12;
      10'd13:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d380 =
	      m_vvrg_ie_1_13;
      10'd14:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d380 =
	      m_vvrg_ie_1_14;
      10'd15:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d380 =
	      m_vvrg_ie_1_15;
      10'd16:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d380 =
	      m_vvrg_ie_1_16;
      default: SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d380 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(source_id__h21877 or
	  m_vvrg_ie_0_0 or
	  m_vvrg_ie_0_1 or
	  m_vvrg_ie_0_2 or
	  m_vvrg_ie_0_3 or
	  m_vvrg_ie_0_4 or
	  m_vvrg_ie_0_5 or
	  m_vvrg_ie_0_6 or
	  m_vvrg_ie_0_7 or
	  m_vvrg_ie_0_8 or
	  m_vvrg_ie_0_9 or
	  m_vvrg_ie_0_10 or
	  m_vvrg_ie_0_11 or
	  m_vvrg_ie_0_12 or
	  m_vvrg_ie_0_13 or
	  m_vvrg_ie_0_14 or m_vvrg_ie_0_15 or m_vvrg_ie_0_16)
  begin
    case (source_id__h21877)
      10'd0:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d386 =
	      m_vvrg_ie_0_0;
      10'd1:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d386 =
	      m_vvrg_ie_0_1;
      10'd2:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d386 =
	      m_vvrg_ie_0_2;
      10'd3:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d386 =
	      m_vvrg_ie_0_3;
      10'd4:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d386 =
	      m_vvrg_ie_0_4;
      10'd5:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d386 =
	      m_vvrg_ie_0_5;
      10'd6:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d386 =
	      m_vvrg_ie_0_6;
      10'd7:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d386 =
	      m_vvrg_ie_0_7;
      10'd8:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d386 =
	      m_vvrg_ie_0_8;
      10'd9:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d386 =
	      m_vvrg_ie_0_9;
      10'd10:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d386 =
	      m_vvrg_ie_0_10;
      10'd11:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d386 =
	      m_vvrg_ie_0_11;
      10'd12:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d386 =
	      m_vvrg_ie_0_12;
      10'd13:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d386 =
	      m_vvrg_ie_0_13;
      10'd14:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d386 =
	      m_vvrg_ie_0_14;
      10'd15:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d386 =
	      m_vvrg_ie_0_15;
      10'd16:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d386 =
	      m_vvrg_ie_0_16;
      default: SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d386 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(source_id__h16701 or
	  m_vrg_source_ip_0 or
	  m_vrg_source_ip_1 or
	  m_vrg_source_ip_2 or
	  m_vrg_source_ip_3 or
	  m_vrg_source_ip_4 or
	  m_vrg_source_ip_5 or
	  m_vrg_source_ip_6 or
	  m_vrg_source_ip_7 or
	  m_vrg_source_ip_8 or
	  m_vrg_source_ip_9 or
	  m_vrg_source_ip_10 or
	  m_vrg_source_ip_11 or
	  m_vrg_source_ip_12 or
	  m_vrg_source_ip_13 or
	  m_vrg_source_ip_14 or m_vrg_source_ip_15 or m_vrg_source_ip_16)
  begin
    case (source_id__h16701)
      10'd0:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d143 =
	      m_vrg_source_ip_0;
      10'd1:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d143 =
	      m_vrg_source_ip_1;
      10'd2:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d143 =
	      m_vrg_source_ip_2;
      10'd3:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d143 =
	      m_vrg_source_ip_3;
      10'd4:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d143 =
	      m_vrg_source_ip_4;
      10'd5:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d143 =
	      m_vrg_source_ip_5;
      10'd6:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d143 =
	      m_vrg_source_ip_6;
      10'd7:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d143 =
	      m_vrg_source_ip_7;
      10'd8:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d143 =
	      m_vrg_source_ip_8;
      10'd9:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d143 =
	      m_vrg_source_ip_9;
      10'd10:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d143 =
	      m_vrg_source_ip_10;
      10'd11:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d143 =
	      m_vrg_source_ip_11;
      10'd12:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d143 =
	      m_vrg_source_ip_12;
      10'd13:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d143 =
	      m_vrg_source_ip_13;
      10'd14:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d143 =
	      m_vrg_source_ip_14;
      10'd15:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d143 =
	      m_vrg_source_ip_15;
      10'd16:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d143 =
	      m_vrg_source_ip_16;
      default: SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d143 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(source_id__h21877 or
	  m_vvrg_ie_1_0 or
	  m_vvrg_ie_1_1 or
	  m_vvrg_ie_1_2 or
	  m_vvrg_ie_1_3 or
	  m_vvrg_ie_1_4 or
	  m_vvrg_ie_1_5 or
	  m_vvrg_ie_1_6 or
	  m_vvrg_ie_1_7 or
	  m_vvrg_ie_1_8 or
	  m_vvrg_ie_1_9 or
	  m_vvrg_ie_1_10 or
	  m_vvrg_ie_1_11 or
	  m_vvrg_ie_1_12 or
	  m_vvrg_ie_1_13 or
	  m_vvrg_ie_1_14 or m_vvrg_ie_1_15 or m_vvrg_ie_1_16)
  begin
    case (source_id__h21877)
      10'd0:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d387 =
	      m_vvrg_ie_1_0;
      10'd1:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d387 =
	      m_vvrg_ie_1_1;
      10'd2:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d387 =
	      m_vvrg_ie_1_2;
      10'd3:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d387 =
	      m_vvrg_ie_1_3;
      10'd4:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d387 =
	      m_vvrg_ie_1_4;
      10'd5:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d387 =
	      m_vvrg_ie_1_5;
      10'd6:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d387 =
	      m_vvrg_ie_1_6;
      10'd7:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d387 =
	      m_vvrg_ie_1_7;
      10'd8:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d387 =
	      m_vvrg_ie_1_8;
      10'd9:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d387 =
	      m_vvrg_ie_1_9;
      10'd10:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d387 =
	      m_vvrg_ie_1_10;
      10'd11:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d387 =
	      m_vvrg_ie_1_11;
      10'd12:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d387 =
	      m_vvrg_ie_1_12;
      10'd13:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d387 =
	      m_vvrg_ie_1_13;
      10'd14:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d387 =
	      m_vvrg_ie_1_14;
      10'd15:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d387 =
	      m_vvrg_ie_1_15;
      10'd16:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d387 =
	      m_vvrg_ie_1_16;
      default: SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d387 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(source_id__h17358 or
	  m_vrg_source_ip_0 or
	  m_vrg_source_ip_1 or
	  m_vrg_source_ip_2 or
	  m_vrg_source_ip_3 or
	  m_vrg_source_ip_4 or
	  m_vrg_source_ip_5 or
	  m_vrg_source_ip_6 or
	  m_vrg_source_ip_7 or
	  m_vrg_source_ip_8 or
	  m_vrg_source_ip_9 or
	  m_vrg_source_ip_10 or
	  m_vrg_source_ip_11 or
	  m_vrg_source_ip_12 or
	  m_vrg_source_ip_13 or
	  m_vrg_source_ip_14 or m_vrg_source_ip_15 or m_vrg_source_ip_16)
  begin
    case (source_id__h17358)
      10'd0:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d183 =
	      m_vrg_source_ip_0;
      10'd1:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d183 =
	      m_vrg_source_ip_1;
      10'd2:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d183 =
	      m_vrg_source_ip_2;
      10'd3:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d183 =
	      m_vrg_source_ip_3;
      10'd4:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d183 =
	      m_vrg_source_ip_4;
      10'd5:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d183 =
	      m_vrg_source_ip_5;
      10'd6:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d183 =
	      m_vrg_source_ip_6;
      10'd7:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d183 =
	      m_vrg_source_ip_7;
      10'd8:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d183 =
	      m_vrg_source_ip_8;
      10'd9:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d183 =
	      m_vrg_source_ip_9;
      10'd10:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d183 =
	      m_vrg_source_ip_10;
      10'd11:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d183 =
	      m_vrg_source_ip_11;
      10'd12:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d183 =
	      m_vrg_source_ip_12;
      10'd13:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d183 =
	      m_vrg_source_ip_13;
      10'd14:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d183 =
	      m_vrg_source_ip_14;
      10'd15:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d183 =
	      m_vrg_source_ip_15;
      10'd16:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d183 =
	      m_vrg_source_ip_16;
      default: SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d183 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(source_id__h16774 or
	  m_vrg_source_ip_0 or
	  m_vrg_source_ip_1 or
	  m_vrg_source_ip_2 or
	  m_vrg_source_ip_3 or
	  m_vrg_source_ip_4 or
	  m_vrg_source_ip_5 or
	  m_vrg_source_ip_6 or
	  m_vrg_source_ip_7 or
	  m_vrg_source_ip_8 or
	  m_vrg_source_ip_9 or
	  m_vrg_source_ip_10 or
	  m_vrg_source_ip_11 or
	  m_vrg_source_ip_12 or
	  m_vrg_source_ip_13 or
	  m_vrg_source_ip_14 or m_vrg_source_ip_15 or m_vrg_source_ip_16)
  begin
    case (source_id__h16774)
      10'd0:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d147 =
	      m_vrg_source_ip_0;
      10'd1:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d147 =
	      m_vrg_source_ip_1;
      10'd2:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d147 =
	      m_vrg_source_ip_2;
      10'd3:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d147 =
	      m_vrg_source_ip_3;
      10'd4:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d147 =
	      m_vrg_source_ip_4;
      10'd5:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d147 =
	      m_vrg_source_ip_5;
      10'd6:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d147 =
	      m_vrg_source_ip_6;
      10'd7:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d147 =
	      m_vrg_source_ip_7;
      10'd8:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d147 =
	      m_vrg_source_ip_8;
      10'd9:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d147 =
	      m_vrg_source_ip_9;
      10'd10:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d147 =
	      m_vrg_source_ip_10;
      10'd11:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d147 =
	      m_vrg_source_ip_11;
      10'd12:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d147 =
	      m_vrg_source_ip_12;
      10'd13:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d147 =
	      m_vrg_source_ip_13;
      10'd14:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d147 =
	      m_vrg_source_ip_14;
      10'd15:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d147 =
	      m_vrg_source_ip_15;
      10'd16:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d147 =
	      m_vrg_source_ip_16;
      default: SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d147 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(source_id__h21985 or
	  m_vvrg_ie_0_0 or
	  m_vvrg_ie_0_1 or
	  m_vvrg_ie_0_2 or
	  m_vvrg_ie_0_3 or
	  m_vvrg_ie_0_4 or
	  m_vvrg_ie_0_5 or
	  m_vvrg_ie_0_6 or
	  m_vvrg_ie_0_7 or
	  m_vvrg_ie_0_8 or
	  m_vvrg_ie_0_9 or
	  m_vvrg_ie_0_10 or
	  m_vvrg_ie_0_11 or
	  m_vvrg_ie_0_12 or
	  m_vvrg_ie_0_13 or
	  m_vvrg_ie_0_14 or m_vvrg_ie_0_15 or m_vvrg_ie_0_16)
  begin
    case (source_id__h21985)
      10'd0:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d394 =
	      m_vvrg_ie_0_0;
      10'd1:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d394 =
	      m_vvrg_ie_0_1;
      10'd2:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d394 =
	      m_vvrg_ie_0_2;
      10'd3:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d394 =
	      m_vvrg_ie_0_3;
      10'd4:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d394 =
	      m_vvrg_ie_0_4;
      10'd5:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d394 =
	      m_vvrg_ie_0_5;
      10'd6:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d394 =
	      m_vvrg_ie_0_6;
      10'd7:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d394 =
	      m_vvrg_ie_0_7;
      10'd8:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d394 =
	      m_vvrg_ie_0_8;
      10'd9:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d394 =
	      m_vvrg_ie_0_9;
      10'd10:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d394 =
	      m_vvrg_ie_0_10;
      10'd11:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d394 =
	      m_vvrg_ie_0_11;
      10'd12:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d394 =
	      m_vvrg_ie_0_12;
      10'd13:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d394 =
	      m_vvrg_ie_0_13;
      10'd14:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d394 =
	      m_vvrg_ie_0_14;
      10'd15:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d394 =
	      m_vvrg_ie_0_15;
      10'd16:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d394 =
	      m_vvrg_ie_0_16;
      default: SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d394 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(source_id__h21985 or
	  m_vvrg_ie_1_0 or
	  m_vvrg_ie_1_1 or
	  m_vvrg_ie_1_2 or
	  m_vvrg_ie_1_3 or
	  m_vvrg_ie_1_4 or
	  m_vvrg_ie_1_5 or
	  m_vvrg_ie_1_6 or
	  m_vvrg_ie_1_7 or
	  m_vvrg_ie_1_8 or
	  m_vvrg_ie_1_9 or
	  m_vvrg_ie_1_10 or
	  m_vvrg_ie_1_11 or
	  m_vvrg_ie_1_12 or
	  m_vvrg_ie_1_13 or
	  m_vvrg_ie_1_14 or m_vvrg_ie_1_15 or m_vvrg_ie_1_16)
  begin
    case (source_id__h21985)
      10'd0:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d395 =
	      m_vvrg_ie_1_0;
      10'd1:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d395 =
	      m_vvrg_ie_1_1;
      10'd2:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d395 =
	      m_vvrg_ie_1_2;
      10'd3:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d395 =
	      m_vvrg_ie_1_3;
      10'd4:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d395 =
	      m_vvrg_ie_1_4;
      10'd5:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d395 =
	      m_vvrg_ie_1_5;
      10'd6:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d395 =
	      m_vvrg_ie_1_6;
      10'd7:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d395 =
	      m_vvrg_ie_1_7;
      10'd8:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d395 =
	      m_vvrg_ie_1_8;
      10'd9:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d395 =
	      m_vvrg_ie_1_9;
      10'd10:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d395 =
	      m_vvrg_ie_1_10;
      10'd11:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d395 =
	      m_vvrg_ie_1_11;
      10'd12:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d395 =
	      m_vvrg_ie_1_12;
      10'd13:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d395 =
	      m_vvrg_ie_1_13;
      10'd14:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d395 =
	      m_vvrg_ie_1_14;
      10'd15:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d395 =
	      m_vvrg_ie_1_15;
      10'd16:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d395 =
	      m_vvrg_ie_1_16;
      default: SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d395 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(source_id__h22093 or
	  m_vvrg_ie_0_0 or
	  m_vvrg_ie_0_1 or
	  m_vvrg_ie_0_2 or
	  m_vvrg_ie_0_3 or
	  m_vvrg_ie_0_4 or
	  m_vvrg_ie_0_5 or
	  m_vvrg_ie_0_6 or
	  m_vvrg_ie_0_7 or
	  m_vvrg_ie_0_8 or
	  m_vvrg_ie_0_9 or
	  m_vvrg_ie_0_10 or
	  m_vvrg_ie_0_11 or
	  m_vvrg_ie_0_12 or
	  m_vvrg_ie_0_13 or
	  m_vvrg_ie_0_14 or m_vvrg_ie_0_15 or m_vvrg_ie_0_16)
  begin
    case (source_id__h22093)
      10'd0:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d401 =
	      m_vvrg_ie_0_0;
      10'd1:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d401 =
	      m_vvrg_ie_0_1;
      10'd2:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d401 =
	      m_vvrg_ie_0_2;
      10'd3:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d401 =
	      m_vvrg_ie_0_3;
      10'd4:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d401 =
	      m_vvrg_ie_0_4;
      10'd5:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d401 =
	      m_vvrg_ie_0_5;
      10'd6:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d401 =
	      m_vvrg_ie_0_6;
      10'd7:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d401 =
	      m_vvrg_ie_0_7;
      10'd8:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d401 =
	      m_vvrg_ie_0_8;
      10'd9:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d401 =
	      m_vvrg_ie_0_9;
      10'd10:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d401 =
	      m_vvrg_ie_0_10;
      10'd11:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d401 =
	      m_vvrg_ie_0_11;
      10'd12:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d401 =
	      m_vvrg_ie_0_12;
      10'd13:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d401 =
	      m_vvrg_ie_0_13;
      10'd14:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d401 =
	      m_vvrg_ie_0_14;
      10'd15:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d401 =
	      m_vvrg_ie_0_15;
      10'd16:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d401 =
	      m_vvrg_ie_0_16;
      default: SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d401 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(source_id__h16847 or
	  m_vrg_source_ip_0 or
	  m_vrg_source_ip_1 or
	  m_vrg_source_ip_2 or
	  m_vrg_source_ip_3 or
	  m_vrg_source_ip_4 or
	  m_vrg_source_ip_5 or
	  m_vrg_source_ip_6 or
	  m_vrg_source_ip_7 or
	  m_vrg_source_ip_8 or
	  m_vrg_source_ip_9 or
	  m_vrg_source_ip_10 or
	  m_vrg_source_ip_11 or
	  m_vrg_source_ip_12 or
	  m_vrg_source_ip_13 or
	  m_vrg_source_ip_14 or m_vrg_source_ip_15 or m_vrg_source_ip_16)
  begin
    case (source_id__h16847)
      10'd0:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d152 =
	      m_vrg_source_ip_0;
      10'd1:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d152 =
	      m_vrg_source_ip_1;
      10'd2:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d152 =
	      m_vrg_source_ip_2;
      10'd3:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d152 =
	      m_vrg_source_ip_3;
      10'd4:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d152 =
	      m_vrg_source_ip_4;
      10'd5:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d152 =
	      m_vrg_source_ip_5;
      10'd6:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d152 =
	      m_vrg_source_ip_6;
      10'd7:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d152 =
	      m_vrg_source_ip_7;
      10'd8:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d152 =
	      m_vrg_source_ip_8;
      10'd9:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d152 =
	      m_vrg_source_ip_9;
      10'd10:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d152 =
	      m_vrg_source_ip_10;
      10'd11:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d152 =
	      m_vrg_source_ip_11;
      10'd12:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d152 =
	      m_vrg_source_ip_12;
      10'd13:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d152 =
	      m_vrg_source_ip_13;
      10'd14:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d152 =
	      m_vrg_source_ip_14;
      10'd15:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d152 =
	      m_vrg_source_ip_15;
      10'd16:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d152 =
	      m_vrg_source_ip_16;
      default: SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d152 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(source_id__h22093 or
	  m_vvrg_ie_1_0 or
	  m_vvrg_ie_1_1 or
	  m_vvrg_ie_1_2 or
	  m_vvrg_ie_1_3 or
	  m_vvrg_ie_1_4 or
	  m_vvrg_ie_1_5 or
	  m_vvrg_ie_1_6 or
	  m_vvrg_ie_1_7 or
	  m_vvrg_ie_1_8 or
	  m_vvrg_ie_1_9 or
	  m_vvrg_ie_1_10 or
	  m_vvrg_ie_1_11 or
	  m_vvrg_ie_1_12 or
	  m_vvrg_ie_1_13 or
	  m_vvrg_ie_1_14 or m_vvrg_ie_1_15 or m_vvrg_ie_1_16)
  begin
    case (source_id__h22093)
      10'd0:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d402 =
	      m_vvrg_ie_1_0;
      10'd1:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d402 =
	      m_vvrg_ie_1_1;
      10'd2:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d402 =
	      m_vvrg_ie_1_2;
      10'd3:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d402 =
	      m_vvrg_ie_1_3;
      10'd4:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d402 =
	      m_vvrg_ie_1_4;
      10'd5:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d402 =
	      m_vvrg_ie_1_5;
      10'd6:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d402 =
	      m_vvrg_ie_1_6;
      10'd7:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d402 =
	      m_vvrg_ie_1_7;
      10'd8:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d402 =
	      m_vvrg_ie_1_8;
      10'd9:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d402 =
	      m_vvrg_ie_1_9;
      10'd10:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d402 =
	      m_vvrg_ie_1_10;
      10'd11:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d402 =
	      m_vvrg_ie_1_11;
      10'd12:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d402 =
	      m_vvrg_ie_1_12;
      10'd13:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d402 =
	      m_vvrg_ie_1_13;
      10'd14:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d402 =
	      m_vvrg_ie_1_14;
      10'd15:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d402 =
	      m_vvrg_ie_1_15;
      10'd16:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d402 =
	      m_vvrg_ie_1_16;
      default: SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d402 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(source_id__h16920 or
	  m_vrg_source_ip_0 or
	  m_vrg_source_ip_1 or
	  m_vrg_source_ip_2 or
	  m_vrg_source_ip_3 or
	  m_vrg_source_ip_4 or
	  m_vrg_source_ip_5 or
	  m_vrg_source_ip_6 or
	  m_vrg_source_ip_7 or
	  m_vrg_source_ip_8 or
	  m_vrg_source_ip_9 or
	  m_vrg_source_ip_10 or
	  m_vrg_source_ip_11 or
	  m_vrg_source_ip_12 or
	  m_vrg_source_ip_13 or
	  m_vrg_source_ip_14 or m_vrg_source_ip_15 or m_vrg_source_ip_16)
  begin
    case (source_id__h16920)
      10'd0:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d156 =
	      m_vrg_source_ip_0;
      10'd1:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d156 =
	      m_vrg_source_ip_1;
      10'd2:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d156 =
	      m_vrg_source_ip_2;
      10'd3:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d156 =
	      m_vrg_source_ip_3;
      10'd4:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d156 =
	      m_vrg_source_ip_4;
      10'd5:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d156 =
	      m_vrg_source_ip_5;
      10'd6:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d156 =
	      m_vrg_source_ip_6;
      10'd7:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d156 =
	      m_vrg_source_ip_7;
      10'd8:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d156 =
	      m_vrg_source_ip_8;
      10'd9:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d156 =
	      m_vrg_source_ip_9;
      10'd10:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d156 =
	      m_vrg_source_ip_10;
      10'd11:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d156 =
	      m_vrg_source_ip_11;
      10'd12:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d156 =
	      m_vrg_source_ip_12;
      10'd13:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d156 =
	      m_vrg_source_ip_13;
      10'd14:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d156 =
	      m_vrg_source_ip_14;
      10'd15:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d156 =
	      m_vrg_source_ip_15;
      10'd16:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d156 =
	      m_vrg_source_ip_16;
      default: SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d156 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(source_id__h22201 or
	  m_vvrg_ie_0_0 or
	  m_vvrg_ie_0_1 or
	  m_vvrg_ie_0_2 or
	  m_vvrg_ie_0_3 or
	  m_vvrg_ie_0_4 or
	  m_vvrg_ie_0_5 or
	  m_vvrg_ie_0_6 or
	  m_vvrg_ie_0_7 or
	  m_vvrg_ie_0_8 or
	  m_vvrg_ie_0_9 or
	  m_vvrg_ie_0_10 or
	  m_vvrg_ie_0_11 or
	  m_vvrg_ie_0_12 or
	  m_vvrg_ie_0_13 or
	  m_vvrg_ie_0_14 or m_vvrg_ie_0_15 or m_vvrg_ie_0_16)
  begin
    case (source_id__h22201)
      10'd0:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d409 =
	      m_vvrg_ie_0_0;
      10'd1:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d409 =
	      m_vvrg_ie_0_1;
      10'd2:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d409 =
	      m_vvrg_ie_0_2;
      10'd3:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d409 =
	      m_vvrg_ie_0_3;
      10'd4:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d409 =
	      m_vvrg_ie_0_4;
      10'd5:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d409 =
	      m_vvrg_ie_0_5;
      10'd6:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d409 =
	      m_vvrg_ie_0_6;
      10'd7:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d409 =
	      m_vvrg_ie_0_7;
      10'd8:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d409 =
	      m_vvrg_ie_0_8;
      10'd9:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d409 =
	      m_vvrg_ie_0_9;
      10'd10:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d409 =
	      m_vvrg_ie_0_10;
      10'd11:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d409 =
	      m_vvrg_ie_0_11;
      10'd12:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d409 =
	      m_vvrg_ie_0_12;
      10'd13:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d409 =
	      m_vvrg_ie_0_13;
      10'd14:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d409 =
	      m_vvrg_ie_0_14;
      10'd15:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d409 =
	      m_vvrg_ie_0_15;
      10'd16:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d409 =
	      m_vvrg_ie_0_16;
      default: SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d409 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(source_id__h22201 or
	  m_vvrg_ie_1_0 or
	  m_vvrg_ie_1_1 or
	  m_vvrg_ie_1_2 or
	  m_vvrg_ie_1_3 or
	  m_vvrg_ie_1_4 or
	  m_vvrg_ie_1_5 or
	  m_vvrg_ie_1_6 or
	  m_vvrg_ie_1_7 or
	  m_vvrg_ie_1_8 or
	  m_vvrg_ie_1_9 or
	  m_vvrg_ie_1_10 or
	  m_vvrg_ie_1_11 or
	  m_vvrg_ie_1_12 or
	  m_vvrg_ie_1_13 or
	  m_vvrg_ie_1_14 or m_vvrg_ie_1_15 or m_vvrg_ie_1_16)
  begin
    case (source_id__h22201)
      10'd0:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d410 =
	      m_vvrg_ie_1_0;
      10'd1:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d410 =
	      m_vvrg_ie_1_1;
      10'd2:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d410 =
	      m_vvrg_ie_1_2;
      10'd3:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d410 =
	      m_vvrg_ie_1_3;
      10'd4:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d410 =
	      m_vvrg_ie_1_4;
      10'd5:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d410 =
	      m_vvrg_ie_1_5;
      10'd6:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d410 =
	      m_vvrg_ie_1_6;
      10'd7:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d410 =
	      m_vvrg_ie_1_7;
      10'd8:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d410 =
	      m_vvrg_ie_1_8;
      10'd9:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d410 =
	      m_vvrg_ie_1_9;
      10'd10:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d410 =
	      m_vvrg_ie_1_10;
      10'd11:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d410 =
	      m_vvrg_ie_1_11;
      10'd12:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d410 =
	      m_vvrg_ie_1_12;
      10'd13:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d410 =
	      m_vvrg_ie_1_13;
      10'd14:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d410 =
	      m_vvrg_ie_1_14;
      10'd15:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d410 =
	      m_vvrg_ie_1_15;
      10'd16:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d410 =
	      m_vvrg_ie_1_16;
      default: SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d410 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(source_id__h22309 or
	  m_vvrg_ie_0_0 or
	  m_vvrg_ie_0_1 or
	  m_vvrg_ie_0_2 or
	  m_vvrg_ie_0_3 or
	  m_vvrg_ie_0_4 or
	  m_vvrg_ie_0_5 or
	  m_vvrg_ie_0_6 or
	  m_vvrg_ie_0_7 or
	  m_vvrg_ie_0_8 or
	  m_vvrg_ie_0_9 or
	  m_vvrg_ie_0_10 or
	  m_vvrg_ie_0_11 or
	  m_vvrg_ie_0_12 or
	  m_vvrg_ie_0_13 or
	  m_vvrg_ie_0_14 or m_vvrg_ie_0_15 or m_vvrg_ie_0_16)
  begin
    case (source_id__h22309)
      10'd0:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d416 =
	      m_vvrg_ie_0_0;
      10'd1:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d416 =
	      m_vvrg_ie_0_1;
      10'd2:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d416 =
	      m_vvrg_ie_0_2;
      10'd3:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d416 =
	      m_vvrg_ie_0_3;
      10'd4:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d416 =
	      m_vvrg_ie_0_4;
      10'd5:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d416 =
	      m_vvrg_ie_0_5;
      10'd6:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d416 =
	      m_vvrg_ie_0_6;
      10'd7:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d416 =
	      m_vvrg_ie_0_7;
      10'd8:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d416 =
	      m_vvrg_ie_0_8;
      10'd9:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d416 =
	      m_vvrg_ie_0_9;
      10'd10:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d416 =
	      m_vvrg_ie_0_10;
      10'd11:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d416 =
	      m_vvrg_ie_0_11;
      10'd12:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d416 =
	      m_vvrg_ie_0_12;
      10'd13:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d416 =
	      m_vvrg_ie_0_13;
      10'd14:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d416 =
	      m_vvrg_ie_0_14;
      10'd15:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d416 =
	      m_vvrg_ie_0_15;
      10'd16:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d416 =
	      m_vvrg_ie_0_16;
      default: SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d416 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(source_id__h16993 or
	  m_vrg_source_ip_0 or
	  m_vrg_source_ip_1 or
	  m_vrg_source_ip_2 or
	  m_vrg_source_ip_3 or
	  m_vrg_source_ip_4 or
	  m_vrg_source_ip_5 or
	  m_vrg_source_ip_6 or
	  m_vrg_source_ip_7 or
	  m_vrg_source_ip_8 or
	  m_vrg_source_ip_9 or
	  m_vrg_source_ip_10 or
	  m_vrg_source_ip_11 or
	  m_vrg_source_ip_12 or
	  m_vrg_source_ip_13 or
	  m_vrg_source_ip_14 or m_vrg_source_ip_15 or m_vrg_source_ip_16)
  begin
    case (source_id__h16993)
      10'd0:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d161 =
	      m_vrg_source_ip_0;
      10'd1:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d161 =
	      m_vrg_source_ip_1;
      10'd2:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d161 =
	      m_vrg_source_ip_2;
      10'd3:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d161 =
	      m_vrg_source_ip_3;
      10'd4:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d161 =
	      m_vrg_source_ip_4;
      10'd5:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d161 =
	      m_vrg_source_ip_5;
      10'd6:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d161 =
	      m_vrg_source_ip_6;
      10'd7:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d161 =
	      m_vrg_source_ip_7;
      10'd8:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d161 =
	      m_vrg_source_ip_8;
      10'd9:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d161 =
	      m_vrg_source_ip_9;
      10'd10:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d161 =
	      m_vrg_source_ip_10;
      10'd11:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d161 =
	      m_vrg_source_ip_11;
      10'd12:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d161 =
	      m_vrg_source_ip_12;
      10'd13:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d161 =
	      m_vrg_source_ip_13;
      10'd14:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d161 =
	      m_vrg_source_ip_14;
      10'd15:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d161 =
	      m_vrg_source_ip_15;
      10'd16:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d161 =
	      m_vrg_source_ip_16;
      default: SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d161 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(source_id__h22309 or
	  m_vvrg_ie_1_0 or
	  m_vvrg_ie_1_1 or
	  m_vvrg_ie_1_2 or
	  m_vvrg_ie_1_3 or
	  m_vvrg_ie_1_4 or
	  m_vvrg_ie_1_5 or
	  m_vvrg_ie_1_6 or
	  m_vvrg_ie_1_7 or
	  m_vvrg_ie_1_8 or
	  m_vvrg_ie_1_9 or
	  m_vvrg_ie_1_10 or
	  m_vvrg_ie_1_11 or
	  m_vvrg_ie_1_12 or
	  m_vvrg_ie_1_13 or
	  m_vvrg_ie_1_14 or m_vvrg_ie_1_15 or m_vvrg_ie_1_16)
  begin
    case (source_id__h22309)
      10'd0:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d417 =
	      m_vvrg_ie_1_0;
      10'd1:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d417 =
	      m_vvrg_ie_1_1;
      10'd2:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d417 =
	      m_vvrg_ie_1_2;
      10'd3:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d417 =
	      m_vvrg_ie_1_3;
      10'd4:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d417 =
	      m_vvrg_ie_1_4;
      10'd5:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d417 =
	      m_vvrg_ie_1_5;
      10'd6:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d417 =
	      m_vvrg_ie_1_6;
      10'd7:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d417 =
	      m_vvrg_ie_1_7;
      10'd8:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d417 =
	      m_vvrg_ie_1_8;
      10'd9:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d417 =
	      m_vvrg_ie_1_9;
      10'd10:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d417 =
	      m_vvrg_ie_1_10;
      10'd11:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d417 =
	      m_vvrg_ie_1_11;
      10'd12:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d417 =
	      m_vvrg_ie_1_12;
      10'd13:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d417 =
	      m_vvrg_ie_1_13;
      10'd14:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d417 =
	      m_vvrg_ie_1_14;
      10'd15:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d417 =
	      m_vvrg_ie_1_15;
      10'd16:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d417 =
	      m_vvrg_ie_1_16;
      default: SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d417 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(source_id__h17066 or
	  m_vrg_source_ip_0 or
	  m_vrg_source_ip_1 or
	  m_vrg_source_ip_2 or
	  m_vrg_source_ip_3 or
	  m_vrg_source_ip_4 or
	  m_vrg_source_ip_5 or
	  m_vrg_source_ip_6 or
	  m_vrg_source_ip_7 or
	  m_vrg_source_ip_8 or
	  m_vrg_source_ip_9 or
	  m_vrg_source_ip_10 or
	  m_vrg_source_ip_11 or
	  m_vrg_source_ip_12 or
	  m_vrg_source_ip_13 or
	  m_vrg_source_ip_14 or m_vrg_source_ip_15 or m_vrg_source_ip_16)
  begin
    case (source_id__h17066)
      10'd0:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d165 =
	      m_vrg_source_ip_0;
      10'd1:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d165 =
	      m_vrg_source_ip_1;
      10'd2:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d165 =
	      m_vrg_source_ip_2;
      10'd3:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d165 =
	      m_vrg_source_ip_3;
      10'd4:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d165 =
	      m_vrg_source_ip_4;
      10'd5:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d165 =
	      m_vrg_source_ip_5;
      10'd6:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d165 =
	      m_vrg_source_ip_6;
      10'd7:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d165 =
	      m_vrg_source_ip_7;
      10'd8:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d165 =
	      m_vrg_source_ip_8;
      10'd9:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d165 =
	      m_vrg_source_ip_9;
      10'd10:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d165 =
	      m_vrg_source_ip_10;
      10'd11:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d165 =
	      m_vrg_source_ip_11;
      10'd12:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d165 =
	      m_vrg_source_ip_12;
      10'd13:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d165 =
	      m_vrg_source_ip_13;
      10'd14:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d165 =
	      m_vrg_source_ip_14;
      10'd15:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d165 =
	      m_vrg_source_ip_15;
      10'd16:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d165 =
	      m_vrg_source_ip_16;
      default: SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d165 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(source_id__h22417 or
	  m_vvrg_ie_0_0 or
	  m_vvrg_ie_0_1 or
	  m_vvrg_ie_0_2 or
	  m_vvrg_ie_0_3 or
	  m_vvrg_ie_0_4 or
	  m_vvrg_ie_0_5 or
	  m_vvrg_ie_0_6 or
	  m_vvrg_ie_0_7 or
	  m_vvrg_ie_0_8 or
	  m_vvrg_ie_0_9 or
	  m_vvrg_ie_0_10 or
	  m_vvrg_ie_0_11 or
	  m_vvrg_ie_0_12 or
	  m_vvrg_ie_0_13 or
	  m_vvrg_ie_0_14 or m_vvrg_ie_0_15 or m_vvrg_ie_0_16)
  begin
    case (source_id__h22417)
      10'd0:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d424 =
	      m_vvrg_ie_0_0;
      10'd1:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d424 =
	      m_vvrg_ie_0_1;
      10'd2:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d424 =
	      m_vvrg_ie_0_2;
      10'd3:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d424 =
	      m_vvrg_ie_0_3;
      10'd4:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d424 =
	      m_vvrg_ie_0_4;
      10'd5:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d424 =
	      m_vvrg_ie_0_5;
      10'd6:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d424 =
	      m_vvrg_ie_0_6;
      10'd7:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d424 =
	      m_vvrg_ie_0_7;
      10'd8:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d424 =
	      m_vvrg_ie_0_8;
      10'd9:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d424 =
	      m_vvrg_ie_0_9;
      10'd10:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d424 =
	      m_vvrg_ie_0_10;
      10'd11:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d424 =
	      m_vvrg_ie_0_11;
      10'd12:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d424 =
	      m_vvrg_ie_0_12;
      10'd13:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d424 =
	      m_vvrg_ie_0_13;
      10'd14:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d424 =
	      m_vvrg_ie_0_14;
      10'd15:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d424 =
	      m_vvrg_ie_0_15;
      10'd16:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d424 =
	      m_vvrg_ie_0_16;
      default: SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d424 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(source_id__h22417 or
	  m_vvrg_ie_1_0 or
	  m_vvrg_ie_1_1 or
	  m_vvrg_ie_1_2 or
	  m_vvrg_ie_1_3 or
	  m_vvrg_ie_1_4 or
	  m_vvrg_ie_1_5 or
	  m_vvrg_ie_1_6 or
	  m_vvrg_ie_1_7 or
	  m_vvrg_ie_1_8 or
	  m_vvrg_ie_1_9 or
	  m_vvrg_ie_1_10 or
	  m_vvrg_ie_1_11 or
	  m_vvrg_ie_1_12 or
	  m_vvrg_ie_1_13 or
	  m_vvrg_ie_1_14 or m_vvrg_ie_1_15 or m_vvrg_ie_1_16)
  begin
    case (source_id__h22417)
      10'd0:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d425 =
	      m_vvrg_ie_1_0;
      10'd1:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d425 =
	      m_vvrg_ie_1_1;
      10'd2:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d425 =
	      m_vvrg_ie_1_2;
      10'd3:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d425 =
	      m_vvrg_ie_1_3;
      10'd4:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d425 =
	      m_vvrg_ie_1_4;
      10'd5:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d425 =
	      m_vvrg_ie_1_5;
      10'd6:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d425 =
	      m_vvrg_ie_1_6;
      10'd7:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d425 =
	      m_vvrg_ie_1_7;
      10'd8:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d425 =
	      m_vvrg_ie_1_8;
      10'd9:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d425 =
	      m_vvrg_ie_1_9;
      10'd10:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d425 =
	      m_vvrg_ie_1_10;
      10'd11:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d425 =
	      m_vvrg_ie_1_11;
      10'd12:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d425 =
	      m_vvrg_ie_1_12;
      10'd13:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d425 =
	      m_vvrg_ie_1_13;
      10'd14:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d425 =
	      m_vvrg_ie_1_14;
      10'd15:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d425 =
	      m_vvrg_ie_1_15;
      10'd16:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d425 =
	      m_vvrg_ie_1_16;
      default: SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d425 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(source_id__h22525 or
	  m_vvrg_ie_0_0 or
	  m_vvrg_ie_0_1 or
	  m_vvrg_ie_0_2 or
	  m_vvrg_ie_0_3 or
	  m_vvrg_ie_0_4 or
	  m_vvrg_ie_0_5 or
	  m_vvrg_ie_0_6 or
	  m_vvrg_ie_0_7 or
	  m_vvrg_ie_0_8 or
	  m_vvrg_ie_0_9 or
	  m_vvrg_ie_0_10 or
	  m_vvrg_ie_0_11 or
	  m_vvrg_ie_0_12 or
	  m_vvrg_ie_0_13 or
	  m_vvrg_ie_0_14 or m_vvrg_ie_0_15 or m_vvrg_ie_0_16)
  begin
    case (source_id__h22525)
      10'd0:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d431 =
	      m_vvrg_ie_0_0;
      10'd1:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d431 =
	      m_vvrg_ie_0_1;
      10'd2:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d431 =
	      m_vvrg_ie_0_2;
      10'd3:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d431 =
	      m_vvrg_ie_0_3;
      10'd4:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d431 =
	      m_vvrg_ie_0_4;
      10'd5:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d431 =
	      m_vvrg_ie_0_5;
      10'd6:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d431 =
	      m_vvrg_ie_0_6;
      10'd7:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d431 =
	      m_vvrg_ie_0_7;
      10'd8:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d431 =
	      m_vvrg_ie_0_8;
      10'd9:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d431 =
	      m_vvrg_ie_0_9;
      10'd10:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d431 =
	      m_vvrg_ie_0_10;
      10'd11:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d431 =
	      m_vvrg_ie_0_11;
      10'd12:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d431 =
	      m_vvrg_ie_0_12;
      10'd13:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d431 =
	      m_vvrg_ie_0_13;
      10'd14:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d431 =
	      m_vvrg_ie_0_14;
      10'd15:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d431 =
	      m_vvrg_ie_0_15;
      10'd16:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d431 =
	      m_vvrg_ie_0_16;
      default: SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d431 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(source_id__h17139 or
	  m_vrg_source_ip_0 or
	  m_vrg_source_ip_1 or
	  m_vrg_source_ip_2 or
	  m_vrg_source_ip_3 or
	  m_vrg_source_ip_4 or
	  m_vrg_source_ip_5 or
	  m_vrg_source_ip_6 or
	  m_vrg_source_ip_7 or
	  m_vrg_source_ip_8 or
	  m_vrg_source_ip_9 or
	  m_vrg_source_ip_10 or
	  m_vrg_source_ip_11 or
	  m_vrg_source_ip_12 or
	  m_vrg_source_ip_13 or
	  m_vrg_source_ip_14 or m_vrg_source_ip_15 or m_vrg_source_ip_16)
  begin
    case (source_id__h17139)
      10'd0:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d170 =
	      m_vrg_source_ip_0;
      10'd1:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d170 =
	      m_vrg_source_ip_1;
      10'd2:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d170 =
	      m_vrg_source_ip_2;
      10'd3:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d170 =
	      m_vrg_source_ip_3;
      10'd4:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d170 =
	      m_vrg_source_ip_4;
      10'd5:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d170 =
	      m_vrg_source_ip_5;
      10'd6:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d170 =
	      m_vrg_source_ip_6;
      10'd7:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d170 =
	      m_vrg_source_ip_7;
      10'd8:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d170 =
	      m_vrg_source_ip_8;
      10'd9:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d170 =
	      m_vrg_source_ip_9;
      10'd10:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d170 =
	      m_vrg_source_ip_10;
      10'd11:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d170 =
	      m_vrg_source_ip_11;
      10'd12:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d170 =
	      m_vrg_source_ip_12;
      10'd13:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d170 =
	      m_vrg_source_ip_13;
      10'd14:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d170 =
	      m_vrg_source_ip_14;
      10'd15:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d170 =
	      m_vrg_source_ip_15;
      10'd16:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d170 =
	      m_vrg_source_ip_16;
      default: SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d170 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(source_id__h22525 or
	  m_vvrg_ie_1_0 or
	  m_vvrg_ie_1_1 or
	  m_vvrg_ie_1_2 or
	  m_vvrg_ie_1_3 or
	  m_vvrg_ie_1_4 or
	  m_vvrg_ie_1_5 or
	  m_vvrg_ie_1_6 or
	  m_vvrg_ie_1_7 or
	  m_vvrg_ie_1_8 or
	  m_vvrg_ie_1_9 or
	  m_vvrg_ie_1_10 or
	  m_vvrg_ie_1_11 or
	  m_vvrg_ie_1_12 or
	  m_vvrg_ie_1_13 or
	  m_vvrg_ie_1_14 or m_vvrg_ie_1_15 or m_vvrg_ie_1_16)
  begin
    case (source_id__h22525)
      10'd0:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d432 =
	      m_vvrg_ie_1_0;
      10'd1:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d432 =
	      m_vvrg_ie_1_1;
      10'd2:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d432 =
	      m_vvrg_ie_1_2;
      10'd3:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d432 =
	      m_vvrg_ie_1_3;
      10'd4:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d432 =
	      m_vvrg_ie_1_4;
      10'd5:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d432 =
	      m_vvrg_ie_1_5;
      10'd6:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d432 =
	      m_vvrg_ie_1_6;
      10'd7:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d432 =
	      m_vvrg_ie_1_7;
      10'd8:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d432 =
	      m_vvrg_ie_1_8;
      10'd9:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d432 =
	      m_vvrg_ie_1_9;
      10'd10:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d432 =
	      m_vvrg_ie_1_10;
      10'd11:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d432 =
	      m_vvrg_ie_1_11;
      10'd12:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d432 =
	      m_vvrg_ie_1_12;
      10'd13:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d432 =
	      m_vvrg_ie_1_13;
      10'd14:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d432 =
	      m_vvrg_ie_1_14;
      10'd15:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d432 =
	      m_vvrg_ie_1_15;
      10'd16:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d432 =
	      m_vvrg_ie_1_16;
      default: SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d432 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(source_id__h17212 or
	  m_vrg_source_ip_0 or
	  m_vrg_source_ip_1 or
	  m_vrg_source_ip_2 or
	  m_vrg_source_ip_3 or
	  m_vrg_source_ip_4 or
	  m_vrg_source_ip_5 or
	  m_vrg_source_ip_6 or
	  m_vrg_source_ip_7 or
	  m_vrg_source_ip_8 or
	  m_vrg_source_ip_9 or
	  m_vrg_source_ip_10 or
	  m_vrg_source_ip_11 or
	  m_vrg_source_ip_12 or
	  m_vrg_source_ip_13 or
	  m_vrg_source_ip_14 or m_vrg_source_ip_15 or m_vrg_source_ip_16)
  begin
    case (source_id__h17212)
      10'd0:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d174 =
	      m_vrg_source_ip_0;
      10'd1:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d174 =
	      m_vrg_source_ip_1;
      10'd2:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d174 =
	      m_vrg_source_ip_2;
      10'd3:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d174 =
	      m_vrg_source_ip_3;
      10'd4:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d174 =
	      m_vrg_source_ip_4;
      10'd5:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d174 =
	      m_vrg_source_ip_5;
      10'd6:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d174 =
	      m_vrg_source_ip_6;
      10'd7:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d174 =
	      m_vrg_source_ip_7;
      10'd8:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d174 =
	      m_vrg_source_ip_8;
      10'd9:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d174 =
	      m_vrg_source_ip_9;
      10'd10:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d174 =
	      m_vrg_source_ip_10;
      10'd11:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d174 =
	      m_vrg_source_ip_11;
      10'd12:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d174 =
	      m_vrg_source_ip_12;
      10'd13:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d174 =
	      m_vrg_source_ip_13;
      10'd14:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d174 =
	      m_vrg_source_ip_14;
      10'd15:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d174 =
	      m_vrg_source_ip_15;
      10'd16:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d174 =
	      m_vrg_source_ip_16;
      default: SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d174 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(source_id__h22633 or
	  m_vvrg_ie_0_0 or
	  m_vvrg_ie_0_1 or
	  m_vvrg_ie_0_2 or
	  m_vvrg_ie_0_3 or
	  m_vvrg_ie_0_4 or
	  m_vvrg_ie_0_5 or
	  m_vvrg_ie_0_6 or
	  m_vvrg_ie_0_7 or
	  m_vvrg_ie_0_8 or
	  m_vvrg_ie_0_9 or
	  m_vvrg_ie_0_10 or
	  m_vvrg_ie_0_11 or
	  m_vvrg_ie_0_12 or
	  m_vvrg_ie_0_13 or
	  m_vvrg_ie_0_14 or m_vvrg_ie_0_15 or m_vvrg_ie_0_16)
  begin
    case (source_id__h22633)
      10'd0:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d439 =
	      m_vvrg_ie_0_0;
      10'd1:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d439 =
	      m_vvrg_ie_0_1;
      10'd2:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d439 =
	      m_vvrg_ie_0_2;
      10'd3:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d439 =
	      m_vvrg_ie_0_3;
      10'd4:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d439 =
	      m_vvrg_ie_0_4;
      10'd5:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d439 =
	      m_vvrg_ie_0_5;
      10'd6:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d439 =
	      m_vvrg_ie_0_6;
      10'd7:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d439 =
	      m_vvrg_ie_0_7;
      10'd8:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d439 =
	      m_vvrg_ie_0_8;
      10'd9:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d439 =
	      m_vvrg_ie_0_9;
      10'd10:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d439 =
	      m_vvrg_ie_0_10;
      10'd11:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d439 =
	      m_vvrg_ie_0_11;
      10'd12:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d439 =
	      m_vvrg_ie_0_12;
      10'd13:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d439 =
	      m_vvrg_ie_0_13;
      10'd14:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d439 =
	      m_vvrg_ie_0_14;
      10'd15:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d439 =
	      m_vvrg_ie_0_15;
      10'd16:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d439 =
	      m_vvrg_ie_0_16;
      default: SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d439 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(source_id__h22633 or
	  m_vvrg_ie_1_0 or
	  m_vvrg_ie_1_1 or
	  m_vvrg_ie_1_2 or
	  m_vvrg_ie_1_3 or
	  m_vvrg_ie_1_4 or
	  m_vvrg_ie_1_5 or
	  m_vvrg_ie_1_6 or
	  m_vvrg_ie_1_7 or
	  m_vvrg_ie_1_8 or
	  m_vvrg_ie_1_9 or
	  m_vvrg_ie_1_10 or
	  m_vvrg_ie_1_11 or
	  m_vvrg_ie_1_12 or
	  m_vvrg_ie_1_13 or
	  m_vvrg_ie_1_14 or m_vvrg_ie_1_15 or m_vvrg_ie_1_16)
  begin
    case (source_id__h22633)
      10'd0:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d440 =
	      m_vvrg_ie_1_0;
      10'd1:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d440 =
	      m_vvrg_ie_1_1;
      10'd2:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d440 =
	      m_vvrg_ie_1_2;
      10'd3:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d440 =
	      m_vvrg_ie_1_3;
      10'd4:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d440 =
	      m_vvrg_ie_1_4;
      10'd5:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d440 =
	      m_vvrg_ie_1_5;
      10'd6:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d440 =
	      m_vvrg_ie_1_6;
      10'd7:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d440 =
	      m_vvrg_ie_1_7;
      10'd8:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d440 =
	      m_vvrg_ie_1_8;
      10'd9:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d440 =
	      m_vvrg_ie_1_9;
      10'd10:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d440 =
	      m_vvrg_ie_1_10;
      10'd11:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d440 =
	      m_vvrg_ie_1_11;
      10'd12:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d440 =
	      m_vvrg_ie_1_12;
      10'd13:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d440 =
	      m_vvrg_ie_1_13;
      10'd14:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d440 =
	      m_vvrg_ie_1_14;
      10'd15:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d440 =
	      m_vvrg_ie_1_15;
      10'd16:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d440 =
	      m_vvrg_ie_1_16;
      default: SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d440 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(source_id__h22741 or
	  m_vvrg_ie_0_0 or
	  m_vvrg_ie_0_1 or
	  m_vvrg_ie_0_2 or
	  m_vvrg_ie_0_3 or
	  m_vvrg_ie_0_4 or
	  m_vvrg_ie_0_5 or
	  m_vvrg_ie_0_6 or
	  m_vvrg_ie_0_7 or
	  m_vvrg_ie_0_8 or
	  m_vvrg_ie_0_9 or
	  m_vvrg_ie_0_10 or
	  m_vvrg_ie_0_11 or
	  m_vvrg_ie_0_12 or
	  m_vvrg_ie_0_13 or
	  m_vvrg_ie_0_14 or m_vvrg_ie_0_15 or m_vvrg_ie_0_16)
  begin
    case (source_id__h22741)
      10'd0:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d446 =
	      m_vvrg_ie_0_0;
      10'd1:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d446 =
	      m_vvrg_ie_0_1;
      10'd2:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d446 =
	      m_vvrg_ie_0_2;
      10'd3:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d446 =
	      m_vvrg_ie_0_3;
      10'd4:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d446 =
	      m_vvrg_ie_0_4;
      10'd5:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d446 =
	      m_vvrg_ie_0_5;
      10'd6:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d446 =
	      m_vvrg_ie_0_6;
      10'd7:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d446 =
	      m_vvrg_ie_0_7;
      10'd8:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d446 =
	      m_vvrg_ie_0_8;
      10'd9:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d446 =
	      m_vvrg_ie_0_9;
      10'd10:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d446 =
	      m_vvrg_ie_0_10;
      10'd11:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d446 =
	      m_vvrg_ie_0_11;
      10'd12:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d446 =
	      m_vvrg_ie_0_12;
      10'd13:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d446 =
	      m_vvrg_ie_0_13;
      10'd14:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d446 =
	      m_vvrg_ie_0_14;
      10'd15:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d446 =
	      m_vvrg_ie_0_15;
      10'd16:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d446 =
	      m_vvrg_ie_0_16;
      default: SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d446 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(source_id__h17285 or
	  m_vrg_source_ip_0 or
	  m_vrg_source_ip_1 or
	  m_vrg_source_ip_2 or
	  m_vrg_source_ip_3 or
	  m_vrg_source_ip_4 or
	  m_vrg_source_ip_5 or
	  m_vrg_source_ip_6 or
	  m_vrg_source_ip_7 or
	  m_vrg_source_ip_8 or
	  m_vrg_source_ip_9 or
	  m_vrg_source_ip_10 or
	  m_vrg_source_ip_11 or
	  m_vrg_source_ip_12 or
	  m_vrg_source_ip_13 or
	  m_vrg_source_ip_14 or m_vrg_source_ip_15 or m_vrg_source_ip_16)
  begin
    case (source_id__h17285)
      10'd0:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d179 =
	      m_vrg_source_ip_0;
      10'd1:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d179 =
	      m_vrg_source_ip_1;
      10'd2:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d179 =
	      m_vrg_source_ip_2;
      10'd3:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d179 =
	      m_vrg_source_ip_3;
      10'd4:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d179 =
	      m_vrg_source_ip_4;
      10'd5:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d179 =
	      m_vrg_source_ip_5;
      10'd6:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d179 =
	      m_vrg_source_ip_6;
      10'd7:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d179 =
	      m_vrg_source_ip_7;
      10'd8:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d179 =
	      m_vrg_source_ip_8;
      10'd9:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d179 =
	      m_vrg_source_ip_9;
      10'd10:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d179 =
	      m_vrg_source_ip_10;
      10'd11:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d179 =
	      m_vrg_source_ip_11;
      10'd12:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d179 =
	      m_vrg_source_ip_12;
      10'd13:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d179 =
	      m_vrg_source_ip_13;
      10'd14:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d179 =
	      m_vrg_source_ip_14;
      10'd15:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d179 =
	      m_vrg_source_ip_15;
      10'd16:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d179 =
	      m_vrg_source_ip_16;
      default: SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d179 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(source_id__h22741 or
	  m_vvrg_ie_1_0 or
	  m_vvrg_ie_1_1 or
	  m_vvrg_ie_1_2 or
	  m_vvrg_ie_1_3 or
	  m_vvrg_ie_1_4 or
	  m_vvrg_ie_1_5 or
	  m_vvrg_ie_1_6 or
	  m_vvrg_ie_1_7 or
	  m_vvrg_ie_1_8 or
	  m_vvrg_ie_1_9 or
	  m_vvrg_ie_1_10 or
	  m_vvrg_ie_1_11 or
	  m_vvrg_ie_1_12 or
	  m_vvrg_ie_1_13 or
	  m_vvrg_ie_1_14 or m_vvrg_ie_1_15 or m_vvrg_ie_1_16)
  begin
    case (source_id__h22741)
      10'd0:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d447 =
	      m_vvrg_ie_1_0;
      10'd1:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d447 =
	      m_vvrg_ie_1_1;
      10'd2:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d447 =
	      m_vvrg_ie_1_2;
      10'd3:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d447 =
	      m_vvrg_ie_1_3;
      10'd4:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d447 =
	      m_vvrg_ie_1_4;
      10'd5:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d447 =
	      m_vvrg_ie_1_5;
      10'd6:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d447 =
	      m_vvrg_ie_1_6;
      10'd7:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d447 =
	      m_vvrg_ie_1_7;
      10'd8:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d447 =
	      m_vvrg_ie_1_8;
      10'd9:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d447 =
	      m_vvrg_ie_1_9;
      10'd10:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d447 =
	      m_vvrg_ie_1_10;
      10'd11:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d447 =
	      m_vvrg_ie_1_11;
      10'd12:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d447 =
	      m_vvrg_ie_1_12;
      10'd13:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d447 =
	      m_vvrg_ie_1_13;
      10'd14:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d447 =
	      m_vvrg_ie_1_14;
      10'd15:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d447 =
	      m_vvrg_ie_1_15;
      10'd16:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d447 =
	      m_vvrg_ie_1_16;
      default: SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d447 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(source_id__h22849 or
	  m_vvrg_ie_0_0 or
	  m_vvrg_ie_0_1 or
	  m_vvrg_ie_0_2 or
	  m_vvrg_ie_0_3 or
	  m_vvrg_ie_0_4 or
	  m_vvrg_ie_0_5 or
	  m_vvrg_ie_0_6 or
	  m_vvrg_ie_0_7 or
	  m_vvrg_ie_0_8 or
	  m_vvrg_ie_0_9 or
	  m_vvrg_ie_0_10 or
	  m_vvrg_ie_0_11 or
	  m_vvrg_ie_0_12 or
	  m_vvrg_ie_0_13 or
	  m_vvrg_ie_0_14 or m_vvrg_ie_0_15 or m_vvrg_ie_0_16)
  begin
    case (source_id__h22849)
      10'd0:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d454 =
	      m_vvrg_ie_0_0;
      10'd1:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d454 =
	      m_vvrg_ie_0_1;
      10'd2:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d454 =
	      m_vvrg_ie_0_2;
      10'd3:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d454 =
	      m_vvrg_ie_0_3;
      10'd4:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d454 =
	      m_vvrg_ie_0_4;
      10'd5:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d454 =
	      m_vvrg_ie_0_5;
      10'd6:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d454 =
	      m_vvrg_ie_0_6;
      10'd7:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d454 =
	      m_vvrg_ie_0_7;
      10'd8:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d454 =
	      m_vvrg_ie_0_8;
      10'd9:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d454 =
	      m_vvrg_ie_0_9;
      10'd10:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d454 =
	      m_vvrg_ie_0_10;
      10'd11:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d454 =
	      m_vvrg_ie_0_11;
      10'd12:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d454 =
	      m_vvrg_ie_0_12;
      10'd13:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d454 =
	      m_vvrg_ie_0_13;
      10'd14:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d454 =
	      m_vvrg_ie_0_14;
      10'd15:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d454 =
	      m_vvrg_ie_0_15;
      10'd16:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d454 =
	      m_vvrg_ie_0_16;
      default: SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d454 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(source_id__h22849 or
	  m_vvrg_ie_1_0 or
	  m_vvrg_ie_1_1 or
	  m_vvrg_ie_1_2 or
	  m_vvrg_ie_1_3 or
	  m_vvrg_ie_1_4 or
	  m_vvrg_ie_1_5 or
	  m_vvrg_ie_1_6 or
	  m_vvrg_ie_1_7 or
	  m_vvrg_ie_1_8 or
	  m_vvrg_ie_1_9 or
	  m_vvrg_ie_1_10 or
	  m_vvrg_ie_1_11 or
	  m_vvrg_ie_1_12 or
	  m_vvrg_ie_1_13 or
	  m_vvrg_ie_1_14 or m_vvrg_ie_1_15 or m_vvrg_ie_1_16)
  begin
    case (source_id__h22849)
      10'd0:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d455 =
	      m_vvrg_ie_1_0;
      10'd1:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d455 =
	      m_vvrg_ie_1_1;
      10'd2:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d455 =
	      m_vvrg_ie_1_2;
      10'd3:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d455 =
	      m_vvrg_ie_1_3;
      10'd4:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d455 =
	      m_vvrg_ie_1_4;
      10'd5:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d455 =
	      m_vvrg_ie_1_5;
      10'd6:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d455 =
	      m_vvrg_ie_1_6;
      10'd7:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d455 =
	      m_vvrg_ie_1_7;
      10'd8:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d455 =
	      m_vvrg_ie_1_8;
      10'd9:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d455 =
	      m_vvrg_ie_1_9;
      10'd10:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d455 =
	      m_vvrg_ie_1_10;
      10'd11:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d455 =
	      m_vvrg_ie_1_11;
      10'd12:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d455 =
	      m_vvrg_ie_1_12;
      10'd13:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d455 =
	      m_vvrg_ie_1_13;
      10'd14:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d455 =
	      m_vvrg_ie_1_14;
      10'd15:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d455 =
	      m_vvrg_ie_1_15;
      10'd16:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d455 =
	      m_vvrg_ie_1_16;
      default: SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d455 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(source_id__h22957 or
	  m_vvrg_ie_0_0 or
	  m_vvrg_ie_0_1 or
	  m_vvrg_ie_0_2 or
	  m_vvrg_ie_0_3 or
	  m_vvrg_ie_0_4 or
	  m_vvrg_ie_0_5 or
	  m_vvrg_ie_0_6 or
	  m_vvrg_ie_0_7 or
	  m_vvrg_ie_0_8 or
	  m_vvrg_ie_0_9 or
	  m_vvrg_ie_0_10 or
	  m_vvrg_ie_0_11 or
	  m_vvrg_ie_0_12 or
	  m_vvrg_ie_0_13 or
	  m_vvrg_ie_0_14 or m_vvrg_ie_0_15 or m_vvrg_ie_0_16)
  begin
    case (source_id__h22957)
      10'd0:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d461 =
	      m_vvrg_ie_0_0;
      10'd1:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d461 =
	      m_vvrg_ie_0_1;
      10'd2:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d461 =
	      m_vvrg_ie_0_2;
      10'd3:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d461 =
	      m_vvrg_ie_0_3;
      10'd4:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d461 =
	      m_vvrg_ie_0_4;
      10'd5:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d461 =
	      m_vvrg_ie_0_5;
      10'd6:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d461 =
	      m_vvrg_ie_0_6;
      10'd7:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d461 =
	      m_vvrg_ie_0_7;
      10'd8:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d461 =
	      m_vvrg_ie_0_8;
      10'd9:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d461 =
	      m_vvrg_ie_0_9;
      10'd10:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d461 =
	      m_vvrg_ie_0_10;
      10'd11:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d461 =
	      m_vvrg_ie_0_11;
      10'd12:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d461 =
	      m_vvrg_ie_0_12;
      10'd13:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d461 =
	      m_vvrg_ie_0_13;
      10'd14:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d461 =
	      m_vvrg_ie_0_14;
      10'd15:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d461 =
	      m_vvrg_ie_0_15;
      10'd16:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d461 =
	      m_vvrg_ie_0_16;
      default: SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d461 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(source_id__h17431 or
	  m_vrg_source_ip_0 or
	  m_vrg_source_ip_1 or
	  m_vrg_source_ip_2 or
	  m_vrg_source_ip_3 or
	  m_vrg_source_ip_4 or
	  m_vrg_source_ip_5 or
	  m_vrg_source_ip_6 or
	  m_vrg_source_ip_7 or
	  m_vrg_source_ip_8 or
	  m_vrg_source_ip_9 or
	  m_vrg_source_ip_10 or
	  m_vrg_source_ip_11 or
	  m_vrg_source_ip_12 or
	  m_vrg_source_ip_13 or
	  m_vrg_source_ip_14 or m_vrg_source_ip_15 or m_vrg_source_ip_16)
  begin
    case (source_id__h17431)
      10'd0:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d188 =
	      m_vrg_source_ip_0;
      10'd1:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d188 =
	      m_vrg_source_ip_1;
      10'd2:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d188 =
	      m_vrg_source_ip_2;
      10'd3:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d188 =
	      m_vrg_source_ip_3;
      10'd4:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d188 =
	      m_vrg_source_ip_4;
      10'd5:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d188 =
	      m_vrg_source_ip_5;
      10'd6:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d188 =
	      m_vrg_source_ip_6;
      10'd7:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d188 =
	      m_vrg_source_ip_7;
      10'd8:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d188 =
	      m_vrg_source_ip_8;
      10'd9:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d188 =
	      m_vrg_source_ip_9;
      10'd10:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d188 =
	      m_vrg_source_ip_10;
      10'd11:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d188 =
	      m_vrg_source_ip_11;
      10'd12:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d188 =
	      m_vrg_source_ip_12;
      10'd13:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d188 =
	      m_vrg_source_ip_13;
      10'd14:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d188 =
	      m_vrg_source_ip_14;
      10'd15:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d188 =
	      m_vrg_source_ip_15;
      10'd16:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d188 =
	      m_vrg_source_ip_16;
      default: SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d188 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(source_id__h22957 or
	  m_vvrg_ie_1_0 or
	  m_vvrg_ie_1_1 or
	  m_vvrg_ie_1_2 or
	  m_vvrg_ie_1_3 or
	  m_vvrg_ie_1_4 or
	  m_vvrg_ie_1_5 or
	  m_vvrg_ie_1_6 or
	  m_vvrg_ie_1_7 or
	  m_vvrg_ie_1_8 or
	  m_vvrg_ie_1_9 or
	  m_vvrg_ie_1_10 or
	  m_vvrg_ie_1_11 or
	  m_vvrg_ie_1_12 or
	  m_vvrg_ie_1_13 or
	  m_vvrg_ie_1_14 or m_vvrg_ie_1_15 or m_vvrg_ie_1_16)
  begin
    case (source_id__h22957)
      10'd0:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d462 =
	      m_vvrg_ie_1_0;
      10'd1:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d462 =
	      m_vvrg_ie_1_1;
      10'd2:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d462 =
	      m_vvrg_ie_1_2;
      10'd3:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d462 =
	      m_vvrg_ie_1_3;
      10'd4:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d462 =
	      m_vvrg_ie_1_4;
      10'd5:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d462 =
	      m_vvrg_ie_1_5;
      10'd6:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d462 =
	      m_vvrg_ie_1_6;
      10'd7:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d462 =
	      m_vvrg_ie_1_7;
      10'd8:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d462 =
	      m_vvrg_ie_1_8;
      10'd9:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d462 =
	      m_vvrg_ie_1_9;
      10'd10:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d462 =
	      m_vvrg_ie_1_10;
      10'd11:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d462 =
	      m_vvrg_ie_1_11;
      10'd12:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d462 =
	      m_vvrg_ie_1_12;
      10'd13:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d462 =
	      m_vvrg_ie_1_13;
      10'd14:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d462 =
	      m_vvrg_ie_1_14;
      10'd15:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d462 =
	      m_vvrg_ie_1_15;
      10'd16:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d462 =
	      m_vvrg_ie_1_16;
      default: SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d462 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(source_id__h17504 or
	  m_vrg_source_ip_0 or
	  m_vrg_source_ip_1 or
	  m_vrg_source_ip_2 or
	  m_vrg_source_ip_3 or
	  m_vrg_source_ip_4 or
	  m_vrg_source_ip_5 or
	  m_vrg_source_ip_6 or
	  m_vrg_source_ip_7 or
	  m_vrg_source_ip_8 or
	  m_vrg_source_ip_9 or
	  m_vrg_source_ip_10 or
	  m_vrg_source_ip_11 or
	  m_vrg_source_ip_12 or
	  m_vrg_source_ip_13 or
	  m_vrg_source_ip_14 or m_vrg_source_ip_15 or m_vrg_source_ip_16)
  begin
    case (source_id__h17504)
      10'd0:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d192 =
	      m_vrg_source_ip_0;
      10'd1:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d192 =
	      m_vrg_source_ip_1;
      10'd2:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d192 =
	      m_vrg_source_ip_2;
      10'd3:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d192 =
	      m_vrg_source_ip_3;
      10'd4:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d192 =
	      m_vrg_source_ip_4;
      10'd5:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d192 =
	      m_vrg_source_ip_5;
      10'd6:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d192 =
	      m_vrg_source_ip_6;
      10'd7:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d192 =
	      m_vrg_source_ip_7;
      10'd8:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d192 =
	      m_vrg_source_ip_8;
      10'd9:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d192 =
	      m_vrg_source_ip_9;
      10'd10:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d192 =
	      m_vrg_source_ip_10;
      10'd11:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d192 =
	      m_vrg_source_ip_11;
      10'd12:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d192 =
	      m_vrg_source_ip_12;
      10'd13:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d192 =
	      m_vrg_source_ip_13;
      10'd14:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d192 =
	      m_vrg_source_ip_14;
      10'd15:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d192 =
	      m_vrg_source_ip_15;
      10'd16:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d192 =
	      m_vrg_source_ip_16;
      default: SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d192 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(source_id__h23065 or
	  m_vvrg_ie_0_0 or
	  m_vvrg_ie_0_1 or
	  m_vvrg_ie_0_2 or
	  m_vvrg_ie_0_3 or
	  m_vvrg_ie_0_4 or
	  m_vvrg_ie_0_5 or
	  m_vvrg_ie_0_6 or
	  m_vvrg_ie_0_7 or
	  m_vvrg_ie_0_8 or
	  m_vvrg_ie_0_9 or
	  m_vvrg_ie_0_10 or
	  m_vvrg_ie_0_11 or
	  m_vvrg_ie_0_12 or
	  m_vvrg_ie_0_13 or
	  m_vvrg_ie_0_14 or m_vvrg_ie_0_15 or m_vvrg_ie_0_16)
  begin
    case (source_id__h23065)
      10'd0:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d469 =
	      m_vvrg_ie_0_0;
      10'd1:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d469 =
	      m_vvrg_ie_0_1;
      10'd2:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d469 =
	      m_vvrg_ie_0_2;
      10'd3:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d469 =
	      m_vvrg_ie_0_3;
      10'd4:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d469 =
	      m_vvrg_ie_0_4;
      10'd5:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d469 =
	      m_vvrg_ie_0_5;
      10'd6:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d469 =
	      m_vvrg_ie_0_6;
      10'd7:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d469 =
	      m_vvrg_ie_0_7;
      10'd8:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d469 =
	      m_vvrg_ie_0_8;
      10'd9:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d469 =
	      m_vvrg_ie_0_9;
      10'd10:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d469 =
	      m_vvrg_ie_0_10;
      10'd11:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d469 =
	      m_vvrg_ie_0_11;
      10'd12:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d469 =
	      m_vvrg_ie_0_12;
      10'd13:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d469 =
	      m_vvrg_ie_0_13;
      10'd14:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d469 =
	      m_vvrg_ie_0_14;
      10'd15:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d469 =
	      m_vvrg_ie_0_15;
      10'd16:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d469 =
	      m_vvrg_ie_0_16;
      default: SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d469 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(source_id__h23065 or
	  m_vvrg_ie_1_0 or
	  m_vvrg_ie_1_1 or
	  m_vvrg_ie_1_2 or
	  m_vvrg_ie_1_3 or
	  m_vvrg_ie_1_4 or
	  m_vvrg_ie_1_5 or
	  m_vvrg_ie_1_6 or
	  m_vvrg_ie_1_7 or
	  m_vvrg_ie_1_8 or
	  m_vvrg_ie_1_9 or
	  m_vvrg_ie_1_10 or
	  m_vvrg_ie_1_11 or
	  m_vvrg_ie_1_12 or
	  m_vvrg_ie_1_13 or
	  m_vvrg_ie_1_14 or m_vvrg_ie_1_15 or m_vvrg_ie_1_16)
  begin
    case (source_id__h23065)
      10'd0:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d470 =
	      m_vvrg_ie_1_0;
      10'd1:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d470 =
	      m_vvrg_ie_1_1;
      10'd2:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d470 =
	      m_vvrg_ie_1_2;
      10'd3:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d470 =
	      m_vvrg_ie_1_3;
      10'd4:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d470 =
	      m_vvrg_ie_1_4;
      10'd5:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d470 =
	      m_vvrg_ie_1_5;
      10'd6:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d470 =
	      m_vvrg_ie_1_6;
      10'd7:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d470 =
	      m_vvrg_ie_1_7;
      10'd8:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d470 =
	      m_vvrg_ie_1_8;
      10'd9:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d470 =
	      m_vvrg_ie_1_9;
      10'd10:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d470 =
	      m_vvrg_ie_1_10;
      10'd11:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d470 =
	      m_vvrg_ie_1_11;
      10'd12:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d470 =
	      m_vvrg_ie_1_12;
      10'd13:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d470 =
	      m_vvrg_ie_1_13;
      10'd14:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d470 =
	      m_vvrg_ie_1_14;
      10'd15:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d470 =
	      m_vvrg_ie_1_15;
      10'd16:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d470 =
	      m_vvrg_ie_1_16;
      default: SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d470 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(source_id__h23173 or
	  m_vvrg_ie_0_0 or
	  m_vvrg_ie_0_1 or
	  m_vvrg_ie_0_2 or
	  m_vvrg_ie_0_3 or
	  m_vvrg_ie_0_4 or
	  m_vvrg_ie_0_5 or
	  m_vvrg_ie_0_6 or
	  m_vvrg_ie_0_7 or
	  m_vvrg_ie_0_8 or
	  m_vvrg_ie_0_9 or
	  m_vvrg_ie_0_10 or
	  m_vvrg_ie_0_11 or
	  m_vvrg_ie_0_12 or
	  m_vvrg_ie_0_13 or
	  m_vvrg_ie_0_14 or m_vvrg_ie_0_15 or m_vvrg_ie_0_16)
  begin
    case (source_id__h23173)
      10'd0:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d476 =
	      m_vvrg_ie_0_0;
      10'd1:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d476 =
	      m_vvrg_ie_0_1;
      10'd2:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d476 =
	      m_vvrg_ie_0_2;
      10'd3:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d476 =
	      m_vvrg_ie_0_3;
      10'd4:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d476 =
	      m_vvrg_ie_0_4;
      10'd5:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d476 =
	      m_vvrg_ie_0_5;
      10'd6:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d476 =
	      m_vvrg_ie_0_6;
      10'd7:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d476 =
	      m_vvrg_ie_0_7;
      10'd8:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d476 =
	      m_vvrg_ie_0_8;
      10'd9:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d476 =
	      m_vvrg_ie_0_9;
      10'd10:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d476 =
	      m_vvrg_ie_0_10;
      10'd11:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d476 =
	      m_vvrg_ie_0_11;
      10'd12:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d476 =
	      m_vvrg_ie_0_12;
      10'd13:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d476 =
	      m_vvrg_ie_0_13;
      10'd14:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d476 =
	      m_vvrg_ie_0_14;
      10'd15:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d476 =
	      m_vvrg_ie_0_15;
      10'd16:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d476 =
	      m_vvrg_ie_0_16;
      default: SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d476 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(source_id__h17577 or
	  m_vrg_source_ip_0 or
	  m_vrg_source_ip_1 or
	  m_vrg_source_ip_2 or
	  m_vrg_source_ip_3 or
	  m_vrg_source_ip_4 or
	  m_vrg_source_ip_5 or
	  m_vrg_source_ip_6 or
	  m_vrg_source_ip_7 or
	  m_vrg_source_ip_8 or
	  m_vrg_source_ip_9 or
	  m_vrg_source_ip_10 or
	  m_vrg_source_ip_11 or
	  m_vrg_source_ip_12 or
	  m_vrg_source_ip_13 or
	  m_vrg_source_ip_14 or m_vrg_source_ip_15 or m_vrg_source_ip_16)
  begin
    case (source_id__h17577)
      10'd0:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d197 =
	      m_vrg_source_ip_0;
      10'd1:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d197 =
	      m_vrg_source_ip_1;
      10'd2:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d197 =
	      m_vrg_source_ip_2;
      10'd3:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d197 =
	      m_vrg_source_ip_3;
      10'd4:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d197 =
	      m_vrg_source_ip_4;
      10'd5:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d197 =
	      m_vrg_source_ip_5;
      10'd6:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d197 =
	      m_vrg_source_ip_6;
      10'd7:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d197 =
	      m_vrg_source_ip_7;
      10'd8:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d197 =
	      m_vrg_source_ip_8;
      10'd9:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d197 =
	      m_vrg_source_ip_9;
      10'd10:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d197 =
	      m_vrg_source_ip_10;
      10'd11:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d197 =
	      m_vrg_source_ip_11;
      10'd12:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d197 =
	      m_vrg_source_ip_12;
      10'd13:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d197 =
	      m_vrg_source_ip_13;
      10'd14:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d197 =
	      m_vrg_source_ip_14;
      10'd15:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d197 =
	      m_vrg_source_ip_15;
      10'd16:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d197 =
	      m_vrg_source_ip_16;
      default: SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d197 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(source_id__h23173 or
	  m_vvrg_ie_1_0 or
	  m_vvrg_ie_1_1 or
	  m_vvrg_ie_1_2 or
	  m_vvrg_ie_1_3 or
	  m_vvrg_ie_1_4 or
	  m_vvrg_ie_1_5 or
	  m_vvrg_ie_1_6 or
	  m_vvrg_ie_1_7 or
	  m_vvrg_ie_1_8 or
	  m_vvrg_ie_1_9 or
	  m_vvrg_ie_1_10 or
	  m_vvrg_ie_1_11 or
	  m_vvrg_ie_1_12 or
	  m_vvrg_ie_1_13 or
	  m_vvrg_ie_1_14 or m_vvrg_ie_1_15 or m_vvrg_ie_1_16)
  begin
    case (source_id__h23173)
      10'd0:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d477 =
	      m_vvrg_ie_1_0;
      10'd1:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d477 =
	      m_vvrg_ie_1_1;
      10'd2:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d477 =
	      m_vvrg_ie_1_2;
      10'd3:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d477 =
	      m_vvrg_ie_1_3;
      10'd4:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d477 =
	      m_vvrg_ie_1_4;
      10'd5:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d477 =
	      m_vvrg_ie_1_5;
      10'd6:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d477 =
	      m_vvrg_ie_1_6;
      10'd7:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d477 =
	      m_vvrg_ie_1_7;
      10'd8:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d477 =
	      m_vvrg_ie_1_8;
      10'd9:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d477 =
	      m_vvrg_ie_1_9;
      10'd10:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d477 =
	      m_vvrg_ie_1_10;
      10'd11:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d477 =
	      m_vvrg_ie_1_11;
      10'd12:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d477 =
	      m_vvrg_ie_1_12;
      10'd13:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d477 =
	      m_vvrg_ie_1_13;
      10'd14:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d477 =
	      m_vvrg_ie_1_14;
      10'd15:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d477 =
	      m_vvrg_ie_1_15;
      10'd16:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d477 =
	      m_vvrg_ie_1_16;
      default: SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d477 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(source_id__h17650 or
	  m_vrg_source_ip_0 or
	  m_vrg_source_ip_1 or
	  m_vrg_source_ip_2 or
	  m_vrg_source_ip_3 or
	  m_vrg_source_ip_4 or
	  m_vrg_source_ip_5 or
	  m_vrg_source_ip_6 or
	  m_vrg_source_ip_7 or
	  m_vrg_source_ip_8 or
	  m_vrg_source_ip_9 or
	  m_vrg_source_ip_10 or
	  m_vrg_source_ip_11 or
	  m_vrg_source_ip_12 or
	  m_vrg_source_ip_13 or
	  m_vrg_source_ip_14 or m_vrg_source_ip_15 or m_vrg_source_ip_16)
  begin
    case (source_id__h17650)
      10'd0:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d201 =
	      m_vrg_source_ip_0;
      10'd1:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d201 =
	      m_vrg_source_ip_1;
      10'd2:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d201 =
	      m_vrg_source_ip_2;
      10'd3:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d201 =
	      m_vrg_source_ip_3;
      10'd4:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d201 =
	      m_vrg_source_ip_4;
      10'd5:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d201 =
	      m_vrg_source_ip_5;
      10'd6:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d201 =
	      m_vrg_source_ip_6;
      10'd7:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d201 =
	      m_vrg_source_ip_7;
      10'd8:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d201 =
	      m_vrg_source_ip_8;
      10'd9:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d201 =
	      m_vrg_source_ip_9;
      10'd10:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d201 =
	      m_vrg_source_ip_10;
      10'd11:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d201 =
	      m_vrg_source_ip_11;
      10'd12:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d201 =
	      m_vrg_source_ip_12;
      10'd13:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d201 =
	      m_vrg_source_ip_13;
      10'd14:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d201 =
	      m_vrg_source_ip_14;
      10'd15:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d201 =
	      m_vrg_source_ip_15;
      10'd16:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d201 =
	      m_vrg_source_ip_16;
      default: SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d201 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(source_id__h23281 or
	  m_vvrg_ie_1_0 or
	  m_vvrg_ie_1_1 or
	  m_vvrg_ie_1_2 or
	  m_vvrg_ie_1_3 or
	  m_vvrg_ie_1_4 or
	  m_vvrg_ie_1_5 or
	  m_vvrg_ie_1_6 or
	  m_vvrg_ie_1_7 or
	  m_vvrg_ie_1_8 or
	  m_vvrg_ie_1_9 or
	  m_vvrg_ie_1_10 or
	  m_vvrg_ie_1_11 or
	  m_vvrg_ie_1_12 or
	  m_vvrg_ie_1_13 or
	  m_vvrg_ie_1_14 or m_vvrg_ie_1_15 or m_vvrg_ie_1_16)
  begin
    case (source_id__h23281)
      10'd0:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d485 =
	      m_vvrg_ie_1_0;
      10'd1:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d485 =
	      m_vvrg_ie_1_1;
      10'd2:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d485 =
	      m_vvrg_ie_1_2;
      10'd3:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d485 =
	      m_vvrg_ie_1_3;
      10'd4:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d485 =
	      m_vvrg_ie_1_4;
      10'd5:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d485 =
	      m_vvrg_ie_1_5;
      10'd6:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d485 =
	      m_vvrg_ie_1_6;
      10'd7:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d485 =
	      m_vvrg_ie_1_7;
      10'd8:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d485 =
	      m_vvrg_ie_1_8;
      10'd9:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d485 =
	      m_vvrg_ie_1_9;
      10'd10:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d485 =
	      m_vvrg_ie_1_10;
      10'd11:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d485 =
	      m_vvrg_ie_1_11;
      10'd12:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d485 =
	      m_vvrg_ie_1_12;
      10'd13:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d485 =
	      m_vvrg_ie_1_13;
      10'd14:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d485 =
	      m_vvrg_ie_1_14;
      10'd15:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d485 =
	      m_vvrg_ie_1_15;
      10'd16:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d485 =
	      m_vvrg_ie_1_16;
      default: SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d485 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(source_id__h23281 or
	  m_vvrg_ie_0_0 or
	  m_vvrg_ie_0_1 or
	  m_vvrg_ie_0_2 or
	  m_vvrg_ie_0_3 or
	  m_vvrg_ie_0_4 or
	  m_vvrg_ie_0_5 or
	  m_vvrg_ie_0_6 or
	  m_vvrg_ie_0_7 or
	  m_vvrg_ie_0_8 or
	  m_vvrg_ie_0_9 or
	  m_vvrg_ie_0_10 or
	  m_vvrg_ie_0_11 or
	  m_vvrg_ie_0_12 or
	  m_vvrg_ie_0_13 or
	  m_vvrg_ie_0_14 or m_vvrg_ie_0_15 or m_vvrg_ie_0_16)
  begin
    case (source_id__h23281)
      10'd0:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d484 =
	      m_vvrg_ie_0_0;
      10'd1:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d484 =
	      m_vvrg_ie_0_1;
      10'd2:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d484 =
	      m_vvrg_ie_0_2;
      10'd3:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d484 =
	      m_vvrg_ie_0_3;
      10'd4:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d484 =
	      m_vvrg_ie_0_4;
      10'd5:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d484 =
	      m_vvrg_ie_0_5;
      10'd6:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d484 =
	      m_vvrg_ie_0_6;
      10'd7:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d484 =
	      m_vvrg_ie_0_7;
      10'd8:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d484 =
	      m_vvrg_ie_0_8;
      10'd9:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d484 =
	      m_vvrg_ie_0_9;
      10'd10:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d484 =
	      m_vvrg_ie_0_10;
      10'd11:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d484 =
	      m_vvrg_ie_0_11;
      10'd12:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d484 =
	      m_vvrg_ie_0_12;
      10'd13:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d484 =
	      m_vvrg_ie_0_13;
      10'd14:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d484 =
	      m_vvrg_ie_0_14;
      10'd15:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d484 =
	      m_vvrg_ie_0_15;
      10'd16:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d484 =
	      m_vvrg_ie_0_16;
      default: SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d484 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(source_id__h23389 or
	  m_vvrg_ie_0_0 or
	  m_vvrg_ie_0_1 or
	  m_vvrg_ie_0_2 or
	  m_vvrg_ie_0_3 or
	  m_vvrg_ie_0_4 or
	  m_vvrg_ie_0_5 or
	  m_vvrg_ie_0_6 or
	  m_vvrg_ie_0_7 or
	  m_vvrg_ie_0_8 or
	  m_vvrg_ie_0_9 or
	  m_vvrg_ie_0_10 or
	  m_vvrg_ie_0_11 or
	  m_vvrg_ie_0_12 or
	  m_vvrg_ie_0_13 or
	  m_vvrg_ie_0_14 or m_vvrg_ie_0_15 or m_vvrg_ie_0_16)
  begin
    case (source_id__h23389)
      10'd0:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d491 =
	      m_vvrg_ie_0_0;
      10'd1:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d491 =
	      m_vvrg_ie_0_1;
      10'd2:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d491 =
	      m_vvrg_ie_0_2;
      10'd3:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d491 =
	      m_vvrg_ie_0_3;
      10'd4:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d491 =
	      m_vvrg_ie_0_4;
      10'd5:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d491 =
	      m_vvrg_ie_0_5;
      10'd6:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d491 =
	      m_vvrg_ie_0_6;
      10'd7:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d491 =
	      m_vvrg_ie_0_7;
      10'd8:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d491 =
	      m_vvrg_ie_0_8;
      10'd9:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d491 =
	      m_vvrg_ie_0_9;
      10'd10:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d491 =
	      m_vvrg_ie_0_10;
      10'd11:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d491 =
	      m_vvrg_ie_0_11;
      10'd12:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d491 =
	      m_vvrg_ie_0_12;
      10'd13:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d491 =
	      m_vvrg_ie_0_13;
      10'd14:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d491 =
	      m_vvrg_ie_0_14;
      10'd15:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d491 =
	      m_vvrg_ie_0_15;
      10'd16:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d491 =
	      m_vvrg_ie_0_16;
      default: SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d491 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(source_id__h17723 or
	  m_vrg_source_ip_0 or
	  m_vrg_source_ip_1 or
	  m_vrg_source_ip_2 or
	  m_vrg_source_ip_3 or
	  m_vrg_source_ip_4 or
	  m_vrg_source_ip_5 or
	  m_vrg_source_ip_6 or
	  m_vrg_source_ip_7 or
	  m_vrg_source_ip_8 or
	  m_vrg_source_ip_9 or
	  m_vrg_source_ip_10 or
	  m_vrg_source_ip_11 or
	  m_vrg_source_ip_12 or
	  m_vrg_source_ip_13 or
	  m_vrg_source_ip_14 or m_vrg_source_ip_15 or m_vrg_source_ip_16)
  begin
    case (source_id__h17723)
      10'd0:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d206 =
	      m_vrg_source_ip_0;
      10'd1:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d206 =
	      m_vrg_source_ip_1;
      10'd2:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d206 =
	      m_vrg_source_ip_2;
      10'd3:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d206 =
	      m_vrg_source_ip_3;
      10'd4:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d206 =
	      m_vrg_source_ip_4;
      10'd5:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d206 =
	      m_vrg_source_ip_5;
      10'd6:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d206 =
	      m_vrg_source_ip_6;
      10'd7:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d206 =
	      m_vrg_source_ip_7;
      10'd8:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d206 =
	      m_vrg_source_ip_8;
      10'd9:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d206 =
	      m_vrg_source_ip_9;
      10'd10:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d206 =
	      m_vrg_source_ip_10;
      10'd11:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d206 =
	      m_vrg_source_ip_11;
      10'd12:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d206 =
	      m_vrg_source_ip_12;
      10'd13:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d206 =
	      m_vrg_source_ip_13;
      10'd14:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d206 =
	      m_vrg_source_ip_14;
      10'd15:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d206 =
	      m_vrg_source_ip_15;
      10'd16:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d206 =
	      m_vrg_source_ip_16;
      default: SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d206 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(source_id__h23389 or
	  m_vvrg_ie_1_0 or
	  m_vvrg_ie_1_1 or
	  m_vvrg_ie_1_2 or
	  m_vvrg_ie_1_3 or
	  m_vvrg_ie_1_4 or
	  m_vvrg_ie_1_5 or
	  m_vvrg_ie_1_6 or
	  m_vvrg_ie_1_7 or
	  m_vvrg_ie_1_8 or
	  m_vvrg_ie_1_9 or
	  m_vvrg_ie_1_10 or
	  m_vvrg_ie_1_11 or
	  m_vvrg_ie_1_12 or
	  m_vvrg_ie_1_13 or
	  m_vvrg_ie_1_14 or m_vvrg_ie_1_15 or m_vvrg_ie_1_16)
  begin
    case (source_id__h23389)
      10'd0:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d492 =
	      m_vvrg_ie_1_0;
      10'd1:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d492 =
	      m_vvrg_ie_1_1;
      10'd2:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d492 =
	      m_vvrg_ie_1_2;
      10'd3:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d492 =
	      m_vvrg_ie_1_3;
      10'd4:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d492 =
	      m_vvrg_ie_1_4;
      10'd5:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d492 =
	      m_vvrg_ie_1_5;
      10'd6:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d492 =
	      m_vvrg_ie_1_6;
      10'd7:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d492 =
	      m_vvrg_ie_1_7;
      10'd8:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d492 =
	      m_vvrg_ie_1_8;
      10'd9:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d492 =
	      m_vvrg_ie_1_9;
      10'd10:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d492 =
	      m_vvrg_ie_1_10;
      10'd11:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d492 =
	      m_vvrg_ie_1_11;
      10'd12:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d492 =
	      m_vvrg_ie_1_12;
      10'd13:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d492 =
	      m_vvrg_ie_1_13;
      10'd14:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d492 =
	      m_vvrg_ie_1_14;
      10'd15:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d492 =
	      m_vvrg_ie_1_15;
      10'd16:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d492 =
	      m_vvrg_ie_1_16;
      default: SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d492 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(source_id__h17796 or
	  m_vrg_source_ip_0 or
	  m_vrg_source_ip_1 or
	  m_vrg_source_ip_2 or
	  m_vrg_source_ip_3 or
	  m_vrg_source_ip_4 or
	  m_vrg_source_ip_5 or
	  m_vrg_source_ip_6 or
	  m_vrg_source_ip_7 or
	  m_vrg_source_ip_8 or
	  m_vrg_source_ip_9 or
	  m_vrg_source_ip_10 or
	  m_vrg_source_ip_11 or
	  m_vrg_source_ip_12 or
	  m_vrg_source_ip_13 or
	  m_vrg_source_ip_14 or m_vrg_source_ip_15 or m_vrg_source_ip_16)
  begin
    case (source_id__h17796)
      10'd0:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d210 =
	      m_vrg_source_ip_0;
      10'd1:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d210 =
	      m_vrg_source_ip_1;
      10'd2:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d210 =
	      m_vrg_source_ip_2;
      10'd3:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d210 =
	      m_vrg_source_ip_3;
      10'd4:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d210 =
	      m_vrg_source_ip_4;
      10'd5:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d210 =
	      m_vrg_source_ip_5;
      10'd6:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d210 =
	      m_vrg_source_ip_6;
      10'd7:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d210 =
	      m_vrg_source_ip_7;
      10'd8:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d210 =
	      m_vrg_source_ip_8;
      10'd9:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d210 =
	      m_vrg_source_ip_9;
      10'd10:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d210 =
	      m_vrg_source_ip_10;
      10'd11:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d210 =
	      m_vrg_source_ip_11;
      10'd12:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d210 =
	      m_vrg_source_ip_12;
      10'd13:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d210 =
	      m_vrg_source_ip_13;
      10'd14:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d210 =
	      m_vrg_source_ip_14;
      10'd15:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d210 =
	      m_vrg_source_ip_15;
      10'd16:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d210 =
	      m_vrg_source_ip_16;
      default: SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d210 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(source_id__h23497 or
	  m_vvrg_ie_0_0 or
	  m_vvrg_ie_0_1 or
	  m_vvrg_ie_0_2 or
	  m_vvrg_ie_0_3 or
	  m_vvrg_ie_0_4 or
	  m_vvrg_ie_0_5 or
	  m_vvrg_ie_0_6 or
	  m_vvrg_ie_0_7 or
	  m_vvrg_ie_0_8 or
	  m_vvrg_ie_0_9 or
	  m_vvrg_ie_0_10 or
	  m_vvrg_ie_0_11 or
	  m_vvrg_ie_0_12 or
	  m_vvrg_ie_0_13 or
	  m_vvrg_ie_0_14 or m_vvrg_ie_0_15 or m_vvrg_ie_0_16)
  begin
    case (source_id__h23497)
      10'd0:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d499 =
	      m_vvrg_ie_0_0;
      10'd1:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d499 =
	      m_vvrg_ie_0_1;
      10'd2:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d499 =
	      m_vvrg_ie_0_2;
      10'd3:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d499 =
	      m_vvrg_ie_0_3;
      10'd4:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d499 =
	      m_vvrg_ie_0_4;
      10'd5:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d499 =
	      m_vvrg_ie_0_5;
      10'd6:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d499 =
	      m_vvrg_ie_0_6;
      10'd7:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d499 =
	      m_vvrg_ie_0_7;
      10'd8:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d499 =
	      m_vvrg_ie_0_8;
      10'd9:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d499 =
	      m_vvrg_ie_0_9;
      10'd10:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d499 =
	      m_vvrg_ie_0_10;
      10'd11:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d499 =
	      m_vvrg_ie_0_11;
      10'd12:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d499 =
	      m_vvrg_ie_0_12;
      10'd13:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d499 =
	      m_vvrg_ie_0_13;
      10'd14:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d499 =
	      m_vvrg_ie_0_14;
      10'd15:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d499 =
	      m_vvrg_ie_0_15;
      10'd16:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d499 =
	      m_vvrg_ie_0_16;
      default: SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d499 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(source_id__h23497 or
	  m_vvrg_ie_1_0 or
	  m_vvrg_ie_1_1 or
	  m_vvrg_ie_1_2 or
	  m_vvrg_ie_1_3 or
	  m_vvrg_ie_1_4 or
	  m_vvrg_ie_1_5 or
	  m_vvrg_ie_1_6 or
	  m_vvrg_ie_1_7 or
	  m_vvrg_ie_1_8 or
	  m_vvrg_ie_1_9 or
	  m_vvrg_ie_1_10 or
	  m_vvrg_ie_1_11 or
	  m_vvrg_ie_1_12 or
	  m_vvrg_ie_1_13 or
	  m_vvrg_ie_1_14 or m_vvrg_ie_1_15 or m_vvrg_ie_1_16)
  begin
    case (source_id__h23497)
      10'd0:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d500 =
	      m_vvrg_ie_1_0;
      10'd1:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d500 =
	      m_vvrg_ie_1_1;
      10'd2:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d500 =
	      m_vvrg_ie_1_2;
      10'd3:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d500 =
	      m_vvrg_ie_1_3;
      10'd4:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d500 =
	      m_vvrg_ie_1_4;
      10'd5:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d500 =
	      m_vvrg_ie_1_5;
      10'd6:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d500 =
	      m_vvrg_ie_1_6;
      10'd7:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d500 =
	      m_vvrg_ie_1_7;
      10'd8:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d500 =
	      m_vvrg_ie_1_8;
      10'd9:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d500 =
	      m_vvrg_ie_1_9;
      10'd10:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d500 =
	      m_vvrg_ie_1_10;
      10'd11:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d500 =
	      m_vvrg_ie_1_11;
      10'd12:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d500 =
	      m_vvrg_ie_1_12;
      10'd13:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d500 =
	      m_vvrg_ie_1_13;
      10'd14:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d500 =
	      m_vvrg_ie_1_14;
      10'd15:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d500 =
	      m_vvrg_ie_1_15;
      10'd16:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d500 =
	      m_vvrg_ie_1_16;
      default: SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d500 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(source_id__h23605 or
	  m_vvrg_ie_0_0 or
	  m_vvrg_ie_0_1 or
	  m_vvrg_ie_0_2 or
	  m_vvrg_ie_0_3 or
	  m_vvrg_ie_0_4 or
	  m_vvrg_ie_0_5 or
	  m_vvrg_ie_0_6 or
	  m_vvrg_ie_0_7 or
	  m_vvrg_ie_0_8 or
	  m_vvrg_ie_0_9 or
	  m_vvrg_ie_0_10 or
	  m_vvrg_ie_0_11 or
	  m_vvrg_ie_0_12 or
	  m_vvrg_ie_0_13 or
	  m_vvrg_ie_0_14 or m_vvrg_ie_0_15 or m_vvrg_ie_0_16)
  begin
    case (source_id__h23605)
      10'd0:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d506 =
	      m_vvrg_ie_0_0;
      10'd1:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d506 =
	      m_vvrg_ie_0_1;
      10'd2:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d506 =
	      m_vvrg_ie_0_2;
      10'd3:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d506 =
	      m_vvrg_ie_0_3;
      10'd4:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d506 =
	      m_vvrg_ie_0_4;
      10'd5:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d506 =
	      m_vvrg_ie_0_5;
      10'd6:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d506 =
	      m_vvrg_ie_0_6;
      10'd7:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d506 =
	      m_vvrg_ie_0_7;
      10'd8:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d506 =
	      m_vvrg_ie_0_8;
      10'd9:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d506 =
	      m_vvrg_ie_0_9;
      10'd10:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d506 =
	      m_vvrg_ie_0_10;
      10'd11:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d506 =
	      m_vvrg_ie_0_11;
      10'd12:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d506 =
	      m_vvrg_ie_0_12;
      10'd13:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d506 =
	      m_vvrg_ie_0_13;
      10'd14:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d506 =
	      m_vvrg_ie_0_14;
      10'd15:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d506 =
	      m_vvrg_ie_0_15;
      10'd16:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d506 =
	      m_vvrg_ie_0_16;
      default: SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d506 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(source_id__h17869 or
	  m_vrg_source_ip_0 or
	  m_vrg_source_ip_1 or
	  m_vrg_source_ip_2 or
	  m_vrg_source_ip_3 or
	  m_vrg_source_ip_4 or
	  m_vrg_source_ip_5 or
	  m_vrg_source_ip_6 or
	  m_vrg_source_ip_7 or
	  m_vrg_source_ip_8 or
	  m_vrg_source_ip_9 or
	  m_vrg_source_ip_10 or
	  m_vrg_source_ip_11 or
	  m_vrg_source_ip_12 or
	  m_vrg_source_ip_13 or
	  m_vrg_source_ip_14 or m_vrg_source_ip_15 or m_vrg_source_ip_16)
  begin
    case (source_id__h17869)
      10'd0:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d215 =
	      m_vrg_source_ip_0;
      10'd1:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d215 =
	      m_vrg_source_ip_1;
      10'd2:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d215 =
	      m_vrg_source_ip_2;
      10'd3:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d215 =
	      m_vrg_source_ip_3;
      10'd4:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d215 =
	      m_vrg_source_ip_4;
      10'd5:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d215 =
	      m_vrg_source_ip_5;
      10'd6:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d215 =
	      m_vrg_source_ip_6;
      10'd7:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d215 =
	      m_vrg_source_ip_7;
      10'd8:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d215 =
	      m_vrg_source_ip_8;
      10'd9:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d215 =
	      m_vrg_source_ip_9;
      10'd10:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d215 =
	      m_vrg_source_ip_10;
      10'd11:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d215 =
	      m_vrg_source_ip_11;
      10'd12:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d215 =
	      m_vrg_source_ip_12;
      10'd13:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d215 =
	      m_vrg_source_ip_13;
      10'd14:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d215 =
	      m_vrg_source_ip_14;
      10'd15:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d215 =
	      m_vrg_source_ip_15;
      10'd16:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d215 =
	      m_vrg_source_ip_16;
      default: SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d215 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(source_id__h23605 or
	  m_vvrg_ie_1_0 or
	  m_vvrg_ie_1_1 or
	  m_vvrg_ie_1_2 or
	  m_vvrg_ie_1_3 or
	  m_vvrg_ie_1_4 or
	  m_vvrg_ie_1_5 or
	  m_vvrg_ie_1_6 or
	  m_vvrg_ie_1_7 or
	  m_vvrg_ie_1_8 or
	  m_vvrg_ie_1_9 or
	  m_vvrg_ie_1_10 or
	  m_vvrg_ie_1_11 or
	  m_vvrg_ie_1_12 or
	  m_vvrg_ie_1_13 or
	  m_vvrg_ie_1_14 or m_vvrg_ie_1_15 or m_vvrg_ie_1_16)
  begin
    case (source_id__h23605)
      10'd0:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d507 =
	      m_vvrg_ie_1_0;
      10'd1:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d507 =
	      m_vvrg_ie_1_1;
      10'd2:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d507 =
	      m_vvrg_ie_1_2;
      10'd3:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d507 =
	      m_vvrg_ie_1_3;
      10'd4:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d507 =
	      m_vvrg_ie_1_4;
      10'd5:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d507 =
	      m_vvrg_ie_1_5;
      10'd6:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d507 =
	      m_vvrg_ie_1_6;
      10'd7:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d507 =
	      m_vvrg_ie_1_7;
      10'd8:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d507 =
	      m_vvrg_ie_1_8;
      10'd9:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d507 =
	      m_vvrg_ie_1_9;
      10'd10:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d507 =
	      m_vvrg_ie_1_10;
      10'd11:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d507 =
	      m_vvrg_ie_1_11;
      10'd12:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d507 =
	      m_vvrg_ie_1_12;
      10'd13:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d507 =
	      m_vvrg_ie_1_13;
      10'd14:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d507 =
	      m_vvrg_ie_1_14;
      10'd15:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d507 =
	      m_vvrg_ie_1_15;
      10'd16:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d507 =
	      m_vvrg_ie_1_16;
      default: SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d507 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(source_id__h17942 or
	  m_vrg_source_ip_0 or
	  m_vrg_source_ip_1 or
	  m_vrg_source_ip_2 or
	  m_vrg_source_ip_3 or
	  m_vrg_source_ip_4 or
	  m_vrg_source_ip_5 or
	  m_vrg_source_ip_6 or
	  m_vrg_source_ip_7 or
	  m_vrg_source_ip_8 or
	  m_vrg_source_ip_9 or
	  m_vrg_source_ip_10 or
	  m_vrg_source_ip_11 or
	  m_vrg_source_ip_12 or
	  m_vrg_source_ip_13 or
	  m_vrg_source_ip_14 or m_vrg_source_ip_15 or m_vrg_source_ip_16)
  begin
    case (source_id__h17942)
      10'd0:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d219 =
	      m_vrg_source_ip_0;
      10'd1:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d219 =
	      m_vrg_source_ip_1;
      10'd2:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d219 =
	      m_vrg_source_ip_2;
      10'd3:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d219 =
	      m_vrg_source_ip_3;
      10'd4:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d219 =
	      m_vrg_source_ip_4;
      10'd5:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d219 =
	      m_vrg_source_ip_5;
      10'd6:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d219 =
	      m_vrg_source_ip_6;
      10'd7:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d219 =
	      m_vrg_source_ip_7;
      10'd8:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d219 =
	      m_vrg_source_ip_8;
      10'd9:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d219 =
	      m_vrg_source_ip_9;
      10'd10:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d219 =
	      m_vrg_source_ip_10;
      10'd11:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d219 =
	      m_vrg_source_ip_11;
      10'd12:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d219 =
	      m_vrg_source_ip_12;
      10'd13:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d219 =
	      m_vrg_source_ip_13;
      10'd14:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d219 =
	      m_vrg_source_ip_14;
      10'd15:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d219 =
	      m_vrg_source_ip_15;
      10'd16:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d219 =
	      m_vrg_source_ip_16;
      default: SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d219 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(source_id__h23713 or
	  m_vvrg_ie_0_0 or
	  m_vvrg_ie_0_1 or
	  m_vvrg_ie_0_2 or
	  m_vvrg_ie_0_3 or
	  m_vvrg_ie_0_4 or
	  m_vvrg_ie_0_5 or
	  m_vvrg_ie_0_6 or
	  m_vvrg_ie_0_7 or
	  m_vvrg_ie_0_8 or
	  m_vvrg_ie_0_9 or
	  m_vvrg_ie_0_10 or
	  m_vvrg_ie_0_11 or
	  m_vvrg_ie_0_12 or
	  m_vvrg_ie_0_13 or
	  m_vvrg_ie_0_14 or m_vvrg_ie_0_15 or m_vvrg_ie_0_16)
  begin
    case (source_id__h23713)
      10'd0:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d514 =
	      m_vvrg_ie_0_0;
      10'd1:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d514 =
	      m_vvrg_ie_0_1;
      10'd2:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d514 =
	      m_vvrg_ie_0_2;
      10'd3:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d514 =
	      m_vvrg_ie_0_3;
      10'd4:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d514 =
	      m_vvrg_ie_0_4;
      10'd5:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d514 =
	      m_vvrg_ie_0_5;
      10'd6:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d514 =
	      m_vvrg_ie_0_6;
      10'd7:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d514 =
	      m_vvrg_ie_0_7;
      10'd8:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d514 =
	      m_vvrg_ie_0_8;
      10'd9:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d514 =
	      m_vvrg_ie_0_9;
      10'd10:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d514 =
	      m_vvrg_ie_0_10;
      10'd11:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d514 =
	      m_vvrg_ie_0_11;
      10'd12:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d514 =
	      m_vvrg_ie_0_12;
      10'd13:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d514 =
	      m_vvrg_ie_0_13;
      10'd14:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d514 =
	      m_vvrg_ie_0_14;
      10'd15:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d514 =
	      m_vvrg_ie_0_15;
      10'd16:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d514 =
	      m_vvrg_ie_0_16;
      default: SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d514 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(source_id__h23713 or
	  m_vvrg_ie_1_0 or
	  m_vvrg_ie_1_1 or
	  m_vvrg_ie_1_2 or
	  m_vvrg_ie_1_3 or
	  m_vvrg_ie_1_4 or
	  m_vvrg_ie_1_5 or
	  m_vvrg_ie_1_6 or
	  m_vvrg_ie_1_7 or
	  m_vvrg_ie_1_8 or
	  m_vvrg_ie_1_9 or
	  m_vvrg_ie_1_10 or
	  m_vvrg_ie_1_11 or
	  m_vvrg_ie_1_12 or
	  m_vvrg_ie_1_13 or
	  m_vvrg_ie_1_14 or m_vvrg_ie_1_15 or m_vvrg_ie_1_16)
  begin
    case (source_id__h23713)
      10'd0:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d515 =
	      m_vvrg_ie_1_0;
      10'd1:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d515 =
	      m_vvrg_ie_1_1;
      10'd2:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d515 =
	      m_vvrg_ie_1_2;
      10'd3:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d515 =
	      m_vvrg_ie_1_3;
      10'd4:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d515 =
	      m_vvrg_ie_1_4;
      10'd5:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d515 =
	      m_vvrg_ie_1_5;
      10'd6:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d515 =
	      m_vvrg_ie_1_6;
      10'd7:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d515 =
	      m_vvrg_ie_1_7;
      10'd8:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d515 =
	      m_vvrg_ie_1_8;
      10'd9:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d515 =
	      m_vvrg_ie_1_9;
      10'd10:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d515 =
	      m_vvrg_ie_1_10;
      10'd11:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d515 =
	      m_vvrg_ie_1_11;
      10'd12:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d515 =
	      m_vvrg_ie_1_12;
      10'd13:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d515 =
	      m_vvrg_ie_1_13;
      10'd14:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d515 =
	      m_vvrg_ie_1_14;
      10'd15:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d515 =
	      m_vvrg_ie_1_15;
      10'd16:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d515 =
	      m_vvrg_ie_1_16;
      default: SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d515 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(source_id_base__h13893 or
	  m_vvrg_ie_0_0 or
	  m_vvrg_ie_0_1 or
	  m_vvrg_ie_0_2 or
	  m_vvrg_ie_0_3 or
	  m_vvrg_ie_0_4 or
	  m_vvrg_ie_0_5 or
	  m_vvrg_ie_0_6 or
	  m_vvrg_ie_0_7 or
	  m_vvrg_ie_0_8 or
	  m_vvrg_ie_0_9 or
	  m_vvrg_ie_0_10 or
	  m_vvrg_ie_0_11 or
	  m_vvrg_ie_0_12 or
	  m_vvrg_ie_0_13 or
	  m_vvrg_ie_0_14 or m_vvrg_ie_0_15 or m_vvrg_ie_0_16)
  begin
    case (source_id_base__h13893)
      10'd0:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d519 =
	      m_vvrg_ie_0_0;
      10'd1:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d519 =
	      m_vvrg_ie_0_1;
      10'd2:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d519 =
	      m_vvrg_ie_0_2;
      10'd3:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d519 =
	      m_vvrg_ie_0_3;
      10'd4:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d519 =
	      m_vvrg_ie_0_4;
      10'd5:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d519 =
	      m_vvrg_ie_0_5;
      10'd6:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d519 =
	      m_vvrg_ie_0_6;
      10'd7:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d519 =
	      m_vvrg_ie_0_7;
      10'd8:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d519 =
	      m_vvrg_ie_0_8;
      10'd9:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d519 =
	      m_vvrg_ie_0_9;
      10'd10:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d519 =
	      m_vvrg_ie_0_10;
      10'd11:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d519 =
	      m_vvrg_ie_0_11;
      10'd12:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d519 =
	      m_vvrg_ie_0_12;
      10'd13:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d519 =
	      m_vvrg_ie_0_13;
      10'd14:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d519 =
	      m_vvrg_ie_0_14;
      10'd15:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d519 =
	      m_vvrg_ie_0_15;
      10'd16:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d519 =
	      m_vvrg_ie_0_16;
      default: SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d519 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(source_id__h18015 or
	  m_vrg_source_ip_0 or
	  m_vrg_source_ip_1 or
	  m_vrg_source_ip_2 or
	  m_vrg_source_ip_3 or
	  m_vrg_source_ip_4 or
	  m_vrg_source_ip_5 or
	  m_vrg_source_ip_6 or
	  m_vrg_source_ip_7 or
	  m_vrg_source_ip_8 or
	  m_vrg_source_ip_9 or
	  m_vrg_source_ip_10 or
	  m_vrg_source_ip_11 or
	  m_vrg_source_ip_12 or
	  m_vrg_source_ip_13 or
	  m_vrg_source_ip_14 or m_vrg_source_ip_15 or m_vrg_source_ip_16)
  begin
    case (source_id__h18015)
      10'd0:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d224 =
	      m_vrg_source_ip_0;
      10'd1:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d224 =
	      m_vrg_source_ip_1;
      10'd2:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d224 =
	      m_vrg_source_ip_2;
      10'd3:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d224 =
	      m_vrg_source_ip_3;
      10'd4:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d224 =
	      m_vrg_source_ip_4;
      10'd5:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d224 =
	      m_vrg_source_ip_5;
      10'd6:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d224 =
	      m_vrg_source_ip_6;
      10'd7:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d224 =
	      m_vrg_source_ip_7;
      10'd8:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d224 =
	      m_vrg_source_ip_8;
      10'd9:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d224 =
	      m_vrg_source_ip_9;
      10'd10:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d224 =
	      m_vrg_source_ip_10;
      10'd11:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d224 =
	      m_vrg_source_ip_11;
      10'd12:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d224 =
	      m_vrg_source_ip_12;
      10'd13:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d224 =
	      m_vrg_source_ip_13;
      10'd14:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d224 =
	      m_vrg_source_ip_14;
      10'd15:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d224 =
	      m_vrg_source_ip_15;
      10'd16:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d224 =
	      m_vrg_source_ip_16;
      default: SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d224 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(source_id_base__h13893 or
	  m_vvrg_ie_1_0 or
	  m_vvrg_ie_1_1 or
	  m_vvrg_ie_1_2 or
	  m_vvrg_ie_1_3 or
	  m_vvrg_ie_1_4 or
	  m_vvrg_ie_1_5 or
	  m_vvrg_ie_1_6 or
	  m_vvrg_ie_1_7 or
	  m_vvrg_ie_1_8 or
	  m_vvrg_ie_1_9 or
	  m_vvrg_ie_1_10 or
	  m_vvrg_ie_1_11 or
	  m_vvrg_ie_1_12 or
	  m_vvrg_ie_1_13 or
	  m_vvrg_ie_1_14 or m_vvrg_ie_1_15 or m_vvrg_ie_1_16)
  begin
    case (source_id_base__h13893)
      10'd0:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d520 =
	      m_vvrg_ie_1_0;
      10'd1:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d520 =
	      m_vvrg_ie_1_1;
      10'd2:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d520 =
	      m_vvrg_ie_1_2;
      10'd3:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d520 =
	      m_vvrg_ie_1_3;
      10'd4:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d520 =
	      m_vvrg_ie_1_4;
      10'd5:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d520 =
	      m_vvrg_ie_1_5;
      10'd6:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d520 =
	      m_vvrg_ie_1_6;
      10'd7:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d520 =
	      m_vvrg_ie_1_7;
      10'd8:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d520 =
	      m_vvrg_ie_1_8;
      10'd9:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d520 =
	      m_vvrg_ie_1_9;
      10'd10:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d520 =
	      m_vvrg_ie_1_10;
      10'd11:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d520 =
	      m_vvrg_ie_1_11;
      10'd12:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d520 =
	      m_vvrg_ie_1_12;
      10'd13:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d520 =
	      m_vvrg_ie_1_13;
      10'd14:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d520 =
	      m_vvrg_ie_1_14;
      10'd15:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d520 =
	      m_vvrg_ie_1_15;
      10'd16:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d520 =
	      m_vvrg_ie_1_16;
      default: SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d520 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(addr_offset__h13465 or
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d271 or
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d290)
  begin
    case (addr_offset__h13465[11:7])
      5'd0:
	  CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q1 =
	      SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d271;
      5'd1:
	  CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q1 =
	      SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d290;
      default: CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q1 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(addr_offset__h13465 or
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d296 or
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d297)
  begin
    case (addr_offset__h13465[11:7])
      5'd0:
	  CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q2 =
	      SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d296;
      5'd1:
	  CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q2 =
	      SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d297;
      default: CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q2 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(addr_offset__h13465 or
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d304 or
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d305)
  begin
    case (addr_offset__h13465[11:7])
      5'd0:
	  CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q3 =
	      SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d304;
      5'd1:
	  CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q3 =
	      SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d305;
      default: CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q3 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(addr_offset__h13465 or
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d311 or
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d312)
  begin
    case (addr_offset__h13465[11:7])
      5'd0:
	  CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q4 =
	      SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d311;
      5'd1:
	  CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q4 =
	      SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d312;
      default: CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q4 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(addr_offset__h13465 or
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d319 or
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d320)
  begin
    case (addr_offset__h13465[11:7])
      5'd0:
	  CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q5 =
	      SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d319;
      5'd1:
	  CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q5 =
	      SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d320;
      default: CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q5 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(addr_offset__h13465 or
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d326 or
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d327)
  begin
    case (addr_offset__h13465[11:7])
      5'd0:
	  CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q6 =
	      SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d326;
      5'd1:
	  CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q6 =
	      SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d327;
      default: CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q6 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(addr_offset__h13465 or
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d334 or
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d335)
  begin
    case (addr_offset__h13465[11:7])
      5'd0:
	  CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q7 =
	      SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d334;
      5'd1:
	  CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q7 =
	      SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d335;
      default: CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q7 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(addr_offset__h13465 or
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d341 or
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d342)
  begin
    case (addr_offset__h13465[11:7])
      5'd0:
	  CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q8 =
	      SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d341;
      5'd1:
	  CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q8 =
	      SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d342;
      default: CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q8 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(addr_offset__h13465 or
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d349 or
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d350)
  begin
    case (addr_offset__h13465[11:7])
      5'd0:
	  CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q9 =
	      SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d349;
      5'd1:
	  CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q9 =
	      SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d350;
      default: CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q9 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(addr_offset__h13465 or
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d356 or
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d357)
  begin
    case (addr_offset__h13465[11:7])
      5'd0:
	  CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q10 =
	      SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d356;
      5'd1:
	  CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q10 =
	      SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d357;
      default: CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q10 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(addr_offset__h13465 or
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d364 or
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d365)
  begin
    case (addr_offset__h13465[11:7])
      5'd0:
	  CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q11 =
	      SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d364;
      5'd1:
	  CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q11 =
	      SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d365;
      default: CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q11 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(addr_offset__h13465 or
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d371 or
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d372)
  begin
    case (addr_offset__h13465[11:7])
      5'd0:
	  CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q12 =
	      SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d371;
      5'd1:
	  CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q12 =
	      SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d372;
      default: CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q12 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(addr_offset__h13465 or
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d379 or
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d380)
  begin
    case (addr_offset__h13465[11:7])
      5'd0:
	  CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q13 =
	      SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d379;
      5'd1:
	  CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q13 =
	      SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d380;
      default: CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q13 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(addr_offset__h13465 or
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d386 or
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d387)
  begin
    case (addr_offset__h13465[11:7])
      5'd0:
	  CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q14 =
	      SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d386;
      5'd1:
	  CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q14 =
	      SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d387;
      default: CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q14 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(addr_offset__h13465 or
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d394 or
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d395)
  begin
    case (addr_offset__h13465[11:7])
      5'd0:
	  CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q15 =
	      SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d394;
      5'd1:
	  CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q15 =
	      SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d395;
      default: CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q15 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(addr_offset__h13465 or
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d401 or
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d402)
  begin
    case (addr_offset__h13465[11:7])
      5'd0:
	  CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q16 =
	      SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d401;
      5'd1:
	  CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q16 =
	      SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d402;
      default: CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q16 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(addr_offset__h13465 or
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d409 or
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d410)
  begin
    case (addr_offset__h13465[11:7])
      5'd0:
	  CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q17 =
	      SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d409;
      5'd1:
	  CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q17 =
	      SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d410;
      default: CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q17 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(addr_offset__h13465 or
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d416 or
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d417)
  begin
    case (addr_offset__h13465[11:7])
      5'd0:
	  CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q18 =
	      SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d416;
      5'd1:
	  CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q18 =
	      SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d417;
      default: CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q18 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(addr_offset__h13465 or
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d424 or
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d425)
  begin
    case (addr_offset__h13465[11:7])
      5'd0:
	  CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q19 =
	      SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d424;
      5'd1:
	  CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q19 =
	      SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d425;
      default: CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q19 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(addr_offset__h13465 or
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d431 or
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d432)
  begin
    case (addr_offset__h13465[11:7])
      5'd0:
	  CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q20 =
	      SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d431;
      5'd1:
	  CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q20 =
	      SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d432;
      default: CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q20 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(addr_offset__h13465 or
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d439 or
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d440)
  begin
    case (addr_offset__h13465[11:7])
      5'd0:
	  CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q21 =
	      SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d439;
      5'd1:
	  CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q21 =
	      SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d440;
      default: CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q21 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(addr_offset__h13465 or
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d446 or
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d447)
  begin
    case (addr_offset__h13465[11:7])
      5'd0:
	  CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q22 =
	      SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d446;
      5'd1:
	  CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q22 =
	      SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d447;
      default: CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q22 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(addr_offset__h13465 or
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d454 or
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d455)
  begin
    case (addr_offset__h13465[11:7])
      5'd0:
	  CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q23 =
	      SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d454;
      5'd1:
	  CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q23 =
	      SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d455;
      default: CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q23 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(addr_offset__h13465 or
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d461 or
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d462)
  begin
    case (addr_offset__h13465[11:7])
      5'd0:
	  CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q24 =
	      SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d461;
      5'd1:
	  CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q24 =
	      SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d462;
      default: CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q24 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(addr_offset__h13465 or
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d469 or
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d470)
  begin
    case (addr_offset__h13465[11:7])
      5'd0:
	  CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q25 =
	      SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d469;
      5'd1:
	  CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q25 =
	      SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d470;
      default: CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q25 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(addr_offset__h13465 or
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d476 or
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d477)
  begin
    case (addr_offset__h13465[11:7])
      5'd0:
	  CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q26 =
	      SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d476;
      5'd1:
	  CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q26 =
	      SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d477;
      default: CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q26 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(addr_offset__h13465 or
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d484 or
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d485)
  begin
    case (addr_offset__h13465[11:7])
      5'd0:
	  CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q27 =
	      SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d484;
      5'd1:
	  CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q27 =
	      SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d485;
      default: CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q27 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(addr_offset__h13465 or
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d491 or
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d492)
  begin
    case (addr_offset__h13465[11:7])
      5'd0:
	  CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q28 =
	      SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d491;
      5'd1:
	  CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q28 =
	      SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d492;
      default: CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q28 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(addr_offset__h13465 or
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d499 or
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d500)
  begin
    case (addr_offset__h13465[11:7])
      5'd0:
	  CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q29 =
	      SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d499;
      5'd1:
	  CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q29 =
	      SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d500;
      default: CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q29 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(addr_offset__h13465 or
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d506 or
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d507)
  begin
    case (addr_offset__h13465[11:7])
      5'd0:
	  CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q30 =
	      SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d506;
      5'd1:
	  CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q30 =
	      SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d507;
      default: CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q30 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(addr_offset__h13465 or
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d514 or
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d515)
  begin
    case (addr_offset__h13465[11:7])
      5'd0:
	  CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q31 =
	      SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d514;
      5'd1:
	  CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q31 =
	      SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d515;
      default: CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q31 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(addr_offset__h13465 or
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d519 or
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d520)
  begin
    case (addr_offset__h13465[11:7])
      5'd0:
	  CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q32 =
	      SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d519;
      5'd1:
	  CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q32 =
	      SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d520;
      default: CASE_addr_offset3465_BITS_11_TO_7_0_SEL_ARR_m__ETC__q32 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(source_id__h18088 or
	  m_vrg_source_ip_0 or
	  m_vrg_source_ip_1 or
	  m_vrg_source_ip_2 or
	  m_vrg_source_ip_3 or
	  m_vrg_source_ip_4 or
	  m_vrg_source_ip_5 or
	  m_vrg_source_ip_6 or
	  m_vrg_source_ip_7 or
	  m_vrg_source_ip_8 or
	  m_vrg_source_ip_9 or
	  m_vrg_source_ip_10 or
	  m_vrg_source_ip_11 or
	  m_vrg_source_ip_12 or
	  m_vrg_source_ip_13 or
	  m_vrg_source_ip_14 or m_vrg_source_ip_15 or m_vrg_source_ip_16)
  begin
    case (source_id__h18088)
      10'd0:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d228 =
	      m_vrg_source_ip_0;
      10'd1:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d228 =
	      m_vrg_source_ip_1;
      10'd2:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d228 =
	      m_vrg_source_ip_2;
      10'd3:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d228 =
	      m_vrg_source_ip_3;
      10'd4:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d228 =
	      m_vrg_source_ip_4;
      10'd5:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d228 =
	      m_vrg_source_ip_5;
      10'd6:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d228 =
	      m_vrg_source_ip_6;
      10'd7:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d228 =
	      m_vrg_source_ip_7;
      10'd8:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d228 =
	      m_vrg_source_ip_8;
      10'd9:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d228 =
	      m_vrg_source_ip_9;
      10'd10:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d228 =
	      m_vrg_source_ip_10;
      10'd11:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d228 =
	      m_vrg_source_ip_11;
      10'd12:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d228 =
	      m_vrg_source_ip_12;
      10'd13:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d228 =
	      m_vrg_source_ip_13;
      10'd14:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d228 =
	      m_vrg_source_ip_14;
      10'd15:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d228 =
	      m_vrg_source_ip_15;
      10'd16:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d228 =
	      m_vrg_source_ip_16;
      default: SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d228 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(source_id__h18161 or
	  m_vrg_source_ip_0 or
	  m_vrg_source_ip_1 or
	  m_vrg_source_ip_2 or
	  m_vrg_source_ip_3 or
	  m_vrg_source_ip_4 or
	  m_vrg_source_ip_5 or
	  m_vrg_source_ip_6 or
	  m_vrg_source_ip_7 or
	  m_vrg_source_ip_8 or
	  m_vrg_source_ip_9 or
	  m_vrg_source_ip_10 or
	  m_vrg_source_ip_11 or
	  m_vrg_source_ip_12 or
	  m_vrg_source_ip_13 or
	  m_vrg_source_ip_14 or m_vrg_source_ip_15 or m_vrg_source_ip_16)
  begin
    case (source_id__h18161)
      10'd0:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d233 =
	      m_vrg_source_ip_0;
      10'd1:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d233 =
	      m_vrg_source_ip_1;
      10'd2:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d233 =
	      m_vrg_source_ip_2;
      10'd3:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d233 =
	      m_vrg_source_ip_3;
      10'd4:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d233 =
	      m_vrg_source_ip_4;
      10'd5:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d233 =
	      m_vrg_source_ip_5;
      10'd6:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d233 =
	      m_vrg_source_ip_6;
      10'd7:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d233 =
	      m_vrg_source_ip_7;
      10'd8:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d233 =
	      m_vrg_source_ip_8;
      10'd9:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d233 =
	      m_vrg_source_ip_9;
      10'd10:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d233 =
	      m_vrg_source_ip_10;
      10'd11:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d233 =
	      m_vrg_source_ip_11;
      10'd12:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d233 =
	      m_vrg_source_ip_12;
      10'd13:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d233 =
	      m_vrg_source_ip_13;
      10'd14:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d233 =
	      m_vrg_source_ip_14;
      10'd15:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d233 =
	      m_vrg_source_ip_15;
      10'd16:
	  SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d233 =
	      m_vrg_source_ip_16;
      default: SEL_ARR_m_vrg_source_ip_0_read__0_m_vrg_source_ETC___d233 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(x__h23928 or y_avValue_snd__h26446)
  begin
    case (x__h23928)
      32'h00200000, 32'h00200004:
	  y_avValue_snd__h26467 = y_avValue_snd__h26446;
      default: y_avValue_snd__h26467 = 2'b10;
    endcase
  end
  always@(addr_offset__h13465 or m_vvrg_ie_0_1 or m_vvrg_ie_1_1)
  begin
    case (addr_offset__h13465[16:12])
      5'd0:
	  CASE_addr_offset3465_BITS_16_TO_12_0_m_vvrg_ie_ETC__q33 =
	      m_vvrg_ie_0_1;
      5'd1:
	  CASE_addr_offset3465_BITS_16_TO_12_0_m_vvrg_ie_ETC__q33 =
	      m_vvrg_ie_1_1;
      default: CASE_addr_offset3465_BITS_16_TO_12_0_m_vvrg_ie_ETC__q33 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(addr_offset__h13465 or m_vvrg_ie_0_2 or m_vvrg_ie_1_2)
  begin
    case (addr_offset__h13465[16:12])
      5'd0:
	  CASE_addr_offset3465_BITS_16_TO_12_0_m_vvrg_ie_ETC__q34 =
	      m_vvrg_ie_0_2;
      5'd1:
	  CASE_addr_offset3465_BITS_16_TO_12_0_m_vvrg_ie_ETC__q34 =
	      m_vvrg_ie_1_2;
      default: CASE_addr_offset3465_BITS_16_TO_12_0_m_vvrg_ie_ETC__q34 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(addr_offset__h13465 or m_vvrg_ie_0_3 or m_vvrg_ie_1_3)
  begin
    case (addr_offset__h13465[16:12])
      5'd0:
	  CASE_addr_offset3465_BITS_16_TO_12_0_m_vvrg_ie_ETC__q35 =
	      m_vvrg_ie_0_3;
      5'd1:
	  CASE_addr_offset3465_BITS_16_TO_12_0_m_vvrg_ie_ETC__q35 =
	      m_vvrg_ie_1_3;
      default: CASE_addr_offset3465_BITS_16_TO_12_0_m_vvrg_ie_ETC__q35 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(addr_offset__h13465 or m_vvrg_ie_0_4 or m_vvrg_ie_1_4)
  begin
    case (addr_offset__h13465[16:12])
      5'd0:
	  CASE_addr_offset3465_BITS_16_TO_12_0_m_vvrg_ie_ETC__q36 =
	      m_vvrg_ie_0_4;
      5'd1:
	  CASE_addr_offset3465_BITS_16_TO_12_0_m_vvrg_ie_ETC__q36 =
	      m_vvrg_ie_1_4;
      default: CASE_addr_offset3465_BITS_16_TO_12_0_m_vvrg_ie_ETC__q36 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(addr_offset__h13465 or m_vvrg_ie_0_5 or m_vvrg_ie_1_5)
  begin
    case (addr_offset__h13465[16:12])
      5'd0:
	  CASE_addr_offset3465_BITS_16_TO_12_0_m_vvrg_ie_ETC__q37 =
	      m_vvrg_ie_0_5;
      5'd1:
	  CASE_addr_offset3465_BITS_16_TO_12_0_m_vvrg_ie_ETC__q37 =
	      m_vvrg_ie_1_5;
      default: CASE_addr_offset3465_BITS_16_TO_12_0_m_vvrg_ie_ETC__q37 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(addr_offset__h13465 or m_vvrg_ie_0_6 or m_vvrg_ie_1_6)
  begin
    case (addr_offset__h13465[16:12])
      5'd0:
	  CASE_addr_offset3465_BITS_16_TO_12_0_m_vvrg_ie_ETC__q38 =
	      m_vvrg_ie_0_6;
      5'd1:
	  CASE_addr_offset3465_BITS_16_TO_12_0_m_vvrg_ie_ETC__q38 =
	      m_vvrg_ie_1_6;
      default: CASE_addr_offset3465_BITS_16_TO_12_0_m_vvrg_ie_ETC__q38 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(addr_offset__h13465 or m_vvrg_ie_0_7 or m_vvrg_ie_1_7)
  begin
    case (addr_offset__h13465[16:12])
      5'd0:
	  CASE_addr_offset3465_BITS_16_TO_12_0_m_vvrg_ie_ETC__q39 =
	      m_vvrg_ie_0_7;
      5'd1:
	  CASE_addr_offset3465_BITS_16_TO_12_0_m_vvrg_ie_ETC__q39 =
	      m_vvrg_ie_1_7;
      default: CASE_addr_offset3465_BITS_16_TO_12_0_m_vvrg_ie_ETC__q39 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(addr_offset__h13465 or m_vvrg_ie_0_8 or m_vvrg_ie_1_8)
  begin
    case (addr_offset__h13465[16:12])
      5'd0:
	  CASE_addr_offset3465_BITS_16_TO_12_0_m_vvrg_ie_ETC__q40 =
	      m_vvrg_ie_0_8;
      5'd1:
	  CASE_addr_offset3465_BITS_16_TO_12_0_m_vvrg_ie_ETC__q40 =
	      m_vvrg_ie_1_8;
      default: CASE_addr_offset3465_BITS_16_TO_12_0_m_vvrg_ie_ETC__q40 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(addr_offset__h13465 or m_vvrg_ie_0_9 or m_vvrg_ie_1_9)
  begin
    case (addr_offset__h13465[16:12])
      5'd0:
	  CASE_addr_offset3465_BITS_16_TO_12_0_m_vvrg_ie_ETC__q41 =
	      m_vvrg_ie_0_9;
      5'd1:
	  CASE_addr_offset3465_BITS_16_TO_12_0_m_vvrg_ie_ETC__q41 =
	      m_vvrg_ie_1_9;
      default: CASE_addr_offset3465_BITS_16_TO_12_0_m_vvrg_ie_ETC__q41 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(addr_offset__h13465 or m_vvrg_ie_0_10 or m_vvrg_ie_1_10)
  begin
    case (addr_offset__h13465[16:12])
      5'd0:
	  CASE_addr_offset3465_BITS_16_TO_12_0_m_vvrg_ie_ETC__q42 =
	      m_vvrg_ie_0_10;
      5'd1:
	  CASE_addr_offset3465_BITS_16_TO_12_0_m_vvrg_ie_ETC__q42 =
	      m_vvrg_ie_1_10;
      default: CASE_addr_offset3465_BITS_16_TO_12_0_m_vvrg_ie_ETC__q42 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(addr_offset__h13465 or m_vvrg_ie_0_11 or m_vvrg_ie_1_11)
  begin
    case (addr_offset__h13465[16:12])
      5'd0:
	  CASE_addr_offset3465_BITS_16_TO_12_0_m_vvrg_ie_ETC__q43 =
	      m_vvrg_ie_0_11;
      5'd1:
	  CASE_addr_offset3465_BITS_16_TO_12_0_m_vvrg_ie_ETC__q43 =
	      m_vvrg_ie_1_11;
      default: CASE_addr_offset3465_BITS_16_TO_12_0_m_vvrg_ie_ETC__q43 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(addr_offset__h13465 or m_vvrg_ie_0_12 or m_vvrg_ie_1_12)
  begin
    case (addr_offset__h13465[16:12])
      5'd0:
	  CASE_addr_offset3465_BITS_16_TO_12_0_m_vvrg_ie_ETC__q44 =
	      m_vvrg_ie_0_12;
      5'd1:
	  CASE_addr_offset3465_BITS_16_TO_12_0_m_vvrg_ie_ETC__q44 =
	      m_vvrg_ie_1_12;
      default: CASE_addr_offset3465_BITS_16_TO_12_0_m_vvrg_ie_ETC__q44 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(addr_offset__h13465 or m_vvrg_ie_0_13 or m_vvrg_ie_1_13)
  begin
    case (addr_offset__h13465[16:12])
      5'd0:
	  CASE_addr_offset3465_BITS_16_TO_12_0_m_vvrg_ie_ETC__q45 =
	      m_vvrg_ie_0_13;
      5'd1:
	  CASE_addr_offset3465_BITS_16_TO_12_0_m_vvrg_ie_ETC__q45 =
	      m_vvrg_ie_1_13;
      default: CASE_addr_offset3465_BITS_16_TO_12_0_m_vvrg_ie_ETC__q45 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(addr_offset__h13465 or m_vvrg_ie_0_14 or m_vvrg_ie_1_14)
  begin
    case (addr_offset__h13465[16:12])
      5'd0:
	  CASE_addr_offset3465_BITS_16_TO_12_0_m_vvrg_ie_ETC__q46 =
	      m_vvrg_ie_0_14;
      5'd1:
	  CASE_addr_offset3465_BITS_16_TO_12_0_m_vvrg_ie_ETC__q46 =
	      m_vvrg_ie_1_14;
      default: CASE_addr_offset3465_BITS_16_TO_12_0_m_vvrg_ie_ETC__q46 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(addr_offset__h13465 or m_vvrg_ie_0_15 or m_vvrg_ie_1_15)
  begin
    case (addr_offset__h13465[16:12])
      5'd0:
	  CASE_addr_offset3465_BITS_16_TO_12_0_m_vvrg_ie_ETC__q47 =
	      m_vvrg_ie_0_15;
      5'd1:
	  CASE_addr_offset3465_BITS_16_TO_12_0_m_vvrg_ie_ETC__q47 =
	      m_vvrg_ie_1_15;
      default: CASE_addr_offset3465_BITS_16_TO_12_0_m_vvrg_ie_ETC__q47 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(addr_offset__h13465 or m_vvrg_ie_0_16 or m_vvrg_ie_1_16)
  begin
    case (addr_offset__h13465[16:12])
      5'd0:
	  CASE_addr_offset3465_BITS_16_TO_12_0_m_vvrg_ie_ETC__q48 =
	      m_vvrg_ie_0_16;
      5'd1:
	  CASE_addr_offset3465_BITS_16_TO_12_0_m_vvrg_ie_ETC__q48 =
	      m_vvrg_ie_1_16;
      default: CASE_addr_offset3465_BITS_16_TO_12_0_m_vvrg_ie_ETC__q48 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(x__h23928 or y_avValue_fst__h26445 or y_avValue_fst__h26433)
  begin
    case (x__h23928)
      32'h00200000: y_avValue_fst__h26466 = y_avValue_fst__h26445;
      32'h00200004: y_avValue_fst__h26466 = y_avValue_fst__h26433;
      default: y_avValue_fst__h26466 = 64'd0;
    endcase
  end
  always@(x__h76716 or v__h76750)
  begin
    case (x__h76716)
      32'h00200000, 32'h00200004: v__h76713 = v__h76750;
      default: v__h76713 = 2'b10;
    endcase
  end
  always@(wdata32__h27246 or
	  m_vvrg_ie_0_0 or
	  m_vvrg_ie_0_1 or
	  m_vvrg_ie_0_2 or
	  m_vvrg_ie_0_3 or
	  m_vvrg_ie_0_4 or
	  m_vvrg_ie_0_5 or
	  m_vvrg_ie_0_6 or
	  m_vvrg_ie_0_7 or
	  m_vvrg_ie_0_8 or
	  m_vvrg_ie_0_9 or
	  m_vvrg_ie_0_10 or
	  m_vvrg_ie_0_11 or
	  m_vvrg_ie_0_12 or
	  m_vvrg_ie_0_13 or
	  m_vvrg_ie_0_14 or m_vvrg_ie_0_15 or m_vvrg_ie_0_16)
  begin
    case (wdata32__h27246[9:0])
      10'd0:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d2875 =
	      m_vvrg_ie_0_0;
      10'd1:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d2875 =
	      m_vvrg_ie_0_1;
      10'd2:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d2875 =
	      m_vvrg_ie_0_2;
      10'd3:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d2875 =
	      m_vvrg_ie_0_3;
      10'd4:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d2875 =
	      m_vvrg_ie_0_4;
      10'd5:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d2875 =
	      m_vvrg_ie_0_5;
      10'd6:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d2875 =
	      m_vvrg_ie_0_6;
      10'd7:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d2875 =
	      m_vvrg_ie_0_7;
      10'd8:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d2875 =
	      m_vvrg_ie_0_8;
      10'd9:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d2875 =
	      m_vvrg_ie_0_9;
      10'd10:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d2875 =
	      m_vvrg_ie_0_10;
      10'd11:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d2875 =
	      m_vvrg_ie_0_11;
      10'd12:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d2875 =
	      m_vvrg_ie_0_12;
      10'd13:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d2875 =
	      m_vvrg_ie_0_13;
      10'd14:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d2875 =
	      m_vvrg_ie_0_14;
      10'd15:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d2875 =
	      m_vvrg_ie_0_15;
      10'd16:
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d2875 =
	      m_vvrg_ie_0_16;
      default: SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d2875 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(wdata32__h27246 or
	  m_vvrg_ie_1_0 or
	  m_vvrg_ie_1_1 or
	  m_vvrg_ie_1_2 or
	  m_vvrg_ie_1_3 or
	  m_vvrg_ie_1_4 or
	  m_vvrg_ie_1_5 or
	  m_vvrg_ie_1_6 or
	  m_vvrg_ie_1_7 or
	  m_vvrg_ie_1_8 or
	  m_vvrg_ie_1_9 or
	  m_vvrg_ie_1_10 or
	  m_vvrg_ie_1_11 or
	  m_vvrg_ie_1_12 or
	  m_vvrg_ie_1_13 or
	  m_vvrg_ie_1_14 or m_vvrg_ie_1_15 or m_vvrg_ie_1_16)
  begin
    case (wdata32__h27246[9:0])
      10'd0:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d2876 =
	      m_vvrg_ie_1_0;
      10'd1:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d2876 =
	      m_vvrg_ie_1_1;
      10'd2:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d2876 =
	      m_vvrg_ie_1_2;
      10'd3:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d2876 =
	      m_vvrg_ie_1_3;
      10'd4:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d2876 =
	      m_vvrg_ie_1_4;
      10'd5:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d2876 =
	      m_vvrg_ie_1_5;
      10'd6:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d2876 =
	      m_vvrg_ie_1_6;
      10'd7:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d2876 =
	      m_vvrg_ie_1_7;
      10'd8:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d2876 =
	      m_vvrg_ie_1_8;
      10'd9:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d2876 =
	      m_vvrg_ie_1_9;
      10'd10:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d2876 =
	      m_vvrg_ie_1_10;
      10'd11:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d2876 =
	      m_vvrg_ie_1_11;
      10'd12:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d2876 =
	      m_vvrg_ie_1_12;
      10'd13:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d2876 =
	      m_vvrg_ie_1_13;
      10'd14:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d2876 =
	      m_vvrg_ie_1_14;
      10'd15:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d2876 =
	      m_vvrg_ie_1_15;
      10'd16:
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d2876 =
	      m_vvrg_ie_1_16;
      default: SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d2876 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  always@(addr_offset__h27245 or
	  SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d2875 or
	  SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d2876)
  begin
    case (addr_offset__h27245[16:12])
      5'd0:
	  SEL_ARR_SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_ETC___d2878 =
	      SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_54_m_vv_ETC___d2875;
      5'd1:
	  SEL_ARR_SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_ETC___d2878 =
	      SEL_ARR_m_vvrg_ie_1_0_72_m_vvrg_ie_1_1_73_m_vv_ETC___d2876;
      default: SEL_ARR_SEL_ARR_m_vvrg_ie_0_0_53_m_vvrg_ie_0_1_ETC___d2878 =
		   1'b0 /* unspecified value */ ;
    endcase
  end
  // handling of inlined registers
  always@(posedge CLK)
  begin
    if (RST_N == `BSV_RESET_VALUE)
      begin
        m_cfg_verbosity <= `BSV_ASSIGNMENT_DELAY 4'd0;
	m_vrg_source_busy_0 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	m_vrg_source_busy_1 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	m_vrg_source_busy_10 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	m_vrg_source_busy_11 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	m_vrg_source_busy_12 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	m_vrg_source_busy_13 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	m_vrg_source_busy_14 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	m_vrg_source_busy_15 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	m_vrg_source_busy_16 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	m_vrg_source_busy_2 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	m_vrg_source_busy_3 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	m_vrg_source_busy_4 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	m_vrg_source_busy_5 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	m_vrg_source_busy_6 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	m_vrg_source_busy_7 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	m_vrg_source_busy_8 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	m_vrg_source_busy_9 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	m_vrg_source_ip_0 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	m_vrg_source_ip_1 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	m_vrg_source_ip_10 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	m_vrg_source_ip_11 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	m_vrg_source_ip_12 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	m_vrg_source_ip_13 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	m_vrg_source_ip_14 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	m_vrg_source_ip_15 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	m_vrg_source_ip_16 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	m_vrg_source_ip_2 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	m_vrg_source_ip_3 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	m_vrg_source_ip_4 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	m_vrg_source_ip_5 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	m_vrg_source_ip_6 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	m_vrg_source_ip_7 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	m_vrg_source_ip_8 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	m_vrg_source_ip_9 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	m_vrg_source_prio_0 <= `BSV_ASSIGNMENT_DELAY 3'd0;
	m_vrg_source_prio_1 <= `BSV_ASSIGNMENT_DELAY 3'd0;
	m_vrg_source_prio_10 <= `BSV_ASSIGNMENT_DELAY 3'd0;
	m_vrg_source_prio_11 <= `BSV_ASSIGNMENT_DELAY 3'd0;
	m_vrg_source_prio_12 <= `BSV_ASSIGNMENT_DELAY 3'd0;
	m_vrg_source_prio_13 <= `BSV_ASSIGNMENT_DELAY 3'd0;
	m_vrg_source_prio_14 <= `BSV_ASSIGNMENT_DELAY 3'd0;
	m_vrg_source_prio_15 <= `BSV_ASSIGNMENT_DELAY 3'd0;
	m_vrg_source_prio_16 <= `BSV_ASSIGNMENT_DELAY 3'd0;
	m_vrg_source_prio_2 <= `BSV_ASSIGNMENT_DELAY 3'd0;
	m_vrg_source_prio_3 <= `BSV_ASSIGNMENT_DELAY 3'd0;
	m_vrg_source_prio_4 <= `BSV_ASSIGNMENT_DELAY 3'd0;
	m_vrg_source_prio_5 <= `BSV_ASSIGNMENT_DELAY 3'd0;
	m_vrg_source_prio_6 <= `BSV_ASSIGNMENT_DELAY 3'd0;
	m_vrg_source_prio_7 <= `BSV_ASSIGNMENT_DELAY 3'd0;
	m_vrg_source_prio_8 <= `BSV_ASSIGNMENT_DELAY 3'd0;
	m_vrg_source_prio_9 <= `BSV_ASSIGNMENT_DELAY 3'd0;
	m_vrg_target_threshold_0 <= `BSV_ASSIGNMENT_DELAY 3'd7;
	m_vrg_target_threshold_1 <= `BSV_ASSIGNMENT_DELAY 3'd7;
	m_vvrg_ie_0_0 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	m_vvrg_ie_0_1 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	m_vvrg_ie_0_10 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	m_vvrg_ie_0_11 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	m_vvrg_ie_0_12 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	m_vvrg_ie_0_13 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	m_vvrg_ie_0_14 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	m_vvrg_ie_0_15 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	m_vvrg_ie_0_16 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	m_vvrg_ie_0_2 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	m_vvrg_ie_0_3 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	m_vvrg_ie_0_4 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	m_vvrg_ie_0_5 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	m_vvrg_ie_0_6 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	m_vvrg_ie_0_7 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	m_vvrg_ie_0_8 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	m_vvrg_ie_0_9 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	m_vvrg_ie_1_0 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	m_vvrg_ie_1_1 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	m_vvrg_ie_1_10 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	m_vvrg_ie_1_11 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	m_vvrg_ie_1_12 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	m_vvrg_ie_1_13 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	m_vvrg_ie_1_14 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	m_vvrg_ie_1_15 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	m_vvrg_ie_1_16 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	m_vvrg_ie_1_2 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	m_vvrg_ie_1_3 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	m_vvrg_ie_1_4 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	m_vvrg_ie_1_5 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	m_vvrg_ie_1_6 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	m_vvrg_ie_1_7 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	m_vvrg_ie_1_8 <= `BSV_ASSIGNMENT_DELAY 1'd0;
	m_vvrg_ie_1_9 <= `BSV_ASSIGNMENT_DELAY 1'd0;
      end
    else
      begin
        if (m_cfg_verbosity$EN)
	  m_cfg_verbosity <= `BSV_ASSIGNMENT_DELAY m_cfg_verbosity$D_IN;
	if (m_vrg_source_busy_0$EN)
	  m_vrg_source_busy_0 <= `BSV_ASSIGNMENT_DELAY
	      m_vrg_source_busy_0$D_IN;
	if (m_vrg_source_busy_1$EN)
	  m_vrg_source_busy_1 <= `BSV_ASSIGNMENT_DELAY
	      m_vrg_source_busy_1$D_IN;
	if (m_vrg_source_busy_10$EN)
	  m_vrg_source_busy_10 <= `BSV_ASSIGNMENT_DELAY
	      m_vrg_source_busy_10$D_IN;
	if (m_vrg_source_busy_11$EN)
	  m_vrg_source_busy_11 <= `BSV_ASSIGNMENT_DELAY
	      m_vrg_source_busy_11$D_IN;
	if (m_vrg_source_busy_12$EN)
	  m_vrg_source_busy_12 <= `BSV_ASSIGNMENT_DELAY
	      m_vrg_source_busy_12$D_IN;
	if (m_vrg_source_busy_13$EN)
	  m_vrg_source_busy_13 <= `BSV_ASSIGNMENT_DELAY
	      m_vrg_source_busy_13$D_IN;
	if (m_vrg_source_busy_14$EN)
	  m_vrg_source_busy_14 <= `BSV_ASSIGNMENT_DELAY
	      m_vrg_source_busy_14$D_IN;
	if (m_vrg_source_busy_15$EN)
	  m_vrg_source_busy_15 <= `BSV_ASSIGNMENT_DELAY
	      m_vrg_source_busy_15$D_IN;
	if (m_vrg_source_busy_16$EN)
	  m_vrg_source_busy_16 <= `BSV_ASSIGNMENT_DELAY
	      m_vrg_source_busy_16$D_IN;
	if (m_vrg_source_busy_2$EN)
	  m_vrg_source_busy_2 <= `BSV_ASSIGNMENT_DELAY
	      m_vrg_source_busy_2$D_IN;
	if (m_vrg_source_busy_3$EN)
	  m_vrg_source_busy_3 <= `BSV_ASSIGNMENT_DELAY
	      m_vrg_source_busy_3$D_IN;
	if (m_vrg_source_busy_4$EN)
	  m_vrg_source_busy_4 <= `BSV_ASSIGNMENT_DELAY
	      m_vrg_source_busy_4$D_IN;
	if (m_vrg_source_busy_5$EN)
	  m_vrg_source_busy_5 <= `BSV_ASSIGNMENT_DELAY
	      m_vrg_source_busy_5$D_IN;
	if (m_vrg_source_busy_6$EN)
	  m_vrg_source_busy_6 <= `BSV_ASSIGNMENT_DELAY
	      m_vrg_source_busy_6$D_IN;
	if (m_vrg_source_busy_7$EN)
	  m_vrg_source_busy_7 <= `BSV_ASSIGNMENT_DELAY
	      m_vrg_source_busy_7$D_IN;
	if (m_vrg_source_busy_8$EN)
	  m_vrg_source_busy_8 <= `BSV_ASSIGNMENT_DELAY
	      m_vrg_source_busy_8$D_IN;
	if (m_vrg_source_busy_9$EN)
	  m_vrg_source_busy_9 <= `BSV_ASSIGNMENT_DELAY
	      m_vrg_source_busy_9$D_IN;
	if (m_vrg_source_ip_0$EN)
	  m_vrg_source_ip_0 <= `BSV_ASSIGNMENT_DELAY m_vrg_source_ip_0$D_IN;
	if (m_vrg_source_ip_1$EN)
	  m_vrg_source_ip_1 <= `BSV_ASSIGNMENT_DELAY m_vrg_source_ip_1$D_IN;
	if (m_vrg_source_ip_10$EN)
	  m_vrg_source_ip_10 <= `BSV_ASSIGNMENT_DELAY m_vrg_source_ip_10$D_IN;
	if (m_vrg_source_ip_11$EN)
	  m_vrg_source_ip_11 <= `BSV_ASSIGNMENT_DELAY m_vrg_source_ip_11$D_IN;
	if (m_vrg_source_ip_12$EN)
	  m_vrg_source_ip_12 <= `BSV_ASSIGNMENT_DELAY m_vrg_source_ip_12$D_IN;
	if (m_vrg_source_ip_13$EN)
	  m_vrg_source_ip_13 <= `BSV_ASSIGNMENT_DELAY m_vrg_source_ip_13$D_IN;
	if (m_vrg_source_ip_14$EN)
	  m_vrg_source_ip_14 <= `BSV_ASSIGNMENT_DELAY m_vrg_source_ip_14$D_IN;
	if (m_vrg_source_ip_15$EN)
	  m_vrg_source_ip_15 <= `BSV_ASSIGNMENT_DELAY m_vrg_source_ip_15$D_IN;
	if (m_vrg_source_ip_16$EN)
	  m_vrg_source_ip_16 <= `BSV_ASSIGNMENT_DELAY m_vrg_source_ip_16$D_IN;
	if (m_vrg_source_ip_2$EN)
	  m_vrg_source_ip_2 <= `BSV_ASSIGNMENT_DELAY m_vrg_source_ip_2$D_IN;
	if (m_vrg_source_ip_3$EN)
	  m_vrg_source_ip_3 <= `BSV_ASSIGNMENT_DELAY m_vrg_source_ip_3$D_IN;
	if (m_vrg_source_ip_4$EN)
	  m_vrg_source_ip_4 <= `BSV_ASSIGNMENT_DELAY m_vrg_source_ip_4$D_IN;
	if (m_vrg_source_ip_5$EN)
	  m_vrg_source_ip_5 <= `BSV_ASSIGNMENT_DELAY m_vrg_source_ip_5$D_IN;
	if (m_vrg_source_ip_6$EN)
	  m_vrg_source_ip_6 <= `BSV_ASSIGNMENT_DELAY m_vrg_source_ip_6$D_IN;
	if (m_vrg_source_ip_7$EN)
	  m_vrg_source_ip_7 <= `BSV_ASSIGNMENT_DELAY m_vrg_source_ip_7$D_IN;
	if (m_vrg_source_ip_8$EN)
	  m_vrg_source_ip_8 <= `BSV_ASSIGNMENT_DELAY m_vrg_source_ip_8$D_IN;
	if (m_vrg_source_ip_9$EN)
	  m_vrg_source_ip_9 <= `BSV_ASSIGNMENT_DELAY m_vrg_source_ip_9$D_IN;
	if (m_vrg_source_prio_0$EN)
	  m_vrg_source_prio_0 <= `BSV_ASSIGNMENT_DELAY
	      m_vrg_source_prio_0$D_IN;
	if (m_vrg_source_prio_1$EN)
	  m_vrg_source_prio_1 <= `BSV_ASSIGNMENT_DELAY
	      m_vrg_source_prio_1$D_IN;
	if (m_vrg_source_prio_10$EN)
	  m_vrg_source_prio_10 <= `BSV_ASSIGNMENT_DELAY
	      m_vrg_source_prio_10$D_IN;
	if (m_vrg_source_prio_11$EN)
	  m_vrg_source_prio_11 <= `BSV_ASSIGNMENT_DELAY
	      m_vrg_source_prio_11$D_IN;
	if (m_vrg_source_prio_12$EN)
	  m_vrg_source_prio_12 <= `BSV_ASSIGNMENT_DELAY
	      m_vrg_source_prio_12$D_IN;
	if (m_vrg_source_prio_13$EN)
	  m_vrg_source_prio_13 <= `BSV_ASSIGNMENT_DELAY
	      m_vrg_source_prio_13$D_IN;
	if (m_vrg_source_prio_14$EN)
	  m_vrg_source_prio_14 <= `BSV_ASSIGNMENT_DELAY
	      m_vrg_source_prio_14$D_IN;
	if (m_vrg_source_prio_15$EN)
	  m_vrg_source_prio_15 <= `BSV_ASSIGNMENT_DELAY
	      m_vrg_source_prio_15$D_IN;
	if (m_vrg_source_prio_16$EN)
	  m_vrg_source_prio_16 <= `BSV_ASSIGNMENT_DELAY
	      m_vrg_source_prio_16$D_IN;
	if (m_vrg_source_prio_2$EN)
	  m_vrg_source_prio_2 <= `BSV_ASSIGNMENT_DELAY
	      m_vrg_source_prio_2$D_IN;
	if (m_vrg_source_prio_3$EN)
	  m_vrg_source_prio_3 <= `BSV_ASSIGNMENT_DELAY
	      m_vrg_source_prio_3$D_IN;
	if (m_vrg_source_prio_4$EN)
	  m_vrg_source_prio_4 <= `BSV_ASSIGNMENT_DELAY
	      m_vrg_source_prio_4$D_IN;
	if (m_vrg_source_prio_5$EN)
	  m_vrg_source_prio_5 <= `BSV_ASSIGNMENT_DELAY
	      m_vrg_source_prio_5$D_IN;
	if (m_vrg_source_prio_6$EN)
	  m_vrg_source_prio_6 <= `BSV_ASSIGNMENT_DELAY
	      m_vrg_source_prio_6$D_IN;
	if (m_vrg_source_prio_7$EN)
	  m_vrg_source_prio_7 <= `BSV_ASSIGNMENT_DELAY
	      m_vrg_source_prio_7$D_IN;
	if (m_vrg_source_prio_8$EN)
	  m_vrg_source_prio_8 <= `BSV_ASSIGNMENT_DELAY
	      m_vrg_source_prio_8$D_IN;
	if (m_vrg_source_prio_9$EN)
	  m_vrg_source_prio_9 <= `BSV_ASSIGNMENT_DELAY
	      m_vrg_source_prio_9$D_IN;
	if (m_vrg_target_threshold_0$EN)
	  m_vrg_target_threshold_0 <= `BSV_ASSIGNMENT_DELAY
	      m_vrg_target_threshold_0$D_IN;
	if (m_vrg_target_threshold_1$EN)
	  m_vrg_target_threshold_1 <= `BSV_ASSIGNMENT_DELAY
	      m_vrg_target_threshold_1$D_IN;
	if (m_vvrg_ie_0_0$EN)
	  m_vvrg_ie_0_0 <= `BSV_ASSIGNMENT_DELAY m_vvrg_ie_0_0$D_IN;
	if (m_vvrg_ie_0_1$EN)
	  m_vvrg_ie_0_1 <= `BSV_ASSIGNMENT_DELAY m_vvrg_ie_0_1$D_IN;
	if (m_vvrg_ie_0_10$EN)
	  m_vvrg_ie_0_10 <= `BSV_ASSIGNMENT_DELAY m_vvrg_ie_0_10$D_IN;
	if (m_vvrg_ie_0_11$EN)
	  m_vvrg_ie_0_11 <= `BSV_ASSIGNMENT_DELAY m_vvrg_ie_0_11$D_IN;
	if (m_vvrg_ie_0_12$EN)
	  m_vvrg_ie_0_12 <= `BSV_ASSIGNMENT_DELAY m_vvrg_ie_0_12$D_IN;
	if (m_vvrg_ie_0_13$EN)
	  m_vvrg_ie_0_13 <= `BSV_ASSIGNMENT_DELAY m_vvrg_ie_0_13$D_IN;
	if (m_vvrg_ie_0_14$EN)
	  m_vvrg_ie_0_14 <= `BSV_ASSIGNMENT_DELAY m_vvrg_ie_0_14$D_IN;
	if (m_vvrg_ie_0_15$EN)
	  m_vvrg_ie_0_15 <= `BSV_ASSIGNMENT_DELAY m_vvrg_ie_0_15$D_IN;
	if (m_vvrg_ie_0_16$EN)
	  m_vvrg_ie_0_16 <= `BSV_ASSIGNMENT_DELAY m_vvrg_ie_0_16$D_IN;
	if (m_vvrg_ie_0_2$EN)
	  m_vvrg_ie_0_2 <= `BSV_ASSIGNMENT_DELAY m_vvrg_ie_0_2$D_IN;
	if (m_vvrg_ie_0_3$EN)
	  m_vvrg_ie_0_3 <= `BSV_ASSIGNMENT_DELAY m_vvrg_ie_0_3$D_IN;
	if (m_vvrg_ie_0_4$EN)
	  m_vvrg_ie_0_4 <= `BSV_ASSIGNMENT_DELAY m_vvrg_ie_0_4$D_IN;
	if (m_vvrg_ie_0_5$EN)
	  m_vvrg_ie_0_5 <= `BSV_ASSIGNMENT_DELAY m_vvrg_ie_0_5$D_IN;
	if (m_vvrg_ie_0_6$EN)
	  m_vvrg_ie_0_6 <= `BSV_ASSIGNMENT_DELAY m_vvrg_ie_0_6$D_IN;
	if (m_vvrg_ie_0_7$EN)
	  m_vvrg_ie_0_7 <= `BSV_ASSIGNMENT_DELAY m_vvrg_ie_0_7$D_IN;
	if (m_vvrg_ie_0_8$EN)
	  m_vvrg_ie_0_8 <= `BSV_ASSIGNMENT_DELAY m_vvrg_ie_0_8$D_IN;
	if (m_vvrg_ie_0_9$EN)
	  m_vvrg_ie_0_9 <= `BSV_ASSIGNMENT_DELAY m_vvrg_ie_0_9$D_IN;
	if (m_vvrg_ie_1_0$EN)
	  m_vvrg_ie_1_0 <= `BSV_ASSIGNMENT_DELAY m_vvrg_ie_1_0$D_IN;
	if (m_vvrg_ie_1_1$EN)
	  m_vvrg_ie_1_1 <= `BSV_ASSIGNMENT_DELAY m_vvrg_ie_1_1$D_IN;
	if (m_vvrg_ie_1_10$EN)
	  m_vvrg_ie_1_10 <= `BSV_ASSIGNMENT_DELAY m_vvrg_ie_1_10$D_IN;
	if (m_vvrg_ie_1_11$EN)
	  m_vvrg_ie_1_11 <= `BSV_ASSIGNMENT_DELAY m_vvrg_ie_1_11$D_IN;
	if (m_vvrg_ie_1_12$EN)
	  m_vvrg_ie_1_12 <= `BSV_ASSIGNMENT_DELAY m_vvrg_ie_1_12$D_IN;
	if (m_vvrg_ie_1_13$EN)
	  m_vvrg_ie_1_13 <= `BSV_ASSIGNMENT_DELAY m_vvrg_ie_1_13$D_IN;
	if (m_vvrg_ie_1_14$EN)
	  m_vvrg_ie_1_14 <= `BSV_ASSIGNMENT_DELAY m_vvrg_ie_1_14$D_IN;
	if (m_vvrg_ie_1_15$EN)
	  m_vvrg_ie_1_15 <= `BSV_ASSIGNMENT_DELAY m_vvrg_ie_1_15$D_IN;
	if (m_vvrg_ie_1_16$EN)
	  m_vvrg_ie_1_16 <= `BSV_ASSIGNMENT_DELAY m_vvrg_ie_1_16$D_IN;
	if (m_vvrg_ie_1_2$EN)
	  m_vvrg_ie_1_2 <= `BSV_ASSIGNMENT_DELAY m_vvrg_ie_1_2$D_IN;
	if (m_vvrg_ie_1_3$EN)
	  m_vvrg_ie_1_3 <= `BSV_ASSIGNMENT_DELAY m_vvrg_ie_1_3$D_IN;
	if (m_vvrg_ie_1_4$EN)
	  m_vvrg_ie_1_4 <= `BSV_ASSIGNMENT_DELAY m_vvrg_ie_1_4$D_IN;
	if (m_vvrg_ie_1_5$EN)
	  m_vvrg_ie_1_5 <= `BSV_ASSIGNMENT_DELAY m_vvrg_ie_1_5$D_IN;
	if (m_vvrg_ie_1_6$EN)
	  m_vvrg_ie_1_6 <= `BSV_ASSIGNMENT_DELAY m_vvrg_ie_1_6$D_IN;
	if (m_vvrg_ie_1_7$EN)
	  m_vvrg_ie_1_7 <= `BSV_ASSIGNMENT_DELAY m_vvrg_ie_1_7$D_IN;
	if (m_vvrg_ie_1_8$EN)
	  m_vvrg_ie_1_8 <= `BSV_ASSIGNMENT_DELAY m_vvrg_ie_1_8$D_IN;
	if (m_vvrg_ie_1_9$EN)
	  m_vvrg_ie_1_9 <= `BSV_ASSIGNMENT_DELAY m_vvrg_ie_1_9$D_IN;
      end
    if (m_rg_addr_base$EN)
      m_rg_addr_base <= `BSV_ASSIGNMENT_DELAY m_rg_addr_base$D_IN;
    if (m_rg_addr_lim$EN)
      m_rg_addr_lim <= `BSV_ASSIGNMENT_DELAY m_rg_addr_lim$D_IN;
  end
  // synopsys translate_off
  `ifdef BSV_NO_INITIAL_BLOCKS
  `else // not BSV_NO_INITIAL_BLOCKS
  initial
  begin
    m_cfg_verbosity = 4'hA;
    m_rg_addr_base = 64'hAAAAAAAAAAAAAAAA;
    m_rg_addr_lim = 64'hAAAAAAAAAAAAAAAA;
    m_vrg_source_busy_0 = 1'h0;
    m_vrg_source_busy_1 = 1'h0;
    m_vrg_source_busy_10 = 1'h0;
    m_vrg_source_busy_11 = 1'h0;
    m_vrg_source_busy_12 = 1'h0;
    m_vrg_source_busy_13 = 1'h0;
    m_vrg_source_busy_14 = 1'h0;
    m_vrg_source_busy_15 = 1'h0;
    m_vrg_source_busy_16 = 1'h0;
    m_vrg_source_busy_2 = 1'h0;
    m_vrg_source_busy_3 = 1'h0;
    m_vrg_source_busy_4 = 1'h0;
    m_vrg_source_busy_5 = 1'h0;
    m_vrg_source_busy_6 = 1'h0;
    m_vrg_source_busy_7 = 1'h0;
    m_vrg_source_busy_8 = 1'h0;
    m_vrg_source_busy_9 = 1'h0;
    m_vrg_source_ip_0 = 1'h0;
    m_vrg_source_ip_1 = 1'h0;
    m_vrg_source_ip_10 = 1'h0;
    m_vrg_source_ip_11 = 1'h0;
    m_vrg_source_ip_12 = 1'h0;
    m_vrg_source_ip_13 = 1'h0;
    m_vrg_source_ip_14 = 1'h0;
    m_vrg_source_ip_15 = 1'h0;
    m_vrg_source_ip_16 = 1'h0;
    m_vrg_source_ip_2 = 1'h0;
    m_vrg_source_ip_3 = 1'h0;
    m_vrg_source_ip_4 = 1'h0;
    m_vrg_source_ip_5 = 1'h0;
    m_vrg_source_ip_6 = 1'h0;
    m_vrg_source_ip_7 = 1'h0;
    m_vrg_source_ip_8 = 1'h0;
    m_vrg_source_ip_9 = 1'h0;
    m_vrg_source_prio_0 = 3'h2;
    m_vrg_source_prio_1 = 3'h2;
    m_vrg_source_prio_10 = 3'h2;
    m_vrg_source_prio_11 = 3'h2;
    m_vrg_source_prio_12 = 3'h2;
    m_vrg_source_prio_13 = 3'h2;
    m_vrg_source_prio_14 = 3'h2;
    m_vrg_source_prio_15 = 3'h2;
    m_vrg_source_prio_16 = 3'h2;
    m_vrg_source_prio_2 = 3'h2;
    m_vrg_source_prio_3 = 3'h2;
    m_vrg_source_prio_4 = 3'h2;
    m_vrg_source_prio_5 = 3'h2;
    m_vrg_source_prio_6 = 3'h2;
    m_vrg_source_prio_7 = 3'h2;
    m_vrg_source_prio_8 = 3'h2;
    m_vrg_source_prio_9 = 3'h2;
    m_vrg_target_threshold_0 = 3'h2;
    m_vrg_target_threshold_1 = 3'h2;
    m_vvrg_ie_0_0 = 1'h0;
    m_vvrg_ie_0_1 = 1'h0;
    m_vvrg_ie_0_10 = 1'h0;
    m_vvrg_ie_0_11 = 1'h0;
    m_vvrg_ie_0_12 = 1'h0;
    m_vvrg_ie_0_13 = 1'h0;
    m_vvrg_ie_0_14 = 1'h0;
    m_vvrg_ie_0_15 = 1'h0;
    m_vvrg_ie_0_16 = 1'h0;
    m_vvrg_ie_0_2 = 1'h0;
    m_vvrg_ie_0_3 = 1'h0;
    m_vvrg_ie_0_4 = 1'h0;
    m_vvrg_ie_0_5 = 1'h0;
    m_vvrg_ie_0_6 = 1'h0;
    m_vvrg_ie_0_7 = 1'h0;
    m_vvrg_ie_0_8 = 1'h0;
    m_vvrg_ie_0_9 = 1'h0;
    m_vvrg_ie_1_0 = 1'h0;
    m_vvrg_ie_1_1 = 1'h0;
    m_vvrg_ie_1_10 = 1'h0;
    m_vvrg_ie_1_11 = 1'h0;
    m_vvrg_ie_1_12 = 1'h0;
    m_vvrg_ie_1_13 = 1'h0;
    m_vvrg_ie_1_14 = 1'h0;
    m_vvrg_ie_1_15 = 1'h0;
    m_vvrg_ie_1_16 = 1'h0;
    m_vvrg_ie_1_2 = 1'h0;
    m_vvrg_ie_1_3 = 1'h0;
    m_vvrg_ie_1_4 = 1'h0;
    m_vvrg_ie_1_5 = 1'h0;
    m_vvrg_ie_1_6 = 1'h0;
    m_vvrg_ie_1_7 = 1'h0;
    m_vvrg_ie_1_8 = 1'h0;
    m_vvrg_ie_1_9 = 1'h0;
  end
  `endif // BSV_NO_INITIAL_BLOCKS
  // synopsys translate_on
  // handling of system tasks
  // synopsys translate_off
  always@(negedge CLK)
  begin
    #0;
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_show_PLIC_state) $display("----------------");
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_show_PLIC_state) $write("Src IPs  :");
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_show_PLIC_state) $write(" %0d", m_vrg_source_ip_0);
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_show_PLIC_state) $write(" %0d", m_vrg_source_ip_1);
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_show_PLIC_state) $write(" %0d", m_vrg_source_ip_2);
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_show_PLIC_state) $write(" %0d", m_vrg_source_ip_3);
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_show_PLIC_state) $write(" %0d", m_vrg_source_ip_4);
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_show_PLIC_state) $write(" %0d", m_vrg_source_ip_5);
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_show_PLIC_state) $write(" %0d", m_vrg_source_ip_6);
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_show_PLIC_state) $write(" %0d", m_vrg_source_ip_7);
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_show_PLIC_state) $write(" %0d", m_vrg_source_ip_8);
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_show_PLIC_state) $write(" %0d", m_vrg_source_ip_9);
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_show_PLIC_state) $write(" %0d", m_vrg_source_ip_10);
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_show_PLIC_state) $write(" %0d", m_vrg_source_ip_11);
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_show_PLIC_state) $write(" %0d", m_vrg_source_ip_12);
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_show_PLIC_state) $write(" %0d", m_vrg_source_ip_13);
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_show_PLIC_state) $write(" %0d", m_vrg_source_ip_14);
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_show_PLIC_state) $write(" %0d", m_vrg_source_ip_15);
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_show_PLIC_state) $write(" %0d", m_vrg_source_ip_16);
    if (RST_N != `BSV_RESET_VALUE) if (EN_show_PLIC_state) $display("");
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_show_PLIC_state) $write("Src Prios:");
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_show_PLIC_state) $write(" %0d", m_vrg_source_prio_0);
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_show_PLIC_state) $write(" %0d", m_vrg_source_prio_1);
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_show_PLIC_state) $write(" %0d", m_vrg_source_prio_2);
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_show_PLIC_state) $write(" %0d", m_vrg_source_prio_3);
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_show_PLIC_state) $write(" %0d", m_vrg_source_prio_4);
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_show_PLIC_state) $write(" %0d", m_vrg_source_prio_5);
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_show_PLIC_state) $write(" %0d", m_vrg_source_prio_6);
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_show_PLIC_state) $write(" %0d", m_vrg_source_prio_7);
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_show_PLIC_state) $write(" %0d", m_vrg_source_prio_8);
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_show_PLIC_state) $write(" %0d", m_vrg_source_prio_9);
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_show_PLIC_state) $write(" %0d", m_vrg_source_prio_10);
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_show_PLIC_state) $write(" %0d", m_vrg_source_prio_11);
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_show_PLIC_state) $write(" %0d", m_vrg_source_prio_12);
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_show_PLIC_state) $write(" %0d", m_vrg_source_prio_13);
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_show_PLIC_state) $write(" %0d", m_vrg_source_prio_14);
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_show_PLIC_state) $write(" %0d", m_vrg_source_prio_15);
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_show_PLIC_state) $write(" %0d", m_vrg_source_prio_16);
    if (RST_N != `BSV_RESET_VALUE) if (EN_show_PLIC_state) $display("");
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_show_PLIC_state) $write("Src busy :");
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_show_PLIC_state) $write(" %0d", m_vrg_source_busy_0);
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_show_PLIC_state) $write(" %0d", m_vrg_source_busy_1);
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_show_PLIC_state) $write(" %0d", m_vrg_source_busy_2);
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_show_PLIC_state) $write(" %0d", m_vrg_source_busy_3);
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_show_PLIC_state) $write(" %0d", m_vrg_source_busy_4);
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_show_PLIC_state) $write(" %0d", m_vrg_source_busy_5);
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_show_PLIC_state) $write(" %0d", m_vrg_source_busy_6);
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_show_PLIC_state) $write(" %0d", m_vrg_source_busy_7);
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_show_PLIC_state) $write(" %0d", m_vrg_source_busy_8);
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_show_PLIC_state) $write(" %0d", m_vrg_source_busy_9);
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_show_PLIC_state) $write(" %0d", m_vrg_source_busy_10);
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_show_PLIC_state) $write(" %0d", m_vrg_source_busy_11);
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_show_PLIC_state) $write(" %0d", m_vrg_source_busy_12);
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_show_PLIC_state) $write(" %0d", m_vrg_source_busy_13);
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_show_PLIC_state) $write(" %0d", m_vrg_source_busy_14);
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_show_PLIC_state) $write(" %0d", m_vrg_source_busy_15);
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_show_PLIC_state) $write(" %0d", m_vrg_source_busy_16);
    if (RST_N != `BSV_RESET_VALUE) if (EN_show_PLIC_state) $display("");
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_show_PLIC_state) $write("T %0d IEs  :", $signed(32'd0));
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_show_PLIC_state) $write(" %0d", m_vvrg_ie_0_0);
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_show_PLIC_state) $write(" %0d", m_vvrg_ie_0_1);
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_show_PLIC_state) $write(" %0d", m_vvrg_ie_0_2);
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_show_PLIC_state) $write(" %0d", m_vvrg_ie_0_3);
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_show_PLIC_state) $write(" %0d", m_vvrg_ie_0_4);
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_show_PLIC_state) $write(" %0d", m_vvrg_ie_0_5);
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_show_PLIC_state) $write(" %0d", m_vvrg_ie_0_6);
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_show_PLIC_state) $write(" %0d", m_vvrg_ie_0_7);
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_show_PLIC_state) $write(" %0d", m_vvrg_ie_0_8);
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_show_PLIC_state) $write(" %0d", m_vvrg_ie_0_9);
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_show_PLIC_state) $write(" %0d", m_vvrg_ie_0_10);
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_show_PLIC_state) $write(" %0d", m_vvrg_ie_0_11);
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_show_PLIC_state) $write(" %0d", m_vvrg_ie_0_12);
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_show_PLIC_state) $write(" %0d", m_vvrg_ie_0_13);
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_show_PLIC_state) $write(" %0d", m_vvrg_ie_0_14);
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_show_PLIC_state) $write(" %0d", m_vvrg_ie_0_15);
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_show_PLIC_state) $write(" %0d", m_vvrg_ie_0_16);
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_show_PLIC_state)
	$display(" MaxPri %0d, Thresh %0d, MaxId %0d",
		 a__h81740,
		 m_vrg_target_threshold_0,
		 b__h81741);
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_show_PLIC_state) $write("T %0d IEs  :", $signed(32'd1));
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_show_PLIC_state) $write(" %0d", m_vvrg_ie_1_0);
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_show_PLIC_state) $write(" %0d", m_vvrg_ie_1_1);
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_show_PLIC_state) $write(" %0d", m_vvrg_ie_1_2);
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_show_PLIC_state) $write(" %0d", m_vvrg_ie_1_3);
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_show_PLIC_state) $write(" %0d", m_vvrg_ie_1_4);
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_show_PLIC_state) $write(" %0d", m_vvrg_ie_1_5);
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_show_PLIC_state) $write(" %0d", m_vvrg_ie_1_6);
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_show_PLIC_state) $write(" %0d", m_vvrg_ie_1_7);
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_show_PLIC_state) $write(" %0d", m_vvrg_ie_1_8);
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_show_PLIC_state) $write(" %0d", m_vvrg_ie_1_9);
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_show_PLIC_state) $write(" %0d", m_vvrg_ie_1_10);
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_show_PLIC_state) $write(" %0d", m_vvrg_ie_1_11);
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_show_PLIC_state) $write(" %0d", m_vvrg_ie_1_12);
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_show_PLIC_state) $write(" %0d", m_vvrg_ie_1_13);
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_show_PLIC_state) $write(" %0d", m_vvrg_ie_1_14);
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_show_PLIC_state) $write(" %0d", m_vvrg_ie_1_15);
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_show_PLIC_state) $write(" %0d", m_vvrg_ie_1_16);
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_show_PLIC_state)
	$display(" MaxPri %0d, Thresh %0d, MaxId %0d",
		 a__h83894,
		 m_vrg_target_threshold_1,
		 b__h83895);
    if (RST_N != `BSV_RESET_VALUE)
      if (NOT_m_vrg_source_busy_1_974_213_AND_NOT_m_cfg__ETC___d3217)
	begin
	  v__h86248 = $stime;
	  #0;
	end
    v__h86242 = v__h86248 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (NOT_m_vrg_source_busy_1_974_213_AND_NOT_m_cfg__ETC___d3217)
	$display("%0d: %m.m_interrupt_req: changing vrg_source_ip [%0d] to %0d",
		 v__h86242,
		 $signed(32'd1),
		 v_sources_0_m_interrupt_req_set_not_clear);
    if (RST_N != `BSV_RESET_VALUE)
      if (NOT_m_vrg_source_busy_2_975_220_AND_NOT_m_cfg__ETC___d3224)
	begin
	  v__h86443 = $stime;
	  #0;
	end
    v__h86437 = v__h86443 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (NOT_m_vrg_source_busy_2_975_220_AND_NOT_m_cfg__ETC___d3224)
	$display("%0d: %m.m_interrupt_req: changing vrg_source_ip [%0d] to %0d",
		 v__h86437,
		 $signed(32'd2),
		 v_sources_1_m_interrupt_req_set_not_clear);
    if (RST_N != `BSV_RESET_VALUE)
      if (NOT_m_vrg_source_busy_3_976_228_AND_NOT_m_cfg__ETC___d3232)
	begin
	  v__h86638 = $stime;
	  #0;
	end
    v__h86632 = v__h86638 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (NOT_m_vrg_source_busy_3_976_228_AND_NOT_m_cfg__ETC___d3232)
	$display("%0d: %m.m_interrupt_req: changing vrg_source_ip [%0d] to %0d",
		 v__h86632,
		 $signed(32'd3),
		 v_sources_2_m_interrupt_req_set_not_clear);
    if (RST_N != `BSV_RESET_VALUE)
      if (NOT_m_vrg_source_busy_4_977_236_AND_NOT_m_cfg__ETC___d3240)
	begin
	  v__h86833 = $stime;
	  #0;
	end
    v__h86827 = v__h86833 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (NOT_m_vrg_source_busy_4_977_236_AND_NOT_m_cfg__ETC___d3240)
	$display("%0d: %m.m_interrupt_req: changing vrg_source_ip [%0d] to %0d",
		 v__h86827,
		 $signed(32'd4),
		 v_sources_3_m_interrupt_req_set_not_clear);
    if (RST_N != `BSV_RESET_VALUE)
      if (NOT_m_vrg_source_busy_5_978_244_AND_NOT_m_cfg__ETC___d3248)
	begin
	  v__h87028 = $stime;
	  #0;
	end
    v__h87022 = v__h87028 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (NOT_m_vrg_source_busy_5_978_244_AND_NOT_m_cfg__ETC___d3248)
	$display("%0d: %m.m_interrupt_req: changing vrg_source_ip [%0d] to %0d",
		 v__h87022,
		 $signed(32'd5),
		 v_sources_4_m_interrupt_req_set_not_clear);
    if (RST_N != `BSV_RESET_VALUE)
      if (NOT_m_vrg_source_busy_6_979_252_AND_NOT_m_cfg__ETC___d3256)
	begin
	  v__h87223 = $stime;
	  #0;
	end
    v__h87217 = v__h87223 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (NOT_m_vrg_source_busy_6_979_252_AND_NOT_m_cfg__ETC___d3256)
	$display("%0d: %m.m_interrupt_req: changing vrg_source_ip [%0d] to %0d",
		 v__h87217,
		 $signed(32'd6),
		 v_sources_5_m_interrupt_req_set_not_clear);
    if (RST_N != `BSV_RESET_VALUE)
      if (NOT_m_vrg_source_busy_7_980_260_AND_NOT_m_cfg__ETC___d3264)
	begin
	  v__h87418 = $stime;
	  #0;
	end
    v__h87412 = v__h87418 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (NOT_m_vrg_source_busy_7_980_260_AND_NOT_m_cfg__ETC___d3264)
	$display("%0d: %m.m_interrupt_req: changing vrg_source_ip [%0d] to %0d",
		 v__h87412,
		 $signed(32'd7),
		 v_sources_6_m_interrupt_req_set_not_clear);
    if (RST_N != `BSV_RESET_VALUE)
      if (NOT_m_vrg_source_busy_8_981_268_AND_NOT_m_cfg__ETC___d3272)
	begin
	  v__h87613 = $stime;
	  #0;
	end
    v__h87607 = v__h87613 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (NOT_m_vrg_source_busy_8_981_268_AND_NOT_m_cfg__ETC___d3272)
	$display("%0d: %m.m_interrupt_req: changing vrg_source_ip [%0d] to %0d",
		 v__h87607,
		 $signed(32'd8),
		 v_sources_7_m_interrupt_req_set_not_clear);
    if (RST_N != `BSV_RESET_VALUE)
      if (NOT_m_vrg_source_busy_9_982_276_AND_NOT_m_cfg__ETC___d3280)
	begin
	  v__h87808 = $stime;
	  #0;
	end
    v__h87802 = v__h87808 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (NOT_m_vrg_source_busy_9_982_276_AND_NOT_m_cfg__ETC___d3280)
	$display("%0d: %m.m_interrupt_req: changing vrg_source_ip [%0d] to %0d",
		 v__h87802,
		 $signed(32'd9),
		 v_sources_8_m_interrupt_req_set_not_clear);
    if (RST_N != `BSV_RESET_VALUE)
      if (NOT_m_vrg_source_busy_10_983_284_AND_NOT_m_cfg_ETC___d3288)
	begin
	  v__h88003 = $stime;
	  #0;
	end
    v__h87997 = v__h88003 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (NOT_m_vrg_source_busy_10_983_284_AND_NOT_m_cfg_ETC___d3288)
	$display("%0d: %m.m_interrupt_req: changing vrg_source_ip [%0d] to %0d",
		 v__h87997,
		 $signed(32'd10),
		 v_sources_9_m_interrupt_req_set_not_clear);
    if (RST_N != `BSV_RESET_VALUE)
      if (NOT_m_vrg_source_busy_11_984_292_AND_NOT_m_cfg_ETC___d3296)
	begin
	  v__h88198 = $stime;
	  #0;
	end
    v__h88192 = v__h88198 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (NOT_m_vrg_source_busy_11_984_292_AND_NOT_m_cfg_ETC___d3296)
	$display("%0d: %m.m_interrupt_req: changing vrg_source_ip [%0d] to %0d",
		 v__h88192,
		 $signed(32'd11),
		 v_sources_10_m_interrupt_req_set_not_clear);
    if (RST_N != `BSV_RESET_VALUE)
      if (NOT_m_vrg_source_busy_12_985_300_AND_NOT_m_cfg_ETC___d3304)
	begin
	  v__h88393 = $stime;
	  #0;
	end
    v__h88387 = v__h88393 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (NOT_m_vrg_source_busy_12_985_300_AND_NOT_m_cfg_ETC___d3304)
	$display("%0d: %m.m_interrupt_req: changing vrg_source_ip [%0d] to %0d",
		 v__h88387,
		 $signed(32'd12),
		 v_sources_11_m_interrupt_req_set_not_clear);
    if (RST_N != `BSV_RESET_VALUE)
      if (NOT_m_vrg_source_busy_13_986_308_AND_NOT_m_cfg_ETC___d3312)
	begin
	  v__h88588 = $stime;
	  #0;
	end
    v__h88582 = v__h88588 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (NOT_m_vrg_source_busy_13_986_308_AND_NOT_m_cfg_ETC___d3312)
	$display("%0d: %m.m_interrupt_req: changing vrg_source_ip [%0d] to %0d",
		 v__h88582,
		 $signed(32'd13),
		 v_sources_12_m_interrupt_req_set_not_clear);
    if (RST_N != `BSV_RESET_VALUE)
      if (NOT_m_vrg_source_busy_14_987_316_AND_NOT_m_cfg_ETC___d3320)
	begin
	  v__h88783 = $stime;
	  #0;
	end
    v__h88777 = v__h88783 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (NOT_m_vrg_source_busy_14_987_316_AND_NOT_m_cfg_ETC___d3320)
	$display("%0d: %m.m_interrupt_req: changing vrg_source_ip [%0d] to %0d",
		 v__h88777,
		 $signed(32'd14),
		 v_sources_13_m_interrupt_req_set_not_clear);
    if (RST_N != `BSV_RESET_VALUE)
      if (NOT_m_vrg_source_busy_15_988_324_AND_NOT_m_cfg_ETC___d3328)
	begin
	  v__h88978 = $stime;
	  #0;
	end
    v__h88972 = v__h88978 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (NOT_m_vrg_source_busy_15_988_324_AND_NOT_m_cfg_ETC___d3328)
	$display("%0d: %m.m_interrupt_req: changing vrg_source_ip [%0d] to %0d",
		 v__h88972,
		 $signed(32'd15),
		 v_sources_14_m_interrupt_req_set_not_clear);
    if (RST_N != `BSV_RESET_VALUE)
      if (NOT_m_vrg_source_busy_16_989_332_AND_NOT_m_cfg_ETC___d3336)
	begin
	  v__h89173 = $stime;
	  #0;
	end
    v__h89167 = v__h89173 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (NOT_m_vrg_source_busy_16_989_332_AND_NOT_m_cfg_ETC___d3336)
	$display("%0d: %m.m_interrupt_req: changing vrg_source_ip [%0d] to %0d",
		 v__h89167,
		 $signed(32'd16),
		 v_sources_15_m_interrupt_req_set_not_clear);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_reset && m_cfg_verbosity != 4'd0)
	begin
	  v__h5962 = $stime;
	  #0;
	end
    v__h5956 = v__h5962 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_reset && m_cfg_verbosity != 4'd0)
	$display("%0d: PLIC.rl_reset", v__h5956);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	begin
	  v__h13331 = $stime;
	  #0;
	end
    v__h13325 = v__h13331 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$display("%0d: PLIC.rl_process_rd_req:", v__h13325);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write("    ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write("AXI4_Rd_Addr { ", "arid: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write("'h%h", m_slave_xactor_f_rd_addr$D_OUT[96:93]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write(", ", "araddr: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write("'h%h", m_slave_xactor_f_rd_addr$D_OUT[92:29]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write(", ", "arlen: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write("'h%h", m_slave_xactor_f_rd_addr$D_OUT[28:21]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write(", ", "arsize: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write("'h%h", m_slave_xactor_f_rd_addr$D_OUT[20:18]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write(", ", "arburst: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write("'h%h", m_slave_xactor_f_rd_addr$D_OUT[17:16]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write(", ", "arlock: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write("'h%h", m_slave_xactor_f_rd_addr$D_OUT[15]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write(", ", "arcache: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write("'h%h", m_slave_xactor_f_rd_addr$D_OUT[14:11]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write(", ", "arprot: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write("'h%h", m_slave_xactor_f_rd_addr$D_OUT[10:8]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write(", ", "arqos: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write("'h%h", m_slave_xactor_f_rd_addr$D_OUT[7:4]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write(", ", "arregion: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write("'h%h", m_slave_xactor_f_rd_addr$D_OUT[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write(", ", "aruser: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write("'h%h", 1'd0, " }");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write("\n");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d31)
	begin
	  v__h13514 = $stime;
	  #0;
	end
    v__h13508 = v__h13514 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d31)
	$display("%0d: ERROR: PLIC.rl_process_rd_req: unrecognized addr",
		 v__h13508);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d31)
	$write("            ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d31)
	$write("AXI4_Rd_Addr { ", "arid: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d31)
	$write("'h%h", m_slave_xactor_f_rd_addr$D_OUT[96:93]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d31)
	$write(", ", "araddr: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d31)
	$write("'h%h", m_slave_xactor_f_rd_addr$D_OUT[92:29]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d31)
	$write(", ", "arlen: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d31)
	$write("'h%h", m_slave_xactor_f_rd_addr$D_OUT[28:21]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d31)
	$write(", ", "arsize: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d31)
	$write("'h%h", m_slave_xactor_f_rd_addr$D_OUT[20:18]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d31)
	$write(", ", "arburst: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d31)
	$write("'h%h", m_slave_xactor_f_rd_addr$D_OUT[17:16]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d31)
	$write(", ", "arlock: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d31)
	$write("'h%h", m_slave_xactor_f_rd_addr$D_OUT[15]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d31)
	$write(", ", "arcache: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d31)
	$write("'h%h", m_slave_xactor_f_rd_addr$D_OUT[14:11]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d31)
	$write(", ", "arprot: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d31)
	$write("'h%h", m_slave_xactor_f_rd_addr$D_OUT[10:8]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d31)
	$write(", ", "arqos: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d31)
	$write("'h%h", m_slave_xactor_f_rd_addr$D_OUT[7:4]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d31)
	$write(", ", "arregion: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d31)
	$write("'h%h", m_slave_xactor_f_rd_addr$D_OUT[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d31)
	$write(", ", "aruser: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d31)
	$write("'h%h", 1'd0, " }");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d31)
	$write("\n");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  !m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d31 &&
	  m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d43)
	begin
	  v__h13730 = $stime;
	  #0;
	end
    v__h13724 = v__h13730 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  !m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d31 &&
	  m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d43)
	$display("%0d: PLIC.rl_process_rd_req: reading Source Priority: source %0d = 0x%0h",
		 v__h13724,
		 addr_offset__h13465[11:2],
		 v__h13689);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  !m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d31 &&
	  NOT_m_slave_xactor_f_rd_addr_first__9_BITS_92__ETC___d74)
	begin
	  v__h13976 = $stime;
	  #0;
	end
    v__h13970 = v__h13976 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  !m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d31 &&
	  NOT_m_slave_xactor_f_rd_addr_first__9_BITS_92__ETC___d74)
	$display("%0d: PLIC.rl_process_rd_req: reading Intr Pending 32 bits from source %0d = 0x%0h",
		 v__h13970,
		 source_id_base__h13893,
		 v__h13934);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  NOT_m_slave_xactor_f_rd_addr_first__9_BITS_92__ETC___d248)
	begin
	  v__h18445 = $stime;
	  #0;
	end
    v__h18439 = v__h18445 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  NOT_m_slave_xactor_f_rd_addr_first__9_BITS_92__ETC___d248)
	$display("%0d: PLIC.rl_process_rd_req: reading Intr Enable 32 bits from source %0d = 0x%0h",
		 v__h18439,
		 source_id_base__h13893,
		 v__h18403);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  NOT_m_slave_xactor_f_rd_addr_first__9_BITS_92__ETC___d538)
	begin
	  v__h24057 = $stime;
	  #0;
	end
    v__h24051 = v__h24057 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  NOT_m_slave_xactor_f_rd_addr_first__9_BITS_92__ETC___d538)
	$display("%0d: PLIC.rl_process_rd_req: reading Threshold for target %0d = 0x%0h",
		 v__h24051,
		 addr_offset__h13465[16:12],
		 v__h24016);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  NOT_m_slave_xactor_f_rd_addr_first__9_BITS_92__ETC___d733)
	begin
	  v__h26355 = $stime;
	  #0;
	end
    v__h26349 = v__h26355 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  NOT_m_slave_xactor_f_rd_addr_first__9_BITS_92__ETC___d733)
	$display("%0d: PLIC.rl_process_rd_req: reading Claim for target %0d = 0x%0h",
		 v__h26349,
		 addr_offset__h13465[16:12],
		 v__h24251);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  (m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d31 ||
	   IF_m_slave_xactor_f_rd_addr_first__9_BITS_92_T_ETC___d750))
	begin
	  v__h26568 = $stime;
	  #0;
	end
    v__h26562 = v__h26568 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  (m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d31 ||
	   IF_m_slave_xactor_f_rd_addr_first__9_BITS_92_T_ETC___d750))
	$display("%0d: ERROR: PLIC.rl_process_rd_req: unrecognized addr",
		 v__h26562);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  (m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d31 ||
	   IF_m_slave_xactor_f_rd_addr_first__9_BITS_92_T_ETC___d750))
	$write("            ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  (m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d31 ||
	   IF_m_slave_xactor_f_rd_addr_first__9_BITS_92_T_ETC___d750))
	$write("AXI4_Rd_Addr { ", "arid: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  (m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d31 ||
	   IF_m_slave_xactor_f_rd_addr_first__9_BITS_92_T_ETC___d750))
	$write("'h%h", m_slave_xactor_f_rd_addr$D_OUT[96:93]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  (m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d31 ||
	   IF_m_slave_xactor_f_rd_addr_first__9_BITS_92_T_ETC___d750))
	$write(", ", "araddr: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  (m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d31 ||
	   IF_m_slave_xactor_f_rd_addr_first__9_BITS_92_T_ETC___d750))
	$write("'h%h", m_slave_xactor_f_rd_addr$D_OUT[92:29]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  (m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d31 ||
	   IF_m_slave_xactor_f_rd_addr_first__9_BITS_92_T_ETC___d750))
	$write(", ", "arlen: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  (m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d31 ||
	   IF_m_slave_xactor_f_rd_addr_first__9_BITS_92_T_ETC___d750))
	$write("'h%h", m_slave_xactor_f_rd_addr$D_OUT[28:21]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  (m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d31 ||
	   IF_m_slave_xactor_f_rd_addr_first__9_BITS_92_T_ETC___d750))
	$write(", ", "arsize: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  (m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d31 ||
	   IF_m_slave_xactor_f_rd_addr_first__9_BITS_92_T_ETC___d750))
	$write("'h%h", m_slave_xactor_f_rd_addr$D_OUT[20:18]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  (m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d31 ||
	   IF_m_slave_xactor_f_rd_addr_first__9_BITS_92_T_ETC___d750))
	$write(", ", "arburst: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  (m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d31 ||
	   IF_m_slave_xactor_f_rd_addr_first__9_BITS_92_T_ETC___d750))
	$write("'h%h", m_slave_xactor_f_rd_addr$D_OUT[17:16]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  (m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d31 ||
	   IF_m_slave_xactor_f_rd_addr_first__9_BITS_92_T_ETC___d750))
	$write(", ", "arlock: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  (m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d31 ||
	   IF_m_slave_xactor_f_rd_addr_first__9_BITS_92_T_ETC___d750))
	$write("'h%h", m_slave_xactor_f_rd_addr$D_OUT[15]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  (m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d31 ||
	   IF_m_slave_xactor_f_rd_addr_first__9_BITS_92_T_ETC___d750))
	$write(", ", "arcache: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  (m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d31 ||
	   IF_m_slave_xactor_f_rd_addr_first__9_BITS_92_T_ETC___d750))
	$write("'h%h", m_slave_xactor_f_rd_addr$D_OUT[14:11]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  (m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d31 ||
	   IF_m_slave_xactor_f_rd_addr_first__9_BITS_92_T_ETC___d750))
	$write(", ", "arprot: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  (m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d31 ||
	   IF_m_slave_xactor_f_rd_addr_first__9_BITS_92_T_ETC___d750))
	$write("'h%h", m_slave_xactor_f_rd_addr$D_OUT[10:8]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  (m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d31 ||
	   IF_m_slave_xactor_f_rd_addr_first__9_BITS_92_T_ETC___d750))
	$write(", ", "arqos: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  (m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d31 ||
	   IF_m_slave_xactor_f_rd_addr_first__9_BITS_92_T_ETC___d750))
	$write("'h%h", m_slave_xactor_f_rd_addr$D_OUT[7:4]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  (m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d31 ||
	   IF_m_slave_xactor_f_rd_addr_first__9_BITS_92_T_ETC___d750))
	$write(", ", "arregion: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  (m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d31 ||
	   IF_m_slave_xactor_f_rd_addr_first__9_BITS_92_T_ETC___d750))
	$write("'h%h", m_slave_xactor_f_rd_addr$D_OUT[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  (m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d31 ||
	   IF_m_slave_xactor_f_rd_addr_first__9_BITS_92_T_ETC___d750))
	$write(", ", "aruser: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  (m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d31 ||
	   IF_m_slave_xactor_f_rd_addr_first__9_BITS_92_T_ETC___d750))
	$write("'h%h", 1'd0, " }");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  (m_slave_xactor_f_rd_addr_first__9_BITS_92_TO_2_ETC___d31 ||
	   IF_m_slave_xactor_f_rd_addr_first__9_BITS_92_T_ETC___d750))
	$write("\n");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	begin
	  v__h26773 = $stime;
	  #0;
	end
    v__h26767 = v__h26773 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$display("%0d: PLIC.rl_process_rd_req", v__h26767);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write("            ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write("AXI4_Rd_Addr { ", "arid: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write("'h%h", m_slave_xactor_f_rd_addr$D_OUT[96:93]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write(", ", "araddr: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write("'h%h", m_slave_xactor_f_rd_addr$D_OUT[92:29]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write(", ", "arlen: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write("'h%h", m_slave_xactor_f_rd_addr$D_OUT[28:21]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write(", ", "arsize: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write("'h%h", m_slave_xactor_f_rd_addr$D_OUT[20:18]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write(", ", "arburst: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write("'h%h", m_slave_xactor_f_rd_addr$D_OUT[17:16]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write(", ", "arlock: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write("'h%h", m_slave_xactor_f_rd_addr$D_OUT[15]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write(", ", "arcache: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write("'h%h", m_slave_xactor_f_rd_addr$D_OUT[14:11]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write(", ", "arprot: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write("'h%h", m_slave_xactor_f_rd_addr$D_OUT[10:8]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write(", ", "arqos: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write("'h%h", m_slave_xactor_f_rd_addr$D_OUT[7:4]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write(", ", "arregion: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write("'h%h", m_slave_xactor_f_rd_addr$D_OUT[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write(", ", "aruser: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write("'h%h", 1'd0, " }");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write("\n");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write("            ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write("AXI4_Rd_Data { ", "rid: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write("'h%h", m_slave_xactor_f_rd_addr$D_OUT[96:93]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write(", ", "rdata: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write("'h%h", x__h26677);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write(", ", "rresp: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write("'h%h", rresp__h26521);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write(", ", "rlast: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write("True");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write(", ", "ruser: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write("'h%h", 1'd0, " }");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_rd_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write("\n");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	begin
	  v__h27053 = $stime;
	  #0;
	end
    v__h27047 = v__h27053 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$display("%0d: PLIC.rl_process_wr_req", v__h27047);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write("    ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write("AXI4_Wr_Addr { ", "awid: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write("'h%h", m_slave_xactor_f_wr_addr$D_OUT[96:93]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write(", ", "awaddr: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write("'h%h", m_slave_xactor_f_wr_addr$D_OUT[92:29]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write(", ", "awlen: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write("'h%h", m_slave_xactor_f_wr_addr$D_OUT[28:21]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write(", ", "awsize: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write("'h%h", m_slave_xactor_f_wr_addr$D_OUT[20:18]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write(", ", "awburst: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write("'h%h", m_slave_xactor_f_wr_addr$D_OUT[17:16]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write(", ", "awlock: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write("'h%h", m_slave_xactor_f_wr_addr$D_OUT[15]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write(", ", "awcache: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write("'h%h", m_slave_xactor_f_wr_addr$D_OUT[14:11]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write(", ", "awprot: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write("'h%h", m_slave_xactor_f_wr_addr$D_OUT[10:8]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write(", ", "awqos: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write("'h%h", m_slave_xactor_f_wr_addr$D_OUT[7:4]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write(", ", "awregion: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write("'h%h", m_slave_xactor_f_wr_addr$D_OUT[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write(", ", "awuser: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write("'h%h", 1'd0, " }");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write("\n");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write("    ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write("AXI4_Wr_Data { ", "wdata: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write("'h%h", m_slave_xactor_f_wr_data$D_OUT[72:9]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write(", ", "wstrb: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write("'h%h", m_slave_xactor_f_wr_data$D_OUT[8:1]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write(", ", "wlast: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16 &&
	  m_slave_xactor_f_wr_data$D_OUT[0])
	$write("True");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16 &&
	  !m_slave_xactor_f_wr_data$D_OUT[0])
	$write("False");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write(", ", "wuser: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write("'h%h", 1'd0, " }");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write("\n");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812)
	begin
	  v__h27284 = $stime;
	  #0;
	end
    v__h27278 = v__h27284 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812)
	$display("%0d: ERROR: PLIC.rl_process_wr_req: unrecognized addr",
		 v__h27278);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812)
	$write("            ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812)
	$write("AXI4_Wr_Addr { ", "awid: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812)
	$write("'h%h", m_slave_xactor_f_wr_addr$D_OUT[96:93]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812)
	$write(", ", "awaddr: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812)
	$write("'h%h", m_slave_xactor_f_wr_addr$D_OUT[92:29]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812)
	$write(", ", "awlen: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812)
	$write("'h%h", m_slave_xactor_f_wr_addr$D_OUT[28:21]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812)
	$write(", ", "awsize: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812)
	$write("'h%h", m_slave_xactor_f_wr_addr$D_OUT[20:18]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812)
	$write(", ", "awburst: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812)
	$write("'h%h", m_slave_xactor_f_wr_addr$D_OUT[17:16]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812)
	$write(", ", "awlock: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812)
	$write("'h%h", m_slave_xactor_f_wr_addr$D_OUT[15]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812)
	$write(", ", "awcache: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812)
	$write("'h%h", m_slave_xactor_f_wr_addr$D_OUT[14:11]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812)
	$write(", ", "awprot: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812)
	$write("'h%h", m_slave_xactor_f_wr_addr$D_OUT[10:8]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812)
	$write(", ", "awqos: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812)
	$write("'h%h", m_slave_xactor_f_wr_addr$D_OUT[7:4]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812)
	$write(", ", "awregion: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812)
	$write("'h%h", m_slave_xactor_f_wr_addr$D_OUT[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812)
	$write(", ", "awuser: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812)
	$write("'h%h", 1'd0, " }");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812)
	$write("\n");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812)
	$write("            ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812)
	$write("AXI4_Wr_Data { ", "wdata: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812)
	$write("'h%h", m_slave_xactor_f_wr_data$D_OUT[72:9]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812)
	$write(", ", "wstrb: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812)
	$write("'h%h", m_slave_xactor_f_wr_data$D_OUT[8:1]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812)
	$write(", ", "wlast: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 &&
	  m_slave_xactor_f_wr_data$D_OUT[0])
	$write("True");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 &&
	  !m_slave_xactor_f_wr_data$D_OUT[0])
	$write("False");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812)
	$write(", ", "wuser: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812)
	$write("'h%h", 1'd0, " }");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812)
	$write("\n");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 &&
	  m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d869)
	begin
	  v__h28359 = $stime;
	  #0;
	end
    v__h28353 = v__h28359 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 &&
	  m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d869)
	$display("%0d: PLIC.rl_process_wr_req: writing Source Priority: source %0d = 0x%0h",
		 v__h28353,
		 addr_offset__h27245[11:2],
		 wdata32__h27246);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 &&
	  NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d880)
	begin
	  v__h28531 = $stime;
	  #0;
	end
    v__h28525 = v__h28531 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 &&
	  NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d880)
	$display("%0d: PLIC.rl_process_wr_req: Ignoring write to Read-only Intr Pending 32 bits from source %0d",
		 v__h28525,
		 source_id_base__h28620);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2844)
	begin
	  v__h76647 = $stime;
	  #0;
	end
    v__h76641 = v__h76647 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2844)
	$display("%0d: PLIC.rl_process_wr_req: writing Intr Enable 32 bits for target %0d from source %0d = 0x%0h",
		 v__h76641,
		 addr_offset__h27245[11:7],
		 source_id_base__h28620,
		 wdata32__h27246);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2868)
	begin
	  v__h76947 = $stime;
	  #0;
	end
    v__h76941 = v__h76947 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2868)
	$display("%0d: PLIC.rl_process_wr_req: writing threshold for target %0d = 0x%0h",
		 v__h76941,
		 addr_offset__h27245[16:12],
		 wdata32__h27246);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 &&
	  !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d821 &&
	  NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2923)
	begin
	  v__h77579 = $stime;
	  #0;
	end
    v__h77573 = v__h77579 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 &&
	  !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d821 &&
	  NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2923)
	$display("%0d: PLIC.rl_process_wr_req: writing completion for target %0d for source 0x%0h",
		 v__h77573,
		 addr_offset__h27245[16:12],
		 wdata32__h27246[9:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 &&
	  !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d821 &&
	  NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2935)
	begin
	  v__h77673 = $stime;
	  #0;
	end
    v__h77667 = v__h77673 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 &&
	  !m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d821 &&
	  NOT_m_slave_xactor_f_wr_addr_first__94_BITS_92_ETC___d2935)
	$display("%0d: PLIC.rl_process_wr_req: ignoring completion for target %0d for source 0x%0h",
		 v__h77667,
		 addr_offset__h27245[16:12],
		 wdata32__h27246[9:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  (m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 ||
	   IF_m_slave_xactor_f_wr_addr_first__94_BITS_92__ETC___d2952))
	begin
	  v__h77844 = $stime;
	  #0;
	end
    v__h77838 = v__h77844 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  (m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 ||
	   IF_m_slave_xactor_f_wr_addr_first__94_BITS_92__ETC___d2952))
	$display("%0d: ERROR: PLIC.rl_process_wr_req: unrecognized addr",
		 v__h77838);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  (m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 ||
	   IF_m_slave_xactor_f_wr_addr_first__94_BITS_92__ETC___d2952))
	$write("            ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  (m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 ||
	   IF_m_slave_xactor_f_wr_addr_first__94_BITS_92__ETC___d2952))
	$write("AXI4_Wr_Addr { ", "awid: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  (m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 ||
	   IF_m_slave_xactor_f_wr_addr_first__94_BITS_92__ETC___d2952))
	$write("'h%h", m_slave_xactor_f_wr_addr$D_OUT[96:93]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  (m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 ||
	   IF_m_slave_xactor_f_wr_addr_first__94_BITS_92__ETC___d2952))
	$write(", ", "awaddr: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  (m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 ||
	   IF_m_slave_xactor_f_wr_addr_first__94_BITS_92__ETC___d2952))
	$write("'h%h", m_slave_xactor_f_wr_addr$D_OUT[92:29]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  (m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 ||
	   IF_m_slave_xactor_f_wr_addr_first__94_BITS_92__ETC___d2952))
	$write(", ", "awlen: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  (m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 ||
	   IF_m_slave_xactor_f_wr_addr_first__94_BITS_92__ETC___d2952))
	$write("'h%h", m_slave_xactor_f_wr_addr$D_OUT[28:21]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  (m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 ||
	   IF_m_slave_xactor_f_wr_addr_first__94_BITS_92__ETC___d2952))
	$write(", ", "awsize: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  (m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 ||
	   IF_m_slave_xactor_f_wr_addr_first__94_BITS_92__ETC___d2952))
	$write("'h%h", m_slave_xactor_f_wr_addr$D_OUT[20:18]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  (m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 ||
	   IF_m_slave_xactor_f_wr_addr_first__94_BITS_92__ETC___d2952))
	$write(", ", "awburst: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  (m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 ||
	   IF_m_slave_xactor_f_wr_addr_first__94_BITS_92__ETC___d2952))
	$write("'h%h", m_slave_xactor_f_wr_addr$D_OUT[17:16]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  (m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 ||
	   IF_m_slave_xactor_f_wr_addr_first__94_BITS_92__ETC___d2952))
	$write(", ", "awlock: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  (m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 ||
	   IF_m_slave_xactor_f_wr_addr_first__94_BITS_92__ETC___d2952))
	$write("'h%h", m_slave_xactor_f_wr_addr$D_OUT[15]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  (m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 ||
	   IF_m_slave_xactor_f_wr_addr_first__94_BITS_92__ETC___d2952))
	$write(", ", "awcache: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  (m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 ||
	   IF_m_slave_xactor_f_wr_addr_first__94_BITS_92__ETC___d2952))
	$write("'h%h", m_slave_xactor_f_wr_addr$D_OUT[14:11]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  (m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 ||
	   IF_m_slave_xactor_f_wr_addr_first__94_BITS_92__ETC___d2952))
	$write(", ", "awprot: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  (m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 ||
	   IF_m_slave_xactor_f_wr_addr_first__94_BITS_92__ETC___d2952))
	$write("'h%h", m_slave_xactor_f_wr_addr$D_OUT[10:8]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  (m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 ||
	   IF_m_slave_xactor_f_wr_addr_first__94_BITS_92__ETC___d2952))
	$write(", ", "awqos: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  (m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 ||
	   IF_m_slave_xactor_f_wr_addr_first__94_BITS_92__ETC___d2952))
	$write("'h%h", m_slave_xactor_f_wr_addr$D_OUT[7:4]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  (m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 ||
	   IF_m_slave_xactor_f_wr_addr_first__94_BITS_92__ETC___d2952))
	$write(", ", "awregion: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  (m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 ||
	   IF_m_slave_xactor_f_wr_addr_first__94_BITS_92__ETC___d2952))
	$write("'h%h", m_slave_xactor_f_wr_addr$D_OUT[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  (m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 ||
	   IF_m_slave_xactor_f_wr_addr_first__94_BITS_92__ETC___d2952))
	$write(", ", "awuser: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  (m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 ||
	   IF_m_slave_xactor_f_wr_addr_first__94_BITS_92__ETC___d2952))
	$write("'h%h", 1'd0, " }");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  (m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 ||
	   IF_m_slave_xactor_f_wr_addr_first__94_BITS_92__ETC___d2952))
	$write("\n");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  (m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 ||
	   IF_m_slave_xactor_f_wr_addr_first__94_BITS_92__ETC___d2952))
	$write("            ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  (m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 ||
	   IF_m_slave_xactor_f_wr_addr_first__94_BITS_92__ETC___d2952))
	$write("AXI4_Wr_Data { ", "wdata: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  (m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 ||
	   IF_m_slave_xactor_f_wr_addr_first__94_BITS_92__ETC___d2952))
	$write("'h%h", m_slave_xactor_f_wr_data$D_OUT[72:9]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  (m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 ||
	   IF_m_slave_xactor_f_wr_addr_first__94_BITS_92__ETC___d2952))
	$write(", ", "wstrb: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  (m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 ||
	   IF_m_slave_xactor_f_wr_addr_first__94_BITS_92__ETC___d2952))
	$write("'h%h", m_slave_xactor_f_wr_data$D_OUT[8:1]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  (m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 ||
	   IF_m_slave_xactor_f_wr_addr_first__94_BITS_92__ETC___d2952))
	$write(", ", "wlast: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  (m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 ||
	   IF_m_slave_xactor_f_wr_addr_first__94_BITS_92__ETC___d2952) &&
	  m_slave_xactor_f_wr_data$D_OUT[0])
	$write("True");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  (m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 ||
	   IF_m_slave_xactor_f_wr_addr_first__94_BITS_92__ETC___d2952) &&
	  !m_slave_xactor_f_wr_data$D_OUT[0])
	$write("False");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  (m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 ||
	   IF_m_slave_xactor_f_wr_addr_first__94_BITS_92__ETC___d2952))
	$write(", ", "wuser: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  (m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 ||
	   IF_m_slave_xactor_f_wr_addr_first__94_BITS_92__ETC___d2952))
	$write("'h%h", 1'd0, " }");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  (m_slave_xactor_f_wr_addr_first__94_BITS_92_TO__ETC___d812 ||
	   IF_m_slave_xactor_f_wr_addr_first__94_BITS_92__ETC___d2952))
	$write("\n");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	begin
	  v__h78064 = $stime;
	  #0;
	end
    v__h78058 = v__h78064 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$display("%0d: PLIC.AXI4.rl_process_wr_req", v__h78058);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write("            ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write("AXI4_Wr_Addr { ", "awid: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write("'h%h", m_slave_xactor_f_wr_addr$D_OUT[96:93]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write(", ", "awaddr: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write("'h%h", m_slave_xactor_f_wr_addr$D_OUT[92:29]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write(", ", "awlen: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write("'h%h", m_slave_xactor_f_wr_addr$D_OUT[28:21]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write(", ", "awsize: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write("'h%h", m_slave_xactor_f_wr_addr$D_OUT[20:18]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write(", ", "awburst: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write("'h%h", m_slave_xactor_f_wr_addr$D_OUT[17:16]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write(", ", "awlock: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write("'h%h", m_slave_xactor_f_wr_addr$D_OUT[15]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write(", ", "awcache: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write("'h%h", m_slave_xactor_f_wr_addr$D_OUT[14:11]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write(", ", "awprot: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write("'h%h", m_slave_xactor_f_wr_addr$D_OUT[10:8]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write(", ", "awqos: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write("'h%h", m_slave_xactor_f_wr_addr$D_OUT[7:4]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write(", ", "awregion: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write("'h%h", m_slave_xactor_f_wr_addr$D_OUT[3:0]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write(", ", "awuser: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write("'h%h", 1'd0, " }");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write("\n");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write("            ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write("AXI4_Wr_Data { ", "wdata: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write("'h%h", m_slave_xactor_f_wr_data$D_OUT[72:9]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write(", ", "wstrb: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write("'h%h", m_slave_xactor_f_wr_data$D_OUT[8:1]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write(", ", "wlast: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16 &&
	  m_slave_xactor_f_wr_data$D_OUT[0])
	$write("True");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16 &&
	  !m_slave_xactor_f_wr_data$D_OUT[0])
	$write("False");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write(", ", "wuser: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write("'h%h", 1'd0, " }");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write("\n");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write("            ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write("AXI4_Wr_Resp { ", "bid: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write("'h%h", m_slave_xactor_f_wr_addr$D_OUT[96:93]);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write(", ", "bresp: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write("'h%h", v__h27250);
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write(", ", "buser: ");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write("'h%h", 1'd0, " }");
    if (RST_N != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_m_rl_process_wr_req &&
	  NOT_m_cfg_verbosity_read_ULE_1_5___d16)
	$write("\n");
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_set_addr_map && set_addr_map_addr_base[1:0] != 2'd0)
	begin
	  v__h85245 = $stime;
	  #0;
	end
    v__h85239 = v__h85245 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_set_addr_map && set_addr_map_addr_base[1:0] != 2'd0)
	$display("%0d: WARNING: PLIC.set_addr_map: addr_base 0x%0h is not 4-Byte-aligned",
		 v__h85239,
		 set_addr_map_addr_base);
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_set_addr_map && set_addr_map_addr_lim[1:0] != 2'd0)
	begin
	  v__h85351 = $stime;
	  #0;
	end
    v__h85345 = v__h85351 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_set_addr_map && set_addr_map_addr_lim[1:0] != 2'd0)
	$display("%0d: WARNING: PLIC.set_addr_map: addr_lim 0x%0h is not 4-Byte-aligned",
		 v__h85345,
		 set_addr_map_addr_lim);
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_set_addr_map && m_cfg_verbosity != 4'd0)
	begin
	  v__h85478 = $stime;
	  #0;
	end
    v__h85472 = v__h85478 / 32'd10;
    if (RST_N != `BSV_RESET_VALUE)
      if (EN_set_addr_map && m_cfg_verbosity != 4'd0)
	$display("%0d: PLIC.set_addr_map: base 0x%0h limit 0x%0h",
		 v__h85472,
		 set_addr_map_addr_base,
		 set_addr_map_addr_lim);
  end
  // synopsys translate_on
endmodule