module be tested as is.
		reset = 0;
	end
endmodule