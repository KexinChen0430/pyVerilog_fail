module top(
  input [15:0] a,
  input [15:0] b,
  output [15:0] o
  );
  wire [0:0] CLBLL_L_X2Y23_SLICE_X0Y23_A;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X0Y23_A1;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X0Y23_A2;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X0Y23_A3;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X0Y23_A4;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X0Y23_A5;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X0Y23_A6;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X0Y23_AMUX;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X0Y23_AO5;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X0Y23_AO6;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X0Y23_AX;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X0Y23_A_CY;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X0Y23_A_XOR;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X0Y23_B;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X0Y23_B1;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X0Y23_B2;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X0Y23_B3;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X0Y23_B4;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X0Y23_B5;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X0Y23_B6;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X0Y23_BMUX;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X0Y23_BO5;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X0Y23_BO6;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X0Y23_BX;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X0Y23_B_CY;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X0Y23_B_XOR;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X0Y23_C;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X0Y23_C1;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X0Y23_C2;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X0Y23_C3;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X0Y23_C4;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X0Y23_C5;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X0Y23_C6;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X0Y23_CMUX;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X0Y23_CO5;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X0Y23_CO6;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X0Y23_COUT;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X0Y23_CX;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X0Y23_C_CY;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X0Y23_C_XOR;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X0Y23_D;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X0Y23_D1;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X0Y23_D2;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X0Y23_D3;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X0Y23_D4;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X0Y23_D5;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X0Y23_D6;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X0Y23_DMUX;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X0Y23_DO5;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X0Y23_DO6;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X0Y23_DX;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X0Y23_D_CY;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X0Y23_D_XOR;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X1Y23_A;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X1Y23_A1;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X1Y23_A2;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X1Y23_A3;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X1Y23_A4;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X1Y23_A5;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X1Y23_A6;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X1Y23_AO5;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X1Y23_AO6;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X1Y23_A_CY;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X1Y23_A_XOR;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X1Y23_B;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X1Y23_B1;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X1Y23_B2;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X1Y23_B3;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X1Y23_B4;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X1Y23_B5;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X1Y23_B6;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X1Y23_BO5;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X1Y23_BO6;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X1Y23_B_CY;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X1Y23_B_XOR;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X1Y23_C;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X1Y23_C1;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X1Y23_C2;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X1Y23_C3;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X1Y23_C4;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X1Y23_C5;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X1Y23_C6;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X1Y23_CO5;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X1Y23_CO6;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X1Y23_C_CY;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X1Y23_C_XOR;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X1Y23_D;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X1Y23_D1;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X1Y23_D2;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X1Y23_D3;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X1Y23_D4;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X1Y23_D5;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X1Y23_D6;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X1Y23_DO5;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X1Y23_DO6;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X1Y23_D_CY;
  wire [0:0] CLBLL_L_X2Y23_SLICE_X1Y23_D_XOR;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X0Y24_A;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X0Y24_A1;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X0Y24_A2;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X0Y24_A3;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X0Y24_A4;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X0Y24_A5;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X0Y24_A6;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X0Y24_AMUX;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X0Y24_AO5;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X0Y24_AO6;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X0Y24_AX;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X0Y24_A_CY;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X0Y24_A_XOR;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X0Y24_B;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X0Y24_B1;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X0Y24_B2;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X0Y24_B3;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X0Y24_B4;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X0Y24_B5;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X0Y24_B6;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X0Y24_BMUX;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X0Y24_BO5;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X0Y24_BO6;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X0Y24_BX;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X0Y24_B_CY;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X0Y24_B_XOR;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X0Y24_C;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X0Y24_C1;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X0Y24_C2;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X0Y24_C3;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X0Y24_C4;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X0Y24_C5;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X0Y24_C6;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X0Y24_CIN;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X0Y24_CMUX;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X0Y24_CO5;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X0Y24_CO6;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X0Y24_COUT;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X0Y24_CX;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X0Y24_C_CY;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X0Y24_C_XOR;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X0Y24_D;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X0Y24_D1;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X0Y24_D2;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X0Y24_D3;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X0Y24_D4;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X0Y24_D5;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X0Y24_D6;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X0Y24_DMUX;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X0Y24_DO5;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X0Y24_DO6;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X0Y24_DX;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X0Y24_D_CY;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X0Y24_D_XOR;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X1Y24_A;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X1Y24_A1;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X1Y24_A2;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X1Y24_A3;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X1Y24_A4;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X1Y24_A5;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X1Y24_A6;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X1Y24_AO5;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X1Y24_AO6;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X1Y24_A_CY;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X1Y24_A_XOR;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X1Y24_B;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X1Y24_B1;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X1Y24_B2;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X1Y24_B3;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X1Y24_B4;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X1Y24_B5;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X1Y24_B6;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X1Y24_BO5;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X1Y24_BO6;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X1Y24_B_CY;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X1Y24_B_XOR;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X1Y24_C;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X1Y24_C1;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X1Y24_C2;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X1Y24_C3;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X1Y24_C4;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X1Y24_C5;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X1Y24_C6;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X1Y24_CO5;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X1Y24_CO6;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X1Y24_C_CY;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X1Y24_C_XOR;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X1Y24_D;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X1Y24_D1;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X1Y24_D2;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X1Y24_D3;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X1Y24_D4;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X1Y24_D5;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X1Y24_D6;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X1Y24_DO5;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X1Y24_DO6;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X1Y24_D_CY;
  wire [0:0] CLBLL_L_X2Y24_SLICE_X1Y24_D_XOR;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X0Y25_A;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X0Y25_A1;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X0Y25_A2;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X0Y25_A3;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X0Y25_A4;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X0Y25_A5;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X0Y25_A6;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X0Y25_AMUX;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X0Y25_AO5;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X0Y25_AO6;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X0Y25_AX;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X0Y25_A_CY;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X0Y25_A_XOR;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X0Y25_B;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X0Y25_B1;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X0Y25_B2;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X0Y25_B3;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X0Y25_B4;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X0Y25_B5;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X0Y25_B6;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X0Y25_BMUX;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X0Y25_BO5;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X0Y25_BO6;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X0Y25_BX;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X0Y25_B_CY;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X0Y25_B_XOR;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X0Y25_C;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X0Y25_C1;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X0Y25_C2;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X0Y25_C3;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X0Y25_C4;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X0Y25_C5;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X0Y25_C6;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X0Y25_CIN;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X0Y25_CMUX;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X0Y25_CO5;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X0Y25_CO6;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X0Y25_COUT;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X0Y25_CX;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X0Y25_C_CY;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X0Y25_C_XOR;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X0Y25_D;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X0Y25_D1;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X0Y25_D2;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X0Y25_D3;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X0Y25_D4;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X0Y25_D5;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X0Y25_D6;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X0Y25_DMUX;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X0Y25_DO5;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X0Y25_DO6;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X0Y25_DX;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X0Y25_D_CY;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X0Y25_D_XOR;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X1Y25_A;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X1Y25_A1;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X1Y25_A2;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X1Y25_A3;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X1Y25_A4;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X1Y25_A5;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X1Y25_A6;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X1Y25_AO5;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X1Y25_AO6;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X1Y25_A_CY;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X1Y25_A_XOR;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X1Y25_B;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X1Y25_B1;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X1Y25_B2;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X1Y25_B3;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X1Y25_B4;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X1Y25_B5;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X1Y25_B6;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X1Y25_BO5;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X1Y25_BO6;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X1Y25_B_CY;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X1Y25_B_XOR;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X1Y25_C;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X1Y25_C1;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X1Y25_C2;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X1Y25_C3;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X1Y25_C4;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X1Y25_C5;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X1Y25_C6;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X1Y25_CO5;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X1Y25_CO6;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X1Y25_C_CY;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X1Y25_C_XOR;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X1Y25_D;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X1Y25_D1;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X1Y25_D2;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X1Y25_D3;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X1Y25_D4;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X1Y25_D5;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X1Y25_D6;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X1Y25_DO5;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X1Y25_DO6;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X1Y25_D_CY;
  wire [0:0] CLBLL_L_X2Y25_SLICE_X1Y25_D_XOR;
  wire [0:0] CLBLL_L_X2Y26_SLICE_X0Y26_A;
  wire [0:0] CLBLL_L_X2Y26_SLICE_X0Y26_A1;
  wire [0:0] CLBLL_L_X2Y26_SLICE_X0Y26_A2;
  wire [0:0] CLBLL_L_X2Y26_SLICE_X0Y26_A3;
  wire [0:0] CLBLL_L_X2Y26_SLICE_X0Y26_A4;
  wire [0:0] CLBLL_L_X2Y26_SLICE_X0Y26_A5;
  wire [0:0] CLBLL_L_X2Y26_SLICE_X0Y26_A6;
  wire [0:0] CLBLL_L_X2Y26_SLICE_X0Y26_AMUX;
  wire [0:0] CLBLL_L_X2Y26_SLICE_X0Y26_AO5;
  wire [0:0] CLBLL_L_X2Y26_SLICE_X0Y26_AO6;
  wire [0:0] CLBLL_L_X2Y26_SLICE_X0Y26_AX;
  wire [0:0] CLBLL_L_X2Y26_SLICE_X0Y26_A_CY;
  wire [0:0] CLBLL_L_X2Y26_SLICE_X0Y26_A_XOR;
  wire [0:0] CLBLL_L_X2Y26_SLICE_X0Y26_B;
  wire [0:0] CLBLL_L_X2Y26_SLICE_X0Y26_B1;
  wire [0:0] CLBLL_L_X2Y26_SLICE_X0Y26_B2;
  wire [0:0] CLBLL_L_X2Y26_SLICE_X0Y26_B3;
  wire [0:0] CLBLL_L_X2Y26_SLICE_X0Y26_B4;
  wire [0:0] CLBLL_L_X2Y26_SLICE_X0Y26_B5;
  wire [0:0] CLBLL_L_X2Y26_SLICE_X0Y26_B6;
  wire [0:0] CLBLL_L_X2Y26_SLICE_X0Y26_BMUX;
  wire [0:0] CLBLL_L_X2Y26_SLICE_X0Y26_BO5;
  wire [0:0] CLBLL_L_X2Y26_SLICE_X0Y26_BO6;
  wire [0:0] CLBLL_L_X2Y26_SLICE_X0Y26_BX;
  wire [0:0] CLBLL_L_X2Y26_SLICE_X0Y26_B_CY;
  wire [0:0] CLBLL_L_X2Y26_SLICE_X0Y26_B_XOR;
  wire [0:0] CLBLL_L_X2Y26_SLICE_X0Y26_C;
  wire [0:0] CLBLL_L_X2Y26_SLICE_X0Y26_C1;
  wire [0:0] CLBLL_L_X2Y26_SLICE_X0Y26_C2;
  wire [0:0] CLBLL_L_X2Y26_SLICE_X0Y26_C3;
  wire [0:0] CLBLL_L_X2Y26_SLICE_X0Y26_C4;
  wire [0:0] CLBLL_L_X2Y26_SLICE_X0Y26_C5;
  wire [0:0] CLBLL_L_X2Y26_SLICE_X0Y26_C6;
  wire [0:0] CLBLL_L_X2Y26_SLICE_X0Y26_CIN;
  wire [0:0] CLBLL_L_X2Y26_SLICE_X0Y26_CMUX;
  wire [0:0] CLBLL_L_X2Y26_SLICE_X0Y26_CO5;
  wire [0:0] CLBLL_L_X2Y26_SLICE_X0Y26_CO6;
  wire [0:0] CLBLL_L_X2Y26_SLICE_X0Y26_COUT;
  wire [0:0] CLBLL_L_X2Y26_SLICE_X0Y26_CX;
  wire [0:0] CLBLL_L_X2Y26_SLICE_X0Y26_C_CY;
  wire [0:0] CLBLL_L_X2Y26_SLICE_X0Y26_C_XOR;
  wire [0:0] CLBLL_L_X2Y26_SLICE_X0Y26_D;
  wire [0:0] CLBLL_L_X2Y26_SLICE_X0Y26_D1;
  wire [0:0] CLBLL_L_X2Y26_SLICE_X0Y26_D2;
  wire [0:0] CLBLL_L_X2Y26_SLICE_X0Y26_D3;
  wire [0:0] CLBLL_L_X2Y26_SLICE_X0Y26_D4;
  wire [0:0] CLBLL_L_X2Y26_SLICE_X0Y26_D5;
  wire [0:0] CLBLL_L_X2Y26_SLICE_X0Y26_D6;
  wire [0:0] CLBLL_L_X2Y26_SLICE_X0Y26_DMUX;
  wire [0:0] CLBLL_L_X2Y26_SLICE_X0Y26_DO5;
  wire [0:0] CLBLL_L_X2Y26_SLICE_X0Y26_DO6;
  wire [0:0] CLBLL_L_X2Y26_SLICE_X0Y26_DX;
  wire [0:0] CLBLL_L_X2Y26_SLICE_X0Y26_D_CY;
  wire [0:0] CLBLL_L_X2Y26_SLICE_X0Y26_D_XOR;
  wire [0:0] CLBLL_L_X2Y26_SLICE_X1Y26_A;
  wire [0:0] CLBLL_L_X2Y26_SLICE_X1Y26_A1;
  wire [0:0] CLBLL_L_X2Y26_SLICE_X1Y26_A2;
  wire [0:0] CLBLL_L_X2Y26_SLICE_X1Y26_A3;
  wire [0:0] CLBLL_L_X2Y26_SLICE_X1Y26_A4;
  wire [0:0] CLBLL_L_X2Y26_SLICE_X1Y26_A5;
  wire [0:0] CLBLL_L_X2Y26_SLICE_X1Y26_A6;
  wire [0:0] CLBLL_L_X2Y26_SLICE_X1Y26_AO5;
  wire [0:0] CLBLL_L_X2Y26_SLICE_X1Y26_AO6;
  wire [0:0] CLBLL_L_X2Y26_SLICE_X1Y26_A_CY;
  wire [0:0] CLBLL_L_X2Y26_SLICE_X1Y26_A_XOR;
  wire [0:0] CLBLL_L_X2Y26_SLICE_X1Y26_B;
  wire [0:0] CLBLL_L_X2Y26_SLICE_X1Y26_B1;
  wire [0:0] CLBLL_L_X2Y26_SLICE_X1Y26_B2;
  wire [0:0] CLBLL_L_X2Y26_SLICE_X1Y26_B3;
  wire [0:0] CLBLL_L_X2Y26_SLICE_X1Y26_B4;
  wire [0:0] CLBLL_L_X2Y26_SLICE_X1Y26_B5;
  wire [0:0] CLBLL_L_X2Y26_SLICE_X1Y26_B6;
  wire [0:0] CLBLL_L_X2Y26_SLICE_X1Y26_BO5;
  wire [0:0] CLBLL_L_X2Y26_SLICE_X1Y26_BO6;
  wire [0:0] CLBLL_L_X2Y26_SLICE_X1Y26_B_CY;
  wire [0:0] CLBLL_L_X2Y26_SLICE_X1Y26_B_XOR;
  wire [0:0] CLBLL_L_X2Y26_SLICE_X1Y26_C;
  wire [0:0] CLBLL_L_X2Y26_SLICE_X1Y26_C1;
  wire [0:0] CLBLL_L_X2Y26_SLICE_X1Y26_C2;
  wire [0:0] CLBLL_L_X2Y26_SLICE_X1Y26_C3;
  wire [0:0] CLBLL_L_X2Y26_SLICE_X1Y26_C4;
  wire [0:0] CLBLL_L_X2Y26_SLICE_X1Y26_C5;
  wire [0:0] CLBLL_L_X2Y26_SLICE_X1Y26_C6;
  wire [0:0] CLBLL_L_X2Y26_SLICE_X1Y26_CO5;
  wire [0:0] CLBLL_L_X2Y26_SLICE_X1Y26_CO6;
  wire [0:0] CLBLL_L_X2Y26_SLICE_X1Y26_C_CY;
  wire [0:0] CLBLL_L_X2Y26_SLICE_X1Y26_C_XOR;
  wire [0:0] CLBLL_L_X2Y26_SLICE_X1Y26_D;
  wire [0:0] CLBLL_L_X2Y26_SLICE_X1Y26_D1;
  wire [0:0] CLBLL_L_X2Y26_SLICE_X1Y26_D2;
  wire [0:0] CLBLL_L_X2Y26_SLICE_X1Y26_D3;
  wire [0:0] CLBLL_L_X2Y26_SLICE_X1Y26_D4;
  wire [0:0] CLBLL_L_X2Y26_SLICE_X1Y26_D5;
  wire [0:0] CLBLL_L_X2Y26_SLICE_X1Y26_D6;
  wire [0:0] CLBLL_L_X2Y26_SLICE_X1Y26_DO5;
  wire [0:0] CLBLL_L_X2Y26_SLICE_X1Y26_DO6;
  wire [0:0] CLBLL_L_X2Y26_SLICE_X1Y26_D_CY;
  wire [0:0] CLBLL_L_X2Y26_SLICE_X1Y26_D_XOR;
  wire [0:0] LIOB33_SING_X0Y0_IOB_X0Y0_I;
  wire [0:0] LIOB33_X0Y11_IOB_X0Y11_I;
  wire [0:0] LIOB33_X0Y11_IOB_X0Y12_I;
  wire [0:0] LIOB33_X0Y13_IOB_X0Y13_I;
  wire [0:0] LIOB33_X0Y13_IOB_X0Y14_I;
  wire [0:0] LIOB33_X0Y15_IOB_X0Y15_I;
  wire [0:0] LIOB33_X0Y15_IOB_X0Y16_I;
  wire [0:0] LIOB33_X0Y17_IOB_X0Y17_I;
  wire [0:0] LIOB33_X0Y17_IOB_X0Y18_I;
  wire [0:0] LIOB33_X0Y19_IOB_X0Y19_I;
  wire [0:0] LIOB33_X0Y19_IOB_X0Y20_I;
  wire [0:0] LIOB33_X0Y1_IOB_X0Y1_I;
  wire [0:0] LIOB33_X0Y1_IOB_X0Y2_I;
  wire [0:0] LIOB33_X0Y21_IOB_X0Y21_I;
  wire [0:0] LIOB33_X0Y21_IOB_X0Y22_I;
  wire [0:0] LIOB33_X0Y23_IOB_X0Y23_I;
  wire [0:0] LIOB33_X0Y23_IOB_X0Y24_I;
  wire [0:0] LIOB33_X0Y25_IOB_X0Y25_I;
  wire [0:0] LIOB33_X0Y25_IOB_X0Y26_I;
  wire [0:0] LIOB33_X0Y27_IOB_X0Y27_I;
  wire [0:0] LIOB33_X0Y27_IOB_X0Y28_I;
  wire [0:0] LIOB33_X0Y29_IOB_X0Y29_I;
  wire [0:0] LIOB33_X0Y29_IOB_X0Y30_I;
  wire [0:0] LIOB33_X0Y31_IOB_X0Y31_I;
  wire [0:0] LIOB33_X0Y31_IOB_X0Y32_O;
  wire [0:0] LIOB33_X0Y33_IOB_X0Y33_O;
  wire [0:0] LIOB33_X0Y33_IOB_X0Y34_O;
  wire [0:0] LIOB33_X0Y35_IOB_X0Y35_O;
  wire [0:0] LIOB33_X0Y35_IOB_X0Y36_O;
  wire [0:0] LIOB33_X0Y37_IOB_X0Y37_O;
  wire [0:0] LIOB33_X0Y37_IOB_X0Y38_O;
  wire [0:0] LIOB33_X0Y39_IOB_X0Y39_O;
  wire [0:0] LIOB33_X0Y39_IOB_X0Y40_O;
  wire [0:0] LIOB33_X0Y3_IOB_X0Y3_I;
  wire [0:0] LIOB33_X0Y3_IOB_X0Y4_I;
  wire [0:0] LIOB33_X0Y41_IOB_X0Y41_O;
  wire [0:0] LIOB33_X0Y41_IOB_X0Y42_O;
  wire [0:0] LIOB33_X0Y43_IOB_X0Y43_O;
  wire [0:0] LIOB33_X0Y43_IOB_X0Y44_O;
  wire [0:0] LIOB33_X0Y45_IOB_X0Y45_O;
  wire [0:0] LIOB33_X0Y45_IOB_X0Y46_O;
  wire [0:0] LIOB33_X0Y47_IOB_X0Y47_O;
  wire [0:0] LIOB33_X0Y5_IOB_X0Y5_I;
  wire [0:0] LIOB33_X0Y5_IOB_X0Y6_I;
  wire [0:0] LIOB33_X0Y7_IOB_X0Y7_I;
  wire [0:0] LIOB33_X0Y7_IOB_X0Y8_I;
  wire [0:0] LIOB33_X0Y9_IOB_X0Y10_I;
  wire [0:0] LIOB33_X0Y9_IOB_X0Y9_I;
  wire [0:0] LIOI3_SING_X0Y0_ILOGIC_X0Y0_D;
  wire [0:0] LIOI3_SING_X0Y0_ILOGIC_X0Y0_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y19_ILOGIC_X0Y19_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y19_ILOGIC_X0Y19_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y19_ILOGIC_X0Y20_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y19_ILOGIC_X0Y20_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y31_ILOGIC_X0Y31_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y31_ILOGIC_X0Y31_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y31_OLOGIC_X0Y32_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y31_OLOGIC_X0Y32_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y31_OLOGIC_X0Y32_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y31_OLOGIC_X0Y32_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y43_OLOGIC_X0Y43_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y43_OLOGIC_X0Y43_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y43_OLOGIC_X0Y43_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y43_OLOGIC_X0Y43_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y43_OLOGIC_X0Y44_D1;
  wire [0:0] LIOI3_TBYTESRC_X0Y43_OLOGIC_X0Y44_OQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y43_OLOGIC_X0Y44_T1;
  wire [0:0] LIOI3_TBYTESRC_X0Y43_OLOGIC_X0Y44_TQ;
  wire [0:0] LIOI3_TBYTESRC_X0Y7_ILOGIC_X0Y7_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y7_ILOGIC_X0Y7_O;
  wire [0:0] LIOI3_TBYTESRC_X0Y7_ILOGIC_X0Y8_D;
  wire [0:0] LIOI3_TBYTESRC_X0Y7_ILOGIC_X0Y8_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y13_ILOGIC_X0Y13_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y13_ILOGIC_X0Y13_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y13_ILOGIC_X0Y14_D;
  wire [0:0] LIOI3_TBYTETERM_X0Y13_ILOGIC_X0Y14_O;
  wire [0:0] LIOI3_TBYTETERM_X0Y37_OLOGIC_X0Y37_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y37_OLOGIC_X0Y37_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y37_OLOGIC_X0Y37_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y37_OLOGIC_X0Y37_TQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y37_OLOGIC_X0Y38_D1;
  wire [0:0] LIOI3_TBYTETERM_X0Y37_OLOGIC_X0Y38_OQ;
  wire [0:0] LIOI3_TBYTETERM_X0Y37_OLOGIC_X0Y38_T1;
  wire [0:0] LIOI3_TBYTETERM_X0Y37_OLOGIC_X0Y38_TQ;
  wire [0:0] LIOI3_X0Y11_ILOGIC_X0Y11_D;
  wire [0:0] LIOI3_X0Y11_ILOGIC_X0Y11_O;
  wire [0:0] LIOI3_X0Y11_ILOGIC_X0Y12_D;
  wire [0:0] LIOI3_X0Y11_ILOGIC_X0Y12_O;
  wire [0:0] LIOI3_X0Y15_ILOGIC_X0Y15_D;
  wire [0:0] LIOI3_X0Y15_ILOGIC_X0Y15_O;
  wire [0:0] LIOI3_X0Y15_ILOGIC_X0Y16_D;
  wire [0:0] LIOI3_X0Y15_ILOGIC_X0Y16_O;
  wire [0:0] LIOI3_X0Y17_ILOGIC_X0Y17_D;
  wire [0:0] LIOI3_X0Y17_ILOGIC_X0Y17_O;
  wire [0:0] LIOI3_X0Y17_ILOGIC_X0Y18_D;
  wire [0:0] LIOI3_X0Y17_ILOGIC_X0Y18_O;
  wire [0:0] LIOI3_X0Y1_ILOGIC_X0Y1_D;
  wire [0:0] LIOI3_X0Y1_ILOGIC_X0Y1_O;
  wire [0:0] LIOI3_X0Y1_ILOGIC_X0Y2_D;
  wire [0:0] LIOI3_X0Y1_ILOGIC_X0Y2_O;
  wire [0:0] LIOI3_X0Y21_ILOGIC_X0Y21_D;
  wire [0:0] LIOI3_X0Y21_ILOGIC_X0Y21_O;
  wire [0:0] LIOI3_X0Y21_ILOGIC_X0Y22_D;
  wire [0:0] LIOI3_X0Y21_ILOGIC_X0Y22_O;
  wire [0:0] LIOI3_X0Y23_ILOGIC_X0Y23_D;
  wire [0:0] LIOI3_X0Y23_ILOGIC_X0Y23_O;
  wire [0:0] LIOI3_X0Y23_ILOGIC_X0Y24_D;
  wire [0:0] LIOI3_X0Y23_ILOGIC_X0Y24_O;
  wire [0:0] LIOI3_X0Y25_ILOGIC_X0Y25_D;
  wire [0:0] LIOI3_X0Y25_ILOGIC_X0Y25_O;
  wire [0:0] LIOI3_X0Y25_ILOGIC_X0Y26_D;
  wire [0:0] LIOI3_X0Y25_ILOGIC_X0Y26_O;
  wire [0:0] LIOI3_X0Y27_ILOGIC_X0Y27_D;
  wire [0:0] LIOI3_X0Y27_ILOGIC_X0Y27_O;
  wire [0:0] LIOI3_X0Y27_ILOGIC_X0Y28_D;
  wire [0:0] LIOI3_X0Y27_ILOGIC_X0Y28_O;
  wire [0:0] LIOI3_X0Y29_ILOGIC_X0Y29_D;
  wire [0:0] LIOI3_X0Y29_ILOGIC_X0Y29_O;
  wire [0:0] LIOI3_X0Y29_ILOGIC_X0Y30_D;
  wire [0:0] LIOI3_X0Y29_ILOGIC_X0Y30_O;
  wire [0:0] LIOI3_X0Y33_OLOGIC_X0Y33_D1;
  wire [0:0] LIOI3_X0Y33_OLOGIC_X0Y33_OQ;
  wire [0:0] LIOI3_X0Y33_OLOGIC_X0Y33_T1;
  wire [0:0] LIOI3_X0Y33_OLOGIC_X0Y33_TQ;
  wire [0:0] LIOI3_X0Y33_OLOGIC_X0Y34_D1;
  wire [0:0] LIOI3_X0Y33_OLOGIC_X0Y34_OQ;
  wire [0:0] LIOI3_X0Y33_OLOGIC_X0Y34_T1;
  wire [0:0] LIOI3_X0Y33_OLOGIC_X0Y34_TQ;
  wire [0:0] LIOI3_X0Y35_OLOGIC_X0Y35_D1;
  wire [0:0] LIOI3_X0Y35_OLOGIC_X0Y35_OQ;
  wire [0:0] LIOI3_X0Y35_OLOGIC_X0Y35_T1;
  wire [0:0] LIOI3_X0Y35_OLOGIC_X0Y35_TQ;
  wire [0:0] LIOI3_X0Y35_OLOGIC_X0Y36_D1;
  wire [0:0] LIOI3_X0Y35_OLOGIC_X0Y36_OQ;
  wire [0:0] LIOI3_X0Y35_OLOGIC_X0Y36_T1;
  wire [0:0] LIOI3_X0Y35_OLOGIC_X0Y36_TQ;
  wire [0:0] LIOI3_X0Y39_OLOGIC_X0Y39_D1;
  wire [0:0] LIOI3_X0Y39_OLOGIC_X0Y39_OQ;
  wire [0:0] LIOI3_X0Y39_OLOGIC_X0Y39_T1;
  wire [0:0] LIOI3_X0Y39_OLOGIC_X0Y39_TQ;
  wire [0:0] LIOI3_X0Y39_OLOGIC_X0Y40_D1;
  wire [0:0] LIOI3_X0Y39_OLOGIC_X0Y40_OQ;
  wire [0:0] LIOI3_X0Y39_OLOGIC_X0Y40_T1;
  wire [0:0] LIOI3_X0Y39_OLOGIC_X0Y40_TQ;
  wire [0:0] LIOI3_X0Y3_ILOGIC_X0Y3_D;
  wire [0:0] LIOI3_X0Y3_ILOGIC_X0Y3_O;
  wire [0:0] LIOI3_X0Y3_ILOGIC_X0Y4_D;
  wire [0:0] LIOI3_X0Y3_ILOGIC_X0Y4_O;
  wire [0:0] LIOI3_X0Y41_OLOGIC_X0Y41_D1;
  wire [0:0] LIOI3_X0Y41_OLOGIC_X0Y41_OQ;
  wire [0:0] LIOI3_X0Y41_OLOGIC_X0Y41_T1;
  wire [0:0] LIOI3_X0Y41_OLOGIC_X0Y41_TQ;
  wire [0:0] LIOI3_X0Y41_OLOGIC_X0Y42_D1;
  wire [0:0] LIOI3_X0Y41_OLOGIC_X0Y42_OQ;
  wire [0:0] LIOI3_X0Y41_OLOGIC_X0Y42_T1;
  wire [0:0] LIOI3_X0Y41_OLOGIC_X0Y42_TQ;
  wire [0:0] LIOI3_X0Y45_OLOGIC_X0Y45_D1;
  wire [0:0] LIOI3_X0Y45_OLOGIC_X0Y45_OQ;
  wire [0:0] LIOI3_X0Y45_OLOGIC_X0Y45_T1;
  wire [0:0] LIOI3_X0Y45_OLOGIC_X0Y45_TQ;
  wire [0:0] LIOI3_X0Y45_OLOGIC_X0Y46_D1;
  wire [0:0] LIOI3_X0Y45_OLOGIC_X0Y46_OQ;
  wire [0:0] LIOI3_X0Y45_OLOGIC_X0Y46_T1;
  wire [0:0] LIOI3_X0Y45_OLOGIC_X0Y46_TQ;
  wire [0:0] LIOI3_X0Y47_OLOGIC_X0Y47_D1;
  wire [0:0] LIOI3_X0Y47_OLOGIC_X0Y47_OQ;
  wire [0:0] LIOI3_X0Y47_OLOGIC_X0Y47_T1;
  wire [0:0] LIOI3_X0Y47_OLOGIC_X0Y47_TQ;
  wire [0:0] LIOI3_X0Y5_ILOGIC_X0Y5_D;
  wire [0:0] LIOI3_X0Y5_ILOGIC_X0Y5_O;
  wire [0:0] LIOI3_X0Y5_ILOGIC_X0Y6_D;
  wire [0:0] LIOI3_X0Y5_ILOGIC_X0Y6_O;
  wire [0:0] LIOI3_X0Y9_ILOGIC_X0Y10_D;
  wire [0:0] LIOI3_X0Y9_ILOGIC_X0Y10_O;
  wire [0:0] LIOI3_X0Y9_ILOGIC_X0Y9_D;
  wire [0:0] LIOI3_X0Y9_ILOGIC_X0Y9_O;
  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLL_L_X2Y23_SLICE_X0Y23_CARRY4 (
.CI(1'b0),
.CO({CLBLL_L_X2Y23_SLICE_X0Y23_D_CY, CLBLL_L_X2Y23_SLICE_X0Y23_C_CY, CLBLL_L_X2Y23_SLICE_X0Y23_B_CY, CLBLL_L_X2Y23_SLICE_X0Y23_A_CY}),
.CYINIT(1'b0),
.DI({LIOB33_X0Y3_IOB_X0Y3_I, LIOB33_X0Y1_IOB_X0Y2_I, LIOB33_X0Y1_IOB_X0Y1_I, LIOB33_SING_X0Y0_IOB_X0Y0_I}),
.O({CLBLL_L_X2Y23_SLICE_X0Y23_D_XOR, CLBLL_L_X2Y23_SLICE_X0Y23_C_XOR, CLBLL_L_X2Y23_SLICE_X0Y23_B_XOR, CLBLL_L_X2Y23_SLICE_X0Y23_A_XOR}),
.S({CLBLL_L_X2Y23_SLICE_X0Y23_DO6, CLBLL_L_X2Y23_SLICE_X0Y23_CO6, CLBLL_L_X2Y23_SLICE_X0Y23_BO6, CLBLL_L_X2Y23_SLICE_X0Y23_AO6})
  );
  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6666666666666666)
  ) CLBLL_L_X2Y23_SLICE_X0Y23_DLUT (
.I0(LIOB33_X0Y3_IOB_X0Y3_I),
.I1(LIOB33_X0Y19_IOB_X0Y19_I),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y23_SLICE_X0Y23_DO5),
.O6(CLBLL_L_X2Y23_SLICE_X0Y23_DO6)
  );
  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5a5a5a5a5a5a5a5a)
  ) CLBLL_L_X2Y23_SLICE_X0Y23_CLUT (
.I0(LIOB33_X0Y17_IOB_X0Y18_I),
.I1(1'b1),
.I2(LIOB33_X0Y1_IOB_X0Y2_I),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y23_SLICE_X0Y23_CO5),
.O6(CLBLL_L_X2Y23_SLICE_X0Y23_CO6)
  );
  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5a5a5a5a5a5a5a5a)
  ) CLBLL_L_X2Y23_SLICE_X0Y23_BLUT (
.I0(LIOB33_X0Y1_IOB_X0Y1_I),
.I1(1'b1),
.I2(LIOB33_X0Y17_IOB_X0Y17_I),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y23_SLICE_X0Y23_BO5),
.O6(CLBLL_L_X2Y23_SLICE_X0Y23_BO6)
  );
  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5555aaaa5555aaaa)
  ) CLBLL_L_X2Y23_SLICE_X0Y23_ALUT (
.I0(LIOB33_SING_X0Y0_IOB_X0Y0_I),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(LIOB33_X0Y15_IOB_X0Y16_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y23_SLICE_X0Y23_AO5),
.O6(CLBLL_L_X2Y23_SLICE_X0Y23_AO6)
  );
  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y23_SLICE_X1Y23_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y23_SLICE_X1Y23_DO5),
.O6(CLBLL_L_X2Y23_SLICE_X1Y23_DO6)
  );
  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y23_SLICE_X1Y23_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y23_SLICE_X1Y23_CO5),
.O6(CLBLL_L_X2Y23_SLICE_X1Y23_CO6)
  );
  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y23_SLICE_X1Y23_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y23_SLICE_X1Y23_BO5),
.O6(CLBLL_L_X2Y23_SLICE_X1Y23_BO6)
  );
  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y23_SLICE_X1Y23_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y23_SLICE_X1Y23_AO5),
.O6(CLBLL_L_X2Y23_SLICE_X1Y23_AO6)
  );
  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLL_L_X2Y24_SLICE_X0Y24_CARRY4 (
.CI(CLBLL_L_X2Y23_SLICE_X0Y23_D_CY),
.CO({CLBLL_L_X2Y24_SLICE_X0Y24_D_CY, CLBLL_L_X2Y24_SLICE_X0Y24_C_CY, CLBLL_L_X2Y24_SLICE_X0Y24_B_CY, CLBLL_L_X2Y24_SLICE_X0Y24_A_CY}),
.CYINIT(1'b0),
.DI({LIOB33_X0Y7_IOB_X0Y7_I, LIOB33_X0Y5_IOB_X0Y6_I, LIOB33_X0Y5_IOB_X0Y5_I, LIOB33_X0Y3_IOB_X0Y4_I}),
.O({CLBLL_L_X2Y24_SLICE_X0Y24_D_XOR, CLBLL_L_X2Y24_SLICE_X0Y24_C_XOR, CLBLL_L_X2Y24_SLICE_X0Y24_B_XOR, CLBLL_L_X2Y24_SLICE_X0Y24_A_XOR}),
.S({CLBLL_L_X2Y24_SLICE_X0Y24_DO6, CLBLL_L_X2Y24_SLICE_X0Y24_CO6, CLBLL_L_X2Y24_SLICE_X0Y24_BO6, CLBLL_L_X2Y24_SLICE_X0Y24_AO6})
  );
  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h6666666666666666)
  ) CLBLL_L_X2Y24_SLICE_X0Y24_DLUT (
.I0(LIOB33_X0Y23_IOB_X0Y23_I),
.I1(LIOB33_X0Y7_IOB_X0Y7_I),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y24_SLICE_X0Y24_DO5),
.O6(CLBLL_L_X2Y24_SLICE_X0Y24_DO6)
  );
  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h5a5a5a5a5a5a5a5a)
  ) CLBLL_L_X2Y24_SLICE_X0Y24_CLUT (
.I0(LIOB33_X0Y21_IOB_X0Y22_I),
.I1(1'b1),
.I2(LIOB33_X0Y5_IOB_X0Y6_I),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y24_SLICE_X0Y24_CO5),
.O6(CLBLL_L_X2Y24_SLICE_X0Y24_CO6)
  );
  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5a5a5a5a5a5a5a5a)
  ) CLBLL_L_X2Y24_SLICE_X0Y24_BLUT (
.I0(LIOB33_X0Y5_IOB_X0Y5_I),
.I1(1'b1),
.I2(LIOB33_X0Y21_IOB_X0Y21_I),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y24_SLICE_X0Y24_BO5),
.O6(CLBLL_L_X2Y24_SLICE_X0Y24_BO6)
  );
  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h00ffff0000ffff00)
  ) CLBLL_L_X2Y24_SLICE_X0Y24_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(LIOB33_X0Y3_IOB_X0Y4_I),
.I4(LIOB33_X0Y19_IOB_X0Y20_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y24_SLICE_X0Y24_AO5),
.O6(CLBLL_L_X2Y24_SLICE_X0Y24_AO6)
  );
  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y24_SLICE_X1Y24_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y24_SLICE_X1Y24_DO5),
.O6(CLBLL_L_X2Y24_SLICE_X1Y24_DO6)
  );
  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y24_SLICE_X1Y24_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y24_SLICE_X1Y24_CO5),
.O6(CLBLL_L_X2Y24_SLICE_X1Y24_CO6)
  );
  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y24_SLICE_X1Y24_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y24_SLICE_X1Y24_BO5),
.O6(CLBLL_L_X2Y24_SLICE_X1Y24_BO6)
  );
  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y24_SLICE_X1Y24_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y24_SLICE_X1Y24_AO5),
.O6(CLBLL_L_X2Y24_SLICE_X1Y24_AO6)
  );
  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLL_L_X2Y25_SLICE_X0Y25_CARRY4 (
.CI(CLBLL_L_X2Y24_SLICE_X0Y24_D_CY),
.CO({CLBLL_L_X2Y25_SLICE_X0Y25_D_CY, CLBLL_L_X2Y25_SLICE_X0Y25_C_CY, CLBLL_L_X2Y25_SLICE_X0Y25_B_CY, CLBLL_L_X2Y25_SLICE_X0Y25_A_CY}),
.CYINIT(1'b0),
.DI({LIOB33_X0Y11_IOB_X0Y11_I, LIOB33_X0Y9_IOB_X0Y10_I, LIOB33_X0Y9_IOB_X0Y9_I, LIOB33_X0Y7_IOB_X0Y8_I}),
.O({CLBLL_L_X2Y25_SLICE_X0Y25_D_XOR, CLBLL_L_X2Y25_SLICE_X0Y25_C_XOR, CLBLL_L_X2Y25_SLICE_X0Y25_B_XOR, CLBLL_L_X2Y25_SLICE_X0Y25_A_XOR}),
.S({CLBLL_L_X2Y25_SLICE_X0Y25_DO6, CLBLL_L_X2Y25_SLICE_X0Y25_CO6, CLBLL_L_X2Y25_SLICE_X0Y25_BO6, CLBLL_L_X2Y25_SLICE_X0Y25_AO6})
  );
  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5a5a5a5a5a5a5a5a)
  ) CLBLL_L_X2Y25_SLICE_X0Y25_DLUT (
.I0(LIOB33_X0Y11_IOB_X0Y11_I),
.I1(1'b1),
.I2(LIOB33_X0Y27_IOB_X0Y27_I),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y25_SLICE_X0Y25_DO5),
.O6(CLBLL_L_X2Y25_SLICE_X0Y25_DO6)
  );
  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h55555555aaaaaaaa)
  ) CLBLL_L_X2Y25_SLICE_X0Y25_CLUT (
.I0(LIOB33_X0Y9_IOB_X0Y10_I),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(LIOB33_X0Y25_IOB_X0Y26_I),
.O5(CLBLL_L_X2Y25_SLICE_X0Y25_CO5),
.O6(CLBLL_L_X2Y25_SLICE_X0Y25_CO6)
  );
  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h5a5a5a5a5a5a5a5a)
  ) CLBLL_L_X2Y25_SLICE_X0Y25_BLUT (
.I0(LIOB33_X0Y9_IOB_X0Y9_I),
.I1(1'b1),
.I2(LIOB33_X0Y25_IOB_X0Y25_I),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y25_SLICE_X0Y25_BO5),
.O6(CLBLL_L_X2Y25_SLICE_X0Y25_BO6)
  );
  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0f0ff0f00f0ff0f0)
  ) CLBLL_L_X2Y25_SLICE_X0Y25_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(LIOB33_X0Y23_IOB_X0Y24_I),
.I3(1'b1),
.I4(LIOB33_X0Y7_IOB_X0Y8_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y25_SLICE_X0Y25_AO5),
.O6(CLBLL_L_X2Y25_SLICE_X0Y25_AO6)
  );
  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y25_SLICE_X1Y25_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y25_SLICE_X1Y25_DO5),
.O6(CLBLL_L_X2Y25_SLICE_X1Y25_DO6)
  );
  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y25_SLICE_X1Y25_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y25_SLICE_X1Y25_CO5),
.O6(CLBLL_L_X2Y25_SLICE_X1Y25_CO6)
  );
  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y25_SLICE_X1Y25_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y25_SLICE_X1Y25_BO5),
.O6(CLBLL_L_X2Y25_SLICE_X1Y25_BO6)
  );
  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y25_SLICE_X1Y25_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y25_SLICE_X1Y25_AO5),
.O6(CLBLL_L_X2Y25_SLICE_X1Y25_AO6)
  );
  (* KEEP, DONT_TOUCH, BEL = "CARRY4" *)
  CARRY4 #(
  ) CLBLL_L_X2Y26_SLICE_X0Y26_CARRY4 (
.CI(CLBLL_L_X2Y25_SLICE_X0Y25_D_CY),
.CO({CLBLL_L_X2Y26_SLICE_X0Y26_D_CY, CLBLL_L_X2Y26_SLICE_X0Y26_C_CY, CLBLL_L_X2Y26_SLICE_X0Y26_B_CY, CLBLL_L_X2Y26_SLICE_X0Y26_A_CY}),
.CYINIT(1'b0),
.DI({1'b0, LIOB33_X0Y13_IOB_X0Y14_I, LIOB33_X0Y13_IOB_X0Y13_I, LIOB33_X0Y11_IOB_X0Y12_I}),
.O({CLBLL_L_X2Y26_SLICE_X0Y26_D_XOR, CLBLL_L_X2Y26_SLICE_X0Y26_C_XOR, CLBLL_L_X2Y26_SLICE_X0Y26_B_XOR, CLBLL_L_X2Y26_SLICE_X0Y26_A_XOR}),
.S({CLBLL_L_X2Y26_SLICE_X0Y26_DO6, CLBLL_L_X2Y26_SLICE_X0Y26_CO6, CLBLL_L_X2Y26_SLICE_X0Y26_BO6, CLBLL_L_X2Y26_SLICE_X0Y26_AO6})
  );
  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h5a5a5a5a5a5a5a5a)
  ) CLBLL_L_X2Y26_SLICE_X0Y26_DLUT (
.I0(LIOB33_X0Y15_IOB_X0Y15_I),
.I1(1'b1),
.I2(LIOB33_X0Y31_IOB_X0Y31_I),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y26_SLICE_X0Y26_DO5),
.O6(CLBLL_L_X2Y26_SLICE_X0Y26_DO6)
  );
  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h55555555aaaaaaaa)
  ) CLBLL_L_X2Y26_SLICE_X0Y26_CLUT (
.I0(LIOB33_X0Y13_IOB_X0Y14_I),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(LIOB33_X0Y29_IOB_X0Y30_I),
.O5(CLBLL_L_X2Y26_SLICE_X0Y26_CO5),
.O6(CLBLL_L_X2Y26_SLICE_X0Y26_CO6)
  );
  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h3333cccc3333cccc)
  ) CLBLL_L_X2Y26_SLICE_X0Y26_BLUT (
.I0(1'b1),
.I1(LIOB33_X0Y13_IOB_X0Y13_I),
.I2(1'b1),
.I3(1'b1),
.I4(LIOB33_X0Y29_IOB_X0Y29_I),
.I5(1'b1),
.O5(CLBLL_L_X2Y26_SLICE_X0Y26_BO5),
.O6(CLBLL_L_X2Y26_SLICE_X0Y26_BO6)
  );
  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h5a5a5a5a5a5a5a5a)
  ) CLBLL_L_X2Y26_SLICE_X0Y26_ALUT (
.I0(LIOB33_X0Y27_IOB_X0Y28_I),
.I1(1'b1),
.I2(LIOB33_X0Y11_IOB_X0Y12_I),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y26_SLICE_X0Y26_AO5),
.O6(CLBLL_L_X2Y26_SLICE_X0Y26_AO6)
  );
  (* KEEP, DONT_TOUCH, BEL = "D6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y26_SLICE_X1Y26_DLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y26_SLICE_X1Y26_DO5),
.O6(CLBLL_L_X2Y26_SLICE_X1Y26_DO6)
  );
  (* KEEP, DONT_TOUCH, BEL = "C6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y26_SLICE_X1Y26_CLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y26_SLICE_X1Y26_CO5),
.O6(CLBLL_L_X2Y26_SLICE_X1Y26_CO6)
  );
  (* KEEP, DONT_TOUCH, BEL = "B6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y26_SLICE_X1Y26_BLUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y26_SLICE_X1Y26_BO5),
.O6(CLBLL_L_X2Y26_SLICE_X1Y26_BO6)
  );
  (* KEEP, DONT_TOUCH, BEL = "A6LUT" *)
  LUT6_2 #(
    .INIT(64'h0000000000000000)
  ) CLBLL_L_X2Y26_SLICE_X1Y26_ALUT (
.I0(1'b1),
.I1(1'b1),
.I2(1'b1),
.I3(1'b1),
.I4(1'b1),
.I5(1'b1),
.O5(CLBLL_L_X2Y26_SLICE_X1Y26_AO5),
.O6(CLBLL_L_X2Y26_SLICE_X1Y26_AO6)
  );
  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y1_IOB_X0Y1_IBUF (
.I(a[1]),
.O(LIOB33_X0Y1_IOB_X0Y1_I)
  );
  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y1_IOB_X0Y2_IBUF (
.I(a[2]),
.O(LIOB33_X0Y1_IOB_X0Y2_I)
  );
  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y3_IOB_X0Y3_IBUF (
.I(a[3]),
.O(LIOB33_X0Y3_IOB_X0Y3_I)
  );
  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y3_IOB_X0Y4_IBUF (
.I(a[4]),
.O(LIOB33_X0Y3_IOB_X0Y4_I)
  );
  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y5_IOB_X0Y5_IBUF (
.I(a[5]),
.O(LIOB33_X0Y5_IOB_X0Y5_I)
  );
  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y5_IOB_X0Y6_IBUF (
.I(a[6]),
.O(LIOB33_X0Y5_IOB_X0Y6_I)
  );
  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y7_IOB_X0Y7_IBUF (
.I(a[7]),
.O(LIOB33_X0Y7_IOB_X0Y7_I)
  );
  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y7_IOB_X0Y8_IBUF (
.I(a[8]),
.O(LIOB33_X0Y7_IOB_X0Y8_I)
  );
  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y9_IOB_X0Y9_IBUF (
.I(a[9]),
.O(LIOB33_X0Y9_IOB_X0Y9_I)
  );
  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y9_IOB_X0Y10_IBUF (
.I(a[10]),
.O(LIOB33_X0Y9_IOB_X0Y10_I)
  );
  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y11_IOB_X0Y11_IBUF (
.I(a[11]),
.O(LIOB33_X0Y11_IOB_X0Y11_I)
  );
  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y11_IOB_X0Y12_IBUF (
.I(a[12]),
.O(LIOB33_X0Y11_IOB_X0Y12_I)
  );
  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y13_IOB_X0Y13_IBUF (
.I(a[13]),
.O(LIOB33_X0Y13_IOB_X0Y13_I)
  );
  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y13_IOB_X0Y14_IBUF (
.I(a[14]),
.O(LIOB33_X0Y13_IOB_X0Y14_I)
  );
  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y15_IOB_X0Y15_IBUF (
.I(a[15]),
.O(LIOB33_X0Y15_IOB_X0Y15_I)
  );
  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y15_IOB_X0Y16_IBUF (
.I(b[0]),
.O(LIOB33_X0Y15_IOB_X0Y16_I)
  );
  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y17_IOB_X0Y17_IBUF (
.I(b[1]),
.O(LIOB33_X0Y17_IOB_X0Y17_I)
  );
  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y17_IOB_X0Y18_IBUF (
.I(b[2]),
.O(LIOB33_X0Y17_IOB_X0Y18_I)
  );
  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y19_IOB_X0Y19_IBUF (
.I(b[3]),
.O(LIOB33_X0Y19_IOB_X0Y19_I)
  );
  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y19_IOB_X0Y20_IBUF (
.I(b[4]),
.O(LIOB33_X0Y19_IOB_X0Y20_I)
  );
  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y21_IOB_X0Y21_IBUF (
.I(b[5]),
.O(LIOB33_X0Y21_IOB_X0Y21_I)
  );
  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y21_IOB_X0Y22_IBUF (
.I(b[6]),
.O(LIOB33_X0Y21_IOB_X0Y22_I)
  );
  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y23_IOB_X0Y23_IBUF (
.I(b[7]),
.O(LIOB33_X0Y23_IOB_X0Y23_I)
  );
  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y23_IOB_X0Y24_IBUF (
.I(b[8]),
.O(LIOB33_X0Y23_IOB_X0Y24_I)
  );
  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y25_IOB_X0Y25_IBUF (
.I(b[9]),
.O(LIOB33_X0Y25_IOB_X0Y25_I)
  );
  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y25_IOB_X0Y26_IBUF (
.I(b[10]),
.O(LIOB33_X0Y25_IOB_X0Y26_I)
  );
  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y27_IOB_X0Y27_IBUF (
.I(b[11]),
.O(LIOB33_X0Y27_IOB_X0Y27_I)
  );
  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y27_IOB_X0Y28_IBUF (
.I(b[12]),
.O(LIOB33_X0Y27_IOB_X0Y28_I)
  );
  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y29_IOB_X0Y29_IBUF (
.I(b[13]),
.O(LIOB33_X0Y29_IOB_X0Y29_I)
  );
  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y29_IOB_X0Y30_IBUF (
.I(b[14]),
.O(LIOB33_X0Y29_IOB_X0Y30_I)
  );
  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_X0Y31_IOB_X0Y31_IBUF (
.I(b[15]),
.O(LIOB33_X0Y31_IOB_X0Y31_I)
  );
  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_X0Y31_IOB_X0Y32_OBUF (
.I(CLBLL_L_X2Y23_SLICE_X0Y23_A_XOR),
.O(o[0])
  );
  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_X0Y33_IOB_X0Y33_OBUF (
.I(CLBLL_L_X2Y23_SLICE_X0Y23_B_XOR),
.O(o[1])
  );
  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_X0Y33_IOB_X0Y34_OBUF (
.I(CLBLL_L_X2Y23_SLICE_X0Y23_C_XOR),
.O(o[2])
  );
  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_X0Y35_IOB_X0Y35_OBUF (
.I(CLBLL_L_X2Y23_SLICE_X0Y23_D_XOR),
.O(o[3])
  );
  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_X0Y35_IOB_X0Y36_OBUF (
.I(CLBLL_L_X2Y24_SLICE_X0Y24_A_XOR),
.O(o[4])
  );
  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_X0Y37_IOB_X0Y37_OBUF (
.I(CLBLL_L_X2Y24_SLICE_X0Y24_B_XOR),
.O(o[5])
  );
  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_X0Y37_IOB_X0Y38_OBUF (
.I(CLBLL_L_X2Y24_SLICE_X0Y24_C_XOR),
.O(o[6])
  );
  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_X0Y39_IOB_X0Y39_OBUF (
.I(CLBLL_L_X2Y24_SLICE_X0Y24_D_XOR),
.O(o[7])
  );
  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_X0Y39_IOB_X0Y40_OBUF (
.I(CLBLL_L_X2Y25_SLICE_X0Y25_A_XOR),
.O(o[8])
  );
  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_X0Y41_IOB_X0Y41_OBUF (
.I(CLBLL_L_X2Y25_SLICE_X0Y25_B_XOR),
.O(o[9])
  );
  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_X0Y41_IOB_X0Y42_OBUF (
.I(CLBLL_L_X2Y25_SLICE_X0Y25_C_XOR),
.O(o[10])
  );
  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_X0Y43_IOB_X0Y43_OBUF (
.I(CLBLL_L_X2Y25_SLICE_X0Y25_D_XOR),
.O(o[11])
  );
  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_X0Y43_IOB_X0Y44_OBUF (
.I(CLBLL_L_X2Y26_SLICE_X0Y26_A_XOR),
.O(o[12])
  );
  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_X0Y45_IOB_X0Y45_OBUF (
.I(CLBLL_L_X2Y26_SLICE_X0Y26_B_XOR),
.O(o[13])
  );
  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_X0Y45_IOB_X0Y46_OBUF (
.I(CLBLL_L_X2Y26_SLICE_X0Y26_C_XOR),
.O(o[14])
  );
  (* KEEP, DONT_TOUCH, BEL = "OUTBUF" *)
  OBUF #(
    .DRIVE("12"),
    .IOSTANDARD("LVCMOS33"),
    .SLEW("SLOW")
  ) LIOB33_X0Y47_IOB_X0Y47_OBUF (
.I(CLBLL_L_X2Y26_SLICE_X0Y26_D_XOR),
.O(o[15])
  );
  (* KEEP, DONT_TOUCH, BEL = "INBUF_EN" *)
  IBUF #(
    .IOSTANDARD("LVCMOS33")
  ) LIOB33_SING_X0Y0_IOB_X0Y0_IBUF (
.I(a[0]),
.O(LIOB33_SING_X0Y0_IOB_X0Y0_I)
  );
  assign CLBLL_L_X2Y23_SLICE_X0Y23_COUT = CLBLL_L_X2Y23_SLICE_X0Y23_D_CY;
  assign CLBLL_L_X2Y23_SLICE_X0Y23_A = CLBLL_L_X2Y23_SLICE_X0Y23_AO6;
  assign CLBLL_L_X2Y23_SLICE_X0Y23_B = CLBLL_L_X2Y23_SLICE_X0Y23_BO6;
  assign CLBLL_L_X2Y23_SLICE_X0Y23_C = CLBLL_L_X2Y23_SLICE_X0Y23_CO6;
  assign CLBLL_L_X2Y23_SLICE_X0Y23_D = CLBLL_L_X2Y23_SLICE_X0Y23_DO6;
  assign CLBLL_L_X2Y23_SLICE_X0Y23_AMUX = CLBLL_L_X2Y23_SLICE_X0Y23_A_XOR;
  assign CLBLL_L_X2Y23_SLICE_X0Y23_BMUX = CLBLL_L_X2Y23_SLICE_X0Y23_B_XOR;
  assign CLBLL_L_X2Y23_SLICE_X0Y23_CMUX = CLBLL_L_X2Y23_SLICE_X0Y23_C_XOR;
  assign CLBLL_L_X2Y23_SLICE_X0Y23_DMUX = CLBLL_L_X2Y23_SLICE_X0Y23_D_XOR;
  assign CLBLL_L_X2Y23_SLICE_X1Y23_COUT = CLBLL_L_X2Y23_SLICE_X1Y23_D_CY;
  assign CLBLL_L_X2Y23_SLICE_X1Y23_A = CLBLL_L_X2Y23_SLICE_X1Y23_AO6;
  assign CLBLL_L_X2Y23_SLICE_X1Y23_B = CLBLL_L_X2Y23_SLICE_X1Y23_BO6;
  assign CLBLL_L_X2Y23_SLICE_X1Y23_C = CLBLL_L_X2Y23_SLICE_X1Y23_CO6;
  assign CLBLL_L_X2Y23_SLICE_X1Y23_D = CLBLL_L_X2Y23_SLICE_X1Y23_DO6;
  assign CLBLL_L_X2Y24_SLICE_X0Y24_COUT = CLBLL_L_X2Y24_SLICE_X0Y24_D_CY;
  assign CLBLL_L_X2Y24_SLICE_X0Y24_A = CLBLL_L_X2Y24_SLICE_X0Y24_AO6;
  assign CLBLL_L_X2Y24_SLICE_X0Y24_B = CLBLL_L_X2Y24_SLICE_X0Y24_BO6;
  assign CLBLL_L_X2Y24_SLICE_X0Y24_C = CLBLL_L_X2Y24_SLICE_X0Y24_CO6;
  assign CLBLL_L_X2Y24_SLICE_X0Y24_D = CLBLL_L_X2Y24_SLICE_X0Y24_DO6;
  assign CLBLL_L_X2Y24_SLICE_X0Y24_AMUX = CLBLL_L_X2Y24_SLICE_X0Y24_A_XOR;
  assign CLBLL_L_X2Y24_SLICE_X0Y24_BMUX = CLBLL_L_X2Y24_SLICE_X0Y24_B_XOR;
  assign CLBLL_L_X2Y24_SLICE_X0Y24_CMUX = CLBLL_L_X2Y24_SLICE_X0Y24_C_XOR;
  assign CLBLL_L_X2Y24_SLICE_X0Y24_DMUX = CLBLL_L_X2Y24_SLICE_X0Y24_D_XOR;
  assign CLBLL_L_X2Y24_SLICE_X1Y24_COUT = CLBLL_L_X2Y24_SLICE_X1Y24_D_CY;
  assign CLBLL_L_X2Y24_SLICE_X1Y24_A = CLBLL_L_X2Y24_SLICE_X1Y24_AO6;
  assign CLBLL_L_X2Y24_SLICE_X1Y24_B = CLBLL_L_X2Y24_SLICE_X1Y24_BO6;
  assign CLBLL_L_X2Y24_SLICE_X1Y24_C = CLBLL_L_X2Y24_SLICE_X1Y24_CO6;
  assign CLBLL_L_X2Y24_SLICE_X1Y24_D = CLBLL_L_X2Y24_SLICE_X1Y24_DO6;
  assign CLBLL_L_X2Y25_SLICE_X0Y25_COUT = CLBLL_L_X2Y25_SLICE_X0Y25_D_CY;
  assign CLBLL_L_X2Y25_SLICE_X0Y25_A = CLBLL_L_X2Y25_SLICE_X0Y25_AO6;
  assign CLBLL_L_X2Y25_SLICE_X0Y25_B = CLBLL_L_X2Y25_SLICE_X0Y25_BO6;
  assign CLBLL_L_X2Y25_SLICE_X0Y25_C = CLBLL_L_X2Y25_SLICE_X0Y25_CO6;
  assign CLBLL_L_X2Y25_SLICE_X0Y25_D = CLBLL_L_X2Y25_SLICE_X0Y25_DO6;
  assign CLBLL_L_X2Y25_SLICE_X0Y25_AMUX = CLBLL_L_X2Y25_SLICE_X0Y25_A_XOR;
  assign CLBLL_L_X2Y25_SLICE_X0Y25_BMUX = CLBLL_L_X2Y25_SLICE_X0Y25_B_XOR;
  assign CLBLL_L_X2Y25_SLICE_X0Y25_CMUX = CLBLL_L_X2Y25_SLICE_X0Y25_C_XOR;
  assign CLBLL_L_X2Y25_SLICE_X0Y25_DMUX = CLBLL_L_X2Y25_SLICE_X0Y25_D_XOR;
  assign CLBLL_L_X2Y25_SLICE_X1Y25_COUT = CLBLL_L_X2Y25_SLICE_X1Y25_D_CY;
  assign CLBLL_L_X2Y25_SLICE_X1Y25_A = CLBLL_L_X2Y25_SLICE_X1Y25_AO6;
  assign CLBLL_L_X2Y25_SLICE_X1Y25_B = CLBLL_L_X2Y25_SLICE_X1Y25_BO6;
  assign CLBLL_L_X2Y25_SLICE_X1Y25_C = CLBLL_L_X2Y25_SLICE_X1Y25_CO6;
  assign CLBLL_L_X2Y25_SLICE_X1Y25_D = CLBLL_L_X2Y25_SLICE_X1Y25_DO6;
  assign CLBLL_L_X2Y26_SLICE_X0Y26_COUT = CLBLL_L_X2Y26_SLICE_X0Y26_D_CY;
  assign CLBLL_L_X2Y26_SLICE_X0Y26_A = CLBLL_L_X2Y26_SLICE_X0Y26_AO6;
  assign CLBLL_L_X2Y26_SLICE_X0Y26_B = CLBLL_L_X2Y26_SLICE_X0Y26_BO6;
  assign CLBLL_L_X2Y26_SLICE_X0Y26_C = CLBLL_L_X2Y26_SLICE_X0Y26_CO6;
  assign CLBLL_L_X2Y26_SLICE_X0Y26_D = CLBLL_L_X2Y26_SLICE_X0Y26_DO6;
  assign CLBLL_L_X2Y26_SLICE_X0Y26_AMUX = CLBLL_L_X2Y26_SLICE_X0Y26_A_XOR;
  assign CLBLL_L_X2Y26_SLICE_X0Y26_BMUX = CLBLL_L_X2Y26_SLICE_X0Y26_B_XOR;
  assign CLBLL_L_X2Y26_SLICE_X0Y26_CMUX = CLBLL_L_X2Y26_SLICE_X0Y26_C_XOR;
  assign CLBLL_L_X2Y26_SLICE_X0Y26_DMUX = CLBLL_L_X2Y26_SLICE_X0Y26_D_XOR;
  assign CLBLL_L_X2Y26_SLICE_X1Y26_COUT = CLBLL_L_X2Y26_SLICE_X1Y26_D_CY;
  assign CLBLL_L_X2Y26_SLICE_X1Y26_A = CLBLL_L_X2Y26_SLICE_X1Y26_AO6;
  assign CLBLL_L_X2Y26_SLICE_X1Y26_B = CLBLL_L_X2Y26_SLICE_X1Y26_BO6;
  assign CLBLL_L_X2Y26_SLICE_X1Y26_C = CLBLL_L_X2Y26_SLICE_X1Y26_CO6;
  assign CLBLL_L_X2Y26_SLICE_X1Y26_D = CLBLL_L_X2Y26_SLICE_X1Y26_DO6;
  assign LIOI3_X0Y1_ILOGIC_X0Y2_O = LIOB33_X0Y1_IOB_X0Y2_I;
  assign LIOI3_X0Y1_ILOGIC_X0Y1_O = LIOB33_X0Y1_IOB_X0Y1_I;
  assign LIOI3_X0Y3_ILOGIC_X0Y4_O = LIOB33_X0Y3_IOB_X0Y4_I;
  assign LIOI3_X0Y3_ILOGIC_X0Y3_O = LIOB33_X0Y3_IOB_X0Y3_I;
  assign LIOI3_X0Y5_ILOGIC_X0Y6_O = LIOB33_X0Y5_IOB_X0Y6_I;
  assign LIOI3_X0Y5_ILOGIC_X0Y5_O = LIOB33_X0Y5_IOB_X0Y5_I;
  assign LIOI3_X0Y9_ILOGIC_X0Y10_O = LIOB33_X0Y9_IOB_X0Y10_I;
  assign LIOI3_X0Y9_ILOGIC_X0Y9_O = LIOB33_X0Y9_IOB_X0Y9_I;
  assign LIOI3_X0Y11_ILOGIC_X0Y12_O = LIOB33_X0Y11_IOB_X0Y12_I;
  assign LIOI3_X0Y11_ILOGIC_X0Y11_O = LIOB33_X0Y11_IOB_X0Y11_I;
  assign LIOI3_X0Y15_ILOGIC_X0Y16_O = LIOB33_X0Y15_IOB_X0Y16_I;
  assign LIOI3_X0Y15_ILOGIC_X0Y15_O = LIOB33_X0Y15_IOB_X0Y15_I;
  assign LIOI3_X0Y17_ILOGIC_X0Y18_O = LIOB33_X0Y17_IOB_X0Y18_I;
  assign LIOI3_X0Y17_ILOGIC_X0Y17_O = LIOB33_X0Y17_IOB_X0Y17_I;
  assign LIOI3_X0Y21_ILOGIC_X0Y22_O = LIOB33_X0Y21_IOB_X0Y22_I;
  assign LIOI3_X0Y21_ILOGIC_X0Y21_O = LIOB33_X0Y21_IOB_X0Y21_I;
  assign LIOI3_X0Y23_ILOGIC_X0Y24_O = LIOB33_X0Y23_IOB_X0Y24_I;
  assign LIOI3_X0Y23_ILOGIC_X0Y23_O = LIOB33_X0Y23_IOB_X0Y23_I;
  assign LIOI3_X0Y25_ILOGIC_X0Y26_O = LIOB33_X0Y25_IOB_X0Y26_I;
  assign LIOI3_X0Y25_ILOGIC_X0Y25_O = LIOB33_X0Y25_IOB_X0Y25_I;
  assign LIOI3_X0Y27_ILOGIC_X0Y28_O = LIOB33_X0Y27_IOB_X0Y28_I;
  assign LIOI3_X0Y27_ILOGIC_X0Y27_O = LIOB33_X0Y27_IOB_X0Y27_I;
  assign LIOI3_X0Y29_ILOGIC_X0Y30_O = LIOB33_X0Y29_IOB_X0Y30_I;
  assign LIOI3_X0Y29_ILOGIC_X0Y29_O = LIOB33_X0Y29_IOB_X0Y29_I;
  assign LIOI3_X0Y33_OLOGIC_X0Y34_OQ = CLBLL_L_X2Y23_SLICE_X0Y23_C_XOR;
  assign LIOI3_X0Y33_OLOGIC_X0Y34_TQ = 1'b1;
  assign LIOI3_X0Y33_OLOGIC_X0Y33_OQ = CLBLL_L_X2Y23_SLICE_X0Y23_B_XOR;
  assign LIOI3_X0Y33_OLOGIC_X0Y33_TQ = 1'b1;
  assign LIOI3_X0Y35_OLOGIC_X0Y36_OQ = CLBLL_L_X2Y24_SLICE_X0Y24_A_XOR;
  assign LIOI3_X0Y35_OLOGIC_X0Y36_TQ = 1'b1;
  assign LIOI3_X0Y35_OLOGIC_X0Y35_OQ = CLBLL_L_X2Y23_SLICE_X0Y23_D_XOR;
  assign LIOI3_X0Y35_OLOGIC_X0Y35_TQ = 1'b1;
  assign LIOI3_X0Y39_OLOGIC_X0Y40_OQ = CLBLL_L_X2Y25_SLICE_X0Y25_A_XOR;
  assign LIOI3_X0Y39_OLOGIC_X0Y40_TQ = 1'b1;
  assign LIOI3_X0Y39_OLOGIC_X0Y39_OQ = CLBLL_L_X2Y24_SLICE_X0Y24_D_XOR;
  assign LIOI3_X0Y39_OLOGIC_X0Y39_TQ = 1'b1;
  assign LIOI3_X0Y41_OLOGIC_X0Y42_OQ = CLBLL_L_X2Y25_SLICE_X0Y25_C_XOR;
  assign LIOI3_X0Y41_OLOGIC_X0Y42_TQ = 1'b1;
  assign LIOI3_X0Y41_OLOGIC_X0Y41_OQ = CLBLL_L_X2Y25_SLICE_X0Y25_B_XOR;
  assign LIOI3_X0Y41_OLOGIC_X0Y41_TQ = 1'b1;
  assign LIOI3_X0Y45_OLOGIC_X0Y46_OQ = CLBLL_L_X2Y26_SLICE_X0Y26_C_XOR;
  assign LIOI3_X0Y45_OLOGIC_X0Y46_TQ = 1'b1;
  assign LIOI3_X0Y45_OLOGIC_X0Y45_OQ = CLBLL_L_X2Y26_SLICE_X0Y26_B_XOR;
  assign LIOI3_X0Y45_OLOGIC_X0Y45_TQ = 1'b1;
  assign LIOI3_X0Y47_OLOGIC_X0Y47_OQ = CLBLL_L_X2Y26_SLICE_X0Y26_D_XOR;
  assign LIOI3_X0Y47_OLOGIC_X0Y47_TQ = 1'b1;
  assign LIOI3_SING_X0Y0_ILOGIC_X0Y0_O = LIOB33_SING_X0Y0_IOB_X0Y0_I;
  assign LIOI3_TBYTESRC_X0Y7_ILOGIC_X0Y8_O = LIOB33_X0Y7_IOB_X0Y8_I;
  assign LIOI3_TBYTESRC_X0Y7_ILOGIC_X0Y7_O = LIOB33_X0Y7_IOB_X0Y7_I;
  assign LIOI3_TBYTESRC_X0Y19_ILOGIC_X0Y20_O = LIOB33_X0Y19_IOB_X0Y20_I;
  assign LIOI3_TBYTESRC_X0Y19_ILOGIC_X0Y19_O = LIOB33_X0Y19_IOB_X0Y19_I;
  assign LIOI3_TBYTESRC_X0Y31_ILOGIC_X0Y31_O = LIOB33_X0Y31_IOB_X0Y31_I;
  assign LIOI3_TBYTESRC_X0Y31_OLOGIC_X0Y32_OQ = CLBLL_L_X2Y23_SLICE_X0Y23_A_XOR;
  assign LIOI3_TBYTESRC_X0Y31_OLOGIC_X0Y32_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y43_OLOGIC_X0Y44_OQ = CLBLL_L_X2Y26_SLICE_X0Y26_A_XOR;
  assign LIOI3_TBYTESRC_X0Y43_OLOGIC_X0Y44_TQ = 1'b1;
  assign LIOI3_TBYTESRC_X0Y43_OLOGIC_X0Y43_OQ = CLBLL_L_X2Y25_SLICE_X0Y25_D_XOR;
  assign LIOI3_TBYTESRC_X0Y43_OLOGIC_X0Y43_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y13_ILOGIC_X0Y14_O = LIOB33_X0Y13_IOB_X0Y14_I;
  assign LIOI3_TBYTETERM_X0Y13_ILOGIC_X0Y13_O = LIOB33_X0Y13_IOB_X0Y13_I;
  assign LIOI3_TBYTETERM_X0Y37_OLOGIC_X0Y38_OQ = CLBLL_L_X2Y24_SLICE_X0Y24_C_XOR;
  assign LIOI3_TBYTETERM_X0Y37_OLOGIC_X0Y38_TQ = 1'b1;
  assign LIOI3_TBYTETERM_X0Y37_OLOGIC_X0Y37_OQ = CLBLL_L_X2Y24_SLICE_X0Y24_B_XOR;
  assign LIOI3_TBYTETERM_X0Y37_OLOGIC_X0Y37_TQ = 1'b1;
  assign CLBLL_L_X2Y24_SLICE_X1Y24_C4 = 1'b1;
  assign CLBLL_L_X2Y24_SLICE_X1Y24_C5 = 1'b1;
  assign CLBLL_L_X2Y24_SLICE_X1Y24_C6 = 1'b1;
  assign LIOB33_X0Y37_IOB_X0Y38_O = CLBLL_L_X2Y24_SLICE_X0Y24_C_XOR;
  assign LIOB33_X0Y37_IOB_X0Y37_O = CLBLL_L_X2Y24_SLICE_X0Y24_B_XOR;
  assign LIOI3_TBYTETERM_X0Y37_OLOGIC_X0Y38_D1 = CLBLL_L_X2Y24_SLICE_X0Y24_C_XOR;
  assign CLBLL_L_X2Y24_SLICE_X1Y24_D1 = 1'b1;
  assign CLBLL_L_X2Y24_SLICE_X1Y24_D2 = 1'b1;
  assign CLBLL_L_X2Y24_SLICE_X1Y24_D3 = 1'b1;
  assign CLBLL_L_X2Y24_SLICE_X1Y24_D4 = 1'b1;
  assign CLBLL_L_X2Y24_SLICE_X1Y24_D5 = 1'b1;
  assign CLBLL_L_X2Y24_SLICE_X1Y24_D6 = 1'b1;
  assign LIOI3_X0Y9_ILOGIC_X0Y10_D = LIOB33_X0Y9_IOB_X0Y10_I;
  assign LIOI3_X0Y9_ILOGIC_X0Y9_D = LIOB33_X0Y9_IOB_X0Y9_I;
  assign LIOI3_X0Y47_OLOGIC_X0Y47_D1 = CLBLL_L_X2Y26_SLICE_X0Y26_D_XOR;
  assign LIOI3_TBYTETERM_X0Y37_OLOGIC_X0Y38_T1 = 1'b1;
  assign LIOI3_X0Y47_OLOGIC_X0Y47_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y31_OLOGIC_X0Y32_T1 = 1'b1;
  assign LIOI3_TBYTETERM_X0Y37_OLOGIC_X0Y37_D1 = CLBLL_L_X2Y24_SLICE_X0Y24_B_XOR;
  assign LIOI3_TBYTETERM_X0Y37_OLOGIC_X0Y37_T1 = 1'b1;
  assign LIOI3_X0Y35_OLOGIC_X0Y36_D1 = CLBLL_L_X2Y24_SLICE_X0Y24_A_XOR;
  assign LIOI3_X0Y35_OLOGIC_X0Y36_T1 = 1'b1;
  assign LIOI3_X0Y27_ILOGIC_X0Y28_D = LIOB33_X0Y27_IOB_X0Y28_I;
  assign LIOI3_X0Y35_OLOGIC_X0Y35_D1 = CLBLL_L_X2Y23_SLICE_X0Y23_D_XOR;
  assign LIOI3_X0Y27_ILOGIC_X0Y27_D = LIOB33_X0Y27_IOB_X0Y27_I;
  assign LIOB33_X0Y45_IOB_X0Y46_O = CLBLL_L_X2Y26_SLICE_X0Y26_C_XOR;
  assign LIOB33_X0Y45_IOB_X0Y45_O = CLBLL_L_X2Y26_SLICE_X0Y26_B_XOR;
  assign LIOI3_X0Y35_OLOGIC_X0Y35_T1 = 1'b1;
  assign LIOB33_X0Y31_IOB_X0Y32_O = CLBLL_L_X2Y23_SLICE_X0Y23_A_XOR;
  assign CLBLL_L_X2Y26_SLICE_X1Y26_D3 = 1'b1;
  assign CLBLL_L_X2Y26_SLICE_X1Y26_D4 = 1'b1;
  assign CLBLL_L_X2Y26_SLICE_X1Y26_D5 = 1'b1;
  assign CLBLL_L_X2Y26_SLICE_X1Y26_D6 = 1'b1;
  assign LIOI3_X0Y17_ILOGIC_X0Y18_D = LIOB33_X0Y17_IOB_X0Y18_I;
  assign LIOI3_X0Y17_ILOGIC_X0Y17_D = LIOB33_X0Y17_IOB_X0Y17_I;
  assign CLBLL_L_X2Y25_SLICE_X0Y25_A1 = 1'b1;
  assign CLBLL_L_X2Y25_SLICE_X0Y25_A2 = 1'b1;
  assign CLBLL_L_X2Y25_SLICE_X0Y25_A3 = LIOB33_X0Y23_IOB_X0Y24_I;
  assign CLBLL_L_X2Y25_SLICE_X0Y25_A4 = 1'b1;
  assign CLBLL_L_X2Y25_SLICE_X0Y25_A5 = LIOB33_X0Y7_IOB_X0Y8_I;
  assign CLBLL_L_X2Y25_SLICE_X0Y25_A6 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y31_ILOGIC_X0Y31_D = LIOB33_X0Y31_IOB_X0Y31_I;
  assign CLBLL_L_X2Y25_SLICE_X0Y25_AX = LIOB33_X0Y7_IOB_X0Y8_I;
  assign CLBLL_L_X2Y25_SLICE_X0Y25_B1 = LIOB33_X0Y9_IOB_X0Y9_I;
  assign CLBLL_L_X2Y25_SLICE_X0Y25_B2 = 1'b1;
  assign CLBLL_L_X2Y25_SLICE_X0Y25_B3 = LIOB33_X0Y25_IOB_X0Y25_I;
  assign CLBLL_L_X2Y25_SLICE_X0Y25_B4 = 1'b1;
  assign CLBLL_L_X2Y25_SLICE_X0Y25_B5 = 1'b1;
  assign CLBLL_L_X2Y25_SLICE_X0Y25_B6 = 1'b1;
  assign CLBLL_L_X2Y25_SLICE_X0Y25_BX = LIOB33_X0Y9_IOB_X0Y9_I;
  assign CLBLL_L_X2Y25_SLICE_X0Y25_C1 = LIOB33_X0Y9_IOB_X0Y10_I;
  assign CLBLL_L_X2Y25_SLICE_X0Y25_C2 = 1'b1;
  assign CLBLL_L_X2Y25_SLICE_X0Y25_C3 = 1'b1;
  assign CLBLL_L_X2Y25_SLICE_X0Y25_C4 = 1'b1;
  assign CLBLL_L_X2Y25_SLICE_X0Y25_C5 = 1'b1;
  assign CLBLL_L_X2Y25_SLICE_X0Y25_C6 = LIOB33_X0Y25_IOB_X0Y26_I;
  assign CLBLL_L_X2Y25_SLICE_X0Y25_CIN = CLBLL_L_X2Y24_SLICE_X0Y24_D_CY;
  assign CLBLL_L_X2Y25_SLICE_X0Y25_CX = LIOB33_X0Y9_IOB_X0Y10_I;
  assign CLBLL_L_X2Y25_SLICE_X0Y25_D1 = LIOB33_X0Y11_IOB_X0Y11_I;
  assign CLBLL_L_X2Y25_SLICE_X0Y25_D2 = 1'b1;
  assign CLBLL_L_X2Y25_SLICE_X0Y25_D3 = LIOB33_X0Y27_IOB_X0Y27_I;
  assign CLBLL_L_X2Y25_SLICE_X0Y25_D4 = 1'b1;
  assign CLBLL_L_X2Y25_SLICE_X0Y25_D5 = 1'b1;
  assign CLBLL_L_X2Y25_SLICE_X0Y25_D6 = 1'b1;
  assign CLBLL_L_X2Y25_SLICE_X0Y25_DX = LIOB33_X0Y11_IOB_X0Y11_I;
  assign LIOI3_X0Y45_OLOGIC_X0Y46_D1 = CLBLL_L_X2Y26_SLICE_X0Y26_C_XOR;
  assign LIOI3_X0Y45_OLOGIC_X0Y46_T1 = 1'b1;
  assign CLBLL_L_X2Y25_SLICE_X1Y25_A1 = 1'b1;
  assign CLBLL_L_X2Y25_SLICE_X1Y25_A2 = 1'b1;
  assign CLBLL_L_X2Y25_SLICE_X1Y25_A3 = 1'b1;
  assign CLBLL_L_X2Y25_SLICE_X1Y25_A4 = 1'b1;
  assign CLBLL_L_X2Y25_SLICE_X1Y25_A5 = 1'b1;
  assign CLBLL_L_X2Y25_SLICE_X1Y25_A6 = 1'b1;
  assign LIOB33_X0Y39_IOB_X0Y39_O = CLBLL_L_X2Y24_SLICE_X0Y24_D_XOR;
  assign LIOB33_X0Y39_IOB_X0Y40_O = CLBLL_L_X2Y25_SLICE_X0Y25_A_XOR;
  assign LIOI3_X0Y45_OLOGIC_X0Y45_D1 = CLBLL_L_X2Y26_SLICE_X0Y26_B_XOR;
  assign CLBLL_L_X2Y25_SLICE_X1Y25_B1 = 1'b1;
  assign CLBLL_L_X2Y25_SLICE_X1Y25_B2 = 1'b1;
  assign CLBLL_L_X2Y25_SLICE_X1Y25_B3 = 1'b1;
  assign CLBLL_L_X2Y25_SLICE_X1Y25_B4 = 1'b1;
  assign CLBLL_L_X2Y25_SLICE_X1Y25_B5 = 1'b1;
  assign CLBLL_L_X2Y25_SLICE_X1Y25_B6 = 1'b1;
  assign LIOI3_X0Y5_ILOGIC_X0Y6_D = LIOB33_X0Y5_IOB_X0Y6_I;
  assign CLBLL_L_X2Y25_SLICE_X1Y25_C1 = 1'b1;
  assign CLBLL_L_X2Y25_SLICE_X1Y25_C2 = 1'b1;
  assign CLBLL_L_X2Y25_SLICE_X1Y25_C3 = 1'b1;
  assign CLBLL_L_X2Y25_SLICE_X1Y25_C4 = 1'b1;
  assign CLBLL_L_X2Y25_SLICE_X1Y25_C5 = 1'b1;
  assign CLBLL_L_X2Y25_SLICE_X1Y25_C6 = 1'b1;
  assign LIOI3_X0Y45_OLOGIC_X0Y45_T1 = 1'b1;
  assign CLBLL_L_X2Y25_SLICE_X1Y25_D1 = 1'b1;
  assign CLBLL_L_X2Y25_SLICE_X1Y25_D2 = 1'b1;
  assign CLBLL_L_X2Y25_SLICE_X1Y25_D3 = 1'b1;
  assign CLBLL_L_X2Y25_SLICE_X1Y25_D4 = 1'b1;
  assign CLBLL_L_X2Y25_SLICE_X1Y25_D5 = 1'b1;
  assign CLBLL_L_X2Y25_SLICE_X1Y25_D6 = 1'b1;
  assign LIOI3_X0Y33_OLOGIC_X0Y34_D1 = CLBLL_L_X2Y23_SLICE_X0Y23_C_XOR;
  assign LIOI3_X0Y33_OLOGIC_X0Y34_T1 = 1'b1;
  assign LIOI3_X0Y25_ILOGIC_X0Y26_D = LIOB33_X0Y25_IOB_X0Y26_I;
  assign LIOI3_X0Y25_ILOGIC_X0Y25_D = LIOB33_X0Y25_IOB_X0Y25_I;
  assign LIOI3_X0Y33_OLOGIC_X0Y33_D1 = CLBLL_L_X2Y23_SLICE_X0Y23_B_XOR;
  assign LIOB33_X0Y47_IOB_X0Y47_O = CLBLL_L_X2Y26_SLICE_X0Y26_D_XOR;
  assign LIOI3_X0Y33_OLOGIC_X0Y33_T1 = 1'b1;
  assign LIOB33_X0Y33_IOB_X0Y34_O = CLBLL_L_X2Y23_SLICE_X0Y23_C_XOR;
  assign LIOB33_X0Y33_IOB_X0Y33_O = CLBLL_L_X2Y23_SLICE_X0Y23_B_XOR;
  assign LIOI3_X0Y15_ILOGIC_X0Y16_D = LIOB33_X0Y15_IOB_X0Y16_I;
  assign LIOI3_X0Y15_ILOGIC_X0Y15_D = LIOB33_X0Y15_IOB_X0Y15_I;
  assign LIOI3_TBYTETERM_X0Y13_ILOGIC_X0Y14_D = LIOB33_X0Y13_IOB_X0Y14_I;
  assign LIOI3_TBYTETERM_X0Y13_ILOGIC_X0Y13_D = LIOB33_X0Y13_IOB_X0Y13_I;
  assign LIOI3_X0Y5_ILOGIC_X0Y5_D = LIOB33_X0Y5_IOB_X0Y5_I;
  assign LIOI3_TBYTESRC_X0Y19_ILOGIC_X0Y20_D = LIOB33_X0Y19_IOB_X0Y20_I;
  assign LIOI3_TBYTESRC_X0Y19_ILOGIC_X0Y19_D = LIOB33_X0Y19_IOB_X0Y19_I;
  assign CLBLL_L_X2Y26_SLICE_X0Y26_A1 = LIOB33_X0Y27_IOB_X0Y28_I;
  assign CLBLL_L_X2Y26_SLICE_X0Y26_A2 = 1'b1;
  assign CLBLL_L_X2Y26_SLICE_X0Y26_A3 = LIOB33_X0Y11_IOB_X0Y12_I;
  assign CLBLL_L_X2Y26_SLICE_X0Y26_A4 = 1'b1;
  assign CLBLL_L_X2Y26_SLICE_X0Y26_A5 = 1'b1;
  assign CLBLL_L_X2Y26_SLICE_X0Y26_A6 = 1'b1;
  assign CLBLL_L_X2Y26_SLICE_X0Y26_AX = LIOB33_X0Y11_IOB_X0Y12_I;
  assign CLBLL_L_X2Y26_SLICE_X0Y26_B1 = 1'b1;
  assign CLBLL_L_X2Y26_SLICE_X0Y26_B2 = LIOB33_X0Y13_IOB_X0Y13_I;
  assign CLBLL_L_X2Y26_SLICE_X0Y26_B3 = 1'b1;
  assign CLBLL_L_X2Y26_SLICE_X0Y26_B4 = 1'b1;
  assign CLBLL_L_X2Y26_SLICE_X0Y26_B5 = LIOB33_X0Y29_IOB_X0Y29_I;
  assign CLBLL_L_X2Y26_SLICE_X0Y26_B6 = 1'b1;
  assign CLBLL_L_X2Y26_SLICE_X0Y26_BX = LIOB33_X0Y13_IOB_X0Y13_I;
  assign CLBLL_L_X2Y26_SLICE_X0Y26_C1 = LIOB33_X0Y13_IOB_X0Y14_I;
  assign CLBLL_L_X2Y26_SLICE_X0Y26_C2 = 1'b1;
  assign CLBLL_L_X2Y26_SLICE_X0Y26_C3 = 1'b1;
  assign CLBLL_L_X2Y26_SLICE_X0Y26_C4 = 1'b1;
  assign CLBLL_L_X2Y26_SLICE_X0Y26_C5 = 1'b1;
  assign CLBLL_L_X2Y26_SLICE_X0Y26_C6 = LIOB33_X0Y29_IOB_X0Y30_I;
  assign LIOI3_X0Y41_OLOGIC_X0Y42_D1 = CLBLL_L_X2Y25_SLICE_X0Y25_C_XOR;
  assign CLBLL_L_X2Y26_SLICE_X0Y26_CIN = CLBLL_L_X2Y25_SLICE_X0Y25_D_CY;
  assign CLBLL_L_X2Y26_SLICE_X0Y26_CX = LIOB33_X0Y13_IOB_X0Y14_I;
  assign CLBLL_L_X2Y26_SLICE_X0Y26_D1 = LIOB33_X0Y15_IOB_X0Y15_I;
  assign CLBLL_L_X2Y26_SLICE_X0Y26_D2 = 1'b1;
  assign CLBLL_L_X2Y26_SLICE_X0Y26_D3 = LIOB33_X0Y31_IOB_X0Y31_I;
  assign CLBLL_L_X2Y26_SLICE_X0Y26_D4 = 1'b1;
  assign CLBLL_L_X2Y26_SLICE_X0Y26_D5 = 1'b1;
  assign CLBLL_L_X2Y26_SLICE_X0Y26_D6 = 1'b1;
  assign LIOI3_X0Y41_OLOGIC_X0Y42_T1 = 1'b1;
  assign CLBLL_L_X2Y26_SLICE_X0Y26_DX = 1'b0;
  assign LIOB33_X0Y41_IOB_X0Y42_O = CLBLL_L_X2Y25_SLICE_X0Y25_C_XOR;
  assign LIOB33_X0Y41_IOB_X0Y41_O = CLBLL_L_X2Y25_SLICE_X0Y25_B_XOR;
  assign LIOI3_X0Y41_OLOGIC_X0Y41_D1 = CLBLL_L_X2Y25_SLICE_X0Y25_B_XOR;
  assign LIOI3_X0Y3_ILOGIC_X0Y4_D = LIOB33_X0Y3_IOB_X0Y4_I;
  assign LIOI3_X0Y3_ILOGIC_X0Y3_D = LIOB33_X0Y3_IOB_X0Y3_I;
  assign LIOI3_X0Y41_OLOGIC_X0Y41_T1 = 1'b1;
  assign CLBLL_L_X2Y26_SLICE_X1Y26_A1 = 1'b1;
  assign CLBLL_L_X2Y26_SLICE_X1Y26_A2 = 1'b1;
  assign CLBLL_L_X2Y26_SLICE_X1Y26_A3 = 1'b1;
  assign CLBLL_L_X2Y26_SLICE_X1Y26_A4 = 1'b1;
  assign CLBLL_L_X2Y26_SLICE_X1Y26_A5 = 1'b1;
  assign CLBLL_L_X2Y26_SLICE_X1Y26_A6 = 1'b1;
  assign CLBLL_L_X2Y26_SLICE_X1Y26_B1 = 1'b1;
  assign CLBLL_L_X2Y26_SLICE_X1Y26_B2 = 1'b1;
  assign CLBLL_L_X2Y26_SLICE_X1Y26_B3 = 1'b1;
  assign CLBLL_L_X2Y26_SLICE_X1Y26_B4 = 1'b1;
  assign CLBLL_L_X2Y26_SLICE_X1Y26_B5 = 1'b1;
  assign CLBLL_L_X2Y26_SLICE_X1Y26_B6 = 1'b1;
  assign CLBLL_L_X2Y26_SLICE_X1Y26_C1 = 1'b1;
  assign CLBLL_L_X2Y26_SLICE_X1Y26_C2 = 1'b1;
  assign CLBLL_L_X2Y26_SLICE_X1Y26_C3 = 1'b1;
  assign CLBLL_L_X2Y26_SLICE_X1Y26_C4 = 1'b1;
  assign CLBLL_L_X2Y23_SLICE_X0Y23_A1 = LIOB33_SING_X0Y0_IOB_X0Y0_I;
  assign CLBLL_L_X2Y23_SLICE_X0Y23_A2 = 1'b1;
  assign CLBLL_L_X2Y23_SLICE_X0Y23_A3 = 1'b1;
  assign CLBLL_L_X2Y23_SLICE_X0Y23_A4 = 1'b1;
  assign CLBLL_L_X2Y23_SLICE_X0Y23_A5 = LIOB33_X0Y15_IOB_X0Y16_I;
  assign CLBLL_L_X2Y23_SLICE_X0Y23_A6 = 1'b1;
  assign CLBLL_L_X2Y26_SLICE_X1Y26_C5 = 1'b1;
  assign CLBLL_L_X2Y26_SLICE_X1Y26_C6 = 1'b1;
  assign CLBLL_L_X2Y23_SLICE_X0Y23_AX = LIOB33_SING_X0Y0_IOB_X0Y0_I;
  assign CLBLL_L_X2Y23_SLICE_X0Y23_B1 = LIOB33_X0Y1_IOB_X0Y1_I;
  assign CLBLL_L_X2Y23_SLICE_X0Y23_B2 = 1'b1;
  assign CLBLL_L_X2Y23_SLICE_X0Y23_B3 = LIOB33_X0Y17_IOB_X0Y17_I;
  assign CLBLL_L_X2Y23_SLICE_X0Y23_B4 = 1'b1;
  assign CLBLL_L_X2Y23_SLICE_X0Y23_B5 = 1'b1;
  assign CLBLL_L_X2Y23_SLICE_X0Y23_B6 = 1'b1;
  assign CLBLL_L_X2Y26_SLICE_X1Y26_D1 = 1'b1;
  assign CLBLL_L_X2Y26_SLICE_X1Y26_D2 = 1'b1;
  assign CLBLL_L_X2Y23_SLICE_X0Y23_BX = LIOB33_X0Y1_IOB_X0Y1_I;
  assign CLBLL_L_X2Y23_SLICE_X0Y23_C1 = LIOB33_X0Y17_IOB_X0Y18_I;
  assign CLBLL_L_X2Y23_SLICE_X0Y23_C2 = 1'b1;
  assign CLBLL_L_X2Y23_SLICE_X0Y23_C3 = LIOB33_X0Y1_IOB_X0Y2_I;
  assign CLBLL_L_X2Y23_SLICE_X0Y23_C4 = 1'b1;
  assign CLBLL_L_X2Y23_SLICE_X0Y23_C5 = 1'b1;
  assign CLBLL_L_X2Y23_SLICE_X0Y23_C6 = 1'b1;
  assign CLBLL_L_X2Y23_SLICE_X0Y23_CX = LIOB33_X0Y1_IOB_X0Y2_I;
  assign CLBLL_L_X2Y23_SLICE_X0Y23_D1 = LIOB33_X0Y3_IOB_X0Y3_I;
  assign CLBLL_L_X2Y23_SLICE_X0Y23_D2 = LIOB33_X0Y19_IOB_X0Y19_I;
  assign CLBLL_L_X2Y23_SLICE_X0Y23_D3 = 1'b1;
  assign CLBLL_L_X2Y23_SLICE_X0Y23_D4 = 1'b1;
  assign CLBLL_L_X2Y23_SLICE_X0Y23_D5 = 1'b1;
  assign CLBLL_L_X2Y23_SLICE_X0Y23_D6 = 1'b1;
  assign CLBLL_L_X2Y23_SLICE_X0Y23_DX = LIOB33_X0Y3_IOB_X0Y3_I;
  assign LIOI3_X0Y23_ILOGIC_X0Y24_D = LIOB33_X0Y23_IOB_X0Y24_I;
  assign LIOI3_X0Y23_ILOGIC_X0Y23_D = LIOB33_X0Y23_IOB_X0Y23_I;
  assign LIOI3_TBYTESRC_X0Y31_OLOGIC_X0Y32_D1 = CLBLL_L_X2Y23_SLICE_X0Y23_A_XOR;
  assign CLBLL_L_X2Y23_SLICE_X1Y23_A1 = 1'b1;
  assign CLBLL_L_X2Y23_SLICE_X1Y23_A2 = 1'b1;
  assign CLBLL_L_X2Y23_SLICE_X1Y23_A3 = 1'b1;
  assign CLBLL_L_X2Y23_SLICE_X1Y23_A4 = 1'b1;
  assign CLBLL_L_X2Y23_SLICE_X1Y23_A5 = 1'b1;
  assign CLBLL_L_X2Y23_SLICE_X1Y23_A6 = 1'b1;
  assign CLBLL_L_X2Y23_SLICE_X1Y23_B1 = 1'b1;
  assign CLBLL_L_X2Y23_SLICE_X1Y23_B2 = 1'b1;
  assign CLBLL_L_X2Y23_SLICE_X1Y23_B3 = 1'b1;
  assign CLBLL_L_X2Y23_SLICE_X1Y23_B4 = 1'b1;
  assign CLBLL_L_X2Y23_SLICE_X1Y23_B5 = 1'b1;
  assign CLBLL_L_X2Y23_SLICE_X1Y23_B6 = 1'b1;
  assign CLBLL_L_X2Y23_SLICE_X1Y23_C1 = 1'b1;
  assign CLBLL_L_X2Y23_SLICE_X1Y23_C2 = 1'b1;
  assign CLBLL_L_X2Y23_SLICE_X1Y23_C3 = 1'b1;
  assign CLBLL_L_X2Y23_SLICE_X1Y23_C4 = 1'b1;
  assign CLBLL_L_X2Y23_SLICE_X1Y23_C5 = 1'b1;
  assign CLBLL_L_X2Y23_SLICE_X1Y23_C6 = 1'b1;
  assign CLBLL_L_X2Y23_SLICE_X1Y23_D1 = 1'b1;
  assign CLBLL_L_X2Y23_SLICE_X1Y23_D2 = 1'b1;
  assign CLBLL_L_X2Y23_SLICE_X1Y23_D3 = 1'b1;
  assign CLBLL_L_X2Y23_SLICE_X1Y23_D4 = 1'b1;
  assign CLBLL_L_X2Y23_SLICE_X1Y23_D5 = 1'b1;
  assign CLBLL_L_X2Y23_SLICE_X1Y23_D6 = 1'b1;
  assign LIOB33_X0Y35_IOB_X0Y36_O = CLBLL_L_X2Y24_SLICE_X0Y24_A_XOR;
  assign LIOB33_X0Y35_IOB_X0Y35_O = CLBLL_L_X2Y23_SLICE_X0Y23_D_XOR;
  assign LIOI3_TBYTESRC_X0Y43_OLOGIC_X0Y44_D1 = CLBLL_L_X2Y26_SLICE_X0Y26_A_XOR;
  assign LIOI3_X0Y11_ILOGIC_X0Y12_D = LIOB33_X0Y11_IOB_X0Y12_I;
  assign LIOI3_X0Y11_ILOGIC_X0Y11_D = LIOB33_X0Y11_IOB_X0Y11_I;
  assign LIOI3_TBYTESRC_X0Y43_OLOGIC_X0Y44_T1 = 1'b1;
  assign LIOI3_TBYTESRC_X0Y7_ILOGIC_X0Y8_D = LIOB33_X0Y7_IOB_X0Y8_I;
  assign LIOI3_TBYTESRC_X0Y7_ILOGIC_X0Y7_D = LIOB33_X0Y7_IOB_X0Y7_I;
  assign LIOI3_TBYTESRC_X0Y43_OLOGIC_X0Y43_D1 = CLBLL_L_X2Y25_SLICE_X0Y25_D_XOR;
  assign LIOI3_TBYTESRC_X0Y43_OLOGIC_X0Y43_T1 = 1'b1;
  assign LIOI3_X0Y39_OLOGIC_X0Y40_D1 = CLBLL_L_X2Y25_SLICE_X0Y25_A_XOR;
  assign LIOI3_X0Y39_OLOGIC_X0Y40_T1 = 1'b1;
  assign LIOI3_X0Y29_ILOGIC_X0Y30_D = LIOB33_X0Y29_IOB_X0Y30_I;
  assign LIOI3_X0Y29_ILOGIC_X0Y29_D = LIOB33_X0Y29_IOB_X0Y29_I;
  assign LIOI3_X0Y39_OLOGIC_X0Y39_D1 = CLBLL_L_X2Y24_SLICE_X0Y24_D_XOR;
  assign LIOB33_X0Y43_IOB_X0Y44_O = CLBLL_L_X2Y26_SLICE_X0Y26_A_XOR;
  assign LIOB33_X0Y43_IOB_X0Y43_O = CLBLL_L_X2Y25_SLICE_X0Y25_D_XOR;
  assign LIOI3_X0Y1_ILOGIC_X0Y2_D = LIOB33_X0Y1_IOB_X0Y2_I;
  assign LIOI3_X0Y1_ILOGIC_X0Y1_D = LIOB33_X0Y1_IOB_X0Y1_I;
  assign LIOI3_X0Y39_OLOGIC_X0Y39_T1 = 1'b1;
  assign CLBLL_L_X2Y24_SLICE_X0Y24_A1 = 1'b1;
  assign CLBLL_L_X2Y24_SLICE_X0Y24_A2 = 1'b1;
  assign CLBLL_L_X2Y24_SLICE_X0Y24_A3 = 1'b1;
  assign CLBLL_L_X2Y24_SLICE_X0Y24_A4 = LIOB33_X0Y3_IOB_X0Y4_I;
  assign CLBLL_L_X2Y24_SLICE_X0Y24_A5 = LIOB33_X0Y19_IOB_X0Y20_I;
  assign CLBLL_L_X2Y24_SLICE_X0Y24_A6 = 1'b1;
  assign CLBLL_L_X2Y24_SLICE_X0Y24_AX = LIOB33_X0Y3_IOB_X0Y4_I;
  assign CLBLL_L_X2Y24_SLICE_X0Y24_B1 = LIOB33_X0Y5_IOB_X0Y5_I;
  assign CLBLL_L_X2Y24_SLICE_X0Y24_B2 = 1'b1;
  assign CLBLL_L_X2Y24_SLICE_X0Y24_B3 = LIOB33_X0Y21_IOB_X0Y21_I;
  assign CLBLL_L_X2Y24_SLICE_X0Y24_B4 = 1'b1;
  assign CLBLL_L_X2Y24_SLICE_X0Y24_B5 = 1'b1;
  assign CLBLL_L_X2Y24_SLICE_X0Y24_B6 = 1'b1;
  assign LIOI3_X0Y21_ILOGIC_X0Y22_D = LIOB33_X0Y21_IOB_X0Y22_I;
  assign CLBLL_L_X2Y24_SLICE_X0Y24_BX = LIOB33_X0Y5_IOB_X0Y5_I;
  assign LIOI3_X0Y21_ILOGIC_X0Y21_D = LIOB33_X0Y21_IOB_X0Y21_I;
  assign CLBLL_L_X2Y24_SLICE_X0Y24_C1 = LIOB33_X0Y21_IOB_X0Y22_I;
  assign CLBLL_L_X2Y24_SLICE_X0Y24_C2 = 1'b1;
  assign CLBLL_L_X2Y24_SLICE_X0Y24_C3 = LIOB33_X0Y5_IOB_X0Y6_I;
  assign CLBLL_L_X2Y24_SLICE_X0Y24_C4 = 1'b1;
  assign CLBLL_L_X2Y24_SLICE_X0Y24_C5 = 1'b1;
  assign CLBLL_L_X2Y24_SLICE_X0Y24_C6 = 1'b1;
  assign CLBLL_L_X2Y24_SLICE_X0Y24_CIN = CLBLL_L_X2Y23_SLICE_X0Y23_D_CY;
  assign CLBLL_L_X2Y24_SLICE_X0Y24_CX = LIOB33_X0Y5_IOB_X0Y6_I;
  assign CLBLL_L_X2Y24_SLICE_X0Y24_D1 = LIOB33_X0Y23_IOB_X0Y23_I;
  assign CLBLL_L_X2Y24_SLICE_X0Y24_D2 = LIOB33_X0Y7_IOB_X0Y7_I;
  assign CLBLL_L_X2Y24_SLICE_X0Y24_D3 = 1'b1;
  assign CLBLL_L_X2Y24_SLICE_X0Y24_D4 = 1'b1;
  assign CLBLL_L_X2Y24_SLICE_X0Y24_D5 = 1'b1;
  assign CLBLL_L_X2Y24_SLICE_X0Y24_D6 = 1'b1;
  assign LIOI3_SING_X0Y0_ILOGIC_X0Y0_D = LIOB33_SING_X0Y0_IOB_X0Y0_I;
  assign CLBLL_L_X2Y24_SLICE_X0Y24_DX = LIOB33_X0Y7_IOB_X0Y7_I;
  assign CLBLL_L_X2Y24_SLICE_X1Y24_A1 = 1'b1;
  assign CLBLL_L_X2Y24_SLICE_X1Y24_A2 = 1'b1;
  assign CLBLL_L_X2Y24_SLICE_X1Y24_A3 = 1'b1;
  assign CLBLL_L_X2Y24_SLICE_X1Y24_A4 = 1'b1;
  assign CLBLL_L_X2Y24_SLICE_X1Y24_A5 = 1'b1;
  assign CLBLL_L_X2Y24_SLICE_X1Y24_A6 = 1'b1;
  assign CLBLL_L_X2Y24_SLICE_X1Y24_B1 = 1'b1;
  assign CLBLL_L_X2Y24_SLICE_X1Y24_B2 = 1'b1;
  assign CLBLL_L_X2Y24_SLICE_X1Y24_B3 = 1'b1;
  assign CLBLL_L_X2Y24_SLICE_X1Y24_B4 = 1'b1;
  assign CLBLL_L_X2Y24_SLICE_X1Y24_B5 = 1'b1;
  assign CLBLL_L_X2Y24_SLICE_X1Y24_B6 = 1'b1;
  assign CLBLL_L_X2Y24_SLICE_X1Y24_C1 = 1'b1;
  assign CLBLL_L_X2Y24_SLICE_X1Y24_C2 = 1'b1;
  assign CLBLL_L_X2Y24_SLICE_X1Y24_C3 = 1'b1;
endmodule