module times ();
   time x;
   initial x = 33ns;	// Note no space
endmodule