module top ;
          wire  Net_829;
          wire  Net_828;
          wire  Net_827;
          wire  Net_826;
          wire  Net_825;
          wire  Net_824;
          wire  Net_823;
          wire  Net_822;
          wire  Net_821;
          wire  Net_820;
          wire  Net_778;
          wire  Net_777;
          wire  Net_776;
          wire  Net_775;
          wire  Net_774;
          wire  Net_773;
          wire  Net_772;
          wire  Net_771;
          wire  Net_770;
          wire  Net_769;
          wire  Net_757;
          wire  Net_756;
          wire  Net_872;
          wire  Net_864;
          wire  Net_863;
          wire  Net_681;
          wire  Net_862;
          wire  Net_861;
          wire  Net_678;
          wire  Net_676;
          wire  Net_675;
          wire  Net_768;
          wire  Net_767;
          wire  Net_766;
          wire  Net_765;
          wire  Net_764;
          wire  Net_763;
          wire  Net_762;
          wire  Net_761;
          wire  Net_760;
          wire  Net_759;
          wire  Net_505;
          wire  Net_504;
          wire  Net_132;
          wire  Net_609;
          wire  Net_608;
          wire  Net_607;
          wire  Net_606;
          wire  Net_605;
          wire  Net_604;
          wire  Net_603;
          wire  Net_602;
          wire  Net_601;
          wire  Net_519;
          wire  Net_518;
          wire  Net_600;
          wire  Net_599;
          wire  Net_80;
          wire  Net_79;
          wire  Net_78;
          wire  Net_77;
          wire  Net_76;
          wire  Net_75;
          wire  Net_74;
          wire  Net_73;
          wire  Net_72;
          wire  Net_71;
          wire  Net_6;
          wire  Net_4;
          wire  Net_747;
          wire  Net_701;
          wire  Net_496;
          wire  Net_49;
          wire  Net_5;
    SCB_P4_v1_20_0 UART_1 (
        .sclk(Net_4),
        .interrupt(Net_5),
        .clock(1'b0));
	cy_isr_v1_0
		#(.int_type(2'b10))
		isr
		 (.int_signal(Net_49));
    TCPWM_P4_v1_10_1 Timer (
        .stop(1'b0),
        .reload(1'b0),
        .start(1'b0),
        .count(1'b1),
        .capture(1'b0),
        .interrupt(Net_49),
        .ov(Net_76),
        .un(Net_77),
        .cc(Net_78),
        .line(Net_79),
        .line_n(Net_80),
        .clock(Net_496));
    defparam Timer.PWMCountMode = 3;
    defparam Timer.PWMReloadMode = 0;
    defparam Timer.PWMReloadPresent = 0;
    defparam Timer.PWMStartMode = 0;
    defparam Timer.PWMStopMode = 0;
    defparam Timer.PWMSwitchMode = 0;
    defparam Timer.QuadIndexMode = 0;
    defparam Timer.QuadPhiAMode = 3;
    defparam Timer.QuadPhiBMode = 3;
    defparam Timer.QuadStopMode = 0;
    defparam Timer.TCCaptureMode = 0;
    defparam Timer.TCCountMode = 3;
    defparam Timer.TCReloadMode = 0;
    defparam Timer.TCStartMode = 0;
    defparam Timer.TCStopMode = 0;
	cy_isr_v1_0
		#(.int_type(2'b10))
		ISRUART
		 (.int_signal(Net_5));
    PWM_v3_0_2 Gimbal (
        .reset(1'b0),
        .clock(Net_496),
        .tc(Net_600),
        .pwm1(Net_518),
        .pwm2(Net_519),
        .interrupt(Net_601),
        .capture(1'b0),
        .kill(1'b1),
        .enable(1'b1),
        .trigger(1'b0),
        .cmp_sel(1'b0),
        .pwm(Net_607),
        .ph1(Net_608),
        .ph2(Net_609));
    defparam Gimbal.Resolution = 16;
	cy_clock_v1_0
		#(.id("77085c73-d3db-49de-a1ad-2dc98b341901"),
		  .source_clock_id(""),
		  .divisor(0),
		  .period("1000000000"),
		  .is_direct(0),
		  .is_digital(1))
		Clock_2
		 (.clock_out(Net_496));
	wire [0:0] tmpOE__L_Servo_net;
	wire [0:0] tmpFB_0__L_Servo_net;
	wire [0:0] tmpIO_0__L_Servo_net;
	wire [0:0] tmpINTERRUPT_0__L_Servo_net;
	electrical [0:0] tmpSIOVREF__L_Servo_net;
	cy_psoc3_pins_v1_10
		#(.id("52f31aa9-2f0a-497d-9a1f-1424095e13e6"),
		  .drive_mode(3'b110),
		  .ibuf_enabled(1'b1),
		  .init_dr_st(1'b1),
		  .input_clk_en(0),
		  .input_sync(1'b1),
		  .input_sync_mode(1'b0),
		  .intr_mode(2'b00),
		  .invert_in_clock(0),
		  .invert_in_clock_en(0),
		  .invert_in_reset(0),
		  .invert_out_clock(0),
		  .invert_out_clock_en(0),
		  .invert_out_reset(0),
		  .io_voltage(""),
		  .layout_mode("CONTIGUOUS"),
		  .oe_conn(1'b0),
		  .oe_reset(0),
		  .oe_sync(1'b0),
		  .output_clk_en(0),
		  .output_clock_mode(1'b0),
		  .output_conn(1'b1),
		  .output_mode(1'b0),
		  .output_reset(0),
		  .output_sync(1'b0),
		  .pa_in_clock(-1),
		  .pa_in_clock_en(-1),
		  .pa_in_reset(-1),
		  .pa_out_clock(-1),
		  .pa_out_clock_en(-1),
		  .pa_out_reset(-1),
		  .pin_aliases(""),
		  .pin_mode("O"),
		  .por_state(4),
		  .sio_group_cnt(0),
		  .sio_hyst(1'b0),
		  .sio_ibuf(""),
		  .sio_info(2'b00),
		  .sio_obuf(""),
		  .sio_refsel(""),
		  .sio_vtrip(""),
		  .slew_rate(1'b0),
		  .spanning(0),
		  .use_annotation(1'b0),
		  .vtrip(2'b10),
		  .width(1))
		L_Servo
		 (.oe(tmpOE__L_Servo_net),
		  .y({Net_504}),
		  .fb({tmpFB_0__L_Servo_net[0:0]}),
		  .io({tmpIO_0__L_Servo_net[0:0]}),
		  .siovref(tmpSIOVREF__L_Servo_net),
		  .interrupt({tmpINTERRUPT_0__L_Servo_net[0:0]}),
		  .in_clock({1'b0}),
		  .in_clock_en({1'b1}),
		  .in_reset({1'b0}),
		  .out_clock({1'b0}),
		  .out_clock_en({1'b1}),
		  .out_reset({1'b0}));
	assign tmpOE__L_Servo_net = (`CYDEV_CHIP_MEMBER_USED == `CYDEV_CHIP_MEMBER_3A && `CYDEV_CHIP_REVISION_USED < `CYDEV_CHIP_REVISION_3A_ES3) ? ~{1'b1} : {1'b1};
	wire [0:0] tmpOE__R_Servo_net;
	wire [0:0] tmpFB_0__R_Servo_net;
	wire [0:0] tmpIO_0__R_Servo_net;
	wire [0:0] tmpINTERRUPT_0__R_Servo_net;
	electrical [0:0] tmpSIOVREF__R_Servo_net;
	cy_psoc3_pins_v1_10
		#(.id("b2308480-dcd7-4ee5-bbdc-18916ee367be"),
		  .drive_mode(3'b110),
		  .ibuf_enabled(1'b1),
		  .init_dr_st(1'b1),
		  .input_clk_en(0),
		  .input_sync(1'b1),
		  .input_sync_mode(1'b0),
		  .intr_mode(2'b00),
		  .invert_in_clock(0),
		  .invert_in_clock_en(0),
		  .invert_in_reset(0),
		  .invert_out_clock(0),
		  .invert_out_clock_en(0),
		  .invert_out_reset(0),
		  .io_voltage(""),
		  .layout_mode("CONTIGUOUS"),
		  .oe_conn(1'b0),
		  .oe_reset(0),
		  .oe_sync(1'b0),
		  .output_clk_en(0),
		  .output_clock_mode(1'b0),
		  .output_conn(1'b1),
		  .output_mode(1'b0),
		  .output_reset(0),
		  .output_sync(1'b0),
		  .pa_in_clock(-1),
		  .pa_in_clock_en(-1),
		  .pa_in_reset(-1),
		  .pa_out_clock(-1),
		  .pa_out_clock_en(-1),
		  .pa_out_reset(-1),
		  .pin_aliases(""),
		  .pin_mode("O"),
		  .por_state(4),
		  .sio_group_cnt(0),
		  .sio_hyst(1'b0),
		  .sio_ibuf(""),
		  .sio_info(2'b00),
		  .sio_obuf(""),
		  .sio_refsel(""),
		  .sio_vtrip(""),
		  .slew_rate(1'b0),
		  .spanning(0),
		  .use_annotation(1'b0),
		  .vtrip(2'b10),
		  .width(1))
		R_Servo
		 (.oe(tmpOE__R_Servo_net),
		  .y({Net_505}),
		  .fb({tmpFB_0__R_Servo_net[0:0]}),
		  .io({tmpIO_0__R_Servo_net[0:0]}),
		  .siovref(tmpSIOVREF__R_Servo_net),
		  .interrupt({tmpINTERRUPT_0__R_Servo_net[0:0]}),
		  .in_clock({1'b0}),
		  .in_clock_en({1'b1}),
		  .in_reset({1'b0}),
		  .out_clock({1'b0}),
		  .out_clock_en({1'b1}),
		  .out_reset({1'b0}));
	assign tmpOE__R_Servo_net = (`CYDEV_CHIP_MEMBER_USED == `CYDEV_CHIP_MEMBER_3A && `CYDEV_CHIP_REVISION_USED < `CYDEV_CHIP_REVISION_3A_ES3) ? ~{1'b1} : {1'b1};
    TCPWM_P4_v1_10_3 Wheels_1 (
        .stop(1'b0),
        .reload(1'b0),
        .start(1'b0),
        .count(1'b1),
        .capture(1'b0),
        .interrupt(Net_764),
        .ov(Net_765),
        .un(Net_766),
        .cc(Net_767),
        .line(Net_504),
        .line_n(Net_768),
        .clock(Net_496));
    defparam Wheels_1.PWMCountMode = 3;
    defparam Wheels_1.PWMReloadMode = 0;
    defparam Wheels_1.PWMReloadPresent = 0;
    defparam Wheels_1.PWMStartMode = 0;
    defparam Wheels_1.PWMStopMode = 0;
    defparam Wheels_1.PWMSwitchMode = 0;
    defparam Wheels_1.QuadIndexMode = 0;
    defparam Wheels_1.QuadPhiAMode = 3;
    defparam Wheels_1.QuadPhiBMode = 3;
    defparam Wheels_1.QuadStopMode = 0;
    defparam Wheels_1.TCCaptureMode = 0;
    defparam Wheels_1.TCCountMode = 3;
    defparam Wheels_1.TCReloadMode = 0;
    defparam Wheels_1.TCStartMode = 0;
    defparam Wheels_1.TCStopMode = 0;
	wire [0:0] tmpOE__GimbalP_net;
	wire [0:0] tmpFB_0__GimbalP_net;
	wire [0:0] tmpIO_0__GimbalP_net;
	wire [0:0] tmpINTERRUPT_0__GimbalP_net;
	electrical [0:0] tmpSIOVREF__GimbalP_net;
	cy_psoc3_pins_v1_10
		#(.id("8c1b8be6-e5e7-4bce-905a-4cfa28d02e70"),
		  .drive_mode(3'b110),
		  .ibuf_enabled(1'b1),
		  .init_dr_st(1'b1),
		  .input_clk_en(0),
		  .input_sync(1'b1),
		  .input_sync_mode(1'b0),
		  .intr_mode(2'b00),
		  .invert_in_clock(0),
		  .invert_in_clock_en(0),
		  .invert_in_reset(0),
		  .invert_out_clock(0),
		  .invert_out_clock_en(0),
		  .invert_out_reset(0),
		  .io_voltage(""),
		  .layout_mode("CONTIGUOUS"),
		  .oe_conn(1'b0),
		  .oe_reset(0),
		  .oe_sync(1'b0),
		  .output_clk_en(0),
		  .output_clock_mode(1'b0),
		  .output_conn(1'b1),
		  .output_mode(1'b0),
		  .output_reset(0),
		  .output_sync(1'b0),
		  .pa_in_clock(-1),
		  .pa_in_clock_en(-1),
		  .pa_in_reset(-1),
		  .pa_out_clock(-1),
		  .pa_out_clock_en(-1),
		  .pa_out_reset(-1),
		  .pin_aliases(""),
		  .pin_mode("O"),
		  .por_state(4),
		  .sio_group_cnt(0),
		  .sio_hyst(1'b0),
		  .sio_ibuf(""),
		  .sio_info(2'b00),
		  .sio_obuf(""),
		  .sio_refsel(""),
		  .sio_vtrip(""),
		  .slew_rate(1'b0),
		  .spanning(0),
		  .use_annotation(1'b0),
		  .vtrip(2'b10),
		  .width(1))
		GimbalP
		 (.oe(tmpOE__GimbalP_net),
		  .y({Net_518}),
		  .fb({tmpFB_0__GimbalP_net[0:0]}),
		  .io({tmpIO_0__GimbalP_net[0:0]}),
		  .siovref(tmpSIOVREF__GimbalP_net),
		  .interrupt({tmpINTERRUPT_0__GimbalP_net[0:0]}),
		  .in_clock({1'b0}),
		  .in_clock_en({1'b1}),
		  .in_reset({1'b0}),
		  .out_clock({1'b0}),
		  .out_clock_en({1'b1}),
		  .out_reset({1'b0}));
	assign tmpOE__GimbalP_net = (`CYDEV_CHIP_MEMBER_USED == `CYDEV_CHIP_MEMBER_3A && `CYDEV_CHIP_REVISION_USED < `CYDEV_CHIP_REVISION_3A_ES3) ? ~{1'b1} : {1'b1};
	wire [0:0] tmpOE__GimbalT_net;
	wire [0:0] tmpFB_0__GimbalT_net;
	wire [0:0] tmpIO_0__GimbalT_net;
	wire [0:0] tmpINTERRUPT_0__GimbalT_net;
	electrical [0:0] tmpSIOVREF__GimbalT_net;
	cy_psoc3_pins_v1_10
		#(.id("c2106cdb-687e-44ec-9e29-5bc0f817d259"),
		  .drive_mode(3'b110),
		  .ibuf_enabled(1'b1),
		  .init_dr_st(1'b1),
		  .input_clk_en(0),
		  .input_sync(1'b1),
		  .input_sync_mode(1'b0),
		  .intr_mode(2'b00),
		  .invert_in_clock(0),
		  .invert_in_clock_en(0),
		  .invert_in_reset(0),
		  .invert_out_clock(0),
		  .invert_out_clock_en(0),
		  .invert_out_reset(0),
		  .io_voltage(""),
		  .layout_mode("CONTIGUOUS"),
		  .oe_conn(1'b0),
		  .oe_reset(0),
		  .oe_sync(1'b0),
		  .output_clk_en(0),
		  .output_clock_mode(1'b0),
		  .output_conn(1'b1),
		  .output_mode(1'b0),
		  .output_reset(0),
		  .output_sync(1'b0),
		  .pa_in_clock(-1),
		  .pa_in_clock_en(-1),
		  .pa_in_reset(-1),
		  .pa_out_clock(-1),
		  .pa_out_clock_en(-1),
		  .pa_out_reset(-1),
		  .pin_aliases(""),
		  .pin_mode("O"),
		  .por_state(4),
		  .sio_group_cnt(0),
		  .sio_hyst(1'b0),
		  .sio_ibuf(""),
		  .sio_info(2'b00),
		  .sio_obuf(""),
		  .sio_refsel(""),
		  .sio_vtrip(""),
		  .slew_rate(1'b0),
		  .spanning(0),
		  .use_annotation(1'b0),
		  .vtrip(2'b10),
		  .width(1))
		GimbalT
		 (.oe(tmpOE__GimbalT_net),
		  .y({Net_519}),
		  .fb({tmpFB_0__GimbalT_net[0:0]}),
		  .io({tmpIO_0__GimbalT_net[0:0]}),
		  .siovref(tmpSIOVREF__GimbalT_net),
		  .interrupt({tmpINTERRUPT_0__GimbalT_net[0:0]}),
		  .in_clock({1'b0}),
		  .in_clock_en({1'b1}),
		  .in_reset({1'b0}),
		  .out_clock({1'b0}),
		  .out_clock_en({1'b1}),
		  .out_reset({1'b0}));
	assign tmpOE__GimbalT_net = (`CYDEV_CHIP_MEMBER_USED == `CYDEV_CHIP_MEMBER_3A && `CYDEV_CHIP_REVISION_USED < `CYDEV_CHIP_REVISION_3A_ES3) ? ~{1'b1} : {1'b1};
    SPI_Master_v2_40_4 SPIM (
        .mosi(Net_675),
        .sclk(Net_676),
        .ss(Net_747),
        .miso(Net_678),
        .clock(1'b0),
        .reset(1'b0),
        .rx_interrupt(Net_681),
        .sdat(Net_863),
        .tx_interrupt(Net_864));
    defparam SPIM.BidirectMode = 0;
    defparam SPIM.HighSpeedMode = 0;
    defparam SPIM.NumberOfDataBits = 8;
    defparam SPIM.ShiftDir = 0;
	cy_isr_v1_0
		#(.int_type(2'b10))
		ISRSPI
		 (.int_signal(Net_872));
    SCB_P4_v1_20_5 GPS_UART (
        .sclk(Net_756),
        .interrupt(Net_701),
        .clock(1'b0));
	cy_isr_v1_0
		#(.int_type(2'b10))
		ISR_UART_2
		 (.int_signal(Net_701));
	wire [0:0] tmpOE__MISO_net;
	wire [0:0] tmpIO_0__MISO_net;
	wire [0:0] tmpINTERRUPT_0__MISO_net;
	electrical [0:0] tmpSIOVREF__MISO_net;
	cy_psoc3_pins_v1_10
		#(.id("552faf00-97dc-47bf-ad14-15574b2c6e9b"),
		  .drive_mode(3'b001),
		  .ibuf_enabled(1'b1),
		  .init_dr_st(1'b0),
		  .input_clk_en(0),
		  .input_sync(1'b1),
		  .input_sync_mode(1'b0),
		  .intr_mode(2'b00),
		  .invert_in_clock(0),
		  .invert_in_clock_en(0),
		  .invert_in_reset(0),
		  .invert_out_clock(0),
		  .invert_out_clock_en(0),
		  .invert_out_reset(0),
		  .io_voltage(""),
		  .layout_mode("CONTIGUOUS"),
		  .oe_conn(1'b0),
		  .oe_reset(0),
		  .oe_sync(1'b0),
		  .output_clk_en(0),
		  .output_clock_mode(1'b0),
		  .output_conn(1'b0),
		  .output_mode(1'b0),
		  .output_reset(0),
		  .output_sync(1'b0),
		  .pa_in_clock(-1),
		  .pa_in_clock_en(-1),
		  .pa_in_reset(-1),
		  .pa_out_clock(-1),
		  .pa_out_clock_en(-1),
		  .pa_out_reset(-1),
		  .pin_aliases(""),
		  .pin_mode("I"),
		  .por_state(4),
		  .sio_group_cnt(0),
		  .sio_hyst(1'b0),
		  .sio_ibuf(""),
		  .sio_info(2'b00),
		  .sio_obuf(""),
		  .sio_refsel(""),
		  .sio_vtrip(""),
		  .slew_rate(1'b0),
		  .spanning(0),
		  .use_annotation(1'b0),
		  .vtrip(2'b00),
		  .width(1))
		MISO
		 (.oe(tmpOE__MISO_net),
		  .y({1'b0}),
		  .fb({Net_678}),
		  .io({tmpIO_0__MISO_net[0:0]}),
		  .siovref(tmpSIOVREF__MISO_net),
		  .interrupt({tmpINTERRUPT_0__MISO_net[0:0]}),
		  .in_clock({1'b0}),
		  .in_clock_en({1'b1}),
		  .in_reset({1'b0}),
		  .out_clock({1'b0}),
		  .out_clock_en({1'b1}),
		  .out_reset({1'b0}));
	assign tmpOE__MISO_net = (`CYDEV_CHIP_MEMBER_USED == `CYDEV_CHIP_MEMBER_3A && `CYDEV_CHIP_REVISION_USED < `CYDEV_CHIP_REVISION_3A_ES3) ? ~{1'b1} : {1'b1};
	wire [0:0] tmpOE__MOSI_net;
	wire [0:0] tmpFB_0__MOSI_net;
	wire [0:0] tmpIO_0__MOSI_net;
	wire [0:0] tmpINTERRUPT_0__MOSI_net;
	electrical [0:0] tmpSIOVREF__MOSI_net;
	cy_psoc3_pins_v1_10
		#(.id("0e0c9380-6965-4440-8709-ce08a91e474c"),
		  .drive_mode(3'b110),
		  .ibuf_enabled(1'b1),
		  .init_dr_st(1'b1),
		  .input_clk_en(0),
		  .input_sync(1'b1),
		  .input_sync_mode(1'b0),
		  .intr_mode(2'b00),
		  .invert_in_clock(0),
		  .invert_in_clock_en(0),
		  .invert_in_reset(0),
		  .invert_out_clock(0),
		  .invert_out_clock_en(0),
		  .invert_out_reset(0),
		  .io_voltage(""),
		  .layout_mode("CONTIGUOUS"),
		  .oe_conn(1'b0),
		  .oe_reset(0),
		  .oe_sync(1'b0),
		  .output_clk_en(0),
		  .output_clock_mode(1'b0),
		  .output_conn(1'b1),
		  .output_mode(1'b0),
		  .output_reset(0),
		  .output_sync(1'b0),
		  .pa_in_clock(-1),
		  .pa_in_clock_en(-1),
		  .pa_in_reset(-1),
		  .pa_out_clock(-1),
		  .pa_out_clock_en(-1),
		  .pa_out_reset(-1),
		  .pin_aliases(""),
		  .pin_mode("O"),
		  .por_state(4),
		  .sio_group_cnt(0),
		  .sio_hyst(1'b0),
		  .sio_ibuf(""),
		  .sio_info(2'b00),
		  .sio_obuf(""),
		  .sio_refsel(""),
		  .sio_vtrip(""),
		  .slew_rate(1'b0),
		  .spanning(0),
		  .use_annotation(1'b0),
		  .vtrip(2'b10),
		  .width(1))
		MOSI
		 (.oe(tmpOE__MOSI_net),
		  .y({Net_675}),
		  .fb({tmpFB_0__MOSI_net[0:0]}),
		  .io({tmpIO_0__MOSI_net[0:0]}),
		  .siovref(tmpSIOVREF__MOSI_net),
		  .interrupt({tmpINTERRUPT_0__MOSI_net[0:0]}),
		  .in_clock({1'b0}),
		  .in_clock_en({1'b1}),
		  .in_reset({1'b0}),
		  .out_clock({1'b0}),
		  .out_clock_en({1'b1}),
		  .out_reset({1'b0}));
	assign tmpOE__MOSI_net = (`CYDEV_CHIP_MEMBER_USED == `CYDEV_CHIP_MEMBER_3A && `CYDEV_CHIP_REVISION_USED < `CYDEV_CHIP_REVISION_3A_ES3) ? ~{1'b1} : {1'b1};
	wire [0:0] tmpOE__SCLK_net;
	wire [0:0] tmpFB_0__SCLK_net;
	wire [0:0] tmpIO_0__SCLK_net;
	wire [0:0] tmpINTERRUPT_0__SCLK_net;
	electrical [0:0] tmpSIOVREF__SCLK_net;
	cy_psoc3_pins_v1_10
		#(.id("7f71d314-4523-45d3-b07e-62700396d125"),
		  .drive_mode(3'b110),
		  .ibuf_enabled(1'b1),
		  .init_dr_st(1'b1),
		  .input_clk_en(0),
		  .input_sync(1'b1),
		  .input_sync_mode(1'b0),
		  .intr_mode(2'b00),
		  .invert_in_clock(0),
		  .invert_in_clock_en(0),
		  .invert_in_reset(0),
		  .invert_out_clock(0),
		  .invert_out_clock_en(0),
		  .invert_out_reset(0),
		  .io_voltage(""),
		  .layout_mode("CONTIGUOUS"),
		  .oe_conn(1'b0),
		  .oe_reset(0),
		  .oe_sync(1'b0),
		  .output_clk_en(0),
		  .output_clock_mode(1'b0),
		  .output_conn(1'b1),
		  .output_mode(1'b0),
		  .output_reset(0),
		  .output_sync(1'b0),
		  .pa_in_clock(-1),
		  .pa_in_clock_en(-1),
		  .pa_in_reset(-1),
		  .pa_out_clock(-1),
		  .pa_out_clock_en(-1),
		  .pa_out_reset(-1),
		  .pin_aliases(""),
		  .pin_mode("O"),
		  .por_state(4),
		  .sio_group_cnt(0),
		  .sio_hyst(1'b0),
		  .sio_ibuf(""),
		  .sio_info(2'b00),
		  .sio_obuf(""),
		  .sio_refsel(""),
		  .sio_vtrip(""),
		  .slew_rate(1'b0),
		  .spanning(0),
		  .use_annotation(1'b0),
		  .vtrip(2'b10),
		  .width(1))
		SCLK
		 (.oe(tmpOE__SCLK_net),
		  .y({Net_676}),
		  .fb({tmpFB_0__SCLK_net[0:0]}),
		  .io({tmpIO_0__SCLK_net[0:0]}),
		  .siovref(tmpSIOVREF__SCLK_net),
		  .interrupt({tmpINTERRUPT_0__SCLK_net[0:0]}),
		  .in_clock({1'b0}),
		  .in_clock_en({1'b1}),
		  .in_reset({1'b0}),
		  .out_clock({1'b0}),
		  .out_clock_en({1'b1}),
		  .out_reset({1'b0}));
	assign tmpOE__SCLK_net = (`CYDEV_CHIP_MEMBER_USED == `CYDEV_CHIP_MEMBER_3A && `CYDEV_CHIP_REVISION_USED < `CYDEV_CHIP_REVISION_3A_ES3) ? ~{1'b1} : {1'b1};
    TCPWM_P4_v1_10_6 Wheels_2 (
        .stop(1'b0),
        .reload(1'b0),
        .start(1'b0),
        .count(1'b1),
        .capture(1'b0),
        .interrupt(Net_774),
        .ov(Net_775),
        .un(Net_776),
        .cc(Net_777),
        .line(Net_505),
        .line_n(Net_778),
        .clock(Net_496));
    defparam Wheels_2.PWMCountMode = 3;
    defparam Wheels_2.PWMReloadMode = 0;
    defparam Wheels_2.PWMReloadPresent = 0;
    defparam Wheels_2.PWMStartMode = 0;
    defparam Wheels_2.PWMStopMode = 0;
    defparam Wheels_2.PWMSwitchMode = 0;
    defparam Wheels_2.QuadIndexMode = 0;
    defparam Wheels_2.QuadPhiAMode = 3;
    defparam Wheels_2.QuadPhiBMode = 3;
    defparam Wheels_2.QuadStopMode = 0;
    defparam Wheels_2.TCCaptureMode = 0;
    defparam Wheels_2.TCCountMode = 3;
    defparam Wheels_2.TCReloadMode = 0;
    defparam Wheels_2.TCStartMode = 0;
    defparam Wheels_2.TCStopMode = 0;
    CyControlReg_v1_70 VidMux (
        .control_1(Net_820),
        .control_2(Net_821),
        .control_3(Net_822),
        .control_0(Net_823),
        .control_4(Net_824),
        .control_5(Net_825),
        .control_6(Net_826),
        .control_7(Net_827),
        .clock(1'b0),
        .reset(1'b0));
    defparam VidMux.Bit0Mode = 0;
    defparam VidMux.Bit1Mode = 0;
    defparam VidMux.Bit2Mode = 0;
    defparam VidMux.Bit3Mode = 0;
    defparam VidMux.Bit4Mode = 0;
    defparam VidMux.Bit5Mode = 0;
    defparam VidMux.Bit6Mode = 0;
    defparam VidMux.Bit7Mode = 0;
    defparam VidMux.BitValue = 0;
    defparam VidMux.BusDisplay = 0;
    defparam VidMux.ExtrReset = 0;
    defparam VidMux.NumOutputs = 3;
	wire [0:0] tmpOE__WIZ_RST_net;
	wire [0:0] tmpFB_0__WIZ_RST_net;
	wire [0:0] tmpIO_0__WIZ_RST_net;
	wire [0:0] tmpINTERRUPT_0__WIZ_RST_net;
	electrical [0:0] tmpSIOVREF__WIZ_RST_net;
	cy_psoc3_pins_v1_10
		#(.id("0685bd1c-6e36-4e2b-bb80-086b6cfb9431"),
		  .drive_mode(3'b110),
		  .ibuf_enabled(1'b1),
		  .init_dr_st(1'b0),
		  .input_clk_en(0),
		  .input_sync(1'b1),
		  .input_sync_mode(1'b0),
		  .intr_mode(2'b00),
		  .invert_in_clock(0),
		  .invert_in_clock_en(0),
		  .invert_in_reset(0),
		  .invert_out_clock(0),
		  .invert_out_clock_en(0),
		  .invert_out_reset(0),
		  .io_voltage(""),
		  .layout_mode("CONTIGUOUS"),
		  .oe_conn(1'b0),
		  .oe_reset(0),
		  .oe_sync(1'b0),
		  .output_clk_en(0),
		  .output_clock_mode(1'b0),
		  .output_conn(1'b0),
		  .output_mode(1'b0),
		  .output_reset(0),
		  .output_sync(1'b0),
		  .pa_in_clock(-1),
		  .pa_in_clock_en(-1),
		  .pa_in_reset(-1),
		  .pa_out_clock(-1),
		  .pa_out_clock_en(-1),
		  .pa_out_reset(-1),
		  .pin_aliases(""),
		  .pin_mode("O"),
		  .por_state(4),
		  .sio_group_cnt(0),
		  .sio_hyst(1'b0),
		  .sio_ibuf(""),
		  .sio_info(2'b00),
		  .sio_obuf(""),
		  .sio_refsel(""),
		  .sio_vtrip(""),
		  .slew_rate(1'b0),
		  .spanning(0),
		  .use_annotation(1'b0),
		  .vtrip(2'b10),
		  .width(1))
		WIZ_RST
		 (.oe(tmpOE__WIZ_RST_net),
		  .y({1'b0}),
		  .fb({tmpFB_0__WIZ_RST_net[0:0]}),
		  .io({tmpIO_0__WIZ_RST_net[0:0]}),
		  .siovref(tmpSIOVREF__WIZ_RST_net),
		  .interrupt({tmpINTERRUPT_0__WIZ_RST_net[0:0]}),
		  .in_clock({1'b0}),
		  .in_clock_en({1'b1}),
		  .in_reset({1'b0}),
		  .out_clock({1'b0}),
		  .out_clock_en({1'b1}),
		  .out_reset({1'b0}));
	assign tmpOE__WIZ_RST_net = (`CYDEV_CHIP_MEMBER_USED == `CYDEV_CHIP_MEMBER_3A && `CYDEV_CHIP_REVISION_USED < `CYDEV_CHIP_REVISION_3A_ES3) ? ~{1'b1} : {1'b1};
	wire [0:0] tmpOE__WIZ_RDY_net;
	wire [0:0] tmpFB_0__WIZ_RDY_net;
	wire [0:0] tmpIO_0__WIZ_RDY_net;
	wire [0:0] tmpINTERRUPT_0__WIZ_RDY_net;
	electrical [0:0] tmpSIOVREF__WIZ_RDY_net;
	cy_psoc3_pins_v1_10
		#(.id("7f151c7d-1f6c-461e-9c68-16dcffc8e4d8"),
		  .drive_mode(3'b001),
		  .ibuf_enabled(1'b1),
		  .init_dr_st(1'b0),
		  .input_clk_en(0),
		  .input_sync(1'b1),
		  .input_sync_mode(1'b0),
		  .intr_mode(2'b00),
		  .invert_in_clock(0),
		  .invert_in_clock_en(0),
		  .invert_in_reset(0),
		  .invert_out_clock(0),
		  .invert_out_clock_en(0),
		  .invert_out_reset(0),
		  .io_voltage(""),
		  .layout_mode("CONTIGUOUS"),
		  .oe_conn(1'b0),
		  .oe_reset(0),
		  .oe_sync(1'b0),
		  .output_clk_en(0),
		  .output_clock_mode(1'b0),
		  .output_conn(1'b0),
		  .output_mode(1'b0),
		  .output_reset(0),
		  .output_sync(1'b0),
		  .pa_in_clock(-1),
		  .pa_in_clock_en(-1),
		  .pa_in_reset(-1),
		  .pa_out_clock(-1),
		  .pa_out_clock_en(-1),
		  .pa_out_reset(-1),
		  .pin_aliases(""),
		  .pin_mode("I"),
		  .por_state(4),
		  .sio_group_cnt(0),
		  .sio_hyst(1'b0),
		  .sio_ibuf(""),
		  .sio_info(2'b00),
		  .sio_obuf(""),
		  .sio_refsel(""),
		  .sio_vtrip(""),
		  .slew_rate(1'b0),
		  .spanning(0),
		  .use_annotation(1'b0),
		  .vtrip(2'b00),
		  .width(1))
		WIZ_RDY
		 (.oe(tmpOE__WIZ_RDY_net),
		  .y({1'b0}),
		  .fb({tmpFB_0__WIZ_RDY_net[0:0]}),
		  .io({tmpIO_0__WIZ_RDY_net[0:0]}),
		  .siovref(tmpSIOVREF__WIZ_RDY_net),
		  .interrupt({tmpINTERRUPT_0__WIZ_RDY_net[0:0]}),
		  .in_clock({1'b0}),
		  .in_clock_en({1'b1}),
		  .in_reset({1'b0}),
		  .out_clock({1'b0}),
		  .out_clock_en({1'b1}),
		  .out_reset({1'b0}));
	assign tmpOE__WIZ_RDY_net = (`CYDEV_CHIP_MEMBER_USED == `CYDEV_CHIP_MEMBER_3A && `CYDEV_CHIP_REVISION_USED < `CYDEV_CHIP_REVISION_3A_ES3) ? ~{1'b1} : {1'b1};
	wire [0:0] tmpOE__WIZ_INT_net;
	wire [0:0] tmpIO_0__WIZ_INT_net;
	wire [0:0] tmpINTERRUPT_0__WIZ_INT_net;
	electrical [0:0] tmpSIOVREF__WIZ_INT_net;
	cy_psoc3_pins_v1_10
		#(.id("f7e52380-b69e-4bcf-b0e7-b82bec578576"),
		  .drive_mode(3'b001),
		  .ibuf_enabled(1'b1),
		  .init_dr_st(1'b0),
		  .input_clk_en(0),
		  .input_sync(1'b1),
		  .input_sync_mode(1'b0),
		  .intr_mode(2'b00),
		  .invert_in_clock(0),
		  .invert_in_clock_en(0),
		  .invert_in_reset(0),
		  .invert_out_clock(0),
		  .invert_out_clock_en(0),
		  .invert_out_reset(0),
		  .io_voltage(""),
		  .layout_mode("CONTIGUOUS"),
		  .oe_conn(1'b0),
		  .oe_reset(0),
		  .oe_sync(1'b0),
		  .output_clk_en(0),
		  .output_clock_mode(1'b0),
		  .output_conn(1'b0),
		  .output_mode(1'b0),
		  .output_reset(0),
		  .output_sync(1'b0),
		  .pa_in_clock(-1),
		  .pa_in_clock_en(-1),
		  .pa_in_reset(-1),
		  .pa_out_clock(-1),
		  .pa_out_clock_en(-1),
		  .pa_out_reset(-1),
		  .pin_aliases(""),
		  .pin_mode("I"),
		  .por_state(4),
		  .sio_group_cnt(0),
		  .sio_hyst(1'b0),
		  .sio_ibuf(""),
		  .sio_info(2'b00),
		  .sio_obuf(""),
		  .sio_refsel(""),
		  .sio_vtrip(""),
		  .slew_rate(1'b0),
		  .spanning(0),
		  .use_annotation(1'b0),
		  .vtrip(2'b00),
		  .width(1))
		WIZ_INT
		 (.oe(tmpOE__WIZ_INT_net),
		  .y({1'b0}),
		  .fb({Net_872}),
		  .io({tmpIO_0__WIZ_INT_net[0:0]}),
		  .siovref(tmpSIOVREF__WIZ_INT_net),
		  .interrupt({tmpINTERRUPT_0__WIZ_INT_net[0:0]}),
		  .in_clock({1'b0}),
		  .in_clock_en({1'b1}),
		  .in_reset({1'b0}),
		  .out_clock({1'b0}),
		  .out_clock_en({1'b1}),
		  .out_reset({1'b0}));
	assign tmpOE__WIZ_INT_net = (`CYDEV_CHIP_MEMBER_USED == `CYDEV_CHIP_MEMBER_3A && `CYDEV_CHIP_REVISION_USED < `CYDEV_CHIP_REVISION_3A_ES3) ? ~{1'b1} : {1'b1};
	wire [0:0] tmpOE__WIZ_SS_net;
	wire [0:0] tmpFB_0__WIZ_SS_net;
	wire [0:0] tmpIO_0__WIZ_SS_net;
	wire [0:0] tmpINTERRUPT_0__WIZ_SS_net;
	electrical [0:0] tmpSIOVREF__WIZ_SS_net;
	cy_psoc3_pins_v1_10
		#(.id("c5824ab3-47bc-41f7-b4a6-1015f51c5578"),
		  .drive_mode(3'b110),
		  .ibuf_enabled(1'b1),
		  .init_dr_st(1'b1),
		  .input_clk_en(0),
		  .input_sync(1'b1),
		  .input_sync_mode(1'b0),
		  .intr_mode(2'b00),
		  .invert_in_clock(0),
		  .invert_in_clock_en(0),
		  .invert_in_reset(0),
		  .invert_out_clock(0),
		  .invert_out_clock_en(0),
		  .invert_out_reset(0),
		  .io_voltage(""),
		  .layout_mode("CONTIGUOUS"),
		  .oe_conn(1'b0),
		  .oe_reset(0),
		  .oe_sync(1'b0),
		  .output_clk_en(0),
		  .output_clock_mode(1'b0),
		  .output_conn(1'b0),
		  .output_mode(1'b0),
		  .output_reset(0),
		  .output_sync(1'b0),
		  .pa_in_clock(-1),
		  .pa_in_clock_en(-1),
		  .pa_in_reset(-1),
		  .pa_out_clock(-1),
		  .pa_out_clock_en(-1),
		  .pa_out_reset(-1),
		  .pin_aliases(""),
		  .pin_mode("O"),
		  .por_state(4),
		  .sio_group_cnt(0),
		  .sio_hyst(1'b0),
		  .sio_ibuf(""),
		  .sio_info(2'b00),
		  .sio_obuf(""),
		  .sio_refsel(""),
		  .sio_vtrip(""),
		  .slew_rate(1'b0),
		  .spanning(0),
		  .use_annotation(1'b0),
		  .vtrip(2'b10),
		  .width(1))
		WIZ_SS
		 (.oe(tmpOE__WIZ_SS_net),
		  .y({1'b0}),
		  .fb({tmpFB_0__WIZ_SS_net[0:0]}),
		  .io({tmpIO_0__WIZ_SS_net[0:0]}),
		  .siovref(tmpSIOVREF__WIZ_SS_net),
		  .interrupt({tmpINTERRUPT_0__WIZ_SS_net[0:0]}),
		  .in_clock({1'b0}),
		  .in_clock_en({1'b1}),
		  .in_reset({1'b0}),
		  .out_clock({1'b0}),
		  .out_clock_en({1'b1}),
		  .out_reset({1'b0}));
	assign tmpOE__WIZ_SS_net = (`CYDEV_CHIP_MEMBER_USED == `CYDEV_CHIP_MEMBER_3A && `CYDEV_CHIP_REVISION_USED < `CYDEV_CHIP_REVISION_3A_ES3) ? ~{1'b1} : {1'b1};
endmodule