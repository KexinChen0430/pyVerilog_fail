module can be reset
            init_flag <= 1;
        end
    end
endmodule