module header
	// Internal signals
	// Generated Signal List
	// End of Generated Signal List
	// %COMPILER_OPTS%
	// Generated Signal Assignments
udc: Verilog BODY HOOK inst_bc1_i
	// Generated Instances and Port Mappings
endmodule