module's unterminated outputs)
   wire o_B_internal = 1'h0;
   wire o_B_outsideo = 1'h0;
   // End of automatics
endmodule