module FFT_IFFT_IP_CORE (
  clk, start, unload, fwd_inv, fwd_inv_we, rfd, busy, edone, done, dv, xn_re, xn_im, xn_index, xk_index, xk_re, xk_im
)/* synthesis syn_black_box syn_noprune=1 */;
  input clk;
  input start;
  input unload;
  input fwd_inv;
  input fwd_inv_we;
  output rfd;
  output busy;
  output edone;
  output done;
  output dv;
  input [8 : 0] xn_re;
  input [8 : 0] xn_im;
  output [8 : 0] xn_index;
  output [8 : 0] xk_index;
  output [18 : 0] xk_re;
  output [18 : 0] xk_im;
  // synthesis translate_off
  wire \NlwRenamedSig_OI_U0/i_synth/non_floating_point.arch_c.xfft_inst/control/cntrl/loading_state/ORS ;
  wire \NlwRenamedSig_OI_U0/i_synth/non_floating_point.arch_c.xfft_inst/control/cntrl/processing_state/ORS ;
  wire \U0/i_synth/non_floating_point.arch_c.xfft_inst/control/cntrl/done_pr_d_1 ;
  wire sig00000001;
  wire sig00000002;
  wire sig00000003;
  wire sig00000004;
  wire sig00000005;
  wire sig00000006;
  wire sig00000007;
  wire sig00000008;
  wire sig00000009;
  wire sig0000000a;
  wire sig0000000b;
  wire sig0000000c;
  wire sig0000000d;
  wire sig0000000e;
  wire sig0000000f;
  wire sig00000010;
  wire sig00000011;
  wire sig00000012;
  wire sig00000013;
  wire sig00000014;
  wire sig00000015;
  wire sig00000016;
  wire sig00000017;
  wire sig00000018;
  wire sig00000019;
  wire sig0000001a;
  wire sig0000001b;
  wire sig0000001c;
  wire sig0000001d;
  wire sig0000001e;
  wire sig0000001f;
  wire sig00000020;
  wire sig00000021;
  wire sig00000022;
  wire sig00000023;
  wire sig00000024;
  wire sig00000025;
  wire sig00000026;
  wire sig00000027;
  wire sig00000028;
  wire sig00000029;
  wire sig0000002a;
  wire sig0000002b;
  wire sig0000002c;
  wire sig0000002d;
  wire sig0000002e;
  wire sig0000002f;
  wire sig00000030;
  wire sig00000031;
  wire sig00000032;
  wire sig00000033;
  wire sig00000034;
  wire sig00000035;
  wire sig00000036;
  wire sig00000037;
  wire sig00000038;
  wire sig00000039;
  wire sig0000003a;
  wire sig0000003b;
  wire sig0000003c;
  wire sig0000003d;
  wire sig0000003e;
  wire sig0000003f;
  wire sig00000040;
  wire sig00000041;
  wire sig00000042;
  wire sig00000043;
  wire sig00000044;
  wire sig00000045;
  wire sig00000046;
  wire sig00000047;
  wire sig00000048;
  wire sig00000049;
  wire sig0000004a;
  wire sig0000004b;
  wire sig0000004c;
  wire sig0000004d;
  wire sig0000004e;
  wire sig0000004f;
  wire sig00000050;
  wire sig00000051;
  wire sig00000052;
  wire sig00000053;
  wire sig00000054;
  wire sig00000055;
  wire sig00000056;
  wire sig00000057;
  wire sig00000058;
  wire sig00000059;
  wire sig0000005a;
  wire sig0000005b;
  wire sig0000005c;
  wire sig0000005d;
  wire sig0000005e;
  wire sig0000005f;
  wire sig00000060;
  wire sig00000061;
  wire sig00000062;
  wire sig00000063;
  wire sig00000064;
  wire sig00000065;
  wire sig00000066;
  wire sig00000067;
  wire sig00000068;
  wire sig00000069;
  wire sig0000006a;
  wire sig0000006b;
  wire sig0000006c;
  wire sig0000006d;
  wire sig0000006e;
  wire sig0000006f;
  wire sig00000070;
  wire sig00000071;
  wire sig00000072;
  wire sig00000073;
  wire sig00000074;
  wire sig00000075;
  wire sig00000076;
  wire sig00000077;
  wire sig00000078;
  wire sig00000079;
  wire sig0000007a;
  wire sig0000007b;
  wire sig0000007c;
  wire sig0000007d;
  wire sig0000007e;
  wire sig0000007f;
  wire sig00000080;
  wire sig00000081;
  wire sig00000082;
  wire sig00000083;
  wire sig00000084;
  wire sig00000085;
  wire sig00000086;
  wire sig00000087;
  wire sig00000088;
  wire sig00000089;
  wire sig0000008a;
  wire sig0000008b;
  wire sig0000008c;
  wire sig0000008d;
  wire sig0000008e;
  wire sig0000008f;
  wire sig00000090;
  wire sig00000091;
  wire sig00000092;
  wire sig00000093;
  wire sig00000094;
  wire sig00000095;
  wire sig00000096;
  wire sig00000097;
  wire sig00000098;
  wire sig00000099;
  wire sig0000009a;
  wire sig0000009b;
  wire sig0000009c;
  wire sig0000009d;
  wire sig0000009e;
  wire sig0000009f;
  wire sig000000a0;
  wire sig000000a1;
  wire sig000000a2;
  wire sig000000a3;
  wire sig000000a4;
  wire sig000000a5;
  wire sig000000a6;
  wire sig000000a7;
  wire sig000000a8;
  wire sig000000a9;
  wire sig000000aa;
  wire sig000000ab;
  wire sig000000ac;
  wire sig000000ad;
  wire sig000000ae;
  wire sig000000af;
  wire sig000000b0;
  wire sig000000b1;
  wire sig000000b2;
  wire sig000000b3;
  wire sig000000b4;
  wire sig000000b5;
  wire sig000000b6;
  wire sig000000b7;
  wire sig000000b8;
  wire sig000000b9;
  wire sig000000ba;
  wire sig000000bb;
  wire sig000000bc;
  wire sig000000bd;
  wire sig000000be;
  wire sig000000bf;
  wire sig000000c0;
  wire sig000000c1;
  wire sig000000c2;
  wire sig000000c3;
  wire sig000000c4;
  wire sig000000c5;
  wire sig000000c6;
  wire sig000000c7;
  wire sig000000c8;
  wire sig000000c9;
  wire sig000000ca;
  wire sig000000cb;
  wire sig000000cc;
  wire sig000000cd;
  wire sig000000ce;
  wire sig000000cf;
  wire sig000000d0;
  wire sig000000d1;
  wire sig000000d2;
  wire sig000000d3;
  wire sig000000d4;
  wire sig000000d5;
  wire sig000000d6;
  wire sig000000d7;
  wire sig000000d8;
  wire sig000000d9;
  wire sig000000da;
  wire sig000000db;
  wire sig000000dc;
  wire sig000000dd;
  wire sig000000de;
  wire sig000000df;
  wire sig000000e0;
  wire sig000000e1;
  wire sig000000e2;
  wire sig000000e3;
  wire sig000000e4;
  wire sig000000e5;
  wire sig000000e6;
  wire sig000000e7;
  wire sig000000e8;
  wire sig000000e9;
  wire sig000000ea;
  wire sig000000eb;
  wire sig000000ec;
  wire sig000000ed;
  wire sig000000ee;
  wire sig000000ef;
  wire sig000000f0;
  wire sig000000f1;
  wire sig000000f2;
  wire sig000000f3;
  wire sig000000f4;
  wire sig000000f5;
  wire sig000000f6;
  wire sig000000f7;
  wire sig000000f8;
  wire sig000000f9;
  wire sig000000fa;
  wire sig000000fb;
  wire sig000000fc;
  wire sig000000fd;
  wire sig000000fe;
  wire sig000000ff;
  wire sig00000100;
  wire sig00000101;
  wire sig00000102;
  wire sig00000103;
  wire sig00000104;
  wire sig00000105;
  wire sig00000106;
  wire sig00000107;
  wire sig00000108;
  wire sig00000109;
  wire sig0000010a;
  wire sig0000010b;
  wire sig0000010c;
  wire sig0000010d;
  wire sig0000010e;
  wire sig0000010f;
  wire sig00000110;
  wire sig00000111;
  wire sig00000112;
  wire sig00000113;
  wire sig00000114;
  wire sig00000115;
  wire sig00000116;
  wire sig00000117;
  wire sig00000118;
  wire sig00000119;
  wire sig0000011a;
  wire sig0000011b;
  wire sig0000011c;
  wire sig0000011d;
  wire sig0000011e;
  wire sig0000011f;
  wire sig00000120;
  wire sig00000121;
  wire sig00000122;
  wire sig00000123;
  wire sig00000124;
  wire sig00000125;
  wire sig00000126;
  wire sig00000127;
  wire sig00000128;
  wire sig00000129;
  wire sig0000012a;
  wire sig0000012b;
  wire sig0000012c;
  wire sig0000012d;
  wire sig0000012e;
  wire sig0000012f;
  wire sig00000130;
  wire sig00000131;
  wire sig00000132;
  wire sig00000133;
  wire sig00000134;
  wire sig00000135;
  wire sig00000136;
  wire sig00000137;
  wire sig00000138;
  wire sig00000139;
  wire sig0000013a;
  wire sig0000013b;
  wire sig0000013c;
  wire sig0000013d;
  wire sig0000013e;
  wire sig0000013f;
  wire sig00000140;
  wire sig00000141;
  wire sig00000142;
  wire sig00000143;
  wire sig00000144;
  wire sig00000145;
  wire sig00000146;
  wire sig00000147;
  wire sig00000148;
  wire sig00000149;
  wire sig0000014a;
  wire sig0000014b;
  wire sig0000014c;
  wire sig0000014d;
  wire sig0000014e;
  wire sig0000014f;
  wire sig00000150;
  wire sig00000151;
  wire sig00000152;
  wire sig00000153;
  wire sig00000154;
  wire sig00000155;
  wire sig00000156;
  wire sig00000157;
  wire sig00000158;
  wire sig00000159;
  wire sig0000015a;
  wire sig0000015b;
  wire sig0000015c;
  wire sig0000015d;
  wire sig0000015e;
  wire sig0000015f;
  wire sig00000160;
  wire sig00000161;
  wire sig00000162;
  wire sig00000163;
  wire sig00000164;
  wire sig00000165;
  wire sig00000166;
  wire sig00000167;
  wire sig00000168;
  wire sig00000169;
  wire sig0000016a;
  wire sig0000016b;
  wire sig0000016c;
  wire sig0000016d;
  wire sig0000016e;
  wire sig0000016f;
  wire sig00000170;
  wire sig00000171;
  wire sig00000172;
  wire sig00000173;
  wire sig00000174;
  wire sig00000175;
  wire sig00000176;
  wire sig00000177;
  wire sig00000178;
  wire sig00000179;
  wire sig0000017a;
  wire sig0000017b;
  wire sig0000017c;
  wire sig0000017d;
  wire sig0000017e;
  wire sig0000017f;
  wire sig00000180;
  wire sig00000181;
  wire sig00000182;
  wire sig00000183;
  wire sig00000184;
  wire sig00000185;
  wire sig00000186;
  wire sig00000187;
  wire sig00000188;
  wire sig00000189;
  wire sig0000018a;
  wire sig0000018b;
  wire sig0000018c;
  wire sig0000018d;
  wire sig0000018e;
  wire sig0000018f;
  wire sig00000190;
  wire sig00000191;
  wire sig00000192;
  wire sig00000193;
  wire sig00000194;
  wire sig00000195;
  wire sig00000196;
  wire sig00000197;
  wire sig00000198;
  wire sig00000199;
  wire sig0000019a;
  wire sig0000019b;
  wire sig0000019c;
  wire sig0000019d;
  wire sig0000019e;
  wire sig0000019f;
  wire sig000001a0;
  wire sig000001a1;
  wire sig000001a2;
  wire sig000001a3;
  wire sig000001a4;
  wire sig000001a5;
  wire sig000001a6;
  wire sig000001a7;
  wire sig000001a8;
  wire sig000001a9;
  wire sig000001aa;
  wire sig000001ab;
  wire sig000001ac;
  wire sig000001ad;
  wire sig000001ae;
  wire sig000001af;
  wire sig000001b0;
  wire sig000001b1;
  wire sig000001b2;
  wire sig000001b3;
  wire sig000001b4;
  wire sig000001b5;
  wire sig000001b6;
  wire sig000001b7;
  wire sig000001b8;
  wire sig000001b9;
  wire sig000001ba;
  wire sig000001bb;
  wire sig000001bc;
  wire sig000001bd;
  wire sig000001be;
  wire sig000001bf;
  wire sig000001c0;
  wire sig000001c1;
  wire sig000001c2;
  wire sig000001c3;
  wire sig000001c4;
  wire sig000001c5;
  wire sig000001c6;
  wire sig000001c7;
  wire sig000001c8;
  wire sig000001c9;
  wire sig000001ca;
  wire sig000001cb;
  wire sig000001cc;
  wire sig000001cd;
  wire sig000001ce;
  wire sig000001cf;
  wire sig000001d0;
  wire sig000001d1;
  wire sig000001d2;
  wire sig000001d3;
  wire sig000001d4;
  wire sig000001d5;
  wire sig000001d6;
  wire sig000001d7;
  wire sig000001d8;
  wire sig000001d9;
  wire sig000001da;
  wire sig000001db;
  wire sig000001dc;
  wire sig000001dd;
  wire sig000001de;
  wire sig000001df;
  wire sig000001e0;
  wire sig000001e1;
  wire sig000001e2;
  wire sig000001e3;
  wire sig000001e4;
  wire sig000001e5;
  wire sig000001e6;
  wire sig000001e7;
  wire sig000001e8;
  wire sig000001e9;
  wire sig000001ea;
  wire sig000001eb;
  wire sig000001ec;
  wire sig000001ed;
  wire sig000001ee;
  wire sig000001ef;
  wire sig000001f0;
  wire sig000001f1;
  wire sig000001f2;
  wire sig000001f3;
  wire sig000001f4;
  wire sig000001f5;
  wire sig000001f6;
  wire sig000001f7;
  wire sig000001f8;
  wire sig000001f9;
  wire sig000001fa;
  wire sig000001fb;
  wire sig000001fc;
  wire sig000001fd;
  wire sig000001fe;
  wire sig000001ff;
  wire sig00000200;
  wire sig00000201;
  wire sig00000202;
  wire sig00000203;
  wire sig00000204;
  wire sig00000205;
  wire sig00000206;
  wire sig00000207;
  wire sig00000208;
  wire sig00000209;
  wire sig0000020a;
  wire sig0000020b;
  wire sig0000020c;
  wire sig0000020d;
  wire sig0000020e;
  wire sig0000020f;
  wire sig00000210;
  wire sig00000211;
  wire sig00000212;
  wire sig00000213;
  wire sig00000214;
  wire sig00000215;
  wire sig00000216;
  wire sig00000217;
  wire sig00000218;
  wire sig00000219;
  wire sig0000021a;
  wire sig0000021b;
  wire sig0000021c;
  wire sig0000021d;
  wire sig0000021e;
  wire sig0000021f;
  wire sig00000220;
  wire sig00000221;
  wire sig00000222;
  wire sig00000223;
  wire sig00000224;
  wire sig00000225;
  wire sig00000226;
  wire sig00000227;
  wire sig00000228;
  wire sig00000229;
  wire sig0000022a;
  wire sig0000022b;
  wire sig0000022c;
  wire sig0000022d;
  wire sig0000022e;
  wire sig0000022f;
  wire sig00000230;
  wire sig00000231;
  wire sig00000232;
  wire sig00000233;
  wire sig00000234;
  wire sig00000235;
  wire sig00000236;
  wire sig00000237;
  wire sig00000238;
  wire sig00000239;
  wire sig0000023a;
  wire sig0000023b;
  wire sig0000023c;
  wire sig0000023d;
  wire sig0000023e;
  wire sig0000023f;
  wire sig00000240;
  wire sig00000241;
  wire sig00000242;
  wire sig00000243;
  wire sig00000244;
  wire sig00000245;
  wire sig00000246;
  wire sig00000247;
  wire sig00000248;
  wire sig00000249;
  wire sig0000024a;
  wire sig0000024b;
  wire sig0000024c;
  wire sig0000024d;
  wire sig0000024e;
  wire sig0000024f;
  wire sig00000250;
  wire sig00000251;
  wire sig00000252;
  wire sig00000253;
  wire sig00000254;
  wire sig00000255;
  wire sig00000256;
  wire sig00000257;
  wire sig00000258;
  wire sig00000259;
  wire sig0000025a;
  wire sig0000025b;
  wire sig0000025c;
  wire sig0000025d;
  wire sig0000025e;
  wire sig0000025f;
  wire sig00000260;
  wire sig00000261;
  wire sig00000262;
  wire sig00000263;
  wire sig00000264;
  wire sig00000265;
  wire sig00000266;
  wire sig00000267;
  wire sig00000268;
  wire sig00000269;
  wire sig0000026a;
  wire sig0000026b;
  wire sig0000026c;
  wire sig0000026d;
  wire sig0000026e;
  wire sig0000026f;
  wire sig00000270;
  wire sig00000271;
  wire sig00000272;
  wire sig00000273;
  wire sig00000274;
  wire sig00000275;
  wire sig00000276;
  wire sig00000277;
  wire sig00000278;
  wire sig00000279;
  wire sig0000027a;
  wire sig0000027b;
  wire sig0000027c;
  wire sig0000027d;
  wire sig0000027e;
  wire sig0000027f;
  wire sig00000280;
  wire sig00000281;
  wire sig00000282;
  wire sig00000283;
  wire sig00000284;
  wire sig00000285;
  wire sig00000286;
  wire sig00000287;
  wire sig00000288;
  wire sig00000289;
  wire sig0000028a;
  wire sig0000028b;
  wire sig0000028c;
  wire sig0000028d;
  wire sig0000028e;
  wire sig0000028f;
  wire sig00000290;
  wire sig00000291;
  wire sig00000292;
  wire sig00000293;
  wire sig00000294;
  wire sig00000295;
  wire sig00000296;
  wire sig00000297;
  wire sig00000298;
  wire sig00000299;
  wire sig0000029a;
  wire sig0000029b;
  wire sig0000029c;
  wire sig0000029d;
  wire sig0000029e;
  wire sig0000029f;
  wire sig000002a0;
  wire sig000002a1;
  wire sig000002a2;
  wire sig000002a3;
  wire sig000002a4;
  wire sig000002a5;
  wire sig000002a6;
  wire sig000002a7;
  wire sig000002a8;
  wire sig000002a9;
  wire sig000002aa;
  wire sig000002ab;
  wire sig000002ac;
  wire sig000002ad;
  wire sig000002ae;
  wire sig000002af;
  wire sig000002b0;
  wire sig000002b1;
  wire sig000002b2;
  wire sig000002b3;
  wire sig000002b4;
  wire sig000002b5;
  wire sig000002b6;
  wire sig000002b7;
  wire sig000002b8;
  wire sig000002b9;
  wire sig000002ba;
  wire sig000002bb;
  wire sig000002bc;
  wire sig000002bd;
  wire sig000002be;
  wire sig000002bf;
  wire sig000002c0;
  wire sig000002c1;
  wire sig000002c2;
  wire sig000002c3;
  wire sig000002c4;
  wire sig000002c5;
  wire sig000002c6;
  wire sig000002c7;
  wire sig000002c8;
  wire sig000002c9;
  wire sig000002ca;
  wire sig000002cb;
  wire sig000002cc;
  wire sig000002cd;
  wire sig000002ce;
  wire sig000002cf;
  wire sig000002d0;
  wire sig000002d1;
  wire sig000002d2;
  wire sig000002d3;
  wire sig000002d4;
  wire sig000002d5;
  wire sig000002d6;
  wire sig000002d7;
  wire sig000002d8;
  wire sig000002d9;
  wire sig000002da;
  wire sig000002db;
  wire sig000002dc;
  wire sig000002dd;
  wire sig000002de;
  wire sig000002df;
  wire sig000002e0;
  wire sig000002e1;
  wire sig000002e2;
  wire sig000002e3;
  wire sig000002e4;
  wire sig000002e5;
  wire sig000002e6;
  wire sig000002e7;
  wire sig000002e8;
  wire sig000002e9;
  wire sig000002ea;
  wire sig000002eb;
  wire sig000002ec;
  wire sig000002ed;
  wire sig000002ee;
  wire sig000002ef;
  wire sig000002f0;
  wire sig000002f1;
  wire sig000002f2;
  wire sig000002f3;
  wire sig000002f4;
  wire sig000002f5;
  wire sig000002f6;
  wire sig000002f7;
  wire sig000002f8;
  wire sig000002f9;
  wire sig000002fa;
  wire sig000002fb;
  wire sig000002fc;
  wire sig000002fd;
  wire sig000002fe;
  wire sig000002ff;
  wire sig00000300;
  wire sig00000301;
  wire sig00000302;
  wire sig00000303;
  wire sig00000304;
  wire sig00000305;
  wire sig00000306;
  wire sig00000307;
  wire sig00000308;
  wire sig00000309;
  wire sig0000030a;
  wire sig0000030c;
  wire sig0000030d;
  wire sig0000030e;
  wire sig0000030f;
  wire sig00000310;
  wire sig00000311;
  wire sig00000312;
  wire sig00000313;
  wire sig00000314;
  wire sig00000315;
  wire sig00000316;
  wire sig00000317;
  wire sig00000318;
  wire sig00000319;
  wire sig0000031a;
  wire sig0000031b;
  wire sig0000031c;
  wire sig0000031d;
  wire sig0000031e;
  wire sig0000031f;
  wire sig00000320;
  wire sig00000329;
  wire sig0000032a;
  wire sig0000032b;
  wire sig0000032c;
  wire sig0000032d;
  wire sig0000032e;
  wire sig0000032f;
  wire sig00000330;
  wire sig00000331;
  wire sig00000332;
  wire sig00000333;
  wire sig00000334;
  wire sig00000335;
  wire sig00000336;
  wire sig00000337;
  wire sig00000338;
  wire sig00000339;
  wire sig0000033a;
  wire sig0000033b;
  wire sig0000033c;
  wire sig0000033d;
  wire sig0000033e;
  wire sig0000033f;
  wire sig00000340;
  wire sig00000341;
  wire sig00000342;
  wire sig00000343;
  wire sig00000344;
  wire sig00000345;
  wire sig00000346;
  wire sig00000347;
  wire sig00000348;
  wire sig00000349;
  wire sig0000034a;
  wire sig00000356;
  wire sig00000357;
  wire sig00000358;
  wire sig00000359;
  wire sig0000035a;
  wire sig0000035b;
  wire sig0000035c;
  wire sig0000035d;
  wire sig0000035e;
  wire sig0000035f;
  wire sig00000360;
  wire sig00000361;
  wire sig00000362;
  wire sig00000363;
  wire sig00000364;
  wire sig00000365;
  wire sig00000366;
  wire sig00000367;
  wire sig00000368;
  wire sig00000369;
  wire sig0000036a;
  wire sig0000036b;
  wire sig0000036c;
  wire sig0000036d;
  wire sig0000036e;
  wire sig0000036f;
  wire sig00000370;
  wire sig00000371;
  wire sig00000372;
  wire sig00000373;
  wire sig00000374;
  wire sig00000375;
  wire sig00000376;
  wire sig00000377;
  wire sig00000378;
  wire sig00000379;
  wire sig0000037a;
  wire sig0000037b;
  wire sig0000037c;
  wire sig0000037d;
  wire sig0000037e;
  wire sig0000037f;
  wire sig00000380;
  wire sig00000381;
  wire sig00000382;
  wire sig00000383;
  wire sig00000384;
  wire sig00000385;
  wire sig00000386;
  wire sig00000387;
  wire sig00000388;
  wire sig00000389;
  wire sig0000038a;
  wire sig0000038b;
  wire sig0000038c;
  wire sig0000038d;
  wire sig0000038e;
  wire sig0000038f;
  wire sig00000390;
  wire sig00000391;
  wire sig00000392;
  wire sig00000393;
  wire sig00000394;
  wire sig00000395;
  wire sig00000396;
  wire sig00000397;
  wire sig00000398;
  wire sig00000399;
  wire sig0000039a;
  wire sig0000039b;
  wire sig0000039c;
  wire sig0000039d;
  wire sig0000039e;
  wire sig0000039f;
  wire sig000003a0;
  wire sig000003a1;
  wire sig000003a2;
  wire sig000003a3;
  wire sig000003a4;
  wire sig000003a5;
  wire sig000003a6;
  wire sig000003a7;
  wire sig000003a8;
  wire sig000003a9;
  wire sig000003aa;
  wire sig000003ab;
  wire sig000003ac;
  wire sig000003ad;
  wire sig000003ae;
  wire sig000003af;
  wire sig000003b0;
  wire sig000003b1;
  wire sig000003b2;
  wire sig000003b3;
  wire sig000003b4;
  wire sig000003b5;
  wire sig000003b6;
  wire sig000003b7;
  wire sig000003b8;
  wire sig000003b9;
  wire sig000003ba;
  wire sig000003bb;
  wire sig000003bc;
  wire sig000003bd;
  wire sig000003be;
  wire sig000003bf;
  wire sig000003c0;
  wire sig000003c1;
  wire sig000003c2;
  wire sig000003c3;
  wire sig000003c4;
  wire sig000003c5;
  wire sig000003c6;
  wire sig000003c7;
  wire sig000003c9;
  wire sig000003ca;
  wire sig000003cb;
  wire sig000003cc;
  wire sig000003cd;
  wire sig000003ce;
  wire sig000003cf;
  wire sig000003d0;
  wire sig000003d1;
  wire sig000003d2;
  wire sig000003d3;
  wire sig000003d4;
  wire sig000003d5;
  wire sig000003d6;
  wire sig000003d7;
  wire sig000003d8;
  wire sig000003d9;
  wire sig000003da;
  wire sig000003db;
  wire sig000003dc;
  wire sig000003e5;
  wire sig000003e6;
  wire sig000003e7;
  wire sig000003e8;
  wire sig000003e9;
  wire sig000003ea;
  wire sig000003eb;
  wire sig000003ec;
  wire sig000003ed;
  wire sig000003ee;
  wire sig000003ef;
  wire sig000003f0;
  wire sig000003f1;
  wire sig000003f2;
  wire sig000003f3;
  wire sig000003f4;
  wire sig000003f5;
  wire sig000003f6;
  wire sig000003f7;
  wire sig000003f8;
  wire sig000003f9;
  wire sig000003fa;
  wire sig000003fb;
  wire sig000003fc;
  wire sig000003fd;
  wire sig000003fe;
  wire sig000003ff;
  wire sig00000400;
  wire sig00000401;
  wire sig00000402;
  wire sig00000403;
  wire sig00000404;
  wire sig00000405;
  wire sig00000406;
  wire sig00000407;
  wire sig00000408;
  wire sig00000409;
  wire sig0000040a;
  wire sig0000040b;
  wire sig0000040c;
  wire sig0000040d;
  wire sig0000040e;
  wire sig0000040f;
  wire sig00000410;
  wire sig00000411;
  wire sig00000412;
  wire sig00000413;
  wire sig00000414;
  wire sig00000415;
  wire sig00000416;
  wire sig00000417;
  wire sig00000418;
  wire sig00000419;
  wire sig0000041a;
  wire sig0000041b;
  wire sig0000041c;
  wire sig0000041d;
  wire sig0000041e;
  wire sig0000041f;
  wire sig00000420;
  wire sig00000421;
  wire sig00000422;
  wire sig00000423;
  wire sig00000424;
  wire sig00000425;
  wire sig00000426;
  wire sig00000427;
  wire sig00000428;
  wire sig00000429;
  wire sig0000042a;
  wire sig0000042b;
  wire sig0000042c;
  wire sig0000042d;
  wire sig0000042e;
  wire sig0000042f;
  wire sig00000430;
  wire sig00000431;
  wire sig00000432;
  wire sig00000433;
  wire sig00000434;
  wire sig00000435;
  wire sig00000436;
  wire sig00000437;
  wire sig00000438;
  wire sig00000439;
  wire sig0000043a;
  wire sig0000043b;
  wire sig0000043c;
  wire sig0000043d;
  wire sig0000043e;
  wire sig0000043f;
  wire sig00000440;
  wire sig00000441;
  wire sig00000442;
  wire sig00000443;
  wire sig00000444;
  wire sig00000445;
  wire sig00000446;
  wire sig00000447;
  wire sig00000448;
  wire sig00000449;
  wire sig0000044a;
  wire sig0000044b;
  wire sig0000044c;
  wire sig0000044d;
  wire sig0000044e;
  wire sig0000044f;
  wire sig00000450;
  wire sig00000451;
  wire sig00000452;
  wire sig00000453;
  wire sig00000454;
  wire sig00000455;
  wire sig00000456;
  wire sig00000457;
  wire sig00000458;
  wire sig00000459;
  wire sig0000045a;
  wire sig0000045b;
  wire sig0000045c;
  wire sig0000045d;
  wire sig0000045e;
  wire sig0000045f;
  wire sig00000460;
  wire sig00000461;
  wire sig00000462;
  wire sig00000463;
  wire sig00000464;
  wire sig00000465;
  wire sig00000466;
  wire sig00000467;
  wire sig00000468;
  wire sig00000469;
  wire sig0000046a;
  wire sig0000046b;
  wire sig0000046c;
  wire sig0000046d;
  wire sig0000046e;
  wire sig0000046f;
  wire sig00000470;
  wire sig00000471;
  wire sig00000472;
  wire sig00000473;
  wire sig00000474;
  wire sig00000475;
  wire sig00000476;
  wire sig00000477;
  wire sig00000478;
  wire sig00000479;
  wire sig0000047a;
  wire sig0000047b;
  wire sig0000047c;
  wire sig0000047d;
  wire sig0000047e;
  wire sig0000047f;
  wire sig00000480;
  wire sig00000481;
  wire sig00000482;
  wire sig00000483;
  wire sig00000484;
  wire sig00000485;
  wire sig00000486;
  wire sig000004a1;
  wire sig000004a2;
  wire sig000004a3;
  wire sig000004a4;
  wire sig000004a5;
  wire sig000004a6;
  wire sig000004a7;
  wire sig000004a8;
  wire sig000004a9;
  wire sig000004aa;
  wire sig000004ab;
  wire sig000004ac;
  wire sig000004ad;
  wire sig000004ae;
  wire sig000004af;
  wire sig000004b0;
  wire sig000004b1;
  wire sig000004b2;
  wire sig000004b3;
  wire sig000004b4;
  wire sig000004c2;
  wire sig000004c3;
  wire sig000004c4;
  wire sig000004c5;
  wire sig000004c6;
  wire sig000004c7;
  wire sig000004c8;
  wire sig000004c9;
  wire sig000004ca;
  wire sig000004cb;
  wire sig000004cd;
  wire sig000004ce;
  wire sig000004cf;
  wire sig000004d0;
  wire sig000004d1;
  wire sig000004d2;
  wire sig000004d3;
  wire sig000004d4;
  wire sig000004d5;
  wire sig000004d6;
  wire sig000004d7;
  wire sig000004d8;
  wire sig000004d9;
  wire sig000004da;
  wire sig000004db;
  wire sig000004dc;
  wire sig000004dd;
  wire sig000004de;
  wire sig000004df;
  wire sig000004e0;
  wire sig000004e1;
  wire sig000004e2;
  wire sig000004e3;
  wire sig000004e4;
  wire sig000004e5;
  wire sig000004e6;
  wire sig000004e7;
  wire sig000004e8;
  wire sig000004e9;
  wire sig000004f4;
  wire sig000004f5;
  wire sig000004f6;
  wire sig000004f7;
  wire sig000004f8;
  wire sig000004f9;
  wire sig000004fa;
  wire sig000004fb;
  wire sig000004fc;
  wire sig000004fd;
  wire sig000004fe;
  wire sig000004ff;
  wire sig00000500;
  wire sig00000501;
  wire sig00000502;
  wire sig00000503;
  wire sig00000504;
  wire sig00000505;
  wire sig00000506;
  wire sig00000518;
  wire sig00000519;
  wire sig0000051a;
  wire sig0000051b;
  wire sig0000051c;
  wire sig0000051d;
  wire sig0000051e;
  wire sig0000051f;
  wire sig00000520;
  wire sig00000521;
  wire sig00000522;
  wire sig00000523;
  wire sig0000052f;
  wire sig00000530;
  wire sig00000531;
  wire sig00000532;
  wire sig00000533;
  wire sig00000534;
  wire sig00000535;
  wire sig00000536;
  wire sig00000537;
  wire sig00000538;
  wire sig00000539;
  wire sig0000053a;
  wire sig0000053b;
  wire sig0000053c;
  wire sig0000053d;
  wire sig0000053e;
  wire sig0000053f;
  wire sig00000540;
  wire sig00000541;
  wire sig00000542;
  wire sig00000543;
  wire sig00000544;
  wire sig00000545;
  wire sig00000546;
  wire sig00000547;
  wire sig0000055b;
  wire sig0000055c;
  wire sig0000055d;
  wire sig00000570;
  wire sig00000571;
  wire sig00000572;
  wire sig00000573;
  wire sig00000574;
  wire sig00000575;
  wire sig00000576;
  wire sig00000577;
  wire sig00000578;
  wire sig00000579;
  wire sig0000057a;
  wire sig0000057b;
  wire sig0000057c;
  wire sig0000057d;
  wire sig0000057e;
  wire sig0000057f;
  wire sig00000580;
  wire sig00000581;
  wire sig00000582;
  wire sig00000583;
  wire sig00000584;
  wire sig00000585;
  wire sig00000586;
  wire sig00000587;
  wire sig00000588;
  wire sig00000589;
  wire sig0000058a;
  wire sig0000058b;
  wire sig0000058c;
  wire sig0000058d;
  wire sig0000058e;
  wire sig0000058f;
  wire sig00000590;
  wire sig00000591;
  wire sig00000592;
  wire sig00000593;
  wire sig00000594;
  wire sig00000595;
  wire sig00000596;
  wire sig00000597;
  wire sig00000598;
  wire sig00000599;
  wire sig0000059a;
  wire sig0000059b;
  wire sig0000059c;
  wire sig0000059d;
  wire sig0000059e;
  wire sig0000059f;
  wire sig000005a0;
  wire sig000005a1;
  wire sig000005a2;
  wire sig000005a3;
  wire sig000005a4;
  wire sig000005a5;
  wire sig000005a6;
  wire sig000005a7;
  wire sig000005a8;
  wire sig000005a9;
  wire sig000005aa;
  wire sig000005ab;
  wire sig000005ac;
  wire sig000005ad;
  wire sig000005ae;
  wire sig000005af;
  wire sig000005b0;
  wire sig000005b1;
  wire sig000005b2;
  wire sig000005b3;
  wire sig000005b4;
  wire sig000005b5;
  wire sig000005b6;
  wire sig000005b7;
  wire sig000005b8;
  wire sig000005b9;
  wire sig000005ba;
  wire sig000005bb;
  wire sig000005bc;
  wire sig000005bd;
  wire sig000005be;
  wire sig000005bf;
  wire sig000005c0;
  wire sig000005c1;
  wire sig000005c2;
  wire sig000005c3;
  wire sig000005c4;
  wire sig000005c5;
  wire sig000005c6;
  wire sig000005c7;
  wire sig000005c8;
  wire sig000005c9;
  wire sig000005ca;
  wire sig000005cb;
  wire sig000005cc;
  wire sig000005cd;
  wire sig000005ce;
  wire sig000005cf;
  wire sig000005d0;
  wire sig000005d1;
  wire sig000005d2;
  wire sig000005d3;
  wire sig000005d4;
  wire sig000005d5;
  wire sig000005d6;
  wire sig000005d7;
  wire sig000005d8;
  wire sig000005d9;
  wire sig000005da;
  wire sig000005db;
  wire sig000005dc;
  wire sig000005dd;
  wire sig000005de;
  wire sig000005df;
  wire sig000005e0;
  wire sig000005e1;
  wire sig000005e2;
  wire sig000005e3;
  wire sig000005e4;
  wire sig000005e5;
  wire sig000005e6;
  wire sig000005e7;
  wire sig000005e8;
  wire sig000005e9;
  wire sig000005ea;
  wire sig000005eb;
  wire sig000005ec;
  wire sig000005ed;
  wire sig000005ee;
  wire sig000005ef;
  wire sig000005f0;
  wire sig000005f1;
  wire sig000005f2;
  wire sig000005f3;
  wire sig000005f4;
  wire sig000005f5;
  wire sig000005f6;
  wire sig000005f7;
  wire sig000005f8;
  wire sig000005f9;
  wire sig000005fa;
  wire sig000005fb;
  wire sig000005fc;
  wire sig000005fd;
  wire sig000005fe;
  wire sig000005ff;
  wire sig00000600;
  wire sig00000601;
  wire sig00000602;
  wire sig00000603;
  wire sig00000604;
  wire sig00000605;
  wire sig00000606;
  wire sig00000607;
  wire sig00000608;
  wire sig00000609;
  wire sig0000060a;
  wire sig0000060b;
  wire sig0000060c;
  wire sig0000060d;
  wire sig0000060e;
  wire sig0000060f;
  wire sig00000610;
  wire sig00000611;
  wire sig00000612;
  wire sig00000613;
  wire sig00000614;
  wire sig00000615;
  wire sig00000616;
  wire sig00000617;
  wire sig00000618;
  wire sig00000619;
  wire sig0000061a;
  wire sig0000061b;
  wire sig0000061c;
  wire sig0000061d;
  wire sig0000061e;
  wire sig0000061f;
  wire sig00000620;
  wire sig00000621;
  wire sig00000622;
  wire sig00000623;
  wire sig00000624;
  wire sig00000625;
  wire sig00000626;
  wire sig00000627;
  wire sig00000628;
  wire sig00000629;
  wire sig0000062a;
  wire sig0000062b;
  wire sig0000062c;
  wire sig0000062d;
  wire sig0000062e;
  wire sig0000062f;
  wire sig00000630;
  wire sig00000631;
  wire sig00000632;
  wire sig00000633;
  wire sig00000634;
  wire sig00000635;
  wire sig00000636;
  wire sig00000637;
  wire sig00000638;
  wire sig00000639;
  wire sig0000063a;
  wire sig0000063b;
  wire sig0000063c;
  wire sig0000063d;
  wire sig0000063e;
  wire sig0000063f;
  wire sig00000640;
  wire sig00000641;
  wire sig00000642;
  wire sig00000643;
  wire sig00000644;
  wire sig00000645;
  wire sig00000646;
  wire sig00000647;
  wire sig00000648;
  wire sig00000649;
  wire sig0000064a;
  wire sig0000064b;
  wire sig0000064c;
  wire sig0000064d;
  wire sig0000064e;
  wire sig0000064f;
  wire sig00000650;
  wire sig00000651;
  wire sig00000652;
  wire sig00000653;
  wire sig00000654;
  wire sig00000655;
  wire sig00000656;
  wire sig00000657;
  wire sig00000658;
  wire sig00000659;
  wire sig0000065a;
  wire sig0000065b;
  wire sig0000065c;
  wire sig0000065d;
  wire sig0000065e;
  wire sig0000065f;
  wire sig00000660;
  wire sig00000661;
  wire sig00000662;
  wire sig00000663;
  wire sig00000664;
  wire sig00000665;
  wire sig00000666;
  wire sig00000667;
  wire sig00000668;
  wire sig00000669;
  wire sig0000066a;
  wire sig0000066b;
  wire sig0000066c;
  wire sig0000066d;
  wire sig0000066e;
  wire sig0000066f;
  wire sig00000670;
  wire sig00000671;
  wire sig00000672;
  wire sig00000673;
  wire sig00000674;
  wire sig00000675;
  wire sig00000676;
  wire sig00000677;
  wire sig00000678;
  wire sig00000679;
  wire sig0000067a;
  wire sig0000067b;
  wire sig0000067c;
  wire sig0000067d;
  wire sig0000067e;
  wire sig0000067f;
  wire sig00000680;
  wire sig00000681;
  wire sig00000682;
  wire sig00000683;
  wire sig00000684;
  wire sig00000685;
  wire sig00000686;
  wire sig00000687;
  wire sig00000688;
  wire sig00000689;
  wire sig0000068a;
  wire sig0000068b;
  wire sig0000068c;
  wire sig0000068d;
  wire sig0000068e;
  wire sig0000068f;
  wire sig00000690;
  wire sig00000691;
  wire sig00000692;
  wire sig00000693;
  wire sig00000694;
  wire sig00000695;
  wire sig00000696;
  wire sig00000697;
  wire sig00000698;
  wire sig00000699;
  wire sig0000069a;
  wire sig0000069b;
  wire sig0000069c;
  wire sig0000069d;
  wire sig0000069e;
  wire sig0000069f;
  wire sig000006a0;
  wire sig000006a1;
  wire sig000006a2;
  wire sig000006a3;
  wire sig000006a4;
  wire sig000006a5;
  wire sig000006a6;
  wire sig000006a7;
  wire sig000006a8;
  wire sig000006a9;
  wire sig000006aa;
  wire sig000006ab;
  wire sig000006ac;
  wire sig000006ad;
  wire sig000006ae;
  wire sig000006af;
  wire sig000006b0;
  wire sig000006b1;
  wire sig000006b2;
  wire sig000006b3;
  wire sig000006b4;
  wire sig000006b5;
  wire sig000006b6;
  wire sig000006b7;
  wire sig000006b8;
  wire sig000006b9;
  wire sig000006ba;
  wire sig000006bb;
  wire sig000006bc;
  wire sig000006bd;
  wire sig000006be;
  wire sig000006bf;
  wire sig000006c0;
  wire sig000006c1;
  wire sig000006c2;
  wire sig000006c3;
  wire sig000006c4;
  wire sig000006c5;
  wire sig000006c6;
  wire sig000006c7;
  wire sig000006c8;
  wire sig000006c9;
  wire sig000006ca;
  wire sig000006cb;
  wire sig000006cc;
  wire sig000006cd;
  wire sig000006ce;
  wire sig000006cf;
  wire sig000006d0;
  wire sig000006d1;
  wire sig000006d2;
  wire sig000006d3;
  wire sig000006d4;
  wire sig000006d5;
  wire sig000006d6;
  wire sig000006d7;
  wire sig000006d8;
  wire sig000006d9;
  wire sig000006da;
  wire sig000006db;
  wire sig000006dc;
  wire sig000006dd;
  wire sig000006de;
  wire sig000006df;
  wire sig000006e0;
  wire sig000006e1;
  wire sig000006e2;
  wire sig000006e3;
  wire sig000006e4;
  wire sig000006e5;
  wire sig000006e6;
  wire sig000006e7;
  wire sig000006e8;
  wire sig000006e9;
  wire sig000006ea;
  wire sig000006eb;
  wire sig000006ec;
  wire sig000006ed;
  wire sig000006ee;
  wire sig000006ef;
  wire sig000006f0;
  wire sig000006f1;
  wire sig000006f2;
  wire sig000006f3;
  wire sig000006f4;
  wire sig000006f5;
  wire sig000006f6;
  wire sig000006f7;
  wire sig000006f8;
  wire sig000006f9;
  wire sig000006fa;
  wire sig000006fb;
  wire sig000006fc;
  wire sig000006fd;
  wire sig000006fe;
  wire sig000006ff;
  wire sig00000700;
  wire sig00000701;
  wire sig00000702;
  wire sig00000703;
  wire sig00000704;
  wire sig00000705;
  wire sig00000706;
  wire sig00000707;
  wire sig00000708;
  wire sig00000709;
  wire sig0000070a;
  wire sig0000070b;
  wire sig0000070c;
  wire sig0000070d;
  wire sig0000070e;
  wire sig0000070f;
  wire sig00000710;
  wire sig00000711;
  wire sig00000712;
  wire sig00000713;
  wire sig00000714;
  wire sig00000715;
  wire sig00000716;
  wire sig00000717;
  wire sig00000718;
  wire sig00000719;
  wire sig0000071a;
  wire sig0000071b;
  wire sig0000071c;
  wire sig0000071d;
  wire sig0000071e;
  wire sig0000071f;
  wire sig00000720;
  wire sig00000721;
  wire sig00000722;
  wire sig00000723;
  wire sig00000724;
  wire sig00000725;
  wire sig00000726;
  wire sig00000727;
  wire sig00000728;
  wire sig00000729;
  wire sig0000072a;
  wire sig0000072b;
  wire sig0000072c;
  wire sig0000072d;
  wire sig0000072e;
  wire sig0000072f;
  wire sig00000730;
  wire sig00000731;
  wire sig00000732;
  wire sig00000733;
  wire sig00000734;
  wire sig00000735;
  wire sig00000736;
  wire sig00000737;
  wire sig00000738;
  wire sig00000739;
  wire sig0000073a;
  wire sig0000073b;
  wire sig0000073c;
  wire sig0000073d;
  wire sig0000073e;
  wire sig0000073f;
  wire sig00000740;
  wire sig00000741;
  wire sig00000742;
  wire sig00000743;
  wire sig00000744;
  wire sig00000745;
  wire sig00000746;
  wire sig00000747;
  wire sig00000748;
  wire sig00000749;
  wire sig0000074a;
  wire sig0000074b;
  wire sig0000074c;
  wire sig0000074d;
  wire sig0000074e;
  wire sig0000074f;
  wire sig00000750;
  wire sig00000751;
  wire sig00000752;
  wire sig00000753;
  wire sig00000754;
  wire sig00000755;
  wire sig00000756;
  wire sig00000757;
  wire sig00000758;
  wire sig00000759;
  wire sig0000075a;
  wire sig0000075b;
  wire sig0000075c;
  wire sig0000075d;
  wire sig0000075e;
  wire sig0000075f;
  wire sig00000760;
  wire sig00000761;
  wire sig00000762;
  wire sig00000763;
  wire sig00000764;
  wire sig00000765;
  wire sig00000766;
  wire sig00000767;
  wire sig00000768;
  wire sig00000769;
  wire sig0000076a;
  wire sig0000076b;
  wire sig0000076c;
  wire sig0000076d;
  wire sig0000076e;
  wire sig0000076f;
  wire sig00000770;
  wire sig00000771;
  wire sig00000772;
  wire sig00000773;
  wire sig00000774;
  wire sig00000775;
  wire sig00000776;
  wire sig00000777;
  wire sig00000778;
  wire sig00000779;
  wire sig0000077a;
  wire sig0000077b;
  wire sig0000077c;
  wire sig0000077d;
  wire sig0000077e;
  wire sig0000077f;
  wire sig00000780;
  wire sig00000781;
  wire sig00000782;
  wire sig00000783;
  wire sig00000784;
  wire sig00000785;
  wire sig00000786;
  wire sig00000787;
  wire sig00000788;
  wire sig00000789;
  wire sig0000078a;
  wire sig0000078b;
  wire sig0000078c;
  wire sig0000078d;
  wire sig0000078e;
  wire sig0000078f;
  wire sig00000790;
  wire sig00000791;
  wire sig00000792;
  wire sig00000793;
  wire sig00000794;
  wire sig00000795;
  wire sig00000796;
  wire sig00000797;
  wire sig00000798;
  wire sig00000799;
  wire sig0000079a;
  wire sig0000079b;
  wire sig0000079c;
  wire sig0000079d;
  wire sig0000079e;
  wire sig0000079f;
  wire sig000007a0;
  wire sig000007a1;
  wire sig000007a2;
  wire sig000007a3;
  wire sig000007a4;
  wire sig000007a5;
  wire sig000007a6;
  wire sig000007a7;
  wire sig000007a8;
  wire sig000007a9;
  wire sig000007aa;
  wire sig000007ab;
  wire sig000007ac;
  wire sig000007ad;
  wire sig000007ae;
  wire sig000007af;
  wire sig000007b0;
  wire sig000007b1;
  wire sig000007b2;
  wire sig000007b3;
  wire sig000007b4;
  wire sig000007b5;
  wire sig000007b6;
  wire sig000007b7;
  wire sig000007b8;
  wire sig000007b9;
  wire sig000007ba;
  wire sig000007bb;
  wire sig000007bc;
  wire sig000007bd;
  wire sig000007be;
  wire sig000007bf;
  wire sig000007c0;
  wire sig000007c1;
  wire sig000007c2;
  wire sig000007c3;
  wire sig000007c4;
  wire sig000007c5;
  wire sig000007c6;
  wire sig000007c7;
  wire sig000007c8;
  wire sig000007c9;
  wire sig000007ca;
  wire sig000007cb;
  wire sig000007cc;
  wire sig000007cd;
  wire sig000007ce;
  wire sig000007cf;
  wire sig000007d0;
  wire sig000007d1;
  wire sig000007d2;
  wire sig000007d3;
  wire sig000007d4;
  wire sig000007d5;
  wire sig000007d6;
  wire sig000007d7;
  wire sig000007d8;
  wire sig000007d9;
  wire sig000007da;
  wire sig000007db;
  wire sig000007dc;
  wire sig000007dd;
  wire sig000007de;
  wire sig000007df;
  wire sig000007e0;
  wire sig000007e1;
  wire sig000007e2;
  wire sig000007e3;
  wire sig000007e4;
  wire sig000007e5;
  wire sig000007e6;
  wire sig000007e7;
  wire sig000007e8;
  wire sig000007e9;
  wire sig000007ea;
  wire sig000007eb;
  wire sig000007ec;
  wire sig000007ed;
  wire sig000007ee;
  wire sig000007ef;
  wire sig000007f0;
  wire sig000007f1;
  wire sig000007f2;
  wire sig000007f3;
  wire sig000007f4;
  wire sig000007f5;
  wire sig000007f6;
  wire sig000007f7;
  wire sig000007f8;
  wire sig000007f9;
  wire sig000007fa;
  wire sig000007fb;
  wire sig000007fc;
  wire sig000007fd;
  wire sig000007fe;
  wire sig000007ff;
  wire sig00000800;
  wire sig00000801;
  wire sig00000802;
  wire sig00000803;
  wire sig00000804;
  wire sig00000805;
  wire sig00000806;
  wire sig00000807;
  wire sig00000808;
  wire sig00000809;
  wire sig0000080a;
  wire sig0000080b;
  wire sig0000080c;
  wire sig0000080d;
  wire sig0000080e;
  wire sig0000080f;
  wire sig00000810;
  wire sig00000811;
  wire sig00000812;
  wire sig00000813;
  wire sig00000814;
  wire sig00000815;
  wire sig00000816;
  wire sig00000817;
  wire sig00000818;
  wire sig00000819;
  wire sig0000081a;
  wire sig0000081b;
  wire sig0000081c;
  wire sig0000081d;
  wire sig0000081e;
  wire sig0000081f;
  wire sig00000820;
  wire sig00000821;
  wire sig00000822;
  wire sig00000823;
  wire sig00000824;
  wire sig00000825;
  wire sig00000826;
  wire sig00000827;
  wire sig00000828;
  wire sig00000829;
  wire sig0000082a;
  wire sig0000082b;
  wire sig0000082c;
  wire sig0000082d;
  wire sig0000082e;
  wire sig0000082f;
  wire sig00000830;
  wire sig00000831;
  wire sig00000832;
  wire sig00000833;
  wire sig00000834;
  wire sig00000835;
  wire sig00000836;
  wire sig00000837;
  wire sig00000838;
  wire sig00000839;
  wire sig0000083a;
  wire sig0000083b;
  wire sig0000083c;
  wire sig0000083d;
  wire sig0000083e;
  wire sig0000083f;
  wire sig00000840;
  wire sig00000841;
  wire sig00000842;
  wire sig00000843;
  wire sig00000844;
  wire sig00000845;
  wire sig00000846;
  wire sig00000847;
  wire sig00000848;
  wire sig00000849;
  wire sig0000084a;
  wire sig0000084b;
  wire sig0000084c;
  wire sig0000084d;
  wire sig0000084e;
  wire sig0000084f;
  wire sig00000850;
  wire sig00000851;
  wire sig00000852;
  wire sig00000853;
  wire sig00000854;
  wire sig00000855;
  wire sig00000856;
  wire sig00000857;
  wire sig00000858;
  wire sig00000859;
  wire sig0000085a;
  wire sig0000085b;
  wire sig0000085c;
  wire sig0000085d;
  wire sig0000085e;
  wire sig0000085f;
  wire sig00000860;
  wire sig00000861;
  wire sig00000862;
  wire sig00000863;
  wire sig00000864;
  wire sig00000865;
  wire sig00000866;
  wire sig00000867;
  wire sig00000868;
  wire sig00000869;
  wire sig0000086a;
  wire sig0000086b;
  wire sig0000086c;
  wire sig0000086d;
  wire sig0000086e;
  wire sig0000086f;
  wire sig00000870;
  wire sig00000871;
  wire sig00000872;
  wire sig00000873;
  wire sig00000874;
  wire sig00000875;
  wire sig00000876;
  wire sig00000877;
  wire sig00000878;
  wire sig00000879;
  wire sig0000087a;
  wire sig0000087b;
  wire sig0000087c;
  wire sig0000087d;
  wire sig0000087e;
  wire sig0000087f;
  wire sig00000880;
  wire sig00000881;
  wire sig00000882;
  wire sig00000883;
  wire sig00000884;
  wire sig00000885;
  wire sig00000886;
  wire sig00000887;
  wire sig00000888;
  wire sig00000889;
  wire sig0000088a;
  wire sig0000088b;
  wire sig0000088c;
  wire sig0000088d;
  wire sig0000088e;
  wire sig0000088f;
  wire sig00000890;
  wire sig00000891;
  wire sig00000892;
  wire sig00000893;
  wire sig00000894;
  wire sig00000895;
  wire sig00000896;
  wire sig00000897;
  wire sig00000898;
  wire sig00000899;
  wire sig0000089a;
  wire sig0000089b;
  wire sig0000089c;
  wire sig0000089d;
  wire sig0000089e;
  wire sig0000089f;
  wire sig000008a0;
  wire sig000008a1;
  wire sig000008a2;
  wire sig000008a3;
  wire sig000008a4;
  wire sig000008a5;
  wire sig000008a6;
  wire sig000008a7;
  wire sig000008a8;
  wire sig000008a9;
  wire sig000008aa;
  wire sig000008ab;
  wire sig000008ac;
  wire sig000008ad;
  wire sig000008ae;
  wire sig000008af;
  wire sig000008b0;
  wire sig000008b1;
  wire sig000008b2;
  wire sig000008b3;
  wire sig000008b4;
  wire sig000008b5;
  wire sig000008b6;
  wire sig000008b7;
  wire sig000008b8;
  wire sig000008b9;
  wire sig000008ba;
  wire sig000008bb;
  wire sig000008bc;
  wire sig000008bd;
  wire sig000008be;
  wire sig000008bf;
  wire sig000008c0;
  wire sig000008c1;
  wire sig000008c2;
  wire sig000008c3;
  wire sig000008c4;
  wire sig000008c5;
  wire sig000008c6;
  wire sig000008c7;
  wire sig000008c8;
  wire sig000008c9;
  wire sig000008ca;
  wire sig000008cb;
  wire sig000008cc;
  wire sig000008cd;
  wire sig000008ce;
  wire sig000008cf;
  wire sig000008d0;
  wire sig000008d1;
  wire sig000008d2;
  wire sig000008d3;
  wire sig000008d4;
  wire sig000008d5;
  wire sig000008d6;
  wire sig000008d7;
  wire sig000008d8;
  wire sig000008d9;
  wire sig000008da;
  wire sig000008db;
  wire sig000008dc;
  wire sig000008dd;
  wire sig000008de;
  wire sig000008df;
  wire sig000008e0;
  wire sig000008e1;
  wire sig000008e2;
  wire sig000008e3;
  wire sig000008e4;
  wire sig000008e5;
  wire sig000008e6;
  wire sig000008e7;
  wire sig000008e8;
  wire sig000008e9;
  wire sig000008ea;
  wire sig000008eb;
  wire sig000008ec;
  wire sig000008ed;
  wire sig000008ee;
  wire sig000008ef;
  wire sig000008f0;
  wire sig000008f1;
  wire sig000008f2;
  wire sig000008f3;
  wire sig000008f4;
  wire sig000008f5;
  wire sig000008f6;
  wire sig000008f7;
  wire sig000008f8;
  wire sig000008f9;
  wire sig000008fa;
  wire sig000008fb;
  wire sig000008fc;
  wire sig000008fd;
  wire sig000008fe;
  wire sig000008ff;
  wire sig00000900;
  wire sig00000901;
  wire sig00000902;
  wire sig00000903;
  wire sig00000904;
  wire sig00000905;
  wire sig00000906;
  wire sig00000907;
  wire sig00000908;
  wire sig00000909;
  wire sig0000090a;
  wire sig0000090b;
  wire sig0000090c;
  wire sig0000090d;
  wire sig0000090e;
  wire sig0000090f;
  wire sig00000910;
  wire sig00000911;
  wire sig00000912;
  wire sig00000913;
  wire sig00000914;
  wire sig00000915;
  wire sig00000916;
  wire sig00000917;
  wire sig00000918;
  wire sig00000919;
  wire sig0000091a;
  wire sig0000091b;
  wire sig0000091c;
  wire sig0000091d;
  wire sig0000091e;
  wire sig0000091f;
  wire sig00000920;
  wire sig00000921;
  wire sig00000922;
  wire sig00000923;
  wire sig00000924;
  wire sig00000925;
  wire sig00000926;
  wire sig00000927;
  wire sig00000928;
  wire sig00000929;
  wire sig0000092a;
  wire sig0000092b;
  wire sig0000092c;
  wire sig0000092d;
  wire sig0000092e;
  wire sig0000092f;
  wire sig00000930;
  wire sig00000931;
  wire sig00000932;
  wire sig00000933;
  wire sig00000934;
  wire sig00000935;
  wire sig00000936;
  wire sig00000937;
  wire sig00000938;
  wire sig00000939;
  wire sig0000093a;
  wire sig0000093b;
  wire sig0000093c;
  wire sig0000093d;
  wire sig0000093e;
  wire sig0000093f;
  wire sig00000940;
  wire sig00000941;
  wire sig00000942;
  wire sig00000943;
  wire sig00000944;
  wire sig00000945;
  wire sig00000946;
  wire sig00000947;
  wire sig00000948;
  wire sig00000949;
  wire sig0000094a;
  wire sig0000094b;
  wire sig0000094c;
  wire sig0000094d;
  wire sig0000094e;
  wire sig0000094f;
  wire sig00000950;
  wire sig00000951;
  wire sig00000952;
  wire sig00000953;
  wire sig00000954;
  wire sig00000955;
  wire sig00000956;
  wire sig00000957;
  wire sig00000958;
  wire sig00000959;
  wire sig0000095a;
  wire sig0000095b;
  wire sig0000095c;
  wire sig0000095d;
  wire sig0000095e;
  wire sig0000095f;
  wire sig00000960;
  wire sig00000961;
  wire sig00000962;
  wire sig00000963;
  wire sig00000964;
  wire sig00000965;
  wire sig00000966;
  wire sig00000967;
  wire sig00000968;
  wire sig00000969;
  wire sig0000096a;
  wire sig0000096b;
  wire sig0000096c;
  wire sig0000096d;
  wire sig0000096e;
  wire sig0000096f;
  wire sig00000970;
  wire sig00000971;
  wire sig00000972;
  wire sig00000973;
  wire sig00000974;
  wire sig00000975;
  wire sig00000976;
  wire sig00000977;
  wire sig00000978;
  wire sig00000979;
  wire sig0000097a;
  wire sig0000097b;
  wire sig0000097c;
  wire sig0000097d;
  wire sig0000097e;
  wire sig0000097f;
  wire sig00000980;
  wire sig00000981;
  wire sig00000982;
  wire sig00000983;
  wire sig00000984;
  wire sig00000985;
  wire sig00000986;
  wire sig00000987;
  wire sig00000988;
  wire sig00000989;
  wire sig0000098a;
  wire sig0000098b;
  wire sig0000098c;
  wire sig0000098d;
  wire sig0000098e;
  wire sig0000098f;
  wire sig00000990;
  wire sig00000991;
  wire sig00000992;
  wire sig00000993;
  wire sig00000994;
  wire sig00000995;
  wire sig00000996;
  wire sig00000997;
  wire sig00000998;
  wire sig00000999;
  wire \NlwRenamedSig_OI_U0/i_synth/non_floating_point.arch_c.xfft_inst/control/cntrl/process_state_r ;
  wire sig0000099a;
  wire sig0000099b;
  wire sig0000099c;
  wire sig0000099d;
  wire sig0000099e;
  wire sig0000099f;
  wire sig000009a0;
  wire sig000009a1;
  wire sig000009a2;
  wire sig000009a3;
  wire sig000009a4;
  wire sig000009a5;
  wire sig000009a6;
  wire sig000009a7;
  wire sig000009a8;
  wire sig000009a9;
  wire sig000009aa;
  wire sig000009ab;
  wire sig000009ac;
  wire sig000009ad;
  wire sig000009ae;
  wire sig000009af;
  wire sig000009b0;
  wire sig000009b1;
  wire sig000009b2;
  wire sig000009b3;
  wire sig000009b4;
  wire sig000009b5;
  wire sig000009b6;
  wire sig000009b7;
  wire sig000009b8;
  wire sig000009b9;
  wire sig000009ba;
  wire sig000009bb;
  wire sig000009bc;
  wire sig000009bd;
  wire sig000009be;
  wire sig000009bf;
  wire sig000009c0;
  wire sig000009c1;
  wire sig000009c2;
  wire sig000009c3;
  wire sig000009c4;
  wire sig000009c5;
  wire sig000009c6;
  wire sig000009c7;
  wire sig000009c8;
  wire sig000009c9;
  wire sig000009ca;
  wire sig000009cb;
  wire sig000009cc;
  wire sig000009cd;
  wire sig000009ce;
  wire sig000009cf;
  wire sig000009d0;
  wire sig000009d1;
  wire sig000009d2;
  wire sig000009d3;
  wire sig000009d4;
  wire sig000009d5;
  wire sig000009d6;
  wire sig000009d7;
  wire sig000009d8;
  wire sig000009d9;
  wire sig000009da;
  wire sig000009db;
  wire sig000009dc;
  wire sig000009dd;
  wire sig000009de;
  wire sig000009df;
  wire sig000009e0;
  wire sig000009e1;
  wire sig000009e2;
  wire sig000009e3;
  wire sig000009e4;
  wire sig000009e5;
  wire sig000009e6;
  wire sig000009e7;
  wire sig000009e8;
  wire sig000009e9;
  wire sig000009ea;
  wire sig000009eb;
  wire sig000009ec;
  wire sig000009ed;
  wire sig000009ee;
  wire sig000009ef;
  wire sig000009f0;
  wire sig000009f1;
  wire sig000009f2;
  wire sig000009f3;
  wire sig000009f4;
  wire sig000009f5;
  wire sig000009f6;
  wire sig000009f7;
  wire sig000009f8;
  wire sig000009f9;
  wire sig000009fa;
  wire sig000009fb;
  wire sig000009fc;
  wire sig000009fd;
  wire sig000009fe;
  wire sig000009ff;
  wire sig00000a00;
  wire sig00000a01;
  wire sig00000a02;
  wire sig00000a03;
  wire sig00000a04;
  wire sig00000a05;
  wire sig00000a06;
  wire sig00000a07;
  wire sig00000a08;
  wire sig00000a09;
  wire sig00000a0a;
  wire sig00000a0b;
  wire sig00000a0c;
  wire sig00000a0d;
  wire sig00000a0e;
  wire sig00000a0f;
  wire sig00000a10;
  wire sig00000a11;
  wire sig00000a12;
  wire sig00000a13;
  wire sig00000a14;
  wire sig00000a15;
  wire sig00000a16;
  wire sig00000a17;
  wire sig00000a18;
  wire sig00000a19;
  wire sig00000a1a;
  wire sig00000a1b;
  wire sig00000a1c;
  wire sig00000a1d;
  wire sig00000a1e;
  wire sig00000a1f;
  wire sig00000a20;
  wire sig00000a21;
  wire sig00000a22;
  wire sig00000a23;
  wire sig00000a24;
  wire sig00000a25;
  wire sig00000a26;
  wire sig00000a27;
  wire sig00000a28;
  wire sig00000a29;
  wire sig00000a2a;
  wire sig00000a2b;
  wire sig00000a2c;
  wire sig00000a2d;
  wire sig00000a2e;
  wire sig00000a2f;
  wire sig00000a30;
  wire sig00000a31;
  wire sig00000a32;
  wire sig00000a33;
  wire sig00000a34;
  wire sig00000a35;
  wire sig00000a36;
  wire sig00000a37;
  wire sig00000a38;
  wire sig00000a39;
  wire sig00000a3a;
  wire sig00000a3b;
  wire sig00000a3c;
  wire sig00000a3d;
  wire sig00000a3e;
  wire sig00000a3f;
  wire sig00000a40;
  wire sig00000a41;
  wire sig00000a42;
  wire sig00000a43;
  wire sig00000a44;
  wire sig00000a45;
  wire sig00000a46;
  wire \blk00000003/sig00000acd ;
  wire \blk00000003/sig00000aa6 ;
  wire \blk00000003/sig00000aa5 ;
  wire \blk00000003/sig00000aa4 ;
  wire \blk00000003/sig00000aa3 ;
  wire \blk00000003/sig00000aa2 ;
  wire \blk00000003/sig00000aa1 ;
  wire \blk00000003/sig00000aa0 ;
  wire \blk00000003/sig00000a9f ;
  wire \blk00000003/sig00000a9e ;
  wire \blk00000003/sig00000a9d ;
  wire \blk00000003/sig00000a9c ;
  wire \blk00000003/sig00000a9b ;
  wire \blk00000003/sig00000a9a ;
  wire \blk00000003/sig00000a99 ;
  wire \blk00000003/sig00000a98 ;
  wire \blk00000003/sig00000a97 ;
  wire \blk00000003/sig00000a96 ;
  wire \blk00000003/sig00000a95 ;
  wire \blk00000003/sig00000a94 ;
  wire \blk00000003/sig00000a93 ;
  wire \blk00000003/sig00000a92 ;
  wire \blk00000003/sig00000a91 ;
  wire \blk00000003/sig00000a90 ;
  wire \blk00000003/sig00000a8f ;
  wire \blk00000003/sig00000a8e ;
  wire \blk00000003/sig00000a8d ;
  wire \blk00000003/sig00000a8c ;
  wire \blk00000003/sig00000a8b ;
  wire \blk00000003/sig00000a8a ;
  wire \blk00000003/sig00000a89 ;
  wire \blk00000003/sig00000a88 ;
  wire \blk00000003/sig00000a87 ;
  wire \blk00000003/sig00000a86 ;
  wire \blk00000003/sig00000a85 ;
  wire \blk00000003/sig00000a84 ;
  wire \blk00000003/sig00000a83 ;
  wire \blk00000003/sig00000a82 ;
  wire \blk00000003/sig00000a81 ;
  wire \blk0000002d/sig00000b54 ;
  wire \blk0000002d/sig00000b2d ;
  wire \blk0000002d/sig00000b2c ;
  wire \blk0000002d/sig00000b2b ;
  wire \blk0000002d/sig00000b2a ;
  wire \blk0000002d/sig00000b29 ;
  wire \blk0000002d/sig00000b28 ;
  wire \blk0000002d/sig00000b27 ;
  wire \blk0000002d/sig00000b26 ;
  wire \blk0000002d/sig00000b25 ;
  wire \blk0000002d/sig00000b24 ;
  wire \blk0000002d/sig00000b23 ;
  wire \blk0000002d/sig00000b22 ;
  wire \blk0000002d/sig00000b21 ;
  wire \blk0000002d/sig00000b20 ;
  wire \blk0000002d/sig00000b1f ;
  wire \blk0000002d/sig00000b1e ;
  wire \blk0000002d/sig00000b1d ;
  wire \blk0000002d/sig00000b1c ;
  wire \blk0000002d/sig00000b1b ;
  wire \blk0000002d/sig00000b1a ;
  wire \blk0000002d/sig00000b19 ;
  wire \blk0000002d/sig00000b18 ;
  wire \blk0000002d/sig00000b17 ;
  wire \blk0000002d/sig00000b16 ;
  wire \blk0000002d/sig00000b15 ;
  wire \blk0000002d/sig00000b14 ;
  wire \blk0000002d/sig00000b13 ;
  wire \blk0000002d/sig00000b12 ;
  wire \blk0000002d/sig00000b11 ;
  wire \blk0000002d/sig00000b10 ;
  wire \blk0000002d/sig00000b0f ;
  wire \blk0000002d/sig00000b0e ;
  wire \blk0000002d/sig00000b0d ;
  wire \blk0000002d/sig00000b0c ;
  wire \blk0000002d/sig00000b0b ;
  wire \blk0000002d/sig00000b0a ;
  wire \blk0000002d/sig00000b09 ;
  wire \blk0000002d/sig00000b08 ;
  wire \blk0000018c/sig00000bcc ;
  wire \blk0000018c/sig00000bcb ;
  wire \blk0000018c/sig00000bca ;
  wire \blk0000018c/sig00000bc9 ;
  wire \blk00000194/sig00000bd8 ;
  wire \blk00000194/sig00000bd7 ;
  wire \blk00000194/sig00000bd6 ;
  wire \blk00000194/sig00000bd5 ;
  wire \blk0000019d/sig00000c00 ;
  wire \blk0000019d/sig00000bff ;
  wire \blk0000019d/sig00000bfe ;
  wire \blk0000019d/sig00000bfd ;
  wire \blk0000019d/sig00000bfc ;
  wire \blk0000019d/sig00000bfb ;
  wire \blk0000019d/sig00000bfa ;
  wire \blk0000019d/sig00000bf9 ;
  wire \blk0000019d/sig00000bf8 ;
  wire \blk0000019d/sig00000bf7 ;
  wire \blk0000019d/sig00000bf6 ;
  wire \blk0000019d/sig00000bf5 ;
  wire \blk0000019d/sig00000bf4 ;
  wire \blk000001b7/sig00000c27 ;
  wire \blk000001b7/sig00000c26 ;
  wire \blk000001b7/sig00000c25 ;
  wire \blk000001b7/sig00000c24 ;
  wire \blk000001b7/sig00000c23 ;
  wire \blk000001b7/sig00000c22 ;
  wire \blk000001b7/sig00000c21 ;
  wire \blk000001b7/sig00000c20 ;
  wire \blk000001b7/sig00000c1f ;
  wire \blk000001b7/sig00000c1e ;
  wire \blk000001b7/sig00000c1d ;
  wire \blk000001b7/sig00000c1c ;
  wire \blk000001b7/sig00000c1b ;
  wire \blk000001d1/sig00000c5d ;
  wire \blk000001d1/sig00000c5c ;
  wire \blk000001d1/sig00000c5b ;
  wire \blk000001d1/sig00000c5a ;
  wire \blk000001d1/sig00000c59 ;
  wire \blk000001d1/sig00000c58 ;
  wire \blk000001d1/sig00000c57 ;
  wire \blk000001d1/sig00000c56 ;
  wire \blk000001d1/sig00000c55 ;
  wire \blk000001d1/sig00000c54 ;
  wire \blk000001d1/sig00000c53 ;
  wire \blk000001d1/sig00000c52 ;
  wire \blk000001d1/sig00000c51 ;
  wire \blk000001d1/sig00000c50 ;
  wire \blk000001d1/sig00000c4f ;
  wire \blk000001d1/sig00000c4e ;
  wire \blk000001d1/sig00000c4d ;
  wire \blk000001d1/sig00000c4c ;
  wire \blk000001f8/sig00000cd2 ;
  wire \blk000001f8/sig00000cd1 ;
  wire \blk000001f8/sig00000cd0 ;
  wire \blk000001fe/sig00000d5e ;
  wire \blk000001fe/sig00000d5d ;
  wire \blk000001fe/sig00000d5c ;
  wire \blk000001fe/sig00000d5b ;
  wire \blk000001fe/sig00000d5a ;
  wire \blk000001fe/sig00000d59 ;
  wire \blk000001fe/sig00000d58 ;
  wire \blk000001fe/sig00000d57 ;
  wire \blk000001fe/sig00000d56 ;
  wire \blk000001fe/sig00000d55 ;
  wire \blk000001fe/sig00000d54 ;
  wire \blk000001fe/sig00000d53 ;
  wire \blk000001fe/sig00000d52 ;
  wire \blk000001fe/sig00000d51 ;
  wire \blk000001fe/sig00000d50 ;
  wire \blk000001fe/sig00000d4f ;
  wire \blk000001fe/sig00000d4e ;
  wire \blk000001fe/sig00000d4d ;
  wire \blk000001fe/sig00000d4c ;
  wire \blk000001fe/sig00000d4b ;
  wire \blk000001fe/sig00000d4a ;
  wire \blk000001fe/sig00000d49 ;
  wire \blk000001fe/sig00000d48 ;
  wire \blk000001fe/sig00000d47 ;
  wire \blk000001fe/sig00000d46 ;
  wire \blk000001fe/sig00000d45 ;
  wire \blk000001fe/sig00000d44 ;
  wire \blk000001fe/sig00000d43 ;
  wire \blk000001fe/sig00000d42 ;
  wire \blk000001fe/sig00000d41 ;
  wire \blk000001fe/sig00000d40 ;
  wire \blk000001fe/sig00000d3f ;
  wire \blk000001fe/sig00000d3e ;
  wire \blk000001fe/sig00000d3d ;
  wire \blk000001fe/sig00000d3c ;
  wire \blk000001fe/sig00000d3b ;
  wire \blk000001fe/sig00000d3a ;
  wire \blk000001fe/sig00000d39 ;
  wire \blk000001fe/sig00000d38 ;
  wire \blk000001fe/sig00000d37 ;
  wire \blk000001fe/sig00000d36 ;
  wire \blk000001fe/sig00000d35 ;
  wire \blk000001fe/sig00000d34 ;
  wire \blk000001fe/sig00000d33 ;
  wire \blk000001fe/sig00000d32 ;
  wire \blk000001fe/sig00000d31 ;
  wire \blk000001fe/sig00000d30 ;
  wire \blk000001fe/sig00000d2f ;
  wire \blk000001fe/sig00000d2e ;
  wire \blk000001fe/sig00000d2d ;
  wire \blk000001fe/sig00000d2c ;
  wire \blk000001fe/sig00000d2b ;
  wire \blk000001fe/sig00000d2a ;
  wire \blk000001fe/sig00000d29 ;
  wire \blk000001fe/sig00000d28 ;
  wire \blk000001fe/sig00000d27 ;
  wire \blk000001fe/sig00000d26 ;
  wire \blk000001fe/sig00000d25 ;
  wire \blk000001fe/sig00000d24 ;
  wire \blk000001fe/sig00000d23 ;
  wire \blk000001fe/sig00000d22 ;
  wire \blk000001fe/sig00000d21 ;
  wire \blk000001fe/sig00000d20 ;
  wire \blk000001fe/sig00000d1f ;
  wire \blk000001fe/sig00000d1e ;
  wire \blk000001fe/sig00000d1d ;
  wire \blk000001fe/sig00000d1c ;
  wire \blk000001fe/sig00000d1b ;
  wire \blk000001fe/sig00000d1a ;
  wire \blk000001fe/sig00000d19 ;
  wire \blk0000025d/sig00000dea ;
  wire \blk0000025d/sig00000de9 ;
  wire \blk0000025d/sig00000de8 ;
  wire \blk0000025d/sig00000de7 ;
  wire \blk0000025d/sig00000de6 ;
  wire \blk0000025d/sig00000de5 ;
  wire \blk0000025d/sig00000de4 ;
  wire \blk0000025d/sig00000de3 ;
  wire \blk0000025d/sig00000de2 ;
  wire \blk0000025d/sig00000de1 ;
  wire \blk0000025d/sig00000de0 ;
  wire \blk0000025d/sig00000ddf ;
  wire \blk0000025d/sig00000dde ;
  wire \blk0000025d/sig00000ddd ;
  wire \blk0000025d/sig00000ddc ;
  wire \blk0000025d/sig00000ddb ;
  wire \blk0000025d/sig00000dda ;
  wire \blk0000025d/sig00000dd9 ;
  wire \blk0000025d/sig00000dd8 ;
  wire \blk0000025d/sig00000dd7 ;
  wire \blk0000025d/sig00000dd6 ;
  wire \blk0000025d/sig00000dd5 ;
  wire \blk0000025d/sig00000dd4 ;
  wire \blk0000025d/sig00000dd3 ;
  wire \blk0000025d/sig00000dd2 ;
  wire \blk0000025d/sig00000dd1 ;
  wire \blk0000025d/sig00000dd0 ;
  wire \blk0000025d/sig00000dcf ;
  wire \blk0000025d/sig00000dce ;
  wire \blk0000025d/sig00000dcd ;
  wire \blk0000025d/sig00000dcc ;
  wire \blk0000025d/sig00000dcb ;
  wire \blk0000025d/sig00000dca ;
  wire \blk0000025d/sig00000dc9 ;
  wire \blk0000025d/sig00000dc8 ;
  wire \blk0000025d/sig00000dc7 ;
  wire \blk0000025d/sig00000dc6 ;
  wire \blk0000025d/sig00000dc5 ;
  wire \blk0000025d/sig00000dc4 ;
  wire \blk0000025d/sig00000dc3 ;
  wire \blk0000025d/sig00000dc2 ;
  wire \blk0000025d/sig00000dc1 ;
  wire \blk0000025d/sig00000dc0 ;
  wire \blk0000025d/sig00000dbf ;
  wire \blk0000025d/sig00000dbe ;
  wire \blk0000025d/sig00000dbd ;
  wire \blk0000025d/sig00000dbc ;
  wire \blk0000025d/sig00000dbb ;
  wire \blk0000025d/sig00000dba ;
  wire \blk0000025d/sig00000db9 ;
  wire \blk0000025d/sig00000db8 ;
  wire \blk0000025d/sig00000db7 ;
  wire \blk0000025d/sig00000db6 ;
  wire \blk0000025d/sig00000db5 ;
  wire \blk0000025d/sig00000db4 ;
  wire \blk0000025d/sig00000db3 ;
  wire \blk0000025d/sig00000db2 ;
  wire \blk0000025d/sig00000db1 ;
  wire \blk0000025d/sig00000db0 ;
  wire \blk0000025d/sig00000daf ;
  wire \blk0000025d/sig00000dae ;
  wire \blk0000025d/sig00000dad ;
  wire \blk0000025d/sig00000dac ;
  wire \blk0000025d/sig00000dab ;
  wire \blk0000025d/sig00000daa ;
  wire \blk0000025d/sig00000da9 ;
  wire \blk0000025d/sig00000da8 ;
  wire \blk0000025d/sig00000da7 ;
  wire \blk0000025d/sig00000da6 ;
  wire \blk0000025d/sig00000da5 ;
  wire \blk000002bc/sig00000e76 ;
  wire \blk000002bc/sig00000e75 ;
  wire \blk000002bc/sig00000e74 ;
  wire \blk000002bc/sig00000e73 ;
  wire \blk000002bc/sig00000e72 ;
  wire \blk000002bc/sig00000e71 ;
  wire \blk000002bc/sig00000e70 ;
  wire \blk000002bc/sig00000e6f ;
  wire \blk000002bc/sig00000e6e ;
  wire \blk000002bc/sig00000e6d ;
  wire \blk000002bc/sig00000e6c ;
  wire \blk000002bc/sig00000e6b ;
  wire \blk000002bc/sig00000e6a ;
  wire \blk000002bc/sig00000e69 ;
  wire \blk000002bc/sig00000e68 ;
  wire \blk000002bc/sig00000e67 ;
  wire \blk000002bc/sig00000e66 ;
  wire \blk000002bc/sig00000e65 ;
  wire \blk000002bc/sig00000e64 ;
  wire \blk000002bc/sig00000e63 ;
  wire \blk000002bc/sig00000e62 ;
  wire \blk000002bc/sig00000e61 ;
  wire \blk000002bc/sig00000e60 ;
  wire \blk000002bc/sig00000e5f ;
  wire \blk000002bc/sig00000e5e ;
  wire \blk000002bc/sig00000e5d ;
  wire \blk000002bc/sig00000e5c ;
  wire \blk000002bc/sig00000e5b ;
  wire \blk000002bc/sig00000e5a ;
  wire \blk000002bc/sig00000e59 ;
  wire \blk000002bc/sig00000e58 ;
  wire \blk000002bc/sig00000e57 ;
  wire \blk000002bc/sig00000e56 ;
  wire \blk000002bc/sig00000e55 ;
  wire \blk000002bc/sig00000e54 ;
  wire \blk000002bc/sig00000e53 ;
  wire \blk000002bc/sig00000e52 ;
  wire \blk000002bc/sig00000e51 ;
  wire \blk000002bc/sig00000e50 ;
  wire \blk000002bc/sig00000e4f ;
  wire \blk000002bc/sig00000e4e ;
  wire \blk000002bc/sig00000e4d ;
  wire \blk000002bc/sig00000e4c ;
  wire \blk000002bc/sig00000e4b ;
  wire \blk000002bc/sig00000e4a ;
  wire \blk000002bc/sig00000e49 ;
  wire \blk000002bc/sig00000e48 ;
  wire \blk000002bc/sig00000e47 ;
  wire \blk000002bc/sig00000e46 ;
  wire \blk000002bc/sig00000e45 ;
  wire \blk000002bc/sig00000e44 ;
  wire \blk000002bc/sig00000e43 ;
  wire \blk000002bc/sig00000e42 ;
  wire \blk000002bc/sig00000e41 ;
  wire \blk000002bc/sig00000e40 ;
  wire \blk000002bc/sig00000e3f ;
  wire \blk000002bc/sig00000e3e ;
  wire \blk000002bc/sig00000e3d ;
  wire \blk000002bc/sig00000e3c ;
  wire \blk000002bc/sig00000e3b ;
  wire \blk000002bc/sig00000e3a ;
  wire \blk000002bc/sig00000e39 ;
  wire \blk000002bc/sig00000e38 ;
  wire \blk000002bc/sig00000e37 ;
  wire \blk000002bc/sig00000e36 ;
  wire \blk000002bc/sig00000e35 ;
  wire \blk000002bc/sig00000e34 ;
  wire \blk000002bc/sig00000e33 ;
  wire \blk000002bc/sig00000e32 ;
  wire \blk000002bc/sig00000e31 ;
  wire \blk0000031b/sig00000f02 ;
  wire \blk0000031b/sig00000f01 ;
  wire \blk0000031b/sig00000f00 ;
  wire \blk0000031b/sig00000eff ;
  wire \blk0000031b/sig00000efe ;
  wire \blk0000031b/sig00000efd ;
  wire \blk0000031b/sig00000efc ;
  wire \blk0000031b/sig00000efb ;
  wire \blk0000031b/sig00000efa ;
  wire \blk0000031b/sig00000ef9 ;
  wire \blk0000031b/sig00000ef8 ;
  wire \blk0000031b/sig00000ef7 ;
  wire \blk0000031b/sig00000ef6 ;
  wire \blk0000031b/sig00000ef5 ;
  wire \blk0000031b/sig00000ef4 ;
  wire \blk0000031b/sig00000ef3 ;
  wire \blk0000031b/sig00000ef2 ;
  wire \blk0000031b/sig00000ef1 ;
  wire \blk0000031b/sig00000ef0 ;
  wire \blk0000031b/sig00000eef ;
  wire \blk0000031b/sig00000eee ;
  wire \blk0000031b/sig00000eed ;
  wire \blk0000031b/sig00000eec ;
  wire \blk0000031b/sig00000eeb ;
  wire \blk0000031b/sig00000eea ;
  wire \blk0000031b/sig00000ee9 ;
  wire \blk0000031b/sig00000ee8 ;
  wire \blk0000031b/sig00000ee7 ;
  wire \blk0000031b/sig00000ee6 ;
  wire \blk0000031b/sig00000ee5 ;
  wire \blk0000031b/sig00000ee4 ;
  wire \blk0000031b/sig00000ee3 ;
  wire \blk0000031b/sig00000ee2 ;
  wire \blk0000031b/sig00000ee1 ;
  wire \blk0000031b/sig00000ee0 ;
  wire \blk0000031b/sig00000edf ;
  wire \blk0000031b/sig00000ede ;
  wire \blk0000031b/sig00000edd ;
  wire \blk0000031b/sig00000edc ;
  wire \blk0000031b/sig00000edb ;
  wire \blk0000031b/sig00000eda ;
  wire \blk0000031b/sig00000ed9 ;
  wire \blk0000031b/sig00000ed8 ;
  wire \blk0000031b/sig00000ed7 ;
  wire \blk0000031b/sig00000ed6 ;
  wire \blk0000031b/sig00000ed5 ;
  wire \blk0000031b/sig00000ed4 ;
  wire \blk0000031b/sig00000ed3 ;
  wire \blk0000031b/sig00000ed2 ;
  wire \blk0000031b/sig00000ed1 ;
  wire \blk0000031b/sig00000ed0 ;
  wire \blk0000031b/sig00000ecf ;
  wire \blk0000031b/sig00000ece ;
  wire \blk0000031b/sig00000ecd ;
  wire \blk0000031b/sig00000ecc ;
  wire \blk0000031b/sig00000ecb ;
  wire \blk0000031b/sig00000eca ;
  wire \blk0000031b/sig00000ec9 ;
  wire \blk0000031b/sig00000ec8 ;
  wire \blk0000031b/sig00000ec7 ;
  wire \blk0000031b/sig00000ec6 ;
  wire \blk0000031b/sig00000ec5 ;
  wire \blk0000031b/sig00000ec4 ;
  wire \blk0000031b/sig00000ec3 ;
  wire \blk0000031b/sig00000ec2 ;
  wire \blk0000031b/sig00000ec1 ;
  wire \blk0000031b/sig00000ec0 ;
  wire \blk0000031b/sig00000ebf ;
  wire \blk0000031b/sig00000ebe ;
  wire \blk0000031b/sig00000ebd ;
  wire \blk0000049e/sig00000f4e ;
  wire \blk0000049e/sig00000f4d ;
  wire \blk0000049e/sig00000f4c ;
  wire \blk0000049e/sig00000f4b ;
  wire \blk0000049e/sig00000f4a ;
  wire \blk0000049e/sig00000f49 ;
  wire \blk0000049e/sig00000f48 ;
  wire \blk0000049e/sig00000f47 ;
  wire \blk0000049e/sig00000f46 ;
  wire \blk0000049e/sig00000f45 ;
  wire \blk0000049e/sig00000f44 ;
  wire \blk0000049e/sig00000f43 ;
  wire \blk0000049e/sig00000f42 ;
  wire \blk0000049e/sig00000f41 ;
  wire \blk0000049e/sig00000f40 ;
  wire \blk0000049e/sig00000f3f ;
  wire \blk0000049e/sig00000f3e ;
  wire \blk0000049e/sig00000f3d ;
  wire \blk0000049e/sig00000f3c ;
  wire \blk0000049e/sig00000f3b ;
  wire \blk0000049e/sig00000f3a ;
  wire \blk0000049e/sig00000f39 ;
  wire \blk0000049e/sig00000f38 ;
  wire \blk0000049e/sig00000f37 ;
  wire \blk0000049e/sig00000f36 ;
  wire \blk0000049e/sig00000f35 ;
  wire \blk0000049e/sig00000f34 ;
  wire \blk0000049e/sig00000f33 ;
  wire \blk0000049e/sig00000f32 ;
  wire \blk0000049e/sig00000f31 ;
  wire \blk0000049e/sig00000f30 ;
  wire \blk0000049e/sig00000f2f ;
  wire \blk0000049e/sig00000f2e ;
  wire \blk0000049e/sig00000f2d ;
  wire \blk0000049e/sig00000f2c ;
  wire \blk0000049e/sig00000f2b ;
  wire \blk0000049e/sig00000f2a ;
  wire \blk000004d7/sig00000f9a ;
  wire \blk000004d7/sig00000f99 ;
  wire \blk000004d7/sig00000f98 ;
  wire \blk000004d7/sig00000f97 ;
  wire \blk000004d7/sig00000f96 ;
  wire \blk000004d7/sig00000f95 ;
  wire \blk000004d7/sig00000f94 ;
  wire \blk000004d7/sig00000f93 ;
  wire \blk000004d7/sig00000f92 ;
  wire \blk000004d7/sig00000f91 ;
  wire \blk000004d7/sig00000f90 ;
  wire \blk000004d7/sig00000f8f ;
  wire \blk000004d7/sig00000f8e ;
  wire \blk000004d7/sig00000f8d ;
  wire \blk000004d7/sig00000f8c ;
  wire \blk000004d7/sig00000f8b ;
  wire \blk000004d7/sig00000f8a ;
  wire \blk000004d7/sig00000f89 ;
  wire \blk000004d7/sig00000f88 ;
  wire \blk000004d7/sig00000f87 ;
  wire \blk000004d7/sig00000f86 ;
  wire \blk000004d7/sig00000f85 ;
  wire \blk000004d7/sig00000f84 ;
  wire \blk000004d7/sig00000f83 ;
  wire \blk000004d7/sig00000f82 ;
  wire \blk000004d7/sig00000f81 ;
  wire \blk000004d7/sig00000f80 ;
  wire \blk000004d7/sig00000f7f ;
  wire \blk000004d7/sig00000f7e ;
  wire \blk000004d7/sig00000f7d ;
  wire \blk000004d7/sig00000f7c ;
  wire \blk000004d7/sig00000f7b ;
  wire \blk000004d7/sig00000f7a ;
  wire \blk000004d7/sig00000f79 ;
  wire \blk000004d7/sig00000f78 ;
  wire \blk000004d7/sig00000f77 ;
  wire \blk000004d7/sig00000f76 ;
  wire \blk00000510/sig00000fe6 ;
  wire \blk00000510/sig00000fe5 ;
  wire \blk00000510/sig00000fe4 ;
  wire \blk00000510/sig00000fe3 ;
  wire \blk00000510/sig00000fe2 ;
  wire \blk00000510/sig00000fe1 ;
  wire \blk00000510/sig00000fe0 ;
  wire \blk00000510/sig00000fdf ;
  wire \blk00000510/sig00000fde ;
  wire \blk00000510/sig00000fdd ;
  wire \blk00000510/sig00000fdc ;
  wire \blk00000510/sig00000fdb ;
  wire \blk00000510/sig00000fda ;
  wire \blk00000510/sig00000fd9 ;
  wire \blk00000510/sig00000fd8 ;
  wire \blk00000510/sig00000fd7 ;
  wire \blk00000510/sig00000fd6 ;
  wire \blk00000510/sig00000fd5 ;
  wire \blk00000510/sig00000fd4 ;
  wire \blk00000510/sig00000fd3 ;
  wire \blk00000510/sig00000fd2 ;
  wire \blk00000510/sig00000fd1 ;
  wire \blk00000510/sig00000fd0 ;
  wire \blk00000510/sig00000fcf ;
  wire \blk00000510/sig00000fce ;
  wire \blk00000510/sig00000fcd ;
  wire \blk00000510/sig00000fcc ;
  wire \blk00000510/sig00000fcb ;
  wire \blk00000510/sig00000fca ;
  wire \blk00000510/sig00000fc9 ;
  wire \blk00000510/sig00000fc8 ;
  wire \blk00000510/sig00000fc7 ;
  wire \blk00000510/sig00000fc6 ;
  wire \blk00000510/sig00000fc5 ;
  wire \blk00000510/sig00000fc4 ;
  wire \blk00000510/sig00000fc3 ;
  wire \blk00000510/sig00000fc2 ;
  wire \blk00000549/sig00001032 ;
  wire \blk00000549/sig00001031 ;
  wire \blk00000549/sig00001030 ;
  wire \blk00000549/sig0000102f ;
  wire \blk00000549/sig0000102e ;
  wire \blk00000549/sig0000102d ;
  wire \blk00000549/sig0000102c ;
  wire \blk00000549/sig0000102b ;
  wire \blk00000549/sig0000102a ;
  wire \blk00000549/sig00001029 ;
  wire \blk00000549/sig00001028 ;
  wire \blk00000549/sig00001027 ;
  wire \blk00000549/sig00001026 ;
  wire \blk00000549/sig00001025 ;
  wire \blk00000549/sig00001024 ;
  wire \blk00000549/sig00001023 ;
  wire \blk00000549/sig00001022 ;
  wire \blk00000549/sig00001021 ;
  wire \blk00000549/sig00001020 ;
  wire \blk00000549/sig0000101f ;
  wire \blk00000549/sig0000101e ;
  wire \blk00000549/sig0000101d ;
  wire \blk00000549/sig0000101c ;
  wire \blk00000549/sig0000101b ;
  wire \blk00000549/sig0000101a ;
  wire \blk00000549/sig00001019 ;
  wire \blk00000549/sig00001018 ;
  wire \blk00000549/sig00001017 ;
  wire \blk00000549/sig00001016 ;
  wire \blk00000549/sig00001015 ;
  wire \blk00000549/sig00001014 ;
  wire \blk00000549/sig00001013 ;
  wire \blk00000549/sig00001012 ;
  wire \blk00000549/sig00001011 ;
  wire \blk00000549/sig00001010 ;
  wire \blk00000549/sig0000100f ;
  wire \blk00000549/sig0000100e ;
  wire \blk00000751/blk00000752/sig0000103e ;
  wire \blk00000751/blk00000752/sig0000103d ;
  wire \blk00000751/blk00000752/sig0000103c ;
  wire \blk00000757/blk00000758/sig0000104a ;
  wire \blk00000757/blk00000758/sig00001049 ;
  wire \blk00000757/blk00000758/sig00001048 ;
  wire \blk000007ea/blk000007eb/sig00001079 ;
  wire \blk000007ea/blk000007eb/sig00001078 ;
  wire \blk000007ea/blk000007eb/sig00001077 ;
  wire \blk000007ea/blk000007eb/sig00001076 ;
  wire \blk000007ea/blk000007eb/sig00001075 ;
  wire \blk000007ea/blk000007eb/sig00001074 ;
  wire \blk000007ea/blk000007eb/sig00001073 ;
  wire \blk000007ea/blk000007eb/sig00001072 ;
  wire \blk000007ea/blk000007eb/sig00001071 ;
  wire \blk000007ea/blk000007eb/sig00001070 ;
  wire \blk000007fe/blk000007ff/sig000010a8 ;
  wire \blk000007fe/blk000007ff/sig000010a7 ;
  wire \blk000007fe/blk000007ff/sig000010a6 ;
  wire \blk000007fe/blk000007ff/sig000010a5 ;
  wire \blk000007fe/blk000007ff/sig000010a4 ;
  wire \blk000007fe/blk000007ff/sig000010a3 ;
  wire \blk000007fe/blk000007ff/sig000010a2 ;
  wire \blk000007fe/blk000007ff/sig000010a1 ;
  wire \blk000007fe/blk000007ff/sig000010a0 ;
  wire \blk000007fe/blk000007ff/sig0000109f ;
  wire \blk00000852/blk00000853/sig000010bc ;
  wire \blk00000852/blk00000853/sig000010bb ;
  wire \blk00000852/blk00000853/sig000010ba ;
  wire \blk00000858/blk00000859/sig000010c8 ;
  wire \blk00000858/blk00000859/sig000010c7 ;
  wire \blk00000858/blk00000859/sig000010c6 ;
  wire \blk0000085e/blk0000085f/sig000010d4 ;
  wire \blk0000085e/blk0000085f/sig000010d3 ;
  wire \blk0000085e/blk0000085f/sig000010d2 ;
  wire \blk000008e1/blk000008e2/sig000010df ;
  wire \blk000008e1/blk000008e2/sig000010de ;
  wire \blk000008e6/blk000008e7/sig000010ea ;
  wire \blk000008e6/blk000008e7/sig000010e9 ;
  wire \blk00000935/sig0000110a ;
  wire \blk00000935/sig00001109 ;
  wire \blk00000935/sig00001108 ;
  wire \blk00000935/sig00001107 ;
  wire \blk00000935/sig00001106 ;
  wire \blk00000935/sig00001105 ;
  wire \blk00000935/sig00001104 ;
  wire \blk00000935/sig00001103 ;
  wire \blk00000935/sig00001102 ;
  wire \blk00000935/sig00001101 ;
  wire \blk00000935/sig00001100 ;
  wire \blk00000935/sig000010ff ;
  wire \blk00000935/sig000010fe ;
  wire \blk00000935/sig000010fd ;
  wire \blk00000935/sig000010fc ;
  wire \blk00000935/sig000010fb ;
  wire \blk0000095a/sig0000111e ;
  wire \blk0000095a/sig0000111d ;
  wire \blk0000095a/sig0000111c ;
  wire \blk0000095a/sig0000111b ;
  wire \blk0000095a/sig0000111a ;
  wire \blk0000095a/sig00001119 ;
  wire \blk0000095a/sig00001118 ;
  wire \blk0000095a/sig00001117 ;
  wire \blk0000095a/sig00001116 ;
  wire \blk0000095a/sig00001115 ;
  wire \blk00000974/sig0000112e ;
  wire \blk00000974/sig0000112d ;
  wire \blk00000974/sig0000112c ;
  wire \blk00000974/sig0000112b ;
  wire \blk00000974/sig0000112a ;
  wire \blk00000974/sig00001129 ;
  wire \blk00000974/sig00001128 ;
  wire \blk00000974/sig00001127 ;
  wire \blk00000981/sig00001152 ;
  wire \blk00000981/sig00001151 ;
  wire \blk00000981/sig00001150 ;
  wire \blk00000981/sig0000114f ;
  wire \blk00000981/sig0000114e ;
  wire \blk00000981/sig0000114d ;
  wire \blk00000981/sig0000114c ;
  wire \blk00000981/sig0000114b ;
  wire \blk00000981/sig0000114a ;
  wire \blk00000981/sig00001149 ;
  wire \blk00000981/sig00001148 ;
  wire \blk00000981/sig00001147 ;
  wire \blk00000981/sig00001146 ;
  wire \blk00000981/sig00001145 ;
  wire \blk00000981/sig00001144 ;
  wire \blk00000981/sig00001143 ;
  wire \blk00000981/sig00001142 ;
  wire \blk00000981/sig00001141 ;
  wire \blk0000099d/sig00001176 ;
  wire \blk0000099d/sig00001175 ;
  wire \blk0000099d/sig00001174 ;
  wire \blk0000099d/sig00001173 ;
  wire \blk0000099d/sig00001172 ;
  wire \blk0000099d/sig00001171 ;
  wire \blk0000099d/sig00001170 ;
  wire \blk0000099d/sig0000116f ;
  wire \blk0000099d/sig0000116e ;
  wire \blk0000099d/sig0000116d ;
  wire \blk0000099d/sig0000116c ;
  wire \blk0000099d/sig0000116b ;
  wire \blk0000099d/sig0000116a ;
  wire \blk0000099d/sig00001169 ;
  wire \blk0000099d/sig00001168 ;
  wire \blk0000099d/sig00001167 ;
  wire \blk0000099d/sig00001166 ;
  wire \blk0000099d/sig00001165 ;
  wire \blk000009cb/blk000009cc/sig00001183 ;
  wire \blk000009cb/blk000009cc/sig00001182 ;
  wire \blk000009cb/blk000009cc/sig00001181 ;
  wire \blk000009cb/blk000009cc/sig00001180 ;
  wire \blk000009cb/blk000009cc/sig0000117f ;
  wire NLW_blk000000d1_CARRYOUTF_UNCONNECTED;
  wire NLW_blk000000d1_CARRYOUT_UNCONNECTED;
  wire \NLW_blk000000d1_M<35>_UNCONNECTED ;
  wire \NLW_blk000000d1_M<34>_UNCONNECTED ;
  wire \NLW_blk000000d1_M<33>_UNCONNECTED ;
  wire \NLW_blk000000d1_M<32>_UNCONNECTED ;
  wire \NLW_blk000000d1_M<31>_UNCONNECTED ;
  wire \NLW_blk000000d1_M<30>_UNCONNECTED ;
  wire \NLW_blk000000d1_M<29>_UNCONNECTED ;
  wire \NLW_blk000000d1_M<28>_UNCONNECTED ;
  wire \NLW_blk000000d1_M<27>_UNCONNECTED ;
  wire \NLW_blk000000d1_M<26>_UNCONNECTED ;
  wire \NLW_blk000000d1_M<25>_UNCONNECTED ;
  wire \NLW_blk000000d1_M<24>_UNCONNECTED ;
  wire \NLW_blk000000d1_M<23>_UNCONNECTED ;
  wire \NLW_blk000000d1_M<22>_UNCONNECTED ;
  wire \NLW_blk000000d1_M<21>_UNCONNECTED ;
  wire \NLW_blk000000d1_M<20>_UNCONNECTED ;
  wire \NLW_blk000000d1_M<19>_UNCONNECTED ;
  wire \NLW_blk000000d1_M<18>_UNCONNECTED ;
  wire \NLW_blk000000d1_M<17>_UNCONNECTED ;
  wire \NLW_blk000000d1_M<16>_UNCONNECTED ;
  wire \NLW_blk000000d1_M<15>_UNCONNECTED ;
  wire \NLW_blk000000d1_M<14>_UNCONNECTED ;
  wire \NLW_blk000000d1_M<13>_UNCONNECTED ;
  wire \NLW_blk000000d1_M<12>_UNCONNECTED ;
  wire \NLW_blk000000d1_M<11>_UNCONNECTED ;
  wire \NLW_blk000000d1_M<10>_UNCONNECTED ;
  wire \NLW_blk000000d1_M<9>_UNCONNECTED ;
  wire \NLW_blk000000d1_M<8>_UNCONNECTED ;
  wire \NLW_blk000000d1_M<7>_UNCONNECTED ;
  wire \NLW_blk000000d1_M<6>_UNCONNECTED ;
  wire \NLW_blk000000d1_M<5>_UNCONNECTED ;
  wire \NLW_blk000000d1_M<4>_UNCONNECTED ;
  wire \NLW_blk000000d1_M<3>_UNCONNECTED ;
  wire \NLW_blk000000d1_M<2>_UNCONNECTED ;
  wire \NLW_blk000000d1_M<1>_UNCONNECTED ;
  wire \NLW_blk000000d1_M<0>_UNCONNECTED ;
  wire NLW_blk000000d2_CARRYOUTF_UNCONNECTED;
  wire NLW_blk000000d2_CARRYOUT_UNCONNECTED;
  wire \NLW_blk000000d2_BCOUT<17>_UNCONNECTED ;
  wire \NLW_blk000000d2_BCOUT<16>_UNCONNECTED ;
  wire \NLW_blk000000d2_BCOUT<15>_UNCONNECTED ;
  wire \NLW_blk000000d2_BCOUT<14>_UNCONNECTED ;
  wire \NLW_blk000000d2_BCOUT<13>_UNCONNECTED ;
  wire \NLW_blk000000d2_BCOUT<12>_UNCONNECTED ;
  wire \NLW_blk000000d2_BCOUT<11>_UNCONNECTED ;
  wire \NLW_blk000000d2_BCOUT<10>_UNCONNECTED ;
  wire \NLW_blk000000d2_BCOUT<9>_UNCONNECTED ;
  wire \NLW_blk000000d2_BCOUT<8>_UNCONNECTED ;
  wire \NLW_blk000000d2_BCOUT<7>_UNCONNECTED ;
  wire \NLW_blk000000d2_BCOUT<6>_UNCONNECTED ;
  wire \NLW_blk000000d2_BCOUT<5>_UNCONNECTED ;
  wire \NLW_blk000000d2_BCOUT<4>_UNCONNECTED ;
  wire \NLW_blk000000d2_BCOUT<3>_UNCONNECTED ;
  wire \NLW_blk000000d2_BCOUT<2>_UNCONNECTED ;
  wire \NLW_blk000000d2_BCOUT<1>_UNCONNECTED ;
  wire \NLW_blk000000d2_BCOUT<0>_UNCONNECTED ;
  wire \NLW_blk000000d2_P<47>_UNCONNECTED ;
  wire \NLW_blk000000d2_P<46>_UNCONNECTED ;
  wire \NLW_blk000000d2_P<45>_UNCONNECTED ;
  wire \NLW_blk000000d2_P<44>_UNCONNECTED ;
  wire \NLW_blk000000d2_P<43>_UNCONNECTED ;
  wire \NLW_blk000000d2_P<42>_UNCONNECTED ;
  wire \NLW_blk000000d2_P<41>_UNCONNECTED ;
  wire \NLW_blk000000d2_P<40>_UNCONNECTED ;
  wire \NLW_blk000000d2_P<39>_UNCONNECTED ;
  wire \NLW_blk000000d2_P<38>_UNCONNECTED ;
  wire \NLW_blk000000d2_P<37>_UNCONNECTED ;
  wire \NLW_blk000000d2_P<36>_UNCONNECTED ;
  wire \NLW_blk000000d2_PCOUT<47>_UNCONNECTED ;
  wire \NLW_blk000000d2_PCOUT<46>_UNCONNECTED ;
  wire \NLW_blk000000d2_PCOUT<45>_UNCONNECTED ;
  wire \NLW_blk000000d2_PCOUT<44>_UNCONNECTED ;
  wire \NLW_blk000000d2_PCOUT<43>_UNCONNECTED ;
  wire \NLW_blk000000d2_PCOUT<42>_UNCONNECTED ;
  wire \NLW_blk000000d2_PCOUT<41>_UNCONNECTED ;
  wire \NLW_blk000000d2_PCOUT<40>_UNCONNECTED ;
  wire \NLW_blk000000d2_PCOUT<39>_UNCONNECTED ;
  wire \NLW_blk000000d2_PCOUT<38>_UNCONNECTED ;
  wire \NLW_blk000000d2_PCOUT<37>_UNCONNECTED ;
  wire \NLW_blk000000d2_PCOUT<36>_UNCONNECTED ;
  wire \NLW_blk000000d2_PCOUT<35>_UNCONNECTED ;
  wire \NLW_blk000000d2_PCOUT<34>_UNCONNECTED ;
  wire \NLW_blk000000d2_PCOUT<33>_UNCONNECTED ;
  wire \NLW_blk000000d2_PCOUT<32>_UNCONNECTED ;
  wire \NLW_blk000000d2_PCOUT<31>_UNCONNECTED ;
  wire \NLW_blk000000d2_PCOUT<30>_UNCONNECTED ;
  wire \NLW_blk000000d2_PCOUT<29>_UNCONNECTED ;
  wire \NLW_blk000000d2_PCOUT<28>_UNCONNECTED ;
  wire \NLW_blk000000d2_PCOUT<27>_UNCONNECTED ;
  wire \NLW_blk000000d2_PCOUT<26>_UNCONNECTED ;
  wire \NLW_blk000000d2_PCOUT<25>_UNCONNECTED ;
  wire \NLW_blk000000d2_PCOUT<24>_UNCONNECTED ;
  wire \NLW_blk000000d2_PCOUT<23>_UNCONNECTED ;
  wire \NLW_blk000000d2_PCOUT<22>_UNCONNECTED ;
  wire \NLW_blk000000d2_PCOUT<21>_UNCONNECTED ;
  wire \NLW_blk000000d2_PCOUT<20>_UNCONNECTED ;
  wire \NLW_blk000000d2_PCOUT<19>_UNCONNECTED ;
  wire \NLW_blk000000d2_PCOUT<18>_UNCONNECTED ;
  wire \NLW_blk000000d2_PCOUT<17>_UNCONNECTED ;
  wire \NLW_blk000000d2_PCOUT<16>_UNCONNECTED ;
  wire \NLW_blk000000d2_PCOUT<15>_UNCONNECTED ;
  wire \NLW_blk000000d2_PCOUT<14>_UNCONNECTED ;
  wire \NLW_blk000000d2_PCOUT<13>_UNCONNECTED ;
  wire \NLW_blk000000d2_PCOUT<12>_UNCONNECTED ;
  wire \NLW_blk000000d2_PCOUT<11>_UNCONNECTED ;
  wire \NLW_blk000000d2_PCOUT<10>_UNCONNECTED ;
  wire \NLW_blk000000d2_PCOUT<9>_UNCONNECTED ;
  wire \NLW_blk000000d2_PCOUT<8>_UNCONNECTED ;
  wire \NLW_blk000000d2_PCOUT<7>_UNCONNECTED ;
  wire \NLW_blk000000d2_PCOUT<6>_UNCONNECTED ;
  wire \NLW_blk000000d2_PCOUT<5>_UNCONNECTED ;
  wire \NLW_blk000000d2_PCOUT<4>_UNCONNECTED ;
  wire \NLW_blk000000d2_PCOUT<3>_UNCONNECTED ;
  wire \NLW_blk000000d2_PCOUT<2>_UNCONNECTED ;
  wire \NLW_blk000000d2_PCOUT<1>_UNCONNECTED ;
  wire \NLW_blk000000d2_PCOUT<0>_UNCONNECTED ;
  wire \NLW_blk000000d2_M<35>_UNCONNECTED ;
  wire \NLW_blk000000d2_M<34>_UNCONNECTED ;
  wire \NLW_blk000000d2_M<33>_UNCONNECTED ;
  wire \NLW_blk000000d2_M<32>_UNCONNECTED ;
  wire \NLW_blk000000d2_M<31>_UNCONNECTED ;
  wire \NLW_blk000000d2_M<30>_UNCONNECTED ;
  wire \NLW_blk000000d2_M<29>_UNCONNECTED ;
  wire \NLW_blk000000d2_M<28>_UNCONNECTED ;
  wire \NLW_blk000000d2_M<27>_UNCONNECTED ;
  wire \NLW_blk000000d2_M<26>_UNCONNECTED ;
  wire \NLW_blk000000d2_M<25>_UNCONNECTED ;
  wire \NLW_blk000000d2_M<24>_UNCONNECTED ;
  wire \NLW_blk000000d2_M<23>_UNCONNECTED ;
  wire \NLW_blk000000d2_M<22>_UNCONNECTED ;
  wire \NLW_blk000000d2_M<21>_UNCONNECTED ;
  wire \NLW_blk000000d2_M<20>_UNCONNECTED ;
  wire \NLW_blk000000d2_M<19>_UNCONNECTED ;
  wire \NLW_blk000000d2_M<18>_UNCONNECTED ;
  wire \NLW_blk000000d2_M<17>_UNCONNECTED ;
  wire \NLW_blk000000d2_M<16>_UNCONNECTED ;
  wire \NLW_blk000000d2_M<15>_UNCONNECTED ;
  wire \NLW_blk000000d2_M<14>_UNCONNECTED ;
  wire \NLW_blk000000d2_M<13>_UNCONNECTED ;
  wire \NLW_blk000000d2_M<12>_UNCONNECTED ;
  wire \NLW_blk000000d2_M<11>_UNCONNECTED ;
  wire \NLW_blk000000d2_M<10>_UNCONNECTED ;
  wire \NLW_blk000000d2_M<9>_UNCONNECTED ;
  wire \NLW_blk000000d2_M<8>_UNCONNECTED ;
  wire \NLW_blk000000d2_M<7>_UNCONNECTED ;
  wire \NLW_blk000000d2_M<6>_UNCONNECTED ;
  wire \NLW_blk000000d2_M<5>_UNCONNECTED ;
  wire \NLW_blk000000d2_M<4>_UNCONNECTED ;
  wire \NLW_blk000000d2_M<3>_UNCONNECTED ;
  wire \NLW_blk000000d2_M<2>_UNCONNECTED ;
  wire \NLW_blk000000d2_M<1>_UNCONNECTED ;
  wire \NLW_blk000000d2_M<0>_UNCONNECTED ;
  wire NLW_blk000000d3_CARRYOUTF_UNCONNECTED;
  wire NLW_blk000000d3_CARRYOUT_UNCONNECTED;
  wire \NLW_blk000000d3_M<35>_UNCONNECTED ;
  wire \NLW_blk000000d3_M<34>_UNCONNECTED ;
  wire \NLW_blk000000d3_M<33>_UNCONNECTED ;
  wire \NLW_blk000000d3_M<32>_UNCONNECTED ;
  wire \NLW_blk000000d3_M<31>_UNCONNECTED ;
  wire \NLW_blk000000d3_M<30>_UNCONNECTED ;
  wire \NLW_blk000000d3_M<29>_UNCONNECTED ;
  wire \NLW_blk000000d3_M<28>_UNCONNECTED ;
  wire \NLW_blk000000d3_M<27>_UNCONNECTED ;
  wire \NLW_blk000000d3_M<26>_UNCONNECTED ;
  wire \NLW_blk000000d3_M<25>_UNCONNECTED ;
  wire \NLW_blk000000d3_M<24>_UNCONNECTED ;
  wire \NLW_blk000000d3_M<23>_UNCONNECTED ;
  wire \NLW_blk000000d3_M<22>_UNCONNECTED ;
  wire \NLW_blk000000d3_M<21>_UNCONNECTED ;
  wire \NLW_blk000000d3_M<20>_UNCONNECTED ;
  wire \NLW_blk000000d3_M<19>_UNCONNECTED ;
  wire \NLW_blk000000d3_M<18>_UNCONNECTED ;
  wire \NLW_blk000000d3_M<17>_UNCONNECTED ;
  wire \NLW_blk000000d3_M<16>_UNCONNECTED ;
  wire \NLW_blk000000d3_M<15>_UNCONNECTED ;
  wire \NLW_blk000000d3_M<14>_UNCONNECTED ;
  wire \NLW_blk000000d3_M<13>_UNCONNECTED ;
  wire \NLW_blk000000d3_M<12>_UNCONNECTED ;
  wire \NLW_blk000000d3_M<11>_UNCONNECTED ;
  wire \NLW_blk000000d3_M<10>_UNCONNECTED ;
  wire \NLW_blk000000d3_M<9>_UNCONNECTED ;
  wire \NLW_blk000000d3_M<8>_UNCONNECTED ;
  wire \NLW_blk000000d3_M<7>_UNCONNECTED ;
  wire \NLW_blk000000d3_M<6>_UNCONNECTED ;
  wire \NLW_blk000000d3_M<5>_UNCONNECTED ;
  wire \NLW_blk000000d3_M<4>_UNCONNECTED ;
  wire \NLW_blk000000d3_M<3>_UNCONNECTED ;
  wire \NLW_blk000000d3_M<2>_UNCONNECTED ;
  wire \NLW_blk000000d3_M<1>_UNCONNECTED ;
  wire \NLW_blk000000d3_M<0>_UNCONNECTED ;
  wire NLW_blk000000d4_CARRYOUTF_UNCONNECTED;
  wire NLW_blk000000d4_CARRYOUT_UNCONNECTED;
  wire \NLW_blk000000d4_BCOUT<17>_UNCONNECTED ;
  wire \NLW_blk000000d4_BCOUT<16>_UNCONNECTED ;
  wire \NLW_blk000000d4_BCOUT<15>_UNCONNECTED ;
  wire \NLW_blk000000d4_BCOUT<14>_UNCONNECTED ;
  wire \NLW_blk000000d4_BCOUT<13>_UNCONNECTED ;
  wire \NLW_blk000000d4_BCOUT<12>_UNCONNECTED ;
  wire \NLW_blk000000d4_BCOUT<11>_UNCONNECTED ;
  wire \NLW_blk000000d4_BCOUT<10>_UNCONNECTED ;
  wire \NLW_blk000000d4_BCOUT<9>_UNCONNECTED ;
  wire \NLW_blk000000d4_BCOUT<8>_UNCONNECTED ;
  wire \NLW_blk000000d4_BCOUT<7>_UNCONNECTED ;
  wire \NLW_blk000000d4_BCOUT<6>_UNCONNECTED ;
  wire \NLW_blk000000d4_BCOUT<5>_UNCONNECTED ;
  wire \NLW_blk000000d4_BCOUT<4>_UNCONNECTED ;
  wire \NLW_blk000000d4_BCOUT<3>_UNCONNECTED ;
  wire \NLW_blk000000d4_BCOUT<2>_UNCONNECTED ;
  wire \NLW_blk000000d4_BCOUT<1>_UNCONNECTED ;
  wire \NLW_blk000000d4_BCOUT<0>_UNCONNECTED ;
  wire \NLW_blk000000d4_P<47>_UNCONNECTED ;
  wire \NLW_blk000000d4_P<46>_UNCONNECTED ;
  wire \NLW_blk000000d4_P<45>_UNCONNECTED ;
  wire \NLW_blk000000d4_P<44>_UNCONNECTED ;
  wire \NLW_blk000000d4_P<43>_UNCONNECTED ;
  wire \NLW_blk000000d4_P<42>_UNCONNECTED ;
  wire \NLW_blk000000d4_P<41>_UNCONNECTED ;
  wire \NLW_blk000000d4_P<40>_UNCONNECTED ;
  wire \NLW_blk000000d4_P<39>_UNCONNECTED ;
  wire \NLW_blk000000d4_P<38>_UNCONNECTED ;
  wire \NLW_blk000000d4_P<37>_UNCONNECTED ;
  wire \NLW_blk000000d4_P<36>_UNCONNECTED ;
  wire \NLW_blk000000d4_PCOUT<47>_UNCONNECTED ;
  wire \NLW_blk000000d4_PCOUT<46>_UNCONNECTED ;
  wire \NLW_blk000000d4_PCOUT<45>_UNCONNECTED ;
  wire \NLW_blk000000d4_PCOUT<44>_UNCONNECTED ;
  wire \NLW_blk000000d4_PCOUT<43>_UNCONNECTED ;
  wire \NLW_blk000000d4_PCOUT<42>_UNCONNECTED ;
  wire \NLW_blk000000d4_PCOUT<41>_UNCONNECTED ;
  wire \NLW_blk000000d4_PCOUT<40>_UNCONNECTED ;
  wire \NLW_blk000000d4_PCOUT<39>_UNCONNECTED ;
  wire \NLW_blk000000d4_PCOUT<38>_UNCONNECTED ;
  wire \NLW_blk000000d4_PCOUT<37>_UNCONNECTED ;
  wire \NLW_blk000000d4_PCOUT<36>_UNCONNECTED ;
  wire \NLW_blk000000d4_PCOUT<35>_UNCONNECTED ;
  wire \NLW_blk000000d4_PCOUT<34>_UNCONNECTED ;
  wire \NLW_blk000000d4_PCOUT<33>_UNCONNECTED ;
  wire \NLW_blk000000d4_PCOUT<32>_UNCONNECTED ;
  wire \NLW_blk000000d4_PCOUT<31>_UNCONNECTED ;
  wire \NLW_blk000000d4_PCOUT<30>_UNCONNECTED ;
  wire \NLW_blk000000d4_PCOUT<29>_UNCONNECTED ;
  wire \NLW_blk000000d4_PCOUT<28>_UNCONNECTED ;
  wire \NLW_blk000000d4_PCOUT<27>_UNCONNECTED ;
  wire \NLW_blk000000d4_PCOUT<26>_UNCONNECTED ;
  wire \NLW_blk000000d4_PCOUT<25>_UNCONNECTED ;
  wire \NLW_blk000000d4_PCOUT<24>_UNCONNECTED ;
  wire \NLW_blk000000d4_PCOUT<23>_UNCONNECTED ;
  wire \NLW_blk000000d4_PCOUT<22>_UNCONNECTED ;
  wire \NLW_blk000000d4_PCOUT<21>_UNCONNECTED ;
  wire \NLW_blk000000d4_PCOUT<20>_UNCONNECTED ;
  wire \NLW_blk000000d4_PCOUT<19>_UNCONNECTED ;
  wire \NLW_blk000000d4_PCOUT<18>_UNCONNECTED ;
  wire \NLW_blk000000d4_PCOUT<17>_UNCONNECTED ;
  wire \NLW_blk000000d4_PCOUT<16>_UNCONNECTED ;
  wire \NLW_blk000000d4_PCOUT<15>_UNCONNECTED ;
  wire \NLW_blk000000d4_PCOUT<14>_UNCONNECTED ;
  wire \NLW_blk000000d4_PCOUT<13>_UNCONNECTED ;
  wire \NLW_blk000000d4_PCOUT<12>_UNCONNECTED ;
  wire \NLW_blk000000d4_PCOUT<11>_UNCONNECTED ;
  wire \NLW_blk000000d4_PCOUT<10>_UNCONNECTED ;
  wire \NLW_blk000000d4_PCOUT<9>_UNCONNECTED ;
  wire \NLW_blk000000d4_PCOUT<8>_UNCONNECTED ;
  wire \NLW_blk000000d4_PCOUT<7>_UNCONNECTED ;
  wire \NLW_blk000000d4_PCOUT<6>_UNCONNECTED ;
  wire \NLW_blk000000d4_PCOUT<5>_UNCONNECTED ;
  wire \NLW_blk000000d4_PCOUT<4>_UNCONNECTED ;
  wire \NLW_blk000000d4_PCOUT<3>_UNCONNECTED ;
  wire \NLW_blk000000d4_PCOUT<2>_UNCONNECTED ;
  wire \NLW_blk000000d4_PCOUT<1>_UNCONNECTED ;
  wire \NLW_blk000000d4_PCOUT<0>_UNCONNECTED ;
  wire \NLW_blk000000d4_M<35>_UNCONNECTED ;
  wire \NLW_blk000000d4_M<34>_UNCONNECTED ;
  wire \NLW_blk000000d4_M<33>_UNCONNECTED ;
  wire \NLW_blk000000d4_M<32>_UNCONNECTED ;
  wire \NLW_blk000000d4_M<31>_UNCONNECTED ;
  wire \NLW_blk000000d4_M<30>_UNCONNECTED ;
  wire \NLW_blk000000d4_M<29>_UNCONNECTED ;
  wire \NLW_blk000000d4_M<28>_UNCONNECTED ;
  wire \NLW_blk000000d4_M<27>_UNCONNECTED ;
  wire \NLW_blk000000d4_M<26>_UNCONNECTED ;
  wire \NLW_blk000000d4_M<25>_UNCONNECTED ;
  wire \NLW_blk000000d4_M<24>_UNCONNECTED ;
  wire \NLW_blk000000d4_M<23>_UNCONNECTED ;
  wire \NLW_blk000000d4_M<22>_UNCONNECTED ;
  wire \NLW_blk000000d4_M<21>_UNCONNECTED ;
  wire \NLW_blk000000d4_M<20>_UNCONNECTED ;
  wire \NLW_blk000000d4_M<19>_UNCONNECTED ;
  wire \NLW_blk000000d4_M<18>_UNCONNECTED ;
  wire \NLW_blk000000d4_M<17>_UNCONNECTED ;
  wire \NLW_blk000000d4_M<16>_UNCONNECTED ;
  wire \NLW_blk000000d4_M<15>_UNCONNECTED ;
  wire \NLW_blk000000d4_M<14>_UNCONNECTED ;
  wire \NLW_blk000000d4_M<13>_UNCONNECTED ;
  wire \NLW_blk000000d4_M<12>_UNCONNECTED ;
  wire \NLW_blk000000d4_M<11>_UNCONNECTED ;
  wire \NLW_blk000000d4_M<10>_UNCONNECTED ;
  wire \NLW_blk000000d4_M<9>_UNCONNECTED ;
  wire \NLW_blk000000d4_M<8>_UNCONNECTED ;
  wire \NLW_blk000000d4_M<7>_UNCONNECTED ;
  wire \NLW_blk000000d4_M<6>_UNCONNECTED ;
  wire \NLW_blk000000d4_M<5>_UNCONNECTED ;
  wire \NLW_blk000000d4_M<4>_UNCONNECTED ;
  wire \NLW_blk000000d4_M<3>_UNCONNECTED ;
  wire \NLW_blk000000d4_M<2>_UNCONNECTED ;
  wire \NLW_blk000000d4_M<1>_UNCONNECTED ;
  wire \NLW_blk000000d4_M<0>_UNCONNECTED ;
  wire NLW_blk00000184_CARRYOUTF_UNCONNECTED;
  wire NLW_blk00000184_CARRYOUT_UNCONNECTED;
  wire \NLW_blk00000184_BCOUT<17>_UNCONNECTED ;
  wire \NLW_blk00000184_BCOUT<16>_UNCONNECTED ;
  wire \NLW_blk00000184_BCOUT<15>_UNCONNECTED ;
  wire \NLW_blk00000184_BCOUT<14>_UNCONNECTED ;
  wire \NLW_blk00000184_BCOUT<13>_UNCONNECTED ;
  wire \NLW_blk00000184_BCOUT<12>_UNCONNECTED ;
  wire \NLW_blk00000184_BCOUT<11>_UNCONNECTED ;
  wire \NLW_blk00000184_BCOUT<10>_UNCONNECTED ;
  wire \NLW_blk00000184_BCOUT<9>_UNCONNECTED ;
  wire \NLW_blk00000184_BCOUT<8>_UNCONNECTED ;
  wire \NLW_blk00000184_BCOUT<7>_UNCONNECTED ;
  wire \NLW_blk00000184_BCOUT<6>_UNCONNECTED ;
  wire \NLW_blk00000184_BCOUT<5>_UNCONNECTED ;
  wire \NLW_blk00000184_BCOUT<4>_UNCONNECTED ;
  wire \NLW_blk00000184_BCOUT<3>_UNCONNECTED ;
  wire \NLW_blk00000184_BCOUT<2>_UNCONNECTED ;
  wire \NLW_blk00000184_BCOUT<1>_UNCONNECTED ;
  wire \NLW_blk00000184_BCOUT<0>_UNCONNECTED ;
  wire \NLW_blk00000184_P<47>_UNCONNECTED ;
  wire \NLW_blk00000184_P<46>_UNCONNECTED ;
  wire \NLW_blk00000184_P<45>_UNCONNECTED ;
  wire \NLW_blk00000184_P<44>_UNCONNECTED ;
  wire \NLW_blk00000184_P<43>_UNCONNECTED ;
  wire \NLW_blk00000184_P<42>_UNCONNECTED ;
  wire \NLW_blk00000184_P<41>_UNCONNECTED ;
  wire \NLW_blk00000184_P<40>_UNCONNECTED ;
  wire \NLW_blk00000184_P<39>_UNCONNECTED ;
  wire \NLW_blk00000184_P<38>_UNCONNECTED ;
  wire \NLW_blk00000184_P<37>_UNCONNECTED ;
  wire \NLW_blk00000184_P<36>_UNCONNECTED ;
  wire \NLW_blk00000184_PCOUT<47>_UNCONNECTED ;
  wire \NLW_blk00000184_PCOUT<46>_UNCONNECTED ;
  wire \NLW_blk00000184_PCOUT<45>_UNCONNECTED ;
  wire \NLW_blk00000184_PCOUT<44>_UNCONNECTED ;
  wire \NLW_blk00000184_PCOUT<43>_UNCONNECTED ;
  wire \NLW_blk00000184_PCOUT<42>_UNCONNECTED ;
  wire \NLW_blk00000184_PCOUT<41>_UNCONNECTED ;
  wire \NLW_blk00000184_PCOUT<40>_UNCONNECTED ;
  wire \NLW_blk00000184_PCOUT<39>_UNCONNECTED ;
  wire \NLW_blk00000184_PCOUT<38>_UNCONNECTED ;
  wire \NLW_blk00000184_PCOUT<37>_UNCONNECTED ;
  wire \NLW_blk00000184_PCOUT<36>_UNCONNECTED ;
  wire \NLW_blk00000184_PCOUT<35>_UNCONNECTED ;
  wire \NLW_blk00000184_PCOUT<34>_UNCONNECTED ;
  wire \NLW_blk00000184_PCOUT<33>_UNCONNECTED ;
  wire \NLW_blk00000184_PCOUT<32>_UNCONNECTED ;
  wire \NLW_blk00000184_PCOUT<31>_UNCONNECTED ;
  wire \NLW_blk00000184_PCOUT<30>_UNCONNECTED ;
  wire \NLW_blk00000184_PCOUT<29>_UNCONNECTED ;
  wire \NLW_blk00000184_PCOUT<28>_UNCONNECTED ;
  wire \NLW_blk00000184_PCOUT<27>_UNCONNECTED ;
  wire \NLW_blk00000184_PCOUT<26>_UNCONNECTED ;
  wire \NLW_blk00000184_PCOUT<25>_UNCONNECTED ;
  wire \NLW_blk00000184_PCOUT<24>_UNCONNECTED ;
  wire \NLW_blk00000184_PCOUT<23>_UNCONNECTED ;
  wire \NLW_blk00000184_PCOUT<22>_UNCONNECTED ;
  wire \NLW_blk00000184_PCOUT<21>_UNCONNECTED ;
  wire \NLW_blk00000184_PCOUT<20>_UNCONNECTED ;
  wire \NLW_blk00000184_PCOUT<19>_UNCONNECTED ;
  wire \NLW_blk00000184_PCOUT<18>_UNCONNECTED ;
  wire \NLW_blk00000184_PCOUT<17>_UNCONNECTED ;
  wire \NLW_blk00000184_PCOUT<16>_UNCONNECTED ;
  wire \NLW_blk00000184_PCOUT<15>_UNCONNECTED ;
  wire \NLW_blk00000184_PCOUT<14>_UNCONNECTED ;
  wire \NLW_blk00000184_PCOUT<13>_UNCONNECTED ;
  wire \NLW_blk00000184_PCOUT<12>_UNCONNECTED ;
  wire \NLW_blk00000184_PCOUT<11>_UNCONNECTED ;
  wire \NLW_blk00000184_PCOUT<10>_UNCONNECTED ;
  wire \NLW_blk00000184_PCOUT<9>_UNCONNECTED ;
  wire \NLW_blk00000184_PCOUT<8>_UNCONNECTED ;
  wire \NLW_blk00000184_PCOUT<7>_UNCONNECTED ;
  wire \NLW_blk00000184_PCOUT<6>_UNCONNECTED ;
  wire \NLW_blk00000184_PCOUT<5>_UNCONNECTED ;
  wire \NLW_blk00000184_PCOUT<4>_UNCONNECTED ;
  wire \NLW_blk00000184_PCOUT<3>_UNCONNECTED ;
  wire \NLW_blk00000184_PCOUT<2>_UNCONNECTED ;
  wire \NLW_blk00000184_PCOUT<1>_UNCONNECTED ;
  wire \NLW_blk00000184_PCOUT<0>_UNCONNECTED ;
  wire \NLW_blk00000184_M<35>_UNCONNECTED ;
  wire \NLW_blk00000184_M<34>_UNCONNECTED ;
  wire \NLW_blk00000184_M<33>_UNCONNECTED ;
  wire \NLW_blk00000184_M<32>_UNCONNECTED ;
  wire \NLW_blk00000184_M<31>_UNCONNECTED ;
  wire \NLW_blk00000184_M<30>_UNCONNECTED ;
  wire \NLW_blk00000184_M<29>_UNCONNECTED ;
  wire \NLW_blk00000184_M<28>_UNCONNECTED ;
  wire \NLW_blk00000184_M<27>_UNCONNECTED ;
  wire \NLW_blk00000184_M<26>_UNCONNECTED ;
  wire \NLW_blk00000184_M<25>_UNCONNECTED ;
  wire \NLW_blk00000184_M<24>_UNCONNECTED ;
  wire \NLW_blk00000184_M<23>_UNCONNECTED ;
  wire \NLW_blk00000184_M<22>_UNCONNECTED ;
  wire \NLW_blk00000184_M<21>_UNCONNECTED ;
  wire \NLW_blk00000184_M<20>_UNCONNECTED ;
  wire \NLW_blk00000184_M<19>_UNCONNECTED ;
  wire \NLW_blk00000184_M<18>_UNCONNECTED ;
  wire \NLW_blk00000184_M<17>_UNCONNECTED ;
  wire \NLW_blk00000184_M<16>_UNCONNECTED ;
  wire \NLW_blk00000184_M<15>_UNCONNECTED ;
  wire \NLW_blk00000184_M<14>_UNCONNECTED ;
  wire \NLW_blk00000184_M<13>_UNCONNECTED ;
  wire \NLW_blk00000184_M<12>_UNCONNECTED ;
  wire \NLW_blk00000184_M<11>_UNCONNECTED ;
  wire \NLW_blk00000184_M<10>_UNCONNECTED ;
  wire \NLW_blk00000184_M<9>_UNCONNECTED ;
  wire \NLW_blk00000184_M<8>_UNCONNECTED ;
  wire \NLW_blk00000184_M<7>_UNCONNECTED ;
  wire \NLW_blk00000184_M<6>_UNCONNECTED ;
  wire \NLW_blk00000184_M<5>_UNCONNECTED ;
  wire \NLW_blk00000184_M<4>_UNCONNECTED ;
  wire \NLW_blk00000184_M<3>_UNCONNECTED ;
  wire \NLW_blk00000184_M<2>_UNCONNECTED ;
  wire \NLW_blk00000184_M<1>_UNCONNECTED ;
  wire \NLW_blk00000184_M<0>_UNCONNECTED ;
  wire NLW_blk00000185_CARRYOUTF_UNCONNECTED;
  wire NLW_blk00000185_CARRYOUT_UNCONNECTED;
  wire \NLW_blk00000185_M<35>_UNCONNECTED ;
  wire \NLW_blk00000185_M<34>_UNCONNECTED ;
  wire \NLW_blk00000185_M<33>_UNCONNECTED ;
  wire \NLW_blk00000185_M<32>_UNCONNECTED ;
  wire \NLW_blk00000185_M<31>_UNCONNECTED ;
  wire \NLW_blk00000185_M<30>_UNCONNECTED ;
  wire \NLW_blk00000185_M<29>_UNCONNECTED ;
  wire \NLW_blk00000185_M<28>_UNCONNECTED ;
  wire \NLW_blk00000185_M<27>_UNCONNECTED ;
  wire \NLW_blk00000185_M<26>_UNCONNECTED ;
  wire \NLW_blk00000185_M<25>_UNCONNECTED ;
  wire \NLW_blk00000185_M<24>_UNCONNECTED ;
  wire \NLW_blk00000185_M<23>_UNCONNECTED ;
  wire \NLW_blk00000185_M<22>_UNCONNECTED ;
  wire \NLW_blk00000185_M<21>_UNCONNECTED ;
  wire \NLW_blk00000185_M<20>_UNCONNECTED ;
  wire \NLW_blk00000185_M<19>_UNCONNECTED ;
  wire \NLW_blk00000185_M<18>_UNCONNECTED ;
  wire \NLW_blk00000185_M<17>_UNCONNECTED ;
  wire \NLW_blk00000185_M<16>_UNCONNECTED ;
  wire \NLW_blk00000185_M<15>_UNCONNECTED ;
  wire \NLW_blk00000185_M<14>_UNCONNECTED ;
  wire \NLW_blk00000185_M<13>_UNCONNECTED ;
  wire \NLW_blk00000185_M<12>_UNCONNECTED ;
  wire \NLW_blk00000185_M<11>_UNCONNECTED ;
  wire \NLW_blk00000185_M<10>_UNCONNECTED ;
  wire \NLW_blk00000185_M<9>_UNCONNECTED ;
  wire \NLW_blk00000185_M<8>_UNCONNECTED ;
  wire \NLW_blk00000185_M<7>_UNCONNECTED ;
  wire \NLW_blk00000185_M<6>_UNCONNECTED ;
  wire \NLW_blk00000185_M<5>_UNCONNECTED ;
  wire \NLW_blk00000185_M<4>_UNCONNECTED ;
  wire \NLW_blk00000185_M<3>_UNCONNECTED ;
  wire \NLW_blk00000185_M<2>_UNCONNECTED ;
  wire \NLW_blk00000185_M<1>_UNCONNECTED ;
  wire \NLW_blk00000185_M<0>_UNCONNECTED ;
  wire NLW_blk00000425_Q_UNCONNECTED;
  wire NLW_blk0000044d_Q_UNCONNECTED;
  wire NLW_blk00000475_Q_UNCONNECTED;
  wire NLW_blk0000049d_Q_UNCONNECTED;
  wire NLW_blk000008c7_Q_UNCONNECTED;
  wire \NLW_blk00000a47_DOADO<15>_UNCONNECTED ;
  wire \NLW_blk00000a47_DOADO<14>_UNCONNECTED ;
  wire \NLW_blk00000a47_DOADO<13>_UNCONNECTED ;
  wire \NLW_blk00000a47_DOADO<12>_UNCONNECTED ;
  wire \NLW_blk00000a47_DOADO<11>_UNCONNECTED ;
  wire \NLW_blk00000a47_DOADO<10>_UNCONNECTED ;
  wire \NLW_blk00000a47_DOPADOP<1>_UNCONNECTED ;
  wire \NLW_blk00000a47_DOPADOP<0>_UNCONNECTED ;
  wire \NLW_blk00000a47_DOPBDOP<1>_UNCONNECTED ;
  wire \NLW_blk00000a47_DOPBDOP<0>_UNCONNECTED ;
  wire \NLW_blk00000a47_ADDRAWRADDR<3>_UNCONNECTED ;
  wire \NLW_blk00000a47_ADDRAWRADDR<2>_UNCONNECTED ;
  wire \NLW_blk00000a47_ADDRAWRADDR<1>_UNCONNECTED ;
  wire \NLW_blk00000a47_ADDRAWRADDR<0>_UNCONNECTED ;
  wire \NLW_blk00000a47_DIPBDIP<1>_UNCONNECTED ;
  wire \NLW_blk00000a47_DIPBDIP<0>_UNCONNECTED ;
  wire \NLW_blk00000a47_DIBDI<15>_UNCONNECTED ;
  wire \NLW_blk00000a47_DIBDI<14>_UNCONNECTED ;
  wire \NLW_blk00000a47_DIBDI<13>_UNCONNECTED ;
  wire \NLW_blk00000a47_DIBDI<12>_UNCONNECTED ;
  wire \NLW_blk00000a47_DIBDI<11>_UNCONNECTED ;
  wire \NLW_blk00000a47_DIBDI<10>_UNCONNECTED ;
  wire \NLW_blk00000a47_DIBDI<9>_UNCONNECTED ;
  wire \NLW_blk00000a47_DIBDI<8>_UNCONNECTED ;
  wire \NLW_blk00000a47_DIBDI<7>_UNCONNECTED ;
  wire \NLW_blk00000a47_DIBDI<6>_UNCONNECTED ;
  wire \NLW_blk00000a47_DIBDI<5>_UNCONNECTED ;
  wire \NLW_blk00000a47_DIBDI<4>_UNCONNECTED ;
  wire \NLW_blk00000a47_DIBDI<3>_UNCONNECTED ;
  wire \NLW_blk00000a47_DIBDI<2>_UNCONNECTED ;
  wire \NLW_blk00000a47_DIBDI<1>_UNCONNECTED ;
  wire \NLW_blk00000a47_DIBDI<0>_UNCONNECTED ;
  wire \NLW_blk00000a47_ADDRBRDADDR<3>_UNCONNECTED ;
  wire \NLW_blk00000a47_ADDRBRDADDR<2>_UNCONNECTED ;
  wire \NLW_blk00000a47_ADDRBRDADDR<1>_UNCONNECTED ;
  wire \NLW_blk00000a47_ADDRBRDADDR<0>_UNCONNECTED ;
  wire \NLW_blk00000a47_DOBDO<15>_UNCONNECTED ;
  wire \NLW_blk00000a47_DOBDO<14>_UNCONNECTED ;
  wire \NLW_blk00000a47_DOBDO<13>_UNCONNECTED ;
  wire \NLW_blk00000a47_DOBDO<12>_UNCONNECTED ;
  wire \NLW_blk00000a47_DOBDO<11>_UNCONNECTED ;
  wire \NLW_blk00000a47_DOBDO<10>_UNCONNECTED ;
  wire NLW_blk00000a48_Q15_UNCONNECTED;
  wire NLW_blk00000a4a_Q15_UNCONNECTED;
  wire NLW_blk00000a4c_Q15_UNCONNECTED;
  wire NLW_blk00000a4e_Q15_UNCONNECTED;
  wire NLW_blk00000a50_Q15_UNCONNECTED;
  wire NLW_blk00000a52_Q15_UNCONNECTED;
  wire NLW_blk00000a54_Q15_UNCONNECTED;
  wire NLW_blk00000a56_Q15_UNCONNECTED;
  wire NLW_blk00000a58_Q15_UNCONNECTED;
  wire NLW_blk00000a5a_Q15_UNCONNECTED;
  wire NLW_blk00000a5c_Q15_UNCONNECTED;
  wire NLW_blk00000a5e_Q15_UNCONNECTED;
  wire NLW_blk00000a60_Q15_UNCONNECTED;
  wire NLW_blk00000a62_Q15_UNCONNECTED;
  wire NLW_blk00000a64_Q15_UNCONNECTED;
  wire NLW_blk00000a66_Q15_UNCONNECTED;
  wire NLW_blk00000a68_Q15_UNCONNECTED;
  wire NLW_blk00000a6a_Q15_UNCONNECTED;
  wire NLW_blk00000a6c_Q15_UNCONNECTED;
  wire NLW_blk00000a6e_Q15_UNCONNECTED;
  wire NLW_blk00000a70_Q15_UNCONNECTED;
  wire NLW_blk00000a72_Q15_UNCONNECTED;
  wire NLW_blk00000a74_Q15_UNCONNECTED;
  wire NLW_blk00000a76_Q15_UNCONNECTED;
  wire NLW_blk00000a78_Q15_UNCONNECTED;
  wire NLW_blk00000a7a_Q15_UNCONNECTED;
  wire NLW_blk00000a7c_Q15_UNCONNECTED;
  wire NLW_blk00000a7e_Q15_UNCONNECTED;
  wire NLW_blk00000a80_Q15_UNCONNECTED;
  wire NLW_blk00000a82_Q15_UNCONNECTED;
  wire NLW_blk00000a84_Q15_UNCONNECTED;
  wire NLW_blk00000a86_Q15_UNCONNECTED;
  wire NLW_blk00000a88_Q15_UNCONNECTED;
  wire NLW_blk00000a8a_Q15_UNCONNECTED;
  wire NLW_blk00000a8c_Q15_UNCONNECTED;
  wire NLW_blk00000a8e_Q15_UNCONNECTED;
  wire NLW_blk00000a90_Q15_UNCONNECTED;
  wire NLW_blk00000a92_Q15_UNCONNECTED;
  wire NLW_blk00000a94_Q15_UNCONNECTED;
  wire NLW_blk00000a96_Q15_UNCONNECTED;
  wire NLW_blk00000a98_Q15_UNCONNECTED;
  wire NLW_blk00000a9a_Q15_UNCONNECTED;
  wire NLW_blk00000a9c_Q15_UNCONNECTED;
  wire NLW_blk00000a9e_Q15_UNCONNECTED;
  wire NLW_blk00000aa0_Q15_UNCONNECTED;
  wire NLW_blk00000aa2_Q15_UNCONNECTED;
  wire NLW_blk00000aa4_Q15_UNCONNECTED;
  wire NLW_blk00000aa6_Q15_UNCONNECTED;
  wire NLW_blk00000aa8_Q15_UNCONNECTED;
  wire NLW_blk00000aaa_Q15_UNCONNECTED;
  wire NLW_blk00000aac_Q15_UNCONNECTED;
  wire NLW_blk00000aae_Q15_UNCONNECTED;
  wire NLW_blk00000ab0_Q15_UNCONNECTED;
  wire NLW_blk00000ab2_Q15_UNCONNECTED;
  wire NLW_blk00000ab4_Q15_UNCONNECTED;
  wire NLW_blk00000ab6_Q15_UNCONNECTED;
  wire NLW_blk00000ab8_Q15_UNCONNECTED;
  wire NLW_blk00000aba_Q15_UNCONNECTED;
  wire NLW_blk00000abc_Q15_UNCONNECTED;
  wire NLW_blk00000abe_Q15_UNCONNECTED;
  wire \NLW_blk00000003/blk0000002c_DOADO<15>_UNCONNECTED ;
  wire \NLW_blk00000003/blk0000002c_DOADO<14>_UNCONNECTED ;
  wire \NLW_blk00000003/blk0000002c_DOADO<13>_UNCONNECTED ;
  wire \NLW_blk00000003/blk0000002c_DOADO<12>_UNCONNECTED ;
  wire \NLW_blk00000003/blk0000002c_DOADO<11>_UNCONNECTED ;
  wire \NLW_blk00000003/blk0000002c_DOADO<10>_UNCONNECTED ;
  wire \NLW_blk00000003/blk0000002c_DOADO<9>_UNCONNECTED ;
  wire \NLW_blk00000003/blk0000002c_DOADO<8>_UNCONNECTED ;
  wire \NLW_blk00000003/blk0000002c_DOADO<7>_UNCONNECTED ;
  wire \NLW_blk00000003/blk0000002c_DOADO<6>_UNCONNECTED ;
  wire \NLW_blk00000003/blk0000002c_DOADO<5>_UNCONNECTED ;
  wire \NLW_blk00000003/blk0000002c_DOADO<4>_UNCONNECTED ;
  wire \NLW_blk00000003/blk0000002c_DOADO<3>_UNCONNECTED ;
  wire \NLW_blk00000003/blk0000002c_DOADO<2>_UNCONNECTED ;
  wire \NLW_blk00000003/blk0000002c_DOPADOP<1>_UNCONNECTED ;
  wire \NLW_blk00000003/blk0000002c_DOPADOP<0>_UNCONNECTED ;
  wire \NLW_blk00000003/blk0000002c_DOPBDOP<1>_UNCONNECTED ;
  wire \NLW_blk00000003/blk0000002c_DOPBDOP<0>_UNCONNECTED ;
  wire \NLW_blk00000003/blk0000002c_DOBDO<15>_UNCONNECTED ;
  wire \NLW_blk00000003/blk0000002c_DOBDO<14>_UNCONNECTED ;
  wire \NLW_blk00000003/blk0000002c_DOBDO<13>_UNCONNECTED ;
  wire \NLW_blk00000003/blk0000002c_DOBDO<12>_UNCONNECTED ;
  wire \NLW_blk00000003/blk0000002c_DOBDO<11>_UNCONNECTED ;
  wire \NLW_blk00000003/blk0000002c_DOBDO<10>_UNCONNECTED ;
  wire \NLW_blk00000003/blk0000002c_DOBDO<9>_UNCONNECTED ;
  wire \NLW_blk00000003/blk0000002c_DOBDO<8>_UNCONNECTED ;
  wire \NLW_blk00000003/blk0000002c_DOBDO<7>_UNCONNECTED ;
  wire \NLW_blk00000003/blk0000002c_DOBDO<6>_UNCONNECTED ;
  wire \NLW_blk00000003/blk0000002c_DOBDO<5>_UNCONNECTED ;
  wire \NLW_blk00000003/blk0000002c_DOBDO<4>_UNCONNECTED ;
  wire \NLW_blk00000003/blk0000002c_DOBDO<3>_UNCONNECTED ;
  wire \NLW_blk00000003/blk0000002c_DOBDO<2>_UNCONNECTED ;
  wire \NLW_blk00000003/blk0000002c_DOBDO<1>_UNCONNECTED ;
  wire \NLW_blk00000003/blk0000002c_DOBDO<0>_UNCONNECTED ;
  wire \NLW_blk0000002d/blk00000056_DOADO<15>_UNCONNECTED ;
  wire \NLW_blk0000002d/blk00000056_DOADO<14>_UNCONNECTED ;
  wire \NLW_blk0000002d/blk00000056_DOADO<13>_UNCONNECTED ;
  wire \NLW_blk0000002d/blk00000056_DOADO<12>_UNCONNECTED ;
  wire \NLW_blk0000002d/blk00000056_DOADO<11>_UNCONNECTED ;
  wire \NLW_blk0000002d/blk00000056_DOADO<10>_UNCONNECTED ;
  wire \NLW_blk0000002d/blk00000056_DOADO<9>_UNCONNECTED ;
  wire \NLW_blk0000002d/blk00000056_DOADO<8>_UNCONNECTED ;
  wire \NLW_blk0000002d/blk00000056_DOADO<7>_UNCONNECTED ;
  wire \NLW_blk0000002d/blk00000056_DOADO<6>_UNCONNECTED ;
  wire \NLW_blk0000002d/blk00000056_DOADO<5>_UNCONNECTED ;
  wire \NLW_blk0000002d/blk00000056_DOADO<4>_UNCONNECTED ;
  wire \NLW_blk0000002d/blk00000056_DOADO<3>_UNCONNECTED ;
  wire \NLW_blk0000002d/blk00000056_DOADO<2>_UNCONNECTED ;
  wire \NLW_blk0000002d/blk00000056_DOPADOP<1>_UNCONNECTED ;
  wire \NLW_blk0000002d/blk00000056_DOPADOP<0>_UNCONNECTED ;
  wire \NLW_blk0000002d/blk00000056_DOPBDOP<1>_UNCONNECTED ;
  wire \NLW_blk0000002d/blk00000056_DOPBDOP<0>_UNCONNECTED ;
  wire \NLW_blk0000002d/blk00000056_DOBDO<15>_UNCONNECTED ;
  wire \NLW_blk0000002d/blk00000056_DOBDO<14>_UNCONNECTED ;
  wire \NLW_blk0000002d/blk00000056_DOBDO<13>_UNCONNECTED ;
  wire \NLW_blk0000002d/blk00000056_DOBDO<12>_UNCONNECTED ;
  wire \NLW_blk0000002d/blk00000056_DOBDO<11>_UNCONNECTED ;
  wire \NLW_blk0000002d/blk00000056_DOBDO<10>_UNCONNECTED ;
  wire \NLW_blk0000002d/blk00000056_DOBDO<9>_UNCONNECTED ;
  wire \NLW_blk0000002d/blk00000056_DOBDO<8>_UNCONNECTED ;
  wire \NLW_blk0000002d/blk00000056_DOBDO<7>_UNCONNECTED ;
  wire \NLW_blk0000002d/blk00000056_DOBDO<6>_UNCONNECTED ;
  wire \NLW_blk0000002d/blk00000056_DOBDO<5>_UNCONNECTED ;
  wire \NLW_blk0000002d/blk00000056_DOBDO<4>_UNCONNECTED ;
  wire \NLW_blk0000002d/blk00000056_DOBDO<3>_UNCONNECTED ;
  wire \NLW_blk0000002d/blk00000056_DOBDO<2>_UNCONNECTED ;
  wire \NLW_blk0000002d/blk00000056_DOBDO<1>_UNCONNECTED ;
  wire \NLW_blk0000002d/blk00000056_DOBDO<0>_UNCONNECTED ;
  wire \NLW_blk0000018c/blk00000192_Q15_UNCONNECTED ;
  wire \NLW_blk0000018c/blk00000190_Q15_UNCONNECTED ;
  wire \NLW_blk0000018c/blk0000018e_Q15_UNCONNECTED ;
  wire \NLW_blk00000194/blk0000019a_Q15_UNCONNECTED ;
  wire \NLW_blk00000194/blk00000198_Q15_UNCONNECTED ;
  wire \NLW_blk00000194/blk00000196_Q15_UNCONNECTED ;
  wire \NLW_blk0000019d/blk000001b5_Q15_UNCONNECTED ;
  wire \NLW_blk0000019d/blk000001b3_Q15_UNCONNECTED ;
  wire \NLW_blk0000019d/blk000001b1_Q15_UNCONNECTED ;
  wire \NLW_blk0000019d/blk000001af_Q15_UNCONNECTED ;
  wire \NLW_blk0000019d/blk000001ad_Q15_UNCONNECTED ;
  wire \NLW_blk0000019d/blk000001ab_Q15_UNCONNECTED ;
  wire \NLW_blk0000019d/blk000001a9_Q15_UNCONNECTED ;
  wire \NLW_blk0000019d/blk000001a7_Q15_UNCONNECTED ;
  wire \NLW_blk0000019d/blk000001a5_Q15_UNCONNECTED ;
  wire \NLW_blk0000019d/blk000001a3_Q15_UNCONNECTED ;
  wire \NLW_blk0000019d/blk000001a1_Q15_UNCONNECTED ;
  wire \NLW_blk0000019d/blk0000019f_Q15_UNCONNECTED ;
  wire \NLW_blk000001b7/blk000001cf_Q15_UNCONNECTED ;
  wire \NLW_blk000001b7/blk000001cd_Q15_UNCONNECTED ;
  wire \NLW_blk000001b7/blk000001cb_Q15_UNCONNECTED ;
  wire \NLW_blk000001b7/blk000001c9_Q15_UNCONNECTED ;
  wire \NLW_blk000001b7/blk000001c7_Q15_UNCONNECTED ;
  wire \NLW_blk000001b7/blk000001c5_Q15_UNCONNECTED ;
  wire \NLW_blk000001b7/blk000001c3_Q15_UNCONNECTED ;
  wire \NLW_blk000001b7/blk000001c1_Q15_UNCONNECTED ;
  wire \NLW_blk000001b7/blk000001bf_Q15_UNCONNECTED ;
  wire \NLW_blk000001b7/blk000001bd_Q15_UNCONNECTED ;
  wire \NLW_blk000001b7/blk000001bb_Q15_UNCONNECTED ;
  wire \NLW_blk000001b7/blk000001b9_Q15_UNCONNECTED ;
  wire \NLW_blk000001d1/blk000001f3_Q15_UNCONNECTED ;
  wire \NLW_blk000001d1/blk000001f1_Q15_UNCONNECTED ;
  wire \NLW_blk000001d1/blk000001ef_Q15_UNCONNECTED ;
  wire \NLW_blk000001d1/blk000001ed_Q15_UNCONNECTED ;
  wire \NLW_blk000001d1/blk000001eb_Q15_UNCONNECTED ;
  wire \NLW_blk000001d1/blk000001e9_Q15_UNCONNECTED ;
  wire \NLW_blk000001d1/blk000001e7_Q15_UNCONNECTED ;
  wire \NLW_blk000001d1/blk000001e5_Q15_UNCONNECTED ;
  wire \NLW_blk000001d1/blk000001e3_Q15_UNCONNECTED ;
  wire \NLW_blk000001d1/blk000001e1_Q15_UNCONNECTED ;
  wire \NLW_blk000001d1/blk000001df_Q15_UNCONNECTED ;
  wire \NLW_blk000001d1/blk000001dd_Q15_UNCONNECTED ;
  wire \NLW_blk000001d1/blk000001db_Q15_UNCONNECTED ;
  wire \NLW_blk000001d1/blk000001d9_Q15_UNCONNECTED ;
  wire \NLW_blk000001d1/blk000001d7_Q15_UNCONNECTED ;
  wire \NLW_blk000001d1/blk000001d5_Q15_UNCONNECTED ;
  wire \NLW_blk000001d1/blk000001d3_Q15_UNCONNECTED ;
  wire \NLW_blk000001f8/blk000001fc_Q15_UNCONNECTED ;
  wire \NLW_blk000001f8/blk000001fa_Q15_UNCONNECTED ;
  wire \NLW_blk000001fe/blk00000202_O_UNCONNECTED ;
  wire \NLW_blk000001fe/blk00000201_O_UNCONNECTED ;
  wire \NLW_blk0000025d/blk00000261_O_UNCONNECTED ;
  wire \NLW_blk0000025d/blk00000260_O_UNCONNECTED ;
  wire \NLW_blk000002bc/blk000002d6_O_UNCONNECTED ;
  wire \NLW_blk000002bc/blk000002d5_O_UNCONNECTED ;
  wire \NLW_blk0000031b/blk00000335_O_UNCONNECTED ;
  wire \NLW_blk0000031b/blk00000334_O_UNCONNECTED ;
  wire \NLW_blk00000751/blk00000752/blk00000755_Q15_UNCONNECTED ;
  wire \NLW_blk00000757/blk00000758/blk0000075b_Q15_UNCONNECTED ;
  wire \NLW_blk000007ea/blk000007eb/blk000007fc_Q31_UNCONNECTED ;
  wire \NLW_blk000007ea/blk000007eb/blk000007fa_Q31_UNCONNECTED ;
  wire \NLW_blk000007ea/blk000007eb/blk000007f8_Q31_UNCONNECTED ;
  wire \NLW_blk000007ea/blk000007eb/blk000007f6_Q31_UNCONNECTED ;
  wire \NLW_blk000007ea/blk000007eb/blk000007f4_Q31_UNCONNECTED ;
  wire \NLW_blk000007ea/blk000007eb/blk000007f2_Q31_UNCONNECTED ;
  wire \NLW_blk000007ea/blk000007eb/blk000007f0_Q31_UNCONNECTED ;
  wire \NLW_blk000007ea/blk000007eb/blk000007ee_Q31_UNCONNECTED ;
  wire \NLW_blk000007fe/blk000007ff/blk00000810_Q31_UNCONNECTED ;
  wire \NLW_blk000007fe/blk000007ff/blk0000080e_Q31_UNCONNECTED ;
  wire \NLW_blk000007fe/blk000007ff/blk0000080c_Q31_UNCONNECTED ;
  wire \NLW_blk000007fe/blk000007ff/blk0000080a_Q31_UNCONNECTED ;
  wire \NLW_blk000007fe/blk000007ff/blk00000808_Q31_UNCONNECTED ;
  wire \NLW_blk000007fe/blk000007ff/blk00000806_Q31_UNCONNECTED ;
  wire \NLW_blk000007fe/blk000007ff/blk00000804_Q31_UNCONNECTED ;
  wire \NLW_blk000007fe/blk000007ff/blk00000802_Q31_UNCONNECTED ;
  wire \NLW_blk00000852/blk00000853/blk00000856_Q31_UNCONNECTED ;
  wire \NLW_blk00000858/blk00000859/blk0000085c_Q15_UNCONNECTED ;
  wire \NLW_blk0000085e/blk0000085f/blk00000862_Q15_UNCONNECTED ;
  wire \NLW_blk000008e1/blk000008e2/blk000008e4_Q15_UNCONNECTED ;
  wire \NLW_blk000008e6/blk000008e7/blk000008e9_Q15_UNCONNECTED ;
  wire \NLW_blk000009cb/blk000009cc/blk000009d1_Q15_UNCONNECTED ;
  wire [8 : 0] NlwRenamedSig_OI_xn_index;
  wire [18 : 0] \U0/i_synth/non_floating_point.arch_c.xfft_inst/single_channel.datapath/output_selector_re/Q ;
  wire [18 : 0] \U0/i_synth/non_floating_point.arch_c.xfft_inst/single_channel.datapath/output_selector_im/Q ;
  assign
    xn_index[8] = NlwRenamedSig_OI_xn_index[8],
    xn_index[7] = NlwRenamedSig_OI_xn_index[7],
    xn_index[6] = NlwRenamedSig_OI_xn_index[6],
    xn_index[5] = NlwRenamedSig_OI_xn_index[5],
    xn_index[4] = NlwRenamedSig_OI_xn_index[4],
    xn_index[3] = NlwRenamedSig_OI_xn_index[3],
    xn_index[2] = NlwRenamedSig_OI_xn_index[2],
    xn_index[1] = NlwRenamedSig_OI_xn_index[1],
    xn_index[0] = NlwRenamedSig_OI_xn_index[0],
    xk_re[18] = \U0/i_synth/non_floating_point.arch_c.xfft_inst/single_channel.datapath/output_selector_re/Q [18],
    xk_re[17] = \U0/i_synth/non_floating_point.arch_c.xfft_inst/single_channel.datapath/output_selector_re/Q [17],
    xk_re[16] = \U0/i_synth/non_floating_point.arch_c.xfft_inst/single_channel.datapath/output_selector_re/Q [16],
    xk_re[15] = \U0/i_synth/non_floating_point.arch_c.xfft_inst/single_channel.datapath/output_selector_re/Q [15],
    xk_re[14] = \U0/i_synth/non_floating_point.arch_c.xfft_inst/single_channel.datapath/output_selector_re/Q [14],
    xk_re[13] = \U0/i_synth/non_floating_point.arch_c.xfft_inst/single_channel.datapath/output_selector_re/Q [13],
    xk_re[12] = \U0/i_synth/non_floating_point.arch_c.xfft_inst/single_channel.datapath/output_selector_re/Q [12],
    xk_re[11] = \U0/i_synth/non_floating_point.arch_c.xfft_inst/single_channel.datapath/output_selector_re/Q [11],
    xk_re[10] = \U0/i_synth/non_floating_point.arch_c.xfft_inst/single_channel.datapath/output_selector_re/Q [10],
    xk_re[9] = \U0/i_synth/non_floating_point.arch_c.xfft_inst/single_channel.datapath/output_selector_re/Q [9],
    xk_re[8] = \U0/i_synth/non_floating_point.arch_c.xfft_inst/single_channel.datapath/output_selector_re/Q [8],
    xk_re[7] = \U0/i_synth/non_floating_point.arch_c.xfft_inst/single_channel.datapath/output_selector_re/Q [7],
    xk_re[6] = \U0/i_synth/non_floating_point.arch_c.xfft_inst/single_channel.datapath/output_selector_re/Q [6],
    xk_re[5] = \U0/i_synth/non_floating_point.arch_c.xfft_inst/single_channel.datapath/output_selector_re/Q [5],
    xk_re[4] = \U0/i_synth/non_floating_point.arch_c.xfft_inst/single_channel.datapath/output_selector_re/Q [4],
    xk_re[3] = \U0/i_synth/non_floating_point.arch_c.xfft_inst/single_channel.datapath/output_selector_re/Q [3],
    xk_re[2] = \U0/i_synth/non_floating_point.arch_c.xfft_inst/single_channel.datapath/output_selector_re/Q [2],
    xk_re[1] = \U0/i_synth/non_floating_point.arch_c.xfft_inst/single_channel.datapath/output_selector_re/Q [1],
    xk_re[0] = \U0/i_synth/non_floating_point.arch_c.xfft_inst/single_channel.datapath/output_selector_re/Q [0],
    xk_im[18] = \U0/i_synth/non_floating_point.arch_c.xfft_inst/single_channel.datapath/output_selector_im/Q [18],
    xk_im[17] = \U0/i_synth/non_floating_point.arch_c.xfft_inst/single_channel.datapath/output_selector_im/Q [17],
    xk_im[16] = \U0/i_synth/non_floating_point.arch_c.xfft_inst/single_channel.datapath/output_selector_im/Q [16],
    xk_im[15] = \U0/i_synth/non_floating_point.arch_c.xfft_inst/single_channel.datapath/output_selector_im/Q [15],
    xk_im[14] = \U0/i_synth/non_floating_point.arch_c.xfft_inst/single_channel.datapath/output_selector_im/Q [14],
    xk_im[13] = \U0/i_synth/non_floating_point.arch_c.xfft_inst/single_channel.datapath/output_selector_im/Q [13],
    xk_im[12] = \U0/i_synth/non_floating_point.arch_c.xfft_inst/single_channel.datapath/output_selector_im/Q [12],
    xk_im[11] = \U0/i_synth/non_floating_point.arch_c.xfft_inst/single_channel.datapath/output_selector_im/Q [11],
    xk_im[10] = \U0/i_synth/non_floating_point.arch_c.xfft_inst/single_channel.datapath/output_selector_im/Q [10],
    xk_im[9] = \U0/i_synth/non_floating_point.arch_c.xfft_inst/single_channel.datapath/output_selector_im/Q [9],
    xk_im[8] = \U0/i_synth/non_floating_point.arch_c.xfft_inst/single_channel.datapath/output_selector_im/Q [8],
    xk_im[7] = \U0/i_synth/non_floating_point.arch_c.xfft_inst/single_channel.datapath/output_selector_im/Q [7],
    xk_im[6] = \U0/i_synth/non_floating_point.arch_c.xfft_inst/single_channel.datapath/output_selector_im/Q [6],
    xk_im[5] = \U0/i_synth/non_floating_point.arch_c.xfft_inst/single_channel.datapath/output_selector_im/Q [5],
    xk_im[4] = \U0/i_synth/non_floating_point.arch_c.xfft_inst/single_channel.datapath/output_selector_im/Q [4],
    xk_im[3] = \U0/i_synth/non_floating_point.arch_c.xfft_inst/single_channel.datapath/output_selector_im/Q [3],
    xk_im[2] = \U0/i_synth/non_floating_point.arch_c.xfft_inst/single_channel.datapath/output_selector_im/Q [2],
    xk_im[1] = \U0/i_synth/non_floating_point.arch_c.xfft_inst/single_channel.datapath/output_selector_im/Q [1],
    xk_im[0] = \U0/i_synth/non_floating_point.arch_c.xfft_inst/single_channel.datapath/output_selector_im/Q [0],
    rfd = \NlwRenamedSig_OI_U0/i_synth/non_floating_point.arch_c.xfft_inst/control/cntrl/loading_state/ORS ,
    busy = \NlwRenamedSig_OI_U0/i_synth/non_floating_point.arch_c.xfft_inst/control/cntrl/processing_state/ORS ,
    edone = \NlwRenamedSig_OI_U0/i_synth/non_floating_point.arch_c.xfft_inst/control/cntrl/process_state_r ,
    done = \U0/i_synth/non_floating_point.arch_c.xfft_inst/control/cntrl/done_pr_d_1 ;
  VCC   blk00000001 (
    .P(sig00000001)
  );
  GND   blk00000002 (
    .G(sig00000002)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000057 (
    .C(clk),
    .D(sig0000024c),
    .Q(sig000001af)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000058 (
    .C(clk),
    .D(sig0000024b),
    .Q(sig000001ae)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000059 (
    .C(clk),
    .D(sig0000024a),
    .Q(sig000001ad)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000005a (
    .C(clk),
    .D(sig00000249),
    .Q(sig000001ac)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000005b (
    .C(clk),
    .D(sig00000248),
    .Q(sig000001ab)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000005c (
    .C(clk),
    .D(sig00000247),
    .Q(sig000001aa)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000005d (
    .C(clk),
    .D(sig00000246),
    .Q(sig000001a9)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000005e (
    .C(clk),
    .D(sig00000245),
    .Q(sig000001a8)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000005f (
    .C(clk),
    .D(sig00000244),
    .Q(sig000001a7)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000060 (
    .C(clk),
    .D(sig00000243),
    .Q(sig000001a6)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000061 (
    .C(clk),
    .D(sig00000242),
    .Q(sig000001a5)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000062 (
    .C(clk),
    .D(sig00000241),
    .Q(sig000001a4)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000063 (
    .C(clk),
    .D(sig00000240),
    .Q(sig000001a3)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000064 (
    .C(clk),
    .D(sig0000023f),
    .Q(sig000001a2)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000065 (
    .C(clk),
    .D(sig0000023e),
    .Q(sig000001a1)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000066 (
    .C(clk),
    .D(sig0000023d),
    .Q(sig000001a0)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000067 (
    .C(clk),
    .D(sig0000023c),
    .Q(sig0000019f)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000068 (
    .C(clk),
    .D(sig0000023b),
    .Q(sig0000019e)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000069 (
    .C(clk),
    .D(sig0000023a),
    .Q(sig0000019d)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000006a (
    .C(clk),
    .D(sig00000239),
    .Q(sig0000019c)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000006b (
    .C(clk),
    .D(sig00000238),
    .Q(sig0000019b)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000006c (
    .C(clk),
    .D(sig00000237),
    .Q(sig0000019a)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000006d (
    .C(clk),
    .D(sig00000236),
    .Q(sig00000199)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000006e (
    .C(clk),
    .D(sig00000235),
    .Q(sig000001c6)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000006f (
    .C(clk),
    .D(sig00000234),
    .Q(sig000001c5)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000070 (
    .C(clk),
    .D(sig00000233),
    .Q(sig000001c4)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000071 (
    .C(clk),
    .D(sig00000232),
    .Q(sig000001c3)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000072 (
    .C(clk),
    .D(sig00000231),
    .Q(sig000001c2)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000073 (
    .C(clk),
    .D(sig00000230),
    .Q(sig000001c1)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000074 (
    .C(clk),
    .D(sig0000022f),
    .Q(sig000001c0)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000075 (
    .C(clk),
    .D(sig0000022e),
    .Q(sig000001bf)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000076 (
    .C(clk),
    .D(sig0000022d),
    .Q(sig000001be)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000077 (
    .C(clk),
    .D(sig0000022c),
    .Q(sig000001bd)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000078 (
    .C(clk),
    .D(sig0000022b),
    .Q(sig000001bc)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000079 (
    .C(clk),
    .D(sig0000022a),
    .Q(sig000001bb)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000007a (
    .C(clk),
    .D(sig00000229),
    .Q(sig000001ba)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000007b (
    .C(clk),
    .D(sig00000228),
    .Q(sig000001b9)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000007c (
    .C(clk),
    .D(sig00000227),
    .Q(sig000001b8)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000007d (
    .C(clk),
    .D(sig00000226),
    .Q(sig000001b7)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000007e (
    .C(clk),
    .D(sig00000225),
    .Q(sig000001b6)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000007f (
    .C(clk),
    .D(sig00000224),
    .Q(sig000001b5)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000080 (
    .C(clk),
    .D(sig00000223),
    .Q(sig000001b4)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000081 (
    .C(clk),
    .D(sig00000222),
    .Q(sig000001b3)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000082 (
    .C(clk),
    .D(sig00000221),
    .Q(sig000001b2)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000083 (
    .C(clk),
    .D(sig00000220),
    .Q(sig000001b1)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000084 (
    .C(clk),
    .D(sig0000021f),
    .Q(sig000001b0)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000085 (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000001),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig0000008e),
    .Q(sig00000273)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000086 (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000001),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig0000008d),
    .Q(sig00000274)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000087 (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000001),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig0000008c),
    .Q(sig00000275)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000088 (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000001),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig0000008b),
    .Q(sig00000276)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000089 (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000001),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig0000008a),
    .Q(sig00000277)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000008a (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000001),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig00000089),
    .Q(sig00000278)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000008b (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000001),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig00000088),
    .Q(sig00000279)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000008c (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000001),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig00000087),
    .Q(sig0000027a)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000008d (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000001),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig00000086),
    .Q(sig0000027b)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000008e (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000001),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig00000085),
    .Q(sig0000027c)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000008f (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000001),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig00000084),
    .Q(sig0000027d)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000090 (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000001),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig00000083),
    .Q(sig0000027e)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000091 (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000001),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig00000082),
    .Q(sig0000027f)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000092 (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000001),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig00000081),
    .Q(sig00000280)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000093 (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000001),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig00000080),
    .Q(sig00000281)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000094 (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000001),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig0000007f),
    .Q(sig00000282)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000095 (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000001),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig0000007e),
    .Q(sig00000283)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000096 (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000001),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig0000007d),
    .Q(sig00000284)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000097 (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000001),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig0000007c),
    .Q(sig00000285)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000098 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000273),
    .R(sig00000002),
    .Q(sig0000025f)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000099 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000274),
    .R(sig00000002),
    .Q(sig0000025e)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000009a (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000275),
    .R(sig00000002),
    .Q(sig0000025d)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000009b (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000276),
    .R(sig00000002),
    .Q(sig0000025c)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000009c (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000277),
    .R(sig00000002),
    .Q(sig0000025b)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000009d (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000278),
    .R(sig00000002),
    .Q(sig0000025a)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000009e (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000279),
    .R(sig00000002),
    .Q(sig00000259)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000009f (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000027a),
    .R(sig00000002),
    .Q(sig00000258)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000000a0 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000027b),
    .R(sig00000002),
    .Q(sig00000257)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000000a1 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000027c),
    .R(sig00000002),
    .Q(sig00000256)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000000a2 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000027d),
    .R(sig00000002),
    .Q(sig00000255)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000000a3 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000027e),
    .R(sig00000002),
    .Q(sig00000254)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000000a4 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000027f),
    .R(sig00000002),
    .Q(sig00000253)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000000a5 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000280),
    .R(sig00000002),
    .Q(sig00000252)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000000a6 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000281),
    .R(sig00000002),
    .Q(sig00000251)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000000a7 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000282),
    .R(sig00000002),
    .Q(sig00000250)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000000a8 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000283),
    .R(sig00000002),
    .Q(sig0000024f)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000000a9 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000284),
    .R(sig00000002),
    .Q(sig0000024e)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000000aa (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000285),
    .R(sig00000002),
    .Q(sig0000024d)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000000ab (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000001),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig0000007b),
    .Q(sig00000286)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000000ac (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000001),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig0000007a),
    .Q(sig00000287)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000000ad (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000001),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig00000079),
    .Q(sig00000288)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000000ae (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000001),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig00000078),
    .Q(sig00000289)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000000af (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000001),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig00000077),
    .Q(sig0000028a)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000000b0 (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000001),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig00000076),
    .Q(sig0000028b)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000000b1 (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000001),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig00000075),
    .Q(sig0000028c)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000000b2 (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000001),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig00000074),
    .Q(sig0000028d)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000000b3 (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000001),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig00000073),
    .Q(sig0000028e)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000000b4 (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000001),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig00000072),
    .Q(sig0000028f)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000000b5 (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000001),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig00000071),
    .Q(sig00000290)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000000b6 (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000001),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig00000070),
    .Q(sig00000291)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000000b7 (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000001),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig0000006f),
    .Q(sig00000292)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000000b8 (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000001),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig0000006e),
    .Q(sig00000293)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000000b9 (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000001),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig0000006d),
    .Q(sig00000294)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000000ba (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000001),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig0000006c),
    .Q(sig00000295)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000000bb (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000001),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig0000006b),
    .Q(sig00000296)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000000bc (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000001),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig0000006a),
    .Q(sig00000297)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000000bd (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000001),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig00000069),
    .Q(sig00000298)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000000be (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000286),
    .R(sig00000002),
    .Q(sig00000272)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000000bf (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000287),
    .R(sig00000002),
    .Q(sig00000271)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000000c0 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000288),
    .R(sig00000002),
    .Q(sig00000270)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000000c1 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000289),
    .R(sig00000002),
    .Q(sig0000026f)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000000c2 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000028a),
    .R(sig00000002),
    .Q(sig0000026e)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000000c3 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000028b),
    .R(sig00000002),
    .Q(sig0000026d)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000000c4 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000028c),
    .R(sig00000002),
    .Q(sig0000026c)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000000c5 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000028d),
    .R(sig00000002),
    .Q(sig0000026b)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000000c6 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000028e),
    .R(sig00000002),
    .Q(sig0000026a)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000000c7 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000028f),
    .R(sig00000002),
    .Q(sig00000269)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000000c8 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000290),
    .R(sig00000002),
    .Q(sig00000268)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000000c9 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000291),
    .R(sig00000002),
    .Q(sig00000267)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000000ca (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000292),
    .R(sig00000002),
    .Q(sig00000266)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000000cb (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000293),
    .R(sig00000002),
    .Q(sig00000265)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000000cc (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000294),
    .R(sig00000002),
    .Q(sig00000264)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000000cd (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000295),
    .R(sig00000002),
    .Q(sig00000263)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000000ce (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000296),
    .R(sig00000002),
    .Q(sig00000262)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000000cf (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000297),
    .R(sig00000002),
    .Q(sig00000261)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000000d0 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000298),
    .R(sig00000002),
    .Q(sig00000260)
  );
  DSP48A1 #(
    .A0REG ( 1 ),
    .A1REG ( 1 ),
    .B0REG ( 1 ),
    .B1REG ( 1 ),
    .CARRYINREG ( 0 ),
    .CARRYINSEL ( "OPMODE5" ),
    .CREG ( 1 ),
    .DREG ( 0 ),
    .MREG ( 1 ),
    .OPMODEREG ( 0 ),
    .PREG ( 1 ),
    .RSTTYPE ( "SYNC" ),
    .CARRYOUTREG ( 0 ))
  blk000000d1 (
    .CECARRYIN(sig00000002),
    .RSTC(sig00000002),
    .RSTCARRYIN(sig00000002),
    .CED(sig00000002),
    .RSTD(sig00000002),
    .CEOPMODE(sig00000002),
    .CEC(sig00000001),
    .CARRYOUTF(NLW_blk000000d1_CARRYOUTF_UNCONNECTED),
    .RSTOPMODE(sig00000002),
    .RSTM(sig00000002),
    .CLK(clk),
    .RSTB(sig00000002),
    .CEM(sig00000001),
    .CEB(sig00000001),
    .CARRYIN(sig00000002),
    .CEP(sig00000001),
    .CEA(sig00000001),
    .CARRYOUT(NLW_blk000000d1_CARRYOUT_UNCONNECTED),
    .RSTA(sig00000002),
    .RSTP(sig00000002),
    .B({sig00000320, sig00000320, sig00000320, sig00000320, sig00000320, sig00000320, sig00000320, sig00000320, sig00000320, sig00000329, sig0000032a
, sig0000032b, sig0000032c, sig0000032d, sig0000032e, sig0000032f, sig00000330, sig00000331}),
    .BCOUT({sig00000299, sig0000029a, sig0000029b, sig0000029c, sig0000029d, sig0000029e, sig0000029f, sig000002a0, sig000002a1, sig000002a2,
sig000002a3, sig000002a4, sig000002a5, sig000002a6, sig000002a7, sig000002a8, sig000002a9, sig000002aa}),
    .PCIN({sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002,
sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002,
sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002,
sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002,
sig00000002, sig00000002, sig00000002, sig00000002, sig00000002}),
    .C({sig00000405, sig00000405, sig00000405, sig00000405, sig00000405, sig00000405, sig00000405, sig00000405, sig00000405, sig00000405, sig00000405
, sig00000405, sig00000405, sig00000405, sig00000405, sig00000405, sig00000405, sig00000405, sig00000405, sig00000406, sig00000407, sig00000408,
sig00000409, sig0000040a, sig0000040b, sig0000040c, sig0000040d, sig0000040e, sig0000040f, sig00000410, sig00000411, sig000004b4, sig000004b3,
sig000004b2, sig000004b1, sig000004b0, sig000004af, sig000004ae, sig000004ad, sig000004ac, sig000004ab, sig000004aa, sig000004a9, sig000004a8,
sig000004a7, sig000004a6, sig000004a5, sig000004a4}),
    .P({sig000002bc, sig000002bd, sig000002be, sig000002bf, sig000002c0, sig000002c1, sig000002c2, sig000002c3, sig000002c4, sig000002c5, sig000002c6
, sig000002c7, sig000002c8, sig000002c9, sig000002ca, sig000002cb, sig000002cc, sig000002cd, sig000002ce, sig000002cf, sig000002d0, sig000002d1,
sig000002d2, sig000002d3, sig000002d4, sig000002d5, sig000002d6, sig000002d7, sig000002d8, sig000002d9, sig000002da, sig000002ab, sig000002ac,
sig000002ad, sig000002ae, sig000002af, sig000002b0, sig000002b1, sig000002b2, sig000002b3, sig000002b4, sig000002b5, sig000002b6, sig000002b7,
sig000002b8, sig000002b9, sig000002ba, sig000002bb}),
    .OPMODE({sig00000002, sig00000002, sig00000002, sig00000002, sig00000001, sig00000001, sig00000002, sig00000001}),
    .D({sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002
, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002}),
    .PCOUT({sig000002db, sig000002dc, sig000002dd, sig000002de, sig000002df, sig000002e0, sig000002e1, sig000002e2, sig000002e3, sig000002e4,
sig000002e5, sig000002e6, sig000002e7, sig000002e8, sig000002e9, sig000002ea, sig000002eb, sig000002ec, sig000002ed, sig000002ee, sig000002ef,
sig000002f0, sig000002f1, sig000002f2, sig000002f3, sig000002f4, sig000002f5, sig000002f6, sig000002f7, sig000002f8, sig000002f9, sig000002fa,
sig000002fb, sig000002fc, sig000002fd, sig000002fe, sig000002ff, sig00000300, sig00000301, sig00000302, sig00000303, sig00000304, sig00000305,
sig00000306, sig00000307, sig00000308, sig00000309, sig0000030a}),
    .A({sig00000002, sig0000030c, sig0000030d, sig0000030e, sig0000030f, sig00000310, sig00000311, sig00000312, sig00000313, sig00000314, sig00000315
, sig00000316, sig00000317, sig00000318, sig00000319, sig0000031a, sig0000031b, sig0000031c}),
    .M({\NLW_blk000000d1_M<35>_UNCONNECTED , \NLW_blk000000d1_M<34>_UNCONNECTED , \NLW_blk000000d1_M<33>_UNCONNECTED ,
\NLW_blk000000d1_M<32>_UNCONNECTED , \NLW_blk000000d1_M<31>_UNCONNECTED , \NLW_blk000000d1_M<30>_UNCONNECTED , \NLW_blk000000d1_M<29>_UNCONNECTED ,
\NLW_blk000000d1_M<28>_UNCONNECTED , \NLW_blk000000d1_M<27>_UNCONNECTED , \NLW_blk000000d1_M<26>_UNCONNECTED , \NLW_blk000000d1_M<25>_UNCONNECTED ,
\NLW_blk000000d1_M<24>_UNCONNECTED , \NLW_blk000000d1_M<23>_UNCONNECTED , \NLW_blk000000d1_M<22>_UNCONNECTED , \NLW_blk000000d1_M<21>_UNCONNECTED ,
\NLW_blk000000d1_M<20>_UNCONNECTED , \NLW_blk000000d1_M<19>_UNCONNECTED , \NLW_blk000000d1_M<18>_UNCONNECTED , \NLW_blk000000d1_M<17>_UNCONNECTED ,
\NLW_blk000000d1_M<16>_UNCONNECTED , \NLW_blk000000d1_M<15>_UNCONNECTED , \NLW_blk000000d1_M<14>_UNCONNECTED , \NLW_blk000000d1_M<13>_UNCONNECTED ,
\NLW_blk000000d1_M<12>_UNCONNECTED , \NLW_blk000000d1_M<11>_UNCONNECTED , \NLW_blk000000d1_M<10>_UNCONNECTED , \NLW_blk000000d1_M<9>_UNCONNECTED ,
\NLW_blk000000d1_M<8>_UNCONNECTED , \NLW_blk000000d1_M<7>_UNCONNECTED , \NLW_blk000000d1_M<6>_UNCONNECTED , \NLW_blk000000d1_M<5>_UNCONNECTED ,
\NLW_blk000000d1_M<4>_UNCONNECTED , \NLW_blk000000d1_M<3>_UNCONNECTED , \NLW_blk000000d1_M<2>_UNCONNECTED , \NLW_blk000000d1_M<1>_UNCONNECTED ,
\NLW_blk000000d1_M<0>_UNCONNECTED })
  );
  DSP48A1 #(
    .A0REG ( 1 ),
    .A1REG ( 1 ),
    .B0REG ( 1 ),
    .B1REG ( 1 ),
    .CARRYINREG ( 0 ),
    .CARRYINSEL ( "OPMODE5" ),
    .CREG ( 1 ),
    .DREG ( 0 ),
    .MREG ( 1 ),
    .OPMODEREG ( 0 ),
    .PREG ( 1 ),
    .RSTTYPE ( "SYNC" ),
    .CARRYOUTREG ( 0 ))
  blk000000d2 (
    .CECARRYIN(sig00000002),
    .RSTC(sig00000002),
    .RSTCARRYIN(sig00000002),
    .CED(sig00000002),
    .RSTD(sig00000002),
    .CEOPMODE(sig00000002),
    .CEC(sig00000001),
    .CARRYOUTF(NLW_blk000000d2_CARRYOUTF_UNCONNECTED),
    .RSTOPMODE(sig00000002),
    .RSTM(sig00000002),
    .CLK(clk),
    .RSTB(sig00000002),
    .CEM(sig00000001),
    .CEB(sig00000001),
    .CARRYIN(sig00000002),
    .CEP(sig00000001),
    .CEA(sig00000001),
    .CARRYOUT(NLW_blk000000d2_CARRYOUT_UNCONNECTED),
    .RSTA(sig00000002),
    .RSTP(sig00000002),
    .B({sig00000299, sig0000029a, sig0000029b, sig0000029c, sig0000029d, sig0000029e, sig0000029f, sig000002a0, sig000002a1, sig000002a2, sig000002a3
, sig000002a4, sig000002a5, sig000002a6, sig000002a7, sig000002a8, sig000002a9, sig000002aa}),
    .BCOUT({\NLW_blk000000d2_BCOUT<17>_UNCONNECTED , \NLW_blk000000d2_BCOUT<16>_UNCONNECTED , \NLW_blk000000d2_BCOUT<15>_UNCONNECTED ,
\NLW_blk000000d2_BCOUT<14>_UNCONNECTED , \NLW_blk000000d2_BCOUT<13>_UNCONNECTED , \NLW_blk000000d2_BCOUT<12>_UNCONNECTED ,
\NLW_blk000000d2_BCOUT<11>_UNCONNECTED , \NLW_blk000000d2_BCOUT<10>_UNCONNECTED , \NLW_blk000000d2_BCOUT<9>_UNCONNECTED ,
\NLW_blk000000d2_BCOUT<8>_UNCONNECTED , \NLW_blk000000d2_BCOUT<7>_UNCONNECTED , \NLW_blk000000d2_BCOUT<6>_UNCONNECTED ,
\NLW_blk000000d2_BCOUT<5>_UNCONNECTED , \NLW_blk000000d2_BCOUT<4>_UNCONNECTED , \NLW_blk000000d2_BCOUT<3>_UNCONNECTED ,
\NLW_blk000000d2_BCOUT<2>_UNCONNECTED , \NLW_blk000000d2_BCOUT<1>_UNCONNECTED , \NLW_blk000000d2_BCOUT<0>_UNCONNECTED }),
    .PCIN({sig000002db, sig000002dc, sig000002dd, sig000002de, sig000002df, sig000002e0, sig000002e1, sig000002e2, sig000002e3, sig000002e4,
sig000002e5, sig000002e6, sig000002e7, sig000002e8, sig000002e9, sig000002ea, sig000002eb, sig000002ec, sig000002ed, sig000002ee, sig000002ef,
sig000002f0, sig000002f1, sig000002f2, sig000002f3, sig000002f4, sig000002f5, sig000002f6, sig000002f7, sig000002f8, sig000002f9, sig000002fa,
sig000002fb, sig000002fc, sig000002fd, sig000002fe, sig000002ff, sig00000300, sig00000301, sig00000302, sig00000303, sig00000304, sig00000305,
sig00000306, sig00000307, sig00000308, sig00000309, sig0000030a}),
    .C({sig000002bc, sig000002bc, sig000002bc, sig000002bc, sig000002bc, sig000002bc, sig000002bc, sig000002bc, sig000002bc, sig000002bc, sig000002bc
, sig000002bc, sig000002bc, sig000002bc, sig000002bc, sig000002bc, sig000002bc, sig000002bc, sig000002bd, sig000002be, sig000002bf, sig000002c0,
sig000002c1, sig000002c2, sig000002c3, sig000002c4, sig000002c5, sig000002c6, sig000002c7, sig000002c8, sig000002c9, sig000002ca, sig000002cb,
sig000002cc, sig000002cd, sig000002ce, sig000002cf, sig000002d0, sig000002d1, sig000002d2, sig000002d3, sig000002d4, sig000002d5, sig000002d6,
sig000002d7, sig000002d8, sig000002d9, sig000002da}),
    .P({\NLW_blk000000d2_P<47>_UNCONNECTED , \NLW_blk000000d2_P<46>_UNCONNECTED , \NLW_blk000000d2_P<45>_UNCONNECTED ,
\NLW_blk000000d2_P<44>_UNCONNECTED , \NLW_blk000000d2_P<43>_UNCONNECTED , \NLW_blk000000d2_P<42>_UNCONNECTED , \NLW_blk000000d2_P<41>_UNCONNECTED ,
\NLW_blk000000d2_P<40>_UNCONNECTED , \NLW_blk000000d2_P<39>_UNCONNECTED , \NLW_blk000000d2_P<38>_UNCONNECTED , \NLW_blk000000d2_P<37>_UNCONNECTED ,
\NLW_blk000000d2_P<36>_UNCONNECTED , sig00000332, sig00000333, sig00000334, sig00000335, sig00000336, sig00000337, sig00000338, sig00000339,
sig0000033a, sig0000033b, sig0000033c, sig0000033d, sig0000033e, sig0000033f, sig00000340, sig00000341, sig00000342, sig00000343, sig00000344,
sig00000345, sig00000346, sig00000347, sig00000348, sig00000349, sig0000034a, sig00000235, sig00000234, sig00000233, sig00000232, sig00000231,
sig00000230, sig0000022f, sig0000022e, sig0000022d, sig0000022c, sig0000022b}),
    .OPMODE({sig00000002, sig00000002, sig00000002, sig00000002, sig00000001, sig00000001, sig00000002, sig00000001}),
    .D({sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002
, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002}),
    .PCOUT({\NLW_blk000000d2_PCOUT<47>_UNCONNECTED , \NLW_blk000000d2_PCOUT<46>_UNCONNECTED , \NLW_blk000000d2_PCOUT<45>_UNCONNECTED ,
\NLW_blk000000d2_PCOUT<44>_UNCONNECTED , \NLW_blk000000d2_PCOUT<43>_UNCONNECTED , \NLW_blk000000d2_PCOUT<42>_UNCONNECTED ,
\NLW_blk000000d2_PCOUT<41>_UNCONNECTED , \NLW_blk000000d2_PCOUT<40>_UNCONNECTED , \NLW_blk000000d2_PCOUT<39>_UNCONNECTED ,
\NLW_blk000000d2_PCOUT<38>_UNCONNECTED , \NLW_blk000000d2_PCOUT<37>_UNCONNECTED , \NLW_blk000000d2_PCOUT<36>_UNCONNECTED ,
\NLW_blk000000d2_PCOUT<35>_UNCONNECTED , \NLW_blk000000d2_PCOUT<34>_UNCONNECTED , \NLW_blk000000d2_PCOUT<33>_UNCONNECTED ,
\NLW_blk000000d2_PCOUT<32>_UNCONNECTED , \NLW_blk000000d2_PCOUT<31>_UNCONNECTED , \NLW_blk000000d2_PCOUT<30>_UNCONNECTED ,
\NLW_blk000000d2_PCOUT<29>_UNCONNECTED , \NLW_blk000000d2_PCOUT<28>_UNCONNECTED , \NLW_blk000000d2_PCOUT<27>_UNCONNECTED ,
\NLW_blk000000d2_PCOUT<26>_UNCONNECTED , \NLW_blk000000d2_PCOUT<25>_UNCONNECTED , \NLW_blk000000d2_PCOUT<24>_UNCONNECTED ,
\NLW_blk000000d2_PCOUT<23>_UNCONNECTED , \NLW_blk000000d2_PCOUT<22>_UNCONNECTED , \NLW_blk000000d2_PCOUT<21>_UNCONNECTED ,
\NLW_blk000000d2_PCOUT<20>_UNCONNECTED , \NLW_blk000000d2_PCOUT<19>_UNCONNECTED , \NLW_blk000000d2_PCOUT<18>_UNCONNECTED ,
\NLW_blk000000d2_PCOUT<17>_UNCONNECTED , \NLW_blk000000d2_PCOUT<16>_UNCONNECTED , \NLW_blk000000d2_PCOUT<15>_UNCONNECTED ,
\NLW_blk000000d2_PCOUT<14>_UNCONNECTED , \NLW_blk000000d2_PCOUT<13>_UNCONNECTED , \NLW_blk000000d2_PCOUT<12>_UNCONNECTED ,
\NLW_blk000000d2_PCOUT<11>_UNCONNECTED , \NLW_blk000000d2_PCOUT<10>_UNCONNECTED , \NLW_blk000000d2_PCOUT<9>_UNCONNECTED ,
\NLW_blk000000d2_PCOUT<8>_UNCONNECTED , \NLW_blk000000d2_PCOUT<7>_UNCONNECTED , \NLW_blk000000d2_PCOUT<6>_UNCONNECTED ,
\NLW_blk000000d2_PCOUT<5>_UNCONNECTED , \NLW_blk000000d2_PCOUT<4>_UNCONNECTED , \NLW_blk000000d2_PCOUT<3>_UNCONNECTED ,
\NLW_blk000000d2_PCOUT<2>_UNCONNECTED , \NLW_blk000000d2_PCOUT<1>_UNCONNECTED , \NLW_blk000000d2_PCOUT<0>_UNCONNECTED }),
    .A({sig0000031d, sig0000031d, sig0000031d, sig0000031d, sig0000031d, sig0000031d, sig0000031d, sig0000031d, sig0000031d, sig0000031d, sig0000031d
, sig0000031d, sig0000031d, sig0000031d, sig0000031d, sig0000031d, sig0000031e, sig0000031f}),
    .M({\NLW_blk000000d2_M<35>_UNCONNECTED , \NLW_blk000000d2_M<34>_UNCONNECTED , \NLW_blk000000d2_M<33>_UNCONNECTED ,
\NLW_blk000000d2_M<32>_UNCONNECTED , \NLW_blk000000d2_M<31>_UNCONNECTED , \NLW_blk000000d2_M<30>_UNCONNECTED , \NLW_blk000000d2_M<29>_UNCONNECTED ,
\NLW_blk000000d2_M<28>_UNCONNECTED , \NLW_blk000000d2_M<27>_UNCONNECTED , \NLW_blk000000d2_M<26>_UNCONNECTED , \NLW_blk000000d2_M<25>_UNCONNECTED ,
\NLW_blk000000d2_M<24>_UNCONNECTED , \NLW_blk000000d2_M<23>_UNCONNECTED , \NLW_blk000000d2_M<22>_UNCONNECTED , \NLW_blk000000d2_M<21>_UNCONNECTED ,
\NLW_blk000000d2_M<20>_UNCONNECTED , \NLW_blk000000d2_M<19>_UNCONNECTED , \NLW_blk000000d2_M<18>_UNCONNECTED , \NLW_blk000000d2_M<17>_UNCONNECTED ,
\NLW_blk000000d2_M<16>_UNCONNECTED , \NLW_blk000000d2_M<15>_UNCONNECTED , \NLW_blk000000d2_M<14>_UNCONNECTED , \NLW_blk000000d2_M<13>_UNCONNECTED ,
\NLW_blk000000d2_M<12>_UNCONNECTED , \NLW_blk000000d2_M<11>_UNCONNECTED , \NLW_blk000000d2_M<10>_UNCONNECTED , \NLW_blk000000d2_M<9>_UNCONNECTED ,
\NLW_blk000000d2_M<8>_UNCONNECTED , \NLW_blk000000d2_M<7>_UNCONNECTED , \NLW_blk000000d2_M<6>_UNCONNECTED , \NLW_blk000000d2_M<5>_UNCONNECTED ,
\NLW_blk000000d2_M<4>_UNCONNECTED , \NLW_blk000000d2_M<3>_UNCONNECTED , \NLW_blk000000d2_M<2>_UNCONNECTED , \NLW_blk000000d2_M<1>_UNCONNECTED ,
\NLW_blk000000d2_M<0>_UNCONNECTED })
  );
  DSP48A1 #(
    .A0REG ( 1 ),
    .A1REG ( 1 ),
    .B0REG ( 1 ),
    .B1REG ( 1 ),
    .CARRYINREG ( 0 ),
    .CARRYINSEL ( "OPMODE5" ),
    .CREG ( 0 ),
    .DREG ( 1 ),
    .MREG ( 1 ),
    .OPMODEREG ( 0 ),
    .PREG ( 1 ),
    .RSTTYPE ( "SYNC" ),
    .CARRYOUTREG ( 0 ))
  blk000000d3 (
    .CECARRYIN(sig00000002),
    .RSTC(sig00000002),
    .RSTCARRYIN(sig00000002),
    .CED(sig00000001),
    .RSTD(sig00000002),
    .CEOPMODE(sig00000002),
    .CEC(sig00000002),
    .CARRYOUTF(NLW_blk000000d3_CARRYOUTF_UNCONNECTED),
    .RSTOPMODE(sig00000002),
    .RSTM(sig00000002),
    .CLK(clk),
    .RSTB(sig00000002),
    .CEM(sig00000001),
    .CEB(sig00000001),
    .CARRYIN(sig00000002),
    .CEP(sig00000001),
    .CEA(sig00000001),
    .CARRYOUT(NLW_blk000000d3_CARRYOUT_UNCONNECTED),
    .RSTA(sig00000002),
    .RSTP(sig00000002),
    .B({sig000003dc, sig000003dc, sig000003dc, sig000003dc, sig000003dc, sig000003dc, sig000003dc, sig000003dc, sig000003dc, sig000003e5, sig000003e6
, sig000003e7, sig000003e8, sig000003e9, sig000003ea, sig000003eb, sig000003ec, sig000003ed}),
    .BCOUT({sig00000356, sig00000357, sig00000358, sig00000359, sig0000035a, sig0000035b, sig0000035c, sig0000035d, sig0000035e, sig0000035f,
sig00000360, sig00000361, sig00000362, sig00000363, sig00000364, sig00000365, sig00000366, sig00000367}),
    .PCIN({sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002,
sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002,
sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002,
sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002,
sig00000002, sig00000002, sig00000002, sig00000002, sig00000002}),
    .C({sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002
, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002,
sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002,
sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002,
sig00000001, sig00000001, sig00000001, sig00000001}),
    .P({sig00000379, sig0000037a, sig0000037b, sig0000037c, sig0000037d, sig0000037e, sig0000037f, sig00000380, sig00000381, sig00000382, sig00000383
, sig00000384, sig00000385, sig00000386, sig00000387, sig00000388, sig00000389, sig0000038a, sig0000038b, sig0000038c, sig0000038d, sig0000038e,
sig0000038f, sig00000390, sig00000391, sig00000392, sig00000393, sig00000394, sig00000395, sig00000396, sig00000397, sig00000368, sig00000369,
sig0000036a, sig0000036b, sig0000036c, sig0000036d, sig0000036e, sig0000036f, sig00000370, sig00000371, sig00000372, sig00000373, sig00000374,
sig00000375, sig00000376, sig00000377, sig00000378}),
    .OPMODE({sig00000002, sig00000002, sig00000002, sig00000001, sig00000001, sig00000001, sig00000002, sig00000001}),
    .D({sig000004e9, sig000004e9, sig000004e9, sig000004e9, sig000004e9, sig000004e9, sig000004e9, sig000004e9, sig000004e9, sig000004e8, sig000004e7
, sig000004e6, sig000004e5, sig000004e4, sig000004e3, sig000004e2, sig000004e1, sig000004e0}),
    .PCOUT({sig00000398, sig00000399, sig0000039a, sig0000039b, sig0000039c, sig0000039d, sig0000039e, sig0000039f, sig000003a0, sig000003a1,
sig000003a2, sig000003a3, sig000003a4, sig000003a5, sig000003a6, sig000003a7, sig000003a8, sig000003a9, sig000003aa, sig000003ab, sig000003ac,
sig000003ad, sig000003ae, sig000003af, sig000003b0, sig000003b1, sig000003b2, sig000003b3, sig000003b4, sig000003b5, sig000003b6, sig000003b7,
sig000003b8, sig000003b9, sig000003ba, sig000003bb, sig000003bc, sig000003bd, sig000003be, sig000003bf, sig000003c0, sig000003c1, sig000003c2,
sig000003c3, sig000003c4, sig000003c5, sig000003c6, sig000003c7}),
    .A({sig00000002, sig000003c9, sig000003ca, sig000003cb, sig000003cc, sig000003cd, sig000003ce, sig000003cf, sig000003d0, sig000003d1, sig000003d2
, sig000003d3, sig000003d4, sig000003d5, sig000003d6, sig000003d7, sig000003d8, sig000003d9}),
    .M({\NLW_blk000000d3_M<35>_UNCONNECTED , \NLW_blk000000d3_M<34>_UNCONNECTED , \NLW_blk000000d3_M<33>_UNCONNECTED ,
\NLW_blk000000d3_M<32>_UNCONNECTED , \NLW_blk000000d3_M<31>_UNCONNECTED , \NLW_blk000000d3_M<30>_UNCONNECTED , \NLW_blk000000d3_M<29>_UNCONNECTED ,
\NLW_blk000000d3_M<28>_UNCONNECTED , \NLW_blk000000d3_M<27>_UNCONNECTED , \NLW_blk000000d3_M<26>_UNCONNECTED , \NLW_blk000000d3_M<25>_UNCONNECTED ,
\NLW_blk000000d3_M<24>_UNCONNECTED , \NLW_blk000000d3_M<23>_UNCONNECTED , \NLW_blk000000d3_M<22>_UNCONNECTED , \NLW_blk000000d3_M<21>_UNCONNECTED ,
\NLW_blk000000d3_M<20>_UNCONNECTED , \NLW_blk000000d3_M<19>_UNCONNECTED , \NLW_blk000000d3_M<18>_UNCONNECTED , \NLW_blk000000d3_M<17>_UNCONNECTED ,
\NLW_blk000000d3_M<16>_UNCONNECTED , \NLW_blk000000d3_M<15>_UNCONNECTED , \NLW_blk000000d3_M<14>_UNCONNECTED , \NLW_blk000000d3_M<13>_UNCONNECTED ,
\NLW_blk000000d3_M<12>_UNCONNECTED , \NLW_blk000000d3_M<11>_UNCONNECTED , \NLW_blk000000d3_M<10>_UNCONNECTED , \NLW_blk000000d3_M<9>_UNCONNECTED ,
\NLW_blk000000d3_M<8>_UNCONNECTED , \NLW_blk000000d3_M<7>_UNCONNECTED , \NLW_blk000000d3_M<6>_UNCONNECTED , \NLW_blk000000d3_M<5>_UNCONNECTED ,
\NLW_blk000000d3_M<4>_UNCONNECTED , \NLW_blk000000d3_M<3>_UNCONNECTED , \NLW_blk000000d3_M<2>_UNCONNECTED , \NLW_blk000000d3_M<1>_UNCONNECTED ,
\NLW_blk000000d3_M<0>_UNCONNECTED })
  );
  DSP48A1 #(
    .A0REG ( 1 ),
    .A1REG ( 1 ),
    .B0REG ( 1 ),
    .B1REG ( 1 ),
    .CARRYINREG ( 0 ),
    .CARRYINSEL ( "OPMODE5" ),
    .CREG ( 1 ),
    .DREG ( 0 ),
    .MREG ( 1 ),
    .OPMODEREG ( 0 ),
    .PREG ( 1 ),
    .RSTTYPE ( "SYNC" ),
    .CARRYOUTREG ( 0 ))
  blk000000d4 (
    .CECARRYIN(sig00000002),
    .RSTC(sig00000002),
    .RSTCARRYIN(sig00000002),
    .CED(sig00000002),
    .RSTD(sig00000002),
    .CEOPMODE(sig00000002),
    .CEC(sig00000001),
    .CARRYOUTF(NLW_blk000000d4_CARRYOUTF_UNCONNECTED),
    .RSTOPMODE(sig00000002),
    .RSTM(sig00000002),
    .CLK(clk),
    .RSTB(sig00000002),
    .CEM(sig00000001),
    .CEB(sig00000001),
    .CARRYIN(sig00000002),
    .CEP(sig00000001),
    .CEA(sig00000001),
    .CARRYOUT(NLW_blk000000d4_CARRYOUT_UNCONNECTED),
    .RSTA(sig00000002),
    .RSTP(sig00000002),
    .B({sig00000356, sig00000357, sig00000358, sig00000359, sig0000035a, sig0000035b, sig0000035c, sig0000035d, sig0000035e, sig0000035f, sig00000360
, sig00000361, sig00000362, sig00000363, sig00000364, sig00000365, sig00000366, sig00000367}),
    .BCOUT({\NLW_blk000000d4_BCOUT<17>_UNCONNECTED , \NLW_blk000000d4_BCOUT<16>_UNCONNECTED , \NLW_blk000000d4_BCOUT<15>_UNCONNECTED ,
\NLW_blk000000d4_BCOUT<14>_UNCONNECTED , \NLW_blk000000d4_BCOUT<13>_UNCONNECTED , \NLW_blk000000d4_BCOUT<12>_UNCONNECTED ,
\NLW_blk000000d4_BCOUT<11>_UNCONNECTED , \NLW_blk000000d4_BCOUT<10>_UNCONNECTED , \NLW_blk000000d4_BCOUT<9>_UNCONNECTED ,
\NLW_blk000000d4_BCOUT<8>_UNCONNECTED , \NLW_blk000000d4_BCOUT<7>_UNCONNECTED , \NLW_blk000000d4_BCOUT<6>_UNCONNECTED ,
\NLW_blk000000d4_BCOUT<5>_UNCONNECTED , \NLW_blk000000d4_BCOUT<4>_UNCONNECTED , \NLW_blk000000d4_BCOUT<3>_UNCONNECTED ,
\NLW_blk000000d4_BCOUT<2>_UNCONNECTED , \NLW_blk000000d4_BCOUT<1>_UNCONNECTED , \NLW_blk000000d4_BCOUT<0>_UNCONNECTED }),
    .PCIN({sig00000398, sig00000399, sig0000039a, sig0000039b, sig0000039c, sig0000039d, sig0000039e, sig0000039f, sig000003a0, sig000003a1,
sig000003a2, sig000003a3, sig000003a4, sig000003a5, sig000003a6, sig000003a7, sig000003a8, sig000003a9, sig000003aa, sig000003ab, sig000003ac,
sig000003ad, sig000003ae, sig000003af, sig000003b0, sig000003b1, sig000003b2, sig000003b3, sig000003b4, sig000003b5, sig000003b6, sig000003b7,
sig000003b8, sig000003b9, sig000003ba, sig000003bb, sig000003bc, sig000003bd, sig000003be, sig000003bf, sig000003c0, sig000003c1, sig000003c2,
sig000003c3, sig000003c4, sig000003c5, sig000003c6, sig000003c7}),
    .C({sig00000379, sig00000379, sig00000379, sig00000379, sig00000379, sig00000379, sig00000379, sig00000379, sig00000379, sig00000379, sig00000379
, sig00000379, sig00000379, sig00000379, sig00000379, sig00000379, sig00000379, sig00000379, sig0000037a, sig0000037b, sig0000037c, sig0000037d,
sig0000037e, sig0000037f, sig00000380, sig00000381, sig00000382, sig00000383, sig00000384, sig00000385, sig00000386, sig00000387, sig00000388,
sig00000389, sig0000038a, sig0000038b, sig0000038c, sig0000038d, sig0000038e, sig0000038f, sig00000390, sig00000391, sig00000392, sig00000393,
sig00000394, sig00000395, sig00000396, sig00000397}),
    .P({\NLW_blk000000d4_P<47>_UNCONNECTED , \NLW_blk000000d4_P<46>_UNCONNECTED , \NLW_blk000000d4_P<45>_UNCONNECTED ,
\NLW_blk000000d4_P<44>_UNCONNECTED , \NLW_blk000000d4_P<43>_UNCONNECTED , \NLW_blk000000d4_P<42>_UNCONNECTED , \NLW_blk000000d4_P<41>_UNCONNECTED ,
\NLW_blk000000d4_P<40>_UNCONNECTED , \NLW_blk000000d4_P<39>_UNCONNECTED , \NLW_blk000000d4_P<38>_UNCONNECTED , \NLW_blk000000d4_P<37>_UNCONNECTED ,
\NLW_blk000000d4_P<36>_UNCONNECTED , sig000003ee, sig000003ef, sig000003f0, sig000003f1, sig000003f2, sig000003f3, sig000003f4, sig000003f5,
sig000003f6, sig000003f7, sig000003f8, sig000003f9, sig000003fa, sig000003fb, sig000003fc, sig000003fd, sig000003fe, sig000003ff, sig00000400,
sig00000401, sig00000402, sig00000403, sig00000404, sig00000405, sig00000406, sig00000407, sig00000408, sig00000409, sig0000040a, sig0000040b,
sig0000040c, sig0000040d, sig0000040e, sig0000040f, sig00000410, sig00000411}),
    .OPMODE({sig00000002, sig00000002, sig00000002, sig00000002, sig00000001, sig00000001, sig00000002, sig00000001}),
    .D({sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002
, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002}),
    .PCOUT({\NLW_blk000000d4_PCOUT<47>_UNCONNECTED , \NLW_blk000000d4_PCOUT<46>_UNCONNECTED , \NLW_blk000000d4_PCOUT<45>_UNCONNECTED ,
\NLW_blk000000d4_PCOUT<44>_UNCONNECTED , \NLW_blk000000d4_PCOUT<43>_UNCONNECTED , \NLW_blk000000d4_PCOUT<42>_UNCONNECTED ,
\NLW_blk000000d4_PCOUT<41>_UNCONNECTED , \NLW_blk000000d4_PCOUT<40>_UNCONNECTED , \NLW_blk000000d4_PCOUT<39>_UNCONNECTED ,
\NLW_blk000000d4_PCOUT<38>_UNCONNECTED , \NLW_blk000000d4_PCOUT<37>_UNCONNECTED , \NLW_blk000000d4_PCOUT<36>_UNCONNECTED ,
\NLW_blk000000d4_PCOUT<35>_UNCONNECTED , \NLW_blk000000d4_PCOUT<34>_UNCONNECTED , \NLW_blk000000d4_PCOUT<33>_UNCONNECTED ,
\NLW_blk000000d4_PCOUT<32>_UNCONNECTED , \NLW_blk000000d4_PCOUT<31>_UNCONNECTED , \NLW_blk000000d4_PCOUT<30>_UNCONNECTED ,
\NLW_blk000000d4_PCOUT<29>_UNCONNECTED , \NLW_blk000000d4_PCOUT<28>_UNCONNECTED , \NLW_blk000000d4_PCOUT<27>_UNCONNECTED ,
\NLW_blk000000d4_PCOUT<26>_UNCONNECTED , \NLW_blk000000d4_PCOUT<25>_UNCONNECTED , \NLW_blk000000d4_PCOUT<24>_UNCONNECTED ,
\NLW_blk000000d4_PCOUT<23>_UNCONNECTED , \NLW_blk000000d4_PCOUT<22>_UNCONNECTED , \NLW_blk000000d4_PCOUT<21>_UNCONNECTED ,
\NLW_blk000000d4_PCOUT<20>_UNCONNECTED , \NLW_blk000000d4_PCOUT<19>_UNCONNECTED , \NLW_blk000000d4_PCOUT<18>_UNCONNECTED ,
\NLW_blk000000d4_PCOUT<17>_UNCONNECTED , \NLW_blk000000d4_PCOUT<16>_UNCONNECTED , \NLW_blk000000d4_PCOUT<15>_UNCONNECTED ,
\NLW_blk000000d4_PCOUT<14>_UNCONNECTED , \NLW_blk000000d4_PCOUT<13>_UNCONNECTED , \NLW_blk000000d4_PCOUT<12>_UNCONNECTED ,
\NLW_blk000000d4_PCOUT<11>_UNCONNECTED , \NLW_blk000000d4_PCOUT<10>_UNCONNECTED , \NLW_blk000000d4_PCOUT<9>_UNCONNECTED ,
\NLW_blk000000d4_PCOUT<8>_UNCONNECTED , \NLW_blk000000d4_PCOUT<7>_UNCONNECTED , \NLW_blk000000d4_PCOUT<6>_UNCONNECTED ,
\NLW_blk000000d4_PCOUT<5>_UNCONNECTED , \NLW_blk000000d4_PCOUT<4>_UNCONNECTED , \NLW_blk000000d4_PCOUT<3>_UNCONNECTED ,
\NLW_blk000000d4_PCOUT<2>_UNCONNECTED , \NLW_blk000000d4_PCOUT<1>_UNCONNECTED , \NLW_blk000000d4_PCOUT<0>_UNCONNECTED }),
    .A({sig000003da, sig000003da, sig000003da, sig000003da, sig000003da, sig000003da, sig000003da, sig000003da, sig000003da, sig000003da, sig000003da
, sig000003da, sig000003da, sig000003da, sig000003da, sig000003da, sig000003da, sig000003db}),
    .M({\NLW_blk000000d4_M<35>_UNCONNECTED , \NLW_blk000000d4_M<34>_UNCONNECTED , \NLW_blk000000d4_M<33>_UNCONNECTED ,
\NLW_blk000000d4_M<32>_UNCONNECTED , \NLW_blk000000d4_M<31>_UNCONNECTED , \NLW_blk000000d4_M<30>_UNCONNECTED , \NLW_blk000000d4_M<29>_UNCONNECTED ,
\NLW_blk000000d4_M<28>_UNCONNECTED , \NLW_blk000000d4_M<27>_UNCONNECTED , \NLW_blk000000d4_M<26>_UNCONNECTED , \NLW_blk000000d4_M<25>_UNCONNECTED ,
\NLW_blk000000d4_M<24>_UNCONNECTED , \NLW_blk000000d4_M<23>_UNCONNECTED , \NLW_blk000000d4_M<22>_UNCONNECTED , \NLW_blk000000d4_M<21>_UNCONNECTED ,
\NLW_blk000000d4_M<20>_UNCONNECTED , \NLW_blk000000d4_M<19>_UNCONNECTED , \NLW_blk000000d4_M<18>_UNCONNECTED , \NLW_blk000000d4_M<17>_UNCONNECTED ,
\NLW_blk000000d4_M<16>_UNCONNECTED , \NLW_blk000000d4_M<15>_UNCONNECTED , \NLW_blk000000d4_M<14>_UNCONNECTED , \NLW_blk000000d4_M<13>_UNCONNECTED ,
\NLW_blk000000d4_M<12>_UNCONNECTED , \NLW_blk000000d4_M<11>_UNCONNECTED , \NLW_blk000000d4_M<10>_UNCONNECTED , \NLW_blk000000d4_M<9>_UNCONNECTED ,
\NLW_blk000000d4_M<8>_UNCONNECTED , \NLW_blk000000d4_M<7>_UNCONNECTED , \NLW_blk000000d4_M<6>_UNCONNECTED , \NLW_blk000000d4_M<5>_UNCONNECTED ,
\NLW_blk000000d4_M<4>_UNCONNECTED , \NLW_blk000000d4_M<3>_UNCONNECTED , \NLW_blk000000d4_M<2>_UNCONNECTED , \NLW_blk000000d4_M<1>_UNCONNECTED ,
\NLW_blk000000d4_M<0>_UNCONNECTED })
  );
  XORCY   blk000000d5 (
    .CI(sig00000413),
    .LI(sig00000412),
    .O(sig00000472)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk000000d6 (
    .I0(sig00000506),
    .I1(sig00000519),
    .O(sig00000412)
  );
  XORCY   blk000000d7 (
    .CI(sig00000415),
    .LI(sig00000414),
    .O(sig00000471)
  );
  MUXCY   blk000000d8 (
    .CI(sig00000415),
    .DI(sig00000506),
    .S(sig00000414),
    .O(sig00000413)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk000000d9 (
    .I0(sig00000506),
    .I1(sig00000519),
    .O(sig00000414)
  );
  XORCY   blk000000da (
    .CI(sig00000417),
    .LI(sig00000416),
    .O(sig00000470)
  );
  MUXCY   blk000000db (
    .CI(sig00000417),
    .DI(sig00000505),
    .S(sig00000416),
    .O(sig00000415)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk000000dc (
    .I0(sig00000505),
    .I1(sig00000518),
    .O(sig00000416)
  );
  XORCY   blk000000dd (
    .CI(sig00000419),
    .LI(sig00000418),
    .O(sig0000046f)
  );
  MUXCY   blk000000de (
    .CI(sig00000419),
    .DI(sig00000504),
    .S(sig00000418),
    .O(sig00000417)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk000000df (
    .I0(sig00000504),
    .I1(sig000003c9),
    .O(sig00000418)
  );
  XORCY   blk000000e0 (
    .CI(sig0000041b),
    .LI(sig0000041a),
    .O(sig0000046e)
  );
  MUXCY   blk000000e1 (
    .CI(sig0000041b),
    .DI(sig00000503),
    .S(sig0000041a),
    .O(sig00000419)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk000000e2 (
    .I0(sig00000503),
    .I1(sig000003ca),
    .O(sig0000041a)
  );
  XORCY   blk000000e3 (
    .CI(sig0000041d),
    .LI(sig0000041c),
    .O(sig0000046d)
  );
  MUXCY   blk000000e4 (
    .CI(sig0000041d),
    .DI(sig00000502),
    .S(sig0000041c),
    .O(sig0000041b)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk000000e5 (
    .I0(sig00000502),
    .I1(sig000003cb),
    .O(sig0000041c)
  );
  XORCY   blk000000e6 (
    .CI(sig0000041f),
    .LI(sig0000041e),
    .O(sig0000046c)
  );
  MUXCY   blk000000e7 (
    .CI(sig0000041f),
    .DI(sig00000501),
    .S(sig0000041e),
    .O(sig0000041d)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk000000e8 (
    .I0(sig00000501),
    .I1(sig000003cc),
    .O(sig0000041e)
  );
  XORCY   blk000000e9 (
    .CI(sig00000421),
    .LI(sig00000420),
    .O(sig0000046b)
  );
  MUXCY   blk000000ea (
    .CI(sig00000421),
    .DI(sig00000500),
    .S(sig00000420),
    .O(sig0000041f)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk000000eb (
    .I0(sig00000500),
    .I1(sig000003cd),
    .O(sig00000420)
  );
  XORCY   blk000000ec (
    .CI(sig00000423),
    .LI(sig00000422),
    .O(sig0000046a)
  );
  MUXCY   blk000000ed (
    .CI(sig00000423),
    .DI(sig000004ff),
    .S(sig00000422),
    .O(sig00000421)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk000000ee (
    .I0(sig000004ff),
    .I1(sig000003ce),
    .O(sig00000422)
  );
  XORCY   blk000000ef (
    .CI(sig00000425),
    .LI(sig00000424),
    .O(sig00000469)
  );
  MUXCY   blk000000f0 (
    .CI(sig00000425),
    .DI(sig000004fe),
    .S(sig00000424),
    .O(sig00000423)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk000000f1 (
    .I0(sig000004fe),
    .I1(sig000003cf),
    .O(sig00000424)
  );
  XORCY   blk000000f2 (
    .CI(sig00000427),
    .LI(sig00000426),
    .O(sig00000468)
  );
  MUXCY   blk000000f3 (
    .CI(sig00000427),
    .DI(sig000004fd),
    .S(sig00000426),
    .O(sig00000425)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk000000f4 (
    .I0(sig000004fd),
    .I1(sig000003d0),
    .O(sig00000426)
  );
  XORCY   blk000000f5 (
    .CI(sig00000429),
    .LI(sig00000428),
    .O(sig00000467)
  );
  MUXCY   blk000000f6 (
    .CI(sig00000429),
    .DI(sig000004fc),
    .S(sig00000428),
    .O(sig00000427)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk000000f7 (
    .I0(sig000004fc),
    .I1(sig000003d1),
    .O(sig00000428)
  );
  XORCY   blk000000f8 (
    .CI(sig0000042b),
    .LI(sig0000042a),
    .O(sig00000466)
  );
  MUXCY   blk000000f9 (
    .CI(sig0000042b),
    .DI(sig000004fb),
    .S(sig0000042a),
    .O(sig00000429)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk000000fa (
    .I0(sig000004fb),
    .I1(sig000003d2),
    .O(sig0000042a)
  );
  XORCY   blk000000fb (
    .CI(sig0000042d),
    .LI(sig0000042c),
    .O(sig00000465)
  );
  MUXCY   blk000000fc (
    .CI(sig0000042d),
    .DI(sig000004fa),
    .S(sig0000042c),
    .O(sig0000042b)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk000000fd (
    .I0(sig000004fa),
    .I1(sig000003d3),
    .O(sig0000042c)
  );
  XORCY   blk000000fe (
    .CI(sig0000042f),
    .LI(sig0000042e),
    .O(sig00000464)
  );
  MUXCY   blk000000ff (
    .CI(sig0000042f),
    .DI(sig000004f9),
    .S(sig0000042e),
    .O(sig0000042d)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000100 (
    .I0(sig000004f9),
    .I1(sig000003d4),
    .O(sig0000042e)
  );
  XORCY   blk00000101 (
    .CI(sig00000431),
    .LI(sig00000430),
    .O(sig00000463)
  );
  MUXCY   blk00000102 (
    .CI(sig00000431),
    .DI(sig000004f8),
    .S(sig00000430),
    .O(sig0000042f)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000103 (
    .I0(sig000004f8),
    .I1(sig000003d5),
    .O(sig00000430)
  );
  XORCY   blk00000104 (
    .CI(sig00000433),
    .LI(sig00000432),
    .O(sig00000462)
  );
  MUXCY   blk00000105 (
    .CI(sig00000433),
    .DI(sig000004f7),
    .S(sig00000432),
    .O(sig00000431)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000106 (
    .I0(sig000004f7),
    .I1(sig000003d6),
    .O(sig00000432)
  );
  XORCY   blk00000107 (
    .CI(sig00000435),
    .LI(sig00000434),
    .O(sig00000461)
  );
  MUXCY   blk00000108 (
    .CI(sig00000435),
    .DI(sig000004f6),
    .S(sig00000434),
    .O(sig00000433)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk00000109 (
    .I0(sig000004f6),
    .I1(sig000003d7),
    .O(sig00000434)
  );
  XORCY   blk0000010a (
    .CI(sig00000437),
    .LI(sig00000436),
    .O(sig00000460)
  );
  MUXCY   blk0000010b (
    .CI(sig00000437),
    .DI(sig000004f5),
    .S(sig00000436),
    .O(sig00000435)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk0000010c (
    .I0(sig000004f5),
    .I1(sig000003d8),
    .O(sig00000436)
  );
  MUXCY   blk0000010d (
    .CI(sig00000001),
    .DI(sig000004f4),
    .S(sig00000438),
    .O(sig00000437)
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  blk0000010e (
    .I0(sig000004f4),
    .I1(sig000003d9),
    .O(sig00000438)
  );
  XORCY   blk0000010f (
    .CI(sig0000043a),
    .LI(sig00000439),
    .O(sig00000486)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000110 (
    .I0(sig00000519),
    .I1(sig00000506),
    .O(sig00000439)
  );
  XORCY   blk00000111 (
    .CI(sig0000043c),
    .LI(sig0000043b),
    .O(sig00000485)
  );
  MUXCY   blk00000112 (
    .CI(sig0000043c),
    .DI(sig00000519),
    .S(sig0000043b),
    .O(sig0000043a)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000113 (
    .I0(sig00000519),
    .I1(sig00000506),
    .O(sig0000043b)
  );
  XORCY   blk00000114 (
    .CI(sig0000043e),
    .LI(sig0000043d),
    .O(sig00000484)
  );
  MUXCY   blk00000115 (
    .CI(sig0000043e),
    .DI(sig00000518),
    .S(sig0000043d),
    .O(sig0000043c)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000116 (
    .I0(sig00000518),
    .I1(sig00000505),
    .O(sig0000043d)
  );
  XORCY   blk00000117 (
    .CI(sig00000440),
    .LI(sig0000043f),
    .O(sig00000483)
  );
  MUXCY   blk00000118 (
    .CI(sig00000440),
    .DI(sig000003c9),
    .S(sig0000043f),
    .O(sig0000043e)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000119 (
    .I0(sig000003c9),
    .I1(sig00000504),
    .O(sig0000043f)
  );
  XORCY   blk0000011a (
    .CI(sig00000442),
    .LI(sig00000441),
    .O(sig00000482)
  );
  MUXCY   blk0000011b (
    .CI(sig00000442),
    .DI(sig000003ca),
    .S(sig00000441),
    .O(sig00000440)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk0000011c (
    .I0(sig000003ca),
    .I1(sig00000503),
    .O(sig00000441)
  );
  XORCY   blk0000011d (
    .CI(sig00000444),
    .LI(sig00000443),
    .O(sig00000481)
  );
  MUXCY   blk0000011e (
    .CI(sig00000444),
    .DI(sig000003cb),
    .S(sig00000443),
    .O(sig00000442)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk0000011f (
    .I0(sig000003cb),
    .I1(sig00000502),
    .O(sig00000443)
  );
  XORCY   blk00000120 (
    .CI(sig00000446),
    .LI(sig00000445),
    .O(sig00000480)
  );
  MUXCY   blk00000121 (
    .CI(sig00000446),
    .DI(sig000003cc),
    .S(sig00000445),
    .O(sig00000444)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000122 (
    .I0(sig000003cc),
    .I1(sig00000501),
    .O(sig00000445)
  );
  XORCY   blk00000123 (
    .CI(sig00000448),
    .LI(sig00000447),
    .O(sig0000047f)
  );
  MUXCY   blk00000124 (
    .CI(sig00000448),
    .DI(sig000003cd),
    .S(sig00000447),
    .O(sig00000446)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000125 (
    .I0(sig000003cd),
    .I1(sig00000500),
    .O(sig00000447)
  );
  XORCY   blk00000126 (
    .CI(sig0000044a),
    .LI(sig00000449),
    .O(sig0000047e)
  );
  MUXCY   blk00000127 (
    .CI(sig0000044a),
    .DI(sig000003ce),
    .S(sig00000449),
    .O(sig00000448)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000128 (
    .I0(sig000003ce),
    .I1(sig000004ff),
    .O(sig00000449)
  );
  XORCY   blk00000129 (
    .CI(sig0000044c),
    .LI(sig0000044b),
    .O(sig0000047d)
  );
  MUXCY   blk0000012a (
    .CI(sig0000044c),
    .DI(sig000003cf),
    .S(sig0000044b),
    .O(sig0000044a)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk0000012b (
    .I0(sig000003cf),
    .I1(sig000004fe),
    .O(sig0000044b)
  );
  XORCY   blk0000012c (
    .CI(sig0000044e),
    .LI(sig0000044d),
    .O(sig0000047c)
  );
  MUXCY   blk0000012d (
    .CI(sig0000044e),
    .DI(sig000003d0),
    .S(sig0000044d),
    .O(sig0000044c)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk0000012e (
    .I0(sig000003d0),
    .I1(sig000004fd),
    .O(sig0000044d)
  );
  XORCY   blk0000012f (
    .CI(sig00000450),
    .LI(sig0000044f),
    .O(sig0000047b)
  );
  MUXCY   blk00000130 (
    .CI(sig00000450),
    .DI(sig000003d1),
    .S(sig0000044f),
    .O(sig0000044e)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000131 (
    .I0(sig000003d1),
    .I1(sig000004fc),
    .O(sig0000044f)
  );
  XORCY   blk00000132 (
    .CI(sig00000452),
    .LI(sig00000451),
    .O(sig0000047a)
  );
  MUXCY   blk00000133 (
    .CI(sig00000452),
    .DI(sig000003d2),
    .S(sig00000451),
    .O(sig00000450)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000134 (
    .I0(sig000003d2),
    .I1(sig000004fb),
    .O(sig00000451)
  );
  XORCY   blk00000135 (
    .CI(sig00000454),
    .LI(sig00000453),
    .O(sig00000479)
  );
  MUXCY   blk00000136 (
    .CI(sig00000454),
    .DI(sig000003d3),
    .S(sig00000453),
    .O(sig00000452)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000137 (
    .I0(sig000003d3),
    .I1(sig000004fa),
    .O(sig00000453)
  );
  XORCY   blk00000138 (
    .CI(sig00000456),
    .LI(sig00000455),
    .O(sig00000478)
  );
  MUXCY   blk00000139 (
    .CI(sig00000456),
    .DI(sig000003d4),
    .S(sig00000455),
    .O(sig00000454)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk0000013a (
    .I0(sig000003d4),
    .I1(sig000004f9),
    .O(sig00000455)
  );
  XORCY   blk0000013b (
    .CI(sig00000458),
    .LI(sig00000457),
    .O(sig00000477)
  );
  MUXCY   blk0000013c (
    .CI(sig00000458),
    .DI(sig000003d5),
    .S(sig00000457),
    .O(sig00000456)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk0000013d (
    .I0(sig000003d5),
    .I1(sig000004f8),
    .O(sig00000457)
  );
  XORCY   blk0000013e (
    .CI(sig0000045a),
    .LI(sig00000459),
    .O(sig00000476)
  );
  MUXCY   blk0000013f (
    .CI(sig0000045a),
    .DI(sig000003d6),
    .S(sig00000459),
    .O(sig00000458)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000140 (
    .I0(sig000003d6),
    .I1(sig000004f7),
    .O(sig00000459)
  );
  XORCY   blk00000141 (
    .CI(sig0000045c),
    .LI(sig0000045b),
    .O(sig00000475)
  );
  MUXCY   blk00000142 (
    .CI(sig0000045c),
    .DI(sig000003d7),
    .S(sig0000045b),
    .O(sig0000045a)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000143 (
    .I0(sig000003d7),
    .I1(sig000004f6),
    .O(sig0000045b)
  );
  XORCY   blk00000144 (
    .CI(sig0000045e),
    .LI(sig0000045d),
    .O(sig00000474)
  );
  MUXCY   blk00000145 (
    .CI(sig0000045e),
    .DI(sig000003d8),
    .S(sig0000045d),
    .O(sig0000045c)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000146 (
    .I0(sig000003d8),
    .I1(sig000004f5),
    .O(sig0000045d)
  );
  XORCY   blk00000147 (
    .CI(sig00000002),
    .LI(sig0000045f),
    .O(sig00000473)
  );
  MUXCY   blk00000148 (
    .CI(sig00000002),
    .DI(sig000003d9),
    .S(sig0000045f),
    .O(sig0000045e)
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  blk00000149 (
    .I0(sig000003d9),
    .I1(sig000004f4),
    .O(sig0000045f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000014a (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000016),
    .Q(sig000003dc)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000014b (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000015),
    .Q(sig000003e5)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000014c (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000014),
    .Q(sig000003e6)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000014d (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000013),
    .Q(sig000003e7)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000014e (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000012),
    .Q(sig000003e8)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000014f (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000011),
    .Q(sig000003e9)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000150 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000010),
    .Q(sig000003ea)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000151 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000000f),
    .Q(sig000003eb)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000152 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000000e),
    .Q(sig000003ec)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000153 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000000d),
    .Q(sig000003ed)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000154 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000523),
    .Q(sig000004e9)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000155 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000522),
    .Q(sig000004e8)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000156 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000521),
    .Q(sig000004e7)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000157 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000520),
    .Q(sig000004e6)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000158 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000051f),
    .Q(sig000004e5)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000159 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000051e),
    .Q(sig000004e4)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000015a (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000051d),
    .Q(sig000004e3)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000015b (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000051c),
    .Q(sig000004e2)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000015c (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000051b),
    .Q(sig000004e1)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000015d (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000017),
    .Q(sig000004e0)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000015e (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000055),
    .Q(sig00000506)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000015f (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000054),
    .Q(sig00000505)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000160 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000053),
    .Q(sig00000504)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000161 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000052),
    .Q(sig00000503)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000162 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000051),
    .Q(sig00000502)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000163 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000050),
    .Q(sig00000501)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000164 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000004f),
    .Q(sig00000500)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000165 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000004e),
    .Q(sig000004ff)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000166 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000004d),
    .Q(sig000004fe)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000167 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000004c),
    .Q(sig000004fd)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000168 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000004b),
    .Q(sig000004fc)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000169 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000004a),
    .Q(sig000004fb)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000016a (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000049),
    .Q(sig000004fa)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000016b (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000048),
    .Q(sig000004f9)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000016c (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000047),
    .Q(sig000004f8)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000016d (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000046),
    .Q(sig000004f7)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000016e (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000045),
    .Q(sig000004f6)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000016f (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000044),
    .Q(sig000004f5)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000170 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000043),
    .Q(sig000004f4)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000171 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000068),
    .Q(sig00000519)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000172 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000067),
    .Q(sig00000518)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000173 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000066),
    .Q(sig000003c9)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000174 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000065),
    .Q(sig000003ca)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000175 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000064),
    .Q(sig000003cb)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000176 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000063),
    .Q(sig000003cc)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000177 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000062),
    .Q(sig000003cd)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000178 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000061),
    .Q(sig000003ce)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000179 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000060),
    .Q(sig000003cf)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000017a (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000005f),
    .Q(sig000003d0)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000017b (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000005e),
    .Q(sig000003d1)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000017c (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000005d),
    .Q(sig000003d2)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000017d (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000005c),
    .Q(sig000003d3)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000017e (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000005b),
    .Q(sig000003d4)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000017f (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000005a),
    .Q(sig000003d5)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000180 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000059),
    .Q(sig000003d6)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000181 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000058),
    .Q(sig000003d7)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000182 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000057),
    .Q(sig000003d8)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000183 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000056),
    .Q(sig000003d9)
  );
  DSP48A1 #(
    .A0REG ( 1 ),
    .A1REG ( 1 ),
    .B0REG ( 1 ),
    .B1REG ( 1 ),
    .CARRYINREG ( 0 ),
    .CARRYINSEL ( "OPMODE5" ),
    .CREG ( 1 ),
    .DREG ( 0 ),
    .MREG ( 1 ),
    .OPMODEREG ( 0 ),
    .PREG ( 1 ),
    .RSTTYPE ( "SYNC" ),
    .CARRYOUTREG ( 0 ))
  blk00000184 (
    .CECARRYIN(sig00000002),
    .RSTC(sig00000002),
    .RSTCARRYIN(sig00000002),
    .CED(sig00000002),
    .RSTD(sig00000002),
    .CEOPMODE(sig00000002),
    .CEC(sig00000001),
    .CARRYOUTF(NLW_blk00000184_CARRYOUTF_UNCONNECTED),
    .RSTOPMODE(sig00000002),
    .RSTM(sig00000002),
    .CLK(clk),
    .RSTB(sig00000002),
    .CEM(sig00000001),
    .CEB(sig00000001),
    .CARRYIN(sig00000002),
    .CEP(sig00000001),
    .CEA(sig00000001),
    .CARRYOUT(NLW_blk00000184_CARRYOUT_UNCONNECTED),
    .RSTA(sig00000002),
    .RSTP(sig00000002),
    .B({sig000005e1, sig000005e0, sig000005df, sig000005de, sig000005dd, sig000005dc, sig000005db, sig000005da, sig000005d9, sig000005d8, sig000005d7
, sig000005d6, sig000005d5, sig000005d4, sig000005d3, sig000005d2, sig000005d1, sig000005d0}),
    .BCOUT({\NLW_blk00000184_BCOUT<17>_UNCONNECTED , \NLW_blk00000184_BCOUT<16>_UNCONNECTED , \NLW_blk00000184_BCOUT<15>_UNCONNECTED ,
\NLW_blk00000184_BCOUT<14>_UNCONNECTED , \NLW_blk00000184_BCOUT<13>_UNCONNECTED , \NLW_blk00000184_BCOUT<12>_UNCONNECTED ,
\NLW_blk00000184_BCOUT<11>_UNCONNECTED , \NLW_blk00000184_BCOUT<10>_UNCONNECTED , \NLW_blk00000184_BCOUT<9>_UNCONNECTED ,
\NLW_blk00000184_BCOUT<8>_UNCONNECTED , \NLW_blk00000184_BCOUT<7>_UNCONNECTED , \NLW_blk00000184_BCOUT<6>_UNCONNECTED ,
\NLW_blk00000184_BCOUT<5>_UNCONNECTED , \NLW_blk00000184_BCOUT<4>_UNCONNECTED , \NLW_blk00000184_BCOUT<3>_UNCONNECTED ,
\NLW_blk00000184_BCOUT<2>_UNCONNECTED , \NLW_blk00000184_BCOUT<1>_UNCONNECTED , \NLW_blk00000184_BCOUT<0>_UNCONNECTED }),
    .PCIN({sig0000059f, sig0000059e, sig0000059d, sig0000059c, sig0000059b, sig0000059a, sig00000599, sig00000598, sig00000597, sig00000596,
sig00000595, sig00000594, sig00000593, sig00000592, sig00000591, sig00000590, sig0000058f, sig0000058e, sig0000058d, sig0000058c, sig0000058b,
sig0000058a, sig00000589, sig00000588, sig00000587, sig00000586, sig00000585, sig00000584, sig00000583, sig00000582, sig00000581, sig00000580,
sig0000057f, sig0000057e, sig0000057d, sig0000057c, sig0000057b, sig0000057a, sig00000579, sig00000578, sig00000577, sig00000576, sig00000575,
sig00000574, sig00000573, sig00000572, sig00000571, sig00000570}),
    .C({sig000005be, sig000005be, sig000005be, sig000005be, sig000005be, sig000005be, sig000005be, sig000005be, sig000005be, sig000005be, sig000005be
, sig000005be, sig000005be, sig000005be, sig000005be, sig000005be, sig000005be, sig000005be, sig000005bd, sig000005bc, sig000005bb, sig000005ba,
sig000005b9, sig000005b8, sig000005b7, sig000005b6, sig000005b5, sig000005b4, sig000005b3, sig000005b2, sig000005b1, sig000005b0, sig000005af,
sig000005ae, sig000005ad, sig000005ac, sig000005ab, sig000005aa, sig000005a9, sig000005a8, sig000005a7, sig000005a6, sig000005a5, sig000005a4,
sig000005a3, sig000005a2, sig000005a1, sig000005a0}),
    .P({\NLW_blk00000184_P<47>_UNCONNECTED , \NLW_blk00000184_P<46>_UNCONNECTED , \NLW_blk00000184_P<45>_UNCONNECTED ,
\NLW_blk00000184_P<44>_UNCONNECTED , \NLW_blk00000184_P<43>_UNCONNECTED , \NLW_blk00000184_P<42>_UNCONNECTED , \NLW_blk00000184_P<41>_UNCONNECTED ,
\NLW_blk00000184_P<40>_UNCONNECTED , \NLW_blk00000184_P<39>_UNCONNECTED , \NLW_blk00000184_P<38>_UNCONNECTED , \NLW_blk00000184_P<37>_UNCONNECTED ,
\NLW_blk00000184_P<36>_UNCONNECTED , sig00000547, sig00000546, sig00000545, sig00000544, sig00000543, sig00000542, sig00000541, sig00000540,
sig0000053f, sig0000053e, sig0000053d, sig0000053c, sig0000053b, sig0000053a, sig00000539, sig00000538, sig00000537, sig00000536, sig00000535,
sig00000534, sig00000533, sig00000532, sig00000531, sig00000530, sig0000052f, sig0000024c, sig0000024b, sig0000024a, sig00000249, sig00000248,
sig00000247, sig00000246, sig00000245, sig00000244, sig00000243, sig00000242}),
    .OPMODE({sig00000001, sig00000002, sig00000002, sig00000002, sig00000001, sig00000001, sig00000002, sig00000001}),
    .D({sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002
, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002}),
    .PCOUT({\NLW_blk00000184_PCOUT<47>_UNCONNECTED , \NLW_blk00000184_PCOUT<46>_UNCONNECTED , \NLW_blk00000184_PCOUT<45>_UNCONNECTED ,
\NLW_blk00000184_PCOUT<44>_UNCONNECTED , \NLW_blk00000184_PCOUT<43>_UNCONNECTED , \NLW_blk00000184_PCOUT<42>_UNCONNECTED ,
\NLW_blk00000184_PCOUT<41>_UNCONNECTED , \NLW_blk00000184_PCOUT<40>_UNCONNECTED , \NLW_blk00000184_PCOUT<39>_UNCONNECTED ,
\NLW_blk00000184_PCOUT<38>_UNCONNECTED , \NLW_blk00000184_PCOUT<37>_UNCONNECTED , \NLW_blk00000184_PCOUT<36>_UNCONNECTED ,
\NLW_blk00000184_PCOUT<35>_UNCONNECTED , \NLW_blk00000184_PCOUT<34>_UNCONNECTED , \NLW_blk00000184_PCOUT<33>_UNCONNECTED ,
\NLW_blk00000184_PCOUT<32>_UNCONNECTED , \NLW_blk00000184_PCOUT<31>_UNCONNECTED , \NLW_blk00000184_PCOUT<30>_UNCONNECTED ,
\NLW_blk00000184_PCOUT<29>_UNCONNECTED , \NLW_blk00000184_PCOUT<28>_UNCONNECTED , \NLW_blk00000184_PCOUT<27>_UNCONNECTED ,
\NLW_blk00000184_PCOUT<26>_UNCONNECTED , \NLW_blk00000184_PCOUT<25>_UNCONNECTED , \NLW_blk00000184_PCOUT<24>_UNCONNECTED ,
\NLW_blk00000184_PCOUT<23>_UNCONNECTED , \NLW_blk00000184_PCOUT<22>_UNCONNECTED , \NLW_blk00000184_PCOUT<21>_UNCONNECTED ,
\NLW_blk00000184_PCOUT<20>_UNCONNECTED , \NLW_blk00000184_PCOUT<19>_UNCONNECTED , \NLW_blk00000184_PCOUT<18>_UNCONNECTED ,
\NLW_blk00000184_PCOUT<17>_UNCONNECTED , \NLW_blk00000184_PCOUT<16>_UNCONNECTED , \NLW_blk00000184_PCOUT<15>_UNCONNECTED ,
\NLW_blk00000184_PCOUT<14>_UNCONNECTED , \NLW_blk00000184_PCOUT<13>_UNCONNECTED , \NLW_blk00000184_PCOUT<12>_UNCONNECTED ,
\NLW_blk00000184_PCOUT<11>_UNCONNECTED , \NLW_blk00000184_PCOUT<10>_UNCONNECTED , \NLW_blk00000184_PCOUT<9>_UNCONNECTED ,
\NLW_blk00000184_PCOUT<8>_UNCONNECTED , \NLW_blk00000184_PCOUT<7>_UNCONNECTED , \NLW_blk00000184_PCOUT<6>_UNCONNECTED ,
\NLW_blk00000184_PCOUT<5>_UNCONNECTED , \NLW_blk00000184_PCOUT<4>_UNCONNECTED , \NLW_blk00000184_PCOUT<3>_UNCONNECTED ,
\NLW_blk00000184_PCOUT<2>_UNCONNECTED , \NLW_blk00000184_PCOUT<1>_UNCONNECTED , \NLW_blk00000184_PCOUT<0>_UNCONNECTED }),
    .A({sig0000055d, sig0000055d, sig0000055d, sig0000055d, sig0000055d, sig0000055d, sig0000055d, sig0000055d, sig0000055d, sig0000055d, sig0000055d
, sig0000055d, sig0000055d, sig0000055d, sig0000055d, sig0000055d, sig0000055c, sig0000055b}),
    .M({\NLW_blk00000184_M<35>_UNCONNECTED , \NLW_blk00000184_M<34>_UNCONNECTED , \NLW_blk00000184_M<33>_UNCONNECTED ,
\NLW_blk00000184_M<32>_UNCONNECTED , \NLW_blk00000184_M<31>_UNCONNECTED , \NLW_blk00000184_M<30>_UNCONNECTED , \NLW_blk00000184_M<29>_UNCONNECTED ,
\NLW_blk00000184_M<28>_UNCONNECTED , \NLW_blk00000184_M<27>_UNCONNECTED , \NLW_blk00000184_M<26>_UNCONNECTED , \NLW_blk00000184_M<25>_UNCONNECTED ,
\NLW_blk00000184_M<24>_UNCONNECTED , \NLW_blk00000184_M<23>_UNCONNECTED , \NLW_blk00000184_M<22>_UNCONNECTED , \NLW_blk00000184_M<21>_UNCONNECTED ,
\NLW_blk00000184_M<20>_UNCONNECTED , \NLW_blk00000184_M<19>_UNCONNECTED , \NLW_blk00000184_M<18>_UNCONNECTED , \NLW_blk00000184_M<17>_UNCONNECTED ,
\NLW_blk00000184_M<16>_UNCONNECTED , \NLW_blk00000184_M<15>_UNCONNECTED , \NLW_blk00000184_M<14>_UNCONNECTED , \NLW_blk00000184_M<13>_UNCONNECTED ,
\NLW_blk00000184_M<12>_UNCONNECTED , \NLW_blk00000184_M<11>_UNCONNECTED , \NLW_blk00000184_M<10>_UNCONNECTED , \NLW_blk00000184_M<9>_UNCONNECTED ,
\NLW_blk00000184_M<8>_UNCONNECTED , \NLW_blk00000184_M<7>_UNCONNECTED , \NLW_blk00000184_M<6>_UNCONNECTED , \NLW_blk00000184_M<5>_UNCONNECTED ,
\NLW_blk00000184_M<4>_UNCONNECTED , \NLW_blk00000184_M<3>_UNCONNECTED , \NLW_blk00000184_M<2>_UNCONNECTED , \NLW_blk00000184_M<1>_UNCONNECTED ,
\NLW_blk00000184_M<0>_UNCONNECTED })
  );
  DSP48A1 #(
    .A0REG ( 1 ),
    .A1REG ( 1 ),
    .B0REG ( 1 ),
    .B1REG ( 1 ),
    .CARRYINREG ( 0 ),
    .CARRYINSEL ( "OPMODE5" ),
    .CREG ( 1 ),
    .DREG ( 0 ),
    .MREG ( 1 ),
    .OPMODEREG ( 0 ),
    .PREG ( 1 ),
    .RSTTYPE ( "SYNC" ),
    .CARRYOUTREG ( 0 ))
  blk00000185 (
    .CECARRYIN(sig00000002),
    .RSTC(sig00000002),
    .RSTCARRYIN(sig00000002),
    .CED(sig00000002),
    .RSTD(sig00000002),
    .CEOPMODE(sig00000002),
    .CEC(sig00000001),
    .CARRYOUTF(NLW_blk00000185_CARRYOUTF_UNCONNECTED),
    .RSTOPMODE(sig00000002),
    .RSTM(sig00000002),
    .CLK(clk),
    .RSTB(sig00000002),
    .CEM(sig00000001),
    .CEB(sig00000001),
    .CARRYIN(sig00000002),
    .CEP(sig00000001),
    .CEA(sig00000001),
    .CARRYOUT(NLW_blk00000185_CARRYOUT_UNCONNECTED),
    .RSTA(sig00000002),
    .RSTP(sig00000002),
    .B({sig000004cb, sig000004cb, sig000004cb, sig000004cb, sig000004cb, sig000004cb, sig000004cb, sig000004cb, sig000004cb, sig000004ca, sig000004c9
, sig000004c8, sig000004c7, sig000004c6, sig000004c5, sig000004c4, sig000004c3, sig000004c2}),
    .BCOUT({sig000005e1, sig000005e0, sig000005df, sig000005de, sig000005dd, sig000005dc, sig000005db, sig000005da, sig000005d9, sig000005d8,
sig000005d7, sig000005d6, sig000005d5, sig000005d4, sig000005d3, sig000005d2, sig000005d1, sig000005d0}),
    .PCIN({sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002,
sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002,
sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002,
sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002,
sig00000002, sig00000002, sig00000002, sig00000002, sig00000002}),
    .C({sig00000405, sig00000405, sig00000405, sig00000405, sig00000405, sig00000405, sig00000405, sig00000405, sig00000405, sig00000405, sig00000405
, sig00000405, sig00000405, sig00000405, sig00000405, sig00000405, sig00000405, sig00000405, sig00000405, sig00000406, sig00000407, sig00000408,
sig00000409, sig0000040a, sig0000040b, sig0000040c, sig0000040d, sig0000040e, sig0000040f, sig00000410, sig00000411, sig000004b4, sig000004b3,
sig000004b2, sig000004b1, sig000004b0, sig000004af, sig000004ae, sig000004ad, sig000004ac, sig000004ab, sig000004aa, sig000004a9, sig000004a8,
sig000004a7, sig000004a6, sig000004a5, sig000004a4}),
    .P({sig000005be, sig000005bd, sig000005bc, sig000005bb, sig000005ba, sig000005b9, sig000005b8, sig000005b7, sig000005b6, sig000005b5, sig000005b4
, sig000005b3, sig000005b2, sig000005b1, sig000005b0, sig000005af, sig000005ae, sig000005ad, sig000005ac, sig000005ab, sig000005aa, sig000005a9,
sig000005a8, sig000005a7, sig000005a6, sig000005a5, sig000005a4, sig000005a3, sig000005a2, sig000005a1, sig000005a0, sig000005cf, sig000005ce,
sig000005cd, sig000005cc, sig000005cb, sig000005ca, sig000005c9, sig000005c8, sig000005c7, sig000005c6, sig000005c5, sig000005c4, sig000005c3,
sig000005c2, sig000005c1, sig000005c0, sig000005bf}),
    .OPMODE({sig00000001, sig00000002, sig00000002, sig00000002, sig00000001, sig00000001, sig00000002, sig00000001}),
    .D({sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002
, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002}),
    .PCOUT({sig0000059f, sig0000059e, sig0000059d, sig0000059c, sig0000059b, sig0000059a, sig00000599, sig00000598, sig00000597, sig00000596,
sig00000595, sig00000594, sig00000593, sig00000592, sig00000591, sig00000590, sig0000058f, sig0000058e, sig0000058d, sig0000058c, sig0000058b,
sig0000058a, sig00000589, sig00000588, sig00000587, sig00000586, sig00000585, sig00000584, sig00000583, sig00000582, sig00000581, sig00000580,
sig0000057f, sig0000057e, sig0000057d, sig0000057c, sig0000057b, sig0000057a, sig00000579, sig00000578, sig00000577, sig00000576, sig00000575,
sig00000574, sig00000573, sig00000572, sig00000571, sig00000570}),
    .A({sig00000002, sig000004dc, sig000004db, sig000004da, sig000004d9, sig000004d8, sig000004d7, sig000004d6, sig000004d5, sig000004d4, sig000004d3
, sig000004d2, sig000004d1, sig000004d0, sig000004cf, sig000004ce, sig000004cd, sig0000031c}),
    .M({\NLW_blk00000185_M<35>_UNCONNECTED , \NLW_blk00000185_M<34>_UNCONNECTED , \NLW_blk00000185_M<33>_UNCONNECTED ,
\NLW_blk00000185_M<32>_UNCONNECTED , \NLW_blk00000185_M<31>_UNCONNECTED , \NLW_blk00000185_M<30>_UNCONNECTED , \NLW_blk00000185_M<29>_UNCONNECTED ,
\NLW_blk00000185_M<28>_UNCONNECTED , \NLW_blk00000185_M<27>_UNCONNECTED , \NLW_blk00000185_M<26>_UNCONNECTED , \NLW_blk00000185_M<25>_UNCONNECTED ,
\NLW_blk00000185_M<24>_UNCONNECTED , \NLW_blk00000185_M<23>_UNCONNECTED , \NLW_blk00000185_M<22>_UNCONNECTED , \NLW_blk00000185_M<21>_UNCONNECTED ,
\NLW_blk00000185_M<20>_UNCONNECTED , \NLW_blk00000185_M<19>_UNCONNECTED , \NLW_blk00000185_M<18>_UNCONNECTED , \NLW_blk00000185_M<17>_UNCONNECTED ,
\NLW_blk00000185_M<16>_UNCONNECTED , \NLW_blk00000185_M<15>_UNCONNECTED , \NLW_blk00000185_M<14>_UNCONNECTED , \NLW_blk00000185_M<13>_UNCONNECTED ,
\NLW_blk00000185_M<12>_UNCONNECTED , \NLW_blk00000185_M<11>_UNCONNECTED , \NLW_blk00000185_M<10>_UNCONNECTED , \NLW_blk00000185_M<9>_UNCONNECTED ,
\NLW_blk00000185_M<8>_UNCONNECTED , \NLW_blk00000185_M<7>_UNCONNECTED , \NLW_blk00000185_M<6>_UNCONNECTED , \NLW_blk00000185_M<5>_UNCONNECTED ,
\NLW_blk00000185_M<4>_UNCONNECTED , \NLW_blk00000185_M<3>_UNCONNECTED , \NLW_blk00000185_M<2>_UNCONNECTED , \NLW_blk00000185_M<1>_UNCONNECTED ,
\NLW_blk00000185_M<0>_UNCONNECTED })
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000037a (
    .C(clk),
    .CE(sig00000001),
    .D(sig000005e8),
    .Q(sig00000114)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000037b (
    .C(clk),
    .CE(sig00000001),
    .D(sig000005e9),
    .Q(sig00000115)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000037c (
    .C(clk),
    .CE(sig00000001),
    .D(sig000005ea),
    .Q(sig00000116)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000037d (
    .C(clk),
    .CE(sig00000001),
    .D(sig000005eb),
    .Q(sig00000117)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000037e (
    .C(clk),
    .CE(sig00000001),
    .D(sig000005ec),
    .Q(sig00000118)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000037f (
    .C(clk),
    .CE(sig00000001),
    .D(sig000005ed),
    .Q(sig00000119)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000380 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000005ee),
    .Q(sig0000011a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000381 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000005ef),
    .Q(sig0000011b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000382 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000005f0),
    .Q(sig0000011c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000383 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000005f1),
    .Q(sig0000011d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000384 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000005f2),
    .Q(sig0000011e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000385 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000005f3),
    .Q(sig0000011f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000386 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000005f4),
    .Q(sig00000120)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000387 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000005f5),
    .Q(sig00000121)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000388 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000005f6),
    .Q(sig00000122)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000389 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000005f7),
    .Q(sig00000123)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000038a (
    .C(clk),
    .CE(sig00000001),
    .D(sig000005f8),
    .Q(sig00000124)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000038b (
    .C(clk),
    .CE(sig00000001),
    .D(sig000005f9),
    .Q(sig00000125)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000038c (
    .C(clk),
    .CE(sig00000001),
    .D(sig000005fa),
    .Q(sig00000126)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000038d (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000060e),
    .Q(sig000005e5)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000038e (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000060f),
    .Q(sig000005e6)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000038f (
    .C(clk),
    .CE(sig00000001),
    .D(sig000005e2),
    .Q(sig000005e4)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000390 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000001c9),
    .Q(sig000005e3)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000391 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000001ca),
    .Q(sig000005e7)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000392 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000616),
    .Q(sig00000101)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000393 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000617),
    .Q(sig00000102)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000394 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000618),
    .Q(sig00000103)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000395 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000619),
    .Q(sig00000104)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000396 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000061a),
    .Q(sig00000105)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000397 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000061b),
    .Q(sig00000106)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000398 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000061c),
    .Q(sig00000107)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000399 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000061d),
    .Q(sig00000108)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000039a (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000061e),
    .Q(sig00000109)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000039b (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000061f),
    .Q(sig0000010a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000039c (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000620),
    .Q(sig0000010b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000039d (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000621),
    .Q(sig0000010c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000039e (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000622),
    .Q(sig0000010d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000039f (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000623),
    .Q(sig0000010e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003a0 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000624),
    .Q(sig0000010f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003a1 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000625),
    .Q(sig00000110)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003a2 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000626),
    .Q(sig00000111)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003a3 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000627),
    .Q(sig00000112)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003a4 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000628),
    .Q(sig00000113)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003a5 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000063c),
    .Q(sig00000613)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003a6 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000063d),
    .Q(sig00000614)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003a7 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000610),
    .Q(sig00000612)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003a8 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000001df),
    .Q(sig00000611)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003a9 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000001e0),
    .Q(sig00000615)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003aa (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000644),
    .Q(sig0000013a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003ab (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000645),
    .Q(sig0000013b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003ac (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000646),
    .Q(sig0000013c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003ad (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000647),
    .Q(sig0000013d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003ae (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000648),
    .Q(sig0000013e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003af (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000649),
    .Q(sig0000013f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003b0 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000064a),
    .Q(sig00000140)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003b1 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000064b),
    .Q(sig00000141)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003b2 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000064c),
    .Q(sig00000142)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003b3 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000064d),
    .Q(sig00000143)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003b4 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000064e),
    .Q(sig00000144)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003b5 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000064f),
    .Q(sig00000145)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003b6 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000650),
    .Q(sig00000146)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003b7 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000651),
    .Q(sig00000147)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003b8 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000652),
    .Q(sig00000148)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003b9 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000653),
    .Q(sig00000149)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003ba (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000654),
    .Q(sig0000014a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003bb (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000655),
    .Q(sig0000014b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003bc (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000656),
    .Q(sig0000014c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003bd (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000066a),
    .Q(sig00000641)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003be (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000066b),
    .Q(sig00000642)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003bf (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000063e),
    .Q(sig00000640)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003c0 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000001f5),
    .Q(sig0000063f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003c1 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000001f6),
    .Q(sig00000643)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003c2 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000672),
    .Q(sig00000127)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003c3 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000673),
    .Q(sig00000128)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003c4 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000674),
    .Q(sig00000129)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003c5 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000675),
    .Q(sig0000012a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003c6 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000676),
    .Q(sig0000012b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003c7 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000677),
    .Q(sig0000012c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003c8 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000678),
    .Q(sig0000012d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003c9 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000679),
    .Q(sig0000012e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003ca (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000067a),
    .Q(sig0000012f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003cb (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000067b),
    .Q(sig00000130)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003cc (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000067c),
    .Q(sig00000131)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003cd (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000067d),
    .Q(sig00000132)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003ce (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000067e),
    .Q(sig00000133)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003cf (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000067f),
    .Q(sig00000134)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003d0 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000680),
    .Q(sig00000135)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003d1 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000681),
    .Q(sig00000136)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003d2 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000682),
    .Q(sig00000137)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003d3 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000683),
    .Q(sig00000138)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003d4 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000684),
    .Q(sig00000139)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003d5 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000698),
    .Q(sig0000066f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003d6 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000699),
    .Q(sig00000670)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003d7 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000066c),
    .Q(sig0000066e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003d8 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000020b),
    .Q(sig0000066d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk000003d9 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000020c),
    .Q(sig00000671)
  );
  XORCY   blk000003da (
    .CI(sig0000069a),
    .LI(sig00000002),
    .O(sig00000698)
  );
  MUXCY   blk000003db (
    .CI(sig0000069d),
    .DI(sig00000002),
    .S(sig0000069e),
    .O(sig0000069a)
  );
  MUXCY   blk000003dc (
    .CI(sig00000001),
    .DI(sig00000002),
    .S(sig0000069f),
    .O(sig0000069b)
  );
  MUXCY   blk000003dd (
    .CI(sig0000069b),
    .DI(sig00000002),
    .S(sig000006a0),
    .O(sig0000069c)
  );
  MUXCY   blk000003de (
    .CI(sig0000069c),
    .DI(sig00000002),
    .S(sig000006a1),
    .O(sig0000069d)
  );
  LUT6 #(
    .INIT ( 64'h8000000000000000 ))
  blk000003df (
    .I0(sig000006a2),
    .I1(sig00000001),
    .I2(sig00000001),
    .I3(sig00000001),
    .I4(sig00000001),
    .I5(sig00000001),
    .O(sig0000069e)
  );
  LUT6 #(
    .INIT ( 64'h8000000000000000 ))
  blk000003e0 (
    .I0(sig0000020c),
    .I1(sig0000020d),
    .I2(sig0000020e),
    .I3(sig0000020f),
    .I4(sig00000210),
    .I5(sig00000211),
    .O(sig0000069f)
  );
  LUT6 #(
    .INIT ( 64'h8000000000000000 ))
  blk000003e1 (
    .I0(sig00000212),
    .I1(sig00000213),
    .I2(sig00000214),
    .I3(sig00000215),
    .I4(sig00000216),
    .I5(sig00000217),
    .O(sig000006a0)
  );
  LUT6 #(
    .INIT ( 64'h8000000000000000 ))
  blk000003e2 (
    .I0(sig00000218),
    .I1(sig00000219),
    .I2(sig0000021a),
    .I3(sig0000021b),
    .I4(sig0000021c),
    .I5(sig0000021d),
    .O(sig000006a1)
  );
  XORCY   blk000003e3 (
    .CI(sig000006a3),
    .LI(sig00000002),
    .O(sig0000066a)
  );
  MUXCY   blk000003e4 (
    .CI(sig000006a6),
    .DI(sig00000002),
    .S(sig000006a7),
    .O(sig000006a3)
  );
  MUXCY   blk000003e5 (
    .CI(sig00000001),
    .DI(sig00000002),
    .S(sig000006a8),
    .O(sig000006a4)
  );
  MUXCY   blk000003e6 (
    .CI(sig000006a4),
    .DI(sig00000002),
    .S(sig000006a9),
    .O(sig000006a5)
  );
  MUXCY   blk000003e7 (
    .CI(sig000006a5),
    .DI(sig00000002),
    .S(sig000006aa),
    .O(sig000006a6)
  );
  LUT6 #(
    .INIT ( 64'h8000000000000000 ))
  blk000003e8 (
    .I0(sig000006ab),
    .I1(sig00000001),
    .I2(sig00000001),
    .I3(sig00000001),
    .I4(sig00000001),
    .I5(sig00000001),
    .O(sig000006a7)
  );
  LUT6 #(
    .INIT ( 64'h8000000000000000 ))
  blk000003e9 (
    .I0(sig000001f6),
    .I1(sig000001f7),
    .I2(sig000001f8),
    .I3(sig000001f9),
    .I4(sig000001fa),
    .I5(sig000001fb),
    .O(sig000006a8)
  );
  LUT6 #(
    .INIT ( 64'h8000000000000000 ))
  blk000003ea (
    .I0(sig000001fc),
    .I1(sig000001fd),
    .I2(sig000001fe),
    .I3(sig000001ff),
    .I4(sig00000200),
    .I5(sig00000201),
    .O(sig000006a9)
  );
  LUT6 #(
    .INIT ( 64'h8000000000000000 ))
  blk000003eb (
    .I0(sig00000202),
    .I1(sig00000203),
    .I2(sig00000204),
    .I3(sig00000205),
    .I4(sig00000206),
    .I5(sig00000207),
    .O(sig000006aa)
  );
  XORCY   blk000003ec (
    .CI(sig000006ac),
    .LI(sig00000002),
    .O(sig0000063c)
  );
  MUXCY   blk000003ed (
    .CI(sig000006af),
    .DI(sig00000002),
    .S(sig000006b0),
    .O(sig000006ac)
  );
  MUXCY   blk000003ee (
    .CI(sig00000001),
    .DI(sig00000002),
    .S(sig000006b1),
    .O(sig000006ad)
  );
  MUXCY   blk000003ef (
    .CI(sig000006ad),
    .DI(sig00000002),
    .S(sig000006b2),
    .O(sig000006ae)
  );
  MUXCY   blk000003f0 (
    .CI(sig000006ae),
    .DI(sig00000002),
    .S(sig000006b3),
    .O(sig000006af)
  );
  LUT6 #(
    .INIT ( 64'h8000000000000000 ))
  blk000003f1 (
    .I0(sig000006b4),
    .I1(sig00000001),
    .I2(sig00000001),
    .I3(sig00000001),
    .I4(sig00000001),
    .I5(sig00000001),
    .O(sig000006b0)
  );
  LUT6 #(
    .INIT ( 64'h8000000000000000 ))
  blk000003f2 (
    .I0(sig000001e0),
    .I1(sig000001e1),
    .I2(sig000001e2),
    .I3(sig000001e3),
    .I4(sig000001e4),
    .I5(sig000001e5),
    .O(sig000006b1)
  );
  LUT6 #(
    .INIT ( 64'h8000000000000000 ))
  blk000003f3 (
    .I0(sig000001e6),
    .I1(sig000001e7),
    .I2(sig000001e8),
    .I3(sig000001e9),
    .I4(sig000001ea),
    .I5(sig000001eb),
    .O(sig000006b2)
  );
  LUT6 #(
    .INIT ( 64'h8000000000000000 ))
  blk000003f4 (
    .I0(sig000001ec),
    .I1(sig000001ed),
    .I2(sig000001ee),
    .I3(sig000001ef),
    .I4(sig000001f0),
    .I5(sig000001f1),
    .O(sig000006b3)
  );
  XORCY   blk000003f5 (
    .CI(sig000006b5),
    .LI(sig00000002),
    .O(sig0000060e)
  );
  MUXCY   blk000003f6 (
    .CI(sig000006b8),
    .DI(sig00000002),
    .S(sig000006b9),
    .O(sig000006b5)
  );
  MUXCY   blk000003f7 (
    .CI(sig00000001),
    .DI(sig00000002),
    .S(sig000006ba),
    .O(sig000006b6)
  );
  MUXCY   blk000003f8 (
    .CI(sig000006b6),
    .DI(sig00000002),
    .S(sig000006bb),
    .O(sig000006b7)
  );
  MUXCY   blk000003f9 (
    .CI(sig000006b7),
    .DI(sig00000002),
    .S(sig000006bc),
    .O(sig000006b8)
  );
  LUT6 #(
    .INIT ( 64'h8000000000000000 ))
  blk000003fa (
    .I0(sig000006bd),
    .I1(sig00000001),
    .I2(sig00000001),
    .I3(sig00000001),
    .I4(sig00000001),
    .I5(sig00000001),
    .O(sig000006b9)
  );
  LUT6 #(
    .INIT ( 64'h8000000000000000 ))
  blk000003fb (
    .I0(sig000001ca),
    .I1(sig000001cb),
    .I2(sig000001cc),
    .I3(sig000001cd),
    .I4(sig000001ce),
    .I5(sig000001cf),
    .O(sig000006ba)
  );
  LUT6 #(
    .INIT ( 64'h8000000000000000 ))
  blk000003fc (
    .I0(sig000001d0),
    .I1(sig000001d1),
    .I2(sig000001d2),
    .I3(sig000001d3),
    .I4(sig000001d4),
    .I5(sig000001d5),
    .O(sig000006bb)
  );
  LUT6 #(
    .INIT ( 64'h8000000000000000 ))
  blk000003fd (
    .I0(sig000001d6),
    .I1(sig000001d7),
    .I2(sig000001d8),
    .I3(sig000001d9),
    .I4(sig000001da),
    .I5(sig000001db),
    .O(sig000006bc)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000003fe (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig0000021e),
    .Q(sig000006be)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000003ff (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig0000021d),
    .Q(sig000006bf)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000400 (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig0000021c),
    .Q(sig000006c0)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000401 (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig0000021b),
    .Q(sig000006c1)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000402 (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig0000021a),
    .Q(sig000006c2)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000403 (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig00000219),
    .Q(sig000006c3)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000404 (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig00000218),
    .Q(sig000006c4)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000405 (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig00000217),
    .Q(sig000006c5)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000406 (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig00000216),
    .Q(sig000006c6)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000407 (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig00000215),
    .Q(sig000006c7)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000408 (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig00000214),
    .Q(sig000006c8)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000409 (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig00000213),
    .Q(sig000006c9)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000040a (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig00000212),
    .Q(sig000006ca)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000040b (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig00000211),
    .Q(sig000006cb)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000040c (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig00000210),
    .Q(sig000006cc)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000040d (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig0000020f),
    .Q(sig000006cd)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000040e (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig0000020e),
    .Q(sig000006ce)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000040f (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig0000020d),
    .Q(sig000006cf)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000410 (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig0000020c),
    .Q(sig000006d0)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000411 (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig0000020b),
    .Q(sig000006d1)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000412 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000006be),
    .R(sig00000002),
    .Q(sig00000697)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000413 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000006bf),
    .R(sig00000002),
    .Q(sig00000696)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000414 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000006c0),
    .R(sig00000002),
    .Q(sig00000695)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000415 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000006c1),
    .R(sig00000002),
    .Q(sig00000694)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000416 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000006c2),
    .R(sig00000002),
    .Q(sig00000693)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000417 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000006c3),
    .R(sig00000002),
    .Q(sig00000692)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000418 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000006c4),
    .R(sig00000002),
    .Q(sig00000691)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000419 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000006c5),
    .R(sig00000002),
    .Q(sig00000690)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000041a (
    .C(clk),
    .CE(sig00000001),
    .D(sig000006c6),
    .R(sig00000002),
    .Q(sig0000068f)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000041b (
    .C(clk),
    .CE(sig00000001),
    .D(sig000006c7),
    .R(sig00000002),
    .Q(sig0000068e)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000041c (
    .C(clk),
    .CE(sig00000001),
    .D(sig000006c8),
    .R(sig00000002),
    .Q(sig0000068d)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000041d (
    .C(clk),
    .CE(sig00000001),
    .D(sig000006c9),
    .R(sig00000002),
    .Q(sig0000068c)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000041e (
    .C(clk),
    .CE(sig00000001),
    .D(sig000006ca),
    .R(sig00000002),
    .Q(sig0000068b)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000041f (
    .C(clk),
    .CE(sig00000001),
    .D(sig000006cb),
    .R(sig00000002),
    .Q(sig0000068a)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000420 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000006cc),
    .R(sig00000002),
    .Q(sig00000689)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000421 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000006cd),
    .R(sig00000002),
    .Q(sig00000688)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000422 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000006ce),
    .R(sig00000002),
    .Q(sig00000687)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000423 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000006cf),
    .R(sig00000002),
    .Q(sig00000686)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000424 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000006d0),
    .R(sig00000002),
    .Q(sig00000685)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000425 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000006d1),
    .R(sig00000002),
    .Q(NLW_blk00000425_Q_UNCONNECTED)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000426 (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig00000208),
    .Q(sig000006d2)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000427 (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig00000207),
    .Q(sig000006d3)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000428 (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig00000206),
    .Q(sig000006d4)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000429 (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig00000205),
    .Q(sig000006d5)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000042a (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig00000204),
    .Q(sig000006d6)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000042b (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig00000203),
    .Q(sig000006d7)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000042c (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig00000202),
    .Q(sig000006d8)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000042d (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig00000201),
    .Q(sig000006d9)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000042e (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig00000200),
    .Q(sig000006da)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000042f (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000001ff),
    .Q(sig000006db)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000430 (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000001fe),
    .Q(sig000006dc)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000431 (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000001fd),
    .Q(sig000006dd)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000432 (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000001fc),
    .Q(sig000006de)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000433 (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000001fb),
    .Q(sig000006df)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000434 (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000001fa),
    .Q(sig000006e0)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000435 (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000001f9),
    .Q(sig000006e1)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000436 (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000001f8),
    .Q(sig000006e2)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000437 (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000001f7),
    .Q(sig000006e3)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000438 (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000001f6),
    .Q(sig000006e4)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000439 (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000001f5),
    .Q(sig000006e5)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000043a (
    .C(clk),
    .CE(sig00000001),
    .D(sig000006d2),
    .R(sig00000002),
    .Q(sig00000669)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000043b (
    .C(clk),
    .CE(sig00000001),
    .D(sig000006d3),
    .R(sig00000002),
    .Q(sig00000668)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000043c (
    .C(clk),
    .CE(sig00000001),
    .D(sig000006d4),
    .R(sig00000002),
    .Q(sig00000667)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000043d (
    .C(clk),
    .CE(sig00000001),
    .D(sig000006d5),
    .R(sig00000002),
    .Q(sig00000666)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000043e (
    .C(clk),
    .CE(sig00000001),
    .D(sig000006d6),
    .R(sig00000002),
    .Q(sig00000665)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000043f (
    .C(clk),
    .CE(sig00000001),
    .D(sig000006d7),
    .R(sig00000002),
    .Q(sig00000664)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000440 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000006d8),
    .R(sig00000002),
    .Q(sig00000663)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000441 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000006d9),
    .R(sig00000002),
    .Q(sig00000662)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000442 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000006da),
    .R(sig00000002),
    .Q(sig00000661)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000443 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000006db),
    .R(sig00000002),
    .Q(sig00000660)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000444 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000006dc),
    .R(sig00000002),
    .Q(sig0000065f)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000445 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000006dd),
    .R(sig00000002),
    .Q(sig0000065e)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000446 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000006de),
    .R(sig00000002),
    .Q(sig0000065d)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000447 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000006df),
    .R(sig00000002),
    .Q(sig0000065c)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000448 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000006e0),
    .R(sig00000002),
    .Q(sig0000065b)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000449 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000006e1),
    .R(sig00000002),
    .Q(sig0000065a)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000044a (
    .C(clk),
    .CE(sig00000001),
    .D(sig000006e2),
    .R(sig00000002),
    .Q(sig00000659)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000044b (
    .C(clk),
    .CE(sig00000001),
    .D(sig000006e3),
    .R(sig00000002),
    .Q(sig00000658)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000044c (
    .C(clk),
    .CE(sig00000001),
    .D(sig000006e4),
    .R(sig00000002),
    .Q(sig00000657)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000044d (
    .C(clk),
    .CE(sig00000001),
    .D(sig000006e5),
    .R(sig00000002),
    .Q(NLW_blk0000044d_Q_UNCONNECTED)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000044e (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000001f2),
    .Q(sig000006e6)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000044f (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000001f1),
    .Q(sig000006e7)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000450 (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000001f0),
    .Q(sig000006e8)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000451 (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000001ef),
    .Q(sig000006e9)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000452 (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000001ee),
    .Q(sig000006ea)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000453 (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000001ed),
    .Q(sig000006eb)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000454 (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000001ec),
    .Q(sig000006ec)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000455 (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000001eb),
    .Q(sig000006ed)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000456 (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000001ea),
    .Q(sig000006ee)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000457 (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000001e9),
    .Q(sig000006ef)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000458 (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000001e8),
    .Q(sig000006f0)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000459 (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000001e7),
    .Q(sig000006f1)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000045a (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000001e6),
    .Q(sig000006f2)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000045b (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000001e5),
    .Q(sig000006f3)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000045c (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000001e4),
    .Q(sig000006f4)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000045d (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000001e3),
    .Q(sig000006f5)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000045e (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000001e2),
    .Q(sig000006f6)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000045f (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000001e1),
    .Q(sig000006f7)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000460 (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000001e0),
    .Q(sig000006f8)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000461 (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000001df),
    .Q(sig000006f9)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000462 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000006e6),
    .R(sig00000002),
    .Q(sig0000063b)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000463 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000006e7),
    .R(sig00000002),
    .Q(sig0000063a)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000464 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000006e8),
    .R(sig00000002),
    .Q(sig00000639)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000465 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000006e9),
    .R(sig00000002),
    .Q(sig00000638)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000466 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000006ea),
    .R(sig00000002),
    .Q(sig00000637)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000467 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000006eb),
    .R(sig00000002),
    .Q(sig00000636)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000468 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000006ec),
    .R(sig00000002),
    .Q(sig00000635)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000469 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000006ed),
    .R(sig00000002),
    .Q(sig00000634)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000046a (
    .C(clk),
    .CE(sig00000001),
    .D(sig000006ee),
    .R(sig00000002),
    .Q(sig00000633)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000046b (
    .C(clk),
    .CE(sig00000001),
    .D(sig000006ef),
    .R(sig00000002),
    .Q(sig00000632)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000046c (
    .C(clk),
    .CE(sig00000001),
    .D(sig000006f0),
    .R(sig00000002),
    .Q(sig00000631)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000046d (
    .C(clk),
    .CE(sig00000001),
    .D(sig000006f1),
    .R(sig00000002),
    .Q(sig00000630)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000046e (
    .C(clk),
    .CE(sig00000001),
    .D(sig000006f2),
    .R(sig00000002),
    .Q(sig0000062f)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000046f (
    .C(clk),
    .CE(sig00000001),
    .D(sig000006f3),
    .R(sig00000002),
    .Q(sig0000062e)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000470 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000006f4),
    .R(sig00000002),
    .Q(sig0000062d)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000471 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000006f5),
    .R(sig00000002),
    .Q(sig0000062c)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000472 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000006f6),
    .R(sig00000002),
    .Q(sig0000062b)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000473 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000006f7),
    .R(sig00000002),
    .Q(sig0000062a)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000474 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000006f8),
    .R(sig00000002),
    .Q(sig00000629)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000475 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000006f9),
    .R(sig00000002),
    .Q(NLW_blk00000475_Q_UNCONNECTED)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000476 (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000001dc),
    .Q(sig000006fa)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000477 (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000001db),
    .Q(sig000006fb)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000478 (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000001da),
    .Q(sig000006fc)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000479 (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000001d9),
    .Q(sig000006fd)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000047a (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000001d8),
    .Q(sig000006fe)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000047b (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000001d7),
    .Q(sig000006ff)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000047c (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000001d6),
    .Q(sig00000700)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000047d (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000001d5),
    .Q(sig00000701)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000047e (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000001d4),
    .Q(sig00000702)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000047f (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000001d3),
    .Q(sig00000703)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000480 (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000001d2),
    .Q(sig00000704)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000481 (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000001d1),
    .Q(sig00000705)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000482 (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000001d0),
    .Q(sig00000706)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000483 (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000001cf),
    .Q(sig00000707)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000484 (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000001ce),
    .Q(sig00000708)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000485 (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000001cd),
    .Q(sig00000709)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000486 (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000001cc),
    .Q(sig0000070a)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000487 (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000001cb),
    .Q(sig0000070b)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000488 (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000001ca),
    .Q(sig0000070c)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000489 (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000001c9),
    .Q(sig0000070d)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000048a (
    .C(clk),
    .CE(sig00000001),
    .D(sig000006fa),
    .R(sig00000002),
    .Q(sig0000060d)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000048b (
    .C(clk),
    .CE(sig00000001),
    .D(sig000006fb),
    .R(sig00000002),
    .Q(sig0000060c)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000048c (
    .C(clk),
    .CE(sig00000001),
    .D(sig000006fc),
    .R(sig00000002),
    .Q(sig0000060b)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000048d (
    .C(clk),
    .CE(sig00000001),
    .D(sig000006fd),
    .R(sig00000002),
    .Q(sig0000060a)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000048e (
    .C(clk),
    .CE(sig00000001),
    .D(sig000006fe),
    .R(sig00000002),
    .Q(sig00000609)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000048f (
    .C(clk),
    .CE(sig00000001),
    .D(sig000006ff),
    .R(sig00000002),
    .Q(sig00000608)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000490 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000700),
    .R(sig00000002),
    .Q(sig00000607)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000491 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000701),
    .R(sig00000002),
    .Q(sig00000606)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000492 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000702),
    .R(sig00000002),
    .Q(sig00000605)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000493 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000703),
    .R(sig00000002),
    .Q(sig00000604)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000494 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000704),
    .R(sig00000002),
    .Q(sig00000603)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000495 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000705),
    .R(sig00000002),
    .Q(sig00000602)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000496 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000706),
    .R(sig00000002),
    .Q(sig00000601)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000497 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000707),
    .R(sig00000002),
    .Q(sig00000600)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000498 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000708),
    .R(sig00000002),
    .Q(sig000005ff)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000499 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000709),
    .R(sig00000002),
    .Q(sig000005fe)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000049a (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000070a),
    .R(sig00000002),
    .Q(sig000005fd)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000049b (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000070b),
    .R(sig00000002),
    .Q(sig000005fc)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000049c (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000070c),
    .R(sig00000002),
    .Q(sig000005fb)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000049d (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000070d),
    .R(sig00000002),
    .Q(NLW_blk0000049d_Q_UNCONNECTED)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000582 (
    .I0(sig00000185),
    .I1(sig0000015f),
    .I2(sig00000007),
    .O(sig0000070e)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000583 (
    .I0(sig00000184),
    .I1(sig0000015e),
    .I2(sig00000007),
    .O(sig0000070f)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000584 (
    .I0(sig00000183),
    .I1(sig0000015d),
    .I2(sig00000007),
    .O(sig00000710)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000585 (
    .I0(sig00000182),
    .I1(sig0000015c),
    .I2(sig00000007),
    .O(sig00000711)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000586 (
    .I0(sig00000181),
    .I1(sig0000015b),
    .I2(sig00000007),
    .O(sig00000712)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000587 (
    .I0(sig00000180),
    .I1(sig0000015a),
    .I2(sig00000007),
    .O(sig00000713)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000588 (
    .I0(sig0000017f),
    .I1(sig00000159),
    .I2(sig00000007),
    .O(sig00000714)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000589 (
    .I0(sig0000017e),
    .I1(sig00000158),
    .I2(sig00000007),
    .O(sig00000715)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk0000058a (
    .I0(sig0000017d),
    .I1(sig00000157),
    .I2(sig00000007),
    .O(sig00000716)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk0000058b (
    .I0(sig0000017c),
    .I1(sig00000156),
    .I2(sig00000007),
    .O(sig00000717)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk0000058c (
    .I0(sig0000017b),
    .I1(sig00000155),
    .I2(sig00000007),
    .O(sig00000718)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk0000058d (
    .I0(sig0000017a),
    .I1(sig00000154),
    .I2(sig00000007),
    .O(sig00000719)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk0000058e (
    .I0(sig00000179),
    .I1(sig00000153),
    .I2(sig00000007),
    .O(sig0000071a)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk0000058f (
    .I0(sig00000178),
    .I1(sig00000152),
    .I2(sig00000007),
    .O(sig0000071b)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000590 (
    .I0(sig00000177),
    .I1(sig00000151),
    .I2(sig00000007),
    .O(sig0000071c)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000591 (
    .I0(sig00000176),
    .I1(sig00000150),
    .I2(sig00000007),
    .O(sig0000071d)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000592 (
    .I0(sig00000175),
    .I1(sig0000014f),
    .I2(sig00000007),
    .O(sig0000071e)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000593 (
    .I0(sig00000174),
    .I1(sig0000014e),
    .I2(sig00000007),
    .O(sig0000071f)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000594 (
    .I0(sig00000173),
    .I1(sig0000014d),
    .I2(sig00000007),
    .O(sig00000720)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000595 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000070e),
    .R(sig00000002),
    .Q(sig00000055)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000596 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000070f),
    .R(sig00000002),
    .Q(sig00000054)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000597 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000710),
    .R(sig00000002),
    .Q(sig00000053)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000598 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000711),
    .R(sig00000002),
    .Q(sig00000052)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000599 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000712),
    .R(sig00000002),
    .Q(sig00000051)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000059a (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000713),
    .R(sig00000002),
    .Q(sig00000050)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000059b (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000714),
    .R(sig00000002),
    .Q(sig0000004f)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000059c (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000715),
    .R(sig00000002),
    .Q(sig0000004e)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000059d (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000716),
    .R(sig00000002),
    .Q(sig0000004d)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000059e (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000717),
    .R(sig00000002),
    .Q(sig0000004c)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000059f (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000718),
    .R(sig00000002),
    .Q(sig0000004b)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000005a0 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000719),
    .R(sig00000002),
    .Q(sig0000004a)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000005a1 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000071a),
    .R(sig00000002),
    .Q(sig00000049)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000005a2 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000071b),
    .R(sig00000002),
    .Q(sig00000048)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000005a3 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000071c),
    .R(sig00000002),
    .Q(sig00000047)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000005a4 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000071d),
    .R(sig00000002),
    .Q(sig00000046)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000005a5 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000071e),
    .R(sig00000002),
    .Q(sig00000045)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000005a6 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000071f),
    .R(sig00000002),
    .Q(sig00000044)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000005a7 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000720),
    .R(sig00000002),
    .Q(sig00000043)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000005a8 (
    .I0(sig00000198),
    .I1(sig00000172),
    .I2(sig00000007),
    .O(sig00000721)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000005a9 (
    .I0(sig00000197),
    .I1(sig00000171),
    .I2(sig00000007),
    .O(sig00000722)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000005aa (
    .I0(sig00000196),
    .I1(sig00000170),
    .I2(sig00000007),
    .O(sig00000723)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000005ab (
    .I0(sig00000195),
    .I1(sig0000016f),
    .I2(sig00000007),
    .O(sig00000724)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000005ac (
    .I0(sig00000194),
    .I1(sig0000016e),
    .I2(sig00000007),
    .O(sig00000725)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000005ad (
    .I0(sig00000193),
    .I1(sig0000016d),
    .I2(sig00000007),
    .O(sig00000726)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000005ae (
    .I0(sig00000192),
    .I1(sig0000016c),
    .I2(sig00000007),
    .O(sig00000727)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000005af (
    .I0(sig00000191),
    .I1(sig0000016b),
    .I2(sig00000007),
    .O(sig00000728)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000005b0 (
    .I0(sig00000190),
    .I1(sig0000016a),
    .I2(sig00000007),
    .O(sig00000729)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000005b1 (
    .I0(sig0000018f),
    .I1(sig00000169),
    .I2(sig00000007),
    .O(sig0000072a)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000005b2 (
    .I0(sig0000018e),
    .I1(sig00000168),
    .I2(sig00000007),
    .O(sig0000072b)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000005b3 (
    .I0(sig0000018d),
    .I1(sig00000167),
    .I2(sig00000007),
    .O(sig0000072c)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000005b4 (
    .I0(sig0000018c),
    .I1(sig00000166),
    .I2(sig00000007),
    .O(sig0000072d)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000005b5 (
    .I0(sig0000018b),
    .I1(sig00000165),
    .I2(sig00000007),
    .O(sig0000072e)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000005b6 (
    .I0(sig0000018a),
    .I1(sig00000164),
    .I2(sig00000007),
    .O(sig0000072f)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000005b7 (
    .I0(sig00000189),
    .I1(sig00000163),
    .I2(sig00000007),
    .O(sig00000730)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000005b8 (
    .I0(sig00000188),
    .I1(sig00000162),
    .I2(sig00000007),
    .O(sig00000731)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000005b9 (
    .I0(sig00000187),
    .I1(sig00000161),
    .I2(sig00000007),
    .O(sig00000732)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000005ba (
    .I0(sig00000186),
    .I1(sig00000160),
    .I2(sig00000007),
    .O(sig00000733)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000005bb (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000721),
    .R(sig00000002),
    .Q(sig00000068)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000005bc (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000722),
    .R(sig00000002),
    .Q(sig00000067)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000005bd (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000723),
    .R(sig00000002),
    .Q(sig00000066)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000005be (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000724),
    .R(sig00000002),
    .Q(sig00000065)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000005bf (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000725),
    .R(sig00000002),
    .Q(sig00000064)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000005c0 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000726),
    .R(sig00000002),
    .Q(sig00000063)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000005c1 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000727),
    .R(sig00000002),
    .Q(sig00000062)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000005c2 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000728),
    .R(sig00000002),
    .Q(sig00000061)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000005c3 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000729),
    .R(sig00000002),
    .Q(sig00000060)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000005c4 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000072a),
    .R(sig00000002),
    .Q(sig0000005f)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000005c5 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000072b),
    .R(sig00000002),
    .Q(sig0000005e)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000005c6 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000072c),
    .R(sig00000002),
    .Q(sig0000005d)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000005c7 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000072d),
    .R(sig00000002),
    .Q(sig0000005c)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000005c8 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000072e),
    .R(sig00000002),
    .Q(sig0000005b)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000005c9 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000072f),
    .R(sig00000002),
    .Q(sig0000005a)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000005ca (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000730),
    .R(sig00000002),
    .Q(sig00000059)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000005cb (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000731),
    .R(sig00000002),
    .Q(sig00000058)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000005cc (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000732),
    .R(sig00000002),
    .Q(sig00000057)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000005cd (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000733),
    .R(sig00000002),
    .Q(sig00000056)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000005ce (
    .I0(sig00000185),
    .I1(sig0000015f),
    .I2(sig00000008),
    .O(sig00000734)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000005cf (
    .I0(sig00000184),
    .I1(sig0000015e),
    .I2(sig00000008),
    .O(sig00000735)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000005d0 (
    .I0(sig00000183),
    .I1(sig0000015d),
    .I2(sig00000008),
    .O(sig00000736)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000005d1 (
    .I0(sig00000182),
    .I1(sig0000015c),
    .I2(sig00000008),
    .O(sig00000737)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000005d2 (
    .I0(sig00000181),
    .I1(sig0000015b),
    .I2(sig00000008),
    .O(sig00000738)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000005d3 (
    .I0(sig00000180),
    .I1(sig0000015a),
    .I2(sig00000008),
    .O(sig00000739)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000005d4 (
    .I0(sig0000017f),
    .I1(sig00000159),
    .I2(sig00000008),
    .O(sig0000073a)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000005d5 (
    .I0(sig0000017e),
    .I1(sig00000158),
    .I2(sig00000008),
    .O(sig0000073b)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000005d6 (
    .I0(sig0000017d),
    .I1(sig00000157),
    .I2(sig00000008),
    .O(sig0000073c)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000005d7 (
    .I0(sig0000017c),
    .I1(sig00000156),
    .I2(sig00000008),
    .O(sig0000073d)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000005d8 (
    .I0(sig0000017b),
    .I1(sig00000155),
    .I2(sig00000008),
    .O(sig0000073e)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000005d9 (
    .I0(sig0000017a),
    .I1(sig00000154),
    .I2(sig00000008),
    .O(sig0000073f)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000005da (
    .I0(sig00000179),
    .I1(sig00000153),
    .I2(sig00000008),
    .O(sig00000740)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000005db (
    .I0(sig00000178),
    .I1(sig00000152),
    .I2(sig00000008),
    .O(sig00000741)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000005dc (
    .I0(sig00000177),
    .I1(sig00000151),
    .I2(sig00000008),
    .O(sig00000742)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000005dd (
    .I0(sig00000176),
    .I1(sig00000150),
    .I2(sig00000008),
    .O(sig00000743)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000005de (
    .I0(sig00000175),
    .I1(sig0000014f),
    .I2(sig00000008),
    .O(sig00000744)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000005df (
    .I0(sig00000174),
    .I1(sig0000014e),
    .I2(sig00000008),
    .O(sig00000745)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000005e0 (
    .I0(sig00000173),
    .I1(sig0000014d),
    .I2(sig00000008),
    .O(sig00000746)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000005e1 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000734),
    .R(sig00000002),
    .Q(sig0000007b)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000005e2 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000735),
    .R(sig00000002),
    .Q(sig0000007a)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000005e3 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000736),
    .R(sig00000002),
    .Q(sig00000079)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000005e4 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000737),
    .R(sig00000002),
    .Q(sig00000078)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000005e5 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000738),
    .R(sig00000002),
    .Q(sig00000077)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000005e6 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000739),
    .R(sig00000002),
    .Q(sig00000076)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000005e7 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000073a),
    .R(sig00000002),
    .Q(sig00000075)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000005e8 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000073b),
    .R(sig00000002),
    .Q(sig00000074)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000005e9 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000073c),
    .R(sig00000002),
    .Q(sig00000073)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000005ea (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000073d),
    .R(sig00000002),
    .Q(sig00000072)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000005eb (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000073e),
    .R(sig00000002),
    .Q(sig00000071)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000005ec (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000073f),
    .R(sig00000002),
    .Q(sig00000070)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000005ed (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000740),
    .R(sig00000002),
    .Q(sig0000006f)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000005ee (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000741),
    .R(sig00000002),
    .Q(sig0000006e)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000005ef (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000742),
    .R(sig00000002),
    .Q(sig0000006d)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000005f0 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000743),
    .R(sig00000002),
    .Q(sig0000006c)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000005f1 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000744),
    .R(sig00000002),
    .Q(sig0000006b)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000005f2 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000745),
    .R(sig00000002),
    .Q(sig0000006a)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000005f3 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000746),
    .R(sig00000002),
    .Q(sig00000069)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000005f4 (
    .I0(sig00000198),
    .I1(sig00000172),
    .I2(sig00000008),
    .O(sig00000747)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000005f5 (
    .I0(sig00000197),
    .I1(sig00000171),
    .I2(sig00000008),
    .O(sig00000748)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000005f6 (
    .I0(sig00000196),
    .I1(sig00000170),
    .I2(sig00000008),
    .O(sig00000749)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000005f7 (
    .I0(sig00000195),
    .I1(sig0000016f),
    .I2(sig00000008),
    .O(sig0000074a)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000005f8 (
    .I0(sig00000194),
    .I1(sig0000016e),
    .I2(sig00000008),
    .O(sig0000074b)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000005f9 (
    .I0(sig00000193),
    .I1(sig0000016d),
    .I2(sig00000008),
    .O(sig0000074c)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000005fa (
    .I0(sig00000192),
    .I1(sig0000016c),
    .I2(sig00000008),
    .O(sig0000074d)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000005fb (
    .I0(sig00000191),
    .I1(sig0000016b),
    .I2(sig00000008),
    .O(sig0000074e)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000005fc (
    .I0(sig00000190),
    .I1(sig0000016a),
    .I2(sig00000008),
    .O(sig0000074f)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000005fd (
    .I0(sig0000018f),
    .I1(sig00000169),
    .I2(sig00000008),
    .O(sig00000750)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000005fe (
    .I0(sig0000018e),
    .I1(sig00000168),
    .I2(sig00000008),
    .O(sig00000751)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk000005ff (
    .I0(sig0000018d),
    .I1(sig00000167),
    .I2(sig00000008),
    .O(sig00000752)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000600 (
    .I0(sig0000018c),
    .I1(sig00000166),
    .I2(sig00000008),
    .O(sig00000753)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000601 (
    .I0(sig0000018b),
    .I1(sig00000165),
    .I2(sig00000008),
    .O(sig00000754)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000602 (
    .I0(sig0000018a),
    .I1(sig00000164),
    .I2(sig00000008),
    .O(sig00000755)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000603 (
    .I0(sig00000189),
    .I1(sig00000163),
    .I2(sig00000008),
    .O(sig00000756)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000604 (
    .I0(sig00000188),
    .I1(sig00000162),
    .I2(sig00000008),
    .O(sig00000757)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000605 (
    .I0(sig00000187),
    .I1(sig00000161),
    .I2(sig00000008),
    .O(sig00000758)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000606 (
    .I0(sig00000186),
    .I1(sig00000160),
    .I2(sig00000008),
    .O(sig00000759)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000607 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000747),
    .R(sig00000002),
    .Q(sig0000008e)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000608 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000748),
    .R(sig00000002),
    .Q(sig0000008d)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000609 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000749),
    .R(sig00000002),
    .Q(sig0000008c)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000060a (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000074a),
    .R(sig00000002),
    .Q(sig0000008b)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000060b (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000074b),
    .R(sig00000002),
    .Q(sig0000008a)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000060c (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000074c),
    .R(sig00000002),
    .Q(sig00000089)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000060d (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000074d),
    .R(sig00000002),
    .Q(sig00000088)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000060e (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000074e),
    .R(sig00000002),
    .Q(sig00000087)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000060f (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000074f),
    .R(sig00000002),
    .Q(sig00000086)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000610 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000750),
    .R(sig00000002),
    .Q(sig00000085)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000611 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000751),
    .R(sig00000002),
    .Q(sig00000084)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000612 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000752),
    .R(sig00000002),
    .Q(sig00000083)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000613 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000753),
    .R(sig00000002),
    .Q(sig00000082)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000614 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000754),
    .R(sig00000002),
    .Q(sig00000081)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000615 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000755),
    .R(sig00000002),
    .Q(sig00000080)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000616 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000756),
    .R(sig00000002),
    .Q(sig0000007f)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000617 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000757),
    .R(sig00000002),
    .Q(sig0000007e)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000618 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000758),
    .R(sig00000002),
    .Q(sig0000007d)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000619 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000759),
    .R(sig00000002),
    .Q(sig0000007c)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk0000061a (
    .I0(sig00000185),
    .I1(sig0000015f),
    .I2(sig0000000c),
    .O(sig0000075a)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk0000061b (
    .I0(sig00000184),
    .I1(sig0000015e),
    .I2(sig0000000c),
    .O(sig0000075b)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk0000061c (
    .I0(sig00000183),
    .I1(sig0000015d),
    .I2(sig0000000c),
    .O(sig0000075c)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk0000061d (
    .I0(sig00000182),
    .I1(sig0000015c),
    .I2(sig0000000c),
    .O(sig0000075d)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk0000061e (
    .I0(sig00000181),
    .I1(sig0000015b),
    .I2(sig0000000c),
    .O(sig0000075e)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk0000061f (
    .I0(sig00000180),
    .I1(sig0000015a),
    .I2(sig0000000c),
    .O(sig0000075f)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000620 (
    .I0(sig0000017f),
    .I1(sig00000159),
    .I2(sig0000000c),
    .O(sig00000760)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000621 (
    .I0(sig0000017e),
    .I1(sig00000158),
    .I2(sig0000000c),
    .O(sig00000761)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000622 (
    .I0(sig0000017d),
    .I1(sig00000157),
    .I2(sig0000000c),
    .O(sig00000762)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000623 (
    .I0(sig0000017c),
    .I1(sig00000156),
    .I2(sig0000000c),
    .O(sig00000763)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000624 (
    .I0(sig0000017b),
    .I1(sig00000155),
    .I2(sig0000000c),
    .O(sig00000764)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000625 (
    .I0(sig0000017a),
    .I1(sig00000154),
    .I2(sig0000000c),
    .O(sig00000765)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000626 (
    .I0(sig00000179),
    .I1(sig00000153),
    .I2(sig0000000c),
    .O(sig00000766)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000627 (
    .I0(sig00000178),
    .I1(sig00000152),
    .I2(sig0000000c),
    .O(sig00000767)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000628 (
    .I0(sig00000177),
    .I1(sig00000151),
    .I2(sig0000000c),
    .O(sig00000768)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000629 (
    .I0(sig00000176),
    .I1(sig00000150),
    .I2(sig0000000c),
    .O(sig00000769)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk0000062a (
    .I0(sig00000175),
    .I1(sig0000014f),
    .I2(sig0000000c),
    .O(sig0000076a)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk0000062b (
    .I0(sig00000174),
    .I1(sig0000014e),
    .I2(sig0000000c),
    .O(sig0000076b)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk0000062c (
    .I0(sig00000173),
    .I1(sig0000014d),
    .I2(sig0000000c),
    .O(sig0000076c)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000062d (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000075a),
    .R(sig00000002),
    .Q(\U0/i_synth/non_floating_point.arch_c.xfft_inst/single_channel.datapath/output_selector_im/Q [18])
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000062e (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000075b),
    .R(sig00000002),
    .Q(\U0/i_synth/non_floating_point.arch_c.xfft_inst/single_channel.datapath/output_selector_im/Q [17])
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000062f (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000075c),
    .R(sig00000002),
    .Q(\U0/i_synth/non_floating_point.arch_c.xfft_inst/single_channel.datapath/output_selector_im/Q [16])
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000630 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000075d),
    .R(sig00000002),
    .Q(\U0/i_synth/non_floating_point.arch_c.xfft_inst/single_channel.datapath/output_selector_im/Q [15])
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000631 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000075e),
    .R(sig00000002),
    .Q(\U0/i_synth/non_floating_point.arch_c.xfft_inst/single_channel.datapath/output_selector_im/Q [14])
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000632 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000075f),
    .R(sig00000002),
    .Q(\U0/i_synth/non_floating_point.arch_c.xfft_inst/single_channel.datapath/output_selector_im/Q [13])
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000633 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000760),
    .R(sig00000002),
    .Q(\U0/i_synth/non_floating_point.arch_c.xfft_inst/single_channel.datapath/output_selector_im/Q [12])
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000634 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000761),
    .R(sig00000002),
    .Q(\U0/i_synth/non_floating_point.arch_c.xfft_inst/single_channel.datapath/output_selector_im/Q [11])
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000635 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000762),
    .R(sig00000002),
    .Q(\U0/i_synth/non_floating_point.arch_c.xfft_inst/single_channel.datapath/output_selector_im/Q [10])
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000636 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000763),
    .R(sig00000002),
    .Q(\U0/i_synth/non_floating_point.arch_c.xfft_inst/single_channel.datapath/output_selector_im/Q [9])
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000637 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000764),
    .R(sig00000002),
    .Q(\U0/i_synth/non_floating_point.arch_c.xfft_inst/single_channel.datapath/output_selector_im/Q [8])
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000638 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000765),
    .R(sig00000002),
    .Q(\U0/i_synth/non_floating_point.arch_c.xfft_inst/single_channel.datapath/output_selector_im/Q [7])
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000639 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000766),
    .R(sig00000002),
    .Q(\U0/i_synth/non_floating_point.arch_c.xfft_inst/single_channel.datapath/output_selector_im/Q [6])
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000063a (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000767),
    .R(sig00000002),
    .Q(\U0/i_synth/non_floating_point.arch_c.xfft_inst/single_channel.datapath/output_selector_im/Q [5])
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000063b (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000768),
    .R(sig00000002),
    .Q(\U0/i_synth/non_floating_point.arch_c.xfft_inst/single_channel.datapath/output_selector_im/Q [4])
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000063c (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000769),
    .R(sig00000002),
    .Q(\U0/i_synth/non_floating_point.arch_c.xfft_inst/single_channel.datapath/output_selector_im/Q [3])
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000063d (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000076a),
    .R(sig00000002),
    .Q(\U0/i_synth/non_floating_point.arch_c.xfft_inst/single_channel.datapath/output_selector_im/Q [2])
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000063e (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000076b),
    .R(sig00000002),
    .Q(\U0/i_synth/non_floating_point.arch_c.xfft_inst/single_channel.datapath/output_selector_im/Q [1])
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000063f (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000076c),
    .R(sig00000002),
    .Q(\U0/i_synth/non_floating_point.arch_c.xfft_inst/single_channel.datapath/output_selector_im/Q [0])
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000640 (
    .I0(sig00000198),
    .I1(sig00000172),
    .I2(sig0000000c),
    .O(sig0000076d)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000641 (
    .I0(sig00000197),
    .I1(sig00000171),
    .I2(sig0000000c),
    .O(sig0000076e)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000642 (
    .I0(sig00000196),
    .I1(sig00000170),
    .I2(sig0000000c),
    .O(sig0000076f)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000643 (
    .I0(sig00000195),
    .I1(sig0000016f),
    .I2(sig0000000c),
    .O(sig00000770)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000644 (
    .I0(sig00000194),
    .I1(sig0000016e),
    .I2(sig0000000c),
    .O(sig00000771)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000645 (
    .I0(sig00000193),
    .I1(sig0000016d),
    .I2(sig0000000c),
    .O(sig00000772)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000646 (
    .I0(sig00000192),
    .I1(sig0000016c),
    .I2(sig0000000c),
    .O(sig00000773)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000647 (
    .I0(sig00000191),
    .I1(sig0000016b),
    .I2(sig0000000c),
    .O(sig00000774)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000648 (
    .I0(sig00000190),
    .I1(sig0000016a),
    .I2(sig0000000c),
    .O(sig00000775)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000649 (
    .I0(sig0000018f),
    .I1(sig00000169),
    .I2(sig0000000c),
    .O(sig00000776)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk0000064a (
    .I0(sig0000018e),
    .I1(sig00000168),
    .I2(sig0000000c),
    .O(sig00000777)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk0000064b (
    .I0(sig0000018d),
    .I1(sig00000167),
    .I2(sig0000000c),
    .O(sig00000778)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk0000064c (
    .I0(sig0000018c),
    .I1(sig00000166),
    .I2(sig0000000c),
    .O(sig00000779)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk0000064d (
    .I0(sig0000018b),
    .I1(sig00000165),
    .I2(sig0000000c),
    .O(sig0000077a)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk0000064e (
    .I0(sig0000018a),
    .I1(sig00000164),
    .I2(sig0000000c),
    .O(sig0000077b)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk0000064f (
    .I0(sig00000189),
    .I1(sig00000163),
    .I2(sig0000000c),
    .O(sig0000077c)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000650 (
    .I0(sig00000188),
    .I1(sig00000162),
    .I2(sig0000000c),
    .O(sig0000077d)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000651 (
    .I0(sig00000187),
    .I1(sig00000161),
    .I2(sig0000000c),
    .O(sig0000077e)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000652 (
    .I0(sig00000186),
    .I1(sig00000160),
    .I2(sig0000000c),
    .O(sig0000077f)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000653 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000076d),
    .R(sig00000002),
    .Q(\U0/i_synth/non_floating_point.arch_c.xfft_inst/single_channel.datapath/output_selector_re/Q [18])
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000654 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000076e),
    .R(sig00000002),
    .Q(\U0/i_synth/non_floating_point.arch_c.xfft_inst/single_channel.datapath/output_selector_re/Q [17])
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000655 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000076f),
    .R(sig00000002),
    .Q(\U0/i_synth/non_floating_point.arch_c.xfft_inst/single_channel.datapath/output_selector_re/Q [16])
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000656 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000770),
    .R(sig00000002),
    .Q(\U0/i_synth/non_floating_point.arch_c.xfft_inst/single_channel.datapath/output_selector_re/Q [15])
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000657 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000771),
    .R(sig00000002),
    .Q(\U0/i_synth/non_floating_point.arch_c.xfft_inst/single_channel.datapath/output_selector_re/Q [14])
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000658 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000772),
    .R(sig00000002),
    .Q(\U0/i_synth/non_floating_point.arch_c.xfft_inst/single_channel.datapath/output_selector_re/Q [13])
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000659 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000773),
    .R(sig00000002),
    .Q(\U0/i_synth/non_floating_point.arch_c.xfft_inst/single_channel.datapath/output_selector_re/Q [12])
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000065a (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000774),
    .R(sig00000002),
    .Q(\U0/i_synth/non_floating_point.arch_c.xfft_inst/single_channel.datapath/output_selector_re/Q [11])
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000065b (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000775),
    .R(sig00000002),
    .Q(\U0/i_synth/non_floating_point.arch_c.xfft_inst/single_channel.datapath/output_selector_re/Q [10])
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000065c (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000776),
    .R(sig00000002),
    .Q(\U0/i_synth/non_floating_point.arch_c.xfft_inst/single_channel.datapath/output_selector_re/Q [9])
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000065d (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000777),
    .R(sig00000002),
    .Q(\U0/i_synth/non_floating_point.arch_c.xfft_inst/single_channel.datapath/output_selector_re/Q [8])
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000065e (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000778),
    .R(sig00000002),
    .Q(\U0/i_synth/non_floating_point.arch_c.xfft_inst/single_channel.datapath/output_selector_re/Q [7])
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000065f (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000779),
    .R(sig00000002),
    .Q(\U0/i_synth/non_floating_point.arch_c.xfft_inst/single_channel.datapath/output_selector_re/Q [6])
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000660 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000077a),
    .R(sig00000002),
    .Q(\U0/i_synth/non_floating_point.arch_c.xfft_inst/single_channel.datapath/output_selector_re/Q [5])
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000661 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000077b),
    .R(sig00000002),
    .Q(\U0/i_synth/non_floating_point.arch_c.xfft_inst/single_channel.datapath/output_selector_re/Q [4])
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000662 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000077c),
    .R(sig00000002),
    .Q(\U0/i_synth/non_floating_point.arch_c.xfft_inst/single_channel.datapath/output_selector_re/Q [3])
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000663 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000077d),
    .R(sig00000002),
    .Q(\U0/i_synth/non_floating_point.arch_c.xfft_inst/single_channel.datapath/output_selector_re/Q [2])
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000664 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000077e),
    .R(sig00000002),
    .Q(\U0/i_synth/non_floating_point.arch_c.xfft_inst/single_channel.datapath/output_selector_re/Q [1])
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000665 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000077f),
    .R(sig00000002),
    .Q(\U0/i_synth/non_floating_point.arch_c.xfft_inst/single_channel.datapath/output_selector_re/Q [0])
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000666 (
    .A0(sig00000001),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(xn_im[8]),
    .Q(sig00000780)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000667 (
    .A0(sig00000001),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(xn_im[8]),
    .Q(sig00000781)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000668 (
    .A0(sig00000001),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(xn_im[8]),
    .Q(sig00000782)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000669 (
    .A0(sig00000001),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(xn_im[8]),
    .Q(sig00000783)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000066a (
    .A0(sig00000001),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(xn_im[8]),
    .Q(sig00000784)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000066b (
    .A0(sig00000001),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(xn_im[8]),
    .Q(sig00000785)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000066c (
    .A0(sig00000001),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(xn_im[8]),
    .Q(sig00000786)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000066d (
    .A0(sig00000001),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(xn_im[8]),
    .Q(sig00000787)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000066e (
    .A0(sig00000001),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(xn_im[8]),
    .Q(sig00000788)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000066f (
    .A0(sig00000001),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(xn_im[8]),
    .Q(sig00000789)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000670 (
    .A0(sig00000001),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(xn_im[8]),
    .Q(sig0000078a)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000671 (
    .A0(sig00000001),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(xn_im[7]),
    .Q(sig0000078b)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000672 (
    .A0(sig00000001),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(xn_im[6]),
    .Q(sig0000078c)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000673 (
    .A0(sig00000001),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(xn_im[5]),
    .Q(sig0000078d)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000674 (
    .A0(sig00000001),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(xn_im[4]),
    .Q(sig0000078e)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000675 (
    .A0(sig00000001),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(xn_im[3]),
    .Q(sig0000078f)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000676 (
    .A0(sig00000001),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(xn_im[2]),
    .Q(sig00000790)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000677 (
    .A0(sig00000001),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(xn_im[1]),
    .Q(sig00000791)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000678 (
    .A0(sig00000001),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(xn_im[0]),
    .Q(sig00000792)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000679 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000780),
    .R(sig00000002),
    .Q(sig000000ed)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000067a (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000781),
    .R(sig00000002),
    .Q(sig000000ec)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000067b (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000782),
    .R(sig00000002),
    .Q(sig000000eb)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000067c (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000783),
    .R(sig00000002),
    .Q(sig000000ea)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000067d (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000784),
    .R(sig00000002),
    .Q(sig000000e9)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000067e (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000785),
    .R(sig00000002),
    .Q(sig000000e8)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000067f (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000786),
    .R(sig00000002),
    .Q(sig000000e7)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000680 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000787),
    .R(sig00000002),
    .Q(sig000000e6)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000681 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000788),
    .R(sig00000002),
    .Q(sig000000e5)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000682 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000789),
    .R(sig00000002),
    .Q(sig000000e4)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000683 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000078a),
    .R(sig00000002),
    .Q(sig000000e3)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000684 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000078b),
    .R(sig00000002),
    .Q(sig000000e2)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000685 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000078c),
    .R(sig00000002),
    .Q(sig000000e1)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000686 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000078d),
    .R(sig00000002),
    .Q(sig000000e0)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000687 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000078e),
    .R(sig00000002),
    .Q(sig000000df)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000688 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000078f),
    .R(sig00000002),
    .Q(sig000000de)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000689 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000790),
    .R(sig00000002),
    .Q(sig000000dd)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000068a (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000791),
    .R(sig00000002),
    .Q(sig000000dc)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000068b (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000792),
    .R(sig00000002),
    .Q(sig000000db)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000068c (
    .A0(sig00000001),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(xn_re[8]),
    .Q(sig00000793)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000068d (
    .A0(sig00000001),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(xn_re[8]),
    .Q(sig00000794)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000068e (
    .A0(sig00000001),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(xn_re[8]),
    .Q(sig00000795)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000068f (
    .A0(sig00000001),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(xn_re[8]),
    .Q(sig00000796)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000690 (
    .A0(sig00000001),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(xn_re[8]),
    .Q(sig00000797)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000691 (
    .A0(sig00000001),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(xn_re[8]),
    .Q(sig00000798)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000692 (
    .A0(sig00000001),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(xn_re[8]),
    .Q(sig00000799)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000693 (
    .A0(sig00000001),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(xn_re[8]),
    .Q(sig0000079a)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000694 (
    .A0(sig00000001),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(xn_re[8]),
    .Q(sig0000079b)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000695 (
    .A0(sig00000001),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(xn_re[8]),
    .Q(sig0000079c)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000696 (
    .A0(sig00000001),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(xn_re[8]),
    .Q(sig0000079d)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000697 (
    .A0(sig00000001),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(xn_re[7]),
    .Q(sig0000079e)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000698 (
    .A0(sig00000001),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(xn_re[6]),
    .Q(sig0000079f)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk00000699 (
    .A0(sig00000001),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(xn_re[5]),
    .Q(sig000007a0)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000069a (
    .A0(sig00000001),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(xn_re[4]),
    .Q(sig000007a1)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000069b (
    .A0(sig00000001),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(xn_re[3]),
    .Q(sig000007a2)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000069c (
    .A0(sig00000001),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(xn_re[2]),
    .Q(sig000007a3)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000069d (
    .A0(sig00000001),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(xn_re[1]),
    .Q(sig000007a4)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000069e (
    .A0(sig00000001),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(xn_re[0]),
    .Q(sig000007a5)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000069f (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000793),
    .R(sig00000002),
    .Q(sig00000100)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000006a0 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000794),
    .R(sig00000002),
    .Q(sig000000ff)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000006a1 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000795),
    .R(sig00000002),
    .Q(sig000000fe)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000006a2 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000796),
    .R(sig00000002),
    .Q(sig000000fd)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000006a3 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000797),
    .R(sig00000002),
    .Q(sig000000fc)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000006a4 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000798),
    .R(sig00000002),
    .Q(sig000000fb)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000006a5 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000799),
    .R(sig00000002),
    .Q(sig000000fa)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000006a6 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000079a),
    .R(sig00000002),
    .Q(sig000000f9)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000006a7 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000079b),
    .R(sig00000002),
    .Q(sig000000f8)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000006a8 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000079c),
    .R(sig00000002),
    .Q(sig000000f7)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000006a9 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000079d),
    .R(sig00000002),
    .Q(sig000000f6)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000006aa (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000079e),
    .R(sig00000002),
    .Q(sig000000f5)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000006ab (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000079f),
    .R(sig00000002),
    .Q(sig000000f4)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000006ac (
    .C(clk),
    .CE(sig00000001),
    .D(sig000007a0),
    .R(sig00000002),
    .Q(sig000000f3)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000006ad (
    .C(clk),
    .CE(sig00000001),
    .D(sig000007a1),
    .R(sig00000002),
    .Q(sig000000f2)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000006ae (
    .C(clk),
    .CE(sig00000001),
    .D(sig000007a2),
    .R(sig00000002),
    .Q(sig000000f1)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000006af (
    .C(clk),
    .CE(sig00000001),
    .D(sig000007a3),
    .R(sig00000002),
    .Q(sig000000f0)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000006b0 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000007a4),
    .R(sig00000002),
    .Q(sig000000ef)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000006b1 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000007a5),
    .R(sig00000002),
    .Q(sig000000ee)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000006b2 (
    .I0(sig0000013a),
    .I1(sig00000114),
    .I2(sig000000db),
    .I3(sig000000db),
    .I4(sig00000004),
    .I5(sig0000000b),
    .O(sig000007a6)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000006b3 (
    .I0(sig0000013b),
    .I1(sig00000115),
    .I2(sig000000dc),
    .I3(sig000000dc),
    .I4(sig00000004),
    .I5(sig0000000b),
    .O(sig000007a7)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000006b4 (
    .I0(sig0000013c),
    .I1(sig00000116),
    .I2(sig000000dd),
    .I3(sig000000dd),
    .I4(sig00000004),
    .I5(sig0000000b),
    .O(sig000007a8)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000006b5 (
    .I0(sig0000013d),
    .I1(sig00000117),
    .I2(sig000000de),
    .I3(sig000000de),
    .I4(sig00000004),
    .I5(sig0000000b),
    .O(sig000007a9)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000006b6 (
    .I0(sig0000013e),
    .I1(sig00000118),
    .I2(sig000000df),
    .I3(sig000000df),
    .I4(sig00000004),
    .I5(sig0000000b),
    .O(sig000007aa)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000006b7 (
    .I0(sig0000013f),
    .I1(sig00000119),
    .I2(sig000000e0),
    .I3(sig000000e0),
    .I4(sig00000004),
    .I5(sig0000000b),
    .O(sig000007ab)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000006b8 (
    .I0(sig00000140),
    .I1(sig0000011a),
    .I2(sig000000e1),
    .I3(sig000000e1),
    .I4(sig00000004),
    .I5(sig0000000b),
    .O(sig000007ac)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000006b9 (
    .I0(sig00000141),
    .I1(sig0000011b),
    .I2(sig000000e2),
    .I3(sig000000e2),
    .I4(sig00000004),
    .I5(sig0000000b),
    .O(sig000007ad)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000006ba (
    .I0(sig00000142),
    .I1(sig0000011c),
    .I2(sig000000e3),
    .I3(sig000000e3),
    .I4(sig00000004),
    .I5(sig0000000b),
    .O(sig000007ae)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000006bb (
    .I0(sig00000143),
    .I1(sig0000011d),
    .I2(sig000000e4),
    .I3(sig000000e4),
    .I4(sig00000004),
    .I5(sig0000000b),
    .O(sig000007af)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000006bc (
    .I0(sig00000144),
    .I1(sig0000011e),
    .I2(sig000000e5),
    .I3(sig000000e5),
    .I4(sig00000004),
    .I5(sig0000000b),
    .O(sig000007b0)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000006bd (
    .I0(sig00000145),
    .I1(sig0000011f),
    .I2(sig000000e6),
    .I3(sig000000e6),
    .I4(sig00000004),
    .I5(sig0000000b),
    .O(sig000007b1)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000006be (
    .I0(sig00000146),
    .I1(sig00000120),
    .I2(sig000000e7),
    .I3(sig000000e7),
    .I4(sig00000004),
    .I5(sig0000000b),
    .O(sig000007b2)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000006bf (
    .I0(sig00000147),
    .I1(sig00000121),
    .I2(sig000000e8),
    .I3(sig000000e8),
    .I4(sig00000004),
    .I5(sig0000000b),
    .O(sig000007b3)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000006c0 (
    .I0(sig00000148),
    .I1(sig00000122),
    .I2(sig000000e9),
    .I3(sig000000e9),
    .I4(sig00000004),
    .I5(sig0000000b),
    .O(sig000007b4)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000006c1 (
    .I0(sig00000149),
    .I1(sig00000123),
    .I2(sig000000ea),
    .I3(sig000000ea),
    .I4(sig00000004),
    .I5(sig0000000b),
    .O(sig000007b5)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000006c2 (
    .I0(sig0000014a),
    .I1(sig00000124),
    .I2(sig000000eb),
    .I3(sig000000eb),
    .I4(sig00000004),
    .I5(sig0000000b),
    .O(sig000007b6)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000006c3 (
    .I0(sig0000014b),
    .I1(sig00000125),
    .I2(sig000000ec),
    .I3(sig000000ec),
    .I4(sig00000004),
    .I5(sig0000000b),
    .O(sig000007b7)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000006c4 (
    .I0(sig0000014c),
    .I1(sig00000126),
    .I2(sig000000ed),
    .I3(sig000000ed),
    .I4(sig00000004),
    .I5(sig0000000b),
    .O(sig000007b8)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000006c5 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000007a6),
    .R(sig00000002),
    .Q(sig0000008f)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000006c6 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000007a7),
    .R(sig00000002),
    .Q(sig00000090)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000006c7 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000007a8),
    .R(sig00000002),
    .Q(sig00000091)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000006c8 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000007a9),
    .R(sig00000002),
    .Q(sig00000092)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000006c9 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000007aa),
    .R(sig00000002),
    .Q(sig00000093)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000006ca (
    .C(clk),
    .CE(sig00000001),
    .D(sig000007ab),
    .R(sig00000002),
    .Q(sig00000094)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000006cb (
    .C(clk),
    .CE(sig00000001),
    .D(sig000007ac),
    .R(sig00000002),
    .Q(sig00000095)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000006cc (
    .C(clk),
    .CE(sig00000001),
    .D(sig000007ad),
    .R(sig00000002),
    .Q(sig00000096)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000006cd (
    .C(clk),
    .CE(sig00000001),
    .D(sig000007ae),
    .R(sig00000002),
    .Q(sig00000097)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000006ce (
    .C(clk),
    .CE(sig00000001),
    .D(sig000007af),
    .R(sig00000002),
    .Q(sig00000098)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000006cf (
    .C(clk),
    .CE(sig00000001),
    .D(sig000007b0),
    .R(sig00000002),
    .Q(sig00000099)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000006d0 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000007b1),
    .R(sig00000002),
    .Q(sig0000009a)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000006d1 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000007b2),
    .R(sig00000002),
    .Q(sig0000009b)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000006d2 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000007b3),
    .R(sig00000002),
    .Q(sig0000009c)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000006d3 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000007b4),
    .R(sig00000002),
    .Q(sig0000009d)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000006d4 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000007b5),
    .R(sig00000002),
    .Q(sig0000009e)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000006d5 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000007b6),
    .R(sig00000002),
    .Q(sig0000009f)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000006d6 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000007b7),
    .R(sig00000002),
    .Q(sig000000a0)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000006d7 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000007b8),
    .R(sig00000002),
    .Q(sig000000a1)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000006d8 (
    .I0(sig00000127),
    .I1(sig00000101),
    .I2(sig000000ee),
    .I3(sig000000ee),
    .I4(sig00000004),
    .I5(sig0000000b),
    .O(sig000007b9)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000006d9 (
    .I0(sig00000128),
    .I1(sig00000102),
    .I2(sig000000ef),
    .I3(sig000000ef),
    .I4(sig00000004),
    .I5(sig0000000b),
    .O(sig000007ba)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000006da (
    .I0(sig00000129),
    .I1(sig00000103),
    .I2(sig000000f0),
    .I3(sig000000f0),
    .I4(sig00000004),
    .I5(sig0000000b),
    .O(sig000007bb)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000006db (
    .I0(sig0000012a),
    .I1(sig00000104),
    .I2(sig000000f1),
    .I3(sig000000f1),
    .I4(sig00000004),
    .I5(sig0000000b),
    .O(sig000007bc)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000006dc (
    .I0(sig0000012b),
    .I1(sig00000105),
    .I2(sig000000f2),
    .I3(sig000000f2),
    .I4(sig00000004),
    .I5(sig0000000b),
    .O(sig000007bd)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000006dd (
    .I0(sig0000012c),
    .I1(sig00000106),
    .I2(sig000000f3),
    .I3(sig000000f3),
    .I4(sig00000004),
    .I5(sig0000000b),
    .O(sig000007be)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000006de (
    .I0(sig0000012d),
    .I1(sig00000107),
    .I2(sig000000f4),
    .I3(sig000000f4),
    .I4(sig00000004),
    .I5(sig0000000b),
    .O(sig000007bf)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000006df (
    .I0(sig0000012e),
    .I1(sig00000108),
    .I2(sig000000f5),
    .I3(sig000000f5),
    .I4(sig00000004),
    .I5(sig0000000b),
    .O(sig000007c0)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000006e0 (
    .I0(sig0000012f),
    .I1(sig00000109),
    .I2(sig000000f6),
    .I3(sig000000f6),
    .I4(sig00000004),
    .I5(sig0000000b),
    .O(sig000007c1)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000006e1 (
    .I0(sig00000130),
    .I1(sig0000010a),
    .I2(sig000000f7),
    .I3(sig000000f7),
    .I4(sig00000004),
    .I5(sig0000000b),
    .O(sig000007c2)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000006e2 (
    .I0(sig00000131),
    .I1(sig0000010b),
    .I2(sig000000f8),
    .I3(sig000000f8),
    .I4(sig00000004),
    .I5(sig0000000b),
    .O(sig000007c3)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000006e3 (
    .I0(sig00000132),
    .I1(sig0000010c),
    .I2(sig000000f9),
    .I3(sig000000f9),
    .I4(sig00000004),
    .I5(sig0000000b),
    .O(sig000007c4)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000006e4 (
    .I0(sig00000133),
    .I1(sig0000010d),
    .I2(sig000000fa),
    .I3(sig000000fa),
    .I4(sig00000004),
    .I5(sig0000000b),
    .O(sig000007c5)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000006e5 (
    .I0(sig00000134),
    .I1(sig0000010e),
    .I2(sig000000fb),
    .I3(sig000000fb),
    .I4(sig00000004),
    .I5(sig0000000b),
    .O(sig000007c6)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000006e6 (
    .I0(sig00000135),
    .I1(sig0000010f),
    .I2(sig000000fc),
    .I3(sig000000fc),
    .I4(sig00000004),
    .I5(sig0000000b),
    .O(sig000007c7)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000006e7 (
    .I0(sig00000136),
    .I1(sig00000110),
    .I2(sig000000fd),
    .I3(sig000000fd),
    .I4(sig00000004),
    .I5(sig0000000b),
    .O(sig000007c8)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000006e8 (
    .I0(sig00000137),
    .I1(sig00000111),
    .I2(sig000000fe),
    .I3(sig000000fe),
    .I4(sig00000004),
    .I5(sig0000000b),
    .O(sig000007c9)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000006e9 (
    .I0(sig00000138),
    .I1(sig00000112),
    .I2(sig000000ff),
    .I3(sig000000ff),
    .I4(sig00000004),
    .I5(sig0000000b),
    .O(sig000007ca)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000006ea (
    .I0(sig00000139),
    .I1(sig00000113),
    .I2(sig00000100),
    .I3(sig00000100),
    .I4(sig00000004),
    .I5(sig0000000b),
    .O(sig000007cb)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000006eb (
    .C(clk),
    .CE(sig00000001),
    .D(sig000007b9),
    .R(sig00000002),
    .Q(sig000000a2)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000006ec (
    .C(clk),
    .CE(sig00000001),
    .D(sig000007ba),
    .R(sig00000002),
    .Q(sig000000a3)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000006ed (
    .C(clk),
    .CE(sig00000001),
    .D(sig000007bb),
    .R(sig00000002),
    .Q(sig000000a4)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000006ee (
    .C(clk),
    .CE(sig00000001),
    .D(sig000007bc),
    .R(sig00000002),
    .Q(sig000000a5)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000006ef (
    .C(clk),
    .CE(sig00000001),
    .D(sig000007bd),
    .R(sig00000002),
    .Q(sig000000a6)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000006f0 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000007be),
    .R(sig00000002),
    .Q(sig000000a7)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000006f1 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000007bf),
    .R(sig00000002),
    .Q(sig000000a8)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000006f2 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000007c0),
    .R(sig00000002),
    .Q(sig000000a9)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000006f3 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000007c1),
    .R(sig00000002),
    .Q(sig000000aa)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000006f4 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000007c2),
    .R(sig00000002),
    .Q(sig000000ab)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000006f5 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000007c3),
    .R(sig00000002),
    .Q(sig000000ac)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000006f6 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000007c4),
    .R(sig00000002),
    .Q(sig000000ad)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000006f7 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000007c5),
    .R(sig00000002),
    .Q(sig000000ae)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000006f8 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000007c6),
    .R(sig00000002),
    .Q(sig000000af)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000006f9 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000007c7),
    .R(sig00000002),
    .Q(sig000000b0)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000006fa (
    .C(clk),
    .CE(sig00000001),
    .D(sig000007c8),
    .R(sig00000002),
    .Q(sig000000b1)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000006fb (
    .C(clk),
    .CE(sig00000001),
    .D(sig000007c9),
    .R(sig00000002),
    .Q(sig000000b2)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000006fc (
    .C(clk),
    .CE(sig00000001),
    .D(sig000007ca),
    .R(sig00000002),
    .Q(sig000000b3)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000006fd (
    .C(clk),
    .CE(sig00000001),
    .D(sig000007cb),
    .R(sig00000002),
    .Q(sig000000b4)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000006fe (
    .I0(sig0000013a),
    .I1(sig00000114),
    .I2(sig000000db),
    .I3(sig000000db),
    .I4(sig00000005),
    .I5(sig0000000b),
    .O(sig000007cc)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000006ff (
    .I0(sig0000013b),
    .I1(sig00000115),
    .I2(sig000000dc),
    .I3(sig000000dc),
    .I4(sig00000005),
    .I5(sig0000000b),
    .O(sig000007cd)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk00000700 (
    .I0(sig0000013c),
    .I1(sig00000116),
    .I2(sig000000dd),
    .I3(sig000000dd),
    .I4(sig00000005),
    .I5(sig0000000b),
    .O(sig000007ce)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk00000701 (
    .I0(sig0000013d),
    .I1(sig00000117),
    .I2(sig000000de),
    .I3(sig000000de),
    .I4(sig00000005),
    .I5(sig0000000b),
    .O(sig000007cf)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk00000702 (
    .I0(sig0000013e),
    .I1(sig00000118),
    .I2(sig000000df),
    .I3(sig000000df),
    .I4(sig00000005),
    .I5(sig0000000b),
    .O(sig000007d0)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk00000703 (
    .I0(sig0000013f),
    .I1(sig00000119),
    .I2(sig000000e0),
    .I3(sig000000e0),
    .I4(sig00000005),
    .I5(sig0000000b),
    .O(sig000007d1)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk00000704 (
    .I0(sig00000140),
    .I1(sig0000011a),
    .I2(sig000000e1),
    .I3(sig000000e1),
    .I4(sig00000005),
    .I5(sig0000000b),
    .O(sig000007d2)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk00000705 (
    .I0(sig00000141),
    .I1(sig0000011b),
    .I2(sig000000e2),
    .I3(sig000000e2),
    .I4(sig00000005),
    .I5(sig0000000b),
    .O(sig000007d3)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk00000706 (
    .I0(sig00000142),
    .I1(sig0000011c),
    .I2(sig000000e3),
    .I3(sig000000e3),
    .I4(sig00000005),
    .I5(sig0000000b),
    .O(sig000007d4)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk00000707 (
    .I0(sig00000143),
    .I1(sig0000011d),
    .I2(sig000000e4),
    .I3(sig000000e4),
    .I4(sig00000005),
    .I5(sig0000000b),
    .O(sig000007d5)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk00000708 (
    .I0(sig00000144),
    .I1(sig0000011e),
    .I2(sig000000e5),
    .I3(sig000000e5),
    .I4(sig00000005),
    .I5(sig0000000b),
    .O(sig000007d6)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk00000709 (
    .I0(sig00000145),
    .I1(sig0000011f),
    .I2(sig000000e6),
    .I3(sig000000e6),
    .I4(sig00000005),
    .I5(sig0000000b),
    .O(sig000007d7)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk0000070a (
    .I0(sig00000146),
    .I1(sig00000120),
    .I2(sig000000e7),
    .I3(sig000000e7),
    .I4(sig00000005),
    .I5(sig0000000b),
    .O(sig000007d8)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk0000070b (
    .I0(sig00000147),
    .I1(sig00000121),
    .I2(sig000000e8),
    .I3(sig000000e8),
    .I4(sig00000005),
    .I5(sig0000000b),
    .O(sig000007d9)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk0000070c (
    .I0(sig00000148),
    .I1(sig00000122),
    .I2(sig000000e9),
    .I3(sig000000e9),
    .I4(sig00000005),
    .I5(sig0000000b),
    .O(sig000007da)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk0000070d (
    .I0(sig00000149),
    .I1(sig00000123),
    .I2(sig000000ea),
    .I3(sig000000ea),
    .I4(sig00000005),
    .I5(sig0000000b),
    .O(sig000007db)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk0000070e (
    .I0(sig0000014a),
    .I1(sig00000124),
    .I2(sig000000eb),
    .I3(sig000000eb),
    .I4(sig00000005),
    .I5(sig0000000b),
    .O(sig000007dc)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk0000070f (
    .I0(sig0000014b),
    .I1(sig00000125),
    .I2(sig000000ec),
    .I3(sig000000ec),
    .I4(sig00000005),
    .I5(sig0000000b),
    .O(sig000007dd)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk00000710 (
    .I0(sig0000014c),
    .I1(sig00000126),
    .I2(sig000000ed),
    .I3(sig000000ed),
    .I4(sig00000005),
    .I5(sig0000000b),
    .O(sig000007de)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000711 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000007cc),
    .R(sig00000002),
    .Q(sig000000b5)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000712 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000007cd),
    .R(sig00000002),
    .Q(sig000000b6)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000713 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000007ce),
    .R(sig00000002),
    .Q(sig000000b7)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000714 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000007cf),
    .R(sig00000002),
    .Q(sig000000b8)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000715 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000007d0),
    .R(sig00000002),
    .Q(sig000000b9)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000716 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000007d1),
    .R(sig00000002),
    .Q(sig000000ba)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000717 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000007d2),
    .R(sig00000002),
    .Q(sig000000bb)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000718 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000007d3),
    .R(sig00000002),
    .Q(sig000000bc)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000719 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000007d4),
    .R(sig00000002),
    .Q(sig000000bd)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000071a (
    .C(clk),
    .CE(sig00000001),
    .D(sig000007d5),
    .R(sig00000002),
    .Q(sig000000be)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000071b (
    .C(clk),
    .CE(sig00000001),
    .D(sig000007d6),
    .R(sig00000002),
    .Q(sig000000bf)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000071c (
    .C(clk),
    .CE(sig00000001),
    .D(sig000007d7),
    .R(sig00000002),
    .Q(sig000000c0)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000071d (
    .C(clk),
    .CE(sig00000001),
    .D(sig000007d8),
    .R(sig00000002),
    .Q(sig000000c1)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000071e (
    .C(clk),
    .CE(sig00000001),
    .D(sig000007d9),
    .R(sig00000002),
    .Q(sig000000c2)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000071f (
    .C(clk),
    .CE(sig00000001),
    .D(sig000007da),
    .R(sig00000002),
    .Q(sig000000c3)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000720 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000007db),
    .R(sig00000002),
    .Q(sig000000c4)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000721 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000007dc),
    .R(sig00000002),
    .Q(sig000000c5)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000722 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000007dd),
    .R(sig00000002),
    .Q(sig000000c6)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000723 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000007de),
    .R(sig00000002),
    .Q(sig000000c7)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk00000724 (
    .I0(sig00000127),
    .I1(sig00000101),
    .I2(sig000000ee),
    .I3(sig000000ee),
    .I4(sig00000005),
    .I5(sig0000000b),
    .O(sig000007df)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk00000725 (
    .I0(sig00000128),
    .I1(sig00000102),
    .I2(sig000000ef),
    .I3(sig000000ef),
    .I4(sig00000005),
    .I5(sig0000000b),
    .O(sig000007e0)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk00000726 (
    .I0(sig00000129),
    .I1(sig00000103),
    .I2(sig000000f0),
    .I3(sig000000f0),
    .I4(sig00000005),
    .I5(sig0000000b),
    .O(sig000007e1)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk00000727 (
    .I0(sig0000012a),
    .I1(sig00000104),
    .I2(sig000000f1),
    .I3(sig000000f1),
    .I4(sig00000005),
    .I5(sig0000000b),
    .O(sig000007e2)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk00000728 (
    .I0(sig0000012b),
    .I1(sig00000105),
    .I2(sig000000f2),
    .I3(sig000000f2),
    .I4(sig00000005),
    .I5(sig0000000b),
    .O(sig000007e3)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk00000729 (
    .I0(sig0000012c),
    .I1(sig00000106),
    .I2(sig000000f3),
    .I3(sig000000f3),
    .I4(sig00000005),
    .I5(sig0000000b),
    .O(sig000007e4)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk0000072a (
    .I0(sig0000012d),
    .I1(sig00000107),
    .I2(sig000000f4),
    .I3(sig000000f4),
    .I4(sig00000005),
    .I5(sig0000000b),
    .O(sig000007e5)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk0000072b (
    .I0(sig0000012e),
    .I1(sig00000108),
    .I2(sig000000f5),
    .I3(sig000000f5),
    .I4(sig00000005),
    .I5(sig0000000b),
    .O(sig000007e6)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk0000072c (
    .I0(sig0000012f),
    .I1(sig00000109),
    .I2(sig000000f6),
    .I3(sig000000f6),
    .I4(sig00000005),
    .I5(sig0000000b),
    .O(sig000007e7)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk0000072d (
    .I0(sig00000130),
    .I1(sig0000010a),
    .I2(sig000000f7),
    .I3(sig000000f7),
    .I4(sig00000005),
    .I5(sig0000000b),
    .O(sig000007e8)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk0000072e (
    .I0(sig00000131),
    .I1(sig0000010b),
    .I2(sig000000f8),
    .I3(sig000000f8),
    .I4(sig00000005),
    .I5(sig0000000b),
    .O(sig000007e9)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk0000072f (
    .I0(sig00000132),
    .I1(sig0000010c),
    .I2(sig000000f9),
    .I3(sig000000f9),
    .I4(sig00000005),
    .I5(sig0000000b),
    .O(sig000007ea)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk00000730 (
    .I0(sig00000133),
    .I1(sig0000010d),
    .I2(sig000000fa),
    .I3(sig000000fa),
    .I4(sig00000005),
    .I5(sig0000000b),
    .O(sig000007eb)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk00000731 (
    .I0(sig00000134),
    .I1(sig0000010e),
    .I2(sig000000fb),
    .I3(sig000000fb),
    .I4(sig00000005),
    .I5(sig0000000b),
    .O(sig000007ec)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk00000732 (
    .I0(sig00000135),
    .I1(sig0000010f),
    .I2(sig000000fc),
    .I3(sig000000fc),
    .I4(sig00000005),
    .I5(sig0000000b),
    .O(sig000007ed)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk00000733 (
    .I0(sig00000136),
    .I1(sig00000110),
    .I2(sig000000fd),
    .I3(sig000000fd),
    .I4(sig00000005),
    .I5(sig0000000b),
    .O(sig000007ee)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk00000734 (
    .I0(sig00000137),
    .I1(sig00000111),
    .I2(sig000000fe),
    .I3(sig000000fe),
    .I4(sig00000005),
    .I5(sig0000000b),
    .O(sig000007ef)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk00000735 (
    .I0(sig00000138),
    .I1(sig00000112),
    .I2(sig000000ff),
    .I3(sig000000ff),
    .I4(sig00000005),
    .I5(sig0000000b),
    .O(sig000007f0)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk00000736 (
    .I0(sig00000139),
    .I1(sig00000113),
    .I2(sig00000100),
    .I3(sig00000100),
    .I4(sig00000005),
    .I5(sig0000000b),
    .O(sig000007f1)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000737 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000007df),
    .R(sig00000002),
    .Q(sig000000c8)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000738 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000007e0),
    .R(sig00000002),
    .Q(sig000000c9)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000739 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000007e1),
    .R(sig00000002),
    .Q(sig000000ca)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000073a (
    .C(clk),
    .CE(sig00000001),
    .D(sig000007e2),
    .R(sig00000002),
    .Q(sig000000cb)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000073b (
    .C(clk),
    .CE(sig00000001),
    .D(sig000007e3),
    .R(sig00000002),
    .Q(sig000000cc)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000073c (
    .C(clk),
    .CE(sig00000001),
    .D(sig000007e4),
    .R(sig00000002),
    .Q(sig000000cd)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000073d (
    .C(clk),
    .CE(sig00000001),
    .D(sig000007e5),
    .R(sig00000002),
    .Q(sig000000ce)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000073e (
    .C(clk),
    .CE(sig00000001),
    .D(sig000007e6),
    .R(sig00000002),
    .Q(sig000000cf)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000073f (
    .C(clk),
    .CE(sig00000001),
    .D(sig000007e7),
    .R(sig00000002),
    .Q(sig000000d0)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000740 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000007e8),
    .R(sig00000002),
    .Q(sig000000d1)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000741 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000007e9),
    .R(sig00000002),
    .Q(sig000000d2)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000742 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000007ea),
    .R(sig00000002),
    .Q(sig000000d3)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000743 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000007eb),
    .R(sig00000002),
    .Q(sig000000d4)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000744 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000007ec),
    .R(sig00000002),
    .Q(sig000000d5)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000745 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000007ed),
    .R(sig00000002),
    .Q(sig000000d6)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000746 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000007ee),
    .R(sig00000002),
    .Q(sig000000d7)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000747 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000007ef),
    .R(sig00000002),
    .Q(sig000000d8)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000748 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000007f0),
    .R(sig00000002),
    .Q(sig000000d9)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000749 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000007f1),
    .R(sig00000002),
    .Q(sig000000da)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk0000074a (
    .A0(sig00000001),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig0000080f),
    .Q(sig000007f2)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000074b (
    .C(clk),
    .CE(sig00000001),
    .D(sig000007f2),
    .R(sig00000002),
    .Q(sig0000000c)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000074c (
    .C(clk),
    .D(sig000007f9),
    .Q(sig00000824)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000074d (
    .C(clk),
    .CE(sig00000001),
    .D(sig000007f3),
    .Q(sig0000080f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000074e (
    .C(clk),
    .CE(sig00000001),
    .D(sig000007f7),
    .Q(sig000007f6)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000074f (
    .C(clk),
    .D(sig000007f5),
    .Q(sig0000000a)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000750 (
    .C(clk),
    .D(sig000007f4),
    .Q(sig00000009)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000075d (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000859),
    .Q(sig00000850)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000075e (
    .C(clk),
    .D(sig0000084f),
    .Q(sig00000861)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000075f (
    .C(clk),
    .D(sig0000084e),
    .Q(sig00000860)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000760 (
    .C(clk),
    .D(sig0000084d),
    .Q(sig0000085f)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000761 (
    .C(clk),
    .D(sig0000084c),
    .Q(sig0000085e)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000762 (
    .C(clk),
    .D(sig0000084b),
    .Q(sig0000085d)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000763 (
    .C(clk),
    .D(sig0000084a),
    .Q(sig0000085c)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000764 (
    .C(clk),
    .D(sig00000849),
    .Q(sig0000085b)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000765 (
    .C(clk),
    .D(sig00000848),
    .Q(sig0000085a)
  );
  MUXF8   blk00000766 (
    .I0(sig0000086c),
    .I1(sig0000086b),
    .S(sig00000001),
    .O(sig00000863)
  );
  MUXF8   blk00000767 (
    .I0(sig0000086e),
    .I1(sig0000086d),
    .S(sig00000001),
    .O(sig00000864)
  );
  MUXF8   blk00000768 (
    .I0(sig00000870),
    .I1(sig0000086f),
    .S(sig00000001),
    .O(sig00000865)
  );
  MUXF8   blk00000769 (
    .I0(sig00000872),
    .I1(sig00000871),
    .S(sig00000001),
    .O(sig00000866)
  );
  MUXF8   blk0000076a (
    .I0(sig00000874),
    .I1(sig00000873),
    .S(sig00000001),
    .O(sig00000867)
  );
  MUXF8   blk0000076b (
    .I0(sig00000876),
    .I1(sig00000875),
    .S(sig00000001),
    .O(sig00000868)
  );
  MUXF8   blk0000076c (
    .I0(sig00000878),
    .I1(sig00000877),
    .S(sig00000001),
    .O(sig00000869)
  );
  MUXF8   blk0000076d (
    .I0(sig0000087a),
    .I1(sig00000879),
    .S(sig00000001),
    .O(sig0000086a)
  );
  MUXF7   blk0000076e (
    .I0(sig00000883),
    .I1(sig0000087b),
    .S(sig00000002),
    .O(sig0000086b)
  );
  MUXF7   blk0000076f (
    .I0(sig00000893),
    .I1(sig0000088b),
    .S(sig00000002),
    .O(sig0000086c)
  );
  MUXF7   blk00000770 (
    .I0(sig00000884),
    .I1(sig0000087c),
    .S(sig00000002),
    .O(sig0000086d)
  );
  MUXF7   blk00000771 (
    .I0(sig00000894),
    .I1(sig0000088c),
    .S(sig00000002),
    .O(sig0000086e)
  );
  MUXF7   blk00000772 (
    .I0(sig00000885),
    .I1(sig0000087d),
    .S(sig00000002),
    .O(sig0000086f)
  );
  MUXF7   blk00000773 (
    .I0(sig00000895),
    .I1(sig0000088d),
    .S(sig00000002),
    .O(sig00000870)
  );
  MUXF7   blk00000774 (
    .I0(sig00000886),
    .I1(sig0000087e),
    .S(sig00000002),
    .O(sig00000871)
  );
  MUXF7   blk00000775 (
    .I0(sig00000896),
    .I1(sig0000088e),
    .S(sig00000002),
    .O(sig00000872)
  );
  MUXF7   blk00000776 (
    .I0(sig00000887),
    .I1(sig0000087f),
    .S(sig00000002),
    .O(sig00000873)
  );
  MUXF7   blk00000777 (
    .I0(sig00000897),
    .I1(sig0000088f),
    .S(sig00000002),
    .O(sig00000874)
  );
  MUXF7   blk00000778 (
    .I0(sig00000888),
    .I1(sig00000880),
    .S(sig00000002),
    .O(sig00000875)
  );
  MUXF7   blk00000779 (
    .I0(sig00000898),
    .I1(sig00000890),
    .S(sig00000002),
    .O(sig00000876)
  );
  MUXF7   blk0000077a (
    .I0(sig00000889),
    .I1(sig00000881),
    .S(sig00000002),
    .O(sig00000877)
  );
  MUXF7   blk0000077b (
    .I0(sig00000899),
    .I1(sig00000891),
    .S(sig00000002),
    .O(sig00000878)
  );
  MUXF7   blk0000077c (
    .I0(sig0000088a),
    .I1(sig00000882),
    .S(sig00000002),
    .O(sig00000879)
  );
  MUXF7   blk0000077d (
    .I0(sig0000089a),
    .I1(sig00000892),
    .S(sig00000002),
    .O(sig0000087a)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk0000077e (
    .I0(sig00000002),
    .I1(sig00000002),
    .I2(sig00000002),
    .I3(sig00000002),
    .I4(sig00000001),
    .I5(sig00000002),
    .O(sig0000087b)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk0000077f (
    .I0(sig00000002),
    .I1(sig00000002),
    .I2(sig00000002),
    .I3(sig00000002),
    .I4(sig00000001),
    .I5(sig00000002),
    .O(sig0000087c)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk00000780 (
    .I0(sig00000002),
    .I1(sig00000002),
    .I2(sig00000002),
    .I3(sig00000002),
    .I4(sig00000001),
    .I5(sig00000002),
    .O(sig0000087d)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk00000781 (
    .I0(sig0000084f),
    .I1(sig00000002),
    .I2(sig00000002),
    .I3(sig00000002),
    .I4(sig00000001),
    .I5(sig00000002),
    .O(sig0000087e)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk00000782 (
    .I0(sig0000084e),
    .I1(sig0000084f),
    .I2(sig00000002),
    .I3(sig00000002),
    .I4(sig00000001),
    .I5(sig00000002),
    .O(sig0000087f)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk00000783 (
    .I0(sig0000084d),
    .I1(sig0000084e),
    .I2(sig0000084f),
    .I3(sig00000002),
    .I4(sig00000001),
    .I5(sig00000002),
    .O(sig00000880)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk00000784 (
    .I0(sig0000084c),
    .I1(sig0000084d),
    .I2(sig0000084e),
    .I3(sig0000084f),
    .I4(sig00000001),
    .I5(sig00000002),
    .O(sig00000881)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk00000785 (
    .I0(sig0000084b),
    .I1(sig0000084c),
    .I2(sig0000084d),
    .I3(sig0000084e),
    .I4(sig00000001),
    .I5(sig00000002),
    .O(sig00000882)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk00000786 (
    .I0(sig0000084e),
    .I1(sig0000084f),
    .I2(sig00000002),
    .I3(sig00000002),
    .I4(sig00000001),
    .I5(sig00000002),
    .O(sig00000883)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk00000787 (
    .I0(sig0000084d),
    .I1(sig0000084e),
    .I2(sig0000084f),
    .I3(sig00000002),
    .I4(sig00000001),
    .I5(sig00000002),
    .O(sig00000884)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk00000788 (
    .I0(sig0000084c),
    .I1(sig0000084d),
    .I2(sig0000084e),
    .I3(sig0000084f),
    .I4(sig00000001),
    .I5(sig00000002),
    .O(sig00000885)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk00000789 (
    .I0(sig0000084b),
    .I1(sig0000084c),
    .I2(sig0000084d),
    .I3(sig0000084e),
    .I4(sig00000001),
    .I5(sig00000002),
    .O(sig00000886)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk0000078a (
    .I0(sig0000084a),
    .I1(sig0000084b),
    .I2(sig0000084c),
    .I3(sig0000084d),
    .I4(sig00000001),
    .I5(sig00000002),
    .O(sig00000887)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk0000078b (
    .I0(sig00000849),
    .I1(sig0000084a),
    .I2(sig0000084b),
    .I3(sig0000084c),
    .I4(sig00000001),
    .I5(sig00000002),
    .O(sig00000888)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk0000078c (
    .I0(sig00000848),
    .I1(sig00000849),
    .I2(sig0000084a),
    .I3(sig0000084b),
    .I4(sig00000001),
    .I5(sig00000002),
    .O(sig00000889)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk0000078d (
    .I0(sig00000002),
    .I1(sig00000848),
    .I2(sig00000849),
    .I3(sig0000084a),
    .I4(sig00000001),
    .I5(sig00000002),
    .O(sig0000088a)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk0000078e (
    .I0(sig0000084a),
    .I1(sig0000084b),
    .I2(sig0000084c),
    .I3(sig0000084d),
    .I4(sig00000001),
    .I5(sig00000002),
    .O(sig0000088b)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk0000078f (
    .I0(sig00000849),
    .I1(sig0000084a),
    .I2(sig0000084b),
    .I3(sig0000084c),
    .I4(sig00000001),
    .I5(sig00000002),
    .O(sig0000088c)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk00000790 (
    .I0(sig00000848),
    .I1(sig00000849),
    .I2(sig0000084a),
    .I3(sig0000084b),
    .I4(sig00000001),
    .I5(sig00000002),
    .O(sig0000088d)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk00000791 (
    .I0(sig00000002),
    .I1(sig00000848),
    .I2(sig00000849),
    .I3(sig0000084a),
    .I4(sig00000001),
    .I5(sig00000002),
    .O(sig0000088e)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk00000792 (
    .I0(sig00000002),
    .I1(sig00000002),
    .I2(sig00000848),
    .I3(sig00000849),
    .I4(sig00000001),
    .I5(sig00000002),
    .O(sig0000088f)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk00000793 (
    .I0(sig00000002),
    .I1(sig00000002),
    .I2(sig00000002),
    .I3(sig00000848),
    .I4(sig00000001),
    .I5(sig00000002),
    .O(sig00000890)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk00000794 (
    .I0(sig00000002),
    .I1(sig00000002),
    .I2(sig00000002),
    .I3(sig00000002),
    .I4(sig00000001),
    .I5(sig00000002),
    .O(sig00000891)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk00000795 (
    .I0(sig00000002),
    .I1(sig00000002),
    .I2(sig00000002),
    .I3(sig00000002),
    .I4(sig00000001),
    .I5(sig00000002),
    .O(sig00000892)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk00000796 (
    .I0(sig00000002),
    .I1(sig00000002),
    .I2(sig00000002),
    .I3(sig00000849),
    .I4(sig00000001),
    .I5(sig00000002),
    .O(sig00000893)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk00000797 (
    .I0(sig00000002),
    .I1(sig00000002),
    .I2(sig00000002),
    .I3(sig00000848),
    .I4(sig00000001),
    .I5(sig00000002),
    .O(sig00000894)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk00000798 (
    .I0(sig00000002),
    .I1(sig00000002),
    .I2(sig00000002),
    .I3(sig00000002),
    .I4(sig00000001),
    .I5(sig00000002),
    .O(sig00000895)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk00000799 (
    .I0(sig00000002),
    .I1(sig00000002),
    .I2(sig00000002),
    .I3(sig00000002),
    .I4(sig00000001),
    .I5(sig00000002),
    .O(sig00000896)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk0000079a (
    .I0(sig00000002),
    .I1(sig00000002),
    .I2(sig00000002),
    .I3(sig00000002),
    .I4(sig00000001),
    .I5(sig00000002),
    .O(sig00000897)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk0000079b (
    .I0(sig00000002),
    .I1(sig00000002),
    .I2(sig00000002),
    .I3(sig00000002),
    .I4(sig00000001),
    .I5(sig00000002),
    .O(sig00000898)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk0000079c (
    .I0(sig00000002),
    .I1(sig00000002),
    .I2(sig00000002),
    .I3(sig00000002),
    .I4(sig00000001),
    .I5(sig00000002),
    .O(sig00000899)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk0000079d (
    .I0(sig00000002),
    .I1(sig00000002),
    .I2(sig00000002),
    .I3(sig00000002),
    .I4(sig00000001),
    .I5(sig00000002),
    .O(sig0000089a)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000079e (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000089b),
    .R(sig00000002),
    .Q(sig00000851)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000079f (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000863),
    .R(sig00000002),
    .Q(sig0000089b)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000007a0 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000089c),
    .R(sig00000002),
    .Q(sig00000852)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000007a1 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000864),
    .R(sig00000002),
    .Q(sig0000089c)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000007a2 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000089d),
    .R(sig00000002),
    .Q(sig00000853)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000007a3 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000865),
    .R(sig00000002),
    .Q(sig0000089d)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000007a4 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000089e),
    .R(sig00000002),
    .Q(sig00000854)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000007a5 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000866),
    .R(sig00000002),
    .Q(sig0000089e)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000007a6 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000089f),
    .R(sig00000002),
    .Q(sig00000855)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000007a7 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000867),
    .R(sig00000002),
    .Q(sig0000089f)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000007a8 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000008a0),
    .R(sig00000002),
    .Q(sig00000856)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000007a9 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000868),
    .R(sig00000002),
    .Q(sig000008a0)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000007aa (
    .C(clk),
    .CE(sig00000001),
    .D(sig000008a1),
    .R(sig00000002),
    .Q(sig00000857)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000007ab (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000869),
    .R(sig00000002),
    .Q(sig000008a1)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000007ac (
    .C(clk),
    .CE(sig00000001),
    .D(sig000008a2),
    .R(sig00000002),
    .Q(sig00000858)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000007ad (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000086a),
    .R(sig00000002),
    .Q(sig000008a2)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000007ae (
    .C(clk),
    .D(NlwRenamedSig_OI_xn_index[7]),
    .Q(sig0000084f)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000007af (
    .C(clk),
    .D(NlwRenamedSig_OI_xn_index[6]),
    .Q(sig0000084e)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000007b0 (
    .C(clk),
    .D(NlwRenamedSig_OI_xn_index[5]),
    .Q(sig0000084d)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000007b1 (
    .C(clk),
    .D(NlwRenamedSig_OI_xn_index[4]),
    .Q(sig0000084c)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000007b2 (
    .C(clk),
    .D(NlwRenamedSig_OI_xn_index[3]),
    .Q(sig0000084b)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000007b3 (
    .C(clk),
    .D(NlwRenamedSig_OI_xn_index[2]),
    .Q(sig0000084a)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000007b4 (
    .C(clk),
    .D(NlwRenamedSig_OI_xn_index[1]),
    .Q(sig00000849)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000007b5 (
    .C(clk),
    .D(NlwRenamedSig_OI_xn_index[0]),
    .Q(sig00000848)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000007b6 (
    .I0(sig000008cd),
    .I1(sig00000002),
    .I2(sig000008cf),
    .I3(sig000008ce),
    .I4(sig000008c4),
    .I5(sig000008c5),
    .O(sig000008a4)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000007b7 (
    .I0(sig000008cc),
    .I1(sig00000002),
    .I2(sig000008cf),
    .I3(sig000008cd),
    .I4(sig000008c5),
    .I5(sig000008c2),
    .O(sig000008a5)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000007b8 (
    .I0(sig000008cb),
    .I1(sig00000002),
    .I2(sig000008cf),
    .I3(sig000008cc),
    .I4(sig000008c2),
    .I5(sig000008c3),
    .O(sig000008a6)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000007b9 (
    .I0(sig000008ca),
    .I1(sig00000002),
    .I2(sig000008cf),
    .I3(sig000008cb),
    .I4(sig000008c3),
    .I5(sig000008c0),
    .O(sig000008a7)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000007ba (
    .I0(sig000008c9),
    .I1(sig00000002),
    .I2(sig000008cf),
    .I3(sig000008ca),
    .I4(sig000008c0),
    .I5(sig000008c1),
    .O(sig000008a8)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000007bb (
    .I0(sig000008c8),
    .I1(sig00000002),
    .I2(sig000008cf),
    .I3(sig000008c9),
    .I4(sig000008c1),
    .I5(sig000008be),
    .O(sig000008a9)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000007bc (
    .I0(sig000008c7),
    .I1(sig00000002),
    .I2(sig000008cf),
    .I3(sig000008c8),
    .I4(sig000008be),
    .I5(sig000008bf),
    .O(sig000008aa)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000007bd (
    .I0(sig00000002),
    .I1(sig00000002),
    .I2(sig000008cf),
    .I3(sig000008c7),
    .I4(sig000008bf),
    .I5(sig000008c6),
    .O(sig000008ab)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000007be (
    .I0(sig000008cd),
    .I1(sig00000002),
    .I2(sig000008bc),
    .I3(sig000008ce),
    .I4(sig000008c4),
    .I5(sig000008c5),
    .O(sig000008ac)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000007bf (
    .I0(sig000008cc),
    .I1(sig00000002),
    .I2(sig000008bc),
    .I3(sig000008cd),
    .I4(sig000008c5),
    .I5(sig000008c2),
    .O(sig000008ad)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000007c0 (
    .I0(sig000008cb),
    .I1(sig00000002),
    .I2(sig000008bc),
    .I3(sig000008cc),
    .I4(sig000008c2),
    .I5(sig000008c3),
    .O(sig000008ae)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000007c1 (
    .I0(sig000008ca),
    .I1(sig00000002),
    .I2(sig000008bc),
    .I3(sig000008cb),
    .I4(sig000008c3),
    .I5(sig000008c0),
    .O(sig000008af)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000007c2 (
    .I0(sig000008c9),
    .I1(sig00000002),
    .I2(sig000008bc),
    .I3(sig000008ca),
    .I4(sig000008c0),
    .I5(sig000008c1),
    .O(sig000008b0)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000007c3 (
    .I0(sig000008c8),
    .I1(sig00000002),
    .I2(sig000008bc),
    .I3(sig000008c9),
    .I4(sig000008c1),
    .I5(sig000008be),
    .O(sig000008b1)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000007c4 (
    .I0(sig000008c7),
    .I1(sig00000002),
    .I2(sig000008bc),
    .I3(sig000008c8),
    .I4(sig000008be),
    .I5(sig000008bf),
    .O(sig000008b2)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000007c5 (
    .I0(sig00000002),
    .I1(sig00000002),
    .I2(sig000008bc),
    .I3(sig000008c7),
    .I4(sig000008bf),
    .I5(sig000008c6),
    .O(sig000008b3)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000007c6 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000008a4),
    .R(sig00000002),
    .Q(sig00000840)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000007c7 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000008a5),
    .R(sig00000002),
    .Q(sig00000841)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000007c8 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000008a6),
    .R(sig00000002),
    .Q(sig00000842)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000007c9 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000008a7),
    .R(sig00000002),
    .Q(sig00000843)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000007ca (
    .C(clk),
    .CE(sig00000001),
    .D(sig000008a8),
    .R(sig00000002),
    .Q(sig00000844)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000007cb (
    .C(clk),
    .CE(sig00000001),
    .D(sig000008a9),
    .R(sig00000002),
    .Q(sig00000845)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000007cc (
    .C(clk),
    .CE(sig00000001),
    .D(sig000008aa),
    .R(sig00000002),
    .Q(sig00000846)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000007cd (
    .C(clk),
    .CE(sig00000001),
    .D(sig000008ab),
    .R(sig00000002),
    .Q(sig00000847)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000007ce (
    .C(clk),
    .CE(sig00000001),
    .D(sig000008ac),
    .R(sig00000002),
    .Q(sig00000838)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000007cf (
    .C(clk),
    .CE(sig00000001),
    .D(sig000008ad),
    .R(sig00000002),
    .Q(sig00000839)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000007d0 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000008ae),
    .R(sig00000002),
    .Q(sig0000083a)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000007d1 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000008af),
    .R(sig00000002),
    .Q(sig0000083b)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000007d2 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000008b0),
    .R(sig00000002),
    .Q(sig0000083c)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000007d3 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000008b1),
    .R(sig00000002),
    .Q(sig0000083d)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000007d4 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000008b2),
    .R(sig00000002),
    .Q(sig0000083e)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000007d5 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000008b3),
    .R(sig00000002),
    .Q(sig0000083f)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000007d6 (
    .C(clk),
    .D(sig000008b4),
    .Q(sig000008cf)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000007d7 (
    .C(clk),
    .D(sig000008cf),
    .Q(sig00000837)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000007d8 (
    .C(clk),
    .D(sig000008b9),
    .Q(sig000008c1)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000007d9 (
    .C(clk),
    .D(sig000008ba),
    .Q(sig000008c0)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000007da (
    .C(clk),
    .D(sig000008bb),
    .Q(sig000008c3)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000007db (
    .C(clk),
    .D(sig000008b5),
    .Q(sig000008c2)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000007dc (
    .C(clk),
    .D(sig000008bd),
    .Q(sig000008bf)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000007dd (
    .C(clk),
    .D(sig000008b8),
    .Q(sig000008be)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000007de (
    .C(clk),
    .D(sig000008bc),
    .Q(sig00000836)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000007df (
    .C(clk),
    .D(sig000008a3),
    .Q(sig000008c5)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000007e0 (
    .C(clk),
    .D(sig000008b6),
    .Q(sig000008c4)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000007e1 (
    .C(clk),
    .D(sig000008b7),
    .Q(sig000008c6)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000007e2 (
    .C(clk),
    .D(sig0000080e),
    .Q(sig000008c7)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000007e3 (
    .C(clk),
    .D(sig0000080d),
    .Q(sig000008c8)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000007e4 (
    .C(clk),
    .D(sig0000080c),
    .Q(sig000008c9)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000007e5 (
    .C(clk),
    .D(sig0000080b),
    .Q(sig000008ca)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000007e6 (
    .C(clk),
    .D(sig0000080a),
    .Q(sig000008cb)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000007e7 (
    .C(clk),
    .D(sig00000809),
    .Q(sig000008cc)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000007e8 (
    .C(clk),
    .D(sig00000808),
    .Q(sig000008cd)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk000007e9 (
    .C(clk),
    .D(sig00000807),
    .Q(sig000008ce)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000812 (
    .I0(sig0000083f),
    .I1(sig00000802),
    .I2(sig00000824),
    .O(sig000008d0)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000813 (
    .I0(sig0000083e),
    .I1(sig00000801),
    .I2(sig00000824),
    .O(sig000008d1)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000814 (
    .I0(sig0000083d),
    .I1(sig00000800),
    .I2(sig00000824),
    .O(sig000008d2)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000815 (
    .I0(sig0000083c),
    .I1(sig000007ff),
    .I2(sig00000824),
    .O(sig000008d3)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000816 (
    .I0(sig0000083b),
    .I1(sig000007fe),
    .I2(sig00000824),
    .O(sig000008d4)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000817 (
    .I0(sig0000083a),
    .I1(sig000007fd),
    .I2(sig00000824),
    .O(sig000008d5)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000818 (
    .I0(sig00000839),
    .I1(sig000007fc),
    .I2(sig00000824),
    .O(sig000008d6)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000819 (
    .I0(sig00000838),
    .I1(sig000007fb),
    .I2(sig00000824),
    .O(sig000008d7)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000081a (
    .C(clk),
    .CE(sig00000001),
    .D(sig000008d0),
    .R(sig00000002),
    .Q(sig00000028)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000081b (
    .C(clk),
    .CE(sig00000001),
    .D(sig000008d1),
    .R(sig00000002),
    .Q(sig00000027)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000081c (
    .C(clk),
    .CE(sig00000001),
    .D(sig000008d2),
    .R(sig00000002),
    .Q(sig00000026)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000081d (
    .C(clk),
    .CE(sig00000001),
    .D(sig000008d3),
    .R(sig00000002),
    .Q(sig00000025)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000081e (
    .C(clk),
    .CE(sig00000001),
    .D(sig000008d4),
    .R(sig00000002),
    .Q(sig00000024)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000081f (
    .C(clk),
    .CE(sig00000001),
    .D(sig000008d5),
    .R(sig00000002),
    .Q(sig00000023)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000820 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000008d6),
    .R(sig00000002),
    .Q(sig00000022)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000821 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000008d7),
    .R(sig00000002),
    .Q(sig00000021)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000822 (
    .I0(sig00000847),
    .I1(sig00000802),
    .I2(sig00000824),
    .O(sig000008d8)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000823 (
    .I0(sig00000846),
    .I1(sig00000801),
    .I2(sig00000824),
    .O(sig000008d9)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000824 (
    .I0(sig00000845),
    .I1(sig00000800),
    .I2(sig00000824),
    .O(sig000008da)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000825 (
    .I0(sig00000844),
    .I1(sig000007ff),
    .I2(sig00000824),
    .O(sig000008db)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000826 (
    .I0(sig00000843),
    .I1(sig000007fe),
    .I2(sig00000824),
    .O(sig000008dc)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000827 (
    .I0(sig00000842),
    .I1(sig000007fd),
    .I2(sig00000824),
    .O(sig000008dd)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000828 (
    .I0(sig00000841),
    .I1(sig000007fc),
    .I2(sig00000824),
    .O(sig000008de)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000829 (
    .I0(sig00000840),
    .I1(sig000007fb),
    .I2(sig00000824),
    .O(sig000008df)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000082a (
    .C(clk),
    .CE(sig00000001),
    .D(sig000008d8),
    .R(sig00000002),
    .Q(sig00000038)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000082b (
    .C(clk),
    .CE(sig00000001),
    .D(sig000008d9),
    .R(sig00000002),
    .Q(sig00000037)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000082c (
    .C(clk),
    .CE(sig00000001),
    .D(sig000008da),
    .R(sig00000002),
    .Q(sig00000036)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000082d (
    .C(clk),
    .CE(sig00000001),
    .D(sig000008db),
    .R(sig00000002),
    .Q(sig00000035)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000082e (
    .C(clk),
    .CE(sig00000001),
    .D(sig000008dc),
    .R(sig00000002),
    .Q(sig00000034)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000082f (
    .C(clk),
    .CE(sig00000001),
    .D(sig000008dd),
    .R(sig00000002),
    .Q(sig00000033)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000830 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000008de),
    .R(sig00000002),
    .Q(sig00000032)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000831 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000008df),
    .R(sig00000002),
    .Q(sig00000031)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000832 (
    .I0(sig0000082d),
    .I1(sig00000858),
    .I2(sig0000000b),
    .O(sig000008e0)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000833 (
    .I0(sig0000082c),
    .I1(sig00000857),
    .I2(sig0000000b),
    .O(sig000008e1)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000834 (
    .I0(sig0000082b),
    .I1(sig00000856),
    .I2(sig0000000b),
    .O(sig000008e2)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000835 (
    .I0(sig0000082a),
    .I1(sig00000855),
    .I2(sig0000000b),
    .O(sig000008e3)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000836 (
    .I0(sig00000829),
    .I1(sig00000854),
    .I2(sig0000000b),
    .O(sig000008e4)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000837 (
    .I0(sig00000828),
    .I1(sig00000853),
    .I2(sig0000000b),
    .O(sig000008e5)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000838 (
    .I0(sig00000827),
    .I1(sig00000852),
    .I2(sig0000000b),
    .O(sig000008e6)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000839 (
    .I0(sig00000826),
    .I1(sig00000851),
    .I2(sig0000000b),
    .O(sig000008e7)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000083a (
    .C(clk),
    .CE(sig00000001),
    .D(sig000008e0),
    .R(sig00000002),
    .Q(sig00000030)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000083b (
    .C(clk),
    .CE(sig00000001),
    .D(sig000008e1),
    .R(sig00000002),
    .Q(sig0000002f)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000083c (
    .C(clk),
    .CE(sig00000001),
    .D(sig000008e2),
    .R(sig00000002),
    .Q(sig0000002e)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000083d (
    .C(clk),
    .CE(sig00000001),
    .D(sig000008e3),
    .R(sig00000002),
    .Q(sig0000002d)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000083e (
    .C(clk),
    .CE(sig00000001),
    .D(sig000008e4),
    .R(sig00000002),
    .Q(sig0000002c)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000083f (
    .C(clk),
    .CE(sig00000001),
    .D(sig000008e5),
    .R(sig00000002),
    .Q(sig0000002b)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000840 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000008e6),
    .R(sig00000002),
    .Q(sig0000002a)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000841 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000008e7),
    .R(sig00000002),
    .Q(sig00000029)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000842 (
    .I0(sig00000835),
    .I1(sig00000858),
    .I2(sig0000000b),
    .O(sig000008e8)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000843 (
    .I0(sig00000834),
    .I1(sig00000857),
    .I2(sig0000000b),
    .O(sig000008e9)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000844 (
    .I0(sig00000833),
    .I1(sig00000856),
    .I2(sig0000000b),
    .O(sig000008ea)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000845 (
    .I0(sig00000832),
    .I1(sig00000855),
    .I2(sig0000000b),
    .O(sig000008eb)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000846 (
    .I0(sig00000831),
    .I1(sig00000854),
    .I2(sig0000000b),
    .O(sig000008ec)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000847 (
    .I0(sig00000830),
    .I1(sig00000853),
    .I2(sig0000000b),
    .O(sig000008ed)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000848 (
    .I0(sig0000082f),
    .I1(sig00000852),
    .I2(sig0000000b),
    .O(sig000008ee)
  );
  LUT3 #(
    .INIT ( 8'hCA ))
  blk00000849 (
    .I0(sig0000082e),
    .I1(sig00000851),
    .I2(sig0000000b),
    .O(sig000008ef)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000084a (
    .C(clk),
    .CE(sig00000001),
    .D(sig000008e8),
    .R(sig00000002),
    .Q(sig00000040)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000084b (
    .C(clk),
    .CE(sig00000001),
    .D(sig000008e9),
    .R(sig00000002),
    .Q(sig0000003f)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000084c (
    .C(clk),
    .CE(sig00000001),
    .D(sig000008ea),
    .R(sig00000002),
    .Q(sig0000003e)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000084d (
    .C(clk),
    .CE(sig00000001),
    .D(sig000008eb),
    .R(sig00000002),
    .Q(sig0000003d)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000084e (
    .C(clk),
    .CE(sig00000001),
    .D(sig000008ec),
    .R(sig00000002),
    .Q(sig0000003c)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000084f (
    .C(clk),
    .CE(sig00000001),
    .D(sig000008ed),
    .R(sig00000002),
    .Q(sig0000003b)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000850 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000008ee),
    .R(sig00000002),
    .Q(sig0000003a)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000851 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000008ef),
    .R(sig00000002),
    .Q(sig00000039)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000864 (
    .C(clk),
    .D(sig000008f9),
    .Q(sig00000016)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000865 (
    .C(clk),
    .D(sig000008f8),
    .Q(sig00000015)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000866 (
    .C(clk),
    .D(sig000008f7),
    .Q(sig00000014)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000867 (
    .C(clk),
    .D(sig000008f6),
    .Q(sig00000013)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000868 (
    .C(clk),
    .D(sig000008f5),
    .Q(sig00000012)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000869 (
    .C(clk),
    .D(sig000008f4),
    .Q(sig00000011)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000086a (
    .C(clk),
    .D(sig000008f3),
    .Q(sig00000010)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000086b (
    .C(clk),
    .D(sig000008f2),
    .Q(sig0000000f)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000086c (
    .C(clk),
    .D(sig000008f1),
    .Q(sig0000000e)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000086d (
    .C(clk),
    .D(sig000008f0),
    .Q(sig0000000d)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000086e (
    .C(clk),
    .D(sig00000903),
    .Q(sig00000020)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000086f (
    .C(clk),
    .D(sig00000902),
    .Q(sig0000001f)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000870 (
    .C(clk),
    .D(sig00000901),
    .Q(sig0000001e)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000871 (
    .C(clk),
    .D(sig00000900),
    .Q(sig0000001d)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000872 (
    .C(clk),
    .D(sig000008ff),
    .Q(sig0000001c)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000873 (
    .C(clk),
    .D(sig000008fe),
    .Q(sig0000001b)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000874 (
    .C(clk),
    .D(sig000008fd),
    .Q(sig0000001a)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000875 (
    .C(clk),
    .D(sig000008fc),
    .Q(sig00000019)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000876 (
    .C(clk),
    .D(sig000008fb),
    .Q(sig00000018)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000877 (
    .C(clk),
    .D(sig000008fa),
    .Q(sig00000017)
  );
  MUXF8   blk00000878 (
    .I0(sig0000090e),
    .I1(sig0000090d),
    .S(sig00000813),
    .O(sig00000904)
  );
  MUXF8   blk00000879 (
    .I0(sig00000910),
    .I1(sig0000090f),
    .S(sig00000813),
    .O(sig00000905)
  );
  MUXF8   blk0000087a (
    .I0(sig00000912),
    .I1(sig00000911),
    .S(sig00000813),
    .O(sig00000906)
  );
  MUXF8   blk0000087b (
    .I0(sig00000914),
    .I1(sig00000913),
    .S(sig00000813),
    .O(sig00000907)
  );
  MUXF8   blk0000087c (
    .I0(sig00000916),
    .I1(sig00000915),
    .S(sig00000813),
    .O(sig00000908)
  );
  MUXF8   blk0000087d (
    .I0(sig00000918),
    .I1(sig00000917),
    .S(sig00000813),
    .O(sig00000909)
  );
  MUXF8   blk0000087e (
    .I0(sig0000091a),
    .I1(sig00000919),
    .S(sig00000813),
    .O(sig0000090a)
  );
  MUXF8   blk0000087f (
    .I0(sig0000091c),
    .I1(sig0000091b),
    .S(sig00000813),
    .O(sig0000090b)
  );
  MUXF8   blk00000880 (
    .I0(sig0000091e),
    .I1(sig0000091d),
    .S(sig00000813),
    .O(sig0000090c)
  );
  MUXF7   blk00000881 (
    .I0(sig00000928),
    .I1(sig0000091f),
    .S(sig00000812),
    .O(sig0000090d)
  );
  MUXF7   blk00000882 (
    .I0(sig0000093a),
    .I1(sig00000931),
    .S(sig00000812),
    .O(sig0000090e)
  );
  MUXF7   blk00000883 (
    .I0(sig00000929),
    .I1(sig00000920),
    .S(sig00000812),
    .O(sig0000090f)
  );
  MUXF7   blk00000884 (
    .I0(sig0000093b),
    .I1(sig00000932),
    .S(sig00000812),
    .O(sig00000910)
  );
  MUXF7   blk00000885 (
    .I0(sig0000092a),
    .I1(sig00000921),
    .S(sig00000812),
    .O(sig00000911)
  );
  MUXF7   blk00000886 (
    .I0(sig0000093c),
    .I1(sig00000933),
    .S(sig00000812),
    .O(sig00000912)
  );
  MUXF7   blk00000887 (
    .I0(sig0000092b),
    .I1(sig00000922),
    .S(sig00000812),
    .O(sig00000913)
  );
  MUXF7   blk00000888 (
    .I0(sig0000093d),
    .I1(sig00000934),
    .S(sig00000812),
    .O(sig00000914)
  );
  MUXF7   blk00000889 (
    .I0(sig0000092c),
    .I1(sig00000923),
    .S(sig00000812),
    .O(sig00000915)
  );
  MUXF7   blk0000088a (
    .I0(sig0000093e),
    .I1(sig00000935),
    .S(sig00000812),
    .O(sig00000916)
  );
  MUXF7   blk0000088b (
    .I0(sig0000092d),
    .I1(sig00000924),
    .S(sig00000812),
    .O(sig00000917)
  );
  MUXF7   blk0000088c (
    .I0(sig0000093f),
    .I1(sig00000936),
    .S(sig00000812),
    .O(sig00000918)
  );
  MUXF7   blk0000088d (
    .I0(sig0000092e),
    .I1(sig00000925),
    .S(sig00000812),
    .O(sig00000919)
  );
  MUXF7   blk0000088e (
    .I0(sig00000940),
    .I1(sig00000937),
    .S(sig00000812),
    .O(sig0000091a)
  );
  MUXF7   blk0000088f (
    .I0(sig0000092f),
    .I1(sig00000926),
    .S(sig00000812),
    .O(sig0000091b)
  );
  MUXF7   blk00000890 (
    .I0(sig00000941),
    .I1(sig00000938),
    .S(sig00000812),
    .O(sig0000091c)
  );
  MUXF7   blk00000891 (
    .I0(sig00000930),
    .I1(sig00000927),
    .S(sig00000812),
    .O(sig0000091d)
  );
  MUXF7   blk00000892 (
    .I0(sig00000942),
    .I1(sig00000939),
    .S(sig00000812),
    .O(sig0000091e)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk00000893 (
    .I0(sig00000002),
    .I1(sig00000002),
    .I2(sig00000002),
    .I3(sig00000002),
    .I4(sig00000810),
    .I5(sig00000811),
    .O(sig0000091f)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk00000894 (
    .I0(sig00000002),
    .I1(sig00000002),
    .I2(sig00000002),
    .I3(sig00000002),
    .I4(sig00000810),
    .I5(sig00000811),
    .O(sig00000920)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk00000895 (
    .I0(sig00000002),
    .I1(sig00000002),
    .I2(sig00000002),
    .I3(sig00000002),
    .I4(sig00000810),
    .I5(sig00000811),
    .O(sig00000921)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk00000896 (
    .I0(sig00000002),
    .I1(sig00000002),
    .I2(sig00000002),
    .I3(sig00000002),
    .I4(sig00000810),
    .I5(sig00000811),
    .O(sig00000922)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk00000897 (
    .I0(sig00000002),
    .I1(sig00000002),
    .I2(sig00000002),
    .I3(sig00000002),
    .I4(sig00000810),
    .I5(sig00000811),
    .O(sig00000923)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk00000898 (
    .I0(sig00000002),
    .I1(sig00000002),
    .I2(sig00000002),
    .I3(sig00000002),
    .I4(sig00000810),
    .I5(sig00000811),
    .O(sig00000924)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk00000899 (
    .I0(sig00000002),
    .I1(sig00000002),
    .I2(sig00000002),
    .I3(sig00000002),
    .I4(sig00000810),
    .I5(sig00000811),
    .O(sig00000925)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk0000089a (
    .I0(sig00000002),
    .I1(sig00000002),
    .I2(sig00000002),
    .I3(sig00000002),
    .I4(sig00000810),
    .I5(sig00000811),
    .O(sig00000926)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk0000089b (
    .I0(sig00000002),
    .I1(sig00000002),
    .I2(sig00000002),
    .I3(sig00000002),
    .I4(sig00000810),
    .I5(sig00000811),
    .O(sig00000927)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk0000089c (
    .I0(sig00000814),
    .I1(sig00000002),
    .I2(sig00000002),
    .I3(sig00000002),
    .I4(sig00000810),
    .I5(sig00000811),
    .O(sig00000928)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk0000089d (
    .I0(sig00000815),
    .I1(sig00000002),
    .I2(sig00000002),
    .I3(sig00000002),
    .I4(sig00000810),
    .I5(sig00000811),
    .O(sig00000929)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk0000089e (
    .I0(sig00000816),
    .I1(sig00000002),
    .I2(sig00000002),
    .I3(sig00000002),
    .I4(sig00000810),
    .I5(sig00000811),
    .O(sig0000092a)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk0000089f (
    .I0(sig00000817),
    .I1(sig00000002),
    .I2(sig00000002),
    .I3(sig00000002),
    .I4(sig00000810),
    .I5(sig00000811),
    .O(sig0000092b)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000008a0 (
    .I0(sig00000818),
    .I1(sig00000002),
    .I2(sig00000002),
    .I3(sig00000002),
    .I4(sig00000810),
    .I5(sig00000811),
    .O(sig0000092c)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000008a1 (
    .I0(sig00000819),
    .I1(sig00000002),
    .I2(sig00000002),
    .I3(sig00000002),
    .I4(sig00000810),
    .I5(sig00000811),
    .O(sig0000092d)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000008a2 (
    .I0(sig0000081a),
    .I1(sig00000002),
    .I2(sig00000002),
    .I3(sig00000002),
    .I4(sig00000810),
    .I5(sig00000811),
    .O(sig0000092e)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000008a3 (
    .I0(sig0000081b),
    .I1(sig00000002),
    .I2(sig00000002),
    .I3(sig00000002),
    .I4(sig00000810),
    .I5(sig00000811),
    .O(sig0000092f)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000008a4 (
    .I0(sig00000002),
    .I1(sig00000002),
    .I2(sig00000002),
    .I3(sig00000002),
    .I4(sig00000810),
    .I5(sig00000811),
    .O(sig00000930)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000008a5 (
    .I0(sig00000002),
    .I1(sig00000002),
    .I2(sig00000002),
    .I3(sig00000002),
    .I4(sig00000810),
    .I5(sig00000811),
    .O(sig00000931)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000008a6 (
    .I0(sig00000002),
    .I1(sig00000002),
    .I2(sig00000002),
    .I3(sig00000814),
    .I4(sig00000810),
    .I5(sig00000811),
    .O(sig00000932)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000008a7 (
    .I0(sig00000002),
    .I1(sig00000002),
    .I2(sig00000814),
    .I3(sig00000815),
    .I4(sig00000810),
    .I5(sig00000811),
    .O(sig00000933)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000008a8 (
    .I0(sig00000002),
    .I1(sig00000814),
    .I2(sig00000815),
    .I3(sig00000816),
    .I4(sig00000810),
    .I5(sig00000811),
    .O(sig00000934)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000008a9 (
    .I0(sig00000814),
    .I1(sig00000815),
    .I2(sig00000816),
    .I3(sig00000817),
    .I4(sig00000810),
    .I5(sig00000811),
    .O(sig00000935)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000008aa (
    .I0(sig00000815),
    .I1(sig00000816),
    .I2(sig00000817),
    .I3(sig00000818),
    .I4(sig00000810),
    .I5(sig00000811),
    .O(sig00000936)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000008ab (
    .I0(sig00000816),
    .I1(sig00000817),
    .I2(sig00000818),
    .I3(sig00000819),
    .I4(sig00000810),
    .I5(sig00000811),
    .O(sig00000937)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000008ac (
    .I0(sig00000817),
    .I1(sig00000818),
    .I2(sig00000819),
    .I3(sig0000081a),
    .I4(sig00000810),
    .I5(sig00000811),
    .O(sig00000938)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000008ad (
    .I0(sig00000002),
    .I1(sig00000002),
    .I2(sig00000002),
    .I3(sig00000002),
    .I4(sig00000810),
    .I5(sig00000811),
    .O(sig00000939)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000008ae (
    .I0(sig00000002),
    .I1(sig00000002),
    .I2(sig00000002),
    .I3(sig00000002),
    .I4(sig00000810),
    .I5(sig00000811),
    .O(sig0000093a)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000008af (
    .I0(sig00000002),
    .I1(sig00000002),
    .I2(sig00000002),
    .I3(sig00000002),
    .I4(sig00000810),
    .I5(sig00000811),
    .O(sig0000093b)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000008b0 (
    .I0(sig00000002),
    .I1(sig00000002),
    .I2(sig00000002),
    .I3(sig00000002),
    .I4(sig00000810),
    .I5(sig00000811),
    .O(sig0000093c)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000008b1 (
    .I0(sig00000002),
    .I1(sig00000002),
    .I2(sig00000002),
    .I3(sig00000002),
    .I4(sig00000810),
    .I5(sig00000811),
    .O(sig0000093d)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000008b2 (
    .I0(sig00000002),
    .I1(sig00000002),
    .I2(sig00000002),
    .I3(sig00000002),
    .I4(sig00000810),
    .I5(sig00000811),
    .O(sig0000093e)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000008b3 (
    .I0(sig00000002),
    .I1(sig00000002),
    .I2(sig00000002),
    .I3(sig00000814),
    .I4(sig00000810),
    .I5(sig00000811),
    .O(sig0000093f)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000008b4 (
    .I0(sig00000002),
    .I1(sig00000002),
    .I2(sig00000814),
    .I3(sig00000815),
    .I4(sig00000810),
    .I5(sig00000811),
    .O(sig00000940)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000008b5 (
    .I0(sig00000002),
    .I1(sig00000814),
    .I2(sig00000815),
    .I3(sig00000816),
    .I4(sig00000810),
    .I5(sig00000811),
    .O(sig00000941)
  );
  LUT6 #(
    .INIT ( 64'hFF00F0F0CCCCAAAA ))
  blk000008b6 (
    .I0(sig00000002),
    .I1(sig00000002),
    .I2(sig00000002),
    .I3(sig00000002),
    .I4(sig00000810),
    .I5(sig00000811),
    .O(sig00000942)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000008b7 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000943),
    .R(sig00000002),
    .Q(sig0000081c)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000008b8 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000904),
    .R(sig00000002),
    .Q(sig00000943)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000008b9 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000944),
    .R(sig00000002),
    .Q(sig0000081d)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000008ba (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000905),
    .R(sig00000002),
    .Q(sig00000944)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000008bb (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000945),
    .R(sig00000002),
    .Q(sig0000081e)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000008bc (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000906),
    .R(sig00000002),
    .Q(sig00000945)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000008bd (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000946),
    .R(sig00000002),
    .Q(sig0000081f)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000008be (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000907),
    .R(sig00000002),
    .Q(sig00000946)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000008bf (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000947),
    .R(sig00000002),
    .Q(sig00000820)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000008c0 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000908),
    .R(sig00000002),
    .Q(sig00000947)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000008c1 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000948),
    .R(sig00000002),
    .Q(sig00000821)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000008c2 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000909),
    .R(sig00000002),
    .Q(sig00000948)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000008c3 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000949),
    .R(sig00000002),
    .Q(sig00000822)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000008c4 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000090a),
    .R(sig00000002),
    .Q(sig00000949)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000008c5 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000094a),
    .R(sig00000002),
    .Q(sig00000823)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000008c6 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000090b),
    .R(sig00000002),
    .Q(sig0000094a)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000008c7 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000094b),
    .R(sig00000002),
    .Q(NLW_blk000008c7_Q_UNCONNECTED)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000008c8 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000090c),
    .R(sig00000002),
    .Q(sig0000094b)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000008c9 (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig0000080e),
    .Q(sig0000094c)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000008ca (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig0000080d),
    .Q(sig0000094d)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000008cb (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig0000080c),
    .Q(sig0000094e)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000008cc (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig0000080b),
    .Q(sig0000094f)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000008cd (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig0000080a),
    .Q(sig00000950)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000008ce (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig00000809),
    .Q(sig00000951)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000008cf (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig00000808),
    .Q(sig00000952)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000008d0 (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig00000807),
    .Q(sig00000953)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000008d1 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000094c),
    .R(sig00000002),
    .Q(sig0000081b)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000008d2 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000094d),
    .R(sig00000002),
    .Q(sig0000081a)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000008d3 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000094e),
    .R(sig00000002),
    .Q(sig00000819)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000008d4 (
    .C(clk),
    .CE(sig00000001),
    .D(sig0000094f),
    .R(sig00000002),
    .Q(sig00000818)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000008d5 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000950),
    .R(sig00000002),
    .Q(sig00000817)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000008d6 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000951),
    .R(sig00000002),
    .Q(sig00000816)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000008d7 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000952),
    .R(sig00000002),
    .Q(sig00000815)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000008d8 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000953),
    .R(sig00000002),
    .Q(sig00000814)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000008d9 (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig00000806),
    .Q(sig00000954)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000008da (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig00000805),
    .Q(sig00000955)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000008db (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig00000804),
    .Q(sig00000956)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000008dc (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig00000803),
    .Q(sig00000957)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000008dd (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000954),
    .R(sig00000002),
    .Q(sig00000813)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000008de (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000955),
    .R(sig00000002),
    .Q(sig00000812)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000008df (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000956),
    .R(sig00000002),
    .Q(sig00000811)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000008e0 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000957),
    .R(sig00000002),
    .Q(sig00000810)
  );
  LUT6 #(
    .INIT ( 64'h9009000000009009 ))
  blk000008eb (
    .I0(sig000009a3),
    .I1(sig000009b6),
    .I2(sig000009a2),
    .I3(sig000009b7),
    .I4(sig000009a1),
    .I5(sig000009b8),
    .O(sig00000958)
  );
  LUT6 #(
    .INIT ( 64'h9009000000009009 ))
  blk000008ec (
    .I0(sig000009a6),
    .I1(sig000009b3),
    .I2(sig000009a5),
    .I3(sig000009b4),
    .I4(sig000009a4),
    .I5(sig000009b5),
    .O(sig00000959)
  );
  LUT6 #(
    .INIT ( 64'h9009000000009009 ))
  blk000008ed (
    .I0(sig000009a9),
    .I1(sig00000001),
    .I2(sig000009a8),
    .I3(sig00000002),
    .I4(sig000009a7),
    .I5(sig000009b2),
    .O(sig0000095a)
  );
  MUXCY   blk000008ee (
    .CI(sig0000095c),
    .DI(sig00000002),
    .S(sig00000958),
    .O(sig0000095b)
  );
  MUXCY   blk000008ef (
    .CI(sig0000095d),
    .DI(sig00000002),
    .S(sig00000959),
    .O(sig0000095c)
  );
  MUXCY   blk000008f0 (
    .CI(sig00000001),
    .DI(sig00000002),
    .S(sig0000095a),
    .O(sig0000095d)
  );
  XORCY   blk000008f1 (
    .CI(sig0000095b),
    .LI(sig00000002),
    .O(sig00000977)
  );
  LUT6 #(
    .INIT ( 64'h9009000000009009 ))
  blk000008f2 (
    .I0(NlwRenamedSig_OI_xn_index[6]),
    .I1(sig000009b6),
    .I2(NlwRenamedSig_OI_xn_index[7]),
    .I3(sig000009b7),
    .I4(NlwRenamedSig_OI_xn_index[8]),
    .I5(sig000009b8),
    .O(sig0000095e)
  );
  LUT6 #(
    .INIT ( 64'h9009000000009009 ))
  blk000008f3 (
    .I0(NlwRenamedSig_OI_xn_index[3]),
    .I1(sig000009b3),
    .I2(NlwRenamedSig_OI_xn_index[4]),
    .I3(sig000009b4),
    .I4(NlwRenamedSig_OI_xn_index[5]),
    .I5(sig000009b5),
    .O(sig0000095f)
  );
  LUT6 #(
    .INIT ( 64'h9009000000009009 ))
  blk000008f4 (
    .I0(NlwRenamedSig_OI_xn_index[0]),
    .I1(sig00000001),
    .I2(NlwRenamedSig_OI_xn_index[1]),
    .I3(sig00000002),
    .I4(NlwRenamedSig_OI_xn_index[2]),
    .I5(sig000009b2),
    .O(sig00000960)
  );
  MUXCY   blk000008f5 (
    .CI(sig00000962),
    .DI(sig00000002),
    .S(sig0000095e),
    .O(sig00000961)
  );
  MUXCY   blk000008f6 (
    .CI(sig00000963),
    .DI(sig00000002),
    .S(sig0000095f),
    .O(sig00000962)
  );
  MUXCY   blk000008f7 (
    .CI(sig00000001),
    .DI(sig00000002),
    .S(sig00000960),
    .O(sig00000963)
  );
  XORCY   blk000008f8 (
    .CI(sig00000961),
    .LI(sig00000002),
    .O(sig00000964)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000008f9 (
    .C(clk),
    .CE(\NlwRenamedSig_OI_U0/i_synth/non_floating_point.arch_c.xfft_inst/control/cntrl/loading_state/ORS ),
    .D(sig00000964),
    .R(sig00000002),
    .Q(sig000009ab)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000008fa (
    .C(clk),
    .CE(\NlwRenamedSig_OI_U0/i_synth/non_floating_point.arch_c.xfft_inst/control/cntrl/loading_state/ORS ),
    .D(sig000009ab),
    .R(sig00000002),
    .Q(sig000009aa)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000008fb (
    .C(clk),
    .CE(\NlwRenamedSig_OI_U0/i_synth/non_floating_point.arch_c.xfft_inst/control/cntrl/loading_state/ORS ),
    .D(sig0000096e),
    .R(sig00000002),
    .Q(NlwRenamedSig_OI_xn_index[8])
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000008fc (
    .C(clk),
    .CE(\NlwRenamedSig_OI_U0/i_synth/non_floating_point.arch_c.xfft_inst/control/cntrl/loading_state/ORS ),
    .D(sig0000096f),
    .R(sig00000002),
    .Q(NlwRenamedSig_OI_xn_index[7])
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000008fd (
    .C(clk),
    .CE(\NlwRenamedSig_OI_U0/i_synth/non_floating_point.arch_c.xfft_inst/control/cntrl/loading_state/ORS ),
    .D(sig00000970),
    .R(sig00000002),
    .Q(NlwRenamedSig_OI_xn_index[6])
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000008fe (
    .C(clk),
    .CE(\NlwRenamedSig_OI_U0/i_synth/non_floating_point.arch_c.xfft_inst/control/cntrl/loading_state/ORS ),
    .D(sig00000971),
    .R(sig00000002),
    .Q(NlwRenamedSig_OI_xn_index[5])
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000008ff (
    .C(clk),
    .CE(\NlwRenamedSig_OI_U0/i_synth/non_floating_point.arch_c.xfft_inst/control/cntrl/loading_state/ORS ),
    .D(sig00000972),
    .R(sig00000002),
    .Q(NlwRenamedSig_OI_xn_index[4])
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000900 (
    .C(clk),
    .CE(\NlwRenamedSig_OI_U0/i_synth/non_floating_point.arch_c.xfft_inst/control/cntrl/loading_state/ORS ),
    .D(sig00000973),
    .R(sig00000002),
    .Q(NlwRenamedSig_OI_xn_index[3])
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000901 (
    .C(clk),
    .CE(\NlwRenamedSig_OI_U0/i_synth/non_floating_point.arch_c.xfft_inst/control/cntrl/loading_state/ORS ),
    .D(sig00000974),
    .R(sig00000002),
    .Q(NlwRenamedSig_OI_xn_index[2])
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000902 (
    .C(clk),
    .CE(\NlwRenamedSig_OI_U0/i_synth/non_floating_point.arch_c.xfft_inst/control/cntrl/loading_state/ORS ),
    .D(sig00000975),
    .R(sig00000002),
    .Q(NlwRenamedSig_OI_xn_index[1])
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000903 (
    .C(clk),
    .CE(\NlwRenamedSig_OI_U0/i_synth/non_floating_point.arch_c.xfft_inst/control/cntrl/loading_state/ORS ),
    .D(sig00000976),
    .R(sig00000002),
    .Q(NlwRenamedSig_OI_xn_index[0])
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000904 (
    .C(clk),
    .CE(sig000007f9),
    .D(sig00000977),
    .R(sig00000002),
    .Q(sig000009a0)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000905 (
    .C(clk),
    .CE(sig000007f9),
    .D(sig000009a0),
    .R(sig00000002),
    .Q(sig0000099f)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000906 (
    .C(clk),
    .CE(sig000007f9),
    .D(sig00000981),
    .R(sig00000002),
    .Q(sig000009a1)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000907 (
    .C(clk),
    .CE(sig000007f9),
    .D(sig00000982),
    .R(sig00000002),
    .Q(sig000009a2)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000908 (
    .C(clk),
    .CE(sig000007f9),
    .D(sig00000983),
    .R(sig00000002),
    .Q(sig000009a3)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000909 (
    .C(clk),
    .CE(sig000007f9),
    .D(sig00000984),
    .R(sig00000002),
    .Q(sig000009a4)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000090a (
    .C(clk),
    .CE(sig000007f9),
    .D(sig00000985),
    .R(sig00000002),
    .Q(sig000009a5)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000090b (
    .C(clk),
    .CE(sig000007f9),
    .D(sig00000986),
    .R(sig00000002),
    .Q(sig000009a6)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000090c (
    .C(clk),
    .CE(sig000007f9),
    .D(sig00000987),
    .R(sig00000002),
    .Q(sig000009a7)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000090d (
    .C(clk),
    .CE(sig000007f9),
    .D(sig00000988),
    .R(sig00000002),
    .Q(sig000009a8)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000090e (
    .C(clk),
    .CE(sig000007f9),
    .D(sig00000989),
    .R(sig00000002),
    .Q(sig000009a9)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk0000090f (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000001),
    .Q(sig000009ae)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000910 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000001),
    .Q(sig000009af)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000911 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000001),
    .Q(sig000009b0)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000912 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000002),
    .Q(sig000009b1)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000913 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000001),
    .Q(sig000009b2)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000914 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000001),
    .Q(sig000009b3)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000915 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000001),
    .Q(sig000009b4)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000916 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000001),
    .Q(sig000009b5)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000917 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000001),
    .Q(sig000009b6)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000918 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000001),
    .Q(sig000009b7)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000919 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000001),
    .Q(sig000009b8)
  );
  FDR #(
    .INIT ( 1'b0 ))
  blk0000091a (
    .C(clk),
    .D(\NlwRenamedSig_OI_U0/i_synth/non_floating_point.arch_c.xfft_inst/control/cntrl/process_state_r ),
    .R(sig00000002),
    .Q(\U0/i_synth/non_floating_point.arch_c.xfft_inst/control/cntrl/done_pr_d_1 )
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000091b (
    .C(clk),
    .D(sig0000098a),
    .Q(sig0000099e)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000091c (
    .C(clk),
    .D(sig0000098e),
    .Q(sig00000802)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000091d (
    .C(clk),
    .D(sig0000098f),
    .Q(sig00000801)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000091e (
    .C(clk),
    .D(sig00000990),
    .Q(sig00000800)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk0000091f (
    .C(clk),
    .D(sig00000991),
    .Q(sig000007ff)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000920 (
    .C(clk),
    .D(sig00000992),
    .Q(sig000007fe)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000921 (
    .C(clk),
    .D(sig00000993),
    .Q(sig000007fd)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000922 (
    .C(clk),
    .D(sig00000994),
    .Q(sig000007fc)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000923 (
    .C(clk),
    .D(sig00000995),
    .Q(sig000007fb)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000924 (
    .C(clk),
    .D(sig00000996),
    .Q(sig000007fa)
  );
  LUT6 #(
    .INIT ( 64'h9009000000009009 ))
  blk00000925 (
    .I0(sig0000080d),
    .I1(sig000009b7),
    .I2(sig0000080e),
    .I3(sig000009b8),
    .I4(sig00000002),
    .I5(sig00000002),
    .O(sig000009b9)
  );
  LUT6 #(
    .INIT ( 64'h9009000000009009 ))
  blk00000926 (
    .I0(sig0000080a),
    .I1(sig000009b4),
    .I2(sig0000080b),
    .I3(sig000009b5),
    .I4(sig0000080c),
    .I5(sig000009b6),
    .O(sig000009ba)
  );
  LUT6 #(
    .INIT ( 64'h9009000000009009 ))
  blk00000927 (
    .I0(sig00000807),
    .I1(sig00000002),
    .I2(sig00000808),
    .I3(sig000009b2),
    .I4(sig00000809),
    .I5(sig000009b3),
    .O(sig000009bb)
  );
  MUXCY   blk00000928 (
    .CI(sig000009bd),
    .DI(sig00000002),
    .S(sig000009b9),
    .O(sig000009bc)
  );
  MUXCY   blk00000929 (
    .CI(sig000009be),
    .DI(sig00000002),
    .S(sig000009ba),
    .O(sig000009bd)
  );
  MUXCY   blk0000092a (
    .CI(sig00000001),
    .DI(sig00000002),
    .S(sig000009bb),
    .O(sig000009be)
  );
  XORCY   blk0000092b (
    .CI(sig000009bc),
    .LI(sig00000002),
    .O(sig000009cf)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000092c (
    .C(clk),
    .CE(sig000007f8),
    .D(sig000009bf),
    .R(\NlwRenamedSig_OI_U0/i_synth/non_floating_point.arch_c.xfft_inst/control/cntrl/loading_state/ORS ),
    .Q(sig00000807)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000092d (
    .C(clk),
    .CE(sig000007f8),
    .D(sig000009c0),
    .R(\NlwRenamedSig_OI_U0/i_synth/non_floating_point.arch_c.xfft_inst/control/cntrl/loading_state/ORS ),
    .Q(sig00000808)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000092e (
    .C(clk),
    .CE(sig000007f8),
    .D(sig000009c1),
    .R(\NlwRenamedSig_OI_U0/i_synth/non_floating_point.arch_c.xfft_inst/control/cntrl/loading_state/ORS ),
    .Q(sig00000809)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000092f (
    .C(clk),
    .CE(sig000007f8),
    .D(sig000009c2),
    .R(\NlwRenamedSig_OI_U0/i_synth/non_floating_point.arch_c.xfft_inst/control/cntrl/loading_state/ORS ),
    .Q(sig0000080a)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000930 (
    .C(clk),
    .CE(sig000007f8),
    .D(sig000009c3),
    .R(\NlwRenamedSig_OI_U0/i_synth/non_floating_point.arch_c.xfft_inst/control/cntrl/loading_state/ORS ),
    .Q(sig0000080b)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000931 (
    .C(clk),
    .CE(sig000007f8),
    .D(sig000009c4),
    .R(\NlwRenamedSig_OI_U0/i_synth/non_floating_point.arch_c.xfft_inst/control/cntrl/loading_state/ORS ),
    .Q(sig0000080c)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000932 (
    .C(clk),
    .CE(sig000007f8),
    .D(sig000009c5),
    .R(\NlwRenamedSig_OI_U0/i_synth/non_floating_point.arch_c.xfft_inst/control/cntrl/loading_state/ORS ),
    .Q(sig0000080d)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000933 (
    .C(clk),
    .CE(sig000007f8),
    .D(sig000009c6),
    .R(\NlwRenamedSig_OI_U0/i_synth/non_floating_point.arch_c.xfft_inst/control/cntrl/loading_state/ORS ),
    .Q(sig0000080e)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000934 (
    .C(clk),
    .CE(sig000007f8),
    .D(sig000009cf),
    .R(\NlwRenamedSig_OI_U0/i_synth/non_floating_point.arch_c.xfft_inst/control/cntrl/loading_state/ORS ),
    .Q(sig0000098d)
  );
  LUT6 #(
    .INIT ( 64'h9009000000009009 ))
  blk0000094e (
    .I0(sig000009e2),
    .I1(sig00000002),
    .I2(sig000009e3),
    .I3(sig00000001),
    .I4(sig00000002),
    .I5(sig00000002),
    .O(sig000009d0)
  );
  LUT6 #(
    .INIT ( 64'h9009000000009009 ))
  blk0000094f (
    .I0(sig000009df),
    .I1(sig00000001),
    .I2(sig000009e0),
    .I3(sig00000001),
    .I4(sig000009e1),
    .I5(sig00000002),
    .O(sig000009d1)
  );
  MUXCY   blk00000950 (
    .CI(sig000009d3),
    .DI(sig00000002),
    .S(sig000009d0),
    .O(sig000009d2)
  );
  MUXCY   blk00000951 (
    .CI(sig00000001),
    .DI(sig00000002),
    .S(sig000009d1),
    .O(sig000009d3)
  );
  XORCY   blk00000952 (
    .CI(sig000009d2),
    .LI(sig00000002),
    .O(sig000009d9)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000953 (
    .C(clk),
    .CE(sig00000997),
    .D(sig000009d4),
    .R(sig00000002),
    .Q(sig000009df)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000954 (
    .C(clk),
    .CE(sig00000997),
    .D(sig000009d5),
    .R(sig00000002),
    .Q(sig000009e0)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000955 (
    .C(clk),
    .CE(sig00000997),
    .D(sig000009d6),
    .R(sig00000002),
    .Q(sig000009e1)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000956 (
    .C(clk),
    .CE(sig00000997),
    .D(sig000009d7),
    .R(sig00000002),
    .Q(sig000009e2)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000957 (
    .C(clk),
    .CE(sig00000997),
    .D(sig000009d8),
    .R(sig00000002),
    .Q(sig000009e3)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000958 (
    .C(clk),
    .CE(sig00000997),
    .D(sig000009ad),
    .R(sig00000002),
    .Q(sig00000003)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000959 (
    .C(clk),
    .CE(sig00000997),
    .D(sig000009d9),
    .R(sig00000002),
    .Q(sig000009ad)
  );
  LUT6 #(
    .INIT ( 64'h9009000000009009 ))
  blk0000096a (
    .I0(sig00000806),
    .I1(sig000009b1),
    .I2(sig00000002),
    .I3(sig00000002),
    .I4(sig00000002),
    .I5(sig00000002),
    .O(sig000009e4)
  );
  LUT6 #(
    .INIT ( 64'h9009000000009009 ))
  blk0000096b (
    .I0(sig00000803),
    .I1(sig000009ae),
    .I2(sig00000804),
    .I3(sig000009af),
    .I4(sig00000805),
    .I5(sig000009b0),
    .O(sig000009e5)
  );
  MUXCY   blk0000096c (
    .CI(sig000009e7),
    .DI(sig00000002),
    .S(sig000009e4),
    .O(sig000009e6)
  );
  MUXCY   blk0000096d (
    .CI(sig00000001),
    .DI(sig00000002),
    .S(sig000009e5),
    .O(sig000009e7)
  );
  XORCY   blk0000096e (
    .CI(sig000009e6),
    .LI(sig00000002),
    .O(sig000009f0)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk0000096f (
    .C(clk),
    .CE(sig0000098b),
    .D(sig000009e8),
    .R(sig0000099b),
    .Q(sig00000803)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000970 (
    .C(clk),
    .CE(sig0000098b),
    .D(sig000009e9),
    .R(sig0000099b),
    .Q(sig00000804)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000971 (
    .C(clk),
    .CE(sig0000098b),
    .D(sig000009ea),
    .R(sig0000099b),
    .Q(sig00000805)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000972 (
    .C(clk),
    .CE(sig0000098b),
    .D(sig000009eb),
    .R(sig0000099b),
    .Q(sig00000806)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk00000973 (
    .C(clk),
    .CE(sig0000098b),
    .D(sig000009f0),
    .R(sig0000099b),
    .Q(sig000009ac)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000009b9 (
    .A0(sig00000001),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig00000802),
    .Q(sig000009f1)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000009ba (
    .A0(sig00000001),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig00000801),
    .Q(sig000009f2)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000009bb (
    .A0(sig00000001),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig00000800),
    .Q(sig000009f3)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000009bc (
    .A0(sig00000001),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000007ff),
    .Q(sig000009f4)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000009bd (
    .A0(sig00000001),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000007fe),
    .Q(sig000009f5)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000009be (
    .A0(sig00000001),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000007fd),
    .Q(sig000009f6)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000009bf (
    .A0(sig00000001),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000007fc),
    .Q(sig000009f7)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000009c0 (
    .A0(sig00000001),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000007fb),
    .Q(sig000009f8)
  );
  SRL16E #(
    .INIT ( 16'h0000 ))
  blk000009c1 (
    .A0(sig00000001),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000007fa),
    .Q(sig000009f9)
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000009c2 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000009f1),
    .R(sig00000002),
    .Q(xk_index[8])
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000009c3 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000009f2),
    .R(sig00000002),
    .Q(xk_index[7])
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000009c4 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000009f3),
    .R(sig00000002),
    .Q(xk_index[6])
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000009c5 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000009f4),
    .R(sig00000002),
    .Q(xk_index[5])
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000009c6 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000009f5),
    .R(sig00000002),
    .Q(xk_index[4])
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000009c7 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000009f6),
    .R(sig00000002),
    .Q(xk_index[3])
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000009c8 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000009f7),
    .R(sig00000002),
    .Q(xk_index[2])
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000009c9 (
    .C(clk),
    .CE(sig00000001),
    .D(sig000009f8),
    .R(sig00000002),
    .Q(xk_index[1])
  );
  FDRE #(
    .INIT ( 1'b0 ))
  blk000009ca (
    .C(clk),
    .CE(sig00000001),
    .D(sig000009f9),
    .R(sig00000002),
    .Q(xk_index[0])
  );
  LUT5 #(
    .INIT ( 32'h6666666A ))
  blk000009d3 (
    .I0(sig0000001a),
    .I1(sig00000042),
    .I2(sig00000017),
    .I3(sig00000018),
    .I4(sig00000019),
    .O(sig0000051d)
  );
  LUT6 #(
    .INIT ( 64'h666666666666666A ))
  blk000009d4 (
    .I0(sig0000001b),
    .I1(sig00000042),
    .I2(sig00000017),
    .I3(sig00000018),
    .I4(sig00000019),
    .I5(sig0000001a),
    .O(sig0000051e)
  );
  LUT5 #(
    .INIT ( 32'hFFFFFFFE ))
  blk000009d5 (
    .I0(sig0000001b),
    .I1(sig00000017),
    .I2(sig00000018),
    .I3(sig00000019),
    .I4(sig0000001a),
    .O(sig0000051a)
  );
  LUT4 #(
    .INIT ( 16'h666A ))
  blk000009d6 (
    .I0(sig0000001d),
    .I1(sig00000042),
    .I2(sig0000001c),
    .I3(sig0000051a),
    .O(sig00000520)
  );
  LUT4 #(
    .INIT ( 16'h666A ))
  blk000009d7 (
    .I0(sig00000019),
    .I1(sig00000042),
    .I2(sig00000017),
    .I3(sig00000018),
    .O(sig0000051c)
  );
  LUT3 #(
    .INIT ( 8'h6A ))
  blk000009d8 (
    .I0(sig0000001c),
    .I1(sig00000042),
    .I2(sig0000051a),
    .O(sig0000051f)
  );
  LUT3 #(
    .INIT ( 8'h6A ))
  blk000009d9 (
    .I0(sig00000018),
    .I1(sig00000017),
    .I2(sig00000042),
    .O(sig0000051b)
  );
  LUT4 #(
    .INIT ( 16'h2220 ))
  blk000009da (
    .I0(sig000005e3),
    .I1(sig000005e5),
    .I2(sig000005e7),
    .I3(sig000005e6),
    .O(sig000005e2)
  );
  LUT2 #(
    .INIT ( 4'hE ))
  blk000009db (
    .I0(sig000001c8),
    .I1(sig000001c7),
    .O(sig0000060f)
  );
  LUT4 #(
    .INIT ( 16'h2220 ))
  blk000009dc (
    .I0(sig00000611),
    .I1(sig00000613),
    .I2(sig00000615),
    .I3(sig00000614),
    .O(sig00000610)
  );
  LUT2 #(
    .INIT ( 4'hE ))
  blk000009dd (
    .I0(sig000001de),
    .I1(sig000001dd),
    .O(sig0000063d)
  );
  LUT4 #(
    .INIT ( 16'h2220 ))
  blk000009de (
    .I0(sig0000063f),
    .I1(sig00000641),
    .I2(sig00000643),
    .I3(sig00000642),
    .O(sig0000063e)
  );
  LUT2 #(
    .INIT ( 4'hE ))
  blk000009df (
    .I0(sig000001f4),
    .I1(sig000001f3),
    .O(sig0000066b)
  );
  LUT4 #(
    .INIT ( 16'h2220 ))
  blk000009e0 (
    .I0(sig0000066d),
    .I1(sig0000066f),
    .I2(sig00000671),
    .I3(sig00000670),
    .O(sig0000066c)
  );
  LUT2 #(
    .INIT ( 4'hE ))
  blk000009e1 (
    .I0(sig0000020a),
    .I1(sig00000209),
    .O(sig00000699)
  );
  LUT3 #(
    .INIT ( 8'hAC ))
  blk000009e2 (
    .I0(sig00000850),
    .I1(sig00000825),
    .I2(sig0000000b),
    .O(sig000007f4)
  );
  LUT3 #(
    .INIT ( 8'h5C ))
  blk000009e3 (
    .I0(sig00000850),
    .I1(sig00000825),
    .I2(sig0000000b),
    .O(sig000007f5)
  );
  LUT3 #(
    .INIT ( 8'h01 ))
  blk000009e4 (
    .I0(sig00000804),
    .I1(sig00000805),
    .I2(sig00000806),
    .O(sig000008a3)
  );
  LUT4 #(
    .INIT ( 16'h0001 ))
  blk000009e5 (
    .I0(sig00000803),
    .I1(sig00000804),
    .I2(sig00000805),
    .I3(sig00000806),
    .O(sig000008b6)
  );
  LUT3 #(
    .INIT ( 8'h15 ))
  blk000009e6 (
    .I0(sig00000806),
    .I1(sig00000804),
    .I2(sig00000805),
    .O(sig000008b9)
  );
  LUT4 #(
    .INIT ( 16'h0155 ))
  blk000009e7 (
    .I0(sig00000806),
    .I1(sig00000804),
    .I2(sig00000803),
    .I3(sig00000805),
    .O(sig000008ba)
  );
  LUT4 #(
    .INIT ( 16'h0111 ))
  blk000009e8 (
    .I0(sig00000805),
    .I1(sig00000806),
    .I2(sig00000803),
    .I3(sig00000804),
    .O(sig000008b5)
  );
  LUT4 #(
    .INIT ( 16'h1555 ))
  blk000009e9 (
    .I0(sig00000806),
    .I1(sig00000803),
    .I2(sig00000804),
    .I3(sig00000805),
    .O(sig000008b8)
  );
  LUT4 #(
    .INIT ( 16'h01FF ))
  blk000009ea (
    .I0(sig00000805),
    .I1(sig00000803),
    .I2(sig00000804),
    .I3(sig00000806),
    .O(sig000008b7)
  );
  LUT2 #(
    .INIT ( 4'h1 ))
  blk000009eb (
    .I0(sig00000806),
    .I1(sig00000805),
    .O(sig000008bb)
  );
  LUT5 #(
    .INIT ( 32'h0000AAA8 ))
  blk000009ec (
    .I0(start),
    .I1(sig0000099d),
    .I2(sig0000099c),
    .I3(sig00000999),
    .I4(sig0000099a),
    .O(sig000007f7)
  );
  LUT2 #(
    .INIT ( 4'hE ))
  blk000009ed (
    .I0(sig0000099b),
    .I1(sig00000003),
    .O(sig0000098b)
  );
  LUT2 #(
    .INIT ( 4'h8 ))
  blk000009ee (
    .I0(sig000009ac),
    .I1(sig000009ad),
    .O(sig0000098c)
  );
  LUT2 #(
    .INIT ( 4'h8 ))
  blk000009ef (
    .I0(sig000009a1),
    .I1(sig000007f9),
    .O(sig0000098e)
  );
  LUT2 #(
    .INIT ( 4'h8 ))
  blk000009f0 (
    .I0(sig000009a2),
    .I1(sig000007f9),
    .O(sig0000098f)
  );
  LUT2 #(
    .INIT ( 4'h8 ))
  blk000009f1 (
    .I0(sig000009a3),
    .I1(sig000007f9),
    .O(sig00000990)
  );
  LUT2 #(
    .INIT ( 4'h8 ))
  blk000009f2 (
    .I0(sig000009a4),
    .I1(sig000007f9),
    .O(sig00000991)
  );
  LUT2 #(
    .INIT ( 4'h8 ))
  blk000009f3 (
    .I0(sig000009a5),
    .I1(sig000007f9),
    .O(sig00000992)
  );
  LUT2 #(
    .INIT ( 4'h8 ))
  blk000009f4 (
    .I0(sig000009a6),
    .I1(sig000007f9),
    .O(sig00000993)
  );
  LUT2 #(
    .INIT ( 4'h8 ))
  blk000009f5 (
    .I0(sig000009a7),
    .I1(sig000007f9),
    .O(sig00000994)
  );
  LUT2 #(
    .INIT ( 4'h8 ))
  blk000009f6 (
    .I0(sig000009a8),
    .I1(sig000007f9),
    .O(sig00000995)
  );
  LUT2 #(
    .INIT ( 4'h8 ))
  blk000009f7 (
    .I0(sig000009a9),
    .I1(sig000007f9),
    .O(sig00000996)
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  blk000009f8 (
    .I0(sig00000998),
    .I1(\NlwRenamedSig_OI_U0/i_synth/non_floating_point.arch_c.xfft_inst/control/cntrl/processing_state/ORS ),
    .O(sig00000997)
  );
  LUT2 #(
    .INIT ( 4'h8 ))
  blk000009f9 (
    .I0(sig00000998),
    .I1(\NlwRenamedSig_OI_U0/i_synth/non_floating_point.arch_c.xfft_inst/control/cntrl/processing_state/ORS ),
    .O(sig000007f8)
  );
  LUT4 #(
    .INIT ( 16'h6996 ))
  blk000009fa (
    .I0(sig00000800),
    .I1(sig000007ff),
    .I2(sig00000802),
    .I3(sig00000801),
    .O(sig000009fa)
  );
  LUT6 #(
    .INIT ( 64'h6996966996696996 ))
  blk000009fb (
    .I0(sig000007fc),
    .I1(sig000007fb),
    .I2(sig000007fe),
    .I3(sig000007fd),
    .I4(sig000007fa),
    .I5(sig000009fa),
    .O(sig000007f3)
  );
  LUT4 #(
    .INIT ( 16'h6996 ))
  blk000009fc (
    .I0(sig00000860),
    .I1(sig0000085f),
    .I2(sig00000862),
    .I3(sig00000861),
    .O(sig000009fb)
  );
  LUT6 #(
    .INIT ( 64'h6996966996696996 ))
  blk000009fd (
    .I0(sig0000085c),
    .I1(sig0000085b),
    .I2(sig0000085e),
    .I3(sig0000085d),
    .I4(sig0000085a),
    .I5(sig000009fb),
    .O(sig00000859)
  );
  LUT3 #(
    .INIT ( 8'h69 ))
  blk000009fe (
    .I0(sig0000080a),
    .I1(sig0000080e),
    .I2(sig0000080d),
    .O(sig000009fc)
  );
  LUT6 #(
    .INIT ( 64'h9669699669969669 ))
  blk000009ff (
    .I0(sig00000809),
    .I1(sig00000808),
    .I2(sig00000807),
    .I3(sig0000080c),
    .I4(sig0000080b),
    .I5(sig000009fc),
    .O(sig000008b4)
  );
  FD #(
    .INIT ( 1'b1 ))
  blk00000a00 (
    .C(clk),
    .D(sig000009fd),
    .Q(sig00000999)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000a01 (
    .C(clk),
    .D(sig0000098c),
    .Q(\NlwRenamedSig_OI_U0/i_synth/non_floating_point.arch_c.xfft_inst/control/cntrl/process_state_r )
  );
  FD #(
    .INIT ( 1'b1 ))
  blk00000a02 (
    .C(clk),
    .D(sig000009fe),
    .Q(sig00000998)
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  blk00000a03 (
    .I0(fwd_inv_we),
    .I1(sig00000041),
    .I2(fwd_inv),
    .O(sig000009ff)
  );
  FDS #(
    .INIT ( 1'b1 ))
  blk00000a04 (
    .C(clk),
    .D(sig000009ff),
    .S(sig00000002),
    .Q(sig00000041)
  );
  LUT3 #(
    .INIT ( 8'hE4 ))
  blk00000a05 (
    .I0(sig00000006),
    .I1(sig00000042),
    .I2(sig00000041),
    .O(sig00000a00)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000a06 (
    .C(clk),
    .D(sig00000a00),
    .Q(sig00000042)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000a07 (
    .C(clk),
    .D(sig00000a01),
    .Q(sig0000099a)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000a08 (
    .C(clk),
    .D(sig00000a02),
    .Q(sig0000099c)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000a09 (
    .C(clk),
    .D(sig00000a03),
    .Q(sig0000099d)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000a0a (
    .C(clk),
    .D(sig00000a04),
    .Q(sig0000099b)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000a0b (
    .C(clk),
    .D(sig00000a05),
    .Q(\NlwRenamedSig_OI_U0/i_synth/non_floating_point.arch_c.xfft_inst/control/cntrl/loading_state/ORS )
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000a0c (
    .C(clk),
    .D(sig00000a06),
    .Q(\NlwRenamedSig_OI_U0/i_synth/non_floating_point.arch_c.xfft_inst/control/cntrl/processing_state/ORS )
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000a0d (
    .C(clk),
    .D(sig00000a07),
    .Q(sig000007f9)
  );
  LUT3 #(
    .INIT ( 8'hEA ))
  blk00000a0e (
    .I0(NlwRenamedSig_OI_xn_index[0]),
    .I1(sig00000a0a),
    .I2(sig000009aa),
    .O(sig0000096d)
  );
  LUT3 #(
    .INIT ( 8'hEA ))
  blk00000a0f (
    .I0(sig000009a9),
    .I1(sig00000a09),
    .I2(sig0000099f),
    .O(sig00000980)
  );
  LUT4 #(
    .INIT ( 16'hEAAA ))
  blk00000a10 (
    .I0(sig00000807),
    .I1(sig0000098d),
    .I2(sig00000998),
    .I3(\NlwRenamedSig_OI_U0/i_synth/non_floating_point.arch_c.xfft_inst/control/cntrl/processing_state/ORS ),
    .O(sig000009c7)
  );
  LUT4 #(
    .INIT ( 16'hAEAA ))
  blk00000a11 (
    .I0(sig000009df),
    .I1(sig00000003),
    .I2(sig00000998),
    .I3(\NlwRenamedSig_OI_U0/i_synth/non_floating_point.arch_c.xfft_inst/control/cntrl/processing_state/ORS ),
    .O(sig000009da)
  );
  LUT4 #(
    .INIT ( 16'hEEEA ))
  blk00000a12 (
    .I0(sig00000803),
    .I1(sig000009ac),
    .I2(sig00000003),
    .I3(sig0000099b),
    .O(sig000009ec)
  );
  LUT3 #(
    .INIT ( 8'h54 ))
  blk00000a13 (
    .I0(sig000009aa),
    .I1(\NlwRenamedSig_OI_U0/i_synth/non_floating_point.arch_c.xfft_inst/control/cntrl/loading_state/ORS ),
    .I2(sig000007f7),
    .O(sig00000a05)
  );
  LUT6 #(
    .INIT ( 64'h5555AAAA5556AAAA ))
  blk00000a14 (
    .I0(sig0000001f),
    .I1(sig0000001e),
    .I2(sig0000001d),
    .I3(sig0000001c),
    .I4(sig00000042),
    .I5(sig0000051a),
    .O(sig00000522)
  );
  LUT5 #(
    .INIT ( 32'h55AA56AA ))
  blk00000a15 (
    .I0(sig0000001e),
    .I1(sig0000001d),
    .I2(sig0000001c),
    .I3(sig00000042),
    .I4(sig0000051a),
    .O(sig00000521)
  );
  LUT3 #(
    .INIT ( 8'hEA ))
  blk00000a16 (
    .I0(NlwRenamedSig_OI_xn_index[1]),
    .I1(sig00000a0a),
    .I2(sig000009aa),
    .O(sig0000096c)
  );
  LUT3 #(
    .INIT ( 8'hEA ))
  blk00000a17 (
    .I0(sig000009a8),
    .I1(sig00000a09),
    .I2(sig0000099f),
    .O(sig0000097f)
  );
  LUT3 #(
    .INIT ( 8'hEA ))
  blk00000a18 (
    .I0(NlwRenamedSig_OI_xn_index[2]),
    .I1(sig00000a0a),
    .I2(sig000009aa),
    .O(sig0000096b)
  );
  LUT3 #(
    .INIT ( 8'hEA ))
  blk00000a19 (
    .I0(sig000009a7),
    .I1(sig00000a09),
    .I2(sig0000099f),
    .O(sig0000097e)
  );
  LUT4 #(
    .INIT ( 16'hEAAA ))
  blk00000a1a (
    .I0(sig00000808),
    .I1(sig0000098d),
    .I2(sig00000998),
    .I3(\NlwRenamedSig_OI_U0/i_synth/non_floating_point.arch_c.xfft_inst/control/cntrl/processing_state/ORS ),
    .O(sig000009c8)
  );
  LUT3 #(
    .INIT ( 8'hEA ))
  blk00000a1b (
    .I0(NlwRenamedSig_OI_xn_index[3]),
    .I1(sig00000a0a),
    .I2(sig000009aa),
    .O(sig0000096a)
  );
  LUT3 #(
    .INIT ( 8'hEA ))
  blk00000a1c (
    .I0(sig000009a6),
    .I1(sig00000a09),
    .I2(sig0000099f),
    .O(sig0000097d)
  );
  LUT4 #(
    .INIT ( 16'hEAAA ))
  blk00000a1d (
    .I0(sig00000809),
    .I1(sig0000098d),
    .I2(sig00000998),
    .I3(\NlwRenamedSig_OI_U0/i_synth/non_floating_point.arch_c.xfft_inst/control/cntrl/processing_state/ORS ),
    .O(sig000009c9)
  );
  LUT3 #(
    .INIT ( 8'hEA ))
  blk00000a1e (
    .I0(NlwRenamedSig_OI_xn_index[4]),
    .I1(sig00000a0a),
    .I2(sig000009aa),
    .O(sig00000969)
  );
  LUT3 #(
    .INIT ( 8'hEA ))
  blk00000a1f (
    .I0(sig000009a5),
    .I1(sig00000a09),
    .I2(sig0000099f),
    .O(sig0000097c)
  );
  LUT4 #(
    .INIT ( 16'hEAAA ))
  blk00000a20 (
    .I0(sig0000080a),
    .I1(sig0000098d),
    .I2(sig00000998),
    .I3(\NlwRenamedSig_OI_U0/i_synth/non_floating_point.arch_c.xfft_inst/control/cntrl/processing_state/ORS ),
    .O(sig000009ca)
  );
  LUT3 #(
    .INIT ( 8'hEA ))
  blk00000a21 (
    .I0(NlwRenamedSig_OI_xn_index[5]),
    .I1(sig00000a0a),
    .I2(sig000009aa),
    .O(sig00000968)
  );
  LUT3 #(
    .INIT ( 8'hEA ))
  blk00000a22 (
    .I0(sig000009a4),
    .I1(sig00000a09),
    .I2(sig0000099f),
    .O(sig0000097b)
  );
  LUT4 #(
    .INIT ( 16'hEAAA ))
  blk00000a23 (
    .I0(sig0000080b),
    .I1(sig0000098d),
    .I2(sig00000998),
    .I3(\NlwRenamedSig_OI_U0/i_synth/non_floating_point.arch_c.xfft_inst/control/cntrl/processing_state/ORS ),
    .O(sig000009cb)
  );
  LUT4 #(
    .INIT ( 16'hAEAA ))
  blk00000a24 (
    .I0(sig000009e0),
    .I1(sig00000003),
    .I2(sig00000998),
    .I3(\NlwRenamedSig_OI_U0/i_synth/non_floating_point.arch_c.xfft_inst/control/cntrl/processing_state/ORS ),
    .O(sig000009db)
  );
  LUT3 #(
    .INIT ( 8'hEA ))
  blk00000a25 (
    .I0(NlwRenamedSig_OI_xn_index[6]),
    .I1(sig00000a0a),
    .I2(sig000009aa),
    .O(sig00000967)
  );
  LUT3 #(
    .INIT ( 8'hEA ))
  blk00000a26 (
    .I0(sig000009a3),
    .I1(sig00000a09),
    .I2(sig0000099f),
    .O(sig0000097a)
  );
  LUT4 #(
    .INIT ( 16'hEAAA ))
  blk00000a27 (
    .I0(sig0000080c),
    .I1(sig0000098d),
    .I2(sig00000998),
    .I3(\NlwRenamedSig_OI_U0/i_synth/non_floating_point.arch_c.xfft_inst/control/cntrl/processing_state/ORS ),
    .O(sig000009cc)
  );
  LUT4 #(
    .INIT ( 16'hAEAA ))
  blk00000a28 (
    .I0(sig000009e1),
    .I1(sig00000003),
    .I2(sig00000998),
    .I3(\NlwRenamedSig_OI_U0/i_synth/non_floating_point.arch_c.xfft_inst/control/cntrl/processing_state/ORS ),
    .O(sig000009dc)
  );
  LUT4 #(
    .INIT ( 16'hEEEC ))
  blk00000a29 (
    .I0(sig000009ac),
    .I1(sig00000804),
    .I2(sig00000003),
    .I3(sig0000099b),
    .O(sig000009ed)
  );
  LUT3 #(
    .INIT ( 8'hEA ))
  blk00000a2a (
    .I0(NlwRenamedSig_OI_xn_index[7]),
    .I1(sig00000a0a),
    .I2(sig000009aa),
    .O(sig00000966)
  );
  LUT3 #(
    .INIT ( 8'hEA ))
  blk00000a2b (
    .I0(sig000009a2),
    .I1(sig00000a09),
    .I2(sig0000099f),
    .O(sig00000979)
  );
  LUT4 #(
    .INIT ( 16'hEAAA ))
  blk00000a2c (
    .I0(sig0000080d),
    .I1(sig0000098d),
    .I2(sig00000998),
    .I3(\NlwRenamedSig_OI_U0/i_synth/non_floating_point.arch_c.xfft_inst/control/cntrl/processing_state/ORS ),
    .O(sig000009cd)
  );
  LUT4 #(
    .INIT ( 16'hAEAA ))
  blk00000a2d (
    .I0(sig000009e2),
    .I1(sig00000003),
    .I2(sig00000998),
    .I3(\NlwRenamedSig_OI_U0/i_synth/non_floating_point.arch_c.xfft_inst/control/cntrl/processing_state/ORS ),
    .O(sig000009dd)
  );
  LUT4 #(
    .INIT ( 16'hFFA8 ))
  blk00000a2e (
    .I0(sig000009ac),
    .I1(sig0000099b),
    .I2(sig00000003),
    .I3(sig00000805),
    .O(sig000009ee)
  );
  LUT2 #(
    .INIT ( 4'h1 ))
  blk00000a2f (
    .I0(sig0000001f),
    .I1(sig0000001e),
    .O(sig00000a08)
  );
  LUT6 #(
    .INIT ( 64'h55AA55AA56AA55AA ))
  blk00000a30 (
    .I0(sig00000020),
    .I1(sig0000001d),
    .I2(sig0000001c),
    .I3(sig00000042),
    .I4(sig00000a08),
    .I5(sig0000051a),
    .O(sig00000523)
  );
  LUT3 #(
    .INIT ( 8'hF8 ))
  blk00000a31 (
    .I0(\NlwRenamedSig_OI_U0/i_synth/non_floating_point.arch_c.xfft_inst/control/cntrl/loading_state/ORS ),
    .I1(sig000009aa),
    .I2(NlwRenamedSig_OI_xn_index[8]),
    .O(sig00000965)
  );
  LUT3 #(
    .INIT ( 8'hF8 ))
  blk00000a32 (
    .I0(sig000007f9),
    .I1(sig0000099f),
    .I2(sig000009a1),
    .O(sig00000978)
  );
  LUT4 #(
    .INIT ( 16'hEAAA ))
  blk00000a33 (
    .I0(sig0000080e),
    .I1(sig00000998),
    .I2(\NlwRenamedSig_OI_U0/i_synth/non_floating_point.arch_c.xfft_inst/control/cntrl/processing_state/ORS ),
    .I3(sig0000098d),
    .O(sig000009ce)
  );
  LUT4 #(
    .INIT ( 16'hAEAA ))
  blk00000a34 (
    .I0(sig000009e3),
    .I1(\NlwRenamedSig_OI_U0/i_synth/non_floating_point.arch_c.xfft_inst/control/cntrl/processing_state/ORS ),
    .I2(sig00000998),
    .I3(sig00000003),
    .O(sig000009de)
  );
  LUT4 #(
    .INIT ( 16'hFFA8 ))
  blk00000a35 (
    .I0(sig000009ac),
    .I1(sig0000099b),
    .I2(sig00000003),
    .I3(sig00000806),
    .O(sig000009ef)
  );
  LUT5 #(
    .INIT ( 32'h1B1B1B00 ))
  blk00000a36 (
    .I0(sig0000099a),
    .I1(start),
    .I2(unload),
    .I3(sig00000999),
    .I4(sig0000099e),
    .O(sig000009fd)
  );
  LUT3 #(
    .INIT ( 8'h80 ))
  blk00000a37 (
    .I0(sig000009ad),
    .I1(\NlwRenamedSig_OI_U0/i_synth/non_floating_point.arch_c.xfft_inst/control/cntrl/processing_state/ORS ),
    .I2(sig000009ac),
    .O(sig00000a02)
  );
  LUT3 #(
    .INIT ( 8'h54 ))
  blk00000a38 (
    .I0(sig0000098d),
    .I1(sig00000998),
    .I2(sig00000003),
    .O(sig000009fe)
  );
  LUT2 #(
    .INIT ( 4'h8 ))
  blk00000a39 (
    .I0(sig000007f9),
    .I1(sig000009a0),
    .O(sig00000a03)
  );
  LUT2 #(
    .INIT ( 4'h8 ))
  blk00000a3a (
    .I0(\NlwRenamedSig_OI_U0/i_synth/non_floating_point.arch_c.xfft_inst/control/cntrl/loading_state/ORS ),
    .I1(sig000009ab),
    .O(sig00000a04)
  );
  LUT3 #(
    .INIT ( 8'h54 ))
  blk00000a3b (
    .I0(\NlwRenamedSig_OI_U0/i_synth/non_floating_point.arch_c.xfft_inst/control/cntrl/process_state_r ),
    .I1(\NlwRenamedSig_OI_U0/i_synth/non_floating_point.arch_c.xfft_inst/control/cntrl/processing_state/ORS ),
    .I2(sig0000099b),
    .O(sig00000a06)
  );
  LUT6 #(
    .INIT ( 64'h5555555540404000 ))
  blk00000a3c (
    .I0(sig0000099f),
    .I1(sig0000099a),
    .I2(unload),
    .I3(sig0000099c),
    .I4(sig00000999),
    .I5(sig000007f9),
    .O(sig00000a07)
  );
  LUT5 #(
    .INIT ( 32'hFF808080 ))
  blk00000a3d (
    .I0(\NlwRenamedSig_OI_U0/i_synth/non_floating_point.arch_c.xfft_inst/control/cntrl/processing_state/ORS ),
    .I1(sig000009ac),
    .I2(sig000009ad),
    .I3(sig000009a0),
    .I4(sig000007f9),
    .O(sig0000098a)
  );
  LUT4 #(
    .INIT ( 16'h5540 ))
  blk00000a3e (
    .I0(sig000009a0),
    .I1(sig000009ac),
    .I2(sig000009ad),
    .I3(sig0000099a),
    .O(sig00000a01)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000a3f (
    .C(clk),
    .D(sig00000a07),
    .Q(sig00000a09)
  );
  FD #(
    .INIT ( 1'b0 ))
  blk00000a40 (
    .C(clk),
    .D(sig00000a05),
    .Q(sig00000a0a)
  );
  INV   blk00000a41 (
    .I(sig0000021e),
    .O(sig000006a2)
  );
  INV   blk00000a42 (
    .I(sig00000208),
    .O(sig000006ab)
  );
  INV   blk00000a43 (
    .I(sig000001f2),
    .O(sig000006b4)
  );
  INV   blk00000a44 (
    .I(sig000001dc),
    .O(sig000006bd)
  );
  INV   blk00000a45 (
    .I(sig000008cf),
    .O(sig000008bc)
  );
  INV   blk00000a46 (
    .I(sig00000806),
    .O(sig000008bd)
  );
  RAMB8BWER #(
    .INIT_00 ( 256'h002F002C002900260022001F001C0019001600130010000D0009000600030000 ),
    .INIT_01 ( 256'h005F005C0059005600530050004D004A004700440041003E003B003800350032 ),
    .INIT_02 ( 256'h008C0089008600840081007E007B0079007600730070006D006B006800650062 ),
    .INIT_03 ( 256'h00B300B100AE00AC00AA00A700A500A200A0009D009B0098009600930091008E ),
    .INIT_04 ( 256'h00D300D100CF00CE00CC00CA00C800C600C400C200C000BE00BC00B900B700B5 ),
    .INIT_05 ( 256'h00EB00EA00E900E700E600E500E300E200E000DF00DD00DC00DA00D800D700D5 ),
    .INIT_06 ( 256'h00FA00FA00F900F800F800F700F600F500F400F300F200F100F000EF00EE00ED ),
    .INIT_07 ( 256'h0100010001000100010000FF00FF00FF00FE00FE00FE00FD00FD00FC00FC00FB ),
    .INIT_08 ( 256'h00FC00FC00FD00FD00FE00FE00FE00FF00FF00FF010001000100010001000100 ),
    .INIT_09 ( 256'h00EE00EF00F000F100F200F300F400F500F600F700F800F800F900FA00FA00FB ),
    .INIT_0A ( 256'h00D700D800DA00DC00DD00DF00E000E200E300E500E600E700E900EA00EB00ED ),
    .INIT_0B ( 256'h00B700B900BC00BE00C000C200C400C600C800CA00CC00CE00CF00D100D300D5 ),
    .INIT_0C ( 256'h0091009300960098009B009D00A000A200A500A700AA00AC00AE00B100B300B5 ),
    .INIT_0D ( 256'h00650068006B006D0070007300760079007B007E0081008400860089008C008E ),
    .INIT_0E ( 256'h00350038003B003E004100440047004A004D0050005300560059005C005F0062 ),
    .INIT_0F ( 256'h000300060009000D0010001300160019001C001F002200260029002C002F0032 ),
    .INIT_10 ( 256'h00FC00FC00FD00FD00FE00FE00FE00FF00FF00FF010001000100010001000100 ),
    .INIT_11 ( 256'h00EE00EF00F000F100F200F300F400F500F600F700F800F800F900FA00FA00FB ),
    .INIT_12 ( 256'h00D700D800DA00DC00DD00DF00E000E200E300E500E600E700E900EA00EB00ED ),
    .INIT_13 ( 256'h00B700B900BC00BE00C000C200C400C600C800CA00CC00CE00CF00D100D300D5 ),
    .INIT_14 ( 256'h0091009300960098009B009D00A000A200A500A700AA00AC00AE00B100B300B5 ),
    .INIT_15 ( 256'h00650068006B006D0070007300760079007B007E0081008400860089008C008E ),
    .INIT_16 ( 256'h00350038003B003E004100440047004A004D0050005300560059005C005F0062 ),
    .INIT_17 ( 256'h000300060009000D0010001300160019001C001F002200260029002C002F0032 ),
    .INIT_18 ( 256'h03D103D403D703DA03DE03E103E403E703EA03ED03F003F303F703FA03FD0000 ),
    .INIT_19 ( 256'h03A103A403A703AA03AD03B003B303B603B903BC03BF03C203C503C803CB03CE ),
    .INIT_1A ( 256'h03740377037A037C037F038203850387038A038D0390039303950398039B039E ),
    .INIT_1B ( 256'h034D034F0352035403560359035B035E0360036303650368036A036D036F0372 ),
    .INIT_1C ( 256'h032D032F03310332033403360338033A033C033E03400342034403470349034B ),
    .INIT_1D ( 256'h0315031603170319031A031B031D031E0320032103230324032603280329032B ),
    .INIT_1E ( 256'h030603060307030803080309030A030B030C030D030E030F0310031103120313 ),
    .INIT_1F ( 256'h0300030003000300030003010301030103020302030203030303030403040305 ),
    .INIT_A ( 18'h00000 ),
    .INIT_B ( 18'h00000 ),
    .WRITE_MODE_A ( "WRITE_FIRST" ),
    .WRITE_MODE_B ( "WRITE_FIRST" ),
    .DATA_WIDTH_A ( 18 ),
    .DATA_WIDTH_B ( 18 ),
    .DOA_REG ( 1 ),
    .DOB_REG ( 1 ),
    .EN_RSTRAM_A ( "TRUE" ),
    .EN_RSTRAM_B ( "TRUE" ),
    .INITP_00 ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INITP_01 ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INITP_02 ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INITP_03 ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .RAM_MODE ( "TDP" ),
    .RST_PRIORITY_A ( "CE" ),
    .RST_PRIORITY_B ( "CE" ),
    .RSTTYPE ( "SYNC" ),
    .SRVAL_A ( 18'h00000 ),
    .SRVAL_B ( 18'h00000 ),
    .INIT_FILE ( "NONE" ),
    .SIM_COLLISION_CHECK ( "ALL" ))
  blk00000a47 (
    .RSTBRST(sig00000002),
    .ENBRDEN(sig00000001),
    .REGCEA(sig00000001),
    .ENAWREN(sig00000001),
    .CLKAWRCLK(clk),
    .CLKBRDCLK(clk),
    .REGCEBREGCE(sig00000001),
    .RSTA(sig00000002),
    .WEAWEL({sig00000002, sig00000002}),
    .DOADO({\NLW_blk00000a47_DOADO<15>_UNCONNECTED , \NLW_blk00000a47_DOADO<14>_UNCONNECTED , \NLW_blk00000a47_DOADO<13>_UNCONNECTED ,
\NLW_blk00000a47_DOADO<12>_UNCONNECTED , \NLW_blk00000a47_DOADO<11>_UNCONNECTED , \NLW_blk00000a47_DOADO<10>_UNCONNECTED , sig00000903, sig00000902,
sig00000901, sig00000900, sig000008ff, sig000008fe, sig000008fd, sig000008fc, sig000008fb, sig000008fa}),
    .DOPADOP({\NLW_blk00000a47_DOPADOP<1>_UNCONNECTED , \NLW_blk00000a47_DOPADOP<0>_UNCONNECTED }),
    .DOPBDOP({\NLW_blk00000a47_DOPBDOP<1>_UNCONNECTED , \NLW_blk00000a47_DOPBDOP<0>_UNCONNECTED }),
    .WEBWEU({sig00000002, sig00000002}),
    .ADDRAWRADDR({sig00000002, sig00000823, sig00000822, sig00000821, sig00000820, sig0000081f, sig0000081e, sig0000081d, sig0000081c,
\NLW_blk00000a47_ADDRAWRADDR<3>_UNCONNECTED , \NLW_blk00000a47_ADDRAWRADDR<2>_UNCONNECTED , \NLW_blk00000a47_ADDRAWRADDR<1>_UNCONNECTED ,
\NLW_blk00000a47_ADDRAWRADDR<0>_UNCONNECTED }),
    .DIPBDIP({\NLW_blk00000a47_DIPBDIP<1>_UNCONNECTED , \NLW_blk00000a47_DIPBDIP<0>_UNCONNECTED }),
    .DIBDI({\NLW_blk00000a47_DIBDI<15>_UNCONNECTED , \NLW_blk00000a47_DIBDI<14>_UNCONNECTED , \NLW_blk00000a47_DIBDI<13>_UNCONNECTED ,
\NLW_blk00000a47_DIBDI<12>_UNCONNECTED , \NLW_blk00000a47_DIBDI<11>_UNCONNECTED , \NLW_blk00000a47_DIBDI<10>_UNCONNECTED ,
\NLW_blk00000a47_DIBDI<9>_UNCONNECTED , \NLW_blk00000a47_DIBDI<8>_UNCONNECTED , \NLW_blk00000a47_DIBDI<7>_UNCONNECTED ,
\NLW_blk00000a47_DIBDI<6>_UNCONNECTED , \NLW_blk00000a47_DIBDI<5>_UNCONNECTED , \NLW_blk00000a47_DIBDI<4>_UNCONNECTED ,
\NLW_blk00000a47_DIBDI<3>_UNCONNECTED , \NLW_blk00000a47_DIBDI<2>_UNCONNECTED , \NLW_blk00000a47_DIBDI<1>_UNCONNECTED ,
\NLW_blk00000a47_DIBDI<0>_UNCONNECTED }),
    .DIADI({sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002,
sig00000002, sig00000002, sig00000002, sig00000002, sig00000002, sig00000002}),
    .ADDRBRDADDR({sig00000001, sig00000823, sig00000822, sig00000821, sig00000820, sig0000081f, sig0000081e, sig0000081d, sig0000081c,
\NLW_blk00000a47_ADDRBRDADDR<3>_UNCONNECTED , \NLW_blk00000a47_ADDRBRDADDR<2>_UNCONNECTED , \NLW_blk00000a47_ADDRBRDADDR<1>_UNCONNECTED ,
\NLW_blk00000a47_ADDRBRDADDR<0>_UNCONNECTED }),
    .DOBDO({\NLW_blk00000a47_DOBDO<15>_UNCONNECTED , \NLW_blk00000a47_DOBDO<14>_UNCONNECTED , \NLW_blk00000a47_DOBDO<13>_UNCONNECTED ,
\NLW_blk00000a47_DOBDO<12>_UNCONNECTED , \NLW_blk00000a47_DOBDO<11>_UNCONNECTED , \NLW_blk00000a47_DOBDO<10>_UNCONNECTED , sig000008f9, sig000008f8,
sig000008f7, sig000008f6, sig000008f5, sig000008f4, sig000008f3, sig000008f2, sig000008f1, sig000008f0}),
    .DIPADIP({sig00000002, sig00000002})
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000a48 (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig00000472),
    .Q(sig00000a0b),
    .Q15(NLW_blk00000a48_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000a49 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000a0b),
    .Q(sig000004a3)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000a4a (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig00000471),
    .Q(sig00000a0c),
    .Q15(NLW_blk00000a4a_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000a4b (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000a0c),
    .Q(sig000004a2)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000a4c (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig00000470),
    .Q(sig00000a0d),
    .Q15(NLW_blk00000a4c_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000a4d (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000a0d),
    .Q(sig000004a1)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000a4e (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig0000046f),
    .Q(sig00000a0e),
    .Q15(NLW_blk00000a4e_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000a4f (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000a0e),
    .Q(sig0000030c)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000a50 (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig0000046e),
    .Q(sig00000a0f),
    .Q15(NLW_blk00000a50_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000a51 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000a0f),
    .Q(sig0000030d)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000a52 (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig0000046d),
    .Q(sig00000a10),
    .Q15(NLW_blk00000a52_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000a53 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000a10),
    .Q(sig0000030e)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000a54 (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig0000046c),
    .Q(sig00000a11),
    .Q15(NLW_blk00000a54_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000a55 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000a11),
    .Q(sig0000030f)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000a56 (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig0000046b),
    .Q(sig00000a12),
    .Q15(NLW_blk00000a56_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000a57 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000a12),
    .Q(sig00000310)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000a58 (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig0000046a),
    .Q(sig00000a13),
    .Q15(NLW_blk00000a58_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000a59 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000a13),
    .Q(sig00000311)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000a5a (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig00000469),
    .Q(sig00000a14),
    .Q15(NLW_blk00000a5a_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000a5b (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000a14),
    .Q(sig00000312)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000a5c (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig00000468),
    .Q(sig00000a15),
    .Q15(NLW_blk00000a5c_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000a5d (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000a15),
    .Q(sig00000313)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000a5e (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig00000467),
    .Q(sig00000a16),
    .Q15(NLW_blk00000a5e_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000a5f (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000a16),
    .Q(sig00000314)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000a60 (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig00000464),
    .Q(sig00000a17),
    .Q15(NLW_blk00000a60_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000a61 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000a17),
    .Q(sig00000317)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000a62 (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig00000466),
    .Q(sig00000a18),
    .Q15(NLW_blk00000a62_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000a63 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000a18),
    .Q(sig00000315)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000a64 (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig00000465),
    .Q(sig00000a19),
    .Q15(NLW_blk00000a64_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000a65 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000a19),
    .Q(sig00000316)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000a66 (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig00000463),
    .Q(sig00000a1a),
    .Q15(NLW_blk00000a66_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000a67 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000a1a),
    .Q(sig00000318)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000a68 (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig00000462),
    .Q(sig00000a1b),
    .Q15(NLW_blk00000a68_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000a69 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000a1b),
    .Q(sig00000319)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000a6a (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig00000461),
    .Q(sig00000a1c),
    .Q15(NLW_blk00000a6a_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000a6b (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000a1c),
    .Q(sig0000031a)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000a6c (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig00000460),
    .Q(sig00000a1d),
    .Q15(NLW_blk00000a6c_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000a6d (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000a1d),
    .Q(sig0000031b)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000a6e (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig00000473),
    .Q(sig00000a1e),
    .Q15(NLW_blk00000a6e_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000a6f (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000a1e),
    .Q(sig0000031c)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000a70 (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig00000486),
    .Q(sig00000a1f),
    .Q15(NLW_blk00000a70_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000a71 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000a1f),
    .Q(sig000004df)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000a72 (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig00000485),
    .Q(sig00000a20),
    .Q15(NLW_blk00000a72_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000a73 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000a20),
    .Q(sig000004de)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000a74 (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig00000484),
    .Q(sig00000a21),
    .Q15(NLW_blk00000a74_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000a75 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000a21),
    .Q(sig000004dd)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000a76 (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig00000483),
    .Q(sig00000a22),
    .Q15(NLW_blk00000a76_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000a77 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000a22),
    .Q(sig000004dc)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000a78 (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig00000482),
    .Q(sig00000a23),
    .Q15(NLW_blk00000a78_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000a79 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000a23),
    .Q(sig000004db)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000a7a (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig00000481),
    .Q(sig00000a24),
    .Q15(NLW_blk00000a7a_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000a7b (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000a24),
    .Q(sig000004da)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000a7c (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig00000480),
    .Q(sig00000a25),
    .Q15(NLW_blk00000a7c_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000a7d (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000a25),
    .Q(sig000004d9)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000a7e (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig0000047d),
    .Q(sig00000a26),
    .Q15(NLW_blk00000a7e_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000a7f (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000a26),
    .Q(sig000004d6)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000a80 (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig0000047f),
    .Q(sig00000a27),
    .Q15(NLW_blk00000a80_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000a81 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000a27),
    .Q(sig000004d8)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000a82 (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig0000047e),
    .Q(sig00000a28),
    .Q15(NLW_blk00000a82_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000a83 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000a28),
    .Q(sig000004d7)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000a84 (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig0000047c),
    .Q(sig00000a29),
    .Q15(NLW_blk00000a84_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000a85 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000a29),
    .Q(sig000004d5)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000a86 (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig0000047b),
    .Q(sig00000a2a),
    .Q15(NLW_blk00000a86_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000a87 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000a2a),
    .Q(sig000004d4)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000a88 (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig0000047a),
    .Q(sig00000a2b),
    .Q15(NLW_blk00000a88_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000a89 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000a2b),
    .Q(sig000004d3)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000a8a (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig00000479),
    .Q(sig00000a2c),
    .Q15(NLW_blk00000a8a_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000a8b (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000a2c),
    .Q(sig000004d2)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000a8c (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig00000478),
    .Q(sig00000a2d),
    .Q15(NLW_blk00000a8c_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000a8d (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000a2d),
    .Q(sig000004d1)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000a8e (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig00000477),
    .Q(sig00000a2e),
    .Q15(NLW_blk00000a8e_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000a8f (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000a2e),
    .Q(sig000004d0)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000a90 (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig00000476),
    .Q(sig00000a2f),
    .Q15(NLW_blk00000a90_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000a91 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000a2f),
    .Q(sig000004cf)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000a92 (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig00000475),
    .Q(sig00000a30),
    .Q15(NLW_blk00000a92_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000a93 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000a30),
    .Q(sig000004ce)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000a94 (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig00000474),
    .Q(sig00000a31),
    .Q15(NLW_blk00000a94_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000a95 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000a31),
    .Q(sig000004cd)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000a96 (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000003dc),
    .Q(sig00000a32),
    .Q15(NLW_blk00000a96_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000a97 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000a32),
    .Q(sig00000320)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000a98 (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000003e5),
    .Q(sig00000a33),
    .Q15(NLW_blk00000a98_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000a99 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000a33),
    .Q(sig00000329)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000a9a (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000003e6),
    .Q(sig00000a34),
    .Q15(NLW_blk00000a9a_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000a9b (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000a34),
    .Q(sig0000032a)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000a9c (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000003e9),
    .Q(sig00000a35),
    .Q15(NLW_blk00000a9c_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000a9d (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000a35),
    .Q(sig0000032d)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000a9e (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000003e7),
    .Q(sig00000a36),
    .Q15(NLW_blk00000a9e_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000a9f (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000a36),
    .Q(sig0000032b)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000aa0 (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000003e8),
    .Q(sig00000a37),
    .Q15(NLW_blk00000aa0_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000aa1 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000a37),
    .Q(sig0000032c)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000aa2 (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000003ea),
    .Q(sig00000a38),
    .Q15(NLW_blk00000aa2_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000aa3 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000a38),
    .Q(sig0000032e)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000aa4 (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000003eb),
    .Q(sig00000a39),
    .Q15(NLW_blk00000aa4_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000aa5 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000a39),
    .Q(sig0000032f)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000aa6 (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000003ec),
    .Q(sig00000a3a),
    .Q15(NLW_blk00000aa6_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000aa7 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000a3a),
    .Q(sig00000330)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000aa8 (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000003ed),
    .Q(sig00000a3b),
    .Q15(NLW_blk00000aa8_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000aa9 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000a3b),
    .Q(sig00000331)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000aaa (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000004e9),
    .Q(sig00000a3c),
    .Q15(NLW_blk00000aaa_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000aab (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000a3c),
    .Q(sig000004cb)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000aac (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000004e8),
    .Q(sig00000a3d),
    .Q15(NLW_blk00000aac_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000aad (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000a3d),
    .Q(sig000004ca)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000aae (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000004e7),
    .Q(sig00000a3e),
    .Q15(NLW_blk00000aae_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000aaf (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000a3e),
    .Q(sig000004c9)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000ab0 (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000004e6),
    .Q(sig00000a3f),
    .Q15(NLW_blk00000ab0_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000ab1 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000a3f),
    .Q(sig000004c8)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000ab2 (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000004e5),
    .Q(sig00000a40),
    .Q15(NLW_blk00000ab2_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000ab3 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000a40),
    .Q(sig000004c7)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000ab4 (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000004e4),
    .Q(sig00000a41),
    .Q15(NLW_blk00000ab4_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000ab5 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000a41),
    .Q(sig000004c6)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000ab6 (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000004e3),
    .Q(sig00000a42),
    .Q15(NLW_blk00000ab6_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000ab7 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000a42),
    .Q(sig000004c5)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000ab8 (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000004e2),
    .Q(sig00000a43),
    .Q15(NLW_blk00000ab8_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000ab9 (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000a43),
    .Q(sig000004c4)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000aba (
    .A0(sig00000002),
    .A1(sig00000002),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(NlwRenamedSig_OI_xn_index[8]),
    .Q(sig00000a44),
    .Q15(NLW_blk00000aba_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000abb (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000a44),
    .Q(sig00000862)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000abc (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000004e1),
    .Q(sig00000a45),
    .Q15(NLW_blk00000abc_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000abd (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000a45),
    .Q(sig000004c3)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  blk00000abe (
    .A0(sig00000002),
    .A1(sig00000001),
    .A2(sig00000002),
    .A3(sig00000002),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000004e0),
    .Q(sig00000a46),
    .Q15(NLW_blk00000abe_Q15_UNCONNECTED)
  );
  FDE #(
    .INIT ( 1'b0 ))
  blk00000abf (
    .C(clk),
    .CE(sig00000001),
    .D(sig00000a46),
    .Q(sig000004c2)
  );
  RAMB8BWER #(
    .DATA_WIDTH_A ( 36 ),
    .DATA_WIDTH_B ( 36 ),
    .DOA_REG ( 0 ),
    .DOB_REG ( 1 ),
    .EN_RSTRAM_A ( "FALSE" ),
    .EN_RSTRAM_B ( "FALSE" ),
    .INITP_00 ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INITP_01 ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INITP_02 ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INITP_03 ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_00 ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_01 ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_02 ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_03 ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_04 ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_05 ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_06 ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_07 ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_08 ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_09 ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_0A ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_0B ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_0C ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_0D ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_0E ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_0F ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_10 ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_11 ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_12 ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_13 ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_14 ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_15 ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_16 ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_17 ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_18 ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_19 ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_1A ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_1B ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_1C ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_1D ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_1E ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_1F ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_A ( 18'h00000 ),
    .INIT_B ( 18'h00000 ),
    .INIT_FILE ( "NONE" ),
    .RAM_MODE ( "SDP" ),
    .RSTTYPE ( "SYNC" ),
    .RST_PRIORITY_A ( "CE" ),
    .RST_PRIORITY_B ( "CE" ),
    .SIM_COLLISION_CHECK ( "GENERATE_X_ONLY" ),
    .SRVAL_A ( 18'h00000 ),
    .SRVAL_B ( 18'h00000 ),
    .WRITE_MODE_A ( "READ_FIRST" ),
    .WRITE_MODE_B ( "READ_FIRST" ))
  \blk00000003/blk0000002c  (
    .RSTBRST(\blk00000003/sig00000acd ),
    .ENBRDEN(sig00000001),
    .REGCEA(\blk00000003/sig00000acd ),
    .ENAWREN(sig00000001),
    .CLKAWRCLK(clk),
    .CLKBRDCLK(clk),
    .REGCEBREGCE(sig00000001),
    .RSTA(\blk00000003/sig00000acd ),
    .WEAWEL({sig00000009, sig00000009}),
    .DOADO({\NLW_blk00000003/blk0000002c_DOADO<15>_UNCONNECTED , \NLW_blk00000003/blk0000002c_DOADO<14>_UNCONNECTED ,
\NLW_blk00000003/blk0000002c_DOADO<13>_UNCONNECTED , \NLW_blk00000003/blk0000002c_DOADO<12>_UNCONNECTED ,
\NLW_blk00000003/blk0000002c_DOADO<11>_UNCONNECTED , \NLW_blk00000003/blk0000002c_DOADO<10>_UNCONNECTED ,
\NLW_blk00000003/blk0000002c_DOADO<9>_UNCONNECTED , \NLW_blk00000003/blk0000002c_DOADO<8>_UNCONNECTED ,
\NLW_blk00000003/blk0000002c_DOADO<7>_UNCONNECTED , \NLW_blk00000003/blk0000002c_DOADO<6>_UNCONNECTED ,
\NLW_blk00000003/blk0000002c_DOADO<5>_UNCONNECTED , \NLW_blk00000003/blk0000002c_DOADO<4>_UNCONNECTED ,
\NLW_blk00000003/blk0000002c_DOADO<3>_UNCONNECTED , \NLW_blk00000003/blk0000002c_DOADO<2>_UNCONNECTED , \blk00000003/sig00000aa5 ,
\blk00000003/sig00000aa6 }),
    .DOPADOP({\NLW_blk00000003/blk0000002c_DOPADOP<1>_UNCONNECTED , \NLW_blk00000003/blk0000002c_DOPADOP<0>_UNCONNECTED }),
    .DOPBDOP({\NLW_blk00000003/blk0000002c_DOPBDOP<1>_UNCONNECTED , \NLW_blk00000003/blk0000002c_DOPBDOP<0>_UNCONNECTED }),
    .WEBWEU({sig00000009, sig00000009}),
    .ADDRAWRADDR({sig00000030, sig0000002f, sig0000002e, sig0000002d, sig0000002c, sig0000002b, sig0000002a, sig00000029, \blk00000003/sig00000acd ,
\blk00000003/sig00000acd , \blk00000003/sig00000acd , \blk00000003/sig00000acd , \blk00000003/sig00000acd }),
    .DIPBDIP({\blk00000003/sig00000acd , \blk00000003/sig00000acd }),
    .DIBDI({\blk00000003/sig00000acd , \blk00000003/sig00000acd , \blk00000003/sig00000acd , \blk00000003/sig00000acd , \blk00000003/sig00000acd ,
\blk00000003/sig00000acd , \blk00000003/sig00000acd , \blk00000003/sig00000acd , \blk00000003/sig00000acd , \blk00000003/sig00000acd ,
\blk00000003/sig00000acd , \blk00000003/sig00000acd , \blk00000003/sig00000acd , \blk00000003/sig00000acd , \blk00000003/sig00000acd ,
\blk00000003/sig00000acd }),
    .DIADI({\blk00000003/sig00000acd , \blk00000003/sig00000acd , \blk00000003/sig00000acd , \blk00000003/sig00000acd , \blk00000003/sig00000acd ,
\blk00000003/sig00000acd , \blk00000003/sig00000acd , \blk00000003/sig00000acd , \blk00000003/sig00000acd , \blk00000003/sig00000acd ,
\blk00000003/sig00000acd , \blk00000003/sig00000acd , \blk00000003/sig00000acd , \blk00000003/sig00000acd , sig000000b4, sig000000b3}),
    .ADDRBRDADDR({sig00000028, sig00000027, sig00000026, sig00000025, sig00000024, sig00000023, sig00000022, sig00000021, \blk00000003/sig00000acd ,
\blk00000003/sig00000acd , \blk00000003/sig00000acd , \blk00000003/sig00000acd , \blk00000003/sig00000acd }),
    .DOBDO({\NLW_blk00000003/blk0000002c_DOBDO<15>_UNCONNECTED , \NLW_blk00000003/blk0000002c_DOBDO<14>_UNCONNECTED ,
\NLW_blk00000003/blk0000002c_DOBDO<13>_UNCONNECTED , \NLW_blk00000003/blk0000002c_DOBDO<12>_UNCONNECTED ,
\NLW_blk00000003/blk0000002c_DOBDO<11>_UNCONNECTED , \NLW_blk00000003/blk0000002c_DOBDO<10>_UNCONNECTED ,
\NLW_blk00000003/blk0000002c_DOBDO<9>_UNCONNECTED , \NLW_blk00000003/blk0000002c_DOBDO<8>_UNCONNECTED ,
\NLW_blk00000003/blk0000002c_DOBDO<7>_UNCONNECTED , \NLW_blk00000003/blk0000002c_DOBDO<6>_UNCONNECTED ,
\NLW_blk00000003/blk0000002c_DOBDO<5>_UNCONNECTED , \NLW_blk00000003/blk0000002c_DOBDO<4>_UNCONNECTED ,
\NLW_blk00000003/blk0000002c_DOBDO<3>_UNCONNECTED , \NLW_blk00000003/blk0000002c_DOBDO<2>_UNCONNECTED ,
\NLW_blk00000003/blk0000002c_DOBDO<1>_UNCONNECTED , \NLW_blk00000003/blk0000002c_DOBDO<0>_UNCONNECTED }),
    .DIPADIP({\blk00000003/sig00000acd , \blk00000003/sig00000acd })
  );
  RAMB8BWER #(
    .DATA_WIDTH_A ( 36 ),
    .DATA_WIDTH_B ( 36 ),
    .DOA_REG ( 0 ),
    .DOB_REG ( 1 ),
    .EN_RSTRAM_A ( "FALSE" ),
    .EN_RSTRAM_B ( "FALSE" ),
    .INITP_00 ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INITP_01 ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INITP_02 ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INITP_03 ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_00 ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_01 ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_02 ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_03 ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_04 ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_05 ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_06 ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_07 ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_08 ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_09 ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_0A ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_0B ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_0C ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_0D ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_0E ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_0F ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_10 ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_11 ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_12 ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_13 ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_14 ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_15 ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_16 ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_17 ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_18 ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_19 ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_1A ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_1B ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_1C ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_1D ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_1E ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_1F ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_A ( 18'h00000 ),
    .INIT_B ( 18'h00000 ),
    .INIT_FILE ( "NONE" ),
    .RAM_MODE ( "SDP" ),
    .RSTTYPE ( "SYNC" ),
    .RST_PRIORITY_A ( "CE" ),
    .RST_PRIORITY_B ( "CE" ),
    .SIM_COLLISION_CHECK ( "GENERATE_X_ONLY" ),
    .SRVAL_A ( 18'h00000 ),
    .SRVAL_B ( 18'h00000 ),
    .WRITE_MODE_A ( "READ_FIRST" ),
    .WRITE_MODE_B ( "READ_FIRST" ))
  \blk00000003/blk0000002b  (
    .RSTBRST(\blk00000003/sig00000acd ),
    .ENBRDEN(sig00000001),
    .REGCEA(\blk00000003/sig00000acd ),
    .ENAWREN(sig00000001),
    .CLKAWRCLK(clk),
    .CLKBRDCLK(clk),
    .REGCEBREGCE(sig00000001),
    .RSTA(\blk00000003/sig00000acd ),
    .WEAWEL({sig00000009, sig00000009}),
    .DOADO({\blk00000003/sig00000a89 , \blk00000003/sig00000a8a , \blk00000003/sig00000a8b , \blk00000003/sig00000a8c , \blk00000003/sig00000a8d ,
\blk00000003/sig00000a8e , \blk00000003/sig00000a8f , \blk00000003/sig00000a90 , \blk00000003/sig00000a81 , \blk00000003/sig00000a82 ,
\blk00000003/sig00000a83 , \blk00000003/sig00000a84 , \blk00000003/sig00000a85 , \blk00000003/sig00000a86 , \blk00000003/sig00000a87 ,
\blk00000003/sig00000a88 }),
    .DOPADOP({\blk00000003/sig00000aa2 , \blk00000003/sig00000aa1 }),
    .DOPBDOP({\blk00000003/sig00000aa4 , \blk00000003/sig00000aa3 }),
    .WEBWEU({sig00000009, sig00000009}),
    .ADDRAWRADDR({sig00000030, sig0000002f, sig0000002e, sig0000002d, sig0000002c, sig0000002b, sig0000002a, sig00000029, \blk00000003/sig00000acd ,
\blk00000003/sig00000acd , \blk00000003/sig00000acd , \blk00000003/sig00000acd , \blk00000003/sig00000acd }),
    .DIPBDIP({sig000000b2, sig000000a9}),
    .DIBDI({sig000000b1, sig000000b0, sig000000af, sig000000ae, sig000000ad, sig000000ac, sig000000ab, sig000000aa, sig000000a8, sig000000a7,
sig000000a6, sig000000a5, sig000000a4, sig000000a3, sig000000a2, sig000000a1}),
    .DIADI({sig0000009f, sig0000009e, sig0000009d, sig0000009c, sig0000009b, sig0000009a, sig00000099, sig00000098, sig00000096, sig00000095,
sig00000094, sig00000093, sig00000092, sig00000091, sig00000090, sig0000008f}),
    .ADDRBRDADDR({sig00000028, sig00000027, sig00000026, sig00000025, sig00000024, sig00000023, sig00000022, sig00000021, \blk00000003/sig00000acd ,
\blk00000003/sig00000acd , \blk00000003/sig00000acd , \blk00000003/sig00000acd , \blk00000003/sig00000acd }),
    .DOBDO({\blk00000003/sig00000a99 , \blk00000003/sig00000a9a , \blk00000003/sig00000a9b , \blk00000003/sig00000a9c , \blk00000003/sig00000a9d ,
\blk00000003/sig00000a9e , \blk00000003/sig00000a9f , \blk00000003/sig00000aa0 , \blk00000003/sig00000a91 , \blk00000003/sig00000a92 ,
\blk00000003/sig00000a93 , \blk00000003/sig00000a94 , \blk00000003/sig00000a95 , \blk00000003/sig00000a96 , \blk00000003/sig00000a97 ,
\blk00000003/sig00000a98 }),
    .DIPADIP({sig000000a0, sig00000097})
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000003/blk0000002a  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk00000003/sig00000aa5 ),
    .Q(sig00000172)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000003/blk00000029  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk00000003/sig00000aa6 ),
    .Q(sig00000171)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000003/blk00000028  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk00000003/sig00000aa4 ),
    .Q(sig00000170)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000003/blk00000027  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk00000003/sig00000a99 ),
    .Q(sig0000016f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000003/blk00000026  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk00000003/sig00000a9a ),
    .Q(sig0000016e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000003/blk00000025  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk00000003/sig00000a9b ),
    .Q(sig0000016d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000003/blk00000024  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk00000003/sig00000a9c ),
    .Q(sig0000016c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000003/blk00000023  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk00000003/sig00000a9d ),
    .Q(sig0000016b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000003/blk00000022  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk00000003/sig00000a9e ),
    .Q(sig0000016a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000003/blk00000021  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk00000003/sig00000a9f ),
    .Q(sig00000169)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000003/blk00000020  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk00000003/sig00000aa0 ),
    .Q(sig00000168)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000003/blk0000001f  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk00000003/sig00000aa3 ),
    .Q(sig00000167)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000003/blk0000001e  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk00000003/sig00000a91 ),
    .Q(sig00000166)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000003/blk0000001d  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk00000003/sig00000a92 ),
    .Q(sig00000165)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000003/blk0000001c  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk00000003/sig00000a93 ),
    .Q(sig00000164)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000003/blk0000001b  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk00000003/sig00000a94 ),
    .Q(sig00000163)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000003/blk0000001a  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk00000003/sig00000a95 ),
    .Q(sig00000162)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000003/blk00000019  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk00000003/sig00000a96 ),
    .Q(sig00000161)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000003/blk00000018  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk00000003/sig00000a97 ),
    .Q(sig00000160)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000003/blk00000017  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk00000003/sig00000a98 ),
    .Q(sig0000015f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000003/blk00000016  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk00000003/sig00000aa2 ),
    .Q(sig0000015e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000003/blk00000015  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk00000003/sig00000a89 ),
    .Q(sig0000015d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000003/blk00000014  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk00000003/sig00000a8a ),
    .Q(sig0000015c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000003/blk00000013  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk00000003/sig00000a8b ),
    .Q(sig0000015b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000003/blk00000012  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk00000003/sig00000a8c ),
    .Q(sig0000015a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000003/blk00000011  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk00000003/sig00000a8d ),
    .Q(sig00000159)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000003/blk00000010  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk00000003/sig00000a8e ),
    .Q(sig00000158)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000003/blk0000000f  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk00000003/sig00000a8f ),
    .Q(sig00000157)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000003/blk0000000e  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk00000003/sig00000a90 ),
    .Q(sig00000156)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000003/blk0000000d  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk00000003/sig00000aa1 ),
    .Q(sig00000155)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000003/blk0000000c  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk00000003/sig00000a81 ),
    .Q(sig00000154)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000003/blk0000000b  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk00000003/sig00000a82 ),
    .Q(sig00000153)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000003/blk0000000a  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk00000003/sig00000a83 ),
    .Q(sig00000152)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000003/blk00000009  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk00000003/sig00000a84 ),
    .Q(sig00000151)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000003/blk00000008  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk00000003/sig00000a85 ),
    .Q(sig00000150)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000003/blk00000007  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk00000003/sig00000a86 ),
    .Q(sig0000014f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000003/blk00000006  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk00000003/sig00000a87 ),
    .Q(sig0000014e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000003/blk00000005  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk00000003/sig00000a88 ),
    .Q(sig0000014d)
  );
  GND   \blk00000003/blk00000004  (
    .G(\blk00000003/sig00000acd )
  );
  RAMB8BWER #(
    .DATA_WIDTH_A ( 36 ),
    .DATA_WIDTH_B ( 36 ),
    .DOA_REG ( 0 ),
    .DOB_REG ( 1 ),
    .EN_RSTRAM_A ( "FALSE" ),
    .EN_RSTRAM_B ( "FALSE" ),
    .INITP_00 ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INITP_01 ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INITP_02 ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INITP_03 ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_00 ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_01 ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_02 ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_03 ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_04 ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_05 ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_06 ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_07 ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_08 ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_09 ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_0A ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_0B ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_0C ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_0D ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_0E ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_0F ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_10 ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_11 ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_12 ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_13 ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_14 ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_15 ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_16 ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_17 ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_18 ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_19 ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_1A ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_1B ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_1C ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_1D ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_1E ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_1F ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_A ( 18'h00000 ),
    .INIT_B ( 18'h00000 ),
    .INIT_FILE ( "NONE" ),
    .RAM_MODE ( "SDP" ),
    .RSTTYPE ( "SYNC" ),
    .RST_PRIORITY_A ( "CE" ),
    .RST_PRIORITY_B ( "CE" ),
    .SIM_COLLISION_CHECK ( "GENERATE_X_ONLY" ),
    .SRVAL_A ( 18'h00000 ),
    .SRVAL_B ( 18'h00000 ),
    .WRITE_MODE_A ( "READ_FIRST" ),
    .WRITE_MODE_B ( "READ_FIRST" ))
  \blk0000002d/blk00000056  (
    .RSTBRST(\blk0000002d/sig00000b54 ),
    .ENBRDEN(sig00000001),
    .REGCEA(\blk0000002d/sig00000b54 ),
    .ENAWREN(sig00000001),
    .CLKAWRCLK(clk),
    .CLKBRDCLK(clk),
    .REGCEBREGCE(sig00000001),
    .RSTA(\blk0000002d/sig00000b54 ),
    .WEAWEL({sig0000000a, sig0000000a}),
    .DOADO({\NLW_blk0000002d/blk00000056_DOADO<15>_UNCONNECTED , \NLW_blk0000002d/blk00000056_DOADO<14>_UNCONNECTED ,
\NLW_blk0000002d/blk00000056_DOADO<13>_UNCONNECTED , \NLW_blk0000002d/blk00000056_DOADO<12>_UNCONNECTED ,
\NLW_blk0000002d/blk00000056_DOADO<11>_UNCONNECTED , \NLW_blk0000002d/blk00000056_DOADO<10>_UNCONNECTED ,
\NLW_blk0000002d/blk00000056_DOADO<9>_UNCONNECTED , \NLW_blk0000002d/blk00000056_DOADO<8>_UNCONNECTED ,
\NLW_blk0000002d/blk00000056_DOADO<7>_UNCONNECTED , \NLW_blk0000002d/blk00000056_DOADO<6>_UNCONNECTED ,
\NLW_blk0000002d/blk00000056_DOADO<5>_UNCONNECTED , \NLW_blk0000002d/blk00000056_DOADO<4>_UNCONNECTED ,
\NLW_blk0000002d/blk00000056_DOADO<3>_UNCONNECTED , \NLW_blk0000002d/blk00000056_DOADO<2>_UNCONNECTED , \blk0000002d/sig00000b2c ,
\blk0000002d/sig00000b2d }),
    .DOPADOP({\NLW_blk0000002d/blk00000056_DOPADOP<1>_UNCONNECTED , \NLW_blk0000002d/blk00000056_DOPADOP<0>_UNCONNECTED }),
    .DOPBDOP({\NLW_blk0000002d/blk00000056_DOPBDOP<1>_UNCONNECTED , \NLW_blk0000002d/blk00000056_DOPBDOP<0>_UNCONNECTED }),
    .WEBWEU({sig0000000a, sig0000000a}),
    .ADDRAWRADDR({sig00000040, sig0000003f, sig0000003e, sig0000003d, sig0000003c, sig0000003b, sig0000003a, sig00000039, \blk0000002d/sig00000b54 ,
\blk0000002d/sig00000b54 , \blk0000002d/sig00000b54 , \blk0000002d/sig00000b54 , \blk0000002d/sig00000b54 }),
    .DIPBDIP({\blk0000002d/sig00000b54 , \blk0000002d/sig00000b54 }),
    .DIBDI({\blk0000002d/sig00000b54 , \blk0000002d/sig00000b54 , \blk0000002d/sig00000b54 , \blk0000002d/sig00000b54 , \blk0000002d/sig00000b54 ,
\blk0000002d/sig00000b54 , \blk0000002d/sig00000b54 , \blk0000002d/sig00000b54 , \blk0000002d/sig00000b54 , \blk0000002d/sig00000b54 ,
\blk0000002d/sig00000b54 , \blk0000002d/sig00000b54 , \blk0000002d/sig00000b54 , \blk0000002d/sig00000b54 , \blk0000002d/sig00000b54 ,
\blk0000002d/sig00000b54 }),
    .DIADI({\blk0000002d/sig00000b54 , \blk0000002d/sig00000b54 , \blk0000002d/sig00000b54 , \blk0000002d/sig00000b54 , \blk0000002d/sig00000b54 ,
\blk0000002d/sig00000b54 , \blk0000002d/sig00000b54 , \blk0000002d/sig00000b54 , \blk0000002d/sig00000b54 , \blk0000002d/sig00000b54 ,
\blk0000002d/sig00000b54 , \blk0000002d/sig00000b54 , \blk0000002d/sig00000b54 , \blk0000002d/sig00000b54 , sig000000da, sig000000d9}),
    .ADDRBRDADDR({sig00000038, sig00000037, sig00000036, sig00000035, sig00000034, sig00000033, sig00000032, sig00000031, \blk0000002d/sig00000b54 ,
\blk0000002d/sig00000b54 , \blk0000002d/sig00000b54 , \blk0000002d/sig00000b54 , \blk0000002d/sig00000b54 }),
    .DOBDO({\NLW_blk0000002d/blk00000056_DOBDO<15>_UNCONNECTED , \NLW_blk0000002d/blk00000056_DOBDO<14>_UNCONNECTED ,
\NLW_blk0000002d/blk00000056_DOBDO<13>_UNCONNECTED , \NLW_blk0000002d/blk00000056_DOBDO<12>_UNCONNECTED ,
\NLW_blk0000002d/blk00000056_DOBDO<11>_UNCONNECTED , \NLW_blk0000002d/blk00000056_DOBDO<10>_UNCONNECTED ,
\NLW_blk0000002d/blk00000056_DOBDO<9>_UNCONNECTED , \NLW_blk0000002d/blk00000056_DOBDO<8>_UNCONNECTED ,
\NLW_blk0000002d/blk00000056_DOBDO<7>_UNCONNECTED , \NLW_blk0000002d/blk00000056_DOBDO<6>_UNCONNECTED ,
\NLW_blk0000002d/blk00000056_DOBDO<5>_UNCONNECTED , \NLW_blk0000002d/blk00000056_DOBDO<4>_UNCONNECTED ,
\NLW_blk0000002d/blk00000056_DOBDO<3>_UNCONNECTED , \NLW_blk0000002d/blk00000056_DOBDO<2>_UNCONNECTED ,
\NLW_blk0000002d/blk00000056_DOBDO<1>_UNCONNECTED , \NLW_blk0000002d/blk00000056_DOBDO<0>_UNCONNECTED }),
    .DIPADIP({\blk0000002d/sig00000b54 , \blk0000002d/sig00000b54 })
  );
  RAMB8BWER #(
    .DATA_WIDTH_A ( 36 ),
    .DATA_WIDTH_B ( 36 ),
    .DOA_REG ( 0 ),
    .DOB_REG ( 1 ),
    .EN_RSTRAM_A ( "FALSE" ),
    .EN_RSTRAM_B ( "FALSE" ),
    .INITP_00 ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INITP_01 ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INITP_02 ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INITP_03 ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_00 ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_01 ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_02 ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_03 ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_04 ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_05 ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_06 ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_07 ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_08 ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_09 ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_0A ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_0B ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_0C ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_0D ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_0E ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_0F ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_10 ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_11 ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_12 ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_13 ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_14 ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_15 ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_16 ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_17 ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_18 ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_19 ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_1A ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_1B ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_1C ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_1D ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_1E ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_1F ( 256'h0000000000000000000000000000000000000000000000000000000000000000 ),
    .INIT_A ( 18'h00000 ),
    .INIT_B ( 18'h00000 ),
    .INIT_FILE ( "NONE" ),
    .RAM_MODE ( "SDP" ),
    .RSTTYPE ( "SYNC" ),
    .RST_PRIORITY_A ( "CE" ),
    .RST_PRIORITY_B ( "CE" ),
    .SIM_COLLISION_CHECK ( "GENERATE_X_ONLY" ),
    .SRVAL_A ( 18'h00000 ),
    .SRVAL_B ( 18'h00000 ),
    .WRITE_MODE_A ( "READ_FIRST" ),
    .WRITE_MODE_B ( "READ_FIRST" ))
  \blk0000002d/blk00000055  (
    .RSTBRST(\blk0000002d/sig00000b54 ),
    .ENBRDEN(sig00000001),
    .REGCEA(\blk0000002d/sig00000b54 ),
    .ENAWREN(sig00000001),
    .CLKAWRCLK(clk),
    .CLKBRDCLK(clk),
    .REGCEBREGCE(sig00000001),
    .RSTA(\blk0000002d/sig00000b54 ),
    .WEAWEL({sig0000000a, sig0000000a}),
    .DOADO({\blk0000002d/sig00000b10 , \blk0000002d/sig00000b11 , \blk0000002d/sig00000b12 , \blk0000002d/sig00000b13 , \blk0000002d/sig00000b14 ,
\blk0000002d/sig00000b15 , \blk0000002d/sig00000b16 , \blk0000002d/sig00000b17 , \blk0000002d/sig00000b08 , \blk0000002d/sig00000b09 ,
\blk0000002d/sig00000b0a , \blk0000002d/sig00000b0b , \blk0000002d/sig00000b0c , \blk0000002d/sig00000b0d , \blk0000002d/sig00000b0e ,
\blk0000002d/sig00000b0f }),
    .DOPADOP({\blk0000002d/sig00000b29 , \blk0000002d/sig00000b28 }),
    .DOPBDOP({\blk0000002d/sig00000b2b , \blk0000002d/sig00000b2a }),
    .WEBWEU({sig0000000a, sig0000000a}),
    .ADDRAWRADDR({sig00000040, sig0000003f, sig0000003e, sig0000003d, sig0000003c, sig0000003b, sig0000003a, sig00000039, \blk0000002d/sig00000b54 ,
\blk0000002d/sig00000b54 , \blk0000002d/sig00000b54 , \blk0000002d/sig00000b54 , \blk0000002d/sig00000b54 }),
    .DIPBDIP({sig000000d8, sig000000cf}),
    .DIBDI({sig000000d7, sig000000d6, sig000000d5, sig000000d4, sig000000d3, sig000000d2, sig000000d1, sig000000d0, sig000000ce, sig000000cd,
sig000000cc, sig000000cb, sig000000ca, sig000000c9, sig000000c8, sig000000c7}),
    .DIADI({sig000000c5, sig000000c4, sig000000c3, sig000000c2, sig000000c1, sig000000c0, sig000000bf, sig000000be, sig000000bc, sig000000bb,
sig000000ba, sig000000b9, sig000000b8, sig000000b7, sig000000b6, sig000000b5}),
    .ADDRBRDADDR({sig00000038, sig00000037, sig00000036, sig00000035, sig00000034, sig00000033, sig00000032, sig00000031, \blk0000002d/sig00000b54 ,
\blk0000002d/sig00000b54 , \blk0000002d/sig00000b54 , \blk0000002d/sig00000b54 , \blk0000002d/sig00000b54 }),
    .DOBDO({\blk0000002d/sig00000b20 , \blk0000002d/sig00000b21 , \blk0000002d/sig00000b22 , \blk0000002d/sig00000b23 , \blk0000002d/sig00000b24 ,
\blk0000002d/sig00000b25 , \blk0000002d/sig00000b26 , \blk0000002d/sig00000b27 , \blk0000002d/sig00000b18 , \blk0000002d/sig00000b19 ,
\blk0000002d/sig00000b1a , \blk0000002d/sig00000b1b , \blk0000002d/sig00000b1c , \blk0000002d/sig00000b1d , \blk0000002d/sig00000b1e ,
\blk0000002d/sig00000b1f }),
    .DIPADIP({sig000000c6, sig000000bd})
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk0000002d/blk00000054  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk0000002d/sig00000b2c ),
    .Q(sig00000198)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk0000002d/blk00000053  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk0000002d/sig00000b2d ),
    .Q(sig00000197)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk0000002d/blk00000052  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk0000002d/sig00000b2b ),
    .Q(sig00000196)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk0000002d/blk00000051  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk0000002d/sig00000b20 ),
    .Q(sig00000195)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk0000002d/blk00000050  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk0000002d/sig00000b21 ),
    .Q(sig00000194)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk0000002d/blk0000004f  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk0000002d/sig00000b22 ),
    .Q(sig00000193)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk0000002d/blk0000004e  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk0000002d/sig00000b23 ),
    .Q(sig00000192)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk0000002d/blk0000004d  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk0000002d/sig00000b24 ),
    .Q(sig00000191)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk0000002d/blk0000004c  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk0000002d/sig00000b25 ),
    .Q(sig00000190)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk0000002d/blk0000004b  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk0000002d/sig00000b26 ),
    .Q(sig0000018f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk0000002d/blk0000004a  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk0000002d/sig00000b27 ),
    .Q(sig0000018e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk0000002d/blk00000049  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk0000002d/sig00000b2a ),
    .Q(sig0000018d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk0000002d/blk00000048  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk0000002d/sig00000b18 ),
    .Q(sig0000018c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk0000002d/blk00000047  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk0000002d/sig00000b19 ),
    .Q(sig0000018b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk0000002d/blk00000046  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk0000002d/sig00000b1a ),
    .Q(sig0000018a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk0000002d/blk00000045  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk0000002d/sig00000b1b ),
    .Q(sig00000189)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk0000002d/blk00000044  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk0000002d/sig00000b1c ),
    .Q(sig00000188)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk0000002d/blk00000043  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk0000002d/sig00000b1d ),
    .Q(sig00000187)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk0000002d/blk00000042  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk0000002d/sig00000b1e ),
    .Q(sig00000186)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk0000002d/blk00000041  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk0000002d/sig00000b1f ),
    .Q(sig00000185)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk0000002d/blk00000040  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk0000002d/sig00000b29 ),
    .Q(sig00000184)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk0000002d/blk0000003f  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk0000002d/sig00000b10 ),
    .Q(sig00000183)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk0000002d/blk0000003e  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk0000002d/sig00000b11 ),
    .Q(sig00000182)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk0000002d/blk0000003d  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk0000002d/sig00000b12 ),
    .Q(sig00000181)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk0000002d/blk0000003c  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk0000002d/sig00000b13 ),
    .Q(sig00000180)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk0000002d/blk0000003b  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk0000002d/sig00000b14 ),
    .Q(sig0000017f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk0000002d/blk0000003a  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk0000002d/sig00000b15 ),
    .Q(sig0000017e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk0000002d/blk00000039  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk0000002d/sig00000b16 ),
    .Q(sig0000017d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk0000002d/blk00000038  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk0000002d/sig00000b17 ),
    .Q(sig0000017c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk0000002d/blk00000037  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk0000002d/sig00000b28 ),
    .Q(sig0000017b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk0000002d/blk00000036  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk0000002d/sig00000b08 ),
    .Q(sig0000017a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk0000002d/blk00000035  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk0000002d/sig00000b09 ),
    .Q(sig00000179)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk0000002d/blk00000034  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk0000002d/sig00000b0a ),
    .Q(sig00000178)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk0000002d/blk00000033  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk0000002d/sig00000b0b ),
    .Q(sig00000177)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk0000002d/blk00000032  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk0000002d/sig00000b0c ),
    .Q(sig00000176)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk0000002d/blk00000031  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk0000002d/sig00000b0d ),
    .Q(sig00000175)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk0000002d/blk00000030  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk0000002d/sig00000b0e ),
    .Q(sig00000174)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk0000002d/blk0000002f  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk0000002d/sig00000b0f ),
    .Q(sig00000173)
  );
  GND   \blk0000002d/blk0000002e  (
    .G(\blk0000002d/sig00000b54 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk0000018c/blk00000193  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk0000018c/sig00000bcc ),
    .Q(sig0000055c)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk0000018c/blk00000192  (
    .A0(\blk0000018c/sig00000bc9 ),
    .A1(\blk0000018c/sig00000bc9 ),
    .A2(\blk0000018c/sig00000bc9 ),
    .A3(\blk0000018c/sig00000bc9 ),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000004de),
    .Q(\blk0000018c/sig00000bcc ),
    .Q15(\NLW_blk0000018c/blk00000192_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk0000018c/blk00000191  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk0000018c/sig00000bcb ),
    .Q(sig0000055b)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk0000018c/blk00000190  (
    .A0(\blk0000018c/sig00000bc9 ),
    .A1(\blk0000018c/sig00000bc9 ),
    .A2(\blk0000018c/sig00000bc9 ),
    .A3(\blk0000018c/sig00000bc9 ),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000004dd),
    .Q(\blk0000018c/sig00000bcb ),
    .Q15(\NLW_blk0000018c/blk00000190_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk0000018c/blk0000018f  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk0000018c/sig00000bca ),
    .Q(sig0000055d)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk0000018c/blk0000018e  (
    .A0(\blk0000018c/sig00000bc9 ),
    .A1(\blk0000018c/sig00000bc9 ),
    .A2(\blk0000018c/sig00000bc9 ),
    .A3(\blk0000018c/sig00000bc9 ),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000004df),
    .Q(\blk0000018c/sig00000bca ),
    .Q15(\NLW_blk0000018c/blk0000018e_Q15_UNCONNECTED )
  );
  GND   \blk0000018c/blk0000018d  (
    .G(\blk0000018c/sig00000bc9 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000194/blk0000019b  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk00000194/sig00000bd8 ),
    .Q(sig0000031e)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000194/blk0000019a  (
    .A0(\blk00000194/sig00000bd5 ),
    .A1(\blk00000194/sig00000bd5 ),
    .A2(\blk00000194/sig00000bd5 ),
    .A3(\blk00000194/sig00000bd5 ),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000004a2),
    .Q(\blk00000194/sig00000bd8 ),
    .Q15(\NLW_blk00000194/blk0000019a_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000194/blk00000199  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk00000194/sig00000bd7 ),
    .Q(sig0000031f)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000194/blk00000198  (
    .A0(\blk00000194/sig00000bd5 ),
    .A1(\blk00000194/sig00000bd5 ),
    .A2(\blk00000194/sig00000bd5 ),
    .A3(\blk00000194/sig00000bd5 ),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000004a1),
    .Q(\blk00000194/sig00000bd7 ),
    .Q15(\NLW_blk00000194/blk00000198_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000194/blk00000197  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk00000194/sig00000bd6 ),
    .Q(sig0000031d)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000194/blk00000196  (
    .A0(\blk00000194/sig00000bd5 ),
    .A1(\blk00000194/sig00000bd5 ),
    .A2(\blk00000194/sig00000bd5 ),
    .A3(\blk00000194/sig00000bd5 ),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000004a3),
    .Q(\blk00000194/sig00000bd6 ),
    .Q15(\NLW_blk00000194/blk00000196_Q15_UNCONNECTED )
  );
  GND   \blk00000194/blk00000195  (
    .G(\blk00000194/sig00000bd5 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk0000019d/blk000001b6  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk0000019d/sig00000c00 ),
    .Q(sig00000240)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk0000019d/blk000001b5  (
    .A0(\blk0000019d/sig00000bf4 ),
    .A1(\blk0000019d/sig00000bf4 ),
    .A2(\blk0000019d/sig00000bf4 ),
    .A3(\blk0000019d/sig00000bf4 ),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000005ce),
    .Q(\blk0000019d/sig00000c00 ),
    .Q15(\NLW_blk0000019d/blk000001b5_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk0000019d/blk000001b4  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk0000019d/sig00000bff ),
    .Q(sig0000023f)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk0000019d/blk000001b3  (
    .A0(\blk0000019d/sig00000bf4 ),
    .A1(\blk0000019d/sig00000bf4 ),
    .A2(\blk0000019d/sig00000bf4 ),
    .A3(\blk0000019d/sig00000bf4 ),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000005cd),
    .Q(\blk0000019d/sig00000bff ),
    .Q15(\NLW_blk0000019d/blk000001b3_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk0000019d/blk000001b2  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk0000019d/sig00000bfe ),
    .Q(sig00000241)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk0000019d/blk000001b1  (
    .A0(\blk0000019d/sig00000bf4 ),
    .A1(\blk0000019d/sig00000bf4 ),
    .A2(\blk0000019d/sig00000bf4 ),
    .A3(\blk0000019d/sig00000bf4 ),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000005cf),
    .Q(\blk0000019d/sig00000bfe ),
    .Q15(\NLW_blk0000019d/blk000001b1_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk0000019d/blk000001b0  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk0000019d/sig00000bfd ),
    .Q(sig0000023d)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk0000019d/blk000001af  (
    .A0(\blk0000019d/sig00000bf4 ),
    .A1(\blk0000019d/sig00000bf4 ),
    .A2(\blk0000019d/sig00000bf4 ),
    .A3(\blk0000019d/sig00000bf4 ),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000005cb),
    .Q(\blk0000019d/sig00000bfd ),
    .Q15(\NLW_blk0000019d/blk000001af_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk0000019d/blk000001ae  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk0000019d/sig00000bfc ),
    .Q(sig0000023c)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk0000019d/blk000001ad  (
    .A0(\blk0000019d/sig00000bf4 ),
    .A1(\blk0000019d/sig00000bf4 ),
    .A2(\blk0000019d/sig00000bf4 ),
    .A3(\blk0000019d/sig00000bf4 ),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000005ca),
    .Q(\blk0000019d/sig00000bfc ),
    .Q15(\NLW_blk0000019d/blk000001ad_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk0000019d/blk000001ac  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk0000019d/sig00000bfb ),
    .Q(sig0000023e)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk0000019d/blk000001ab  (
    .A0(\blk0000019d/sig00000bf4 ),
    .A1(\blk0000019d/sig00000bf4 ),
    .A2(\blk0000019d/sig00000bf4 ),
    .A3(\blk0000019d/sig00000bf4 ),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000005cc),
    .Q(\blk0000019d/sig00000bfb ),
    .Q15(\NLW_blk0000019d/blk000001ab_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk0000019d/blk000001aa  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk0000019d/sig00000bfa ),
    .Q(sig0000023a)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk0000019d/blk000001a9  (
    .A0(\blk0000019d/sig00000bf4 ),
    .A1(\blk0000019d/sig00000bf4 ),
    .A2(\blk0000019d/sig00000bf4 ),
    .A3(\blk0000019d/sig00000bf4 ),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000005c8),
    .Q(\blk0000019d/sig00000bfa ),
    .Q15(\NLW_blk0000019d/blk000001a9_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk0000019d/blk000001a8  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk0000019d/sig00000bf9 ),
    .Q(sig00000239)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk0000019d/blk000001a7  (
    .A0(\blk0000019d/sig00000bf4 ),
    .A1(\blk0000019d/sig00000bf4 ),
    .A2(\blk0000019d/sig00000bf4 ),
    .A3(\blk0000019d/sig00000bf4 ),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000005c7),
    .Q(\blk0000019d/sig00000bf9 ),
    .Q15(\NLW_blk0000019d/blk000001a7_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk0000019d/blk000001a6  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk0000019d/sig00000bf8 ),
    .Q(sig0000023b)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk0000019d/blk000001a5  (
    .A0(\blk0000019d/sig00000bf4 ),
    .A1(\blk0000019d/sig00000bf4 ),
    .A2(\blk0000019d/sig00000bf4 ),
    .A3(\blk0000019d/sig00000bf4 ),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000005c9),
    .Q(\blk0000019d/sig00000bf8 ),
    .Q15(\NLW_blk0000019d/blk000001a5_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk0000019d/blk000001a4  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk0000019d/sig00000bf7 ),
    .Q(sig00000237)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk0000019d/blk000001a3  (
    .A0(\blk0000019d/sig00000bf4 ),
    .A1(\blk0000019d/sig00000bf4 ),
    .A2(\blk0000019d/sig00000bf4 ),
    .A3(\blk0000019d/sig00000bf4 ),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000005c5),
    .Q(\blk0000019d/sig00000bf7 ),
    .Q15(\NLW_blk0000019d/blk000001a3_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk0000019d/blk000001a2  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk0000019d/sig00000bf6 ),
    .Q(sig00000236)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk0000019d/blk000001a1  (
    .A0(\blk0000019d/sig00000bf4 ),
    .A1(\blk0000019d/sig00000bf4 ),
    .A2(\blk0000019d/sig00000bf4 ),
    .A3(\blk0000019d/sig00000bf4 ),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000005c4),
    .Q(\blk0000019d/sig00000bf6 ),
    .Q15(\NLW_blk0000019d/blk000001a1_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk0000019d/blk000001a0  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk0000019d/sig00000bf5 ),
    .Q(sig00000238)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk0000019d/blk0000019f  (
    .A0(\blk0000019d/sig00000bf4 ),
    .A1(\blk0000019d/sig00000bf4 ),
    .A2(\blk0000019d/sig00000bf4 ),
    .A3(\blk0000019d/sig00000bf4 ),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000005c6),
    .Q(\blk0000019d/sig00000bf5 ),
    .Q15(\NLW_blk0000019d/blk0000019f_Q15_UNCONNECTED )
  );
  GND   \blk0000019d/blk0000019e  (
    .G(\blk0000019d/sig00000bf4 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000001b7/blk000001d0  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk000001b7/sig00000c27 ),
    .Q(sig00000229)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk000001b7/blk000001cf  (
    .A0(\blk000001b7/sig00000c1b ),
    .A1(\blk000001b7/sig00000c1b ),
    .A2(\blk000001b7/sig00000c1b ),
    .A3(\blk000001b7/sig00000c1b ),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000002ac),
    .Q(\blk000001b7/sig00000c27 ),
    .Q15(\NLW_blk000001b7/blk000001cf_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000001b7/blk000001ce  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk000001b7/sig00000c26 ),
    .Q(sig00000228)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk000001b7/blk000001cd  (
    .A0(\blk000001b7/sig00000c1b ),
    .A1(\blk000001b7/sig00000c1b ),
    .A2(\blk000001b7/sig00000c1b ),
    .A3(\blk000001b7/sig00000c1b ),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000002ad),
    .Q(\blk000001b7/sig00000c26 ),
    .Q15(\NLW_blk000001b7/blk000001cd_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000001b7/blk000001cc  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk000001b7/sig00000c25 ),
    .Q(sig0000022a)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk000001b7/blk000001cb  (
    .A0(\blk000001b7/sig00000c1b ),
    .A1(\blk000001b7/sig00000c1b ),
    .A2(\blk000001b7/sig00000c1b ),
    .A3(\blk000001b7/sig00000c1b ),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000002ab),
    .Q(\blk000001b7/sig00000c25 ),
    .Q15(\NLW_blk000001b7/blk000001cb_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000001b7/blk000001ca  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk000001b7/sig00000c24 ),
    .Q(sig00000226)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk000001b7/blk000001c9  (
    .A0(\blk000001b7/sig00000c1b ),
    .A1(\blk000001b7/sig00000c1b ),
    .A2(\blk000001b7/sig00000c1b ),
    .A3(\blk000001b7/sig00000c1b ),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000002af),
    .Q(\blk000001b7/sig00000c24 ),
    .Q15(\NLW_blk000001b7/blk000001c9_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000001b7/blk000001c8  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk000001b7/sig00000c23 ),
    .Q(sig00000225)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk000001b7/blk000001c7  (
    .A0(\blk000001b7/sig00000c1b ),
    .A1(\blk000001b7/sig00000c1b ),
    .A2(\blk000001b7/sig00000c1b ),
    .A3(\blk000001b7/sig00000c1b ),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000002b0),
    .Q(\blk000001b7/sig00000c23 ),
    .Q15(\NLW_blk000001b7/blk000001c7_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000001b7/blk000001c6  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk000001b7/sig00000c22 ),
    .Q(sig00000227)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk000001b7/blk000001c5  (
    .A0(\blk000001b7/sig00000c1b ),
    .A1(\blk000001b7/sig00000c1b ),
    .A2(\blk000001b7/sig00000c1b ),
    .A3(\blk000001b7/sig00000c1b ),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000002ae),
    .Q(\blk000001b7/sig00000c22 ),
    .Q15(\NLW_blk000001b7/blk000001c5_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000001b7/blk000001c4  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk000001b7/sig00000c21 ),
    .Q(sig00000223)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk000001b7/blk000001c3  (
    .A0(\blk000001b7/sig00000c1b ),
    .A1(\blk000001b7/sig00000c1b ),
    .A2(\blk000001b7/sig00000c1b ),
    .A3(\blk000001b7/sig00000c1b ),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000002b2),
    .Q(\blk000001b7/sig00000c21 ),
    .Q15(\NLW_blk000001b7/blk000001c3_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000001b7/blk000001c2  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk000001b7/sig00000c20 ),
    .Q(sig00000222)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk000001b7/blk000001c1  (
    .A0(\blk000001b7/sig00000c1b ),
    .A1(\blk000001b7/sig00000c1b ),
    .A2(\blk000001b7/sig00000c1b ),
    .A3(\blk000001b7/sig00000c1b ),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000002b3),
    .Q(\blk000001b7/sig00000c20 ),
    .Q15(\NLW_blk000001b7/blk000001c1_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000001b7/blk000001c0  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk000001b7/sig00000c1f ),
    .Q(sig00000224)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk000001b7/blk000001bf  (
    .A0(\blk000001b7/sig00000c1b ),
    .A1(\blk000001b7/sig00000c1b ),
    .A2(\blk000001b7/sig00000c1b ),
    .A3(\blk000001b7/sig00000c1b ),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000002b1),
    .Q(\blk000001b7/sig00000c1f ),
    .Q15(\NLW_blk000001b7/blk000001bf_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000001b7/blk000001be  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk000001b7/sig00000c1e ),
    .Q(sig00000220)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk000001b7/blk000001bd  (
    .A0(\blk000001b7/sig00000c1b ),
    .A1(\blk000001b7/sig00000c1b ),
    .A2(\blk000001b7/sig00000c1b ),
    .A3(\blk000001b7/sig00000c1b ),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000002b5),
    .Q(\blk000001b7/sig00000c1e ),
    .Q15(\NLW_blk000001b7/blk000001bd_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000001b7/blk000001bc  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk000001b7/sig00000c1d ),
    .Q(sig0000021f)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk000001b7/blk000001bb  (
    .A0(\blk000001b7/sig00000c1b ),
    .A1(\blk000001b7/sig00000c1b ),
    .A2(\blk000001b7/sig00000c1b ),
    .A3(\blk000001b7/sig00000c1b ),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000002b6),
    .Q(\blk000001b7/sig00000c1d ),
    .Q15(\NLW_blk000001b7/blk000001bb_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000001b7/blk000001ba  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk000001b7/sig00000c1c ),
    .Q(sig00000221)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk000001b7/blk000001b9  (
    .A0(\blk000001b7/sig00000c1b ),
    .A1(\blk000001b7/sig00000c1b ),
    .A2(\blk000001b7/sig00000c1b ),
    .A3(\blk000001b7/sig00000c1b ),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000002b4),
    .Q(\blk000001b7/sig00000c1c ),
    .Q15(\NLW_blk000001b7/blk000001b9_Q15_UNCONNECTED )
  );
  GND   \blk000001b7/blk000001b8  (
    .G(\blk000001b7/sig00000c1b )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000001d1/blk000001f4  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk000001d1/sig00000c5d ),
    .Q(sig000004b4)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk000001d1/blk000001f3  (
    .A0(\blk000001d1/sig00000c4c ),
    .A1(\blk000001d1/sig00000c4c ),
    .A2(\blk000001d1/sig00000c4c ),
    .A3(\blk000001d1/sig00000c4c ),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig00000368),
    .Q(\blk000001d1/sig00000c5d ),
    .Q15(\NLW_blk000001d1/blk000001f3_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000001d1/blk000001f2  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk000001d1/sig00000c5c ),
    .Q(sig000004b3)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk000001d1/blk000001f1  (
    .A0(\blk000001d1/sig00000c4c ),
    .A1(\blk000001d1/sig00000c4c ),
    .A2(\blk000001d1/sig00000c4c ),
    .A3(\blk000001d1/sig00000c4c ),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig00000369),
    .Q(\blk000001d1/sig00000c5c ),
    .Q15(\NLW_blk000001d1/blk000001f1_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000001d1/blk000001f0  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk000001d1/sig00000c5b ),
    .Q(sig000004b2)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk000001d1/blk000001ef  (
    .A0(\blk000001d1/sig00000c4c ),
    .A1(\blk000001d1/sig00000c4c ),
    .A2(\blk000001d1/sig00000c4c ),
    .A3(\blk000001d1/sig00000c4c ),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig0000036a),
    .Q(\blk000001d1/sig00000c5b ),
    .Q15(\NLW_blk000001d1/blk000001ef_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000001d1/blk000001ee  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk000001d1/sig00000c5a ),
    .Q(sig000004b1)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk000001d1/blk000001ed  (
    .A0(\blk000001d1/sig00000c4c ),
    .A1(\blk000001d1/sig00000c4c ),
    .A2(\blk000001d1/sig00000c4c ),
    .A3(\blk000001d1/sig00000c4c ),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig0000036b),
    .Q(\blk000001d1/sig00000c5a ),
    .Q15(\NLW_blk000001d1/blk000001ed_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000001d1/blk000001ec  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk000001d1/sig00000c59 ),
    .Q(sig000004b0)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk000001d1/blk000001eb  (
    .A0(\blk000001d1/sig00000c4c ),
    .A1(\blk000001d1/sig00000c4c ),
    .A2(\blk000001d1/sig00000c4c ),
    .A3(\blk000001d1/sig00000c4c ),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig0000036c),
    .Q(\blk000001d1/sig00000c59 ),
    .Q15(\NLW_blk000001d1/blk000001eb_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000001d1/blk000001ea  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk000001d1/sig00000c58 ),
    .Q(sig000004af)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk000001d1/blk000001e9  (
    .A0(\blk000001d1/sig00000c4c ),
    .A1(\blk000001d1/sig00000c4c ),
    .A2(\blk000001d1/sig00000c4c ),
    .A3(\blk000001d1/sig00000c4c ),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig0000036d),
    .Q(\blk000001d1/sig00000c58 ),
    .Q15(\NLW_blk000001d1/blk000001e9_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000001d1/blk000001e8  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk000001d1/sig00000c57 ),
    .Q(sig000004ae)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk000001d1/blk000001e7  (
    .A0(\blk000001d1/sig00000c4c ),
    .A1(\blk000001d1/sig00000c4c ),
    .A2(\blk000001d1/sig00000c4c ),
    .A3(\blk000001d1/sig00000c4c ),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig0000036e),
    .Q(\blk000001d1/sig00000c57 ),
    .Q15(\NLW_blk000001d1/blk000001e7_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000001d1/blk000001e6  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk000001d1/sig00000c56 ),
    .Q(sig000004ad)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk000001d1/blk000001e5  (
    .A0(\blk000001d1/sig00000c4c ),
    .A1(\blk000001d1/sig00000c4c ),
    .A2(\blk000001d1/sig00000c4c ),
    .A3(\blk000001d1/sig00000c4c ),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig0000036f),
    .Q(\blk000001d1/sig00000c56 ),
    .Q15(\NLW_blk000001d1/blk000001e5_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000001d1/blk000001e4  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk000001d1/sig00000c55 ),
    .Q(sig000004ac)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk000001d1/blk000001e3  (
    .A0(\blk000001d1/sig00000c4c ),
    .A1(\blk000001d1/sig00000c4c ),
    .A2(\blk000001d1/sig00000c4c ),
    .A3(\blk000001d1/sig00000c4c ),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig00000370),
    .Q(\blk000001d1/sig00000c55 ),
    .Q15(\NLW_blk000001d1/blk000001e3_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000001d1/blk000001e2  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk000001d1/sig00000c54 ),
    .Q(sig000004ab)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk000001d1/blk000001e1  (
    .A0(\blk000001d1/sig00000c4c ),
    .A1(\blk000001d1/sig00000c4c ),
    .A2(\blk000001d1/sig00000c4c ),
    .A3(\blk000001d1/sig00000c4c ),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig00000371),
    .Q(\blk000001d1/sig00000c54 ),
    .Q15(\NLW_blk000001d1/blk000001e1_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000001d1/blk000001e0  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk000001d1/sig00000c53 ),
    .Q(sig000004aa)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk000001d1/blk000001df  (
    .A0(\blk000001d1/sig00000c4c ),
    .A1(\blk000001d1/sig00000c4c ),
    .A2(\blk000001d1/sig00000c4c ),
    .A3(\blk000001d1/sig00000c4c ),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig00000372),
    .Q(\blk000001d1/sig00000c53 ),
    .Q15(\NLW_blk000001d1/blk000001df_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000001d1/blk000001de  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk000001d1/sig00000c52 ),
    .Q(sig000004a9)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk000001d1/blk000001dd  (
    .A0(\blk000001d1/sig00000c4c ),
    .A1(\blk000001d1/sig00000c4c ),
    .A2(\blk000001d1/sig00000c4c ),
    .A3(\blk000001d1/sig00000c4c ),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig00000373),
    .Q(\blk000001d1/sig00000c52 ),
    .Q15(\NLW_blk000001d1/blk000001dd_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000001d1/blk000001dc  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk000001d1/sig00000c51 ),
    .Q(sig000004a8)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk000001d1/blk000001db  (
    .A0(\blk000001d1/sig00000c4c ),
    .A1(\blk000001d1/sig00000c4c ),
    .A2(\blk000001d1/sig00000c4c ),
    .A3(\blk000001d1/sig00000c4c ),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig00000374),
    .Q(\blk000001d1/sig00000c51 ),
    .Q15(\NLW_blk000001d1/blk000001db_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000001d1/blk000001da  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk000001d1/sig00000c50 ),
    .Q(sig000004a7)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk000001d1/blk000001d9  (
    .A0(\blk000001d1/sig00000c4c ),
    .A1(\blk000001d1/sig00000c4c ),
    .A2(\blk000001d1/sig00000c4c ),
    .A3(\blk000001d1/sig00000c4c ),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig00000375),
    .Q(\blk000001d1/sig00000c50 ),
    .Q15(\NLW_blk000001d1/blk000001d9_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000001d1/blk000001d8  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk000001d1/sig00000c4f ),
    .Q(sig000004a5)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk000001d1/blk000001d7  (
    .A0(\blk000001d1/sig00000c4c ),
    .A1(\blk000001d1/sig00000c4c ),
    .A2(\blk000001d1/sig00000c4c ),
    .A3(\blk000001d1/sig00000c4c ),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig00000377),
    .Q(\blk000001d1/sig00000c4f ),
    .Q15(\NLW_blk000001d1/blk000001d7_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000001d1/blk000001d6  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk000001d1/sig00000c4e ),
    .Q(sig000004a4)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk000001d1/blk000001d5  (
    .A0(\blk000001d1/sig00000c4c ),
    .A1(\blk000001d1/sig00000c4c ),
    .A2(\blk000001d1/sig00000c4c ),
    .A3(\blk000001d1/sig00000c4c ),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig00000378),
    .Q(\blk000001d1/sig00000c4e ),
    .Q15(\NLW_blk000001d1/blk000001d5_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000001d1/blk000001d4  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk000001d1/sig00000c4d ),
    .Q(sig000004a6)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk000001d1/blk000001d3  (
    .A0(\blk000001d1/sig00000c4c ),
    .A1(\blk000001d1/sig00000c4c ),
    .A2(\blk000001d1/sig00000c4c ),
    .A3(\blk000001d1/sig00000c4c ),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig00000376),
    .Q(\blk000001d1/sig00000c4d ),
    .Q15(\NLW_blk000001d1/blk000001d3_Q15_UNCONNECTED )
  );
  GND   \blk000001d1/blk000001d2  (
    .G(\blk000001d1/sig00000c4c )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000001f8/blk000001fd  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk000001f8/sig00000cd2 ),
    .Q(sig000003da)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk000001f8/blk000001fc  (
    .A0(\blk000001f8/sig00000cd0 ),
    .A1(\blk000001f8/sig00000cd0 ),
    .A2(\blk000001f8/sig00000cd0 ),
    .A3(\blk000001f8/sig00000cd0 ),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig00000519),
    .Q(\blk000001f8/sig00000cd2 ),
    .Q15(\NLW_blk000001f8/blk000001fc_Q15_UNCONNECTED )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000001f8/blk000001fb  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk000001f8/sig00000cd1 ),
    .Q(sig000003db)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk000001f8/blk000001fa  (
    .A0(\blk000001f8/sig00000cd0 ),
    .A1(\blk000001f8/sig00000cd0 ),
    .A2(\blk000001f8/sig00000cd0 ),
    .A3(\blk000001f8/sig00000cd0 ),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig00000518),
    .Q(\blk000001f8/sig00000cd1 ),
    .Q15(\NLW_blk000001f8/blk000001fa_Q15_UNCONNECTED )
  );
  GND   \blk000001f8/blk000001f9  (
    .G(\blk000001f8/sig00000cd0 )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk000001fe/blk0000025c  (
    .I0(sig00000199),
    .O(\blk000001fe/sig00000d5e )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk000001fe/blk0000025b  (
    .I0(sig0000019a),
    .O(\blk000001fe/sig00000d5d )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk000001fe/blk0000025a  (
    .I0(sig0000019b),
    .O(\blk000001fe/sig00000d5c )
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  \blk000001fe/blk00000259  (
    .I0(sig0000025f),
    .I1(sig000001af),
    .O(\blk000001fe/sig00000d5b )
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  \blk000001fe/blk00000258  (
    .I0(sig0000025f),
    .I1(sig000001af),
    .O(\blk000001fe/sig00000d30 )
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  \blk000001fe/blk00000257  (
    .I0(sig0000025f),
    .I1(sig000001ae),
    .O(\blk000001fe/sig00000d31 )
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  \blk000001fe/blk00000256  (
    .I0(sig0000025e),
    .I1(sig000001ad),
    .O(\blk000001fe/sig00000d32 )
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  \blk000001fe/blk00000255  (
    .I0(sig0000025d),
    .I1(sig000001ac),
    .O(\blk000001fe/sig00000d33 )
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  \blk000001fe/blk00000254  (
    .I0(sig0000025c),
    .I1(sig000001ab),
    .O(\blk000001fe/sig00000d34 )
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  \blk000001fe/blk00000253  (
    .I0(sig0000025b),
    .I1(sig000001aa),
    .O(\blk000001fe/sig00000d35 )
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  \blk000001fe/blk00000252  (
    .I0(sig0000025a),
    .I1(sig000001a9),
    .O(\blk000001fe/sig00000d36 )
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  \blk000001fe/blk00000251  (
    .I0(sig00000259),
    .I1(sig000001a8),
    .O(\blk000001fe/sig00000d37 )
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  \blk000001fe/blk00000250  (
    .I0(sig00000258),
    .I1(sig000001a7),
    .O(\blk000001fe/sig00000d38 )
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  \blk000001fe/blk0000024f  (
    .I0(sig00000257),
    .I1(sig000001a6),
    .O(\blk000001fe/sig00000d39 )
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  \blk000001fe/blk0000024e  (
    .I0(sig00000256),
    .I1(sig000001a5),
    .O(\blk000001fe/sig00000d3a )
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  \blk000001fe/blk0000024d  (
    .I0(sig00000255),
    .I1(sig000001a4),
    .O(\blk000001fe/sig00000d3b )
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  \blk000001fe/blk0000024c  (
    .I0(sig00000254),
    .I1(sig000001a3),
    .O(\blk000001fe/sig00000d3c )
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  \blk000001fe/blk0000024b  (
    .I0(sig00000253),
    .I1(sig000001a2),
    .O(\blk000001fe/sig00000d3d )
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  \blk000001fe/blk0000024a  (
    .I0(sig00000252),
    .I1(sig000001a1),
    .O(\blk000001fe/sig00000d3e )
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  \blk000001fe/blk00000249  (
    .I0(sig00000251),
    .I1(sig000001a0),
    .O(\blk000001fe/sig00000d3f )
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  \blk000001fe/blk00000248  (
    .I0(sig00000250),
    .I1(sig0000019f),
    .O(\blk000001fe/sig00000d40 )
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  \blk000001fe/blk00000247  (
    .I0(sig0000024f),
    .I1(sig0000019e),
    .O(\blk000001fe/sig00000d41 )
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  \blk000001fe/blk00000246  (
    .I0(sig0000024e),
    .I1(sig0000019d),
    .O(\blk000001fe/sig00000d42 )
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  \blk000001fe/blk00000245  (
    .I0(sig0000024d),
    .I1(sig0000019c),
    .O(\blk000001fe/sig00000d43 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000001fe/blk00000244  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk000001fe/sig00000d1a ),
    .Q(sig00000209)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000001fe/blk00000243  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk000001fe/sig00000d2f ),
    .Q(sig0000020a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000001fe/blk00000242  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk000001fe/sig00000d2e ),
    .Q(sig0000020b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000001fe/blk00000241  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk000001fe/sig00000d2d ),
    .Q(sig0000020c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000001fe/blk00000240  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk000001fe/sig00000d2c ),
    .Q(sig0000020d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000001fe/blk0000023f  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk000001fe/sig00000d2b ),
    .Q(sig0000020e)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000001fe/blk0000023e  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk000001fe/sig00000d2a ),
    .Q(sig0000020f)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000001fe/blk0000023d  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk000001fe/sig00000d29 ),
    .Q(sig00000210)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000001fe/blk0000023c  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk000001fe/sig00000d28 ),
    .Q(sig00000211)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000001fe/blk0000023b  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk000001fe/sig00000d27 ),
    .Q(sig00000212)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000001fe/blk0000023a  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk000001fe/sig00000d26 ),
    .Q(sig00000213)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000001fe/blk00000239  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk000001fe/sig00000d25 ),
    .Q(sig00000214)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000001fe/blk00000238  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk000001fe/sig00000d24 ),
    .Q(sig00000215)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000001fe/blk00000237  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk000001fe/sig00000d23 ),
    .Q(sig00000216)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000001fe/blk00000236  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk000001fe/sig00000d22 ),
    .Q(sig00000217)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000001fe/blk00000235  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk000001fe/sig00000d21 ),
    .Q(sig00000218)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000001fe/blk00000234  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk000001fe/sig00000d20 ),
    .Q(sig00000219)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000001fe/blk00000233  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk000001fe/sig00000d1f ),
    .Q(sig0000021a)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000001fe/blk00000232  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk000001fe/sig00000d1e ),
    .Q(sig0000021b)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000001fe/blk00000231  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk000001fe/sig00000d1d ),
    .Q(sig0000021c)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000001fe/blk00000230  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk000001fe/sig00000d1c ),
    .Q(sig0000021d)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000001fe/blk0000022f  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk000001fe/sig00000d1b ),
    .Q(sig0000021e)
  );
  MUXCY   \blk000001fe/blk0000022e  (
    .CI(\blk000001fe/sig00000d19 ),
    .DI(sig00000002),
    .S(\blk000001fe/sig00000d5e ),
    .O(\blk000001fe/sig00000d5a )
  );
  MUXCY   \blk000001fe/blk0000022d  (
    .CI(\blk000001fe/sig00000d5a ),
    .DI(sig00000002),
    .S(\blk000001fe/sig00000d5d ),
    .O(\blk000001fe/sig00000d59 )
  );
  MUXCY   \blk000001fe/blk0000022c  (
    .CI(\blk000001fe/sig00000d59 ),
    .DI(sig00000002),
    .S(\blk000001fe/sig00000d5c ),
    .O(\blk000001fe/sig00000d58 )
  );
  MUXCY   \blk000001fe/blk0000022b  (
    .CI(\blk000001fe/sig00000d58 ),
    .DI(sig0000024d),
    .S(\blk000001fe/sig00000d43 ),
    .O(\blk000001fe/sig00000d57 )
  );
  MUXCY   \blk000001fe/blk0000022a  (
    .CI(\blk000001fe/sig00000d57 ),
    .DI(sig0000024e),
    .S(\blk000001fe/sig00000d42 ),
    .O(\blk000001fe/sig00000d56 )
  );
  MUXCY   \blk000001fe/blk00000229  (
    .CI(\blk000001fe/sig00000d56 ),
    .DI(sig0000024f),
    .S(\blk000001fe/sig00000d41 ),
    .O(\blk000001fe/sig00000d55 )
  );
  MUXCY   \blk000001fe/blk00000228  (
    .CI(\blk000001fe/sig00000d55 ),
    .DI(sig00000250),
    .S(\blk000001fe/sig00000d40 ),
    .O(\blk000001fe/sig00000d54 )
  );
  MUXCY   \blk000001fe/blk00000227  (
    .CI(\blk000001fe/sig00000d54 ),
    .DI(sig00000251),
    .S(\blk000001fe/sig00000d3f ),
    .O(\blk000001fe/sig00000d53 )
  );
  MUXCY   \blk000001fe/blk00000226  (
    .CI(\blk000001fe/sig00000d53 ),
    .DI(sig00000252),
    .S(\blk000001fe/sig00000d3e ),
    .O(\blk000001fe/sig00000d52 )
  );
  MUXCY   \blk000001fe/blk00000225  (
    .CI(\blk000001fe/sig00000d52 ),
    .DI(sig00000253),
    .S(\blk000001fe/sig00000d3d ),
    .O(\blk000001fe/sig00000d51 )
  );
  MUXCY   \blk000001fe/blk00000224  (
    .CI(\blk000001fe/sig00000d51 ),
    .DI(sig00000254),
    .S(\blk000001fe/sig00000d3c ),
    .O(\blk000001fe/sig00000d50 )
  );
  MUXCY   \blk000001fe/blk00000223  (
    .CI(\blk000001fe/sig00000d50 ),
    .DI(sig00000255),
    .S(\blk000001fe/sig00000d3b ),
    .O(\blk000001fe/sig00000d4f )
  );
  MUXCY   \blk000001fe/blk00000222  (
    .CI(\blk000001fe/sig00000d4f ),
    .DI(sig00000256),
    .S(\blk000001fe/sig00000d3a ),
    .O(\blk000001fe/sig00000d4e )
  );
  MUXCY   \blk000001fe/blk00000221  (
    .CI(\blk000001fe/sig00000d4e ),
    .DI(sig00000257),
    .S(\blk000001fe/sig00000d39 ),
    .O(\blk000001fe/sig00000d4d )
  );
  MUXCY   \blk000001fe/blk00000220  (
    .CI(\blk000001fe/sig00000d4d ),
    .DI(sig00000258),
    .S(\blk000001fe/sig00000d38 ),
    .O(\blk000001fe/sig00000d4c )
  );
  MUXCY   \blk000001fe/blk0000021f  (
    .CI(\blk000001fe/sig00000d4c ),
    .DI(sig00000259),
    .S(\blk000001fe/sig00000d37 ),
    .O(\blk000001fe/sig00000d4b )
  );
  MUXCY   \blk000001fe/blk0000021e  (
    .CI(\blk000001fe/sig00000d4b ),
    .DI(sig0000025a),
    .S(\blk000001fe/sig00000d36 ),
    .O(\blk000001fe/sig00000d4a )
  );
  MUXCY   \blk000001fe/blk0000021d  (
    .CI(\blk000001fe/sig00000d4a ),
    .DI(sig0000025b),
    .S(\blk000001fe/sig00000d35 ),
    .O(\blk000001fe/sig00000d49 )
  );
  MUXCY   \blk000001fe/blk0000021c  (
    .CI(\blk000001fe/sig00000d49 ),
    .DI(sig0000025c),
    .S(\blk000001fe/sig00000d34 ),
    .O(\blk000001fe/sig00000d48 )
  );
  MUXCY   \blk000001fe/blk0000021b  (
    .CI(\blk000001fe/sig00000d48 ),
    .DI(sig0000025d),
    .S(\blk000001fe/sig00000d33 ),
    .O(\blk000001fe/sig00000d47 )
  );
  MUXCY   \blk000001fe/blk0000021a  (
    .CI(\blk000001fe/sig00000d47 ),
    .DI(sig0000025e),
    .S(\blk000001fe/sig00000d32 ),
    .O(\blk000001fe/sig00000d46 )
  );
  MUXCY   \blk000001fe/blk00000219  (
    .CI(\blk000001fe/sig00000d46 ),
    .DI(sig0000025f),
    .S(\blk000001fe/sig00000d31 ),
    .O(\blk000001fe/sig00000d45 )
  );
  MUXCY   \blk000001fe/blk00000218  (
    .CI(\blk000001fe/sig00000d45 ),
    .DI(sig0000025f),
    .S(\blk000001fe/sig00000d5b ),
    .O(\blk000001fe/sig00000d44 )
  );
  XORCY   \blk000001fe/blk00000217  (
    .CI(\blk000001fe/sig00000d5a ),
    .LI(\blk000001fe/sig00000d5d ),
    .O(\blk000001fe/sig00000d2f )
  );
  XORCY   \blk000001fe/blk00000216  (
    .CI(\blk000001fe/sig00000d59 ),
    .LI(\blk000001fe/sig00000d5c ),
    .O(\blk000001fe/sig00000d2e )
  );
  XORCY   \blk000001fe/blk00000215  (
    .CI(\blk000001fe/sig00000d58 ),
    .LI(\blk000001fe/sig00000d43 ),
    .O(\blk000001fe/sig00000d2d )
  );
  XORCY   \blk000001fe/blk00000214  (
    .CI(\blk000001fe/sig00000d57 ),
    .LI(\blk000001fe/sig00000d42 ),
    .O(\blk000001fe/sig00000d2c )
  );
  XORCY   \blk000001fe/blk00000213  (
    .CI(\blk000001fe/sig00000d56 ),
    .LI(\blk000001fe/sig00000d41 ),
    .O(\blk000001fe/sig00000d2b )
  );
  XORCY   \blk000001fe/blk00000212  (
    .CI(\blk000001fe/sig00000d55 ),
    .LI(\blk000001fe/sig00000d40 ),
    .O(\blk000001fe/sig00000d2a )
  );
  XORCY   \blk000001fe/blk00000211  (
    .CI(\blk000001fe/sig00000d54 ),
    .LI(\blk000001fe/sig00000d3f ),
    .O(\blk000001fe/sig00000d29 )
  );
  XORCY   \blk000001fe/blk00000210  (
    .CI(\blk000001fe/sig00000d53 ),
    .LI(\blk000001fe/sig00000d3e ),
    .O(\blk000001fe/sig00000d28 )
  );
  XORCY   \blk000001fe/blk0000020f  (
    .CI(\blk000001fe/sig00000d52 ),
    .LI(\blk000001fe/sig00000d3d ),
    .O(\blk000001fe/sig00000d27 )
  );
  XORCY   \blk000001fe/blk0000020e  (
    .CI(\blk000001fe/sig00000d51 ),
    .LI(\blk000001fe/sig00000d3c ),
    .O(\blk000001fe/sig00000d26 )
  );
  XORCY   \blk000001fe/blk0000020d  (
    .CI(\blk000001fe/sig00000d50 ),
    .LI(\blk000001fe/sig00000d3b ),
    .O(\blk000001fe/sig00000d25 )
  );
  XORCY   \blk000001fe/blk0000020c  (
    .CI(\blk000001fe/sig00000d4f ),
    .LI(\blk000001fe/sig00000d3a ),
    .O(\blk000001fe/sig00000d24 )
  );
  XORCY   \blk000001fe/blk0000020b  (
    .CI(\blk000001fe/sig00000d4e ),
    .LI(\blk000001fe/sig00000d39 ),
    .O(\blk000001fe/sig00000d23 )
  );
  XORCY   \blk000001fe/blk0000020a  (
    .CI(\blk000001fe/sig00000d4d ),
    .LI(\blk000001fe/sig00000d38 ),
    .O(\blk000001fe/sig00000d22 )
  );
  XORCY   \blk000001fe/blk00000209  (
    .CI(\blk000001fe/sig00000d4c ),
    .LI(\blk000001fe/sig00000d37 ),
    .O(\blk000001fe/sig00000d21 )
  );
  XORCY   \blk000001fe/blk00000208  (
    .CI(\blk000001fe/sig00000d4b ),
    .LI(\blk000001fe/sig00000d36 ),
    .O(\blk000001fe/sig00000d20 )
  );
  XORCY   \blk000001fe/blk00000207  (
    .CI(\blk000001fe/sig00000d4a ),
    .LI(\blk000001fe/sig00000d35 ),
    .O(\blk000001fe/sig00000d1f )
  );
  XORCY   \blk000001fe/blk00000206  (
    .CI(\blk000001fe/sig00000d49 ),
    .LI(\blk000001fe/sig00000d34 ),
    .O(\blk000001fe/sig00000d1e )
  );
  XORCY   \blk000001fe/blk00000205  (
    .CI(\blk000001fe/sig00000d48 ),
    .LI(\blk000001fe/sig00000d33 ),
    .O(\blk000001fe/sig00000d1d )
  );
  XORCY   \blk000001fe/blk00000204  (
    .CI(\blk000001fe/sig00000d47 ),
    .LI(\blk000001fe/sig00000d32 ),
    .O(\blk000001fe/sig00000d1c )
  );
  XORCY   \blk000001fe/blk00000203  (
    .CI(\blk000001fe/sig00000d46 ),
    .LI(\blk000001fe/sig00000d31 ),
    .O(\blk000001fe/sig00000d1b )
  );
  XORCY   \blk000001fe/blk00000202  (
    .CI(\blk000001fe/sig00000d45 ),
    .LI(\blk000001fe/sig00000d5b ),
    .O(\NLW_blk000001fe/blk00000202_O_UNCONNECTED )
  );
  XORCY   \blk000001fe/blk00000201  (
    .CI(\blk000001fe/sig00000d44 ),
    .LI(\blk000001fe/sig00000d30 ),
    .O(\NLW_blk000001fe/blk00000201_O_UNCONNECTED )
  );
  XORCY   \blk000001fe/blk00000200  (
    .CI(\blk000001fe/sig00000d19 ),
    .LI(\blk000001fe/sig00000d5e ),
    .O(\blk000001fe/sig00000d1a )
  );
  GND   \blk000001fe/blk000001ff  (
    .G(\blk000001fe/sig00000d19 )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk0000025d/blk000002bb  (
    .I0(sig000001b0),
    .O(\blk0000025d/sig00000dea )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk0000025d/blk000002ba  (
    .I0(sig000001b1),
    .O(\blk0000025d/sig00000de9 )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk0000025d/blk000002b9  (
    .I0(sig000001b2),
    .O(\blk0000025d/sig00000de8 )
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  \blk0000025d/blk000002b8  (
    .I0(sig00000272),
    .I1(sig000001c6),
    .O(\blk0000025d/sig00000de7 )
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  \blk0000025d/blk000002b7  (
    .I0(sig00000272),
    .I1(sig000001c6),
    .O(\blk0000025d/sig00000dbc )
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  \blk0000025d/blk000002b6  (
    .I0(sig00000272),
    .I1(sig000001c5),
    .O(\blk0000025d/sig00000dbd )
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  \blk0000025d/blk000002b5  (
    .I0(sig00000271),
    .I1(sig000001c4),
    .O(\blk0000025d/sig00000dbe )
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  \blk0000025d/blk000002b4  (
    .I0(sig00000270),
    .I1(sig000001c3),
    .O(\blk0000025d/sig00000dbf )
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  \blk0000025d/blk000002b3  (
    .I0(sig0000026f),
    .I1(sig000001c2),
    .O(\blk0000025d/sig00000dc0 )
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  \blk0000025d/blk000002b2  (
    .I0(sig0000026e),
    .I1(sig000001c1),
    .O(\blk0000025d/sig00000dc1 )
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  \blk0000025d/blk000002b1  (
    .I0(sig0000026d),
    .I1(sig000001c0),
    .O(\blk0000025d/sig00000dc2 )
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  \blk0000025d/blk000002b0  (
    .I0(sig0000026c),
    .I1(sig000001bf),
    .O(\blk0000025d/sig00000dc3 )
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  \blk0000025d/blk000002af  (
    .I0(sig0000026b),
    .I1(sig000001be),
    .O(\blk0000025d/sig00000dc4 )
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  \blk0000025d/blk000002ae  (
    .I0(sig0000026a),
    .I1(sig000001bd),
    .O(\blk0000025d/sig00000dc5 )
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  \blk0000025d/blk000002ad  (
    .I0(sig00000269),
    .I1(sig000001bc),
    .O(\blk0000025d/sig00000dc6 )
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  \blk0000025d/blk000002ac  (
    .I0(sig00000268),
    .I1(sig000001bb),
    .O(\blk0000025d/sig00000dc7 )
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  \blk0000025d/blk000002ab  (
    .I0(sig00000267),
    .I1(sig000001ba),
    .O(\blk0000025d/sig00000dc8 )
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  \blk0000025d/blk000002aa  (
    .I0(sig00000266),
    .I1(sig000001b9),
    .O(\blk0000025d/sig00000dc9 )
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  \blk0000025d/blk000002a9  (
    .I0(sig00000265),
    .I1(sig000001b8),
    .O(\blk0000025d/sig00000dca )
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  \blk0000025d/blk000002a8  (
    .I0(sig00000264),
    .I1(sig000001b7),
    .O(\blk0000025d/sig00000dcb )
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  \blk0000025d/blk000002a7  (
    .I0(sig00000263),
    .I1(sig000001b6),
    .O(\blk0000025d/sig00000dcc )
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  \blk0000025d/blk000002a6  (
    .I0(sig00000262),
    .I1(sig000001b5),
    .O(\blk0000025d/sig00000dcd )
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  \blk0000025d/blk000002a5  (
    .I0(sig00000261),
    .I1(sig000001b4),
    .O(\blk0000025d/sig00000dce )
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  \blk0000025d/blk000002a4  (
    .I0(sig00000260),
    .I1(sig000001b3),
    .O(\blk0000025d/sig00000dcf )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk0000025d/blk000002a3  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk0000025d/sig00000da6 ),
    .Q(sig000001f3)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk0000025d/blk000002a2  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk0000025d/sig00000dbb ),
    .Q(sig000001f4)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk0000025d/blk000002a1  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk0000025d/sig00000dba ),
    .Q(sig000001f5)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk0000025d/blk000002a0  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk0000025d/sig00000db9 ),
    .Q(sig000001f6)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk0000025d/blk0000029f  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk0000025d/sig00000db8 ),
    .Q(sig000001f7)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk0000025d/blk0000029e  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk0000025d/sig00000db7 ),
    .Q(sig000001f8)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk0000025d/blk0000029d  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk0000025d/sig00000db6 ),
    .Q(sig000001f9)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk0000025d/blk0000029c  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk0000025d/sig00000db5 ),
    .Q(sig000001fa)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk0000025d/blk0000029b  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk0000025d/sig00000db4 ),
    .Q(sig000001fb)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk0000025d/blk0000029a  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk0000025d/sig00000db3 ),
    .Q(sig000001fc)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk0000025d/blk00000299  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk0000025d/sig00000db2 ),
    .Q(sig000001fd)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk0000025d/blk00000298  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk0000025d/sig00000db1 ),
    .Q(sig000001fe)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk0000025d/blk00000297  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk0000025d/sig00000db0 ),
    .Q(sig000001ff)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk0000025d/blk00000296  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk0000025d/sig00000daf ),
    .Q(sig00000200)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk0000025d/blk00000295  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk0000025d/sig00000dae ),
    .Q(sig00000201)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk0000025d/blk00000294  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk0000025d/sig00000dad ),
    .Q(sig00000202)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk0000025d/blk00000293  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk0000025d/sig00000dac ),
    .Q(sig00000203)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk0000025d/blk00000292  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk0000025d/sig00000dab ),
    .Q(sig00000204)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk0000025d/blk00000291  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk0000025d/sig00000daa ),
    .Q(sig00000205)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk0000025d/blk00000290  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk0000025d/sig00000da9 ),
    .Q(sig00000206)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk0000025d/blk0000028f  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk0000025d/sig00000da8 ),
    .Q(sig00000207)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk0000025d/blk0000028e  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk0000025d/sig00000da7 ),
    .Q(sig00000208)
  );
  MUXCY   \blk0000025d/blk0000028d  (
    .CI(\blk0000025d/sig00000da5 ),
    .DI(sig00000002),
    .S(\blk0000025d/sig00000dea ),
    .O(\blk0000025d/sig00000de6 )
  );
  MUXCY   \blk0000025d/blk0000028c  (
    .CI(\blk0000025d/sig00000de6 ),
    .DI(sig00000002),
    .S(\blk0000025d/sig00000de9 ),
    .O(\blk0000025d/sig00000de5 )
  );
  MUXCY   \blk0000025d/blk0000028b  (
    .CI(\blk0000025d/sig00000de5 ),
    .DI(sig00000002),
    .S(\blk0000025d/sig00000de8 ),
    .O(\blk0000025d/sig00000de4 )
  );
  MUXCY   \blk0000025d/blk0000028a  (
    .CI(\blk0000025d/sig00000de4 ),
    .DI(sig00000260),
    .S(\blk0000025d/sig00000dcf ),
    .O(\blk0000025d/sig00000de3 )
  );
  MUXCY   \blk0000025d/blk00000289  (
    .CI(\blk0000025d/sig00000de3 ),
    .DI(sig00000261),
    .S(\blk0000025d/sig00000dce ),
    .O(\blk0000025d/sig00000de2 )
  );
  MUXCY   \blk0000025d/blk00000288  (
    .CI(\blk0000025d/sig00000de2 ),
    .DI(sig00000262),
    .S(\blk0000025d/sig00000dcd ),
    .O(\blk0000025d/sig00000de1 )
  );
  MUXCY   \blk0000025d/blk00000287  (
    .CI(\blk0000025d/sig00000de1 ),
    .DI(sig00000263),
    .S(\blk0000025d/sig00000dcc ),
    .O(\blk0000025d/sig00000de0 )
  );
  MUXCY   \blk0000025d/blk00000286  (
    .CI(\blk0000025d/sig00000de0 ),
    .DI(sig00000264),
    .S(\blk0000025d/sig00000dcb ),
    .O(\blk0000025d/sig00000ddf )
  );
  MUXCY   \blk0000025d/blk00000285  (
    .CI(\blk0000025d/sig00000ddf ),
    .DI(sig00000265),
    .S(\blk0000025d/sig00000dca ),
    .O(\blk0000025d/sig00000dde )
  );
  MUXCY   \blk0000025d/blk00000284  (
    .CI(\blk0000025d/sig00000dde ),
    .DI(sig00000266),
    .S(\blk0000025d/sig00000dc9 ),
    .O(\blk0000025d/sig00000ddd )
  );
  MUXCY   \blk0000025d/blk00000283  (
    .CI(\blk0000025d/sig00000ddd ),
    .DI(sig00000267),
    .S(\blk0000025d/sig00000dc8 ),
    .O(\blk0000025d/sig00000ddc )
  );
  MUXCY   \blk0000025d/blk00000282  (
    .CI(\blk0000025d/sig00000ddc ),
    .DI(sig00000268),
    .S(\blk0000025d/sig00000dc7 ),
    .O(\blk0000025d/sig00000ddb )
  );
  MUXCY   \blk0000025d/blk00000281  (
    .CI(\blk0000025d/sig00000ddb ),
    .DI(sig00000269),
    .S(\blk0000025d/sig00000dc6 ),
    .O(\blk0000025d/sig00000dda )
  );
  MUXCY   \blk0000025d/blk00000280  (
    .CI(\blk0000025d/sig00000dda ),
    .DI(sig0000026a),
    .S(\blk0000025d/sig00000dc5 ),
    .O(\blk0000025d/sig00000dd9 )
  );
  MUXCY   \blk0000025d/blk0000027f  (
    .CI(\blk0000025d/sig00000dd9 ),
    .DI(sig0000026b),
    .S(\blk0000025d/sig00000dc4 ),
    .O(\blk0000025d/sig00000dd8 )
  );
  MUXCY   \blk0000025d/blk0000027e  (
    .CI(\blk0000025d/sig00000dd8 ),
    .DI(sig0000026c),
    .S(\blk0000025d/sig00000dc3 ),
    .O(\blk0000025d/sig00000dd7 )
  );
  MUXCY   \blk0000025d/blk0000027d  (
    .CI(\blk0000025d/sig00000dd7 ),
    .DI(sig0000026d),
    .S(\blk0000025d/sig00000dc2 ),
    .O(\blk0000025d/sig00000dd6 )
  );
  MUXCY   \blk0000025d/blk0000027c  (
    .CI(\blk0000025d/sig00000dd6 ),
    .DI(sig0000026e),
    .S(\blk0000025d/sig00000dc1 ),
    .O(\blk0000025d/sig00000dd5 )
  );
  MUXCY   \blk0000025d/blk0000027b  (
    .CI(\blk0000025d/sig00000dd5 ),
    .DI(sig0000026f),
    .S(\blk0000025d/sig00000dc0 ),
    .O(\blk0000025d/sig00000dd4 )
  );
  MUXCY   \blk0000025d/blk0000027a  (
    .CI(\blk0000025d/sig00000dd4 ),
    .DI(sig00000270),
    .S(\blk0000025d/sig00000dbf ),
    .O(\blk0000025d/sig00000dd3 )
  );
  MUXCY   \blk0000025d/blk00000279  (
    .CI(\blk0000025d/sig00000dd3 ),
    .DI(sig00000271),
    .S(\blk0000025d/sig00000dbe ),
    .O(\blk0000025d/sig00000dd2 )
  );
  MUXCY   \blk0000025d/blk00000278  (
    .CI(\blk0000025d/sig00000dd2 ),
    .DI(sig00000272),
    .S(\blk0000025d/sig00000dbd ),
    .O(\blk0000025d/sig00000dd1 )
  );
  MUXCY   \blk0000025d/blk00000277  (
    .CI(\blk0000025d/sig00000dd1 ),
    .DI(sig00000272),
    .S(\blk0000025d/sig00000de7 ),
    .O(\blk0000025d/sig00000dd0 )
  );
  XORCY   \blk0000025d/blk00000276  (
    .CI(\blk0000025d/sig00000de6 ),
    .LI(\blk0000025d/sig00000de9 ),
    .O(\blk0000025d/sig00000dbb )
  );
  XORCY   \blk0000025d/blk00000275  (
    .CI(\blk0000025d/sig00000de5 ),
    .LI(\blk0000025d/sig00000de8 ),
    .O(\blk0000025d/sig00000dba )
  );
  XORCY   \blk0000025d/blk00000274  (
    .CI(\blk0000025d/sig00000de4 ),
    .LI(\blk0000025d/sig00000dcf ),
    .O(\blk0000025d/sig00000db9 )
  );
  XORCY   \blk0000025d/blk00000273  (
    .CI(\blk0000025d/sig00000de3 ),
    .LI(\blk0000025d/sig00000dce ),
    .O(\blk0000025d/sig00000db8 )
  );
  XORCY   \blk0000025d/blk00000272  (
    .CI(\blk0000025d/sig00000de2 ),
    .LI(\blk0000025d/sig00000dcd ),
    .O(\blk0000025d/sig00000db7 )
  );
  XORCY   \blk0000025d/blk00000271  (
    .CI(\blk0000025d/sig00000de1 ),
    .LI(\blk0000025d/sig00000dcc ),
    .O(\blk0000025d/sig00000db6 )
  );
  XORCY   \blk0000025d/blk00000270  (
    .CI(\blk0000025d/sig00000de0 ),
    .LI(\blk0000025d/sig00000dcb ),
    .O(\blk0000025d/sig00000db5 )
  );
  XORCY   \blk0000025d/blk0000026f  (
    .CI(\blk0000025d/sig00000ddf ),
    .LI(\blk0000025d/sig00000dca ),
    .O(\blk0000025d/sig00000db4 )
  );
  XORCY   \blk0000025d/blk0000026e  (
    .CI(\blk0000025d/sig00000dde ),
    .LI(\blk0000025d/sig00000dc9 ),
    .O(\blk0000025d/sig00000db3 )
  );
  XORCY   \blk0000025d/blk0000026d  (
    .CI(\blk0000025d/sig00000ddd ),
    .LI(\blk0000025d/sig00000dc8 ),
    .O(\blk0000025d/sig00000db2 )
  );
  XORCY   \blk0000025d/blk0000026c  (
    .CI(\blk0000025d/sig00000ddc ),
    .LI(\blk0000025d/sig00000dc7 ),
    .O(\blk0000025d/sig00000db1 )
  );
  XORCY   \blk0000025d/blk0000026b  (
    .CI(\blk0000025d/sig00000ddb ),
    .LI(\blk0000025d/sig00000dc6 ),
    .O(\blk0000025d/sig00000db0 )
  );
  XORCY   \blk0000025d/blk0000026a  (
    .CI(\blk0000025d/sig00000dda ),
    .LI(\blk0000025d/sig00000dc5 ),
    .O(\blk0000025d/sig00000daf )
  );
  XORCY   \blk0000025d/blk00000269  (
    .CI(\blk0000025d/sig00000dd9 ),
    .LI(\blk0000025d/sig00000dc4 ),
    .O(\blk0000025d/sig00000dae )
  );
  XORCY   \blk0000025d/blk00000268  (
    .CI(\blk0000025d/sig00000dd8 ),
    .LI(\blk0000025d/sig00000dc3 ),
    .O(\blk0000025d/sig00000dad )
  );
  XORCY   \blk0000025d/blk00000267  (
    .CI(\blk0000025d/sig00000dd7 ),
    .LI(\blk0000025d/sig00000dc2 ),
    .O(\blk0000025d/sig00000dac )
  );
  XORCY   \blk0000025d/blk00000266  (
    .CI(\blk0000025d/sig00000dd6 ),
    .LI(\blk0000025d/sig00000dc1 ),
    .O(\blk0000025d/sig00000dab )
  );
  XORCY   \blk0000025d/blk00000265  (
    .CI(\blk0000025d/sig00000dd5 ),
    .LI(\blk0000025d/sig00000dc0 ),
    .O(\blk0000025d/sig00000daa )
  );
  XORCY   \blk0000025d/blk00000264  (
    .CI(\blk0000025d/sig00000dd4 ),
    .LI(\blk0000025d/sig00000dbf ),
    .O(\blk0000025d/sig00000da9 )
  );
  XORCY   \blk0000025d/blk00000263  (
    .CI(\blk0000025d/sig00000dd3 ),
    .LI(\blk0000025d/sig00000dbe ),
    .O(\blk0000025d/sig00000da8 )
  );
  XORCY   \blk0000025d/blk00000262  (
    .CI(\blk0000025d/sig00000dd2 ),
    .LI(\blk0000025d/sig00000dbd ),
    .O(\blk0000025d/sig00000da7 )
  );
  XORCY   \blk0000025d/blk00000261  (
    .CI(\blk0000025d/sig00000dd1 ),
    .LI(\blk0000025d/sig00000de7 ),
    .O(\NLW_blk0000025d/blk00000261_O_UNCONNECTED )
  );
  XORCY   \blk0000025d/blk00000260  (
    .CI(\blk0000025d/sig00000dd0 ),
    .LI(\blk0000025d/sig00000dbc ),
    .O(\NLW_blk0000025d/blk00000260_O_UNCONNECTED )
  );
  XORCY   \blk0000025d/blk0000025f  (
    .CI(\blk0000025d/sig00000da5 ),
    .LI(\blk0000025d/sig00000dea ),
    .O(\blk0000025d/sig00000da6 )
  );
  GND   \blk0000025d/blk0000025e  (
    .G(\blk0000025d/sig00000da5 )
  );
  INV   \blk000002bc/blk0000031a  (
    .I(sig0000019b),
    .O(\blk000002bc/sig00000e5c )
  );
  INV   \blk000002bc/blk00000319  (
    .I(sig0000019a),
    .O(\blk000002bc/sig00000e5d )
  );
  INV   \blk000002bc/blk00000318  (
    .I(sig00000199),
    .O(\blk000002bc/sig00000e5e )
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  \blk000002bc/blk00000317  (
    .I0(sig0000025f),
    .I1(sig000001af),
    .O(\blk000002bc/sig00000e76 )
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  \blk000002bc/blk00000316  (
    .I0(sig0000025f),
    .I1(sig000001af),
    .O(\blk000002bc/sig00000e48 )
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  \blk000002bc/blk00000315  (
    .I0(sig0000025f),
    .I1(sig000001ae),
    .O(\blk000002bc/sig00000e49 )
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  \blk000002bc/blk00000314  (
    .I0(sig0000025e),
    .I1(sig000001ad),
    .O(\blk000002bc/sig00000e4a )
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  \blk000002bc/blk00000313  (
    .I0(sig0000025d),
    .I1(sig000001ac),
    .O(\blk000002bc/sig00000e4b )
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  \blk000002bc/blk00000312  (
    .I0(sig0000025c),
    .I1(sig000001ab),
    .O(\blk000002bc/sig00000e4c )
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  \blk000002bc/blk00000311  (
    .I0(sig0000025b),
    .I1(sig000001aa),
    .O(\blk000002bc/sig00000e4d )
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  \blk000002bc/blk00000310  (
    .I0(sig0000025a),
    .I1(sig000001a9),
    .O(\blk000002bc/sig00000e4e )
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  \blk000002bc/blk0000030f  (
    .I0(sig00000259),
    .I1(sig000001a8),
    .O(\blk000002bc/sig00000e4f )
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  \blk000002bc/blk0000030e  (
    .I0(sig00000258),
    .I1(sig000001a7),
    .O(\blk000002bc/sig00000e50 )
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  \blk000002bc/blk0000030d  (
    .I0(sig00000257),
    .I1(sig000001a6),
    .O(\blk000002bc/sig00000e51 )
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  \blk000002bc/blk0000030c  (
    .I0(sig00000256),
    .I1(sig000001a5),
    .O(\blk000002bc/sig00000e52 )
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  \blk000002bc/blk0000030b  (
    .I0(sig00000255),
    .I1(sig000001a4),
    .O(\blk000002bc/sig00000e53 )
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  \blk000002bc/blk0000030a  (
    .I0(sig00000254),
    .I1(sig000001a3),
    .O(\blk000002bc/sig00000e54 )
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  \blk000002bc/blk00000309  (
    .I0(sig00000253),
    .I1(sig000001a2),
    .O(\blk000002bc/sig00000e55 )
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  \blk000002bc/blk00000308  (
    .I0(sig00000252),
    .I1(sig000001a1),
    .O(\blk000002bc/sig00000e56 )
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  \blk000002bc/blk00000307  (
    .I0(sig00000251),
    .I1(sig000001a0),
    .O(\blk000002bc/sig00000e57 )
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  \blk000002bc/blk00000306  (
    .I0(sig00000250),
    .I1(sig0000019f),
    .O(\blk000002bc/sig00000e58 )
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  \blk000002bc/blk00000305  (
    .I0(sig0000024f),
    .I1(sig0000019e),
    .O(\blk000002bc/sig00000e59 )
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  \blk000002bc/blk00000304  (
    .I0(sig0000024e),
    .I1(sig0000019d),
    .O(\blk000002bc/sig00000e5a )
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  \blk000002bc/blk00000303  (
    .I0(sig0000024d),
    .I1(sig0000019c),
    .O(\blk000002bc/sig00000e5b )
  );
  MUXCY   \blk000002bc/blk00000302  (
    .CI(\blk000002bc/sig00000e31 ),
    .DI(sig00000002),
    .S(\blk000002bc/sig00000e5e ),
    .O(\blk000002bc/sig00000e75 )
  );
  MUXCY   \blk000002bc/blk00000301  (
    .CI(\blk000002bc/sig00000e75 ),
    .DI(sig00000002),
    .S(\blk000002bc/sig00000e5d ),
    .O(\blk000002bc/sig00000e74 )
  );
  MUXCY   \blk000002bc/blk00000300  (
    .CI(\blk000002bc/sig00000e74 ),
    .DI(sig00000002),
    .S(\blk000002bc/sig00000e5c ),
    .O(\blk000002bc/sig00000e73 )
  );
  MUXCY   \blk000002bc/blk000002ff  (
    .CI(\blk000002bc/sig00000e73 ),
    .DI(sig0000024d),
    .S(\blk000002bc/sig00000e5b ),
    .O(\blk000002bc/sig00000e72 )
  );
  MUXCY   \blk000002bc/blk000002fe  (
    .CI(\blk000002bc/sig00000e72 ),
    .DI(sig0000024e),
    .S(\blk000002bc/sig00000e5a ),
    .O(\blk000002bc/sig00000e71 )
  );
  MUXCY   \blk000002bc/blk000002fd  (
    .CI(\blk000002bc/sig00000e71 ),
    .DI(sig0000024f),
    .S(\blk000002bc/sig00000e59 ),
    .O(\blk000002bc/sig00000e70 )
  );
  MUXCY   \blk000002bc/blk000002fc  (
    .CI(\blk000002bc/sig00000e70 ),
    .DI(sig00000250),
    .S(\blk000002bc/sig00000e58 ),
    .O(\blk000002bc/sig00000e6f )
  );
  MUXCY   \blk000002bc/blk000002fb  (
    .CI(\blk000002bc/sig00000e6f ),
    .DI(sig00000251),
    .S(\blk000002bc/sig00000e57 ),
    .O(\blk000002bc/sig00000e6e )
  );
  MUXCY   \blk000002bc/blk000002fa  (
    .CI(\blk000002bc/sig00000e6e ),
    .DI(sig00000252),
    .S(\blk000002bc/sig00000e56 ),
    .O(\blk000002bc/sig00000e6d )
  );
  MUXCY   \blk000002bc/blk000002f9  (
    .CI(\blk000002bc/sig00000e6d ),
    .DI(sig00000253),
    .S(\blk000002bc/sig00000e55 ),
    .O(\blk000002bc/sig00000e6c )
  );
  MUXCY   \blk000002bc/blk000002f8  (
    .CI(\blk000002bc/sig00000e6c ),
    .DI(sig00000254),
    .S(\blk000002bc/sig00000e54 ),
    .O(\blk000002bc/sig00000e6b )
  );
  MUXCY   \blk000002bc/blk000002f7  (
    .CI(\blk000002bc/sig00000e6b ),
    .DI(sig00000255),
    .S(\blk000002bc/sig00000e53 ),
    .O(\blk000002bc/sig00000e6a )
  );
  MUXCY   \blk000002bc/blk000002f6  (
    .CI(\blk000002bc/sig00000e6a ),
    .DI(sig00000256),
    .S(\blk000002bc/sig00000e52 ),
    .O(\blk000002bc/sig00000e69 )
  );
  MUXCY   \blk000002bc/blk000002f5  (
    .CI(\blk000002bc/sig00000e69 ),
    .DI(sig00000257),
    .S(\blk000002bc/sig00000e51 ),
    .O(\blk000002bc/sig00000e68 )
  );
  MUXCY   \blk000002bc/blk000002f4  (
    .CI(\blk000002bc/sig00000e68 ),
    .DI(sig00000258),
    .S(\blk000002bc/sig00000e50 ),
    .O(\blk000002bc/sig00000e67 )
  );
  MUXCY   \blk000002bc/blk000002f3  (
    .CI(\blk000002bc/sig00000e67 ),
    .DI(sig00000259),
    .S(\blk000002bc/sig00000e4f ),
    .O(\blk000002bc/sig00000e66 )
  );
  MUXCY   \blk000002bc/blk000002f2  (
    .CI(\blk000002bc/sig00000e66 ),
    .DI(sig0000025a),
    .S(\blk000002bc/sig00000e4e ),
    .O(\blk000002bc/sig00000e65 )
  );
  MUXCY   \blk000002bc/blk000002f1  (
    .CI(\blk000002bc/sig00000e65 ),
    .DI(sig0000025b),
    .S(\blk000002bc/sig00000e4d ),
    .O(\blk000002bc/sig00000e64 )
  );
  MUXCY   \blk000002bc/blk000002f0  (
    .CI(\blk000002bc/sig00000e64 ),
    .DI(sig0000025c),
    .S(\blk000002bc/sig00000e4c ),
    .O(\blk000002bc/sig00000e63 )
  );
  MUXCY   \blk000002bc/blk000002ef  (
    .CI(\blk000002bc/sig00000e63 ),
    .DI(sig0000025d),
    .S(\blk000002bc/sig00000e4b ),
    .O(\blk000002bc/sig00000e62 )
  );
  MUXCY   \blk000002bc/blk000002ee  (
    .CI(\blk000002bc/sig00000e62 ),
    .DI(sig0000025e),
    .S(\blk000002bc/sig00000e4a ),
    .O(\blk000002bc/sig00000e61 )
  );
  MUXCY   \blk000002bc/blk000002ed  (
    .CI(\blk000002bc/sig00000e61 ),
    .DI(sig0000025f),
    .S(\blk000002bc/sig00000e49 ),
    .O(\blk000002bc/sig00000e60 )
  );
  MUXCY   \blk000002bc/blk000002ec  (
    .CI(\blk000002bc/sig00000e60 ),
    .DI(sig0000025f),
    .S(\blk000002bc/sig00000e76 ),
    .O(\blk000002bc/sig00000e5f )
  );
  XORCY   \blk000002bc/blk000002eb  (
    .CI(\blk000002bc/sig00000e75 ),
    .LI(\blk000002bc/sig00000e5d ),
    .O(\blk000002bc/sig00000e47 )
  );
  XORCY   \blk000002bc/blk000002ea  (
    .CI(\blk000002bc/sig00000e74 ),
    .LI(\blk000002bc/sig00000e5c ),
    .O(\blk000002bc/sig00000e46 )
  );
  XORCY   \blk000002bc/blk000002e9  (
    .CI(\blk000002bc/sig00000e73 ),
    .LI(\blk000002bc/sig00000e5b ),
    .O(\blk000002bc/sig00000e45 )
  );
  XORCY   \blk000002bc/blk000002e8  (
    .CI(\blk000002bc/sig00000e72 ),
    .LI(\blk000002bc/sig00000e5a ),
    .O(\blk000002bc/sig00000e44 )
  );
  XORCY   \blk000002bc/blk000002e7  (
    .CI(\blk000002bc/sig00000e71 ),
    .LI(\blk000002bc/sig00000e59 ),
    .O(\blk000002bc/sig00000e43 )
  );
  XORCY   \blk000002bc/blk000002e6  (
    .CI(\blk000002bc/sig00000e70 ),
    .LI(\blk000002bc/sig00000e58 ),
    .O(\blk000002bc/sig00000e42 )
  );
  XORCY   \blk000002bc/blk000002e5  (
    .CI(\blk000002bc/sig00000e6f ),
    .LI(\blk000002bc/sig00000e57 ),
    .O(\blk000002bc/sig00000e41 )
  );
  XORCY   \blk000002bc/blk000002e4  (
    .CI(\blk000002bc/sig00000e6e ),
    .LI(\blk000002bc/sig00000e56 ),
    .O(\blk000002bc/sig00000e40 )
  );
  XORCY   \blk000002bc/blk000002e3  (
    .CI(\blk000002bc/sig00000e6d ),
    .LI(\blk000002bc/sig00000e55 ),
    .O(\blk000002bc/sig00000e3f )
  );
  XORCY   \blk000002bc/blk000002e2  (
    .CI(\blk000002bc/sig00000e6c ),
    .LI(\blk000002bc/sig00000e54 ),
    .O(\blk000002bc/sig00000e3e )
  );
  XORCY   \blk000002bc/blk000002e1  (
    .CI(\blk000002bc/sig00000e6b ),
    .LI(\blk000002bc/sig00000e53 ),
    .O(\blk000002bc/sig00000e3d )
  );
  XORCY   \blk000002bc/blk000002e0  (
    .CI(\blk000002bc/sig00000e6a ),
    .LI(\blk000002bc/sig00000e52 ),
    .O(\blk000002bc/sig00000e3c )
  );
  XORCY   \blk000002bc/blk000002df  (
    .CI(\blk000002bc/sig00000e69 ),
    .LI(\blk000002bc/sig00000e51 ),
    .O(\blk000002bc/sig00000e3b )
  );
  XORCY   \blk000002bc/blk000002de  (
    .CI(\blk000002bc/sig00000e68 ),
    .LI(\blk000002bc/sig00000e50 ),
    .O(\blk000002bc/sig00000e3a )
  );
  XORCY   \blk000002bc/blk000002dd  (
    .CI(\blk000002bc/sig00000e67 ),
    .LI(\blk000002bc/sig00000e4f ),
    .O(\blk000002bc/sig00000e39 )
  );
  XORCY   \blk000002bc/blk000002dc  (
    .CI(\blk000002bc/sig00000e66 ),
    .LI(\blk000002bc/sig00000e4e ),
    .O(\blk000002bc/sig00000e38 )
  );
  XORCY   \blk000002bc/blk000002db  (
    .CI(\blk000002bc/sig00000e65 ),
    .LI(\blk000002bc/sig00000e4d ),
    .O(\blk000002bc/sig00000e37 )
  );
  XORCY   \blk000002bc/blk000002da  (
    .CI(\blk000002bc/sig00000e64 ),
    .LI(\blk000002bc/sig00000e4c ),
    .O(\blk000002bc/sig00000e36 )
  );
  XORCY   \blk000002bc/blk000002d9  (
    .CI(\blk000002bc/sig00000e63 ),
    .LI(\blk000002bc/sig00000e4b ),
    .O(\blk000002bc/sig00000e35 )
  );
  XORCY   \blk000002bc/blk000002d8  (
    .CI(\blk000002bc/sig00000e62 ),
    .LI(\blk000002bc/sig00000e4a ),
    .O(\blk000002bc/sig00000e34 )
  );
  XORCY   \blk000002bc/blk000002d7  (
    .CI(\blk000002bc/sig00000e61 ),
    .LI(\blk000002bc/sig00000e49 ),
    .O(\blk000002bc/sig00000e33 )
  );
  XORCY   \blk000002bc/blk000002d6  (
    .CI(\blk000002bc/sig00000e60 ),
    .LI(\blk000002bc/sig00000e76 ),
    .O(\NLW_blk000002bc/blk000002d6_O_UNCONNECTED )
  );
  XORCY   \blk000002bc/blk000002d5  (
    .CI(\blk000002bc/sig00000e5f ),
    .LI(\blk000002bc/sig00000e48 ),
    .O(\NLW_blk000002bc/blk000002d5_O_UNCONNECTED )
  );
  XORCY   \blk000002bc/blk000002d4  (
    .CI(\blk000002bc/sig00000e31 ),
    .LI(\blk000002bc/sig00000e5e ),
    .O(\blk000002bc/sig00000e32 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000002bc/blk000002d3  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk000002bc/sig00000e33 ),
    .Q(sig000001f2)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000002bc/blk000002d2  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk000002bc/sig00000e34 ),
    .Q(sig000001f1)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000002bc/blk000002d1  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk000002bc/sig00000e35 ),
    .Q(sig000001f0)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000002bc/blk000002d0  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk000002bc/sig00000e36 ),
    .Q(sig000001ef)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000002bc/blk000002cf  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk000002bc/sig00000e37 ),
    .Q(sig000001ee)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000002bc/blk000002ce  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk000002bc/sig00000e38 ),
    .Q(sig000001ed)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000002bc/blk000002cd  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk000002bc/sig00000e39 ),
    .Q(sig000001ec)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000002bc/blk000002cc  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk000002bc/sig00000e3a ),
    .Q(sig000001eb)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000002bc/blk000002cb  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk000002bc/sig00000e3b ),
    .Q(sig000001ea)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000002bc/blk000002ca  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk000002bc/sig00000e3c ),
    .Q(sig000001e9)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000002bc/blk000002c9  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk000002bc/sig00000e3d ),
    .Q(sig000001e8)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000002bc/blk000002c8  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk000002bc/sig00000e3e ),
    .Q(sig000001e7)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000002bc/blk000002c7  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk000002bc/sig00000e3f ),
    .Q(sig000001e6)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000002bc/blk000002c6  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk000002bc/sig00000e40 ),
    .Q(sig000001e5)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000002bc/blk000002c5  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk000002bc/sig00000e41 ),
    .Q(sig000001e4)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000002bc/blk000002c4  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk000002bc/sig00000e42 ),
    .Q(sig000001e3)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000002bc/blk000002c3  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk000002bc/sig00000e43 ),
    .Q(sig000001e2)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000002bc/blk000002c2  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk000002bc/sig00000e44 ),
    .Q(sig000001e1)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000002bc/blk000002c1  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk000002bc/sig00000e45 ),
    .Q(sig000001e0)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000002bc/blk000002c0  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk000002bc/sig00000e46 ),
    .Q(sig000001df)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000002bc/blk000002bf  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk000002bc/sig00000e47 ),
    .Q(sig000001de)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000002bc/blk000002be  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk000002bc/sig00000e32 ),
    .Q(sig000001dd)
  );
  VCC   \blk000002bc/blk000002bd  (
    .P(\blk000002bc/sig00000e31 )
  );
  INV   \blk0000031b/blk00000379  (
    .I(sig000001b2),
    .O(\blk0000031b/sig00000ee8 )
  );
  INV   \blk0000031b/blk00000378  (
    .I(sig000001b1),
    .O(\blk0000031b/sig00000ee9 )
  );
  INV   \blk0000031b/blk00000377  (
    .I(sig000001b0),
    .O(\blk0000031b/sig00000eea )
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  \blk0000031b/blk00000376  (
    .I0(sig00000272),
    .I1(sig000001c6),
    .O(\blk0000031b/sig00000f02 )
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  \blk0000031b/blk00000375  (
    .I0(sig00000272),
    .I1(sig000001c6),
    .O(\blk0000031b/sig00000ed4 )
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  \blk0000031b/blk00000374  (
    .I0(sig00000272),
    .I1(sig000001c5),
    .O(\blk0000031b/sig00000ed5 )
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  \blk0000031b/blk00000373  (
    .I0(sig00000271),
    .I1(sig000001c4),
    .O(\blk0000031b/sig00000ed6 )
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  \blk0000031b/blk00000372  (
    .I0(sig00000270),
    .I1(sig000001c3),
    .O(\blk0000031b/sig00000ed7 )
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  \blk0000031b/blk00000371  (
    .I0(sig0000026f),
    .I1(sig000001c2),
    .O(\blk0000031b/sig00000ed8 )
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  \blk0000031b/blk00000370  (
    .I0(sig0000026e),
    .I1(sig000001c1),
    .O(\blk0000031b/sig00000ed9 )
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  \blk0000031b/blk0000036f  (
    .I0(sig0000026d),
    .I1(sig000001c0),
    .O(\blk0000031b/sig00000eda )
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  \blk0000031b/blk0000036e  (
    .I0(sig0000026c),
    .I1(sig000001bf),
    .O(\blk0000031b/sig00000edb )
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  \blk0000031b/blk0000036d  (
    .I0(sig0000026b),
    .I1(sig000001be),
    .O(\blk0000031b/sig00000edc )
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  \blk0000031b/blk0000036c  (
    .I0(sig0000026a),
    .I1(sig000001bd),
    .O(\blk0000031b/sig00000edd )
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  \blk0000031b/blk0000036b  (
    .I0(sig00000269),
    .I1(sig000001bc),
    .O(\blk0000031b/sig00000ede )
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  \blk0000031b/blk0000036a  (
    .I0(sig00000268),
    .I1(sig000001bb),
    .O(\blk0000031b/sig00000edf )
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  \blk0000031b/blk00000369  (
    .I0(sig00000267),
    .I1(sig000001ba),
    .O(\blk0000031b/sig00000ee0 )
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  \blk0000031b/blk00000368  (
    .I0(sig00000266),
    .I1(sig000001b9),
    .O(\blk0000031b/sig00000ee1 )
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  \blk0000031b/blk00000367  (
    .I0(sig00000265),
    .I1(sig000001b8),
    .O(\blk0000031b/sig00000ee2 )
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  \blk0000031b/blk00000366  (
    .I0(sig00000264),
    .I1(sig000001b7),
    .O(\blk0000031b/sig00000ee3 )
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  \blk0000031b/blk00000365  (
    .I0(sig00000263),
    .I1(sig000001b6),
    .O(\blk0000031b/sig00000ee4 )
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  \blk0000031b/blk00000364  (
    .I0(sig00000262),
    .I1(sig000001b5),
    .O(\blk0000031b/sig00000ee5 )
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  \blk0000031b/blk00000363  (
    .I0(sig00000261),
    .I1(sig000001b4),
    .O(\blk0000031b/sig00000ee6 )
  );
  LUT2 #(
    .INIT ( 4'h9 ))
  \blk0000031b/blk00000362  (
    .I0(sig00000260),
    .I1(sig000001b3),
    .O(\blk0000031b/sig00000ee7 )
  );
  MUXCY   \blk0000031b/blk00000361  (
    .CI(\blk0000031b/sig00000ebd ),
    .DI(sig00000002),
    .S(\blk0000031b/sig00000eea ),
    .O(\blk0000031b/sig00000f01 )
  );
  MUXCY   \blk0000031b/blk00000360  (
    .CI(\blk0000031b/sig00000f01 ),
    .DI(sig00000002),
    .S(\blk0000031b/sig00000ee9 ),
    .O(\blk0000031b/sig00000f00 )
  );
  MUXCY   \blk0000031b/blk0000035f  (
    .CI(\blk0000031b/sig00000f00 ),
    .DI(sig00000002),
    .S(\blk0000031b/sig00000ee8 ),
    .O(\blk0000031b/sig00000eff )
  );
  MUXCY   \blk0000031b/blk0000035e  (
    .CI(\blk0000031b/sig00000eff ),
    .DI(sig00000260),
    .S(\blk0000031b/sig00000ee7 ),
    .O(\blk0000031b/sig00000efe )
  );
  MUXCY   \blk0000031b/blk0000035d  (
    .CI(\blk0000031b/sig00000efe ),
    .DI(sig00000261),
    .S(\blk0000031b/sig00000ee6 ),
    .O(\blk0000031b/sig00000efd )
  );
  MUXCY   \blk0000031b/blk0000035c  (
    .CI(\blk0000031b/sig00000efd ),
    .DI(sig00000262),
    .S(\blk0000031b/sig00000ee5 ),
    .O(\blk0000031b/sig00000efc )
  );
  MUXCY   \blk0000031b/blk0000035b  (
    .CI(\blk0000031b/sig00000efc ),
    .DI(sig00000263),
    .S(\blk0000031b/sig00000ee4 ),
    .O(\blk0000031b/sig00000efb )
  );
  MUXCY   \blk0000031b/blk0000035a  (
    .CI(\blk0000031b/sig00000efb ),
    .DI(sig00000264),
    .S(\blk0000031b/sig00000ee3 ),
    .O(\blk0000031b/sig00000efa )
  );
  MUXCY   \blk0000031b/blk00000359  (
    .CI(\blk0000031b/sig00000efa ),
    .DI(sig00000265),
    .S(\blk0000031b/sig00000ee2 ),
    .O(\blk0000031b/sig00000ef9 )
  );
  MUXCY   \blk0000031b/blk00000358  (
    .CI(\blk0000031b/sig00000ef9 ),
    .DI(sig00000266),
    .S(\blk0000031b/sig00000ee1 ),
    .O(\blk0000031b/sig00000ef8 )
  );
  MUXCY   \blk0000031b/blk00000357  (
    .CI(\blk0000031b/sig00000ef8 ),
    .DI(sig00000267),
    .S(\blk0000031b/sig00000ee0 ),
    .O(\blk0000031b/sig00000ef7 )
  );
  MUXCY   \blk0000031b/blk00000356  (
    .CI(\blk0000031b/sig00000ef7 ),
    .DI(sig00000268),
    .S(\blk0000031b/sig00000edf ),
    .O(\blk0000031b/sig00000ef6 )
  );
  MUXCY   \blk0000031b/blk00000355  (
    .CI(\blk0000031b/sig00000ef6 ),
    .DI(sig00000269),
    .S(\blk0000031b/sig00000ede ),
    .O(\blk0000031b/sig00000ef5 )
  );
  MUXCY   \blk0000031b/blk00000354  (
    .CI(\blk0000031b/sig00000ef5 ),
    .DI(sig0000026a),
    .S(\blk0000031b/sig00000edd ),
    .O(\blk0000031b/sig00000ef4 )
  );
  MUXCY   \blk0000031b/blk00000353  (
    .CI(\blk0000031b/sig00000ef4 ),
    .DI(sig0000026b),
    .S(\blk0000031b/sig00000edc ),
    .O(\blk0000031b/sig00000ef3 )
  );
  MUXCY   \blk0000031b/blk00000352  (
    .CI(\blk0000031b/sig00000ef3 ),
    .DI(sig0000026c),
    .S(\blk0000031b/sig00000edb ),
    .O(\blk0000031b/sig00000ef2 )
  );
  MUXCY   \blk0000031b/blk00000351  (
    .CI(\blk0000031b/sig00000ef2 ),
    .DI(sig0000026d),
    .S(\blk0000031b/sig00000eda ),
    .O(\blk0000031b/sig00000ef1 )
  );
  MUXCY   \blk0000031b/blk00000350  (
    .CI(\blk0000031b/sig00000ef1 ),
    .DI(sig0000026e),
    .S(\blk0000031b/sig00000ed9 ),
    .O(\blk0000031b/sig00000ef0 )
  );
  MUXCY   \blk0000031b/blk0000034f  (
    .CI(\blk0000031b/sig00000ef0 ),
    .DI(sig0000026f),
    .S(\blk0000031b/sig00000ed8 ),
    .O(\blk0000031b/sig00000eef )
  );
  MUXCY   \blk0000031b/blk0000034e  (
    .CI(\blk0000031b/sig00000eef ),
    .DI(sig00000270),
    .S(\blk0000031b/sig00000ed7 ),
    .O(\blk0000031b/sig00000eee )
  );
  MUXCY   \blk0000031b/blk0000034d  (
    .CI(\blk0000031b/sig00000eee ),
    .DI(sig00000271),
    .S(\blk0000031b/sig00000ed6 ),
    .O(\blk0000031b/sig00000eed )
  );
  MUXCY   \blk0000031b/blk0000034c  (
    .CI(\blk0000031b/sig00000eed ),
    .DI(sig00000272),
    .S(\blk0000031b/sig00000ed5 ),
    .O(\blk0000031b/sig00000eec )
  );
  MUXCY   \blk0000031b/blk0000034b  (
    .CI(\blk0000031b/sig00000eec ),
    .DI(sig00000272),
    .S(\blk0000031b/sig00000f02 ),
    .O(\blk0000031b/sig00000eeb )
  );
  XORCY   \blk0000031b/blk0000034a  (
    .CI(\blk0000031b/sig00000f01 ),
    .LI(\blk0000031b/sig00000ee9 ),
    .O(\blk0000031b/sig00000ed3 )
  );
  XORCY   \blk0000031b/blk00000349  (
    .CI(\blk0000031b/sig00000f00 ),
    .LI(\blk0000031b/sig00000ee8 ),
    .O(\blk0000031b/sig00000ed2 )
  );
  XORCY   \blk0000031b/blk00000348  (
    .CI(\blk0000031b/sig00000eff ),
    .LI(\blk0000031b/sig00000ee7 ),
    .O(\blk0000031b/sig00000ed1 )
  );
  XORCY   \blk0000031b/blk00000347  (
    .CI(\blk0000031b/sig00000efe ),
    .LI(\blk0000031b/sig00000ee6 ),
    .O(\blk0000031b/sig00000ed0 )
  );
  XORCY   \blk0000031b/blk00000346  (
    .CI(\blk0000031b/sig00000efd ),
    .LI(\blk0000031b/sig00000ee5 ),
    .O(\blk0000031b/sig00000ecf )
  );
  XORCY   \blk0000031b/blk00000345  (
    .CI(\blk0000031b/sig00000efc ),
    .LI(\blk0000031b/sig00000ee4 ),
    .O(\blk0000031b/sig00000ece )
  );
  XORCY   \blk0000031b/blk00000344  (
    .CI(\blk0000031b/sig00000efb ),
    .LI(\blk0000031b/sig00000ee3 ),
    .O(\blk0000031b/sig00000ecd )
  );
  XORCY   \blk0000031b/blk00000343  (
    .CI(\blk0000031b/sig00000efa ),
    .LI(\blk0000031b/sig00000ee2 ),
    .O(\blk0000031b/sig00000ecc )
  );
  XORCY   \blk0000031b/blk00000342  (
    .CI(\blk0000031b/sig00000ef9 ),
    .LI(\blk0000031b/sig00000ee1 ),
    .O(\blk0000031b/sig00000ecb )
  );
  XORCY   \blk0000031b/blk00000341  (
    .CI(\blk0000031b/sig00000ef8 ),
    .LI(\blk0000031b/sig00000ee0 ),
    .O(\blk0000031b/sig00000eca )
  );
  XORCY   \blk0000031b/blk00000340  (
    .CI(\blk0000031b/sig00000ef7 ),
    .LI(\blk0000031b/sig00000edf ),
    .O(\blk0000031b/sig00000ec9 )
  );
  XORCY   \blk0000031b/blk0000033f  (
    .CI(\blk0000031b/sig00000ef6 ),
    .LI(\blk0000031b/sig00000ede ),
    .O(\blk0000031b/sig00000ec8 )
  );
  XORCY   \blk0000031b/blk0000033e  (
    .CI(\blk0000031b/sig00000ef5 ),
    .LI(\blk0000031b/sig00000edd ),
    .O(\blk0000031b/sig00000ec7 )
  );
  XORCY   \blk0000031b/blk0000033d  (
    .CI(\blk0000031b/sig00000ef4 ),
    .LI(\blk0000031b/sig00000edc ),
    .O(\blk0000031b/sig00000ec6 )
  );
  XORCY   \blk0000031b/blk0000033c  (
    .CI(\blk0000031b/sig00000ef3 ),
    .LI(\blk0000031b/sig00000edb ),
    .O(\blk0000031b/sig00000ec5 )
  );
  XORCY   \blk0000031b/blk0000033b  (
    .CI(\blk0000031b/sig00000ef2 ),
    .LI(\blk0000031b/sig00000eda ),
    .O(\blk0000031b/sig00000ec4 )
  );
  XORCY   \blk0000031b/blk0000033a  (
    .CI(\blk0000031b/sig00000ef1 ),
    .LI(\blk0000031b/sig00000ed9 ),
    .O(\blk0000031b/sig00000ec3 )
  );
  XORCY   \blk0000031b/blk00000339  (
    .CI(\blk0000031b/sig00000ef0 ),
    .LI(\blk0000031b/sig00000ed8 ),
    .O(\blk0000031b/sig00000ec2 )
  );
  XORCY   \blk0000031b/blk00000338  (
    .CI(\blk0000031b/sig00000eef ),
    .LI(\blk0000031b/sig00000ed7 ),
    .O(\blk0000031b/sig00000ec1 )
  );
  XORCY   \blk0000031b/blk00000337  (
    .CI(\blk0000031b/sig00000eee ),
    .LI(\blk0000031b/sig00000ed6 ),
    .O(\blk0000031b/sig00000ec0 )
  );
  XORCY   \blk0000031b/blk00000336  (
    .CI(\blk0000031b/sig00000eed ),
    .LI(\blk0000031b/sig00000ed5 ),
    .O(\blk0000031b/sig00000ebf )
  );
  XORCY   \blk0000031b/blk00000335  (
    .CI(\blk0000031b/sig00000eec ),
    .LI(\blk0000031b/sig00000f02 ),
    .O(\NLW_blk0000031b/blk00000335_O_UNCONNECTED )
  );
  XORCY   \blk0000031b/blk00000334  (
    .CI(\blk0000031b/sig00000eeb ),
    .LI(\blk0000031b/sig00000ed4 ),
    .O(\NLW_blk0000031b/blk00000334_O_UNCONNECTED )
  );
  XORCY   \blk0000031b/blk00000333  (
    .CI(\blk0000031b/sig00000ebd ),
    .LI(\blk0000031b/sig00000eea ),
    .O(\blk0000031b/sig00000ebe )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk0000031b/blk00000332  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk0000031b/sig00000ebf ),
    .Q(sig000001dc)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk0000031b/blk00000331  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk0000031b/sig00000ec0 ),
    .Q(sig000001db)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk0000031b/blk00000330  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk0000031b/sig00000ec1 ),
    .Q(sig000001da)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk0000031b/blk0000032f  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk0000031b/sig00000ec2 ),
    .Q(sig000001d9)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk0000031b/blk0000032e  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk0000031b/sig00000ec3 ),
    .Q(sig000001d8)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk0000031b/blk0000032d  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk0000031b/sig00000ec4 ),
    .Q(sig000001d7)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk0000031b/blk0000032c  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk0000031b/sig00000ec5 ),
    .Q(sig000001d6)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk0000031b/blk0000032b  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk0000031b/sig00000ec6 ),
    .Q(sig000001d5)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk0000031b/blk0000032a  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk0000031b/sig00000ec7 ),
    .Q(sig000001d4)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk0000031b/blk00000329  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk0000031b/sig00000ec8 ),
    .Q(sig000001d3)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk0000031b/blk00000328  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk0000031b/sig00000ec9 ),
    .Q(sig000001d2)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk0000031b/blk00000327  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk0000031b/sig00000eca ),
    .Q(sig000001d1)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk0000031b/blk00000326  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk0000031b/sig00000ecb ),
    .Q(sig000001d0)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk0000031b/blk00000325  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk0000031b/sig00000ecc ),
    .Q(sig000001cf)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk0000031b/blk00000324  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk0000031b/sig00000ecd ),
    .Q(sig000001ce)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk0000031b/blk00000323  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk0000031b/sig00000ece ),
    .Q(sig000001cd)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk0000031b/blk00000322  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk0000031b/sig00000ecf ),
    .Q(sig000001cc)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk0000031b/blk00000321  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk0000031b/sig00000ed0 ),
    .Q(sig000001cb)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk0000031b/blk00000320  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk0000031b/sig00000ed1 ),
    .Q(sig000001ca)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk0000031b/blk0000031f  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk0000031b/sig00000ed2 ),
    .Q(sig000001c9)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk0000031b/blk0000031e  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk0000031b/sig00000ed3 ),
    .Q(sig000001c8)
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk0000031b/blk0000031d  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk0000031b/sig00000ebe ),
    .Q(sig000001c7)
  );
  VCC   \blk0000031b/blk0000031c  (
    .P(\blk0000031b/sig00000ebd )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk0000049e/blk000004d6  (
    .I0(sig00000686),
    .O(\blk0000049e/sig00000f4e )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk0000049e/blk000004d5  (
    .I0(sig00000687),
    .O(\blk0000049e/sig00000f4d )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk0000049e/blk000004d4  (
    .I0(sig00000688),
    .O(\blk0000049e/sig00000f4c )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk0000049e/blk000004d3  (
    .I0(sig00000689),
    .O(\blk0000049e/sig00000f4b )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk0000049e/blk000004d2  (
    .I0(sig0000068a),
    .O(\blk0000049e/sig00000f4a )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk0000049e/blk000004d1  (
    .I0(sig0000068b),
    .O(\blk0000049e/sig00000f49 )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk0000049e/blk000004d0  (
    .I0(sig0000068c),
    .O(\blk0000049e/sig00000f48 )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk0000049e/blk000004cf  (
    .I0(sig0000068d),
    .O(\blk0000049e/sig00000f47 )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk0000049e/blk000004ce  (
    .I0(sig0000068e),
    .O(\blk0000049e/sig00000f46 )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk0000049e/blk000004cd  (
    .I0(sig0000068f),
    .O(\blk0000049e/sig00000f45 )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk0000049e/blk000004cc  (
    .I0(sig00000690),
    .O(\blk0000049e/sig00000f44 )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk0000049e/blk000004cb  (
    .I0(sig00000691),
    .O(\blk0000049e/sig00000f43 )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk0000049e/blk000004ca  (
    .I0(sig00000692),
    .O(\blk0000049e/sig00000f42 )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk0000049e/blk000004c9  (
    .I0(sig00000693),
    .O(\blk0000049e/sig00000f41 )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk0000049e/blk000004c8  (
    .I0(sig00000694),
    .O(\blk0000049e/sig00000f40 )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk0000049e/blk000004c7  (
    .I0(sig00000695),
    .O(\blk0000049e/sig00000f3f )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk0000049e/blk000004c6  (
    .I0(sig00000696),
    .O(\blk0000049e/sig00000f3e )
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  \blk0000049e/blk000004c5  (
    .I0(sig00000685),
    .I1(sig0000066e),
    .O(\blk0000049e/sig00000f2b )
  );
  MUXCY   \blk0000049e/blk000004c4  (
    .CI(\blk0000049e/sig00000f2a ),
    .DI(sig00000685),
    .S(\blk0000049e/sig00000f2b ),
    .O(\blk0000049e/sig00000f3d )
  );
  MUXCY   \blk0000049e/blk000004c3  (
    .CI(\blk0000049e/sig00000f3d ),
    .DI(sig00000686),
    .S(\blk0000049e/sig00000f4e ),
    .O(\blk0000049e/sig00000f3c )
  );
  MUXCY   \blk0000049e/blk000004c2  (
    .CI(\blk0000049e/sig00000f3c ),
    .DI(sig00000687),
    .S(\blk0000049e/sig00000f4d ),
    .O(\blk0000049e/sig00000f3b )
  );
  MUXCY   \blk0000049e/blk000004c1  (
    .CI(\blk0000049e/sig00000f3b ),
    .DI(sig00000688),
    .S(\blk0000049e/sig00000f4c ),
    .O(\blk0000049e/sig00000f3a )
  );
  MUXCY   \blk0000049e/blk000004c0  (
    .CI(\blk0000049e/sig00000f3a ),
    .DI(sig00000689),
    .S(\blk0000049e/sig00000f4b ),
    .O(\blk0000049e/sig00000f39 )
  );
  MUXCY   \blk0000049e/blk000004bf  (
    .CI(\blk0000049e/sig00000f39 ),
    .DI(sig0000068a),
    .S(\blk0000049e/sig00000f4a ),
    .O(\blk0000049e/sig00000f38 )
  );
  MUXCY   \blk0000049e/blk000004be  (
    .CI(\blk0000049e/sig00000f38 ),
    .DI(sig0000068b),
    .S(\blk0000049e/sig00000f49 ),
    .O(\blk0000049e/sig00000f37 )
  );
  MUXCY   \blk0000049e/blk000004bd  (
    .CI(\blk0000049e/sig00000f37 ),
    .DI(sig0000068c),
    .S(\blk0000049e/sig00000f48 ),
    .O(\blk0000049e/sig00000f36 )
  );
  MUXCY   \blk0000049e/blk000004bc  (
    .CI(\blk0000049e/sig00000f36 ),
    .DI(sig0000068d),
    .S(\blk0000049e/sig00000f47 ),
    .O(\blk0000049e/sig00000f35 )
  );
  MUXCY   \blk0000049e/blk000004bb  (
    .CI(\blk0000049e/sig00000f35 ),
    .DI(sig0000068e),
    .S(\blk0000049e/sig00000f46 ),
    .O(\blk0000049e/sig00000f34 )
  );
  MUXCY   \blk0000049e/blk000004ba  (
    .CI(\blk0000049e/sig00000f34 ),
    .DI(sig0000068f),
    .S(\blk0000049e/sig00000f45 ),
    .O(\blk0000049e/sig00000f33 )
  );
  MUXCY   \blk0000049e/blk000004b9  (
    .CI(\blk0000049e/sig00000f33 ),
    .DI(sig00000690),
    .S(\blk0000049e/sig00000f44 ),
    .O(\blk0000049e/sig00000f32 )
  );
  MUXCY   \blk0000049e/blk000004b8  (
    .CI(\blk0000049e/sig00000f32 ),
    .DI(sig00000691),
    .S(\blk0000049e/sig00000f43 ),
    .O(\blk0000049e/sig00000f31 )
  );
  MUXCY   \blk0000049e/blk000004b7  (
    .CI(\blk0000049e/sig00000f31 ),
    .DI(sig00000692),
    .S(\blk0000049e/sig00000f42 ),
    .O(\blk0000049e/sig00000f30 )
  );
  MUXCY   \blk0000049e/blk000004b6  (
    .CI(\blk0000049e/sig00000f30 ),
    .DI(sig00000693),
    .S(\blk0000049e/sig00000f41 ),
    .O(\blk0000049e/sig00000f2f )
  );
  MUXCY   \blk0000049e/blk000004b5  (
    .CI(\blk0000049e/sig00000f2f ),
    .DI(sig00000694),
    .S(\blk0000049e/sig00000f40 ),
    .O(\blk0000049e/sig00000f2e )
  );
  MUXCY   \blk0000049e/blk000004b4  (
    .CI(\blk0000049e/sig00000f2e ),
    .DI(sig00000695),
    .S(\blk0000049e/sig00000f3f ),
    .O(\blk0000049e/sig00000f2d )
  );
  MUXCY   \blk0000049e/blk000004b3  (
    .CI(\blk0000049e/sig00000f2d ),
    .DI(sig00000696),
    .S(\blk0000049e/sig00000f3e ),
    .O(\blk0000049e/sig00000f2c )
  );
  XORCY   \blk0000049e/blk000004b2  (
    .CI(\blk0000049e/sig00000f3d ),
    .LI(\blk0000049e/sig00000f4e ),
    .O(sig00000673)
  );
  XORCY   \blk0000049e/blk000004b1  (
    .CI(\blk0000049e/sig00000f3c ),
    .LI(\blk0000049e/sig00000f4d ),
    .O(sig00000674)
  );
  XORCY   \blk0000049e/blk000004b0  (
    .CI(\blk0000049e/sig00000f3b ),
    .LI(\blk0000049e/sig00000f4c ),
    .O(sig00000675)
  );
  XORCY   \blk0000049e/blk000004af  (
    .CI(\blk0000049e/sig00000f3a ),
    .LI(\blk0000049e/sig00000f4b ),
    .O(sig00000676)
  );
  XORCY   \blk0000049e/blk000004ae  (
    .CI(\blk0000049e/sig00000f39 ),
    .LI(\blk0000049e/sig00000f4a ),
    .O(sig00000677)
  );
  XORCY   \blk0000049e/blk000004ad  (
    .CI(\blk0000049e/sig00000f38 ),
    .LI(\blk0000049e/sig00000f49 ),
    .O(sig00000678)
  );
  XORCY   \blk0000049e/blk000004ac  (
    .CI(\blk0000049e/sig00000f37 ),
    .LI(\blk0000049e/sig00000f48 ),
    .O(sig00000679)
  );
  XORCY   \blk0000049e/blk000004ab  (
    .CI(\blk0000049e/sig00000f36 ),
    .LI(\blk0000049e/sig00000f47 ),
    .O(sig0000067a)
  );
  XORCY   \blk0000049e/blk000004aa  (
    .CI(\blk0000049e/sig00000f35 ),
    .LI(\blk0000049e/sig00000f46 ),
    .O(sig0000067b)
  );
  XORCY   \blk0000049e/blk000004a9  (
    .CI(\blk0000049e/sig00000f34 ),
    .LI(\blk0000049e/sig00000f45 ),
    .O(sig0000067c)
  );
  XORCY   \blk0000049e/blk000004a8  (
    .CI(\blk0000049e/sig00000f33 ),
    .LI(\blk0000049e/sig00000f44 ),
    .O(sig0000067d)
  );
  XORCY   \blk0000049e/blk000004a7  (
    .CI(\blk0000049e/sig00000f32 ),
    .LI(\blk0000049e/sig00000f43 ),
    .O(sig0000067e)
  );
  XORCY   \blk0000049e/blk000004a6  (
    .CI(\blk0000049e/sig00000f31 ),
    .LI(\blk0000049e/sig00000f42 ),
    .O(sig0000067f)
  );
  XORCY   \blk0000049e/blk000004a5  (
    .CI(\blk0000049e/sig00000f30 ),
    .LI(\blk0000049e/sig00000f41 ),
    .O(sig00000680)
  );
  XORCY   \blk0000049e/blk000004a4  (
    .CI(\blk0000049e/sig00000f2f ),
    .LI(\blk0000049e/sig00000f40 ),
    .O(sig00000681)
  );
  XORCY   \blk0000049e/blk000004a3  (
    .CI(\blk0000049e/sig00000f2e ),
    .LI(\blk0000049e/sig00000f3f ),
    .O(sig00000682)
  );
  XORCY   \blk0000049e/blk000004a2  (
    .CI(\blk0000049e/sig00000f2d ),
    .LI(\blk0000049e/sig00000f3e ),
    .O(sig00000683)
  );
  XORCY   \blk0000049e/blk000004a1  (
    .CI(\blk0000049e/sig00000f2c ),
    .LI(sig00000697),
    .O(sig00000684)
  );
  XORCY   \blk0000049e/blk000004a0  (
    .CI(\blk0000049e/sig00000f2a ),
    .LI(\blk0000049e/sig00000f2b ),
    .O(sig00000672)
  );
  GND   \blk0000049e/blk0000049f  (
    .G(\blk0000049e/sig00000f2a )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk000004d7/blk0000050f  (
    .I0(sig00000658),
    .O(\blk000004d7/sig00000f9a )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk000004d7/blk0000050e  (
    .I0(sig00000659),
    .O(\blk000004d7/sig00000f99 )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk000004d7/blk0000050d  (
    .I0(sig0000065a),
    .O(\blk000004d7/sig00000f98 )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk000004d7/blk0000050c  (
    .I0(sig0000065b),
    .O(\blk000004d7/sig00000f97 )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk000004d7/blk0000050b  (
    .I0(sig0000065c),
    .O(\blk000004d7/sig00000f96 )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk000004d7/blk0000050a  (
    .I0(sig0000065d),
    .O(\blk000004d7/sig00000f95 )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk000004d7/blk00000509  (
    .I0(sig0000065e),
    .O(\blk000004d7/sig00000f94 )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk000004d7/blk00000508  (
    .I0(sig0000065f),
    .O(\blk000004d7/sig00000f93 )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk000004d7/blk00000507  (
    .I0(sig00000660),
    .O(\blk000004d7/sig00000f92 )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk000004d7/blk00000506  (
    .I0(sig00000661),
    .O(\blk000004d7/sig00000f91 )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk000004d7/blk00000505  (
    .I0(sig00000662),
    .O(\blk000004d7/sig00000f90 )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk000004d7/blk00000504  (
    .I0(sig00000663),
    .O(\blk000004d7/sig00000f8f )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk000004d7/blk00000503  (
    .I0(sig00000664),
    .O(\blk000004d7/sig00000f8e )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk000004d7/blk00000502  (
    .I0(sig00000665),
    .O(\blk000004d7/sig00000f8d )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk000004d7/blk00000501  (
    .I0(sig00000666),
    .O(\blk000004d7/sig00000f8c )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk000004d7/blk00000500  (
    .I0(sig00000667),
    .O(\blk000004d7/sig00000f8b )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk000004d7/blk000004ff  (
    .I0(sig00000668),
    .O(\blk000004d7/sig00000f8a )
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  \blk000004d7/blk000004fe  (
    .I0(sig00000657),
    .I1(sig00000640),
    .O(\blk000004d7/sig00000f77 )
  );
  MUXCY   \blk000004d7/blk000004fd  (
    .CI(\blk000004d7/sig00000f76 ),
    .DI(sig00000657),
    .S(\blk000004d7/sig00000f77 ),
    .O(\blk000004d7/sig00000f89 )
  );
  MUXCY   \blk000004d7/blk000004fc  (
    .CI(\blk000004d7/sig00000f89 ),
    .DI(sig00000658),
    .S(\blk000004d7/sig00000f9a ),
    .O(\blk000004d7/sig00000f88 )
  );
  MUXCY   \blk000004d7/blk000004fb  (
    .CI(\blk000004d7/sig00000f88 ),
    .DI(sig00000659),
    .S(\blk000004d7/sig00000f99 ),
    .O(\blk000004d7/sig00000f87 )
  );
  MUXCY   \blk000004d7/blk000004fa  (
    .CI(\blk000004d7/sig00000f87 ),
    .DI(sig0000065a),
    .S(\blk000004d7/sig00000f98 ),
    .O(\blk000004d7/sig00000f86 )
  );
  MUXCY   \blk000004d7/blk000004f9  (
    .CI(\blk000004d7/sig00000f86 ),
    .DI(sig0000065b),
    .S(\blk000004d7/sig00000f97 ),
    .O(\blk000004d7/sig00000f85 )
  );
  MUXCY   \blk000004d7/blk000004f8  (
    .CI(\blk000004d7/sig00000f85 ),
    .DI(sig0000065c),
    .S(\blk000004d7/sig00000f96 ),
    .O(\blk000004d7/sig00000f84 )
  );
  MUXCY   \blk000004d7/blk000004f7  (
    .CI(\blk000004d7/sig00000f84 ),
    .DI(sig0000065d),
    .S(\blk000004d7/sig00000f95 ),
    .O(\blk000004d7/sig00000f83 )
  );
  MUXCY   \blk000004d7/blk000004f6  (
    .CI(\blk000004d7/sig00000f83 ),
    .DI(sig0000065e),
    .S(\blk000004d7/sig00000f94 ),
    .O(\blk000004d7/sig00000f82 )
  );
  MUXCY   \blk000004d7/blk000004f5  (
    .CI(\blk000004d7/sig00000f82 ),
    .DI(sig0000065f),
    .S(\blk000004d7/sig00000f93 ),
    .O(\blk000004d7/sig00000f81 )
  );
  MUXCY   \blk000004d7/blk000004f4  (
    .CI(\blk000004d7/sig00000f81 ),
    .DI(sig00000660),
    .S(\blk000004d7/sig00000f92 ),
    .O(\blk000004d7/sig00000f80 )
  );
  MUXCY   \blk000004d7/blk000004f3  (
    .CI(\blk000004d7/sig00000f80 ),
    .DI(sig00000661),
    .S(\blk000004d7/sig00000f91 ),
    .O(\blk000004d7/sig00000f7f )
  );
  MUXCY   \blk000004d7/blk000004f2  (
    .CI(\blk000004d7/sig00000f7f ),
    .DI(sig00000662),
    .S(\blk000004d7/sig00000f90 ),
    .O(\blk000004d7/sig00000f7e )
  );
  MUXCY   \blk000004d7/blk000004f1  (
    .CI(\blk000004d7/sig00000f7e ),
    .DI(sig00000663),
    .S(\blk000004d7/sig00000f8f ),
    .O(\blk000004d7/sig00000f7d )
  );
  MUXCY   \blk000004d7/blk000004f0  (
    .CI(\blk000004d7/sig00000f7d ),
    .DI(sig00000664),
    .S(\blk000004d7/sig00000f8e ),
    .O(\blk000004d7/sig00000f7c )
  );
  MUXCY   \blk000004d7/blk000004ef  (
    .CI(\blk000004d7/sig00000f7c ),
    .DI(sig00000665),
    .S(\blk000004d7/sig00000f8d ),
    .O(\blk000004d7/sig00000f7b )
  );
  MUXCY   \blk000004d7/blk000004ee  (
    .CI(\blk000004d7/sig00000f7b ),
    .DI(sig00000666),
    .S(\blk000004d7/sig00000f8c ),
    .O(\blk000004d7/sig00000f7a )
  );
  MUXCY   \blk000004d7/blk000004ed  (
    .CI(\blk000004d7/sig00000f7a ),
    .DI(sig00000667),
    .S(\blk000004d7/sig00000f8b ),
    .O(\blk000004d7/sig00000f79 )
  );
  MUXCY   \blk000004d7/blk000004ec  (
    .CI(\blk000004d7/sig00000f79 ),
    .DI(sig00000668),
    .S(\blk000004d7/sig00000f8a ),
    .O(\blk000004d7/sig00000f78 )
  );
  XORCY   \blk000004d7/blk000004eb  (
    .CI(\blk000004d7/sig00000f89 ),
    .LI(\blk000004d7/sig00000f9a ),
    .O(sig00000645)
  );
  XORCY   \blk000004d7/blk000004ea  (
    .CI(\blk000004d7/sig00000f88 ),
    .LI(\blk000004d7/sig00000f99 ),
    .O(sig00000646)
  );
  XORCY   \blk000004d7/blk000004e9  (
    .CI(\blk000004d7/sig00000f87 ),
    .LI(\blk000004d7/sig00000f98 ),
    .O(sig00000647)
  );
  XORCY   \blk000004d7/blk000004e8  (
    .CI(\blk000004d7/sig00000f86 ),
    .LI(\blk000004d7/sig00000f97 ),
    .O(sig00000648)
  );
  XORCY   \blk000004d7/blk000004e7  (
    .CI(\blk000004d7/sig00000f85 ),
    .LI(\blk000004d7/sig00000f96 ),
    .O(sig00000649)
  );
  XORCY   \blk000004d7/blk000004e6  (
    .CI(\blk000004d7/sig00000f84 ),
    .LI(\blk000004d7/sig00000f95 ),
    .O(sig0000064a)
  );
  XORCY   \blk000004d7/blk000004e5  (
    .CI(\blk000004d7/sig00000f83 ),
    .LI(\blk000004d7/sig00000f94 ),
    .O(sig0000064b)
  );
  XORCY   \blk000004d7/blk000004e4  (
    .CI(\blk000004d7/sig00000f82 ),
    .LI(\blk000004d7/sig00000f93 ),
    .O(sig0000064c)
  );
  XORCY   \blk000004d7/blk000004e3  (
    .CI(\blk000004d7/sig00000f81 ),
    .LI(\blk000004d7/sig00000f92 ),
    .O(sig0000064d)
  );
  XORCY   \blk000004d7/blk000004e2  (
    .CI(\blk000004d7/sig00000f80 ),
    .LI(\blk000004d7/sig00000f91 ),
    .O(sig0000064e)
  );
  XORCY   \blk000004d7/blk000004e1  (
    .CI(\blk000004d7/sig00000f7f ),
    .LI(\blk000004d7/sig00000f90 ),
    .O(sig0000064f)
  );
  XORCY   \blk000004d7/blk000004e0  (
    .CI(\blk000004d7/sig00000f7e ),
    .LI(\blk000004d7/sig00000f8f ),
    .O(sig00000650)
  );
  XORCY   \blk000004d7/blk000004df  (
    .CI(\blk000004d7/sig00000f7d ),
    .LI(\blk000004d7/sig00000f8e ),
    .O(sig00000651)
  );
  XORCY   \blk000004d7/blk000004de  (
    .CI(\blk000004d7/sig00000f7c ),
    .LI(\blk000004d7/sig00000f8d ),
    .O(sig00000652)
  );
  XORCY   \blk000004d7/blk000004dd  (
    .CI(\blk000004d7/sig00000f7b ),
    .LI(\blk000004d7/sig00000f8c ),
    .O(sig00000653)
  );
  XORCY   \blk000004d7/blk000004dc  (
    .CI(\blk000004d7/sig00000f7a ),
    .LI(\blk000004d7/sig00000f8b ),
    .O(sig00000654)
  );
  XORCY   \blk000004d7/blk000004db  (
    .CI(\blk000004d7/sig00000f79 ),
    .LI(\blk000004d7/sig00000f8a ),
    .O(sig00000655)
  );
  XORCY   \blk000004d7/blk000004da  (
    .CI(\blk000004d7/sig00000f78 ),
    .LI(sig00000669),
    .O(sig00000656)
  );
  XORCY   \blk000004d7/blk000004d9  (
    .CI(\blk000004d7/sig00000f76 ),
    .LI(\blk000004d7/sig00000f77 ),
    .O(sig00000644)
  );
  GND   \blk000004d7/blk000004d8  (
    .G(\blk000004d7/sig00000f76 )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk00000510/blk00000548  (
    .I0(sig0000062a),
    .O(\blk00000510/sig00000fe6 )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk00000510/blk00000547  (
    .I0(sig0000062b),
    .O(\blk00000510/sig00000fe5 )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk00000510/blk00000546  (
    .I0(sig0000062c),
    .O(\blk00000510/sig00000fe4 )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk00000510/blk00000545  (
    .I0(sig0000062d),
    .O(\blk00000510/sig00000fe3 )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk00000510/blk00000544  (
    .I0(sig0000062e),
    .O(\blk00000510/sig00000fe2 )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk00000510/blk00000543  (
    .I0(sig0000062f),
    .O(\blk00000510/sig00000fe1 )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk00000510/blk00000542  (
    .I0(sig00000630),
    .O(\blk00000510/sig00000fe0 )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk00000510/blk00000541  (
    .I0(sig00000631),
    .O(\blk00000510/sig00000fdf )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk00000510/blk00000540  (
    .I0(sig00000632),
    .O(\blk00000510/sig00000fde )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk00000510/blk0000053f  (
    .I0(sig00000633),
    .O(\blk00000510/sig00000fdd )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk00000510/blk0000053e  (
    .I0(sig00000634),
    .O(\blk00000510/sig00000fdc )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk00000510/blk0000053d  (
    .I0(sig00000635),
    .O(\blk00000510/sig00000fdb )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk00000510/blk0000053c  (
    .I0(sig00000636),
    .O(\blk00000510/sig00000fda )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk00000510/blk0000053b  (
    .I0(sig00000637),
    .O(\blk00000510/sig00000fd9 )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk00000510/blk0000053a  (
    .I0(sig00000638),
    .O(\blk00000510/sig00000fd8 )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk00000510/blk00000539  (
    .I0(sig00000639),
    .O(\blk00000510/sig00000fd7 )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk00000510/blk00000538  (
    .I0(sig0000063a),
    .O(\blk00000510/sig00000fd6 )
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  \blk00000510/blk00000537  (
    .I0(sig00000629),
    .I1(sig00000612),
    .O(\blk00000510/sig00000fc3 )
  );
  MUXCY   \blk00000510/blk00000536  (
    .CI(\blk00000510/sig00000fc2 ),
    .DI(sig00000629),
    .S(\blk00000510/sig00000fc3 ),
    .O(\blk00000510/sig00000fd5 )
  );
  MUXCY   \blk00000510/blk00000535  (
    .CI(\blk00000510/sig00000fd5 ),
    .DI(sig0000062a),
    .S(\blk00000510/sig00000fe6 ),
    .O(\blk00000510/sig00000fd4 )
  );
  MUXCY   \blk00000510/blk00000534  (
    .CI(\blk00000510/sig00000fd4 ),
    .DI(sig0000062b),
    .S(\blk00000510/sig00000fe5 ),
    .O(\blk00000510/sig00000fd3 )
  );
  MUXCY   \blk00000510/blk00000533  (
    .CI(\blk00000510/sig00000fd3 ),
    .DI(sig0000062c),
    .S(\blk00000510/sig00000fe4 ),
    .O(\blk00000510/sig00000fd2 )
  );
  MUXCY   \blk00000510/blk00000532  (
    .CI(\blk00000510/sig00000fd2 ),
    .DI(sig0000062d),
    .S(\blk00000510/sig00000fe3 ),
    .O(\blk00000510/sig00000fd1 )
  );
  MUXCY   \blk00000510/blk00000531  (
    .CI(\blk00000510/sig00000fd1 ),
    .DI(sig0000062e),
    .S(\blk00000510/sig00000fe2 ),
    .O(\blk00000510/sig00000fd0 )
  );
  MUXCY   \blk00000510/blk00000530  (
    .CI(\blk00000510/sig00000fd0 ),
    .DI(sig0000062f),
    .S(\blk00000510/sig00000fe1 ),
    .O(\blk00000510/sig00000fcf )
  );
  MUXCY   \blk00000510/blk0000052f  (
    .CI(\blk00000510/sig00000fcf ),
    .DI(sig00000630),
    .S(\blk00000510/sig00000fe0 ),
    .O(\blk00000510/sig00000fce )
  );
  MUXCY   \blk00000510/blk0000052e  (
    .CI(\blk00000510/sig00000fce ),
    .DI(sig00000631),
    .S(\blk00000510/sig00000fdf ),
    .O(\blk00000510/sig00000fcd )
  );
  MUXCY   \blk00000510/blk0000052d  (
    .CI(\blk00000510/sig00000fcd ),
    .DI(sig00000632),
    .S(\blk00000510/sig00000fde ),
    .O(\blk00000510/sig00000fcc )
  );
  MUXCY   \blk00000510/blk0000052c  (
    .CI(\blk00000510/sig00000fcc ),
    .DI(sig00000633),
    .S(\blk00000510/sig00000fdd ),
    .O(\blk00000510/sig00000fcb )
  );
  MUXCY   \blk00000510/blk0000052b  (
    .CI(\blk00000510/sig00000fcb ),
    .DI(sig00000634),
    .S(\blk00000510/sig00000fdc ),
    .O(\blk00000510/sig00000fca )
  );
  MUXCY   \blk00000510/blk0000052a  (
    .CI(\blk00000510/sig00000fca ),
    .DI(sig00000635),
    .S(\blk00000510/sig00000fdb ),
    .O(\blk00000510/sig00000fc9 )
  );
  MUXCY   \blk00000510/blk00000529  (
    .CI(\blk00000510/sig00000fc9 ),
    .DI(sig00000636),
    .S(\blk00000510/sig00000fda ),
    .O(\blk00000510/sig00000fc8 )
  );
  MUXCY   \blk00000510/blk00000528  (
    .CI(\blk00000510/sig00000fc8 ),
    .DI(sig00000637),
    .S(\blk00000510/sig00000fd9 ),
    .O(\blk00000510/sig00000fc7 )
  );
  MUXCY   \blk00000510/blk00000527  (
    .CI(\blk00000510/sig00000fc7 ),
    .DI(sig00000638),
    .S(\blk00000510/sig00000fd8 ),
    .O(\blk00000510/sig00000fc6 )
  );
  MUXCY   \blk00000510/blk00000526  (
    .CI(\blk00000510/sig00000fc6 ),
    .DI(sig00000639),
    .S(\blk00000510/sig00000fd7 ),
    .O(\blk00000510/sig00000fc5 )
  );
  MUXCY   \blk00000510/blk00000525  (
    .CI(\blk00000510/sig00000fc5 ),
    .DI(sig0000063a),
    .S(\blk00000510/sig00000fd6 ),
    .O(\blk00000510/sig00000fc4 )
  );
  XORCY   \blk00000510/blk00000524  (
    .CI(\blk00000510/sig00000fd5 ),
    .LI(\blk00000510/sig00000fe6 ),
    .O(sig00000617)
  );
  XORCY   \blk00000510/blk00000523  (
    .CI(\blk00000510/sig00000fd4 ),
    .LI(\blk00000510/sig00000fe5 ),
    .O(sig00000618)
  );
  XORCY   \blk00000510/blk00000522  (
    .CI(\blk00000510/sig00000fd3 ),
    .LI(\blk00000510/sig00000fe4 ),
    .O(sig00000619)
  );
  XORCY   \blk00000510/blk00000521  (
    .CI(\blk00000510/sig00000fd2 ),
    .LI(\blk00000510/sig00000fe3 ),
    .O(sig0000061a)
  );
  XORCY   \blk00000510/blk00000520  (
    .CI(\blk00000510/sig00000fd1 ),
    .LI(\blk00000510/sig00000fe2 ),
    .O(sig0000061b)
  );
  XORCY   \blk00000510/blk0000051f  (
    .CI(\blk00000510/sig00000fd0 ),
    .LI(\blk00000510/sig00000fe1 ),
    .O(sig0000061c)
  );
  XORCY   \blk00000510/blk0000051e  (
    .CI(\blk00000510/sig00000fcf ),
    .LI(\blk00000510/sig00000fe0 ),
    .O(sig0000061d)
  );
  XORCY   \blk00000510/blk0000051d  (
    .CI(\blk00000510/sig00000fce ),
    .LI(\blk00000510/sig00000fdf ),
    .O(sig0000061e)
  );
  XORCY   \blk00000510/blk0000051c  (
    .CI(\blk00000510/sig00000fcd ),
    .LI(\blk00000510/sig00000fde ),
    .O(sig0000061f)
  );
  XORCY   \blk00000510/blk0000051b  (
    .CI(\blk00000510/sig00000fcc ),
    .LI(\blk00000510/sig00000fdd ),
    .O(sig00000620)
  );
  XORCY   \blk00000510/blk0000051a  (
    .CI(\blk00000510/sig00000fcb ),
    .LI(\blk00000510/sig00000fdc ),
    .O(sig00000621)
  );
  XORCY   \blk00000510/blk00000519  (
    .CI(\blk00000510/sig00000fca ),
    .LI(\blk00000510/sig00000fdb ),
    .O(sig00000622)
  );
  XORCY   \blk00000510/blk00000518  (
    .CI(\blk00000510/sig00000fc9 ),
    .LI(\blk00000510/sig00000fda ),
    .O(sig00000623)
  );
  XORCY   \blk00000510/blk00000517  (
    .CI(\blk00000510/sig00000fc8 ),
    .LI(\blk00000510/sig00000fd9 ),
    .O(sig00000624)
  );
  XORCY   \blk00000510/blk00000516  (
    .CI(\blk00000510/sig00000fc7 ),
    .LI(\blk00000510/sig00000fd8 ),
    .O(sig00000625)
  );
  XORCY   \blk00000510/blk00000515  (
    .CI(\blk00000510/sig00000fc6 ),
    .LI(\blk00000510/sig00000fd7 ),
    .O(sig00000626)
  );
  XORCY   \blk00000510/blk00000514  (
    .CI(\blk00000510/sig00000fc5 ),
    .LI(\blk00000510/sig00000fd6 ),
    .O(sig00000627)
  );
  XORCY   \blk00000510/blk00000513  (
    .CI(\blk00000510/sig00000fc4 ),
    .LI(sig0000063b),
    .O(sig00000628)
  );
  XORCY   \blk00000510/blk00000512  (
    .CI(\blk00000510/sig00000fc2 ),
    .LI(\blk00000510/sig00000fc3 ),
    .O(sig00000616)
  );
  GND   \blk00000510/blk00000511  (
    .G(\blk00000510/sig00000fc2 )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk00000549/blk00000581  (
    .I0(sig000005fc),
    .O(\blk00000549/sig00001032 )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk00000549/blk00000580  (
    .I0(sig000005fd),
    .O(\blk00000549/sig00001031 )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk00000549/blk0000057f  (
    .I0(sig000005fe),
    .O(\blk00000549/sig00001030 )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk00000549/blk0000057e  (
    .I0(sig000005ff),
    .O(\blk00000549/sig0000102f )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk00000549/blk0000057d  (
    .I0(sig00000600),
    .O(\blk00000549/sig0000102e )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk00000549/blk0000057c  (
    .I0(sig00000601),
    .O(\blk00000549/sig0000102d )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk00000549/blk0000057b  (
    .I0(sig00000602),
    .O(\blk00000549/sig0000102c )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk00000549/blk0000057a  (
    .I0(sig00000603),
    .O(\blk00000549/sig0000102b )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk00000549/blk00000579  (
    .I0(sig00000604),
    .O(\blk00000549/sig0000102a )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk00000549/blk00000578  (
    .I0(sig00000605),
    .O(\blk00000549/sig00001029 )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk00000549/blk00000577  (
    .I0(sig00000606),
    .O(\blk00000549/sig00001028 )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk00000549/blk00000576  (
    .I0(sig00000607),
    .O(\blk00000549/sig00001027 )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk00000549/blk00000575  (
    .I0(sig00000608),
    .O(\blk00000549/sig00001026 )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk00000549/blk00000574  (
    .I0(sig00000609),
    .O(\blk00000549/sig00001025 )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk00000549/blk00000573  (
    .I0(sig0000060a),
    .O(\blk00000549/sig00001024 )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk00000549/blk00000572  (
    .I0(sig0000060b),
    .O(\blk00000549/sig00001023 )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk00000549/blk00000571  (
    .I0(sig0000060c),
    .O(\blk00000549/sig00001022 )
  );
  LUT2 #(
    .INIT ( 4'h6 ))
  \blk00000549/blk00000570  (
    .I0(sig000005fb),
    .I1(sig000005e4),
    .O(\blk00000549/sig0000100f )
  );
  MUXCY   \blk00000549/blk0000056f  (
    .CI(\blk00000549/sig0000100e ),
    .DI(sig000005fb),
    .S(\blk00000549/sig0000100f ),
    .O(\blk00000549/sig00001021 )
  );
  MUXCY   \blk00000549/blk0000056e  (
    .CI(\blk00000549/sig00001021 ),
    .DI(sig000005fc),
    .S(\blk00000549/sig00001032 ),
    .O(\blk00000549/sig00001020 )
  );
  MUXCY   \blk00000549/blk0000056d  (
    .CI(\blk00000549/sig00001020 ),
    .DI(sig000005fd),
    .S(\blk00000549/sig00001031 ),
    .O(\blk00000549/sig0000101f )
  );
  MUXCY   \blk00000549/blk0000056c  (
    .CI(\blk00000549/sig0000101f ),
    .DI(sig000005fe),
    .S(\blk00000549/sig00001030 ),
    .O(\blk00000549/sig0000101e )
  );
  MUXCY   \blk00000549/blk0000056b  (
    .CI(\blk00000549/sig0000101e ),
    .DI(sig000005ff),
    .S(\blk00000549/sig0000102f ),
    .O(\blk00000549/sig0000101d )
  );
  MUXCY   \blk00000549/blk0000056a  (
    .CI(\blk00000549/sig0000101d ),
    .DI(sig00000600),
    .S(\blk00000549/sig0000102e ),
    .O(\blk00000549/sig0000101c )
  );
  MUXCY   \blk00000549/blk00000569  (
    .CI(\blk00000549/sig0000101c ),
    .DI(sig00000601),
    .S(\blk00000549/sig0000102d ),
    .O(\blk00000549/sig0000101b )
  );
  MUXCY   \blk00000549/blk00000568  (
    .CI(\blk00000549/sig0000101b ),
    .DI(sig00000602),
    .S(\blk00000549/sig0000102c ),
    .O(\blk00000549/sig0000101a )
  );
  MUXCY   \blk00000549/blk00000567  (
    .CI(\blk00000549/sig0000101a ),
    .DI(sig00000603),
    .S(\blk00000549/sig0000102b ),
    .O(\blk00000549/sig00001019 )
  );
  MUXCY   \blk00000549/blk00000566  (
    .CI(\blk00000549/sig00001019 ),
    .DI(sig00000604),
    .S(\blk00000549/sig0000102a ),
    .O(\blk00000549/sig00001018 )
  );
  MUXCY   \blk00000549/blk00000565  (
    .CI(\blk00000549/sig00001018 ),
    .DI(sig00000605),
    .S(\blk00000549/sig00001029 ),
    .O(\blk00000549/sig00001017 )
  );
  MUXCY   \blk00000549/blk00000564  (
    .CI(\blk00000549/sig00001017 ),
    .DI(sig00000606),
    .S(\blk00000549/sig00001028 ),
    .O(\blk00000549/sig00001016 )
  );
  MUXCY   \blk00000549/blk00000563  (
    .CI(\blk00000549/sig00001016 ),
    .DI(sig00000607),
    .S(\blk00000549/sig00001027 ),
    .O(\blk00000549/sig00001015 )
  );
  MUXCY   \blk00000549/blk00000562  (
    .CI(\blk00000549/sig00001015 ),
    .DI(sig00000608),
    .S(\blk00000549/sig00001026 ),
    .O(\blk00000549/sig00001014 )
  );
  MUXCY   \blk00000549/blk00000561  (
    .CI(\blk00000549/sig00001014 ),
    .DI(sig00000609),
    .S(\blk00000549/sig00001025 ),
    .O(\blk00000549/sig00001013 )
  );
  MUXCY   \blk00000549/blk00000560  (
    .CI(\blk00000549/sig00001013 ),
    .DI(sig0000060a),
    .S(\blk00000549/sig00001024 ),
    .O(\blk00000549/sig00001012 )
  );
  MUXCY   \blk00000549/blk0000055f  (
    .CI(\blk00000549/sig00001012 ),
    .DI(sig0000060b),
    .S(\blk00000549/sig00001023 ),
    .O(\blk00000549/sig00001011 )
  );
  MUXCY   \blk00000549/blk0000055e  (
    .CI(\blk00000549/sig00001011 ),
    .DI(sig0000060c),
    .S(\blk00000549/sig00001022 ),
    .O(\blk00000549/sig00001010 )
  );
  XORCY   \blk00000549/blk0000055d  (
    .CI(\blk00000549/sig00001021 ),
    .LI(\blk00000549/sig00001032 ),
    .O(sig000005e9)
  );
  XORCY   \blk00000549/blk0000055c  (
    .CI(\blk00000549/sig00001020 ),
    .LI(\blk00000549/sig00001031 ),
    .O(sig000005ea)
  );
  XORCY   \blk00000549/blk0000055b  (
    .CI(\blk00000549/sig0000101f ),
    .LI(\blk00000549/sig00001030 ),
    .O(sig000005eb)
  );
  XORCY   \blk00000549/blk0000055a  (
    .CI(\blk00000549/sig0000101e ),
    .LI(\blk00000549/sig0000102f ),
    .O(sig000005ec)
  );
  XORCY   \blk00000549/blk00000559  (
    .CI(\blk00000549/sig0000101d ),
    .LI(\blk00000549/sig0000102e ),
    .O(sig000005ed)
  );
  XORCY   \blk00000549/blk00000558  (
    .CI(\blk00000549/sig0000101c ),
    .LI(\blk00000549/sig0000102d ),
    .O(sig000005ee)
  );
  XORCY   \blk00000549/blk00000557  (
    .CI(\blk00000549/sig0000101b ),
    .LI(\blk00000549/sig0000102c ),
    .O(sig000005ef)
  );
  XORCY   \blk00000549/blk00000556  (
    .CI(\blk00000549/sig0000101a ),
    .LI(\blk00000549/sig0000102b ),
    .O(sig000005f0)
  );
  XORCY   \blk00000549/blk00000555  (
    .CI(\blk00000549/sig00001019 ),
    .LI(\blk00000549/sig0000102a ),
    .O(sig000005f1)
  );
  XORCY   \blk00000549/blk00000554  (
    .CI(\blk00000549/sig00001018 ),
    .LI(\blk00000549/sig00001029 ),
    .O(sig000005f2)
  );
  XORCY   \blk00000549/blk00000553  (
    .CI(\blk00000549/sig00001017 ),
    .LI(\blk00000549/sig00001028 ),
    .O(sig000005f3)
  );
  XORCY   \blk00000549/blk00000552  (
    .CI(\blk00000549/sig00001016 ),
    .LI(\blk00000549/sig00001027 ),
    .O(sig000005f4)
  );
  XORCY   \blk00000549/blk00000551  (
    .CI(\blk00000549/sig00001015 ),
    .LI(\blk00000549/sig00001026 ),
    .O(sig000005f5)
  );
  XORCY   \blk00000549/blk00000550  (
    .CI(\blk00000549/sig00001014 ),
    .LI(\blk00000549/sig00001025 ),
    .O(sig000005f6)
  );
  XORCY   \blk00000549/blk0000054f  (
    .CI(\blk00000549/sig00001013 ),
    .LI(\blk00000549/sig00001024 ),
    .O(sig000005f7)
  );
  XORCY   \blk00000549/blk0000054e  (
    .CI(\blk00000549/sig00001012 ),
    .LI(\blk00000549/sig00001023 ),
    .O(sig000005f8)
  );
  XORCY   \blk00000549/blk0000054d  (
    .CI(\blk00000549/sig00001011 ),
    .LI(\blk00000549/sig00001022 ),
    .O(sig000005f9)
  );
  XORCY   \blk00000549/blk0000054c  (
    .CI(\blk00000549/sig00001010 ),
    .LI(sig0000060d),
    .O(sig000005fa)
  );
  XORCY   \blk00000549/blk0000054b  (
    .CI(\blk00000549/sig0000100e ),
    .LI(\blk00000549/sig0000100f ),
    .O(sig000005e8)
  );
  GND   \blk00000549/blk0000054a  (
    .G(\blk00000549/sig0000100e )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000751/blk00000752/blk00000756  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk00000751/blk00000752/sig0000103e ),
    .Q(sig0000000b)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000751/blk00000752/blk00000755  (
    .A0(\blk00000751/blk00000752/sig0000103d ),
    .A1(\blk00000751/blk00000752/sig0000103c ),
    .A2(\blk00000751/blk00000752/sig0000103c ),
    .A3(\blk00000751/blk00000752/sig0000103c ),
    .CE(sig00000001),
    .CLK(clk),
    .D(\NlwRenamedSig_OI_U0/i_synth/non_floating_point.arch_c.xfft_inst/control/cntrl/loading_state/ORS ),
    .Q(\blk00000751/blk00000752/sig0000103e ),
    .Q15(\NLW_blk00000751/blk00000752/blk00000755_Q15_UNCONNECTED )
  );
  VCC   \blk00000751/blk00000752/blk00000754  (
    .P(\blk00000751/blk00000752/sig0000103d )
  );
  GND   \blk00000751/blk00000752/blk00000753  (
    .G(\blk00000751/blk00000752/sig0000103c )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000757/blk00000758/blk0000075c  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk00000757/blk00000758/sig0000104a ),
    .Q(sig00000006)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000757/blk00000758/blk0000075b  (
    .A0(\blk00000757/blk00000758/sig00001049 ),
    .A1(\blk00000757/blk00000758/sig00001048 ),
    .A2(\blk00000757/blk00000758/sig00001048 ),
    .A3(\blk00000757/blk00000758/sig00001048 ),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig000007f6),
    .Q(\blk00000757/blk00000758/sig0000104a ),
    .Q15(\NLW_blk00000757/blk00000758/blk0000075b_Q15_UNCONNECTED )
  );
  VCC   \blk00000757/blk00000758/blk0000075a  (
    .P(\blk00000757/blk00000758/sig00001049 )
  );
  GND   \blk00000757/blk00000758/blk00000759  (
    .G(\blk00000757/blk00000758/sig00001048 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000007ea/blk000007eb/blk000007fd  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk000007ea/blk000007eb/sig00001079 ),
    .Q(sig00000835)
  );
  SRLC32E #(
    .INIT ( 32'h00000000 ))
  \blk000007ea/blk000007eb/blk000007fc  (
    .CLK(clk),
    .D(sig00000847),
    .CE(sig00000001),
    .Q(\blk000007ea/blk000007eb/sig00001079 ),
    .Q31(\NLW_blk000007ea/blk000007eb/blk000007fc_Q31_UNCONNECTED ),
    .A({\blk000007ea/blk000007eb/sig00001071 , \blk000007ea/blk000007eb/sig00001070 , \blk000007ea/blk000007eb/sig00001070 ,
\blk000007ea/blk000007eb/sig00001071 , \blk000007ea/blk000007eb/sig00001071 })
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000007ea/blk000007eb/blk000007fb  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk000007ea/blk000007eb/sig00001078 ),
    .Q(sig00000834)
  );
  SRLC32E #(
    .INIT ( 32'h00000000 ))
  \blk000007ea/blk000007eb/blk000007fa  (
    .CLK(clk),
    .D(sig00000846),
    .CE(sig00000001),
    .Q(\blk000007ea/blk000007eb/sig00001078 ),
    .Q31(\NLW_blk000007ea/blk000007eb/blk000007fa_Q31_UNCONNECTED ),
    .A({\blk000007ea/blk000007eb/sig00001071 , \blk000007ea/blk000007eb/sig00001070 , \blk000007ea/blk000007eb/sig00001070 ,
\blk000007ea/blk000007eb/sig00001071 , \blk000007ea/blk000007eb/sig00001071 })
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000007ea/blk000007eb/blk000007f9  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk000007ea/blk000007eb/sig00001077 ),
    .Q(sig00000833)
  );
  SRLC32E #(
    .INIT ( 32'h00000000 ))
  \blk000007ea/blk000007eb/blk000007f8  (
    .CLK(clk),
    .D(sig00000845),
    .CE(sig00000001),
    .Q(\blk000007ea/blk000007eb/sig00001077 ),
    .Q31(\NLW_blk000007ea/blk000007eb/blk000007f8_Q31_UNCONNECTED ),
    .A({\blk000007ea/blk000007eb/sig00001071 , \blk000007ea/blk000007eb/sig00001070 , \blk000007ea/blk000007eb/sig00001070 ,
\blk000007ea/blk000007eb/sig00001071 , \blk000007ea/blk000007eb/sig00001071 })
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000007ea/blk000007eb/blk000007f7  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk000007ea/blk000007eb/sig00001076 ),
    .Q(sig00000832)
  );
  SRLC32E #(
    .INIT ( 32'h00000000 ))
  \blk000007ea/blk000007eb/blk000007f6  (
    .CLK(clk),
    .D(sig00000844),
    .CE(sig00000001),
    .Q(\blk000007ea/blk000007eb/sig00001076 ),
    .Q31(\NLW_blk000007ea/blk000007eb/blk000007f6_Q31_UNCONNECTED ),
    .A({\blk000007ea/blk000007eb/sig00001071 , \blk000007ea/blk000007eb/sig00001070 , \blk000007ea/blk000007eb/sig00001070 ,
\blk000007ea/blk000007eb/sig00001071 , \blk000007ea/blk000007eb/sig00001071 })
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000007ea/blk000007eb/blk000007f5  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk000007ea/blk000007eb/sig00001075 ),
    .Q(sig00000831)
  );
  SRLC32E #(
    .INIT ( 32'h00000000 ))
  \blk000007ea/blk000007eb/blk000007f4  (
    .CLK(clk),
    .D(sig00000843),
    .CE(sig00000001),
    .Q(\blk000007ea/blk000007eb/sig00001075 ),
    .Q31(\NLW_blk000007ea/blk000007eb/blk000007f4_Q31_UNCONNECTED ),
    .A({\blk000007ea/blk000007eb/sig00001071 , \blk000007ea/blk000007eb/sig00001070 , \blk000007ea/blk000007eb/sig00001070 ,
\blk000007ea/blk000007eb/sig00001071 , \blk000007ea/blk000007eb/sig00001071 })
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000007ea/blk000007eb/blk000007f3  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk000007ea/blk000007eb/sig00001074 ),
    .Q(sig00000830)
  );
  SRLC32E #(
    .INIT ( 32'h00000000 ))
  \blk000007ea/blk000007eb/blk000007f2  (
    .CLK(clk),
    .D(sig00000842),
    .CE(sig00000001),
    .Q(\blk000007ea/blk000007eb/sig00001074 ),
    .Q31(\NLW_blk000007ea/blk000007eb/blk000007f2_Q31_UNCONNECTED ),
    .A({\blk000007ea/blk000007eb/sig00001071 , \blk000007ea/blk000007eb/sig00001070 , \blk000007ea/blk000007eb/sig00001070 ,
\blk000007ea/blk000007eb/sig00001071 , \blk000007ea/blk000007eb/sig00001071 })
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000007ea/blk000007eb/blk000007f1  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk000007ea/blk000007eb/sig00001073 ),
    .Q(sig0000082f)
  );
  SRLC32E #(
    .INIT ( 32'h00000000 ))
  \blk000007ea/blk000007eb/blk000007f0  (
    .CLK(clk),
    .D(sig00000841),
    .CE(sig00000001),
    .Q(\blk000007ea/blk000007eb/sig00001073 ),
    .Q31(\NLW_blk000007ea/blk000007eb/blk000007f0_Q31_UNCONNECTED ),
    .A({\blk000007ea/blk000007eb/sig00001071 , \blk000007ea/blk000007eb/sig00001070 , \blk000007ea/blk000007eb/sig00001070 ,
\blk000007ea/blk000007eb/sig00001071 , \blk000007ea/blk000007eb/sig00001071 })
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000007ea/blk000007eb/blk000007ef  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk000007ea/blk000007eb/sig00001072 ),
    .Q(sig0000082e)
  );
  SRLC32E #(
    .INIT ( 32'h00000000 ))
  \blk000007ea/blk000007eb/blk000007ee  (
    .CLK(clk),
    .D(sig00000840),
    .CE(sig00000001),
    .Q(\blk000007ea/blk000007eb/sig00001072 ),
    .Q31(\NLW_blk000007ea/blk000007eb/blk000007ee_Q31_UNCONNECTED ),
    .A({\blk000007ea/blk000007eb/sig00001071 , \blk000007ea/blk000007eb/sig00001070 , \blk000007ea/blk000007eb/sig00001070 ,
\blk000007ea/blk000007eb/sig00001071 , \blk000007ea/blk000007eb/sig00001071 })
  );
  VCC   \blk000007ea/blk000007eb/blk000007ed  (
    .P(\blk000007ea/blk000007eb/sig00001071 )
  );
  GND   \blk000007ea/blk000007eb/blk000007ec  (
    .G(\blk000007ea/blk000007eb/sig00001070 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000007fe/blk000007ff/blk00000811  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk000007fe/blk000007ff/sig000010a8 ),
    .Q(sig0000082d)
  );
  SRLC32E #(
    .INIT ( 32'h00000000 ))
  \blk000007fe/blk000007ff/blk00000810  (
    .CLK(clk),
    .D(sig0000083f),
    .CE(sig00000001),
    .Q(\blk000007fe/blk000007ff/sig000010a8 ),
    .Q31(\NLW_blk000007fe/blk000007ff/blk00000810_Q31_UNCONNECTED ),
    .A({\blk000007fe/blk000007ff/sig000010a0 , \blk000007fe/blk000007ff/sig0000109f , \blk000007fe/blk000007ff/sig0000109f ,
\blk000007fe/blk000007ff/sig000010a0 , \blk000007fe/blk000007ff/sig000010a0 })
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000007fe/blk000007ff/blk0000080f  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk000007fe/blk000007ff/sig000010a7 ),
    .Q(sig0000082c)
  );
  SRLC32E #(
    .INIT ( 32'h00000000 ))
  \blk000007fe/blk000007ff/blk0000080e  (
    .CLK(clk),
    .D(sig0000083e),
    .CE(sig00000001),
    .Q(\blk000007fe/blk000007ff/sig000010a7 ),
    .Q31(\NLW_blk000007fe/blk000007ff/blk0000080e_Q31_UNCONNECTED ),
    .A({\blk000007fe/blk000007ff/sig000010a0 , \blk000007fe/blk000007ff/sig0000109f , \blk000007fe/blk000007ff/sig0000109f ,
\blk000007fe/blk000007ff/sig000010a0 , \blk000007fe/blk000007ff/sig000010a0 })
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000007fe/blk000007ff/blk0000080d  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk000007fe/blk000007ff/sig000010a6 ),
    .Q(sig0000082b)
  );
  SRLC32E #(
    .INIT ( 32'h00000000 ))
  \blk000007fe/blk000007ff/blk0000080c  (
    .CLK(clk),
    .D(sig0000083d),
    .CE(sig00000001),
    .Q(\blk000007fe/blk000007ff/sig000010a6 ),
    .Q31(\NLW_blk000007fe/blk000007ff/blk0000080c_Q31_UNCONNECTED ),
    .A({\blk000007fe/blk000007ff/sig000010a0 , \blk000007fe/blk000007ff/sig0000109f , \blk000007fe/blk000007ff/sig0000109f ,
\blk000007fe/blk000007ff/sig000010a0 , \blk000007fe/blk000007ff/sig000010a0 })
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000007fe/blk000007ff/blk0000080b  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk000007fe/blk000007ff/sig000010a5 ),
    .Q(sig0000082a)
  );
  SRLC32E #(
    .INIT ( 32'h00000000 ))
  \blk000007fe/blk000007ff/blk0000080a  (
    .CLK(clk),
    .D(sig0000083c),
    .CE(sig00000001),
    .Q(\blk000007fe/blk000007ff/sig000010a5 ),
    .Q31(\NLW_blk000007fe/blk000007ff/blk0000080a_Q31_UNCONNECTED ),
    .A({\blk000007fe/blk000007ff/sig000010a0 , \blk000007fe/blk000007ff/sig0000109f , \blk000007fe/blk000007ff/sig0000109f ,
\blk000007fe/blk000007ff/sig000010a0 , \blk000007fe/blk000007ff/sig000010a0 })
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000007fe/blk000007ff/blk00000809  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk000007fe/blk000007ff/sig000010a4 ),
    .Q(sig00000829)
  );
  SRLC32E #(
    .INIT ( 32'h00000000 ))
  \blk000007fe/blk000007ff/blk00000808  (
    .CLK(clk),
    .D(sig0000083b),
    .CE(sig00000001),
    .Q(\blk000007fe/blk000007ff/sig000010a4 ),
    .Q31(\NLW_blk000007fe/blk000007ff/blk00000808_Q31_UNCONNECTED ),
    .A({\blk000007fe/blk000007ff/sig000010a0 , \blk000007fe/blk000007ff/sig0000109f , \blk000007fe/blk000007ff/sig0000109f ,
\blk000007fe/blk000007ff/sig000010a0 , \blk000007fe/blk000007ff/sig000010a0 })
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000007fe/blk000007ff/blk00000807  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk000007fe/blk000007ff/sig000010a3 ),
    .Q(sig00000828)
  );
  SRLC32E #(
    .INIT ( 32'h00000000 ))
  \blk000007fe/blk000007ff/blk00000806  (
    .CLK(clk),
    .D(sig0000083a),
    .CE(sig00000001),
    .Q(\blk000007fe/blk000007ff/sig000010a3 ),
    .Q31(\NLW_blk000007fe/blk000007ff/blk00000806_Q31_UNCONNECTED ),
    .A({\blk000007fe/blk000007ff/sig000010a0 , \blk000007fe/blk000007ff/sig0000109f , \blk000007fe/blk000007ff/sig0000109f ,
\blk000007fe/blk000007ff/sig000010a0 , \blk000007fe/blk000007ff/sig000010a0 })
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000007fe/blk000007ff/blk00000805  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk000007fe/blk000007ff/sig000010a2 ),
    .Q(sig00000827)
  );
  SRLC32E #(
    .INIT ( 32'h00000000 ))
  \blk000007fe/blk000007ff/blk00000804  (
    .CLK(clk),
    .D(sig00000839),
    .CE(sig00000001),
    .Q(\blk000007fe/blk000007ff/sig000010a2 ),
    .Q31(\NLW_blk000007fe/blk000007ff/blk00000804_Q31_UNCONNECTED ),
    .A({\blk000007fe/blk000007ff/sig000010a0 , \blk000007fe/blk000007ff/sig0000109f , \blk000007fe/blk000007ff/sig0000109f ,
\blk000007fe/blk000007ff/sig000010a0 , \blk000007fe/blk000007ff/sig000010a0 })
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000007fe/blk000007ff/blk00000803  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk000007fe/blk000007ff/sig000010a1 ),
    .Q(sig00000826)
  );
  SRLC32E #(
    .INIT ( 32'h00000000 ))
  \blk000007fe/blk000007ff/blk00000802  (
    .CLK(clk),
    .D(sig00000838),
    .CE(sig00000001),
    .Q(\blk000007fe/blk000007ff/sig000010a1 ),
    .Q31(\NLW_blk000007fe/blk000007ff/blk00000802_Q31_UNCONNECTED ),
    .A({\blk000007fe/blk000007ff/sig000010a0 , \blk000007fe/blk000007ff/sig0000109f , \blk000007fe/blk000007ff/sig0000109f ,
\blk000007fe/blk000007ff/sig000010a0 , \blk000007fe/blk000007ff/sig000010a0 })
  );
  VCC   \blk000007fe/blk000007ff/blk00000801  (
    .P(\blk000007fe/blk000007ff/sig000010a0 )
  );
  GND   \blk000007fe/blk000007ff/blk00000800  (
    .G(\blk000007fe/blk000007ff/sig0000109f )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000852/blk00000853/blk00000857  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk00000852/blk00000853/sig000010bc ),
    .Q(sig00000825)
  );
  SRLC32E #(
    .INIT ( 32'h00000000 ))
  \blk00000852/blk00000853/blk00000856  (
    .CLK(clk),
    .D(sig000007f8),
    .CE(sig00000001),
    .Q(\blk00000852/blk00000853/sig000010bc ),
    .Q31(\NLW_blk00000852/blk00000853/blk00000856_Q31_UNCONNECTED ),
    .A({\blk00000852/blk00000853/sig000010bb , \blk00000852/blk00000853/sig000010ba , \blk00000852/blk00000853/sig000010bb ,
\blk00000852/blk00000853/sig000010ba , \blk00000852/blk00000853/sig000010bb })
  );
  VCC   \blk00000852/blk00000853/blk00000855  (
    .P(\blk00000852/blk00000853/sig000010bb )
  );
  GND   \blk00000852/blk00000853/blk00000854  (
    .G(\blk00000852/blk00000853/sig000010ba )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk00000858/blk00000859/blk0000085d  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk00000858/blk00000859/sig000010c8 ),
    .Q(sig00000008)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk00000858/blk00000859/blk0000085c  (
    .A0(\blk00000858/blk00000859/sig000010c6 ),
    .A1(\blk00000858/blk00000859/sig000010c7 ),
    .A2(\blk00000858/blk00000859/sig000010c6 ),
    .A3(\blk00000858/blk00000859/sig000010c6 ),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig00000837),
    .Q(\blk00000858/blk00000859/sig000010c8 ),
    .Q15(\NLW_blk00000858/blk00000859/blk0000085c_Q15_UNCONNECTED )
  );
  VCC   \blk00000858/blk00000859/blk0000085b  (
    .P(\blk00000858/blk00000859/sig000010c7 )
  );
  GND   \blk00000858/blk00000859/blk0000085a  (
    .G(\blk00000858/blk00000859/sig000010c6 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk0000085e/blk0000085f/blk00000863  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk0000085e/blk0000085f/sig000010d4 ),
    .Q(sig00000007)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk0000085e/blk0000085f/blk00000862  (
    .A0(\blk0000085e/blk0000085f/sig000010d2 ),
    .A1(\blk0000085e/blk0000085f/sig000010d3 ),
    .A2(\blk0000085e/blk0000085f/sig000010d2 ),
    .A3(\blk0000085e/blk0000085f/sig000010d2 ),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig00000836),
    .Q(\blk0000085e/blk0000085f/sig000010d4 ),
    .Q15(\NLW_blk0000085e/blk0000085f/blk00000862_Q15_UNCONNECTED )
  );
  VCC   \blk0000085e/blk0000085f/blk00000861  (
    .P(\blk0000085e/blk0000085f/sig000010d3 )
  );
  GND   \blk0000085e/blk0000085f/blk00000860  (
    .G(\blk0000085e/blk0000085f/sig000010d2 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000008e1/blk000008e2/blk000008e5  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk000008e1/blk000008e2/sig000010df ),
    .Q(sig00000005)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk000008e1/blk000008e2/blk000008e4  (
    .A0(\blk000008e1/blk000008e2/sig000010de ),
    .A1(\blk000008e1/blk000008e2/sig000010de ),
    .A2(\blk000008e1/blk000008e2/sig000010de ),
    .A3(\blk000008e1/blk000008e2/sig000010de ),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig00000008),
    .Q(\blk000008e1/blk000008e2/sig000010df ),
    .Q15(\NLW_blk000008e1/blk000008e2/blk000008e4_Q15_UNCONNECTED )
  );
  VCC   \blk000008e1/blk000008e2/blk000008e3  (
    .P(\blk000008e1/blk000008e2/sig000010de )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000008e6/blk000008e7/blk000008ea  (
    .C(clk),
    .CE(sig00000001),
    .D(\blk000008e6/blk000008e7/sig000010ea ),
    .Q(sig00000004)
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk000008e6/blk000008e7/blk000008e9  (
    .A0(\blk000008e6/blk000008e7/sig000010e9 ),
    .A1(\blk000008e6/blk000008e7/sig000010e9 ),
    .A2(\blk000008e6/blk000008e7/sig000010e9 ),
    .A3(\blk000008e6/blk000008e7/sig000010e9 ),
    .CE(sig00000001),
    .CLK(clk),
    .D(sig00000007),
    .Q(\blk000008e6/blk000008e7/sig000010ea ),
    .Q15(\NLW_blk000008e6/blk000008e7/blk000008e9_Q15_UNCONNECTED )
  );
  VCC   \blk000008e6/blk000008e7/blk000008e8  (
    .P(\blk000008e6/blk000008e7/sig000010e9 )
  );
  INV   \blk00000935/blk0000094d  (
    .I(sig000009c7),
    .O(\blk00000935/sig00001104 )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk00000935/blk0000094c  (
    .I0(sig000009c8),
    .O(\blk00000935/sig0000110a )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk00000935/blk0000094b  (
    .I0(sig000009c9),
    .O(\blk00000935/sig00001109 )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk00000935/blk0000094a  (
    .I0(sig000009ca),
    .O(\blk00000935/sig00001108 )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk00000935/blk00000949  (
    .I0(sig000009cb),
    .O(\blk00000935/sig00001107 )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk00000935/blk00000948  (
    .I0(sig000009cc),
    .O(\blk00000935/sig00001106 )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk00000935/blk00000947  (
    .I0(sig000009cd),
    .O(\blk00000935/sig00001105 )
  );
  MUXCY   \blk00000935/blk00000946  (
    .CI(\blk00000935/sig000010fc ),
    .DI(\blk00000935/sig000010fb ),
    .S(\blk00000935/sig00001104 ),
    .O(\blk00000935/sig00001103 )
  );
  XORCY   \blk00000935/blk00000945  (
    .CI(\blk00000935/sig000010fc ),
    .LI(\blk00000935/sig00001104 ),
    .O(sig000009bf)
  );
  XORCY   \blk00000935/blk00000944  (
    .CI(\blk00000935/sig000010fd ),
    .LI(sig000009ce),
    .O(sig000009c6)
  );
  MUXCY   \blk00000935/blk00000943  (
    .CI(\blk00000935/sig00001103 ),
    .DI(\blk00000935/sig000010fc ),
    .S(\blk00000935/sig0000110a ),
    .O(\blk00000935/sig00001102 )
  );
  XORCY   \blk00000935/blk00000942  (
    .CI(\blk00000935/sig00001103 ),
    .LI(\blk00000935/sig0000110a ),
    .O(sig000009c0)
  );
  MUXCY   \blk00000935/blk00000941  (
    .CI(\blk00000935/sig00001102 ),
    .DI(\blk00000935/sig000010fc ),
    .S(\blk00000935/sig00001109 ),
    .O(\blk00000935/sig00001101 )
  );
  XORCY   \blk00000935/blk00000940  (
    .CI(\blk00000935/sig00001102 ),
    .LI(\blk00000935/sig00001109 ),
    .O(sig000009c1)
  );
  MUXCY   \blk00000935/blk0000093f  (
    .CI(\blk00000935/sig00001101 ),
    .DI(\blk00000935/sig000010fc ),
    .S(\blk00000935/sig00001108 ),
    .O(\blk00000935/sig00001100 )
  );
  XORCY   \blk00000935/blk0000093e  (
    .CI(\blk00000935/sig00001101 ),
    .LI(\blk00000935/sig00001108 ),
    .O(sig000009c2)
  );
  MUXCY   \blk00000935/blk0000093d  (
    .CI(\blk00000935/sig00001100 ),
    .DI(\blk00000935/sig000010fc ),
    .S(\blk00000935/sig00001107 ),
    .O(\blk00000935/sig000010ff )
  );
  XORCY   \blk00000935/blk0000093c  (
    .CI(\blk00000935/sig00001100 ),
    .LI(\blk00000935/sig00001107 ),
    .O(sig000009c3)
  );
  MUXCY   \blk00000935/blk0000093b  (
    .CI(\blk00000935/sig000010ff ),
    .DI(\blk00000935/sig000010fc ),
    .S(\blk00000935/sig00001106 ),
    .O(\blk00000935/sig000010fe )
  );
  XORCY   \blk00000935/blk0000093a  (
    .CI(\blk00000935/sig000010ff ),
    .LI(\blk00000935/sig00001106 ),
    .O(sig000009c4)
  );
  MUXCY   \blk00000935/blk00000939  (
    .CI(\blk00000935/sig000010fe ),
    .DI(\blk00000935/sig000010fc ),
    .S(\blk00000935/sig00001105 ),
    .O(\blk00000935/sig000010fd )
  );
  XORCY   \blk00000935/blk00000938  (
    .CI(\blk00000935/sig000010fe ),
    .LI(\blk00000935/sig00001105 ),
    .O(sig000009c5)
  );
  GND   \blk00000935/blk00000937  (
    .G(\blk00000935/sig000010fc )
  );
  VCC   \blk00000935/blk00000936  (
    .P(\blk00000935/sig000010fb )
  );
  INV   \blk0000095a/blk00000969  (
    .I(sig000009da),
    .O(\blk0000095a/sig0000111b )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk0000095a/blk00000968  (
    .I0(sig000009db),
    .O(\blk0000095a/sig0000111e )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk0000095a/blk00000967  (
    .I0(sig000009dc),
    .O(\blk0000095a/sig0000111d )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk0000095a/blk00000966  (
    .I0(sig000009dd),
    .O(\blk0000095a/sig0000111c )
  );
  MUXCY   \blk0000095a/blk00000965  (
    .CI(\blk0000095a/sig00001116 ),
    .DI(\blk0000095a/sig00001115 ),
    .S(\blk0000095a/sig0000111b ),
    .O(\blk0000095a/sig0000111a )
  );
  XORCY   \blk0000095a/blk00000964  (
    .CI(\blk0000095a/sig00001116 ),
    .LI(\blk0000095a/sig0000111b ),
    .O(sig000009d4)
  );
  XORCY   \blk0000095a/blk00000963  (
    .CI(\blk0000095a/sig00001117 ),
    .LI(sig000009de),
    .O(sig000009d8)
  );
  MUXCY   \blk0000095a/blk00000962  (
    .CI(\blk0000095a/sig0000111a ),
    .DI(\blk0000095a/sig00001116 ),
    .S(\blk0000095a/sig0000111e ),
    .O(\blk0000095a/sig00001119 )
  );
  XORCY   \blk0000095a/blk00000961  (
    .CI(\blk0000095a/sig0000111a ),
    .LI(\blk0000095a/sig0000111e ),
    .O(sig000009d5)
  );
  MUXCY   \blk0000095a/blk00000960  (
    .CI(\blk0000095a/sig00001119 ),
    .DI(\blk0000095a/sig00001116 ),
    .S(\blk0000095a/sig0000111d ),
    .O(\blk0000095a/sig00001118 )
  );
  XORCY   \blk0000095a/blk0000095f  (
    .CI(\blk0000095a/sig00001119 ),
    .LI(\blk0000095a/sig0000111d ),
    .O(sig000009d6)
  );
  MUXCY   \blk0000095a/blk0000095e  (
    .CI(\blk0000095a/sig00001118 ),
    .DI(\blk0000095a/sig00001116 ),
    .S(\blk0000095a/sig0000111c ),
    .O(\blk0000095a/sig00001117 )
  );
  XORCY   \blk0000095a/blk0000095d  (
    .CI(\blk0000095a/sig00001118 ),
    .LI(\blk0000095a/sig0000111c ),
    .O(sig000009d7)
  );
  GND   \blk0000095a/blk0000095c  (
    .G(\blk0000095a/sig00001116 )
  );
  VCC   \blk0000095a/blk0000095b  (
    .P(\blk0000095a/sig00001115 )
  );
  INV   \blk00000974/blk00000980  (
    .I(sig000009ec),
    .O(\blk00000974/sig0000112c )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk00000974/blk0000097f  (
    .I0(sig000009ed),
    .O(\blk00000974/sig0000112e )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk00000974/blk0000097e  (
    .I0(sig000009ee),
    .O(\blk00000974/sig0000112d )
  );
  MUXCY   \blk00000974/blk0000097d  (
    .CI(\blk00000974/sig00001128 ),
    .DI(\blk00000974/sig00001127 ),
    .S(\blk00000974/sig0000112c ),
    .O(\blk00000974/sig0000112b )
  );
  XORCY   \blk00000974/blk0000097c  (
    .CI(\blk00000974/sig00001128 ),
    .LI(\blk00000974/sig0000112c ),
    .O(sig000009e8)
  );
  XORCY   \blk00000974/blk0000097b  (
    .CI(\blk00000974/sig00001129 ),
    .LI(sig000009ef),
    .O(sig000009eb)
  );
  MUXCY   \blk00000974/blk0000097a  (
    .CI(\blk00000974/sig0000112b ),
    .DI(\blk00000974/sig00001128 ),
    .S(\blk00000974/sig0000112e ),
    .O(\blk00000974/sig0000112a )
  );
  XORCY   \blk00000974/blk00000979  (
    .CI(\blk00000974/sig0000112b ),
    .LI(\blk00000974/sig0000112e ),
    .O(sig000009e9)
  );
  MUXCY   \blk00000974/blk00000978  (
    .CI(\blk00000974/sig0000112a ),
    .DI(\blk00000974/sig00001128 ),
    .S(\blk00000974/sig0000112d ),
    .O(\blk00000974/sig00001129 )
  );
  XORCY   \blk00000974/blk00000977  (
    .CI(\blk00000974/sig0000112a ),
    .LI(\blk00000974/sig0000112d ),
    .O(sig000009ea)
  );
  GND   \blk00000974/blk00000976  (
    .G(\blk00000974/sig00001128 )
  );
  VCC   \blk00000974/blk00000975  (
    .P(\blk00000974/sig00001127 )
  );
  INV   \blk00000981/blk0000099c  (
    .I(sig0000096d),
    .O(\blk00000981/sig0000114b )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk00000981/blk0000099b  (
    .I0(sig0000096c),
    .O(\blk00000981/sig00001152 )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk00000981/blk0000099a  (
    .I0(sig0000096b),
    .O(\blk00000981/sig00001151 )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk00000981/blk00000999  (
    .I0(sig0000096a),
    .O(\blk00000981/sig00001150 )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk00000981/blk00000998  (
    .I0(sig00000969),
    .O(\blk00000981/sig0000114f )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk00000981/blk00000997  (
    .I0(sig00000968),
    .O(\blk00000981/sig0000114e )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk00000981/blk00000996  (
    .I0(sig00000967),
    .O(\blk00000981/sig0000114d )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk00000981/blk00000995  (
    .I0(sig00000966),
    .O(\blk00000981/sig0000114c )
  );
  MUXCY   \blk00000981/blk00000994  (
    .CI(\blk00000981/sig00001142 ),
    .DI(\blk00000981/sig00001141 ),
    .S(\blk00000981/sig0000114b ),
    .O(\blk00000981/sig0000114a )
  );
  XORCY   \blk00000981/blk00000993  (
    .CI(\blk00000981/sig00001142 ),
    .LI(\blk00000981/sig0000114b ),
    .O(sig00000976)
  );
  XORCY   \blk00000981/blk00000992  (
    .CI(\blk00000981/sig00001143 ),
    .LI(sig00000965),
    .O(sig0000096e)
  );
  MUXCY   \blk00000981/blk00000991  (
    .CI(\blk00000981/sig0000114a ),
    .DI(\blk00000981/sig00001142 ),
    .S(\blk00000981/sig00001152 ),
    .O(\blk00000981/sig00001149 )
  );
  XORCY   \blk00000981/blk00000990  (
    .CI(\blk00000981/sig0000114a ),
    .LI(\blk00000981/sig00001152 ),
    .O(sig00000975)
  );
  MUXCY   \blk00000981/blk0000098f  (
    .CI(\blk00000981/sig00001149 ),
    .DI(\blk00000981/sig00001142 ),
    .S(\blk00000981/sig00001151 ),
    .O(\blk00000981/sig00001148 )
  );
  XORCY   \blk00000981/blk0000098e  (
    .CI(\blk00000981/sig00001149 ),
    .LI(\blk00000981/sig00001151 ),
    .O(sig00000974)
  );
  MUXCY   \blk00000981/blk0000098d  (
    .CI(\blk00000981/sig00001148 ),
    .DI(\blk00000981/sig00001142 ),
    .S(\blk00000981/sig00001150 ),
    .O(\blk00000981/sig00001147 )
  );
  XORCY   \blk00000981/blk0000098c  (
    .CI(\blk00000981/sig00001148 ),
    .LI(\blk00000981/sig00001150 ),
    .O(sig00000973)
  );
  MUXCY   \blk00000981/blk0000098b  (
    .CI(\blk00000981/sig00001147 ),
    .DI(\blk00000981/sig00001142 ),
    .S(\blk00000981/sig0000114f ),
    .O(\blk00000981/sig00001146 )
  );
  XORCY   \blk00000981/blk0000098a  (
    .CI(\blk00000981/sig00001147 ),
    .LI(\blk00000981/sig0000114f ),
    .O(sig00000972)
  );
  MUXCY   \blk00000981/blk00000989  (
    .CI(\blk00000981/sig00001146 ),
    .DI(\blk00000981/sig00001142 ),
    .S(\blk00000981/sig0000114e ),
    .O(\blk00000981/sig00001145 )
  );
  XORCY   \blk00000981/blk00000988  (
    .CI(\blk00000981/sig00001146 ),
    .LI(\blk00000981/sig0000114e ),
    .O(sig00000971)
  );
  MUXCY   \blk00000981/blk00000987  (
    .CI(\blk00000981/sig00001145 ),
    .DI(\blk00000981/sig00001142 ),
    .S(\blk00000981/sig0000114d ),
    .O(\blk00000981/sig00001144 )
  );
  XORCY   \blk00000981/blk00000986  (
    .CI(\blk00000981/sig00001145 ),
    .LI(\blk00000981/sig0000114d ),
    .O(sig00000970)
  );
  MUXCY   \blk00000981/blk00000985  (
    .CI(\blk00000981/sig00001144 ),
    .DI(\blk00000981/sig00001142 ),
    .S(\blk00000981/sig0000114c ),
    .O(\blk00000981/sig00001143 )
  );
  XORCY   \blk00000981/blk00000984  (
    .CI(\blk00000981/sig00001144 ),
    .LI(\blk00000981/sig0000114c ),
    .O(sig0000096f)
  );
  GND   \blk00000981/blk00000983  (
    .G(\blk00000981/sig00001142 )
  );
  VCC   \blk00000981/blk00000982  (
    .P(\blk00000981/sig00001141 )
  );
  INV   \blk0000099d/blk000009b8  (
    .I(sig00000980),
    .O(\blk0000099d/sig0000116f )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk0000099d/blk000009b7  (
    .I0(sig0000097f),
    .O(\blk0000099d/sig00001176 )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk0000099d/blk000009b6  (
    .I0(sig0000097e),
    .O(\blk0000099d/sig00001175 )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk0000099d/blk000009b5  (
    .I0(sig0000097d),
    .O(\blk0000099d/sig00001174 )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk0000099d/blk000009b4  (
    .I0(sig0000097c),
    .O(\blk0000099d/sig00001173 )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk0000099d/blk000009b3  (
    .I0(sig0000097b),
    .O(\blk0000099d/sig00001172 )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk0000099d/blk000009b2  (
    .I0(sig0000097a),
    .O(\blk0000099d/sig00001171 )
  );
  LUT1 #(
    .INIT ( 2'h2 ))
  \blk0000099d/blk000009b1  (
    .I0(sig00000979),
    .O(\blk0000099d/sig00001170 )
  );
  MUXCY   \blk0000099d/blk000009b0  (
    .CI(\blk0000099d/sig00001166 ),
    .DI(\blk0000099d/sig00001165 ),
    .S(\blk0000099d/sig0000116f ),
    .O(\blk0000099d/sig0000116e )
  );
  XORCY   \blk0000099d/blk000009af  (
    .CI(\blk0000099d/sig00001166 ),
    .LI(\blk0000099d/sig0000116f ),
    .O(sig00000989)
  );
  XORCY   \blk0000099d/blk000009ae  (
    .CI(\blk0000099d/sig00001167 ),
    .LI(sig00000978),
    .O(sig00000981)
  );
  MUXCY   \blk0000099d/blk000009ad  (
    .CI(\blk0000099d/sig0000116e ),
    .DI(\blk0000099d/sig00001166 ),
    .S(\blk0000099d/sig00001176 ),
    .O(\blk0000099d/sig0000116d )
  );
  XORCY   \blk0000099d/blk000009ac  (
    .CI(\blk0000099d/sig0000116e ),
    .LI(\blk0000099d/sig00001176 ),
    .O(sig00000988)
  );
  MUXCY   \blk0000099d/blk000009ab  (
    .CI(\blk0000099d/sig0000116d ),
    .DI(\blk0000099d/sig00001166 ),
    .S(\blk0000099d/sig00001175 ),
    .O(\blk0000099d/sig0000116c )
  );
  XORCY   \blk0000099d/blk000009aa  (
    .CI(\blk0000099d/sig0000116d ),
    .LI(\blk0000099d/sig00001175 ),
    .O(sig00000987)
  );
  MUXCY   \blk0000099d/blk000009a9  (
    .CI(\blk0000099d/sig0000116c ),
    .DI(\blk0000099d/sig00001166 ),
    .S(\blk0000099d/sig00001174 ),
    .O(\blk0000099d/sig0000116b )
  );
  XORCY   \blk0000099d/blk000009a8  (
    .CI(\blk0000099d/sig0000116c ),
    .LI(\blk0000099d/sig00001174 ),
    .O(sig00000986)
  );
  MUXCY   \blk0000099d/blk000009a7  (
    .CI(\blk0000099d/sig0000116b ),
    .DI(\blk0000099d/sig00001166 ),
    .S(\blk0000099d/sig00001173 ),
    .O(\blk0000099d/sig0000116a )
  );
  XORCY   \blk0000099d/blk000009a6  (
    .CI(\blk0000099d/sig0000116b ),
    .LI(\blk0000099d/sig00001173 ),
    .O(sig00000985)
  );
  MUXCY   \blk0000099d/blk000009a5  (
    .CI(\blk0000099d/sig0000116a ),
    .DI(\blk0000099d/sig00001166 ),
    .S(\blk0000099d/sig00001172 ),
    .O(\blk0000099d/sig00001169 )
  );
  XORCY   \blk0000099d/blk000009a4  (
    .CI(\blk0000099d/sig0000116a ),
    .LI(\blk0000099d/sig00001172 ),
    .O(sig00000984)
  );
  MUXCY   \blk0000099d/blk000009a3  (
    .CI(\blk0000099d/sig00001169 ),
    .DI(\blk0000099d/sig00001166 ),
    .S(\blk0000099d/sig00001171 ),
    .O(\blk0000099d/sig00001168 )
  );
  XORCY   \blk0000099d/blk000009a2  (
    .CI(\blk0000099d/sig00001169 ),
    .LI(\blk0000099d/sig00001171 ),
    .O(sig00000983)
  );
  MUXCY   \blk0000099d/blk000009a1  (
    .CI(\blk0000099d/sig00001168 ),
    .DI(\blk0000099d/sig00001166 ),
    .S(\blk0000099d/sig00001170 ),
    .O(\blk0000099d/sig00001167 )
  );
  XORCY   \blk0000099d/blk000009a0  (
    .CI(\blk0000099d/sig00001168 ),
    .LI(\blk0000099d/sig00001170 ),
    .O(sig00000982)
  );
  GND   \blk0000099d/blk0000099f  (
    .G(\blk0000099d/sig00001166 )
  );
  VCC   \blk0000099d/blk0000099e  (
    .P(\blk0000099d/sig00001165 )
  );
  FDE #(
    .INIT ( 1'b0 ))
  \blk000009cb/blk000009cc/blk000009d2  (
    .C(clk),
    .CE(\blk000009cb/blk000009cc/sig00001182 ),
    .D(\blk000009cb/blk000009cc/sig00001183 ),
    .Q(\blk000009cb/blk000009cc/sig0000117f )
  );
  SRLC16E #(
    .INIT ( 16'h0000 ))
  \blk000009cb/blk000009cc/blk000009d1  (
    .A0(\blk000009cb/blk000009cc/sig00001182 ),
    .A1(\blk000009cb/blk000009cc/sig00001182 ),
    .A2(\blk000009cb/blk000009cc/sig00001181 ),
    .A3(\blk000009cb/blk000009cc/sig00001181 ),
    .CE(\blk000009cb/blk000009cc/sig00001182 ),
    .CLK(clk),
    .D(sig000007f9),
    .Q(\blk000009cb/blk000009cc/sig00001183 ),
    .Q15(\NLW_blk000009cb/blk000009cc/blk000009d1_Q15_UNCONNECTED )
  );
  VCC   \blk000009cb/blk000009cc/blk000009d0  (
    .P(\blk000009cb/blk000009cc/sig00001182 )
  );
  GND   \blk000009cb/blk000009cc/blk000009cf  (
    .G(\blk000009cb/blk000009cc/sig00001181 )
  );
  FD #(
    .INIT ( 1'b0 ))
  \blk000009cb/blk000009cc/blk000009ce  (
    .C(clk),
    .D(\blk000009cb/blk000009cc/sig00001180 ),
    .Q(dv)
  );
  LUT2 #(
    .INIT ( 4'h4 ))
  \blk000009cb/blk000009cc/blk000009cd  (
    .I0(sig00000002),
    .I1(\blk000009cb/blk000009cc/sig0000117f ),
    .O(\blk000009cb/blk000009cc/sig00001180 )
  );
// synthesis translate_on
endmodule