module header
	// Internal signals
	// Generated Signal List
		wire		mix_logic0_0;
	// End of Generated Signal List
	// %COMPILER_OPTS%
	// Generated Signal Assignments
		assign	mix_logic0_0 = 1'b0;
	// Generated Instances and Port Mappings
		// Generated Instance Port Map for inst_a
		ent_a inst_a (
			.low_bit_a(mix_logic0_0)	// Ground bit port
		);
		// End of Generated Instance Port Map for inst_a
		// Generated Instance Port Map for inst_b
		ent_b inst_b (
		);
		// End of Generated Instance Port Map for inst_b
endmodule