module main;
   test tt();
   defparam tt.foo = 4;
endmodule