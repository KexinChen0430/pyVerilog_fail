module
assign daisy_p_o = 1'bz;
assign daisy_n_o = 1'bz;
endmodule