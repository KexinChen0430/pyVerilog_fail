module
         .sys_reset_out                   (sys_reset_out),
         .tx_out_clk                      (tx_out_clk)
     );
 endmodule