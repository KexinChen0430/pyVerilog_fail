module b14_inj (clock,reset,addr,datai,datao,rd,wr,p_b_Z_p_O_FDC,p_desc52_p_O_FDC,p_desc53_p_O_FDC,p_desc54_p_O_FDC,p_desc55_p_O_FDC,p_desc56_p_O_FDC,p_desc57_p_O_FDC,p_desc58_p_O_FDC,p_desc59_p_O_FDC,p_desc60_p_O_FDC,p_desc61_p_O_FDC,p_desc62_p_O_FDC,p_desc63_p_O_FDC,p_desc64_p_O_FDC,p_desc65_p_O_FDC,p_desc66_p_O_FDC,p_desc67_p_O_FDC,p_desc68_p_O_FDC,p_desc69_p_O_FDC,p_desc70_p_O_FDC,p_desc71_p_O_FDC,p_desc72_p_O_FDC,p_desc73_p_O_FDC,p_desc74_p_O_FDC,p_desc75_p_O_FDC,p_desc76_p_O_FDC,p_desc77_p_O_FDC,p_desc78_p_O_FDC,p_desc79_p_O_FDC,p_desc80_p_O_FDC,p_desc81_p_O_FDC,p_desc82_p_O_FDC,p_desc83_p_O_FDC,p_rd_Z_p_O_FDC,p_desc261_p_O_FDC,p_wr_Z_p_O_FDC,p_desc262_p_O_FDC,p_desc50_p_O_FDCE,p_desc51_p_O_FDCE,p_desc84_p_O_FDCE,p_desc85_p_O_FDCE,p_desc86_p_O_FDCE,p_desc87_p_O_FDCE,p_desc88_p_O_FDCE,p_desc89_p_O_FDCE,p_desc90_p_O_FDCE,p_desc91_p_O_FDCE,p_desc92_p_O_FDCE,p_desc93_p_O_FDCE,p_desc94_p_O_FDCE,p_desc95_p_O_FDCE,p_desc96_p_O_FDCE,p_desc97_p_O_FDCE,p_desc98_p_O_FDCE,p_desc99_p_O_FDCE,p_desc100_p_O_FDCE,p_desc101_p_O_FDCE,p_desc102_p_O_FDCE,p_desc103_p_O_FDCE,p_desc104_p_O_FDCE,p_desc105_p_O_FDCE,p_desc106_p_O_FDCE,p_desc107_p_O_FDCE,p_desc108_p_O_FDCE,p_desc109_p_O_FDCE,p_desc110_p_O_FDCE,p_desc111_p_O_FDCE,p_desc112_p_O_FDCE,p_desc113_p_O_FDCE,p_desc114_p_O_FDCE,p_desc115_p_O_FDCE,p_desc116_p_O_FDCE,p_desc117_p_O_FDCE,p_desc118_p_O_FDCE,p_desc119_p_O_FDCE,p_desc120_p_O_FDCE,p_desc121_p_O_FDCE,p_desc122_p_O_FDCE,p_desc123_p_O_FDCE,p_desc124_p_O_FDCE,p_desc125_p_O_FDCE,p_desc126_p_O_FDCE,p_desc127_p_O_FDCE,p_desc128_p_O_FDCE,p_desc129_p_O_FDCE,p_desc130_p_O_FDCE,p_desc131_p_O_FDCE,p_desc132_p_O_FDCE,p_desc133_p_O_FDCE,p_desc134_p_O_FDCE,p_desc135_p_O_FDCE,p_desc136_p_O_FDCE,p_desc137_p_O_FDCE,p_desc138_p_O_FDCE,p_desc139_p_O_FDCE,p_desc140_p_O_FDCE,p_desc141_p_O_FDCE,p_desc142_p_O_FDCE,p_desc143_p_O_FDCE,p_desc144_p_O_FDCE,p_desc145_p_O_FDCE,p_desc146_p_O_FDCE,p_desc147_p_O_FDCE,p_desc148_p_O_FDCE,p_desc149_p_O_FDCE,p_desc150_p_O_FDCE,p_desc151_p_O_FDCE,p_desc152_p_O_FDCE,p_desc153_p_O_FDCE,p_desc154_p_O_FDCE,p_desc155_p_O_FDCE,p_desc156_p_O_FDCE,p_desc157_p_O_FDCE,p_desc158_p_O_FDCE,p_desc159_p_O_FDCE,p_desc160_p_O_FDCE,p_desc161_p_O_FDCE,p_desc162_p_O_FDCE,p_desc163_p_O_FDCE,p_desc164_p_O_FDCE,p_desc165_p_O_FDCE,p_desc166_p_O_FDCE,p_desc167_p_O_FDCE,p_desc168_p_O_FDCE,p_desc169_p_O_FDCE,p_desc170_p_O_FDCE,p_desc171_p_O_FDCE,p_desc172_p_O_FDCE,p_desc173_p_O_FDCE,p_desc174_p_O_FDCE,p_desc175_p_O_FDCE,p_desc176_p_O_FDCE,p_desc177_p_O_FDCE,p_desc178_p_O_FDCE,p_desc179_p_O_FDCE,p_desc180_p_O_FDCE,p_desc181_p_O_FDCE,p_desc182_p_O_FDCE,p_desc183_p_O_FDCE,p_desc184_p_O_FDCE,p_desc185_p_O_FDCE,p_desc186_p_O_FDCE,p_desc187_p_O_FDCE,p_desc188_p_O_FDCE,p_desc189_p_O_FDCE,p_desc190_p_O_FDCE,p_desc191_p_O_FDCE,p_desc192_p_O_FDCE,p_desc193_p_O_FDCE,p_desc194_p_O_FDCE,p_desc195_p_O_FDCE,p_desc196_p_O_FDCE,p_desc197_p_O_FDCE,p_desc198_p_O_FDCE,p_desc199_p_O_FDCE,p_desc200_p_O_FDCE,p_desc201_p_O_FDCE,p_desc202_p_O_FDCE,p_desc203_p_O_FDCE,p_desc204_p_O_FDCE,p_desc205_p_O_FDCE,p_desc206_p_O_FDCE,p_desc207_p_O_FDCE,p_desc208_p_O_FDCE,p_desc209_p_O_FDCE,p_desc210_p_O_FDCE,p_desc211_p_O_FDCE,p_desc212_p_O_FDCE,p_desc213_p_O_FDCE,p_desc214_p_O_FDCE,p_desc215_p_O_FDCE,p_desc216_p_O_FDCE,p_desc217_p_O_FDCE,p_desc218_p_O_FDCE,p_desc219_p_O_FDCE,p_desc220_p_O_FDCE,p_desc221_p_O_FDCE,p_desc222_p_O_FDCE,p_desc223_p_O_FDCE,p_desc224_p_O_FDCE,p_desc225_p_O_FDCE,p_desc226_p_O_FDCE,p_desc227_p_O_FDCE,p_desc228_p_O_FDCE,p_desc229_p_O_FDCE,p_desc230_p_O_FDCE,p_desc231_p_O_FDCE,p_desc232_p_O_FDCE,p_desc233_p_O_FDCE,p_desc234_p_O_FDCE,p_desc235_p_O_FDCE,p_desc236_p_O_FDCE,p_desc237_p_O_FDCE,p_desc238_p_O_FDCE,p_desc239_p_O_FDCE,p_desc240_p_O_FDCE,p_desc241_p_O_FDCE,p_desc242_p_O_FDCE,p_desc243_p_O_FDCE,p_desc244_p_O_FDCE,p_desc245_p_O_FDCE,p_desc246_p_O_FDCE,p_desc247_p_O_FDCE,p_desc248_p_O_FDCE,p_desc249_p_O_FDCE,p_desc250_p_O_FDCE,p_desc251_p_O_FDCE,p_desc252_p_O_FDCE,p_desc253_p_O_FDCE,p_desc254_p_O_FDCE,p_desc255_p_O_FDCE,p_desc256_p_O_FDCE,p_desc257_p_O_FDCE,p_desc258_p_O_FDCE,p_desc259_p_O_FDCE,p_desc260_p_O_FDCE);
input clock ;
input reset ;
output [19:0] addr ;
input [31:0] datai ;
output [31:0] datao ;
output rd ;
output wr ;
wire clock ;
wire reset ;
wire rd ;
wire wr ;
wire state ;
wire [31:0] ir ;
wire [28:0] reg3 ;
wire [31:0] ir_3 ;
wire [31:0] reg2 ;
wire [31:0] m_2 ;
wire [31:0] reg1 ;
wire [31:0] r_4 ;
wire [31:0] reg0 ;
wire [30:0] un11_r_cry ;
wire [1:0] d ;
wire [30:30] r_6 ;
wire [30:0] un26_r_cry ;
wire [31:0] reg2_16 ;
wire [19:0] un1_inf_abs0_10 ;
wire [19:0] un1_inf_abs0_11 ;
wire [18:0] reg0_28 ;
wire [18:0] reg1_16 ;
wire [28:0] reg3_17 ;
wire [28:0] b18_cry ;
wire [30:30] r_4_3_lut6_2_O5 ;
wire [9:0] un14_r_0_data_tmp ;
wire [16:1] t_6 ;
wire d_cnst ;
wire dce ;
wire [31:0] inf_abs0_2 ;
wire [31:1] reg3_1_1 ;
wire [31:0] t_1 ;
wire [18:17] reg0_28_7_a1 ;
wire [24:24] reg0_28_7_d ;
wire [24:21] reg3_17_a0 ;
wire [29:29] reg2_16_11_a1 ;
wire [29:17] reg2_16_11_a2 ;
wire [29:17] reg2_16_11_a3 ;
wire [1:0] r_4_2_a0 ;
wire [13:13] reg3_17_4_a2 ;
wire [10:10] r_4_1_RNIDBOH1 ;
wire [25:21] reg2_16_11_a4 ;
wire [9:9] r_4_1_RNIS3K91 ;
wire [7:7] r_4_1_RNIFO731 ;
wire [8:8] r_4_1_RNIIQ731 ;
wire [5:5] r_4_1_RNI9K731 ;
wire [6:6] r_4_1_RNICM731 ;
wire [3:3] r_4_2_a1_lut6_2_RNI5V8R3 ;
wire [3:3] r_4_2_a1_lut6_2_RNI2T8R3 ;
wire [24:21] \d_cnst_sn.reg3_17_0_tz  ;
wire [4:0] \d_cnst_sn.r_4_0_0  ;
wire [20:20] reg2_16_2_d ;
wire [3:3] r_4_2_a1_lut6_2_O6 ;
wire [3:3] r_4_2_a1_lut6_2_O5 ;
wire [28:28] \d_cnst_sn.reg2_16_0_1_tz  ;
wire [28:28] \d_cnst_sn.reg2_16_11_1_tz  ;
wire [7:7] \d_cnst_sn.reg0_28_a0_1  ;
wire [5:5] \d_cnst_sn.reg1_16_a2_0  ;
wire [4:4] \d_cnst_sn.reg0_28_a1_1  ;
wire [3:3] \d_cnst_sn.reg1_16_a0_1  ;
wire [9:9] \d_cnst_sn.reg0_28_7_a0_0  ;
wire [24:24] \d_cnst_sn.reg3_17_a1_2  ;
wire state_i ;
wire [31:31] r_4_i ;
wire [31:0] m_2_i ;
wire [28:20] \d_cnst_sn.reg3_17_4_a2_0  ;
wire [21:21] \d_cnst_sn.reg3_17_a2_2_0  ;
wire [8:2] \d_cnst_sn.reg0_1  ;
wire [8:3] \d_cnst_sn.reg1_1  ;
wire [28:12] \d_cnst_sn.reg3_17_6_0  ;
wire [19:12] \d_cnst_sn.reg3_17_6_1  ;
wire [20:19] \d_cnst_sn.reg0_28_0  ;
wire [25:20] \d_cnst_sn.reg2_16_0  ;
wire [29:20] \d_cnst_sn.reg2_16_1  ;
wire [17:17] \d_cnst_sn.reg0_0  ;
wire [18:18] \d_cnst_sn.reg1_0  ;
wire [28:26] \d_cnst_sn.reg2_16_0_1_0  ;
wire [31:31] r_4_3_ci ;
wire [31:31] ir_fast ;
wire [31:31] ir_3_fast ;
wire [31:31] inf_abs0_2_0 ;
wire [31:31] inf_abs0_2_1 ;
wire [1:1] \d_cnst_sn.reg2_16_11muxnet_0  ;
wire [1:1] \d_cnst_sn.reg2_16_11muxnet_1  ;
wire b ;
wire VCC ;
wire GND ;
wire addr_4_sqmuxa_1 ;
wire un14_r_0_I_83 ;
wire b18 ;
wire un11_reg0_s_1 ;
wire un11_reg0_s_2 ;
wire un11_reg0_s_3 ;
wire un11_reg0_s_4 ;
wire un11_reg0_s_5 ;
wire un11_reg0_s_6 ;
wire un11_reg0_s_7 ;
wire un11_reg0_s_8 ;
wire un11_reg0_s_9 ;
wire un11_reg0_s_10 ;
wire un11_reg0_s_11 ;
wire un11_reg0_s_12 ;
wire un11_reg0_s_13 ;
wire un11_reg0_s_14 ;
wire un11_reg0_s_15 ;
wire un11_reg0_s_16 ;
wire un11_reg0_s_17 ;
wire un11_reg0_s_18 ;
wire un11_reg0_s_19 ;
wire un11_reg0_s_20 ;
wire un11_reg0_s_21 ;
wire un11_reg0_s_22 ;
wire un11_reg0_s_23 ;
wire un11_reg0_s_24 ;
wire un11_reg0_s_25 ;
wire un11_reg0_s_26 ;
wire un11_reg0_s_27 ;
wire un11_reg0_s_28 ;
wire un11_reg0_s_29 ;
wire rd_18 ;
wire un11_r_df0 ;
wire un11_r_lt0 ;
wire un11_r_df2 ;
wire un11_r_lt2 ;
wire un11_r_df4 ;
wire un11_r_lt4 ;
wire un11_r_df6 ;
wire un11_r_lt6 ;
wire un11_r_df8 ;
wire un11_r_lt8 ;
wire un11_r_df10 ;
wire un11_r_lt10 ;
wire un11_r_df12 ;
wire un11_r_lt12 ;
wire un11_r_df14 ;
wire un11_r_lt14 ;
wire un11_r_df16 ;
wire un11_r_lt16 ;
wire un11_r_df18 ;
wire un11_r_lt18 ;
wire un11_r_df20 ;
wire un11_r_lt20 ;
wire un11_r_df22 ;
wire un11_r_lt22 ;
wire un11_r_df24 ;
wire un11_r_lt24 ;
wire un11_r_df26 ;
wire un11_r_lt26 ;
wire un11_r_df28 ;
wire un11_r_lt28 ;
wire un11_r_df30 ;
wire un11_r_lt30 ;
wire b18_df0 ;
wire b18_lt0 ;
wire b18_df2 ;
wire b18_lt2 ;
wire b18_df4 ;
wire b18_lt4 ;
wire b18_df6 ;
wire b18_lt6 ;
wire b18_df8 ;
wire b18_lt8 ;
wire b18_df10 ;
wire b18_lt10 ;
wire b18_df12 ;
wire b18_lt12 ;
wire b18_df14 ;
wire b18_lt14 ;
wire b18_df16 ;
wire b18_lt16 ;
wire b18_df18 ;
wire b18_lt18 ;
wire b18_df20 ;
wire b18_lt20 ;
wire b18_df22 ;
wire b18_lt22 ;
wire b18_df24 ;
wire b18_lt24 ;
wire b18_df26 ;
wire b18_lt26 ;
wire b18_df28 ;
wire b18_lt28 ;
wire b18_df30 ;
wire b18_lt30 ;
wire un26_r_df0 ;
wire un26_r_lt0 ;
wire un26_r_df2 ;
wire un26_r_lt2 ;
wire un26_r_df4 ;
wire un26_r_lt4 ;
wire un26_r_df6 ;
wire un26_r_lt6 ;
wire un26_r_df8 ;
wire un26_r_lt8 ;
wire un26_r_df10 ;
wire un26_r_lt10 ;
wire un26_r_df12 ;
wire un26_r_lt12 ;
wire un26_r_df14 ;
wire un26_r_lt14 ;
wire un26_r_df16 ;
wire un26_r_lt16 ;
wire un26_r_df18 ;
wire un26_r_lt18 ;
wire un26_r_df20 ;
wire un26_r_lt20 ;
wire un26_r_df22 ;
wire un26_r_lt22 ;
wire un26_r_df24 ;
wire un26_r_lt24 ;
wire un26_r_df26 ;
wire un26_r_lt26 ;
wire un26_r_df28 ;
wire un26_r_lt28 ;
wire un26_r_df30 ;
wire un26_r_lt30 ;
wire r_4_3_30_680_i_m2 ;
wire r_4_3_29_706_i_m2 ;
wire r_4_3_28_732_i_m2 ;
wire r_4_3_27_758_i_m2 ;
wire r_4_3_25_810_i_m2 ;
wire r_4_3_24_836_i_m2 ;
wire r_4_3_23_1078_i_m2 ;
wire r_4_3_22_1104_i_m2 ;
wire r_4_3_20_1156_i_m2 ;
wire r_4_3_19_1182_i_m2 ;
wire r_4_3_18_1208_i_m2 ;
wire r_4_3_17_1234_i_m2 ;
wire r_4_3_16_1260_i_m2 ;
wire r_4_3_15_1286_i_m2 ;
wire r_4_3_14_1312_i_m2 ;
wire r_4_3_13_1338_i_m2 ;
wire r_4_3_12_1364_i_m2 ;
wire r_4_3_11_1390_i_m2 ;
wire r_4_3_10_1416_i_m2 ;
wire r_4_3_9_1442_i_m2 ;
wire r_4_3_8_1467 ;
wire r_4_3_6_1508_i_m2 ;
wire r_4_3_5_1534_i_m2 ;
wire r_4_3_4_1560_i_m2 ;
wire r_4_3_3_1586_i_m2 ;
wire r_4_3_2_1612_i_m2 ;
wire r_4_3_1_1638_i_m2 ;
wire r_4_3_0_1664_i_m2 ;
wire r_4_3_1690_i_m2 ;
wire reg1_16_9 ;
wire reg1_16_8_1837 ;
wire reg1_16_7_1870 ;
wire reg0_28_10_2261_a6_3_2_lut6_2_RNIOK9O5 ;
wire reg0_28_8_2327 ;
wire reg0_28_7_2360 ;
wire reg0_28_6_2393 ;
wire reg0_28_5_2426 ;
wire reg0_28_4_2459 ;
wire reg0_28_3_2492 ;
wire un14_r_0_N_2 ;
wire un14_r_0_N_7 ;
wire un14_r_0_N_14 ;
wire un14_r_0_N_21 ;
wire un14_r_0_N_28 ;
wire un14_r_0_N_35 ;
wire un14_r_0_N_42 ;
wire un14_r_0_N_49 ;
wire un14_r_0_N_56 ;
wire un14_r_0_N_63 ;
wire un14_r_0_N_70 ;
wire N_28 ;
wire N_3550 ;
wire N_3856 ;
wire N_2724 ;
wire N_3673 ;
wire N_939 ;
wire N_3_0 ;
wire N_971 ;
wire N_13 ;
wire un1_cf ;
wire N_1688 ;
wire reg3_1_sqmuxa ;
wire un1_df_16 ;
wire N_1750 ;
wire reg3_14_sqmuxa ;
wire N_1812 ;
wire N_1810 ;
wire N_1841 ;
wire N_1661 ;
wire N_1816 ;
wire N_1681 ;
wire N_1743 ;
wire N_938 ;
wire N_970 ;
wire N_1033 ;
wire N_513_i ;
wire N_3873_2 ;
wire N_512_i ;
wire un1_df_1 ;
wire un36_df ;
wire d_cnst_sm0 ;
wire N_3913 ;
wire N_1342 ;
wire N_1374 ;
wire N_514_i ;
wire N_1566 ;
wire N_1584 ;
wire N_1890 ;
wire un86_df ;
wire N_1664 ;
wire N_1819 ;
wire N_1682 ;
wire N_1837 ;
wire N_527_i ;
wire N_1042 ;
wire N_3916 ;
wire N_1270 ;
wire N_1132 ;
wire N_1892 ;
wire N_2641 ;
wire un87_df ;
wire N_7_i ;
wire N_1043 ;
wire b_2_sqmuxa ;
wire N_3912 ;
wire N_895 ;
wire N_526_i ;
wire un1_df_17_2 ;
wire N_1493 ;
wire N_1337 ;
wire N_1343 ;
wire N_1369 ;
wire N_1375 ;
wire N_1561 ;
wire N_1567 ;
wire N_934 ;
wire N_2722 ;
wire N_45 ;
wire N_54 ;
wire m7 ;
wire N_1901 ;
wire addr_4_sqmuxa_1_1 ;
wire un1_b57 ;
wire rd_4_sqmuxa ;
wire N_1740 ;
wire N_2240_i ;
wire N_3568 ;
wire N_2660_2 ;
wire N_915 ;
wire N_919 ;
wire N_918 ;
wire N_1076 ;
wire N_1044 ;
wire N_953 ;
wire N_921 ;
wire N_959 ;
wire N_927 ;
wire N_969 ;
wire N_937 ;
wire N_1084 ;
wire N_1052 ;
wire N_965 ;
wire N_933 ;
wire N_1741 ;
wire N_1679 ;
wire N_1742 ;
wire N_1680 ;
wire N_3614 ;
wire N_974 ;
wire N_942 ;
wire N_1838 ;
wire N_1683 ;
wire N_1039 ;
wire N_1085 ;
wire N_1053 ;
wire N_1083 ;
wire N_1051 ;
wire N_1040 ;
wire N_1038 ;
wire N_952 ;
wire N_920 ;
wire N_1077 ;
wire N_1045 ;
wire N_1081 ;
wire N_1049 ;
wire N_1827 ;
wire N_1672 ;
wire N_1082 ;
wire N_1050 ;
wire N_964 ;
wire N_932 ;
wire N_962 ;
wire N_930 ;
wire N_967 ;
wire N_935 ;
wire N_1079 ;
wire N_1047 ;
wire N_1068 ;
wire N_1036 ;
wire N_1078 ;
wire N_1046 ;
wire N_968 ;
wire N_936 ;
wire N_1069 ;
wire N_1037 ;
wire N_916 ;
wire N_1080 ;
wire N_1048 ;
wire N_1815 ;
wire N_1660 ;
wire N_1820 ;
wire N_1818 ;
wire N_1814 ;
wire N_1665 ;
wire N_1663 ;
wire N_1659 ;
wire N_1752 ;
wire N_1690 ;
wire N_955 ;
wire N_923 ;
wire N_954 ;
wire N_922 ;
wire N_1823 ;
wire N_1668 ;
wire N_956 ;
wire N_924 ;
wire N_1822 ;
wire N_1667 ;
wire N_957 ;
wire N_925 ;
wire N_1829 ;
wire N_1824 ;
wire N_1674 ;
wire N_1669 ;
wire N_961 ;
wire N_929 ;
wire N_1817 ;
wire N_1662 ;
wire N_963 ;
wire N_931 ;
wire N_1830 ;
wire N_1826 ;
wire N_1675 ;
wire N_1671 ;
wire N_960 ;
wire N_928 ;
wire N_1832 ;
wire N_1677 ;
wire N_1831 ;
wire N_1821 ;
wire N_1676 ;
wire N_1666 ;
wire N_1041 ;
wire N_1828 ;
wire N_1673 ;
wire N_972 ;
wire N_940 ;
wire N_1840 ;
wire N_1685 ;
wire N_975 ;
wire N_943 ;
wire N_1839 ;
wire N_1684 ;
wire N_973 ;
wire N_941 ;
wire N_958 ;
wire N_926 ;
wire un1_b59 ;
wire N_1813 ;
wire N_1732 ;
wire N_1670 ;
wire N_1658 ;
wire N_1751 ;
wire N_1689 ;
wire N_1583 ;
wire N_1582 ;
wire N_1581 ;
wire N_1580 ;
wire N_1575 ;
wire N_1574 ;
wire N_1573 ;
wire N_1572 ;
wire N_1571 ;
wire N_1570 ;
wire N_1569 ;
wire N_1568 ;
wire N_1565 ;
wire N_1564 ;
wire N_1563 ;
wire N_1562 ;
wire N_1560 ;
wire N_1035 ;
wire N_1363 ;
wire N_1362 ;
wire N_1361 ;
wire N_1354 ;
wire N_1353 ;
wire N_1352 ;
wire N_1351 ;
wire N_1383 ;
wire N_1350 ;
wire N_1382 ;
wire N_1349 ;
wire N_1381 ;
wire N_1348 ;
wire N_1380 ;
wire N_1347 ;
wire N_1379 ;
wire N_1346 ;
wire N_1378 ;
wire N_1345 ;
wire N_1377 ;
wire N_1344 ;
wire N_1376 ;
wire N_1341 ;
wire N_1373 ;
wire N_1340 ;
wire N_1372 ;
wire N_1339 ;
wire N_1371 ;
wire N_1338 ;
wire N_1370 ;
wire N_1336 ;
wire N_1368 ;
wire N_1335 ;
wire inf_abs0_2_axb_0 ;
wire inf_abs0_2_cry_0 ;
wire inf_abs0_2_axb_1 ;
wire inf_abs0_2_cry_1 ;
wire inf_abs0_2_axb_2 ;
wire inf_abs0_2_cry_2 ;
wire inf_abs0_2_axb_3 ;
wire inf_abs0_2_cry_3 ;
wire inf_abs0_2_axb_4 ;
wire inf_abs0_2_cry_4 ;
wire inf_abs0_2_axb_5 ;
wire inf_abs0_2_cry_5 ;
wire inf_abs0_2_axb_6 ;
wire inf_abs0_2_cry_6 ;
wire inf_abs0_2_axb_7 ;
wire inf_abs0_2_cry_7 ;
wire inf_abs0_2_axb_8 ;
wire inf_abs0_2_cry_8 ;
wire inf_abs0_2_axb_9 ;
wire inf_abs0_2_cry_9 ;
wire inf_abs0_2_axb_10 ;
wire inf_abs0_2_cry_10 ;
wire inf_abs0_2_axb_11 ;
wire inf_abs0_2_cry_11 ;
wire inf_abs0_2_axb_12 ;
wire inf_abs0_2_cry_12 ;
wire inf_abs0_2_axb_13 ;
wire inf_abs0_2_cry_13 ;
wire inf_abs0_2_axb_14 ;
wire inf_abs0_2_cry_14 ;
wire inf_abs0_2_axb_15 ;
wire inf_abs0_2_cry_15 ;
wire inf_abs0_2_axb_16 ;
wire inf_abs0_2_cry_16 ;
wire inf_abs0_2_axb_17 ;
wire inf_abs0_2_cry_17 ;
wire inf_abs0_2_axb_18 ;
wire inf_abs0_2_cry_18 ;
wire inf_abs0_2_axb_19 ;
wire inf_abs0_2_cry_19 ;
wire inf_abs0_2_axb_20 ;
wire inf_abs0_2_cry_20 ;
wire inf_abs0_2_axb_21 ;
wire inf_abs0_2_cry_21 ;
wire inf_abs0_2_axb_22 ;
wire inf_abs0_2_cry_22 ;
wire inf_abs0_2_axb_23 ;
wire inf_abs0_2_cry_23 ;
wire inf_abs0_2_axb_24 ;
wire inf_abs0_2_cry_24 ;
wire inf_abs0_2_axb_25 ;
wire inf_abs0_2_cry_25 ;
wire inf_abs0_2_axb_26 ;
wire inf_abs0_2_cry_26 ;
wire inf_abs0_2_axb_27 ;
wire inf_abs0_2_cry_27 ;
wire inf_abs0_2_axb_28 ;
wire inf_abs0_2_cry_28 ;
wire inf_abs0_2_axb_29 ;
wire inf_abs0_2_cry_29 ;
wire inf_abs0_2_axb_30 ;
wire reg3_1_1_axb_0 ;
wire reg3_1_1_cry_0 ;
wire reg3_1_1_axb_1 ;
wire reg3_1_1_cry_1 ;
wire reg3_1_1_axb_2 ;
wire reg3_1_1_cry_2 ;
wire reg3_1_1_axb_3 ;
wire reg3_1_1_cry_3 ;
wire reg3_1_1_axb_4 ;
wire reg3_1_1_cry_4 ;
wire reg3_1_1_axb_5 ;
wire reg3_1_1_cry_5 ;
wire reg3_1_1_axb_6 ;
wire reg3_1_1_cry_6 ;
wire reg3_1_1_axb_7 ;
wire reg3_1_1_cry_7 ;
wire reg3_1_1_axb_8 ;
wire reg3_1_1_cry_8 ;
wire reg3_1_1_axb_9 ;
wire reg3_1_1_cry_9 ;
wire reg3_1_1_axb_10 ;
wire reg3_1_1_cry_10 ;
wire reg3_1_1_axb_11 ;
wire reg3_1_1_cry_11 ;
wire reg3_1_1_axb_12 ;
wire reg3_1_1_cry_12 ;
wire reg3_1_1_axb_13 ;
wire reg3_1_1_cry_13 ;
wire reg3_1_1_axb_14 ;
wire reg3_1_1_cry_14 ;
wire reg3_1_1_axb_15 ;
wire reg3_1_1_cry_15 ;
wire reg3_1_1_axb_16 ;
wire reg3_1_1_cry_16 ;
wire reg3_1_1_axb_17 ;
wire reg3_1_1_cry_17 ;
wire reg3_1_1_axb_18 ;
wire reg3_1_1_cry_18 ;
wire reg3_1_1_axb_19 ;
wire reg3_1_1_cry_19 ;
wire reg3_1_1_cry_20 ;
wire reg3_1_1_cry_21 ;
wire reg3_1_1_cry_22 ;
wire reg3_1_1_cry_23 ;
wire reg3_1_1_cry_24 ;
wire reg3_1_1_cry_25 ;
wire reg3_1_1_cry_26 ;
wire reg3_1_1_cry_27 ;
wire reg3_1_1_cry_28 ;
wire reg3_1_1_axb_29 ;
wire reg3_1_1_cry_29 ;
wire reg3_1_1_axb_30 ;
wire reg3_1_1_cry_30 ;
wire reg3_1_1_axb_31 ;
wire un3_t_s_1 ;
wire un3_t_s_2 ;
wire un3_t_s_3 ;
wire un3_t_s_4 ;
wire un3_t_s_5 ;
wire un3_t_s_6 ;
wire un3_t_s_7 ;
wire un3_t_s_8 ;
wire un3_t_s_9 ;
wire un3_t_s_10 ;
wire un3_t_s_11 ;
wire un3_t_s_12 ;
wire un3_t_s_13 ;
wire un3_t_s_14 ;
wire un3_t_s_15 ;
wire un3_t_s_16 ;
wire un3_t_s_17 ;
wire un3_t_s_18 ;
wire un3_t_s_19 ;
wire un3_t_s_20 ;
wire un3_t_s_21 ;
wire un3_t_s_22 ;
wire un3_t_s_23 ;
wire un3_t_s_24 ;
wire un3_t_s_25 ;
wire un3_t_s_26 ;
wire un3_t_s_27 ;
wire un3_t_s_28 ;
wire un3_t_s_29 ;
wire un3_t_s_30 ;
wire un3_t_s_31 ;
wire un3_t_cry_0 ;
wire un3_t_cry_1 ;
wire un3_t_axb_2 ;
wire un3_t_cry_2 ;
wire un3_t_cry_3 ;
wire un3_t_cry_4 ;
wire un3_t_cry_5 ;
wire un3_t_cry_6 ;
wire un3_t_cry_7 ;
wire un3_t_cry_8 ;
wire un3_t_cry_9 ;
wire un3_t_cry_10 ;
wire un3_t_cry_11 ;
wire un3_t_cry_12 ;
wire un3_t_cry_13 ;
wire un3_t_cry_14 ;
wire un3_t_cry_15 ;
wire un3_t_cry_16 ;
wire un3_t_cry_17 ;
wire un3_t_cry_18 ;
wire un3_t_cry_19 ;
wire un3_t_cry_20 ;
wire un3_t_cry_21 ;
wire un3_t_cry_22 ;
wire un3_t_cry_23 ;
wire un3_t_cry_24 ;
wire un3_t_cry_25 ;
wire un3_t_cry_26 ;
wire un3_t_cry_27 ;
wire un3_t_cry_28 ;
wire un3_t_axb_29 ;
wire un3_t_cry_29 ;
wire un3_t_axb_30 ;
wire un3_t_cry_30 ;
wire un3_t_axb_31 ;
wire un11_reg0_axb_0 ;
wire un11_reg0_cry_0 ;
wire un11_reg0_axb_1 ;
wire un11_reg0_cry_1 ;
wire un11_reg0_axb_2 ;
wire un11_reg0_cry_2 ;
wire un11_reg0_axb_3 ;
wire un11_reg0_cry_3 ;
wire un11_reg0_axb_4 ;
wire un11_reg0_cry_4 ;
wire un11_reg0_axb_5 ;
wire un11_reg0_cry_5 ;
wire un11_reg0_axb_6 ;
wire un11_reg0_cry_6 ;
wire un11_reg0_axb_7 ;
wire un11_reg0_cry_7 ;
wire un11_reg0_axb_8 ;
wire un11_reg0_cry_8 ;
wire un11_reg0_axb_9 ;
wire un11_reg0_cry_9 ;
wire un11_reg0_axb_10 ;
wire un11_reg0_cry_10 ;
wire un11_reg0_axb_11 ;
wire un11_reg0_cry_11 ;
wire un11_reg0_axb_12 ;
wire un11_reg0_cry_12 ;
wire un11_reg0_axb_13 ;
wire un11_reg0_cry_13 ;
wire un11_reg0_axb_14 ;
wire un11_reg0_cry_14 ;
wire un11_reg0_axb_15 ;
wire un11_reg0_cry_15 ;
wire un11_reg0_axb_16 ;
wire un11_reg0_cry_16 ;
wire un11_reg0_axb_17 ;
wire un11_reg0_cry_17 ;
wire un11_reg0_axb_18 ;
wire un11_reg0_cry_18 ;
wire un11_reg0_axb_19 ;
wire un11_reg0_cry_19 ;
wire un11_reg0_axb_20 ;
wire un11_reg0_cry_20 ;
wire un11_reg0_axb_21 ;
wire un11_reg0_cry_21 ;
wire un11_reg0_axb_22 ;
wire un11_reg0_cry_22 ;
wire un11_reg0_axb_23 ;
wire un11_reg0_cry_23 ;
wire un11_reg0_axb_24 ;
wire un11_reg0_cry_24 ;
wire un11_reg0_axb_25 ;
wire un11_reg0_cry_25 ;
wire un11_reg0_axb_26 ;
wire un11_reg0_cry_26 ;
wire un11_reg0_axb_27 ;
wire un11_reg0_cry_27 ;
wire un11_reg0_axb_28 ;
wire un11_reg0_cry_28 ;
wire un11_reg0_axb_29 ;
wire un32_reg0_s_1 ;
wire un32_reg0_s_2 ;
wire un32_reg0_s_3 ;
wire un32_reg0_s_4 ;
wire un32_reg0_s_5 ;
wire un32_reg0_s_6 ;
wire un32_reg0_s_7 ;
wire un32_reg0_s_8 ;
wire un32_reg0_s_9 ;
wire un32_reg0_s_10 ;
wire un32_reg0_s_11 ;
wire un32_reg0_s_12 ;
wire un32_reg0_s_13 ;
wire un32_reg0_s_14 ;
wire un32_reg0_s_15 ;
wire un32_reg0_s_16 ;
wire un32_reg0_s_17 ;
wire un32_reg0_s_18 ;
wire un32_reg0_s_19 ;
wire un32_reg0_s_20 ;
wire un32_reg0_s_21 ;
wire un32_reg0_s_22 ;
wire un32_reg0_s_23 ;
wire un32_reg0_s_24 ;
wire un32_reg0_s_25 ;
wire un32_reg0_s_26 ;
wire un32_reg0_s_27 ;
wire un32_reg0_s_28 ;
wire un32_reg0_s_29 ;
wire un32_reg0_cry_0 ;
wire un32_reg0_axb_1 ;
wire un32_reg0_cry_1 ;
wire un32_reg0_axb_2 ;
wire un32_reg0_cry_2 ;
wire un32_reg0_axb_3 ;
wire un32_reg0_cry_3 ;
wire un32_reg0_axb_4 ;
wire un32_reg0_cry_4 ;
wire un32_reg0_axb_5 ;
wire un32_reg0_cry_5 ;
wire un32_reg0_axb_6 ;
wire un32_reg0_cry_6 ;
wire un32_reg0_axb_7 ;
wire un32_reg0_cry_7 ;
wire un32_reg0_axb_8 ;
wire un32_reg0_cry_8 ;
wire un32_reg0_axb_9 ;
wire un32_reg0_cry_9 ;
wire un32_reg0_axb_10 ;
wire un32_reg0_cry_10 ;
wire un32_reg0_axb_11 ;
wire un32_reg0_cry_11 ;
wire un32_reg0_axb_12 ;
wire un32_reg0_cry_12 ;
wire un32_reg0_axb_13 ;
wire un32_reg0_cry_13 ;
wire un32_reg0_axb_14 ;
wire un32_reg0_cry_14 ;
wire un32_reg0_axb_15 ;
wire un32_reg0_cry_15 ;
wire un32_reg0_axb_16 ;
wire un32_reg0_cry_16 ;
wire un32_reg0_axb_17 ;
wire un32_reg0_cry_17 ;
wire un32_reg0_axb_18 ;
wire un32_reg0_cry_18 ;
wire un32_reg0_axb_19 ;
wire un32_reg0_cry_19 ;
wire un32_reg0_axb_20 ;
wire un32_reg0_cry_20 ;
wire un32_reg0_axb_21 ;
wire un32_reg0_cry_21 ;
wire un32_reg0_axb_22 ;
wire un32_reg0_cry_22 ;
wire un32_reg0_axb_23 ;
wire un32_reg0_cry_23 ;
wire un32_reg0_axb_24 ;
wire un32_reg0_cry_24 ;
wire un32_reg0_axb_25 ;
wire un32_reg0_cry_25 ;
wire un32_reg0_axb_26 ;
wire un32_reg0_cry_26 ;
wire un32_reg0_axb_27 ;
wire un32_reg0_cry_27 ;
wire un32_reg0_axb_28 ;
wire un32_reg0_cry_28 ;
wire un32_reg0_axb_29 ;
wire un1_inf_abs0_cry_0 ;
wire un1_inf_abs0_axb_1 ;
wire un1_inf_abs0_cry_1 ;
wire un1_inf_abs0_axb_2 ;
wire un1_inf_abs0_cry_2 ;
wire un1_inf_abs0_axb_3 ;
wire un1_inf_abs0_cry_3 ;
wire un1_inf_abs0_axb_4 ;
wire un1_inf_abs0_cry_4 ;
wire un1_inf_abs0_axb_5 ;
wire un1_inf_abs0_cry_5 ;
wire un1_inf_abs0_axb_6 ;
wire un1_inf_abs0_cry_6 ;
wire un1_inf_abs0_axb_7 ;
wire un1_inf_abs0_cry_7 ;
wire un1_inf_abs0_axb_8 ;
wire un1_inf_abs0_cry_8 ;
wire un1_inf_abs0_axb_9 ;
wire un1_inf_abs0_cry_9 ;
wire un1_inf_abs0_axb_10 ;
wire un1_inf_abs0_cry_10 ;
wire un1_inf_abs0_axb_11 ;
wire un1_inf_abs0_cry_11 ;
wire un1_inf_abs0_axb_12 ;
wire un1_inf_abs0_cry_12 ;
wire un1_inf_abs0_axb_13 ;
wire un1_inf_abs0_cry_13 ;
wire un1_inf_abs0_axb_14 ;
wire un1_inf_abs0_cry_14 ;
wire un1_inf_abs0_axb_15 ;
wire un1_inf_abs0_cry_15 ;
wire un1_inf_abs0_axb_16 ;
wire un1_inf_abs0_cry_16 ;
wire un1_inf_abs0_axb_17 ;
wire un1_inf_abs0_cry_17 ;
wire un1_inf_abs0_axb_18 ;
wire un1_inf_abs0_cry_18 ;
wire un1_inf_abs0_axb_19 ;
wire un1_inf_abs0_0_cry_0 ;
wire un1_inf_abs0_0_axb_1 ;
wire un1_inf_abs0_0_cry_1 ;
wire un1_inf_abs0_0_axb_2 ;
wire un1_inf_abs0_0_cry_2 ;
wire un1_inf_abs0_0_axb_3 ;
wire un1_inf_abs0_0_cry_3 ;
wire un1_inf_abs0_0_axb_4 ;
wire un1_inf_abs0_0_cry_4 ;
wire un1_inf_abs0_0_axb_5 ;
wire un1_inf_abs0_0_cry_5 ;
wire un1_inf_abs0_0_axb_6 ;
wire un1_inf_abs0_0_cry_6 ;
wire un1_inf_abs0_0_axb_7 ;
wire un1_inf_abs0_0_cry_7 ;
wire un1_inf_abs0_0_axb_8 ;
wire un1_inf_abs0_0_cry_8 ;
wire un1_inf_abs0_0_axb_9 ;
wire un1_inf_abs0_0_cry_9 ;
wire un1_inf_abs0_0_axb_10 ;
wire un1_inf_abs0_0_cry_10 ;
wire un1_inf_abs0_0_axb_11 ;
wire un1_inf_abs0_0_cry_11 ;
wire un1_inf_abs0_0_axb_12 ;
wire un1_inf_abs0_0_cry_12 ;
wire un1_inf_abs0_0_axb_13 ;
wire un1_inf_abs0_0_cry_13 ;
wire un1_inf_abs0_0_axb_14 ;
wire un1_inf_abs0_0_cry_14 ;
wire un1_inf_abs0_0_axb_15 ;
wire un1_inf_abs0_0_cry_15 ;
wire un1_inf_abs0_0_axb_16 ;
wire un1_inf_abs0_0_cry_16 ;
wire un1_inf_abs0_0_axb_17 ;
wire un1_inf_abs0_0_cry_17 ;
wire un1_inf_abs0_0_axb_18 ;
wire un1_inf_abs0_0_cry_18 ;
wire un1_inf_abs0_0_axb_19 ;
wire un3_reg3_s_1 ;
wire un3_reg3_s_2 ;
wire un3_reg3_s_3 ;
wire un3_reg3_s_4 ;
wire un3_reg3_s_5 ;
wire un3_reg3_s_6 ;
wire un3_reg3_s_7 ;
wire un3_reg3_s_8 ;
wire un3_reg3_s_9 ;
wire un3_reg3_s_10 ;
wire un3_reg3_s_11 ;
wire un3_reg3_s_12 ;
wire un3_reg3_s_13 ;
wire un3_reg3_s_14 ;
wire un3_reg3_s_15 ;
wire un3_reg3_s_16 ;
wire un3_reg3_s_17 ;
wire un3_reg3_s_18 ;
wire un3_reg3_s_19 ;
wire un3_reg3_s_20 ;
wire un3_reg3_s_21 ;
wire un3_reg3_s_22 ;
wire un3_reg3_s_23 ;
wire un3_reg3_s_24 ;
wire un3_reg3_s_25 ;
wire un3_reg3_cry_25 ;
wire un3_reg3_axb_1 ;
wire un3_reg3_cry_1 ;
wire un3_reg3_axb_2 ;
wire un3_reg3_cry_2 ;
wire un3_reg3_axb_3 ;
wire un3_reg3_cry_3 ;
wire un3_reg3_axb_4 ;
wire un3_reg3_cry_4 ;
wire un3_reg3_axb_5 ;
wire un3_reg3_cry_5 ;
wire un3_reg3_axb_6 ;
wire un3_reg3_cry_6 ;
wire un3_reg3_axb_7 ;
wire un3_reg3_cry_7 ;
wire un3_reg3_axb_8 ;
wire un3_reg3_cry_8 ;
wire un3_reg3_axb_9 ;
wire un3_reg3_cry_9 ;
wire un3_reg3_axb_10 ;
wire un3_reg3_cry_10 ;
wire un3_reg3_axb_11 ;
wire un3_reg3_cry_11 ;
wire un3_reg3_axb_12 ;
wire un3_reg3_cry_12 ;
wire un3_reg3_axb_13 ;
wire un3_reg3_cry_13 ;
wire un3_reg3_axb_14 ;
wire un3_reg3_cry_14 ;
wire un3_reg3_axb_15 ;
wire un3_reg3_cry_15 ;
wire un3_reg3_axb_16 ;
wire un3_reg3_cry_16 ;
wire un3_reg3_axb_17 ;
wire un3_reg3_cry_17 ;
wire un3_reg3_axb_18 ;
wire un3_reg3_cry_18 ;
wire un3_reg3_axb_19 ;
wire un3_reg3_cry_19 ;
wire un3_reg3_axb_20 ;
wire un3_reg3_cry_20 ;
wire un3_reg3_axb_21 ;
wire un3_reg3_cry_21 ;
wire un3_reg3_axb_22 ;
wire un3_reg3_cry_22 ;
wire un3_reg3_axb_23 ;
wire un3_reg3_cry_23 ;
wire un3_reg3_axb_24 ;
wire un3_reg3_cry_24 ;
wire un3_reg3_axb_25 ;
wire t_1_cry_0 ;
wire t_1_cry_1 ;
wire t_1_cry_2 ;
wire t_1_cry_3 ;
wire t_1_cry_4 ;
wire t_1_cry_5 ;
wire t_1_cry_6 ;
wire t_1_cry_7 ;
wire t_1_cry_8 ;
wire t_1_cry_9 ;
wire t_1_cry_10 ;
wire t_1_cry_11 ;
wire t_1_cry_12 ;
wire t_1_cry_13 ;
wire t_1_cry_14 ;
wire t_1_cry_15 ;
wire t_1_cry_16 ;
wire t_1_cry_17 ;
wire t_1_cry_18 ;
wire t_1_cry_19 ;
wire t_1_cry_20 ;
wire t_1_cry_21 ;
wire t_1_cry_22 ;
wire t_1_cry_23 ;
wire t_1_cry_24 ;
wire t_1_cry_25 ;
wire t_1_cry_26 ;
wire t_1_cry_27 ;
wire t_1_cry_28 ;
wire t_1_cry_29 ;
wire t_1_cry_30 ;
wire \d_cnst_sn.reg1_16_8_1837_2_tz  ;
wire reg0_28_sn_m6_lut6_2_O5 ;
wire \d_cnst_sn.reg3_17_sn_m7_0  ;
wire reg3_1_sqmuxa_RNIH1DM1 ;
wire reg3_1_sqmuxa_RNIE1DM1 ;
wire reg3_1_sqmuxa_RNIQMUH1 ;
wire reg3_1_sqmuxa_RNITMUH1 ;
wire reg3_1_sqmuxa_RNIKMUH1 ;
wire reg3_1_sqmuxa_RNINMUH1 ;
wire reg3_1_sqmuxa_RNIHMUH1 ;
wire reg3_1_sqmuxa_RNIEMUH1 ;
wire reg0_m9_i_a1 ;
wire \d_cnst_sn.reg2_N_3_mux  ;
wire g0_2_0_i2_lut6_2_O6 ;
wire reg3_N_7_i_RNO ;
wire \d_cnst_sn.reg1_16_9_1804_3_tz  ;
wire \d_cnst_sn.addr_20_iv_1052_i_a6_1_0  ;
wire \d_cnst_sn.reg0_m8_e_0  ;
wire \d_cnst_sn.reg3_5_sqmuxa_2_1  ;
wire \d_cnst_sn.reg0_28_9_2294_a6_3_0  ;
wire N_3910 ;
wire \d_cnst_sn.un1_state_3_1  ;
wire \d_cnst_sn.b60_0  ;
wire \d_cnst_sn.b64_0  ;
wire \d_cnst_sn.reg0_m9_i_a3_0  ;
wire reg3_17_sn_N_5 ;
wire \d_cnst_sn.reg0_28_2526_a5_1_0  ;
wire N_4571_i ;
wire N_4570_i ;
wire N_4569_i ;
wire N_4568_i ;
wire N_4567_i ;
wire N_4566_i ;
wire N_4565_i ;
wire N_4564_i ;
wire N_4563_i ;
wire N_4562_i ;
wire N_4561_i ;
wire N_4560_i ;
wire N_4559_i ;
wire N_4558_i ;
wire N_4557_i ;
wire N_4556_i ;
wire N_4555_i ;
wire N_4554_i ;
wire N_4553_i ;
wire N_4552_i ;
wire N_4551_i ;
wire N_4550_i ;
wire N_4549_i ;
wire N_4548_i ;
wire N_4547_i ;
wire N_4546_i ;
wire N_4545_i ;
wire N_4544_i ;
wire N_4543_i ;
wire N_4542_i ;
wire N_4541_i ;
wire \d_cnst_sn.reg3_N_7_i  ;
wire N_2099_i ;
wire addr_0_sqmuxa_1_i ;
wire N_2119_i ;
wire N_2139_i ;
wire N_2159_i ;
wire N_2179_i ;
wire N_2199_i ;
wire N_2219_i ;
wire N_56_i ;
wire N_2267_i ;
wire N_47_i ;
wire N_2315_i ;
wire N_2335_i ;
wire N_36_i ;
wire N_2516_i ;
wire N_2536_i ;
wire N_2556_i ;
wire N_2576_i ;
wire N_2596_i ;
wire N_2616_i ;
wire N_2636_i ;
wire N_2656_i ;
wire un1_state_1_0_i ;
wire un1_state_3_i ;
wire un1_state_4_i ;
wire \d_cnst_sn.addr_20_iv_1052_i_a6_2_0  ;
wire \d_cnst_sn.m26_0_1  ;
wire \d_cnst_sn.m19_0_1  ;
wire \d_cnst_sn.addr_20_iv_7_654_i_1  ;
wire \d_cnst_sn.addr_20_iv_8_627_i_1  ;
wire \d_cnst_sn.addr_20_iv_16_389_i_1  ;
wire \d_cnst_sn.addr_20_iv_12_497_i_1  ;
wire \d_cnst_sn.addr_20_iv_10_562_i_1  ;
wire \d_cnst_sn.addr_20_iv_14_443_i_2  ;
wire \d_cnst_sn.addr_20_iv_15_416_i_1  ;
wire \d_cnst_sn.addr_20_iv_17_362_i_1  ;
wire \d_cnst_sn.addr_20_iv_13_470_i_1  ;
wire \d_cnst_sn.addr_20_iv_18_335_i_1  ;
wire \d_cnst_sn.addr_20_iv_2_971_i_0  ;
wire \d_cnst_sn.addr_20_iv_1_998_i_0  ;
wire \d_cnst_sn.addr_20_iv_1052_i_0  ;
wire \d_cnst_sn.addr_20_iv_0_1025_i_0  ;
wire \d_cnst_sn.addr_20_iv_3_944_i_0  ;
wire \d_cnst_sn.addr_20_iv_4_917_i_0  ;
wire \d_cnst_sn.addr_20_iv_5_890_i_0  ;
wire \d_cnst_sn.addr_20_iv_6_863_i_0  ;
wire \d_cnst_sn.reg0_28_12_2195_a6_1_2_0  ;
wire \d_cnst_sn.reg0_m9_i_a0_0  ;
wire \d_cnst_sn.reg0_28_5_2426_a6_1_1  ;
wire \d_cnst_sn.reg0_28_5_2426_3_1  ;
wire \d_cnst_sn.reg0_28_8_2327_a6_1_1  ;
wire \d_cnst_sn.reg0_28_6_2393_3_1  ;
wire \d_cnst_sn.reg0_28_6_2393_a6_1_1  ;
wire \d_cnst_sn.reg0_28_7_2360_3_1  ;
wire \d_cnst_sn.reg0_28_7_2360_a6_1_1  ;
wire \d_cnst_sn.reg0_28_14_2135_1_a0_2  ;
wire \d_cnst_sn.reg0_28_9_2294_a6_1_1  ;
wire \d_cnst_sn.reg0_28_9_2294_3_1  ;
wire \d_cnst_sn.reg1_16_7_1870_3_1  ;
wire \d_cnst_sn.reg0_28_10_2261_a6_1_1  ;
wire \d_cnst_sn.reg1_16_8_1837_3_1  ;
wire \d_cnst_sn.reg0_28_11_2228_a6_1_1  ;
wire \d_cnst_sn.reg0_28_3_2492_0  ;
wire \d_cnst_sn.reg0_28_3_2492_1  ;
wire \d_cnst_sn.reg0_28_4_2459_0  ;
wire \d_cnst_sn.reg0_28_8_2327_0  ;
wire \d_cnst_sn.reg0_28_5_2426_0  ;
wire \d_cnst_sn.reg0_28_6_2393_0  ;
wire \d_cnst_sn.reg0_28_7_2360_0  ;
wire \d_cnst_sn.reg0_28_14_0  ;
wire \d_cnst_sn.reg0_28_9_2294_0  ;
wire \d_cnst_sn.reg1_16_7_1870_0  ;
wire \d_cnst_sn.reg1_16_8_1837_0  ;
wire b_0 ;
wire un3_t_axb_28 ;
wire un3_t_axb_27 ;
wire un3_t_axb_26 ;
wire un3_t_axb_25 ;
wire un3_t_axb_24 ;
wire un3_t_axb_23 ;
wire un3_t_axb_22 ;
wire un3_t_axb_21 ;
wire un3_t_axb_20 ;
wire un3_t_axb_19 ;
wire un3_t_axb_18 ;
wire un3_t_axb_17 ;
wire un3_t_axb_16 ;
wire un3_t_axb_15 ;
wire un3_t_axb_14 ;
wire un3_t_axb_13 ;
wire un3_t_axb_12 ;
wire un3_t_axb_11 ;
wire un3_t_axb_10 ;
wire un3_t_axb_9 ;
wire un3_t_axb_8 ;
wire un3_t_axb_7 ;
wire un3_t_axb_6 ;
wire un3_t_axb_5 ;
wire un3_t_axb_4 ;
wire un3_t_axb_3 ;
wire un3_t_axb_1 ;
wire un3_t_axb_0 ;
wire reg3_1_1_axb_28 ;
wire reg3_1_1_axb_27 ;
wire reg3_1_1_axb_26 ;
wire reg3_1_1_axb_25 ;
wire reg3_1_1_axb_24 ;
wire reg3_1_1_axb_23 ;
wire reg3_1_1_axb_22 ;
wire reg3_1_1_axb_21 ;
wire reg3_1_1_axb_20 ;
wire t_1_cry_0_cy ;
wire un3_t_cry_0_cy ;
wire N_7 ;
wire N_12 ;
wire \d_cnst_sn.g0_3_a2_2  ;
wire \d_cnst_sn.g0_3_1  ;
wire \d_cnst_sn.g3  ;
wire \d_cnst_sn.reg0_N_13_0  ;
wire \d_cnst_sn.g0_0_2  ;
wire \d_cnst_sn.g0_1  ;
wire N_7_0 ;
wire \d_cnst_sn.g0_0_0_a5_0_0  ;
wire \d_cnst_sn.g0_0_0_a5_2  ;
wire \d_cnst_sn.g0_0_0_1  ;
wire N_3856_rep1 ;
wire N_3569_rep1 ;
wire N_3289_rep1 ;
wire N_3315_rep1 ;
wire N_3550_rep1 ;
wire N_3341_rep1 ;
wire N_3673_rep1 ;
wire N_3699_rep1 ;
wire N_3725_rep1 ;
wire N_3751_rep1 ;
wire N_3777_rep1 ;
wire N_3803_rep1 ;
wire N_3829_rep1 ;
wire \d_cnst_sn.g0_rn_1  ;
wire reg0_28_7_rep1 ;
wire d_cnst_ss0_x ;
wire un1_cf_x ;
wire un3_reg3_cry_25_0 ;
wire un3_reg3_cry_25_1 ;
wire inf_abs0_2_cry_29_0 ;
wire inf_abs0_2_cry_29_1 ;
input p_b_Z_p_O_FDC ;
input p_desc52_p_O_FDC ;
input p_desc53_p_O_FDC ;
input p_desc54_p_O_FDC ;
input p_desc55_p_O_FDC ;
input p_desc56_p_O_FDC ;
input p_desc57_p_O_FDC ;
input p_desc58_p_O_FDC ;
input p_desc59_p_O_FDC ;
input p_desc60_p_O_FDC ;
input p_desc61_p_O_FDC ;
input p_desc62_p_O_FDC ;
input p_desc63_p_O_FDC ;
input p_desc64_p_O_FDC ;
input p_desc65_p_O_FDC ;
input p_desc66_p_O_FDC ;
input p_desc67_p_O_FDC ;
input p_desc68_p_O_FDC ;
input p_desc69_p_O_FDC ;
input p_desc70_p_O_FDC ;
input p_desc71_p_O_FDC ;
input p_desc72_p_O_FDC ;
input p_desc73_p_O_FDC ;
input p_desc74_p_O_FDC ;
input p_desc75_p_O_FDC ;
input p_desc76_p_O_FDC ;
input p_desc77_p_O_FDC ;
input p_desc78_p_O_FDC ;
input p_desc79_p_O_FDC ;
input p_desc80_p_O_FDC ;
input p_desc81_p_O_FDC ;
input p_desc82_p_O_FDC ;
input p_desc83_p_O_FDC ;
input p_rd_Z_p_O_FDC ;
input p_desc261_p_O_FDC ;
input p_wr_Z_p_O_FDC ;
input p_desc262_p_O_FDC ;
input p_desc50_p_O_FDCE ;
input p_desc51_p_O_FDCE ;
input p_desc84_p_O_FDCE ;
input p_desc85_p_O_FDCE ;
input p_desc86_p_O_FDCE ;
input p_desc87_p_O_FDCE ;
input p_desc88_p_O_FDCE ;
input p_desc89_p_O_FDCE ;
input p_desc90_p_O_FDCE ;
input p_desc91_p_O_FDCE ;
input p_desc92_p_O_FDCE ;
input p_desc93_p_O_FDCE ;
input p_desc94_p_O_FDCE ;
input p_desc95_p_O_FDCE ;
input p_desc96_p_O_FDCE ;
input p_desc97_p_O_FDCE ;
input p_desc98_p_O_FDCE ;
input p_desc99_p_O_FDCE ;
input p_desc100_p_O_FDCE ;
input p_desc101_p_O_FDCE ;
input p_desc102_p_O_FDCE ;
input p_desc103_p_O_FDCE ;
input p_desc104_p_O_FDCE ;
input p_desc105_p_O_FDCE ;
input p_desc106_p_O_FDCE ;
input p_desc107_p_O_FDCE ;
input p_desc108_p_O_FDCE ;
input p_desc109_p_O_FDCE ;
input p_desc110_p_O_FDCE ;
input p_desc111_p_O_FDCE ;
input p_desc112_p_O_FDCE ;
input p_desc113_p_O_FDCE ;
input p_desc114_p_O_FDCE ;
input p_desc115_p_O_FDCE ;
input p_desc116_p_O_FDCE ;
input p_desc117_p_O_FDCE ;
input p_desc118_p_O_FDCE ;
input p_desc119_p_O_FDCE ;
input p_desc120_p_O_FDCE ;
input p_desc121_p_O_FDCE ;
input p_desc122_p_O_FDCE ;
input p_desc123_p_O_FDCE ;
input p_desc124_p_O_FDCE ;
input p_desc125_p_O_FDCE ;
input p_desc126_p_O_FDCE ;
input p_desc127_p_O_FDCE ;
input p_desc128_p_O_FDCE ;
input p_desc129_p_O_FDCE ;
input p_desc130_p_O_FDCE ;
input p_desc131_p_O_FDCE ;
input p_desc132_p_O_FDCE ;
input p_desc133_p_O_FDCE ;
input p_desc134_p_O_FDCE ;
input p_desc135_p_O_FDCE ;
input p_desc136_p_O_FDCE ;
input p_desc137_p_O_FDCE ;
input p_desc138_p_O_FDCE ;
input p_desc139_p_O_FDCE ;
input p_desc140_p_O_FDCE ;
input p_desc141_p_O_FDCE ;
input p_desc142_p_O_FDCE ;
input p_desc143_p_O_FDCE ;
input p_desc144_p_O_FDCE ;
input p_desc145_p_O_FDCE ;
input p_desc146_p_O_FDCE ;
input p_desc147_p_O_FDCE ;
input p_desc148_p_O_FDCE ;
input p_desc149_p_O_FDCE ;
input p_desc150_p_O_FDCE ;
input p_desc151_p_O_FDCE ;
input p_desc152_p_O_FDCE ;
input p_desc153_p_O_FDCE ;
input p_desc154_p_O_FDCE ;
input p_desc155_p_O_FDCE ;
input p_desc156_p_O_FDCE ;
input p_desc157_p_O_FDCE ;
input p_desc158_p_O_FDCE ;
input p_desc159_p_O_FDCE ;
input p_desc160_p_O_FDCE ;
input p_desc161_p_O_FDCE ;
input p_desc162_p_O_FDCE ;
input p_desc163_p_O_FDCE ;
input p_desc164_p_O_FDCE ;
input p_desc165_p_O_FDCE ;
input p_desc166_p_O_FDCE ;
input p_desc167_p_O_FDCE ;
input p_desc168_p_O_FDCE ;
input p_desc169_p_O_FDCE ;
input p_desc170_p_O_FDCE ;
input p_desc171_p_O_FDCE ;
input p_desc172_p_O_FDCE ;
input p_desc173_p_O_FDCE ;
input p_desc174_p_O_FDCE ;
input p_desc175_p_O_FDCE ;
input p_desc176_p_O_FDCE ;
input p_desc177_p_O_FDCE ;
input p_desc178_p_O_FDCE ;
input p_desc179_p_O_FDCE ;
input p_desc180_p_O_FDCE ;
input p_desc181_p_O_FDCE ;
input p_desc182_p_O_FDCE ;
input p_desc183_p_O_FDCE ;
input p_desc184_p_O_FDCE ;
input p_desc185_p_O_FDCE ;
input p_desc186_p_O_FDCE ;
input p_desc187_p_O_FDCE ;
input p_desc188_p_O_FDCE ;
input p_desc189_p_O_FDCE ;
input p_desc190_p_O_FDCE ;
input p_desc191_p_O_FDCE ;
input p_desc192_p_O_FDCE ;
input p_desc193_p_O_FDCE ;
input p_desc194_p_O_FDCE ;
input p_desc195_p_O_FDCE ;
input p_desc196_p_O_FDCE ;
input p_desc197_p_O_FDCE ;
input p_desc198_p_O_FDCE ;
input p_desc199_p_O_FDCE ;
input p_desc200_p_O_FDCE ;
input p_desc201_p_O_FDCE ;
input p_desc202_p_O_FDCE ;
input p_desc203_p_O_FDCE ;
input p_desc204_p_O_FDCE ;
input p_desc205_p_O_FDCE ;
input p_desc206_p_O_FDCE ;
input p_desc207_p_O_FDCE ;
input p_desc208_p_O_FDCE ;
input p_desc209_p_O_FDCE ;
input p_desc210_p_O_FDCE ;
input p_desc211_p_O_FDCE ;
input p_desc212_p_O_FDCE ;
input p_desc213_p_O_FDCE ;
input p_desc214_p_O_FDCE ;
input p_desc215_p_O_FDCE ;
input p_desc216_p_O_FDCE ;
input p_desc217_p_O_FDCE ;
input p_desc218_p_O_FDCE ;
input p_desc219_p_O_FDCE ;
input p_desc220_p_O_FDCE ;
input p_desc221_p_O_FDCE ;
input p_desc222_p_O_FDCE ;
input p_desc223_p_O_FDCE ;
input p_desc224_p_O_FDCE ;
input p_desc225_p_O_FDCE ;
input p_desc226_p_O_FDCE ;
input p_desc227_p_O_FDCE ;
input p_desc228_p_O_FDCE ;
input p_desc229_p_O_FDCE ;
input p_desc230_p_O_FDCE ;
input p_desc231_p_O_FDCE ;
input p_desc232_p_O_FDCE ;
input p_desc233_p_O_FDCE ;
input p_desc234_p_O_FDCE ;
input p_desc235_p_O_FDCE ;
input p_desc236_p_O_FDCE ;
input p_desc237_p_O_FDCE ;
input p_desc238_p_O_FDCE ;
input p_desc239_p_O_FDCE ;
input p_desc240_p_O_FDCE ;
input p_desc241_p_O_FDCE ;
input p_desc242_p_O_FDCE ;
input p_desc243_p_O_FDCE ;
input p_desc244_p_O_FDCE ;
input p_desc245_p_O_FDCE ;
input p_desc246_p_O_FDCE ;
input p_desc247_p_O_FDCE ;
input p_desc248_p_O_FDCE ;
input p_desc249_p_O_FDCE ;
input p_desc250_p_O_FDCE ;
input p_desc251_p_O_FDCE ;
input p_desc252_p_O_FDCE ;
input p_desc253_p_O_FDCE ;
input p_desc254_p_O_FDCE ;
input p_desc255_p_O_FDCE ;
input p_desc256_p_O_FDCE ;
input p_desc257_p_O_FDCE ;
input p_desc258_p_O_FDCE ;
input p_desc259_p_O_FDCE ;
input p_desc260_p_O_FDCE ;
// instances
  GND GND_cZ(.G(GND));
  VCC VCC_cZ(.P(VCC));
  MUXF8 desc0(.I0(\d_cnst_sn.reg2_16_11muxnet_0 [1:1]),.I1(\d_cnst_sn.reg2_16_11muxnet_1 [1:1]),.S(N_513_i),.O(reg2_16[1:1]));
  MUXF7 desc1(.I0(N_1560),.I1(t_6[1:1]),.S(N_514_i),.O(\d_cnst_sn.reg2_16_11muxnet_1 [1:1]));
  MUXF7 desc2(.I0(N_1336),.I1(N_1368),.S(N_514_i),.O(\d_cnst_sn.reg2_16_11muxnet_0 [1:1]));
  LUT1 inf_abs0_2_cry_29_outextlut(.I0(VCC),.O(inf_abs0_2_cry_29_1));
defparam inf_abs0_2_cry_29_outextlut.INIT=2'h3;
  LUT1 un3_reg3_cry_25_outextlut(.I0(VCC),.O(un3_reg3_cry_25_1));
defparam un3_reg3_cry_25_outextlut.INIT=2'h3;
  LUT1 inf_abs0_2_cry_30_outextlut(.I0(VCC),.O(inf_abs0_2_1[31:31]));
defparam inf_abs0_2_cry_30_outextlut.INIT=2'h3;
  LUT6_2 desc3(.I0(reg0[30:30]),.I1(reg1[30:30]),.I2(reg2[30:30]),.I3(inf_abs0_2[29:29]),.I4(inf_abs0_2[30:30]),.I5(inf_abs0_2[31:31]),.O6(r_4[30:30]),.O5(r_4_3_lut6_2_O5[30:30]));
defparam desc3.INIT=64'hAAAAAAAA00F0CCAA;
  LUT4 un11_r_df0_cZ(.I0(m_2[0:0]),.I1(m_2[1:1]),.I2(r_4[0:0]),.I3(r_4[1:1]),.O(un11_r_df0));
defparam un11_r_df0_cZ.INIT=16'h8421;
  LUT4 un11_r_df2_cZ(.I0(N_28),.I1(m_2[2:2]),.I2(m_2[3:3]),.I3(r_4[3:3]),.O(un11_r_df2));
defparam un11_r_df2_cZ.INIT=16'h9009;
  LUT4 un11_r_df4_cZ(.I0(m_2[4:4]),.I1(m_2[5:5]),.I2(r_4[4:4]),.I3(r_4[5:5]),.O(un11_r_df4));
defparam un11_r_df4_cZ.INIT=16'h8421;
  LUT4 un11_r_df6_cZ(.I0(m_2[6:6]),.I1(m_2[7:7]),.I2(r_4[6:6]),.I3(r_4[7:7]),.O(un11_r_df6));
defparam un11_r_df6_cZ.INIT=16'h8421;
  LUT4 un11_r_df8_cZ(.I0(m_2[8:8]),.I1(m_2[9:9]),.I2(r_4[8:8]),.I3(r_4[9:9]),.O(un11_r_df8));
defparam un11_r_df8_cZ.INIT=16'h8421;
  LUT4 un11_r_df10_cZ(.I0(m_2[10:10]),.I1(m_2[11:11]),.I2(r_4[10:10]),.I3(r_4[11:11]),.O(un11_r_df10));
defparam un11_r_df10_cZ.INIT=16'h8421;
  LUT4 un11_r_df12_cZ(.I0(m_2[12:12]),.I1(m_2[13:13]),.I2(r_4[12:12]),.I3(r_4[13:13]),.O(un11_r_df12));
defparam un11_r_df12_cZ.INIT=16'h8421;
  LUT4 un11_r_df14_cZ(.I0(m_2[14:14]),.I1(m_2[15:15]),.I2(r_4[14:14]),.I3(r_4[15:15]),.O(un11_r_df14));
defparam un11_r_df14_cZ.INIT=16'h8421;
  LUT4 un11_r_df16_cZ(.I0(m_2[16:16]),.I1(m_2[17:17]),.I2(r_4[16:16]),.I3(r_4[17:17]),.O(un11_r_df16));
defparam un11_r_df16_cZ.INIT=16'h8421;
  LUT4 un11_r_df18_cZ(.I0(m_2[18:18]),.I1(m_2[19:19]),.I2(r_4[18:18]),.I3(r_4[19:19]),.O(un11_r_df18));
defparam un11_r_df18_cZ.INIT=16'h8421;
  LUT4 b18_df0_cZ(.I0(m_2[0:0]),.I1(m_2[1:1]),.I2(r_4[0:0]),.I3(r_4[1:1]),.O(b18_df0));
defparam b18_df0_cZ.INIT=16'h8421;
  LUT4 b18_df2_cZ(.I0(N_28),.I1(m_2[2:2]),.I2(m_2[3:3]),.I3(r_4[3:3]),.O(b18_df2));
defparam b18_df2_cZ.INIT=16'h9009;
  LUT4 b18_df4_cZ(.I0(m_2[4:4]),.I1(m_2[5:5]),.I2(r_4[4:4]),.I3(r_4[5:5]),.O(b18_df4));
defparam b18_df4_cZ.INIT=16'h8421;
  LUT4 b18_df6_cZ(.I0(m_2[6:6]),.I1(m_2[7:7]),.I2(r_4[6:6]),.I3(r_4[7:7]),.O(b18_df6));
defparam b18_df6_cZ.INIT=16'h8421;
  LUT4 b18_df8_cZ(.I0(m_2[8:8]),.I1(m_2[9:9]),.I2(r_4[8:8]),.I3(r_4[9:9]),.O(b18_df8));
defparam b18_df8_cZ.INIT=16'h8421;
  LUT4 b18_df10_cZ(.I0(m_2[10:10]),.I1(m_2[11:11]),.I2(r_4[10:10]),.I3(r_4[11:11]),.O(b18_df10));
defparam b18_df10_cZ.INIT=16'h8421;
  LUT4 b18_df12_cZ(.I0(m_2[12:12]),.I1(m_2[13:13]),.I2(r_4[12:12]),.I3(r_4[13:13]),.O(b18_df12));
defparam b18_df12_cZ.INIT=16'h8421;
  LUT4 b18_df14_cZ(.I0(m_2[14:14]),.I1(m_2[15:15]),.I2(r_4[14:14]),.I3(r_4[15:15]),.O(b18_df14));
defparam b18_df14_cZ.INIT=16'h8421;
  LUT4 b18_df16_cZ(.I0(m_2[16:16]),.I1(m_2[17:17]),.I2(r_4[16:16]),.I3(r_4[17:17]),.O(b18_df16));
defparam b18_df16_cZ.INIT=16'h8421;
  LUT4 b18_df18_cZ(.I0(m_2[18:18]),.I1(m_2[19:19]),.I2(r_4[18:18]),.I3(r_4[19:19]),.O(b18_df18));
defparam b18_df18_cZ.INIT=16'h8421;
  LUT4 un26_r_df0_cZ(.I0(m_2[0:0]),.I1(m_2[1:1]),.I2(r_4[0:0]),.I3(r_4[1:1]),.O(un26_r_df0));
defparam un26_r_df0_cZ.INIT=16'h8421;
  LUT4 un26_r_df2_cZ(.I0(N_28),.I1(m_2[2:2]),.I2(m_2[3:3]),.I3(r_4[3:3]),.O(un26_r_df2));
defparam un26_r_df2_cZ.INIT=16'h9009;
  LUT4 un26_r_df4_cZ(.I0(m_2[4:4]),.I1(m_2[5:5]),.I2(r_4[4:4]),.I3(r_4[5:5]),.O(un26_r_df4));
defparam un26_r_df4_cZ.INIT=16'h8421;
  LUT4 un26_r_df6_cZ(.I0(m_2[6:6]),.I1(m_2[7:7]),.I2(r_4[6:6]),.I3(r_4[7:7]),.O(un26_r_df6));
defparam un26_r_df6_cZ.INIT=16'h8421;
  LUT4 un26_r_df8_cZ(.I0(m_2[8:8]),.I1(m_2[9:9]),.I2(r_4[8:8]),.I3(r_4[9:9]),.O(un26_r_df8));
defparam un26_r_df8_cZ.INIT=16'h8421;
  LUT4 un26_r_df10_cZ(.I0(m_2[10:10]),.I1(m_2[11:11]),.I2(r_4[10:10]),.I3(r_4[11:11]),.O(un26_r_df10));
defparam un26_r_df10_cZ.INIT=16'h8421;
  LUT4 un26_r_df12_cZ(.I0(m_2[12:12]),.I1(m_2[13:13]),.I2(r_4[12:12]),.I3(r_4[13:13]),.O(un26_r_df12));
defparam un26_r_df12_cZ.INIT=16'h8421;
  LUT4 un26_r_df14_cZ(.I0(m_2[14:14]),.I1(m_2[15:15]),.I2(r_4[14:14]),.I3(r_4[15:15]),.O(un26_r_df14));
defparam un26_r_df14_cZ.INIT=16'h8421;
  LUT4 un26_r_df16_cZ(.I0(m_2[16:16]),.I1(m_2[17:17]),.I2(r_4[16:16]),.I3(r_4[17:17]),.O(un26_r_df16));
defparam un26_r_df16_cZ.INIT=16'h8421;
  LUT4 un26_r_df18_cZ(.I0(m_2[18:18]),.I1(m_2[19:19]),.I2(r_4[18:18]),.I3(r_4[19:19]),.O(un26_r_df18));
defparam un26_r_df18_cZ.INIT=16'h8421;
  LUT2 inf_abs0_2_axb_0_cZ(.I0(ir[0:0]),.I1(ir_fast[31:31]),.O(inf_abs0_2_axb_0));
defparam inf_abs0_2_axb_0_cZ.INIT=4'h6;
  LUT2 inf_abs0_2_axb_1_cZ(.I0(ir[1:1]),.I1(ir_fast[31:31]),.O(inf_abs0_2_axb_1));
defparam inf_abs0_2_axb_1_cZ.INIT=4'h6;
  LUT2 inf_abs0_2_axb_2_cZ(.I0(ir[2:2]),.I1(ir_fast[31:31]),.O(inf_abs0_2_axb_2));
defparam inf_abs0_2_axb_2_cZ.INIT=4'h6;
  LUT2 inf_abs0_2_axb_3_cZ(.I0(ir[3:3]),.I1(ir_fast[31:31]),.O(inf_abs0_2_axb_3));
defparam inf_abs0_2_axb_3_cZ.INIT=4'h6;
  LUT2 inf_abs0_2_axb_4_cZ(.I0(ir[4:4]),.I1(ir_fast[31:31]),.O(inf_abs0_2_axb_4));
defparam inf_abs0_2_axb_4_cZ.INIT=4'h6;
  LUT2 inf_abs0_2_axb_5_cZ(.I0(ir[5:5]),.I1(ir_fast[31:31]),.O(inf_abs0_2_axb_5));
defparam inf_abs0_2_axb_5_cZ.INIT=4'h6;
  LUT2 inf_abs0_2_axb_6_cZ(.I0(ir[6:6]),.I1(ir_fast[31:31]),.O(inf_abs0_2_axb_6));
defparam inf_abs0_2_axb_6_cZ.INIT=4'h6;
  LUT2 inf_abs0_2_axb_7_cZ(.I0(ir[7:7]),.I1(ir_fast[31:31]),.O(inf_abs0_2_axb_7));
defparam inf_abs0_2_axb_7_cZ.INIT=4'h6;
  LUT2 inf_abs0_2_axb_8_cZ(.I0(ir[8:8]),.I1(ir_fast[31:31]),.O(inf_abs0_2_axb_8));
defparam inf_abs0_2_axb_8_cZ.INIT=4'h6;
  LUT2 inf_abs0_2_axb_9_cZ(.I0(ir[9:9]),.I1(ir[31:31]),.O(inf_abs0_2_axb_9));
defparam inf_abs0_2_axb_9_cZ.INIT=4'h6;
  LUT2 inf_abs0_2_axb_10_cZ(.I0(ir[10:10]),.I1(ir[31:31]),.O(inf_abs0_2_axb_10));
defparam inf_abs0_2_axb_10_cZ.INIT=4'h6;
  LUT2 inf_abs0_2_axb_11_cZ(.I0(ir[11:11]),.I1(ir[31:31]),.O(inf_abs0_2_axb_11));
defparam inf_abs0_2_axb_11_cZ.INIT=4'h6;
  LUT2 inf_abs0_2_axb_12_cZ(.I0(ir[12:12]),.I1(ir[31:31]),.O(inf_abs0_2_axb_12));
defparam inf_abs0_2_axb_12_cZ.INIT=4'h6;
  LUT2 inf_abs0_2_axb_13_cZ(.I0(ir[13:13]),.I1(ir[31:31]),.O(inf_abs0_2_axb_13));
defparam inf_abs0_2_axb_13_cZ.INIT=4'h6;
  LUT2 inf_abs0_2_axb_14_cZ(.I0(ir[14:14]),.I1(ir[31:31]),.O(inf_abs0_2_axb_14));
defparam inf_abs0_2_axb_14_cZ.INIT=4'h6;
  LUT2 inf_abs0_2_axb_15_cZ(.I0(ir[15:15]),.I1(ir[31:31]),.O(inf_abs0_2_axb_15));
defparam inf_abs0_2_axb_15_cZ.INIT=4'h6;
  LUT2 inf_abs0_2_axb_16_cZ(.I0(ir[16:16]),.I1(ir[31:31]),.O(inf_abs0_2_axb_16));
defparam inf_abs0_2_axb_16_cZ.INIT=4'h6;
  LUT2 inf_abs0_2_axb_17_cZ(.I0(ir[17:17]),.I1(ir[31:31]),.O(inf_abs0_2_axb_17));
defparam inf_abs0_2_axb_17_cZ.INIT=4'h6;
  LUT2 inf_abs0_2_axb_18_cZ(.I0(ir[18:18]),.I1(ir[31:31]),.O(inf_abs0_2_axb_18));
defparam inf_abs0_2_axb_18_cZ.INIT=4'h6;
  LUT2 inf_abs0_2_axb_19_cZ(.I0(ir[19:19]),.I1(ir[31:31]),.O(inf_abs0_2_axb_19));
defparam inf_abs0_2_axb_19_cZ.INIT=4'h6;
  LUT2 inf_abs0_2_axb_20_cZ(.I0(ir[20:20]),.I1(ir[31:31]),.O(inf_abs0_2_axb_20));
defparam inf_abs0_2_axb_20_cZ.INIT=4'h6;
  LUT2 inf_abs0_2_axb_21_cZ(.I0(ir[21:21]),.I1(ir[31:31]),.O(inf_abs0_2_axb_21));
defparam inf_abs0_2_axb_21_cZ.INIT=4'h6;
  LUT2 inf_abs0_2_axb_22_cZ(.I0(ir[22:22]),.I1(ir[31:31]),.O(inf_abs0_2_axb_22));
defparam inf_abs0_2_axb_22_cZ.INIT=4'h6;
  LUT2 inf_abs0_2_axb_23_cZ(.I0(ir[23:23]),.I1(ir[31:31]),.O(inf_abs0_2_axb_23));
defparam inf_abs0_2_axb_23_cZ.INIT=4'h6;
  LUT2 inf_abs0_2_axb_24_cZ(.I0(ir[24:24]),.I1(ir[31:31]),.O(inf_abs0_2_axb_24));
defparam inf_abs0_2_axb_24_cZ.INIT=4'h6;
  LUT2 inf_abs0_2_axb_25_cZ(.I0(ir[25:25]),.I1(ir[31:31]),.O(inf_abs0_2_axb_25));
defparam inf_abs0_2_axb_25_cZ.INIT=4'h6;
  LUT2 inf_abs0_2_axb_26_cZ(.I0(ir[26:26]),.I1(ir[31:31]),.O(inf_abs0_2_axb_26));
defparam inf_abs0_2_axb_26_cZ.INIT=4'h6;
  LUT2 inf_abs0_2_axb_27_cZ(.I0(ir[27:27]),.I1(ir[31:31]),.O(inf_abs0_2_axb_27));
defparam inf_abs0_2_axb_27_cZ.INIT=4'h6;
  LUT2 inf_abs0_2_axb_28_cZ(.I0(ir[28:28]),.I1(ir[31:31]),.O(inf_abs0_2_axb_28));
defparam inf_abs0_2_axb_28_cZ.INIT=4'h6;
  LUT4 desc4(.I0(datai[20:20]),.I1(inf_abs0_2[27:27]),.I2(inf_abs0_2[28:28]),.I3(inf_abs0_2[31:31]),.O(reg3_1_1_axb_20));
defparam desc4.INIT=16'hFF57;
  LUT4 desc5(.I0(datai[21:21]),.I1(inf_abs0_2[27:27]),.I2(inf_abs0_2[28:28]),.I3(inf_abs0_2[31:31]),.O(reg3_1_1_axb_21));
defparam desc5.INIT=16'hFF57;
  LUT4 desc6(.I0(datai[22:22]),.I1(inf_abs0_2[27:27]),.I2(inf_abs0_2[28:28]),.I3(inf_abs0_2[31:31]),.O(reg3_1_1_axb_22));
defparam desc6.INIT=16'hFF57;
  LUT4 desc7(.I0(datai[23:23]),.I1(inf_abs0_2[27:27]),.I2(inf_abs0_2[28:28]),.I3(inf_abs0_2[31:31]),.O(reg3_1_1_axb_23));
defparam desc7.INIT=16'hFF57;
  LUT4 desc8(.I0(datai[24:24]),.I1(inf_abs0_2[27:27]),.I2(inf_abs0_2[28:28]),.I3(inf_abs0_2[31:31]),.O(reg3_1_1_axb_24));
defparam desc8.INIT=16'hFF57;
  LUT4 desc9(.I0(datai[25:25]),.I1(inf_abs0_2[27:27]),.I2(inf_abs0_2[28:28]),.I3(inf_abs0_2[31:31]),.O(reg3_1_1_axb_25));
defparam desc9.INIT=16'hFF57;
  LUT4 desc10(.I0(datai[26:26]),.I1(inf_abs0_2[27:27]),.I2(inf_abs0_2[28:28]),.I3(inf_abs0_2[31:31]),.O(reg3_1_1_axb_26));
defparam desc10.INIT=16'hFF57;
  LUT4 desc11(.I0(datai[27:27]),.I1(inf_abs0_2[27:27]),.I2(inf_abs0_2[28:28]),.I3(inf_abs0_2[31:31]),.O(reg3_1_1_axb_27));
defparam desc11.INIT=16'hFF57;
  LUT4 desc12(.I0(datai[28:28]),.I1(inf_abs0_2[27:27]),.I2(inf_abs0_2[28:28]),.I3(inf_abs0_2[31:31]),.O(reg3_1_1_axb_28));
defparam desc12.INIT=16'hFF57;
  LUT4 reg3_1_1_axb_29_cZ(.I0(datai[29:29]),.I1(inf_abs0_2[27:27]),.I2(inf_abs0_2[28:28]),.I3(inf_abs0_2[31:31]),.O(reg3_1_1_axb_29));
defparam reg3_1_1_axb_29_cZ.INIT=16'hFF57;
  LUT4 reg3_1_1_axb_30_cZ(.I0(datai[30:30]),.I1(inf_abs0_2[27:27]),.I2(inf_abs0_2[28:28]),.I3(inf_abs0_2[31:31]),.O(reg3_1_1_axb_30));
defparam reg3_1_1_axb_30_cZ.INIT=16'hFF57;
  LUT2 un1_inf_abs0_cry_0_RNO(.I0(inf_abs0_2[0:0]),.I1(reg2[0:0]),.O(un1_inf_abs0_10[0:0]));
defparam un1_inf_abs0_cry_0_RNO.INIT=4'h6;
  LUT2 desc13(.I0(inf_abs0_2[1:1]),.I1(reg2[1:1]),.O(un1_inf_abs0_axb_1));
defparam desc13.INIT=4'h6;
  LUT2 desc14(.I0(inf_abs0_2[2:2]),.I1(reg2[2:2]),.O(un1_inf_abs0_axb_2));
defparam desc14.INIT=4'h6;
  LUT2 desc15(.I0(inf_abs0_2[3:3]),.I1(reg2[3:3]),.O(un1_inf_abs0_axb_3));
defparam desc15.INIT=4'h6;
  LUT2 desc16(.I0(inf_abs0_2[4:4]),.I1(reg2[4:4]),.O(un1_inf_abs0_axb_4));
defparam desc16.INIT=4'h6;
  LUT2 desc17(.I0(inf_abs0_2[5:5]),.I1(reg2[5:5]),.O(un1_inf_abs0_axb_5));
defparam desc17.INIT=4'h6;
  LUT2 desc18(.I0(inf_abs0_2[6:6]),.I1(reg2[6:6]),.O(un1_inf_abs0_axb_6));
defparam desc18.INIT=4'h6;
  LUT2 desc19(.I0(inf_abs0_2[7:7]),.I1(reg2[7:7]),.O(un1_inf_abs0_axb_7));
defparam desc19.INIT=4'h6;
  LUT2 desc20(.I0(inf_abs0_2[8:8]),.I1(reg2[8:8]),.O(un1_inf_abs0_axb_8));
defparam desc20.INIT=4'h6;
  LUT2 desc21(.I0(inf_abs0_2[9:9]),.I1(reg2[9:9]),.O(un1_inf_abs0_axb_9));
defparam desc21.INIT=4'h6;
  LUT2 desc22(.I0(inf_abs0_2[10:10]),.I1(reg2[10:10]),.O(un1_inf_abs0_axb_10));
defparam desc22.INIT=4'h6;
  LUT2 desc23(.I0(inf_abs0_2[11:11]),.I1(reg2[11:11]),.O(un1_inf_abs0_axb_11));
defparam desc23.INIT=4'h6;
  LUT2 desc24(.I0(inf_abs0_2[12:12]),.I1(reg2[12:12]),.O(un1_inf_abs0_axb_12));
defparam desc24.INIT=4'h6;
  LUT2 desc25(.I0(inf_abs0_2[13:13]),.I1(reg2[13:13]),.O(un1_inf_abs0_axb_13));
defparam desc25.INIT=4'h6;
  LUT2 desc26(.I0(inf_abs0_2[14:14]),.I1(reg2[14:14]),.O(un1_inf_abs0_axb_14));
defparam desc26.INIT=4'h6;
  LUT2 desc27(.I0(inf_abs0_2[15:15]),.I1(reg2[15:15]),.O(un1_inf_abs0_axb_15));
defparam desc27.INIT=4'h6;
  LUT2 desc28(.I0(inf_abs0_2[16:16]),.I1(reg2[16:16]),.O(un1_inf_abs0_axb_16));
defparam desc28.INIT=4'h6;
  LUT2 desc29(.I0(inf_abs0_2[17:17]),.I1(reg2[17:17]),.O(un1_inf_abs0_axb_17));
defparam desc29.INIT=4'h6;
  LUT2 desc30(.I0(inf_abs0_2[18:18]),.I1(reg2[18:18]),.O(un1_inf_abs0_axb_18));
defparam desc30.INIT=4'h6;
  LUT2 un1_inf_abs0_0_cry_0_RNO(.I0(inf_abs0_2[0:0]),.I1(reg1[0:0]),.O(un1_inf_abs0_11[0:0]));
defparam un1_inf_abs0_0_cry_0_RNO.INIT=4'h6;
  LUT2 desc31(.I0(inf_abs0_2[1:1]),.I1(reg1[1:1]),.O(un1_inf_abs0_0_axb_1));
defparam desc31.INIT=4'h6;
  LUT2 desc32(.I0(inf_abs0_2[2:2]),.I1(reg1[2:2]),.O(un1_inf_abs0_0_axb_2));
defparam desc32.INIT=4'h6;
  LUT2 desc33(.I0(inf_abs0_2[3:3]),.I1(reg1[3:3]),.O(un1_inf_abs0_0_axb_3));
defparam desc33.INIT=4'h6;
  LUT2 desc34(.I0(inf_abs0_2[4:4]),.I1(reg1[4:4]),.O(un1_inf_abs0_0_axb_4));
defparam desc34.INIT=4'h6;
  LUT2 desc35(.I0(inf_abs0_2[5:5]),.I1(reg1[5:5]),.O(un1_inf_abs0_0_axb_5));
defparam desc35.INIT=4'h6;
  LUT2 desc36(.I0(inf_abs0_2[6:6]),.I1(reg1[6:6]),.O(un1_inf_abs0_0_axb_6));
defparam desc36.INIT=4'h6;
  LUT2 desc37(.I0(inf_abs0_2[7:7]),.I1(reg1[7:7]),.O(un1_inf_abs0_0_axb_7));
defparam desc37.INIT=4'h6;
  LUT2 desc38(.I0(inf_abs0_2[8:8]),.I1(reg1[8:8]),.O(un1_inf_abs0_0_axb_8));
defparam desc38.INIT=4'h6;
  LUT2 desc39(.I0(inf_abs0_2[9:9]),.I1(reg1[9:9]),.O(un1_inf_abs0_0_axb_9));
defparam desc39.INIT=4'h6;
  LUT2 desc40(.I0(inf_abs0_2[10:10]),.I1(reg1[10:10]),.O(un1_inf_abs0_0_axb_10));
defparam desc40.INIT=4'h6;
  LUT2 desc41(.I0(inf_abs0_2[11:11]),.I1(reg1[11:11]),.O(un1_inf_abs0_0_axb_11));
defparam desc41.INIT=4'h6;
  LUT2 desc42(.I0(inf_abs0_2[12:12]),.I1(reg1[12:12]),.O(un1_inf_abs0_0_axb_12));
defparam desc42.INIT=4'h6;
  LUT2 desc43(.I0(inf_abs0_2[13:13]),.I1(reg1[13:13]),.O(un1_inf_abs0_0_axb_13));
defparam desc43.INIT=4'h6;
  LUT2 desc44(.I0(inf_abs0_2[14:14]),.I1(reg1[14:14]),.O(un1_inf_abs0_0_axb_14));
defparam desc44.INIT=4'h6;
  LUT2 desc45(.I0(inf_abs0_2[15:15]),.I1(reg1[15:15]),.O(un1_inf_abs0_0_axb_15));
defparam desc45.INIT=4'h6;
  LUT2 desc46(.I0(inf_abs0_2[16:16]),.I1(reg1[16:16]),.O(un1_inf_abs0_0_axb_16));
defparam desc46.INIT=4'h6;
  LUT2 desc47(.I0(inf_abs0_2[17:17]),.I1(reg1[17:17]),.O(un1_inf_abs0_0_axb_17));
defparam desc47.INIT=4'h6;
  LUT2 desc48(.I0(inf_abs0_2[18:18]),.I1(reg1[18:18]),.O(un1_inf_abs0_0_axb_18));
defparam desc48.INIT=4'h6;
  LUT1 un3_reg3_axb_1_cZ(.I0(reg3[4:4]),.O(un3_reg3_axb_1));
defparam un3_reg3_axb_1_cZ.INIT=2'h2;
  LUT1 un3_reg3_axb_2_cZ(.I0(reg3[5:5]),.O(un3_reg3_axb_2));
defparam un3_reg3_axb_2_cZ.INIT=2'h2;
  LUT1 un3_reg3_axb_3_cZ(.I0(reg3[6:6]),.O(un3_reg3_axb_3));
defparam un3_reg3_axb_3_cZ.INIT=2'h2;
  LUT1 un3_reg3_axb_4_cZ(.I0(reg3[7:7]),.O(un3_reg3_axb_4));
defparam un3_reg3_axb_4_cZ.INIT=2'h2;
  LUT1 un3_reg3_axb_5_cZ(.I0(reg3[8:8]),.O(un3_reg3_axb_5));
defparam un3_reg3_axb_5_cZ.INIT=2'h2;
  LUT1 un3_reg3_axb_6_cZ(.I0(reg3[9:9]),.O(un3_reg3_axb_6));
defparam un3_reg3_axb_6_cZ.INIT=2'h2;
  LUT1 un3_reg3_axb_7_cZ(.I0(reg3[10:10]),.O(un3_reg3_axb_7));
defparam un3_reg3_axb_7_cZ.INIT=2'h2;
  LUT1 un3_reg3_axb_8_cZ(.I0(reg3[11:11]),.O(un3_reg3_axb_8));
defparam un3_reg3_axb_8_cZ.INIT=2'h2;
  LUT1 un3_reg3_axb_9_cZ(.I0(reg3[12:12]),.O(un3_reg3_axb_9));
defparam un3_reg3_axb_9_cZ.INIT=2'h2;
  LUT1 un3_reg3_axb_10_cZ(.I0(reg3[13:13]),.O(un3_reg3_axb_10));
defparam un3_reg3_axb_10_cZ.INIT=2'h2;
  LUT1 un3_reg3_axb_11_cZ(.I0(reg3[14:14]),.O(un3_reg3_axb_11));
defparam un3_reg3_axb_11_cZ.INIT=2'h2;
  LUT1 un3_reg3_axb_12_cZ(.I0(reg3[15:15]),.O(un3_reg3_axb_12));
defparam un3_reg3_axb_12_cZ.INIT=2'h2;
  LUT1 un3_reg3_axb_13_cZ(.I0(reg3[16:16]),.O(un3_reg3_axb_13));
defparam un3_reg3_axb_13_cZ.INIT=2'h2;
  LUT1 un3_reg3_axb_14_cZ(.I0(reg3[17:17]),.O(un3_reg3_axb_14));
defparam un3_reg3_axb_14_cZ.INIT=2'h2;
  LUT1 un3_reg3_axb_15_cZ(.I0(reg3[18:18]),.O(un3_reg3_axb_15));
defparam un3_reg3_axb_15_cZ.INIT=2'h2;
  LUT1 un3_reg3_axb_16_cZ(.I0(reg3[19:19]),.O(un3_reg3_axb_16));
defparam un3_reg3_axb_16_cZ.INIT=2'h2;
  LUT1 un3_reg3_axb_17_cZ(.I0(reg3[20:20]),.O(un3_reg3_axb_17));
defparam un3_reg3_axb_17_cZ.INIT=2'h2;
  LUT1 un3_reg3_axb_18_cZ(.I0(reg3[21:21]),.O(un3_reg3_axb_18));
defparam un3_reg3_axb_18_cZ.INIT=2'h2;
  LUT1 un3_reg3_axb_19_cZ(.I0(reg3[22:22]),.O(un3_reg3_axb_19));
defparam un3_reg3_axb_19_cZ.INIT=2'h2;
  LUT1 un3_reg3_axb_20_cZ(.I0(reg3[23:23]),.O(un3_reg3_axb_20));
defparam un3_reg3_axb_20_cZ.INIT=2'h2;
  LUT1 un3_reg3_axb_21_cZ(.I0(reg3[24:24]),.O(un3_reg3_axb_21));
defparam un3_reg3_axb_21_cZ.INIT=2'h2;
  LUT1 un3_reg3_axb_22_cZ(.I0(reg3[25:25]),.O(un3_reg3_axb_22));
defparam un3_reg3_axb_22_cZ.INIT=2'h2;
  LUT1 un3_reg3_axb_23_cZ(.I0(reg3[26:26]),.O(un3_reg3_axb_23));
defparam un3_reg3_axb_23_cZ.INIT=2'h2;
  LUT1 un3_reg3_axb_24_cZ(.I0(reg3[27:27]),.O(un3_reg3_axb_24));
defparam un3_reg3_axb_24_cZ.INIT=2'h2;
  LUT1 un3_reg3_axb_25_cZ(.I0(reg3[28:28]),.O(un3_reg3_axb_25));
defparam un3_reg3_axb_25_cZ.INIT=2'h2;
  LUT1 un3_t_s_1_RNIB3TC(.I0(un3_t_s_1),.O(N_4541_i));
defparam un3_t_s_1_RNIB3TC.INIT=2'h1;
  LUT1 un3_t_s_2_RNIC3TC(.I0(un3_t_s_2),.O(N_4542_i));
defparam un3_t_s_2_RNIC3TC.INIT=2'h1;
  LUT1 un3_t_s_3_RNID3TC(.I0(un3_t_s_3),.O(N_4543_i));
defparam un3_t_s_3_RNID3TC.INIT=2'h1;
  LUT1 un3_t_s_4_RNIE3TC(.I0(un3_t_s_4),.O(N_4544_i));
defparam un3_t_s_4_RNIE3TC.INIT=2'h1;
  LUT1 un3_t_s_5_RNIF3TC(.I0(un3_t_s_5),.O(N_4545_i));
defparam un3_t_s_5_RNIF3TC.INIT=2'h1;
  LUT1 un3_t_s_6_RNIG3TC(.I0(un3_t_s_6),.O(N_4546_i));
defparam un3_t_s_6_RNIG3TC.INIT=2'h1;
  LUT1 un3_t_s_7_RNIH3TC(.I0(un3_t_s_7),.O(N_4547_i));
defparam un3_t_s_7_RNIH3TC.INIT=2'h1;
  LUT1 un3_t_s_8_RNII3TC(.I0(un3_t_s_8),.O(N_4548_i));
defparam un3_t_s_8_RNII3TC.INIT=2'h1;
  LUT1 un3_t_s_9_RNIJ3TC(.I0(un3_t_s_9),.O(N_4549_i));
defparam un3_t_s_9_RNIJ3TC.INIT=2'h1;
  LUT1 un3_t_s_10_RNIRF0A(.I0(un3_t_s_10),.O(N_4550_i));
defparam un3_t_s_10_RNIRF0A.INIT=2'h1;
  LUT1 un3_t_s_11_RNISF0A(.I0(un3_t_s_11),.O(N_4551_i));
defparam un3_t_s_11_RNISF0A.INIT=2'h1;
  LUT1 un3_t_s_12_RNITF0A(.I0(un3_t_s_12),.O(N_4552_i));
defparam un3_t_s_12_RNITF0A.INIT=2'h1;
  LUT1 un3_t_s_13_RNIUF0A(.I0(un3_t_s_13),.O(N_4553_i));
defparam un3_t_s_13_RNIUF0A.INIT=2'h1;
  LUT1 un3_t_s_14_RNIVF0A(.I0(un3_t_s_14),.O(N_4554_i));
defparam un3_t_s_14_RNIVF0A.INIT=2'h1;
  LUT1 un3_t_s_15_RNI0G0A(.I0(un3_t_s_15),.O(N_4555_i));
defparam un3_t_s_15_RNI0G0A.INIT=2'h1;
  LUT1 un3_t_s_16_RNI1G0A(.I0(un3_t_s_16),.O(N_4556_i));
defparam un3_t_s_16_RNI1G0A.INIT=2'h1;
  LUT1 un3_t_s_17_RNI2G0A(.I0(un3_t_s_17),.O(N_4557_i));
defparam un3_t_s_17_RNI2G0A.INIT=2'h1;
  LUT1 un3_t_s_18_RNI3G0A(.I0(un3_t_s_18),.O(N_4558_i));
defparam un3_t_s_18_RNI3G0A.INIT=2'h1;
  LUT1 un3_t_s_19_RNI4G0A(.I0(un3_t_s_19),.O(N_4559_i));
defparam un3_t_s_19_RNI4G0A.INIT=2'h1;
  LUT1 un3_t_s_20_RNISG0A(.I0(un3_t_s_20),.O(N_4560_i));
defparam un3_t_s_20_RNISG0A.INIT=2'h1;
  LUT1 un3_t_s_21_RNITG0A(.I0(un3_t_s_21),.O(N_4561_i));
defparam un3_t_s_21_RNITG0A.INIT=2'h1;
  LUT1 un3_t_s_22_RNIUG0A(.I0(un3_t_s_22),.O(N_4562_i));
defparam un3_t_s_22_RNIUG0A.INIT=2'h1;
  LUT1 un3_t_s_23_RNIVG0A(.I0(un3_t_s_23),.O(N_4563_i));
defparam un3_t_s_23_RNIVG0A.INIT=2'h1;
  LUT1 un3_t_s_24_RNI0H0A(.I0(un3_t_s_24),.O(N_4564_i));
defparam un3_t_s_24_RNI0H0A.INIT=2'h1;
  LUT1 un3_t_s_25_RNI1H0A(.I0(un3_t_s_25),.O(N_4565_i));
defparam un3_t_s_25_RNI1H0A.INIT=2'h1;
  LUT1 un3_t_s_26_RNI2H0A(.I0(un3_t_s_26),.O(N_4566_i));
defparam un3_t_s_26_RNI2H0A.INIT=2'h1;
  LUT1 un3_t_s_27_RNI3H0A(.I0(un3_t_s_27),.O(N_4567_i));
defparam un3_t_s_27_RNI3H0A.INIT=2'h1;
  LUT1 un3_t_s_28_RNI4H0A(.I0(un3_t_s_28),.O(N_4568_i));
defparam un3_t_s_28_RNI4H0A.INIT=2'h1;
  LUT1 un3_t_s_29_RNI5H0A(.I0(un3_t_s_29),.O(N_4569_i));
defparam un3_t_s_29_RNI5H0A.INIT=2'h1;
  LUT1 un3_t_s_30_RNITH0A(.I0(un3_t_s_30),.O(N_4570_i));
defparam un3_t_s_30_RNITH0A.INIT=2'h1;
  LUT1 un3_t_s_31_RNIUH0A(.I0(un3_t_s_31),.O(N_4571_i));
defparam un3_t_s_31_RNIUH0A.INIT=2'h1;
  LUT2 inf_abs0_2_axb_29_cZ(.I0(ir[29:29]),.I1(ir[31:31]),.O(inf_abs0_2_axb_29));
defparam inf_abs0_2_axb_29_cZ.INIT=4'h6;
  LUT4 un26_r_df30_cZ(.I0(m_2[30:30]),.I1(m_2_i[31:31]),.I2(r_4_i[31:31]),.I3(r_6[30:30]),.O(un26_r_df30));
defparam un26_r_df30_cZ.INIT=16'h8241;
  LUT4 desc49(.I0(m_2[30:30]),.I1(m_2[31:31]),.I2(r_4[30:30]),.I3(r_4[31:31]),.O(un14_r_0_N_2));
defparam desc49.INIT=16'h8421;
  p_O_FDC b_Z(.Q(b),.D(b_0),.C(clock),.CLR(reset),.E(p_b_Z_p_O_FDC));
  p_O_FDCE desc50(.Q(d[0:0]),.D(d_cnst),.C(clock),.CLR(reset),.CE(dce),.E(p_desc50_p_O_FDCE));
  p_O_FDCE desc51(.Q(d[1:1]),.D(d_cnst_sm0),.C(clock),.CLR(reset),.CE(dce),.E(p_desc51_p_O_FDCE));
  p_O_FDC desc52(.Q(ir[22:22]),.D(ir_3[22:22]),.C(clock),.CLR(reset),.E(p_desc52_p_O_FDC));
  p_O_FDC desc53(.Q(ir[23:23]),.D(ir_3[23:23]),.C(clock),.CLR(reset),.E(p_desc53_p_O_FDC));
  p_O_FDC desc54(.Q(ir[24:24]),.D(ir_3[24:24]),.C(clock),.CLR(reset),.E(p_desc54_p_O_FDC));
  p_O_FDC desc55(.Q(ir[25:25]),.D(ir_3[25:25]),.C(clock),.CLR(reset),.E(p_desc55_p_O_FDC));
  p_O_FDC desc56(.Q(ir[26:26]),.D(ir_3[26:26]),.C(clock),.CLR(reset),.E(p_desc56_p_O_FDC));
  p_O_FDC desc57(.Q(ir[27:27]),.D(ir_3[27:27]),.C(clock),.CLR(reset),.E(p_desc57_p_O_FDC));
  p_O_FDC desc58(.Q(ir[28:28]),.D(ir_3[28:28]),.C(clock),.CLR(reset),.E(p_desc58_p_O_FDC));
  p_O_FDC desc59(.Q(ir[29:29]),.D(ir_3[29:29]),.C(clock),.CLR(reset),.E(p_desc59_p_O_FDC));
  p_O_FDC desc60(.Q(ir[30:30]),.D(ir_3[30:30]),.C(clock),.CLR(reset),.E(p_desc60_p_O_FDC));
  p_O_FDC desc61(.Q(ir[31:31]),.D(ir_3[31:31]),.C(clock),.CLR(reset),.E(p_desc61_p_O_FDC));
  p_O_FDC desc62(.Q(ir[7:7]),.D(ir_3[7:7]),.C(clock),.CLR(reset),.E(p_desc62_p_O_FDC));
  p_O_FDC desc63(.Q(ir[8:8]),.D(ir_3[8:8]),.C(clock),.CLR(reset),.E(p_desc63_p_O_FDC));
  p_O_FDC desc64(.Q(ir[9:9]),.D(ir_3[9:9]),.C(clock),.CLR(reset),.E(p_desc64_p_O_FDC));
  p_O_FDC desc65(.Q(ir[10:10]),.D(ir_3[10:10]),.C(clock),.CLR(reset),.E(p_desc65_p_O_FDC));
  p_O_FDC desc66(.Q(ir[11:11]),.D(ir_3[11:11]),.C(clock),.CLR(reset),.E(p_desc66_p_O_FDC));
  p_O_FDC desc67(.Q(ir[12:12]),.D(ir_3[12:12]),.C(clock),.CLR(reset),.E(p_desc67_p_O_FDC));
  p_O_FDC desc68(.Q(ir[13:13]),.D(ir_3[13:13]),.C(clock),.CLR(reset),.E(p_desc68_p_O_FDC));
  p_O_FDC desc69(.Q(ir[14:14]),.D(ir_3[14:14]),.C(clock),.CLR(reset),.E(p_desc69_p_O_FDC));
  p_O_FDC desc70(.Q(ir[15:15]),.D(ir_3[15:15]),.C(clock),.CLR(reset),.E(p_desc70_p_O_FDC));
  p_O_FDC desc71(.Q(ir[16:16]),.D(ir_3[16:16]),.C(clock),.CLR(reset),.E(p_desc71_p_O_FDC));
  p_O_FDC desc72(.Q(ir[17:17]),.D(ir_3[17:17]),.C(clock),.CLR(reset),.E(p_desc72_p_O_FDC));
  p_O_FDC desc73(.Q(ir[18:18]),.D(ir_3[18:18]),.C(clock),.CLR(reset),.E(p_desc73_p_O_FDC));
  p_O_FDC desc74(.Q(ir[19:19]),.D(ir_3[19:19]),.C(clock),.CLR(reset),.E(p_desc74_p_O_FDC));
  p_O_FDC desc75(.Q(ir[20:20]),.D(ir_3[20:20]),.C(clock),.CLR(reset),.E(p_desc75_p_O_FDC));
  p_O_FDC desc76(.Q(ir[21:21]),.D(ir_3[21:21]),.C(clock),.CLR(reset),.E(p_desc76_p_O_FDC));
  p_O_FDC desc77(.Q(ir[0:0]),.D(ir_3[0:0]),.C(clock),.CLR(reset),.E(p_desc77_p_O_FDC));
  p_O_FDC desc78(.Q(ir[1:1]),.D(ir_3[1:1]),.C(clock),.CLR(reset),.E(p_desc78_p_O_FDC));
  p_O_FDC desc79(.Q(ir[2:2]),.D(ir_3[2:2]),.C(clock),.CLR(reset),.E(p_desc79_p_O_FDC));
  p_O_FDC desc80(.Q(ir[3:3]),.D(ir_3[3:3]),.C(clock),.CLR(reset),.E(p_desc80_p_O_FDC));
  p_O_FDC desc81(.Q(ir[4:4]),.D(ir_3[4:4]),.C(clock),.CLR(reset),.E(p_desc81_p_O_FDC));
  p_O_FDC desc82(.Q(ir[5:5]),.D(ir_3[5:5]),.C(clock),.CLR(reset),.E(p_desc82_p_O_FDC));
  p_O_FDC desc83(.Q(ir[6:6]),.D(ir_3[6:6]),.C(clock),.CLR(reset),.E(p_desc83_p_O_FDC));
  p_O_FDCE desc84(.Q(reg0[31:31]),.D(N_3856_rep1),.C(clock),.CLR(reset),.CE(un1_state_4_i),.E(p_desc84_p_O_FDCE));
  p_O_FDCE desc85(.Q(reg0[16:16]),.D(reg0_28[16:16]),.C(clock),.CLR(reset),.CE(un1_state_4_i),.E(p_desc85_p_O_FDCE));
  p_O_FDCE desc86(.Q(reg0[17:17]),.D(reg0_28[17:17]),.C(clock),.CLR(reset),.CE(un1_state_4_i),.E(p_desc86_p_O_FDCE));
  p_O_FDCE desc87(.Q(reg0[18:18]),.D(reg0_28[18:18]),.C(clock),.CLR(reset),.CE(un1_state_4_i),.E(p_desc87_p_O_FDCE));
  p_O_FDCE desc88(.Q(reg0[19:19]),.D(N_3829_rep1),.C(clock),.CLR(reset),.CE(un1_state_4_i),.E(p_desc88_p_O_FDCE));
  p_O_FDCE desc89(.Q(reg0[20:20]),.D(N_3803_rep1),.C(clock),.CLR(reset),.CE(un1_state_4_i),.E(p_desc89_p_O_FDCE));
  p_O_FDCE desc90(.Q(reg0[21:21]),.D(N_3777_rep1),.C(clock),.CLR(reset),.CE(un1_state_4_i),.E(p_desc90_p_O_FDCE));
  p_O_FDCE desc91(.Q(reg0[22:22]),.D(N_3751_rep1),.C(clock),.CLR(reset),.CE(un1_state_4_i),.E(p_desc91_p_O_FDCE));
  p_O_FDCE desc92(.Q(reg0[23:23]),.D(N_3725_rep1),.C(clock),.CLR(reset),.CE(un1_state_4_i),.E(p_desc92_p_O_FDCE));
  p_O_FDCE desc93(.Q(reg0[24:24]),.D(N_3699_rep1),.C(clock),.CLR(reset),.CE(un1_state_4_i),.E(p_desc93_p_O_FDCE));
  p_O_FDCE desc94(.Q(reg0[25:25]),.D(N_3673_rep1),.C(clock),.CLR(reset),.CE(un1_state_4_i),.E(p_desc94_p_O_FDCE));
  p_O_FDCE desc95(.Q(reg0[26:26]),.D(N_3341_rep1),.C(clock),.CLR(reset),.CE(un1_state_4_i),.E(p_desc95_p_O_FDCE));
  p_O_FDCE desc96(.Q(reg0[27:27]),.D(N_3315_rep1),.C(clock),.CLR(reset),.CE(un1_state_4_i),.E(p_desc96_p_O_FDCE));
  p_O_FDCE desc97(.Q(reg0[28:28]),.D(N_3289_rep1),.C(clock),.CLR(reset),.CE(un1_state_4_i),.E(p_desc97_p_O_FDCE));
  p_O_FDCE desc98(.Q(reg0[29:29]),.D(N_3569_rep1),.C(clock),.CLR(reset),.CE(un1_state_4_i),.E(p_desc98_p_O_FDCE));
  p_O_FDCE desc99(.Q(reg0[30:30]),.D(N_3550_rep1),.C(clock),.CLR(reset),.CE(un1_state_4_i),.E(p_desc99_p_O_FDCE));
  p_O_FDCE desc100(.Q(reg0[1:1]),.D(reg0_28[1:1]),.C(clock),.CLR(reset),.CE(un1_state_4_i),.E(p_desc100_p_O_FDCE));
  p_O_FDCE desc101(.Q(reg0[2:2]),.D(reg0_28[2:2]),.C(clock),.CLR(reset),.CE(un1_state_4_i),.E(p_desc101_p_O_FDCE));
  p_O_FDCE desc102(.Q(reg0[3:3]),.D(reg0_28[3:3]),.C(clock),.CLR(reset),.CE(un1_state_4_i),.E(p_desc102_p_O_FDCE));
  p_O_FDCE desc103(.Q(reg0[4:4]),.D(reg0_28[4:4]),.C(clock),.CLR(reset),.CE(un1_state_4_i),.E(p_desc103_p_O_FDCE));
  p_O_FDCE desc104(.Q(reg0[5:5]),.D(reg0_28[5:5]),.C(clock),.CLR(reset),.CE(un1_state_4_i),.E(p_desc104_p_O_FDCE));
  p_O_FDCE desc105(.Q(reg0[6:6]),.D(reg0_28[6:6]),.C(clock),.CLR(reset),.CE(un1_state_4_i),.E(p_desc105_p_O_FDCE));
  p_O_FDCE desc106(.Q(reg0[7:7]),.D(reg0_28_7_rep1),.C(clock),.CLR(reset),.CE(un1_state_4_i),.E(p_desc106_p_O_FDCE));
  p_O_FDCE desc107(.Q(reg0[8:8]),.D(reg0_28[8:8]),.C(clock),.CLR(reset),.CE(un1_state_4_i),.E(p_desc107_p_O_FDCE));
  p_O_FDCE desc108(.Q(reg0[9:9]),.D(reg0_28[9:9]),.C(clock),.CLR(reset),.CE(un1_state_4_i),.E(p_desc108_p_O_FDCE));
  p_O_FDCE desc109(.Q(reg0[10:10]),.D(reg0_28[10:10]),.C(clock),.CLR(reset),.CE(un1_state_4_i),.E(p_desc109_p_O_FDCE));
  p_O_FDCE desc110(.Q(reg0[11:11]),.D(reg0_28[11:11]),.C(clock),.CLR(reset),.CE(un1_state_4_i),.E(p_desc110_p_O_FDCE));
  p_O_FDCE desc111(.Q(reg0[12:12]),.D(reg0_28[12:12]),.C(clock),.CLR(reset),.CE(un1_state_4_i),.E(p_desc111_p_O_FDCE));
  p_O_FDCE desc112(.Q(reg0[13:13]),.D(reg0_28[13:13]),.C(clock),.CLR(reset),.CE(un1_state_4_i),.E(p_desc112_p_O_FDCE));
  p_O_FDCE desc113(.Q(reg0[14:14]),.D(reg0_28[14:14]),.C(clock),.CLR(reset),.CE(un1_state_4_i),.E(p_desc113_p_O_FDCE));
  p_O_FDCE desc114(.Q(reg0[15:15]),.D(reg0_28[15:15]),.C(clock),.CLR(reset),.CE(un1_state_4_i),.E(p_desc114_p_O_FDCE));
  p_O_FDCE desc115(.Q(reg1[18:18]),.D(reg1_16[18:18]),.C(clock),.CLR(reset),.CE(un1_state_3_i),.E(p_desc115_p_O_FDCE));
  p_O_FDCE desc116(.Q(reg1[19:19]),.D(reg0_28_3_2492),.C(clock),.CLR(reset),.CE(un1_state_3_i),.E(p_desc116_p_O_FDCE));
  p_O_FDCE desc117(.Q(reg1[20:20]),.D(reg0_28_4_2459),.C(clock),.CLR(reset),.CE(un1_state_3_i),.E(p_desc117_p_O_FDCE));
  p_O_FDCE desc118(.Q(reg1[21:21]),.D(reg0_28_5_2426),.C(clock),.CLR(reset),.CE(un1_state_3_i),.E(p_desc118_p_O_FDCE));
  p_O_FDCE desc119(.Q(reg1[22:22]),.D(reg0_28_6_2393),.C(clock),.CLR(reset),.CE(un1_state_3_i),.E(p_desc119_p_O_FDCE));
  p_O_FDCE desc120(.Q(reg1[23:23]),.D(reg0_28_7_2360),.C(clock),.CLR(reset),.CE(un1_state_3_i),.E(p_desc120_p_O_FDCE));
  p_O_FDCE desc121(.Q(reg1[24:24]),.D(reg0_28_8_2327),.C(clock),.CLR(reset),.CE(un1_state_3_i),.E(p_desc121_p_O_FDCE));
  p_O_FDCE desc122(.Q(reg1[25:25]),.D(N_3673),.C(clock),.CLR(reset),.CE(un1_state_3_i),.E(p_desc122_p_O_FDCE));
  p_O_FDCE desc123(.Q(reg1[26:26]),.D(reg1_16_7_1870),.C(clock),.CLR(reset),.CE(un1_state_3_i),.E(p_desc123_p_O_FDCE));
  p_O_FDCE desc124(.Q(reg1[27:27]),.D(reg1_16_8_1837),.C(clock),.CLR(reset),.CE(un1_state_3_i),.E(p_desc124_p_O_FDCE));
  p_O_FDCE desc125(.Q(reg1[28:28]),.D(reg1_16_9),.C(clock),.CLR(reset),.CE(un1_state_3_i),.E(p_desc125_p_O_FDCE));
  p_O_FDCE desc126(.Q(reg1[29:29]),.D(reg0_28_10_2261_a6_3_2_lut6_2_RNIOK9O5),.C(clock),.CLR(reset),.CE(un1_state_3_i),.E(p_desc126_p_O_FDCE));
  p_O_FDCE desc127(.Q(reg1[30:30]),.D(N_3550),.C(clock),.CLR(reset),.CE(un1_state_3_i),.E(p_desc127_p_O_FDCE));
  p_O_FDCE desc128(.Q(reg1[31:31]),.D(N_3856),.C(clock),.CLR(reset),.CE(un1_state_3_i),.E(p_desc128_p_O_FDCE));
  p_O_FDCE desc129(.Q(reg0[0:0]),.D(reg0_28[0:0]),.C(clock),.CLR(reset),.CE(un1_state_4_i),.E(p_desc129_p_O_FDCE));
  p_O_FDCE desc130(.Q(reg1[3:3]),.D(reg1_16[3:3]),.C(clock),.CLR(reset),.CE(un1_state_3_i),.E(p_desc130_p_O_FDCE));
  p_O_FDCE desc131(.Q(reg1[4:4]),.D(reg1_16[4:4]),.C(clock),.CLR(reset),.CE(un1_state_3_i),.E(p_desc131_p_O_FDCE));
  p_O_FDCE desc132(.Q(reg1[5:5]),.D(reg1_16[5:5]),.C(clock),.CLR(reset),.CE(un1_state_3_i),.E(p_desc132_p_O_FDCE));
  p_O_FDCE desc133(.Q(reg1[6:6]),.D(reg1_16[6:6]),.C(clock),.CLR(reset),.CE(un1_state_3_i),.E(p_desc133_p_O_FDCE));
  p_O_FDCE desc134(.Q(reg1[7:7]),.D(reg0_28[7:7]),.C(clock),.CLR(reset),.CE(un1_state_3_i),.E(p_desc134_p_O_FDCE));
  p_O_FDCE desc135(.Q(reg1[8:8]),.D(reg1_16[8:8]),.C(clock),.CLR(reset),.CE(un1_state_3_i),.E(p_desc135_p_O_FDCE));
  p_O_FDCE desc136(.Q(reg1[9:9]),.D(reg1_16[9:9]),.C(clock),.CLR(reset),.CE(un1_state_3_i),.E(p_desc136_p_O_FDCE));
  p_O_FDCE desc137(.Q(reg1[10:10]),.D(reg1_16[10:10]),.C(clock),.CLR(reset),.CE(un1_state_3_i),.E(p_desc137_p_O_FDCE));
  p_O_FDCE desc138(.Q(reg1[11:11]),.D(reg1_16[11:11]),.C(clock),.CLR(reset),.CE(un1_state_3_i),.E(p_desc138_p_O_FDCE));
  p_O_FDCE desc139(.Q(reg1[12:12]),.D(reg1_16[12:12]),.C(clock),.CLR(reset),.CE(un1_state_3_i),.E(p_desc139_p_O_FDCE));
  p_O_FDCE desc140(.Q(reg1[13:13]),.D(reg1_16[13:13]),.C(clock),.CLR(reset),.CE(un1_state_3_i),.E(p_desc140_p_O_FDCE));
  p_O_FDCE desc141(.Q(reg1[14:14]),.D(reg1_16[14:14]),.C(clock),.CLR(reset),.CE(un1_state_3_i),.E(p_desc141_p_O_FDCE));
  p_O_FDCE desc142(.Q(reg1[15:15]),.D(reg1_16[15:15]),.C(clock),.CLR(reset),.CE(un1_state_3_i),.E(p_desc142_p_O_FDCE));
  p_O_FDCE desc143(.Q(reg1[16:16]),.D(reg1_16[16:16]),.C(clock),.CLR(reset),.CE(un1_state_3_i),.E(p_desc143_p_O_FDCE));
  p_O_FDCE desc144(.Q(reg1[17:17]),.D(reg1_16[17:17]),.C(clock),.CLR(reset),.CE(un1_state_3_i),.E(p_desc144_p_O_FDCE));
  p_O_FDCE desc145(.Q(reg2[20:20]),.D(reg2_16[20:20]),.C(clock),.CLR(reset),.CE(un1_state_1_0_i),.E(p_desc145_p_O_FDCE));
  p_O_FDCE desc146(.Q(reg2[21:21]),.D(reg2_16[21:21]),.C(clock),.CLR(reset),.CE(un1_state_1_0_i),.E(p_desc146_p_O_FDCE));
  p_O_FDCE desc147(.Q(reg2[22:22]),.D(reg2_16[22:22]),.C(clock),.CLR(reset),.CE(un1_state_1_0_i),.E(p_desc147_p_O_FDCE));
  p_O_FDCE desc148(.Q(reg2[23:23]),.D(reg2_16[23:23]),.C(clock),.CLR(reset),.CE(un1_state_1_0_i),.E(p_desc148_p_O_FDCE));
  p_O_FDCE desc149(.Q(reg2[24:24]),.D(reg2_16[24:24]),.C(clock),.CLR(reset),.CE(un1_state_1_0_i),.E(p_desc149_p_O_FDCE));
  p_O_FDCE desc150(.Q(reg2[25:25]),.D(reg2_16[25:25]),.C(clock),.CLR(reset),.CE(un1_state_1_0_i),.E(p_desc150_p_O_FDCE));
  p_O_FDCE desc151(.Q(reg2[26:26]),.D(reg2_16[26:26]),.C(clock),.CLR(reset),.CE(un1_state_1_0_i),.E(p_desc151_p_O_FDCE));
  p_O_FDCE desc152(.Q(reg2[27:27]),.D(reg2_16[27:27]),.C(clock),.CLR(reset),.CE(un1_state_1_0_i),.E(p_desc152_p_O_FDCE));
  p_O_FDCE desc153(.Q(reg2[28:28]),.D(reg2_16[28:28]),.C(clock),.CLR(reset),.CE(un1_state_1_0_i),.E(p_desc153_p_O_FDCE));
  p_O_FDCE desc154(.Q(reg2[29:29]),.D(reg2_16[29:29]),.C(clock),.CLR(reset),.CE(un1_state_1_0_i),.E(p_desc154_p_O_FDCE));
  p_O_FDCE desc155(.Q(reg2[30:30]),.D(reg2_16[30:30]),.C(clock),.CLR(reset),.CE(un1_state_1_0_i),.E(p_desc155_p_O_FDCE));
  p_O_FDCE desc156(.Q(reg2[31:31]),.D(reg2_16[31:31]),.C(clock),.CLR(reset),.CE(un1_state_1_0_i),.E(p_desc156_p_O_FDCE));
  p_O_FDCE desc157(.Q(reg1[0:0]),.D(reg1_16[0:0]),.C(clock),.CLR(reset),.CE(un1_state_3_i),.E(p_desc157_p_O_FDCE));
  p_O_FDCE desc158(.Q(reg1[1:1]),.D(reg1_16[1:1]),.C(clock),.CLR(reset),.CE(un1_state_3_i),.E(p_desc158_p_O_FDCE));
  p_O_FDCE desc159(.Q(reg1[2:2]),.D(reg1_16[2:2]),.C(clock),.CLR(reset),.CE(un1_state_3_i),.E(p_desc159_p_O_FDCE));
  p_O_FDCE desc160(.Q(reg2[5:5]),.D(reg2_16[5:5]),.C(clock),.CLR(reset),.CE(un1_state_1_0_i),.E(p_desc160_p_O_FDCE));
  p_O_FDCE desc161(.Q(reg2[6:6]),.D(reg2_16[6:6]),.C(clock),.CLR(reset),.CE(un1_state_1_0_i),.E(p_desc161_p_O_FDCE));
  p_O_FDCE desc162(.Q(reg2[7:7]),.D(reg2_16[7:7]),.C(clock),.CLR(reset),.CE(un1_state_1_0_i),.E(p_desc162_p_O_FDCE));
  p_O_FDCE desc163(.Q(reg2[8:8]),.D(reg2_16[8:8]),.C(clock),.CLR(reset),.CE(un1_state_1_0_i),.E(p_desc163_p_O_FDCE));
  p_O_FDCE desc164(.Q(reg2[9:9]),.D(reg2_16[9:9]),.C(clock),.CLR(reset),.CE(un1_state_1_0_i),.E(p_desc164_p_O_FDCE));
  p_O_FDCE desc165(.Q(reg2[10:10]),.D(reg2_16[10:10]),.C(clock),.CLR(reset),.CE(un1_state_1_0_i),.E(p_desc165_p_O_FDCE));
  p_O_FDCE desc166(.Q(reg2[11:11]),.D(reg2_16[11:11]),.C(clock),.CLR(reset),.CE(un1_state_1_0_i),.E(p_desc166_p_O_FDCE));
  p_O_FDCE desc167(.Q(reg2[12:12]),.D(reg2_16[12:12]),.C(clock),.CLR(reset),.CE(un1_state_1_0_i),.E(p_desc167_p_O_FDCE));
  p_O_FDCE desc168(.Q(reg2[13:13]),.D(reg2_16[13:13]),.C(clock),.CLR(reset),.CE(un1_state_1_0_i),.E(p_desc168_p_O_FDCE));
  p_O_FDCE desc169(.Q(reg2[14:14]),.D(reg2_16[14:14]),.C(clock),.CLR(reset),.CE(un1_state_1_0_i),.E(p_desc169_p_O_FDCE));
  p_O_FDCE desc170(.Q(reg2[15:15]),.D(reg2_16[15:15]),.C(clock),.CLR(reset),.CE(un1_state_1_0_i),.E(p_desc170_p_O_FDCE));
  p_O_FDCE desc171(.Q(reg2[16:16]),.D(reg2_16[16:16]),.C(clock),.CLR(reset),.CE(un1_state_1_0_i),.E(p_desc171_p_O_FDCE));
  p_O_FDCE desc172(.Q(reg2[17:17]),.D(reg2_16[17:17]),.C(clock),.CLR(reset),.CE(un1_state_1_0_i),.E(p_desc172_p_O_FDCE));
  p_O_FDCE desc173(.Q(reg2[18:18]),.D(reg2_16[18:18]),.C(clock),.CLR(reset),.CE(un1_state_1_0_i),.E(p_desc173_p_O_FDCE));
  p_O_FDCE desc174(.Q(reg2[19:19]),.D(reg2_16[19:19]),.C(clock),.CLR(reset),.CE(un1_state_1_0_i),.E(p_desc174_p_O_FDCE));
  p_O_FDCE desc175(.Q(datao[22:22]),.D(r_4_3_1690_i_m2),.C(clock),.CLR(reset),.CE(addr_4_sqmuxa_1),.E(p_desc175_p_O_FDCE));
  p_O_FDCE desc176(.Q(datao[23:23]),.D(r_4_3_0_1664_i_m2),.C(clock),.CLR(reset),.CE(addr_4_sqmuxa_1),.E(p_desc176_p_O_FDCE));
  p_O_FDCE desc177(.Q(datao[24:24]),.D(r_4_3_1_1638_i_m2),.C(clock),.CLR(reset),.CE(addr_4_sqmuxa_1),.E(p_desc177_p_O_FDCE));
  p_O_FDCE desc178(.Q(datao[25:25]),.D(r_4_3_2_1612_i_m2),.C(clock),.CLR(reset),.CE(addr_4_sqmuxa_1),.E(p_desc178_p_O_FDCE));
  p_O_FDCE desc179(.Q(datao[26:26]),.D(r_4_3_3_1586_i_m2),.C(clock),.CLR(reset),.CE(addr_4_sqmuxa_1),.E(p_desc179_p_O_FDCE));
  p_O_FDCE desc180(.Q(datao[27:27]),.D(r_4_3_4_1560_i_m2),.C(clock),.CLR(reset),.CE(addr_4_sqmuxa_1),.E(p_desc180_p_O_FDCE));
  p_O_FDCE desc181(.Q(datao[28:28]),.D(r_4_3_5_1534_i_m2),.C(clock),.CLR(reset),.CE(addr_4_sqmuxa_1),.E(p_desc181_p_O_FDCE));
  p_O_FDCE desc182(.Q(datao[29:29]),.D(r_4_3_6_1508_i_m2),.C(clock),.CLR(reset),.CE(addr_4_sqmuxa_1),.E(p_desc182_p_O_FDCE));
  p_O_FDCE desc183(.Q(datao[30:30]),.D(r_4_3_lut6_2_O5[30:30]),.C(clock),.CLR(reset),.CE(addr_4_sqmuxa_1),.E(p_desc183_p_O_FDCE));
  p_O_FDCE desc184(.Q(datao[31:31]),.D(r_4_3_8_1467),.C(clock),.CLR(reset),.CE(addr_4_sqmuxa_1),.E(p_desc184_p_O_FDCE));
  p_O_FDCE desc185(.Q(reg2[0:0]),.D(reg2_16[0:0]),.C(clock),.CLR(reset),.CE(un1_state_1_0_i),.E(p_desc185_p_O_FDCE));
  p_O_FDCE desc186(.Q(reg2[1:1]),.D(reg2_16[1:1]),.C(clock),.CLR(reset),.CE(un1_state_1_0_i),.E(p_desc186_p_O_FDCE));
  p_O_FDCE desc187(.Q(reg2[2:2]),.D(reg2_16[2:2]),.C(clock),.CLR(reset),.CE(un1_state_1_0_i),.E(p_desc187_p_O_FDCE));
  p_O_FDCE desc188(.Q(reg2[3:3]),.D(reg2_16[3:3]),.C(clock),.CLR(reset),.CE(un1_state_1_0_i),.E(p_desc188_p_O_FDCE));
  p_O_FDCE desc189(.Q(reg2[4:4]),.D(reg2_16[4:4]),.C(clock),.CLR(reset),.CE(un1_state_1_0_i),.E(p_desc189_p_O_FDCE));
  p_O_FDCE desc190(.Q(datao[7:7]),.D(r_4_3_9_1442_i_m2),.C(clock),.CLR(reset),.CE(addr_4_sqmuxa_1),.E(p_desc190_p_O_FDCE));
  p_O_FDCE desc191(.Q(datao[8:8]),.D(r_4_3_10_1416_i_m2),.C(clock),.CLR(reset),.CE(addr_4_sqmuxa_1),.E(p_desc191_p_O_FDCE));
  p_O_FDCE desc192(.Q(datao[9:9]),.D(r_4_3_11_1390_i_m2),.C(clock),.CLR(reset),.CE(addr_4_sqmuxa_1),.E(p_desc192_p_O_FDCE));
  p_O_FDCE desc193(.Q(datao[10:10]),.D(r_4_3_12_1364_i_m2),.C(clock),.CLR(reset),.CE(addr_4_sqmuxa_1),.E(p_desc193_p_O_FDCE));
  p_O_FDCE desc194(.Q(datao[11:11]),.D(r_4_3_13_1338_i_m2),.C(clock),.CLR(reset),.CE(addr_4_sqmuxa_1),.E(p_desc194_p_O_FDCE));
  p_O_FDCE desc195(.Q(datao[12:12]),.D(r_4_3_14_1312_i_m2),.C(clock),.CLR(reset),.CE(addr_4_sqmuxa_1),.E(p_desc195_p_O_FDCE));
  p_O_FDCE desc196(.Q(datao[13:13]),.D(r_4_3_15_1286_i_m2),.C(clock),.CLR(reset),.CE(addr_4_sqmuxa_1),.E(p_desc196_p_O_FDCE));
  p_O_FDCE desc197(.Q(datao[14:14]),.D(r_4_3_16_1260_i_m2),.C(clock),.CLR(reset),.CE(addr_4_sqmuxa_1),.E(p_desc197_p_O_FDCE));
  p_O_FDCE desc198(.Q(datao[15:15]),.D(r_4_3_17_1234_i_m2),.C(clock),.CLR(reset),.CE(addr_4_sqmuxa_1),.E(p_desc198_p_O_FDCE));
  p_O_FDCE desc199(.Q(datao[16:16]),.D(r_4_3_18_1208_i_m2),.C(clock),.CLR(reset),.CE(addr_4_sqmuxa_1),.E(p_desc199_p_O_FDCE));
  p_O_FDCE desc200(.Q(datao[17:17]),.D(r_4_3_19_1182_i_m2),.C(clock),.CLR(reset),.CE(addr_4_sqmuxa_1),.E(p_desc200_p_O_FDCE));
  p_O_FDCE desc201(.Q(datao[18:18]),.D(r_4_3_20_1156_i_m2),.C(clock),.CLR(reset),.CE(addr_4_sqmuxa_1),.E(p_desc201_p_O_FDCE));
  p_O_FDCE desc202(.Q(datao[19:19]),.D(N_2724),.C(clock),.CLR(reset),.CE(addr_4_sqmuxa_1),.E(p_desc202_p_O_FDCE));
  p_O_FDCE desc203(.Q(datao[20:20]),.D(r_4_3_22_1104_i_m2),.C(clock),.CLR(reset),.CE(addr_4_sqmuxa_1),.E(p_desc203_p_O_FDCE));
  p_O_FDCE desc204(.Q(datao[21:21]),.D(r_4_3_23_1078_i_m2),.C(clock),.CLR(reset),.CE(addr_4_sqmuxa_1),.E(p_desc204_p_O_FDCE));
  p_O_FDCE desc205(.Q(addr[12:12]),.D(N_2656_i),.C(clock),.CLR(reset),.CE(addr_0_sqmuxa_1_i),.E(p_desc205_p_O_FDCE));
  p_O_FDCE desc206(.Q(addr[13:13]),.D(N_2636_i),.C(clock),.CLR(reset),.CE(addr_0_sqmuxa_1_i),.E(p_desc206_p_O_FDCE));
  p_O_FDCE desc207(.Q(addr[14:14]),.D(N_2616_i),.C(clock),.CLR(reset),.CE(addr_0_sqmuxa_1_i),.E(p_desc207_p_O_FDCE));
  p_O_FDCE desc208(.Q(addr[15:15]),.D(N_2596_i),.C(clock),.CLR(reset),.CE(addr_0_sqmuxa_1_i),.E(p_desc208_p_O_FDCE));
  p_O_FDCE desc209(.Q(addr[16:16]),.D(N_2576_i),.C(clock),.CLR(reset),.CE(addr_0_sqmuxa_1_i),.E(p_desc209_p_O_FDCE));
  p_O_FDCE desc210(.Q(addr[17:17]),.D(N_2556_i),.C(clock),.CLR(reset),.CE(addr_0_sqmuxa_1_i),.E(p_desc210_p_O_FDCE));
  p_O_FDCE desc211(.Q(addr[18:18]),.D(N_2536_i),.C(clock),.CLR(reset),.CE(addr_0_sqmuxa_1_i),.E(p_desc211_p_O_FDCE));
  p_O_FDCE desc212(.Q(addr[19:19]),.D(N_2516_i),.C(clock),.CLR(reset),.CE(addr_0_sqmuxa_1_i),.E(p_desc212_p_O_FDCE));
  p_O_FDCE desc213(.Q(datao[0:0]),.D(r_4_3_24_836_i_m2),.C(clock),.CLR(reset),.CE(addr_4_sqmuxa_1),.E(p_desc213_p_O_FDCE));
  p_O_FDCE desc214(.Q(datao[1:1]),.D(r_4_3_25_810_i_m2),.C(clock),.CLR(reset),.CE(addr_4_sqmuxa_1),.E(p_desc214_p_O_FDCE));
  p_O_FDCE desc215(.Q(datao[2:2]),.D(N_36_i),.C(clock),.CLR(reset),.CE(addr_4_sqmuxa_1),.E(p_desc215_p_O_FDCE));
  p_O_FDCE desc216(.Q(datao[3:3]),.D(r_4_3_27_758_i_m2),.C(clock),.CLR(reset),.CE(addr_4_sqmuxa_1),.E(p_desc216_p_O_FDCE));
  p_O_FDCE desc217(.Q(datao[4:4]),.D(r_4_3_28_732_i_m2),.C(clock),.CLR(reset),.CE(addr_4_sqmuxa_1),.E(p_desc217_p_O_FDCE));
  p_O_FDCE desc218(.Q(datao[5:5]),.D(r_4_3_29_706_i_m2),.C(clock),.CLR(reset),.CE(addr_4_sqmuxa_1),.E(p_desc218_p_O_FDCE));
  p_O_FDCE desc219(.Q(datao[6:6]),.D(r_4_3_30_680_i_m2),.C(clock),.CLR(reset),.CE(addr_4_sqmuxa_1),.E(p_desc219_p_O_FDCE));
  p_O_FDCE desc220(.Q(reg3[26:26]),.D(reg3_17[26:26]),.C(clock),.CLR(reset),.CE(state),.E(p_desc220_p_O_FDCE));
  p_O_FDCE desc221(.Q(reg3[27:27]),.D(reg3_17[27:27]),.C(clock),.CLR(reset),.CE(state),.E(p_desc221_p_O_FDCE));
  p_O_FDCE desc222(.Q(reg3[28:28]),.D(reg3_17[28:28]),.C(clock),.CLR(reset),.CE(state),.E(p_desc222_p_O_FDCE));
  p_O_FDCE desc223(.Q(addr[0:0]),.D(N_2335_i),.C(clock),.CLR(reset),.CE(addr_0_sqmuxa_1_i),.E(p_desc223_p_O_FDCE));
  p_O_FDCE desc224(.Q(addr[1:1]),.D(N_2315_i),.C(clock),.CLR(reset),.CE(addr_0_sqmuxa_1_i),.E(p_desc224_p_O_FDCE));
  p_O_FDCE desc225(.Q(addr[2:2]),.D(N_47_i),.C(clock),.CLR(reset),.CE(addr_0_sqmuxa_1_i),.E(p_desc225_p_O_FDCE));
  p_O_FDCE desc226(.Q(addr[3:3]),.D(N_2267_i),.C(clock),.CLR(reset),.CE(addr_0_sqmuxa_1_i),.E(p_desc226_p_O_FDCE));
  p_O_FDCE desc227(.Q(addr[4:4]),.D(N_56_i),.C(clock),.CLR(reset),.CE(addr_0_sqmuxa_1_i),.E(p_desc227_p_O_FDCE));
  p_O_FDCE desc228(.Q(addr[5:5]),.D(N_2219_i),.C(clock),.CLR(reset),.CE(addr_0_sqmuxa_1_i),.E(p_desc228_p_O_FDCE));
  p_O_FDCE desc229(.Q(addr[6:6]),.D(N_2199_i),.C(clock),.CLR(reset),.CE(addr_0_sqmuxa_1_i),.E(p_desc229_p_O_FDCE));
  p_O_FDCE desc230(.Q(addr[7:7]),.D(N_2179_i),.C(clock),.CLR(reset),.CE(addr_0_sqmuxa_1_i),.E(p_desc230_p_O_FDCE));
  p_O_FDCE desc231(.Q(addr[8:8]),.D(N_2159_i),.C(clock),.CLR(reset),.CE(addr_0_sqmuxa_1_i),.E(p_desc231_p_O_FDCE));
  p_O_FDCE desc232(.Q(addr[9:9]),.D(N_2139_i),.C(clock),.CLR(reset),.CE(addr_0_sqmuxa_1_i),.E(p_desc232_p_O_FDCE));
  p_O_FDCE desc233(.Q(addr[10:10]),.D(N_2119_i),.C(clock),.CLR(reset),.CE(addr_0_sqmuxa_1_i),.E(p_desc233_p_O_FDCE));
  p_O_FDCE desc234(.Q(addr[11:11]),.D(N_2099_i),.C(clock),.CLR(reset),.CE(addr_0_sqmuxa_1_i),.E(p_desc234_p_O_FDCE));
  p_O_FDCE desc235(.Q(reg3[11:11]),.D(reg3_17[11:11]),.C(clock),.CLR(reset),.CE(state),.E(p_desc235_p_O_FDCE));
  p_O_FDCE desc236(.Q(reg3[12:12]),.D(reg3_17[12:12]),.C(clock),.CLR(reset),.CE(state),.E(p_desc236_p_O_FDCE));
  p_O_FDCE desc237(.Q(reg3[13:13]),.D(reg3_17[13:13]),.C(clock),.CLR(reset),.CE(state),.E(p_desc237_p_O_FDCE));
  p_O_FDCE desc238(.Q(reg3[14:14]),.D(reg3_17[14:14]),.C(clock),.CLR(reset),.CE(state),.E(p_desc238_p_O_FDCE));
  p_O_FDCE desc239(.Q(reg3[15:15]),.D(reg3_17[15:15]),.C(clock),.CLR(reset),.CE(state),.E(p_desc239_p_O_FDCE));
  p_O_FDCE desc240(.Q(reg3[16:16]),.D(reg3_17[16:16]),.C(clock),.CLR(reset),.CE(state),.E(p_desc240_p_O_FDCE));
  p_O_FDCE desc241(.Q(reg3[17:17]),.D(reg3_17[17:17]),.C(clock),.CLR(reset),.CE(state),.E(p_desc241_p_O_FDCE));
  p_O_FDCE desc242(.Q(reg3[18:18]),.D(reg3_17[18:18]),.C(clock),.CLR(reset),.CE(state),.E(p_desc242_p_O_FDCE));
  p_O_FDCE desc243(.Q(reg3[19:19]),.D(reg3_17[19:19]),.C(clock),.CLR(reset),.CE(state),.E(p_desc243_p_O_FDCE));
  p_O_FDCE desc244(.Q(reg3[20:20]),.D(reg3_17[20:20]),.C(clock),.CLR(reset),.CE(state),.E(p_desc244_p_O_FDCE));
  p_O_FDCE desc245(.Q(reg3[21:21]),.D(reg3_17[21:21]),.C(clock),.CLR(reset),.CE(state),.E(p_desc245_p_O_FDCE));
  p_O_FDCE desc246(.Q(reg3[22:22]),.D(reg3_17[22:22]),.C(clock),.CLR(reset),.CE(state),.E(p_desc246_p_O_FDCE));
  p_O_FDCE desc247(.Q(reg3[23:23]),.D(reg3_17[23:23]),.C(clock),.CLR(reset),.CE(state),.E(p_desc247_p_O_FDCE));
  p_O_FDCE desc248(.Q(reg3[24:24]),.D(reg3_17[24:24]),.C(clock),.CLR(reset),.CE(state),.E(p_desc248_p_O_FDCE));
  p_O_FDCE desc249(.Q(reg3[25:25]),.D(reg3_17[25:25]),.C(clock),.CLR(reset),.CE(state),.E(p_desc249_p_O_FDCE));
  p_O_FDCE desc250(.Q(reg3[0:0]),.D(reg3_17[0:0]),.C(clock),.CLR(reset),.CE(state),.E(p_desc250_p_O_FDCE));
  p_O_FDCE desc251(.Q(reg3[1:1]),.D(reg3_17[1:1]),.C(clock),.CLR(reset),.CE(state),.E(p_desc251_p_O_FDCE));
  p_O_FDCE desc252(.Q(reg3[2:2]),.D(reg3_17[2:2]),.C(clock),.CLR(reset),.CE(state),.E(p_desc252_p_O_FDCE));
  p_O_FDCE desc253(.Q(reg3[3:3]),.D(\d_cnst_sn.reg3_N_7_i ),.C(clock),.CLR(reset),.CE(state),.E(p_desc253_p_O_FDCE));
  p_O_FDCE desc254(.Q(reg3[4:4]),.D(reg3_17[4:4]),.C(clock),.CLR(reset),.CE(state),.E(p_desc254_p_O_FDCE));
  p_O_FDCE desc255(.Q(reg3[5:5]),.D(reg3_17[5:5]),.C(clock),.CLR(reset),.CE(state),.E(p_desc255_p_O_FDCE));
  p_O_FDCE desc256(.Q(reg3[6:6]),.D(reg3_17[6:6]),.C(clock),.CLR(reset),.CE(state),.E(p_desc256_p_O_FDCE));
  p_O_FDCE desc257(.Q(reg3[7:7]),.D(reg3_17[7:7]),.C(clock),.CLR(reset),.CE(state),.E(p_desc257_p_O_FDCE));
  p_O_FDCE desc258(.Q(reg3[8:8]),.D(reg3_17[8:8]),.C(clock),.CLR(reset),.CE(state),.E(p_desc258_p_O_FDCE));
  p_O_FDCE desc259(.Q(reg3[9:9]),.D(reg3_17[9:9]),.C(clock),.CLR(reset),.CE(state),.E(p_desc259_p_O_FDCE));
  p_O_FDCE desc260(.Q(reg3[10:10]),.D(reg3_17[10:10]),.C(clock),.CLR(reset),.CE(state),.E(p_desc260_p_O_FDCE));
  p_O_FDC rd_Z(.Q(rd),.D(rd_18),.C(clock),.CLR(reset),.E(p_rd_Z_p_O_FDC));
  p_O_FDC desc261(.Q(state),.D(state_i),.C(clock),.CLR(reset),.E(p_desc261_p_O_FDC));
  p_O_FDC wr_Z(.Q(wr),.D(addr_4_sqmuxa_1),.C(clock),.CLR(reset),.E(p_wr_Z_p_O_FDC));
  p_O_FDC desc262(.Q(ir_fast[31:31]),.D(ir_3_fast[31:31]),.C(clock),.CLR(reset),.E(p_desc262_p_O_FDC));
  MUXCY_L inf_abs0_2_cry_29_outext(.DI(GND),.CI(inf_abs0_2_cry_29_0),.S(inf_abs0_2_cry_29_1),.LO(inf_abs0_2_cry_29));
  MUXCY un3_reg3_cry_25_outext(.DI(GND),.CI(un3_reg3_cry_25_0),.S(un3_reg3_cry_25_1),.O(un3_reg3_cry_25));
  MUXCY inf_abs0_2_cry_30_outext(.DI(GND),.CI(inf_abs0_2_0[31:31]),.S(inf_abs0_2_1[31:31]),.O(inf_abs0_2[31:31]));
  MUXCY un14_r_0_I_83_cZ(.DI(GND),.CI(un14_r_0_data_tmp[9:9]),.S(un14_r_0_N_2),.O(un14_r_0_I_83));
  MUXCY desc263(.DI(un11_r_lt30),.CI(un11_r_cry[28:28]),.S(un11_r_df30),.O(un11_r_cry[30:30]));
  MUXCY desc264(.DI(b18_lt30),.CI(b18_cry[28:28]),.S(b18_df30),.O(b18));
  MUXCY desc265(.DI(un26_r_lt30),.CI(un26_r_cry[28:28]),.S(un26_r_df30),.O(un26_r_cry[30:30]));
  MUXCY inf_abs0_2_cry_29_cZ(.DI(GND),.CI(inf_abs0_2_cry_28),.S(inf_abs0_2_axb_29),.O(inf_abs0_2_cry_29_0));
  LUT5 desc266(.I0(d[0:0]),.I1(d[1:1]),.I2(d_cnst_ss0_x),.I3(un1_df_1),.I4(d_cnst_sm0),.O(un87_df));
defparam desc266.INIT=32'h88F08800;
  LUT4_L desc267(.I0(\d_cnst_sn.g0_0_2 ),.I1(\d_cnst_sn.reg0_m9_i_a3_0 ),.I2(t_1[29:29]),.I3(\d_cnst_sn.g0_rn_1 ),.LO(reg0_28_10_2261_a6_3_2_lut6_2_RNIOK9O5));
defparam desc267.INIT=16'hFF02;
  LUT6 desc268(.I0(inf_abs0_2[23:23]),.I1(un36_df),.I2(N_1890),.I3(m7),.I4(un1_cf_x),.I5(un87_df),.O(\d_cnst_sn.reg3_17_sn_m7_0 ));
defparam desc268.INIT=64'h0000FFFEFFFEFFFE;
  LUT4 desc269(.I0(inf_abs0_2[23:23]),.I1(inf_abs0_2[20:20]),.I2(inf_abs0_2[21:21]),.I3(\d_cnst_sn.reg3_5_sqmuxa_2_1 ),.O(un1_cf_x));
defparam desc269.INIT=16'h0400;
  LUT3 desc270(.I0(inf_abs0_2[24:24]),.I1(inf_abs0_2[25:25]),.I2(inf_abs0_2[26:26]),.O(d_cnst_ss0_x));
defparam desc270.INIT=8'hBA;
  LUT6_L desc271(.I0(\d_cnst_sn.b64_0 ),.I1(\d_cnst_sn.b60_0 ),.I2(\d_cnst_sn.reg1_16_a0_1 [3:3]),.I3(\d_cnst_sn.reg0_1 [7:7]),.I4(t_1[7:7]),.I5(N_1042),.LO(reg0_28_7_rep1));
defparam desc271.INIT=64'h0F00FF0001001100;
  LUT6 desc272(.I0(datai[0:0]),.I1(inf_abs0_2_axb_30),.I2(inf_abs0_2[0:0]),.I3(inf_abs0_2_cry_29),.I4(inf_abs0_2[27:27]),.I5(inf_abs0_2[28:28]),.O(m_2_i[0:0]));
defparam desc272.INIT=64'h1D551D551D550F0F;
  LUT5_L desc273(.I0(\d_cnst_sn.reg0_m9_i_a3_0 ),.I1(N_1033),.I2(\d_cnst_sn.g0_1 ),.I3(un32_reg0_s_29),.I4(un11_reg0_s_29),.LO(\d_cnst_sn.g0_rn_1 ));
defparam desc273.INIT=32'hFAF8F2F0;
  LUT6 desc274(.I0(b),.I1(inf_abs0_2_axb_30),.I2(inf_abs0_2_cry_29),.I3(inf_abs0_2[24:24]),.I4(inf_abs0_2[25:25]),.I5(inf_abs0_2[26:26]),.O(un1_df_1));
defparam desc274.INIT=64'h2A3F2A1500000000;
  LUT5_L desc275(.I0(\d_cnst_sn.g0_0_2 ),.I1(\d_cnst_sn.reg0_m9_i_a3_0 ),.I2(\d_cnst_sn.g0_1 ),.I3(t_1[29:29]),.I4(\d_cnst_sn.g3 ),.LO(N_3569_rep1));
defparam desc275.INIT=32'hFCFEF0F2;
  LUT6_L desc276(.I0(\d_cnst_sn.reg0_28_2526_a5_1_0 ),.I1(\d_cnst_sn.reg1_16_8_1837_2_tz ),.I2(\d_cnst_sn.reg0_28_7_a0_0 [9:9]),.I3(\d_cnst_sn.reg0_28_0 [19:19]),.I4(t_1[19:19]),.I5(\d_cnst_sn.reg0_28_3_2492_1 ),.LO(N_3829_rep1));
defparam desc276.INIT=64'hFFFFFFFF0E00EE00;
  LUT6_L desc277(.I0(\d_cnst_sn.reg0_28_2526_a5_1_0 ),.I1(\d_cnst_sn.reg1_16_8_1837_2_tz ),.I2(\d_cnst_sn.reg0_28_7_a0_0 [9:9]),.I3(\d_cnst_sn.reg0_28_0 [20:20]),.I4(t_1[20:20]),.I5(\d_cnst_sn.reg0_28_4_2459_0 ),.LO(N_3803_rep1));
defparam desc277.INIT=64'hFFFFFFFF0E00EE00;
  LUT5_L desc278(.I0(\d_cnst_sn.reg0_28_7_a0_0 [9:9]),.I1(\d_cnst_sn.reg0_28_5_2426_3_1 ),.I2(\d_cnst_sn.reg0_28_5_2426_a6_1_1 ),.I3(t_1[21:21]),.I4(\d_cnst_sn.reg0_28_5_2426_0 ),.LO(N_3777_rep1));
defparam desc278.INIT=32'hFFFF54FC;
  LUT5_L desc279(.I0(\d_cnst_sn.reg0_28_7_a0_0 [9:9]),.I1(\d_cnst_sn.reg0_28_6_2393_3_1 ),.I2(\d_cnst_sn.reg0_28_6_2393_a6_1_1 ),.I3(t_1[22:22]),.I4(\d_cnst_sn.reg0_28_6_2393_0 ),.LO(N_3751_rep1));
defparam desc279.INIT=32'hFFFF54FC;
  LUT5_L desc280(.I0(\d_cnst_sn.reg0_28_7_a0_0 [9:9]),.I1(\d_cnst_sn.reg0_28_7_2360_3_1 ),.I2(\d_cnst_sn.reg0_28_7_2360_a6_1_1 ),.I3(t_1[23:23]),.I4(\d_cnst_sn.reg0_28_7_2360_0 ),.LO(N_3725_rep1));
defparam desc280.INIT=32'hFFFF54FC;
  LUT6_L desc281(.I0(\d_cnst_sn.reg1_16_8_1837_2_tz ),.I1(\d_cnst_sn.reg0_28_7_a0_0 [9:9]),.I2(reg0_28_7_d[24:24]),.I3(\d_cnst_sn.reg0_28_8_2327_a6_1_1 ),.I4(t_1[24:24]),.I5(\d_cnst_sn.reg0_28_8_2327_0 ),.LO(N_3699_rep1));
defparam desc281.INIT=64'hFFFFFFFF3320FFA8;
  LUT5_L desc282(.I0(\d_cnst_sn.reg0_28_7_a0_0 [9:9]),.I1(\d_cnst_sn.reg0_28_9_2294_3_1 ),.I2(\d_cnst_sn.reg0_28_9_2294_a6_1_1 ),.I3(t_1[25:25]),.I4(\d_cnst_sn.reg0_28_9_2294_0 ),.LO(N_3673_rep1));
defparam desc282.INIT=32'hFFFF54FC;
  LUT5_L desc283(.I0(\d_cnst_sn.reg0_28_7_a0_0 [9:9]),.I1(\d_cnst_sn.reg0_28_10_2261_a6_1_1 ),.I2(\d_cnst_sn.reg1_16_7_1870_3_1 ),.I3(t_1[26:26]),.I4(\d_cnst_sn.reg1_16_7_1870_0 ),.LO(N_3341_rep1));
defparam desc283.INIT=32'hFFFF54FC;
  LUT5_L desc284(.I0(inf_abs0_2[31:31]),.I1(\d_cnst_sn.reg0_28_14_2135_1_a0_2 ),.I2(reg3_1_1[30:30]),.I3(\d_cnst_sn.reg0_28_14_0 ),.I4(t_1[30:30]),.LO(N_3550_rep1));
defparam desc284.INIT=32'hFFA0FFEC;
  LUT5_L desc285(.I0(\d_cnst_sn.reg0_28_7_a0_0 [9:9]),.I1(\d_cnst_sn.reg0_28_11_2228_a6_1_1 ),.I2(\d_cnst_sn.reg1_16_8_1837_3_1 ),.I3(t_1[27:27]),.I4(\d_cnst_sn.reg1_16_8_1837_0 ),.LO(N_3315_rep1));
defparam desc285.INIT=32'hFFFF54FC;
  LUT6_L desc286(.I0(\d_cnst_sn.reg0_28_9_2294_a6_3_0 ),.I1(m_2[28:28]),.I2(\d_cnst_sn.reg0_28_7_a0_0 [9:9]),.I3(\d_cnst_sn.reg1_16_9_1804_3_tz ),.I4(t_1[28:28]),.I5(N_3614),.LO(N_3289_rep1));
defparam desc286.INIT=64'hFFFFFFFF8F88FF88;
  LUT6_L desc287(.I0(b),.I1(inf_abs0_2[27:27]),.I2(\d_cnst_sn.g0_3_a2_2 ),.I3(\d_cnst_sn.g0_3_1 ),.I4(t_1[31:31]),.I5(t_1[30:30]),.LO(N_3856_rep1));
defparam desc287.INIT=64'hFF00FF30FF40FF70;
  LUT6 desc288(.I0(inf_abs0_2[21:21]),.I1(inf_abs0_2[22:22]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[27:27]),.I4(inf_abs0_2[28:28]),.I5(\d_cnst_sn.g0_0_0_a5_0_0 ),.O(N_7_0));
defparam desc288.INIT=64'h0101010000000000;
  LUT6 desc289(.I0(inf_abs0_2[19:19]),.I1(inf_abs0_2[20:20]),.I2(inf_abs0_2[31:31]),.I3(N_7_0),.I4(\d_cnst_sn.reg1_16_a2_0 [5:5]),.I5(reg3_1_1[31:31]),.O(\d_cnst_sn.g0_0_0_1 ));
defparam desc289.INIT=64'hFFF1FF00FF00FF00;
  LUT6_L desc290(.I0(b),.I1(inf_abs0_2[27:27]),.I2(\d_cnst_sn.g0_0_0_a5_2 ),.I3(\d_cnst_sn.g0_0_0_1 ),.I4(t_1[31:31]),.I5(t_1[30:30]),.LO(reg2_16[31:31]));
defparam desc290.INIT=64'hFF00FF30FF40FF70;
  LUT3_L desc291(.I0(N_1033),.I1(un32_reg0_s_29),.I2(un11_reg0_s_29),.LO(\d_cnst_sn.g3 ));
defparam desc291.INIT=8'hE4;
  LUT5 desc292(.I0(b),.I1(inf_abs0_2[21:21]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[27:27]),.I4(inf_abs0_2[28:28]),.O(\d_cnst_sn.g0_0_2 ));
defparam desc292.INIT=32'h0000040C;
  LUT6 desc293(.I0(\d_cnst_sn.reg0_N_13_0 ),.I1(\d_cnst_sn.reg0_28_9_2294_a6_3_0 ),.I2(N_513_i),.I3(m_2[29:29]),.I4(reg0_m9_i_a1),.I5(reg3_1_1[29:29]),.O(\d_cnst_sn.g0_1 ));
defparam desc293.INIT=64'hFFFFCD05FFFFCC00;
  LUT6 desc294(.I0(datai[31:31]),.I1(inf_abs0_2[20:20]),.I2(inf_abs0_2[21:21]),.I3(inf_abs0_2[22:22]),.I4(inf_abs0_2[31:31]),.I5(N_7),.O(N_12));
defparam desc294.INIT=64'h0000000800000000;
  LUT6 desc295(.I0(inf_abs0_2[20:20]),.I1(inf_abs0_2[21:21]),.I2(inf_abs0_2[22:22]),.I3(inf_abs0_2[31:31]),.I4(N_12),.I5(reg3_1_1[31:31]),.O(\d_cnst_sn.g0_3_1 ));
defparam desc295.INIT=64'hFFFFFF01FFFF0000;
  LUT6_L desc296(.I0(b),.I1(inf_abs0_2[27:27]),.I2(\d_cnst_sn.g0_3_a2_2 ),.I3(\d_cnst_sn.g0_3_1 ),.I4(t_1[31:31]),.I5(t_1[30:30]),.LO(N_3856));
defparam desc296.INIT=64'hFF00FF30FF40FF70;
  LUT4 desc297(.I0(datai[28:28]),.I1(inf_abs0_2[27:27]),.I2(inf_abs0_2[28:28]),.I3(un1_cf),.O(N_1685));
defparam desc297.INIT=16'hA8AA;
  LUT4 desc298(.I0(datai[27:27]),.I1(inf_abs0_2[27:27]),.I2(inf_abs0_2[28:28]),.I3(un1_cf),.O(N_1684));
defparam desc298.INIT=16'hA8AA;
  LUT4 desc299(.I0(datai[26:26]),.I1(inf_abs0_2[27:27]),.I2(inf_abs0_2[28:28]),.I3(un1_cf),.O(N_1683));
defparam desc299.INIT=16'hA8AA;
  LUT4 desc300(.I0(datai[25:25]),.I1(inf_abs0_2[27:27]),.I2(inf_abs0_2[28:28]),.I3(un1_cf),.O(N_1682));
defparam desc300.INIT=16'hA8AA;
  LUT4_L desc301(.I0(datai[24:24]),.I1(inf_abs0_2[27:27]),.I2(inf_abs0_2[28:28]),.I3(un1_cf),.LO(N_1681));
defparam desc301.INIT=16'hA8AA;
  LUT4_L desc302(.I0(datai[23:23]),.I1(inf_abs0_2[27:27]),.I2(inf_abs0_2[28:28]),.I3(un1_cf),.LO(N_1680));
defparam desc302.INIT=16'hA8AA;
  LUT4_L desc303(.I0(datai[22:22]),.I1(inf_abs0_2[27:27]),.I2(inf_abs0_2[28:28]),.I3(un1_cf),.LO(N_1679));
defparam desc303.INIT=16'hA8AA;
  LUT4 desc304(.I0(datai[20:20]),.I1(inf_abs0_2[27:27]),.I2(inf_abs0_2[28:28]),.I3(un1_cf),.O(N_1677));
defparam desc304.INIT=16'hA8AA;
  LUT5 desc305(.I0(datai[7:7]),.I1(inf_abs0_2[7:7]),.I2(inf_abs0_2[27:27]),.I3(inf_abs0_2[28:28]),.I4(un1_cf),.O(N_1664));
defparam desc305.INIT=32'hAAACAAAA;
  LUT5 desc306(.I0(datai[6:6]),.I1(inf_abs0_2[6:6]),.I2(inf_abs0_2[27:27]),.I3(inf_abs0_2[28:28]),.I4(un1_cf),.O(N_1663));
defparam desc306.INIT=32'hAAACAAAA;
  LUT5_L desc307(.I0(datai[2:2]),.I1(inf_abs0_2[2:2]),.I2(inf_abs0_2[27:27]),.I3(inf_abs0_2[28:28]),.I4(un1_cf),.LO(N_1659));
defparam desc307.INIT=32'hAAACAAAA;
  LUT5 desc308(.I0(datai[9:9]),.I1(inf_abs0_2[9:9]),.I2(inf_abs0_2[27:27]),.I3(inf_abs0_2[28:28]),.I4(un1_cf),.O(N_1666));
defparam desc308.INIT=32'hAAACAAAA;
  LUT5 desc309(.I0(datai[11:11]),.I1(inf_abs0_2[11:11]),.I2(inf_abs0_2[27:27]),.I3(inf_abs0_2[28:28]),.I4(un1_cf),.O(N_1668));
defparam desc309.INIT=32'hAAACAAAA;
  LUT5 desc310(.I0(datai[10:10]),.I1(inf_abs0_2[10:10]),.I2(inf_abs0_2[27:27]),.I3(inf_abs0_2[28:28]),.I4(un1_cf),.O(N_1667));
defparam desc310.INIT=32'hAAACAAAA;
  LUT5 desc311(.I0(datai[17:17]),.I1(inf_abs0_2[17:17]),.I2(inf_abs0_2[27:27]),.I3(inf_abs0_2[28:28]),.I4(un1_cf),.O(N_1674));
defparam desc311.INIT=32'hAAACAAAA;
  LUT5 desc312(.I0(datai[12:12]),.I1(inf_abs0_2[12:12]),.I2(inf_abs0_2[27:27]),.I3(inf_abs0_2[28:28]),.I4(un1_cf),.O(N_1669));
defparam desc312.INIT=32'hAAACAAAA;
  LUT5 desc313(.I0(datai[18:18]),.I1(inf_abs0_2[18:18]),.I2(inf_abs0_2[27:27]),.I3(inf_abs0_2[28:28]),.I4(un1_cf),.O(N_1675));
defparam desc313.INIT=32'hAAACAAAA;
  LUT5 desc314(.I0(datai[14:14]),.I1(inf_abs0_2[14:14]),.I2(inf_abs0_2[27:27]),.I3(inf_abs0_2[28:28]),.I4(un1_cf),.O(N_1671));
defparam desc314.INIT=32'hAAACAAAA;
  LUT5 desc315(.I0(datai[19:19]),.I1(inf_abs0_2[19:19]),.I2(inf_abs0_2[27:27]),.I3(inf_abs0_2[28:28]),.I4(un1_cf),.O(N_1676));
defparam desc315.INIT=32'hAAACAAAA;
  LUT5 desc316(.I0(datai[13:13]),.I1(inf_abs0_2[13:13]),.I2(inf_abs0_2[27:27]),.I3(inf_abs0_2[28:28]),.I4(un1_cf),.O(N_1670));
defparam desc316.INIT=32'hAAACAAAA;
  LUT5_L desc317(.I0(datai[1:1]),.I1(inf_abs0_2[1:1]),.I2(inf_abs0_2[27:27]),.I3(inf_abs0_2[28:28]),.I4(un1_cf),.LO(N_1658));
defparam desc317.INIT=32'hAAACAAAA;
  LUT5 desc318(.I0(datai[16:16]),.I1(inf_abs0_2[16:16]),.I2(inf_abs0_2[27:27]),.I3(inf_abs0_2[28:28]),.I4(un1_cf),.O(N_1673));
defparam desc318.INIT=32'hAAACAAAA;
  LUT5 desc319(.I0(datai[15:15]),.I1(inf_abs0_2[15:15]),.I2(inf_abs0_2[27:27]),.I3(inf_abs0_2[28:28]),.I4(un1_cf),.O(N_1672));
defparam desc319.INIT=32'hAAACAAAA;
  LUT5 desc320(.I0(datai[8:8]),.I1(inf_abs0_2[8:8]),.I2(inf_abs0_2[27:27]),.I3(inf_abs0_2[28:28]),.I4(un1_cf),.O(N_1665));
defparam desc320.INIT=32'hAAACAAAA;
  LUT5 desc321(.I0(inf_abs0_2[23:23]),.I1(inf_abs0_2[20:20]),.I2(inf_abs0_2[21:21]),.I3(\d_cnst_sn.reg3_5_sqmuxa_2_1 ),.I4(un87_df),.O(un1_cf));
defparam desc321.INIT=32'h04000000;
  LUT5 desc322(.I0(inf_abs0_2[23:23]),.I1(inf_abs0_2[27:27]),.I2(inf_abs0_2[28:28]),.I3(un36_df),.I4(N_1890),.O(rd_4_sqmuxa));
defparam desc322.INIT=32'h00000001;
  LUT5 desc323(.I0(inf_abs0_2[23:23]),.I1(un1_b57),.I2(un1_df_17_2),.I3(un1_df_16),.I4(\d_cnst_sn.reg3_17_sn_m7_0 ),.O(N_1841));
defparam desc323.INIT=32'h00BF0000;
  LUT4 desc324(.I0(inf_abs0_2[23:23]),.I1(un36_df),.I2(un1_b59),.I3(un87_df),.O(un1_df_16));
defparam desc324.INIT=16'h1000;
  LUT5 desc325(.I0(inf_abs0_2[23:23]),.I1(un1_b57),.I2(un36_df),.I3(un1_b59),.I4(un87_df),.O(N_1810));
defparam desc325.INIT=32'hFAFBFFFF;
  LUT5_L desc326(.I0(inf_abs0_2[28:28]),.I1(inf_abs0_2[29:29]),.I2(N_933),.I3(N_965),.I4(reg3_14_sqmuxa),.LO(\d_cnst_sn.reg3_17_6_0 [19:19]));
defparam desc326.INIT=32'hFD75FFFF;
  LUT3_L desc327(.I0(inf_abs0_2[28:28]),.I1(reg3_14_sqmuxa),.I2(t_1[13:13]),.LO(reg3_17_4_a2[13:13]));
defparam desc327.INIT=8'h40;
  LUT5 desc328(.I0(inf_abs0_2[2:2]),.I1(inf_abs0_2[28:28]),.I2(r_4[1:1]),.I3(reg3_14_sqmuxa),.I4(t_1[2:2]),.O(N_1752));
defparam desc328.INIT=32'hC0AAF3AA;
  LUT5 desc329(.I0(inf_abs0_2[1:1]),.I1(inf_abs0_2[28:28]),.I2(r_4[0:0]),.I3(reg3_14_sqmuxa),.I4(t_1[1:1]),.O(N_1751));
defparam desc329.INIT=32'hC0AAF3AA;
  LUT4_L desc330(.I0(inf_abs0_2[0:0]),.I1(inf_abs0_2[28:28]),.I2(reg3_14_sqmuxa),.I3(t_1[0:0]),.LO(N_1750));
defparam desc330.INIT=16'h0A3A;
  LUT5 desc331(.I0(inf_abs0_2[28:28]),.I1(r_4[23:23]),.I2(\d_cnst_sn.reg3_17_sn_m7_0 ),.I3(reg3_14_sqmuxa),.I4(N_1681),.O(\d_cnst_sn.reg3_17_0_tz [24:24]));
defparam desc331.INIT=32'h8F0F8000;
  LUT5 desc332(.I0(inf_abs0_2[28:28]),.I1(r_4[21:21]),.I2(\d_cnst_sn.reg3_17_sn_m7_0 ),.I3(reg3_14_sqmuxa),.I4(N_1679),.O(\d_cnst_sn.reg3_17_0_tz [22:22]));
defparam desc332.INIT=32'h8F0F8000;
  LUT5 desc333(.I0(inf_abs0_2[28:28]),.I1(r_4[22:22]),.I2(\d_cnst_sn.reg3_17_sn_m7_0 ),.I3(reg3_14_sqmuxa),.I4(N_1680),.O(\d_cnst_sn.reg3_17_0_tz [23:23]));
defparam desc333.INIT=32'h8F0F8000;
  LUT5_L desc334(.I0(inf_abs0_2[17:17]),.I1(inf_abs0_2[28:28]),.I2(r_4[16:16]),.I3(rd_4_sqmuxa),.I4(reg3_14_sqmuxa),.LO(\d_cnst_sn.reg3_17_6_0 [17:17]));
defparam desc334.INIT=32'hF3F3AAFF;
  LUT5_L desc335(.I0(inf_abs0_2[16:16]),.I1(inf_abs0_2[28:28]),.I2(r_4[15:15]),.I3(rd_4_sqmuxa),.I4(reg3_14_sqmuxa),.LO(\d_cnst_sn.reg3_17_6_0 [16:16]));
defparam desc335.INIT=32'hF3F3AAFF;
  LUT5_L desc336(.I0(inf_abs0_2[14:14]),.I1(inf_abs0_2[28:28]),.I2(r_4[13:13]),.I3(rd_4_sqmuxa),.I4(reg3_14_sqmuxa),.LO(\d_cnst_sn.reg3_17_6_0 [14:14]));
defparam desc336.INIT=32'hF3F3AAFF;
  LUT5_L desc337(.I0(inf_abs0_2[15:15]),.I1(inf_abs0_2[28:28]),.I2(r_4[14:14]),.I3(rd_4_sqmuxa),.I4(reg3_14_sqmuxa),.LO(\d_cnst_sn.reg3_17_6_0 [15:15]));
defparam desc337.INIT=32'hF3F3AAFF;
  LUT5_L desc338(.I0(inf_abs0_2[12:12]),.I1(inf_abs0_2[28:28]),.I2(r_4[11:11]),.I3(rd_4_sqmuxa),.I4(reg3_14_sqmuxa),.LO(\d_cnst_sn.reg3_17_6_0 [12:12]));
defparam desc338.INIT=32'hF3F3AAFF;
  LUT5_L desc339(.I0(inf_abs0_2[13:13]),.I1(inf_abs0_2[28:28]),.I2(r_4[12:12]),.I3(rd_4_sqmuxa),.I4(reg3_14_sqmuxa),.LO(\d_cnst_sn.reg3_17_6_0 [13:13]));
defparam desc339.INIT=32'hF3F3AAFF;
  LUT5_L desc340(.I0(inf_abs0_2[18:18]),.I1(inf_abs0_2[28:28]),.I2(r_4[17:17]),.I3(rd_4_sqmuxa),.I4(reg3_14_sqmuxa),.LO(\d_cnst_sn.reg3_17_6_0 [18:18]));
defparam desc340.INIT=32'hF3F3AAFF;
  LUT2 desc341(.I0(inf_abs0_2[28:28]),.I1(reg3_14_sqmuxa),.O(\d_cnst_sn.reg3_17_a1_2 [24:24]));
defparam desc341.INIT=4'h4;
  LUT5 desc342(.I0(datai[4:4]),.I1(inf_abs0_2[4:4]),.I2(inf_abs0_2[27:27]),.I3(inf_abs0_2[28:28]),.I4(un1_cf),.O(N_1661));
defparam desc342.INIT=32'hAAACAAAA;
  LUT5_L desc343(.I0(datai[3:3]),.I1(inf_abs0_2[3:3]),.I2(inf_abs0_2[27:27]),.I3(inf_abs0_2[28:28]),.I4(un1_cf),.LO(N_1660));
defparam desc343.INIT=32'hAAACAAAA;
  LUT5 desc344(.I0(datai[5:5]),.I1(inf_abs0_2[5:5]),.I2(inf_abs0_2[27:27]),.I3(inf_abs0_2[28:28]),.I4(un1_cf),.O(N_1662));
defparam desc344.INIT=32'hAAACAAAA;
  LUT6 desc345(.I0(inf_abs0_2[21:21]),.I1(inf_abs0_2[22:22]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[28:28]),.I4(r_4[26:26]),.I5(reg3_1_1[27:27]),.O(\d_cnst_sn.reg1_16_8_1837_3_1 ));
defparam desc345.INIT=64'hF8F8F0F808080008;
  LUT6 desc346(.I0(inf_abs0_2[21:21]),.I1(inf_abs0_2[22:22]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[28:28]),.I4(r_4[25:25]),.I5(reg3_1_1[26:26]),.O(\d_cnst_sn.reg1_16_7_1870_3_1 ));
defparam desc346.INIT=64'hF8F8F0F808080008;
  LUT6 desc347(.I0(inf_abs0_2[21:21]),.I1(inf_abs0_2[22:22]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[28:28]),.I4(r_4[24:24]),.I5(reg3_1_1[25:25]),.O(\d_cnst_sn.reg0_28_9_2294_3_1 ));
defparam desc347.INIT=64'hF8F8F0F808080008;
  LUT6 desc348(.I0(inf_abs0_2[21:21]),.I1(inf_abs0_2[22:22]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[28:28]),.I4(r_4[22:22]),.I5(reg3_1_1[23:23]),.O(\d_cnst_sn.reg0_28_7_2360_3_1 ));
defparam desc348.INIT=64'hF8F8F0F808080008;
  LUT6 desc349(.I0(inf_abs0_2[21:21]),.I1(inf_abs0_2[22:22]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[28:28]),.I4(r_4[21:21]),.I5(reg3_1_1[22:22]),.O(\d_cnst_sn.reg0_28_6_2393_3_1 ));
defparam desc349.INIT=64'hF8F8F0F808080008;
  LUT6 desc350(.I0(inf_abs0_2[21:21]),.I1(inf_abs0_2[22:22]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[28:28]),.I4(r_4[20:20]),.I5(reg3_1_1[21:21]),.O(\d_cnst_sn.reg0_28_5_2426_3_1 ));
defparam desc350.INIT=64'hF8F8F0F808080008;
  LUT6 desc351(.I0(reg0[18:18]),.I1(reg2[18:18]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[29:29]),.I4(inf_abs0_2[30:30]),.I5(N_965),.O(r_4[18:18]));
defparam desc351.INIT=64'hAFACAFAAA0ACA0AA;
  LUT6 desc352(.I0(reg0[18:18]),.I1(reg2[18:18]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[29:29]),.I4(inf_abs0_2[30:30]),.I5(N_965),.O(un3_t_axb_18));
defparam desc352.INIT=64'h505350555F535F55;
  LUT6 desc353(.I0(reg0[21:21]),.I1(reg2[21:21]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[29:29]),.I4(inf_abs0_2[30:30]),.I5(N_968),.O(un3_t_axb_21));
defparam desc353.INIT=64'h505350555F535F55;
  LUT6 desc354(.I0(reg0[21:21]),.I1(reg2[21:21]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[29:29]),.I4(inf_abs0_2[30:30]),.I5(N_968),.O(r_4[21:21]));
defparam desc354.INIT=64'hAFACAFAAA0ACA0AA;
  LUT5 un32_reg0_axb_29_cZ(.I0(datai[29:29]),.I1(inf_abs0_2[31:31]),.I2(inf_abs0_2[27:27]),.I3(inf_abs0_2[28:28]),.I4(r_4[29:29]),.O(un32_reg0_axb_29));
defparam un32_reg0_axb_29_cZ.INIT=32'h2220DDDF;
  LUT6 desc355(.I0(inf_abs0_2[19:19]),.I1(inf_abs0_2[20:20]),.I2(inf_abs0_2[22:22]),.I3(inf_abs0_2[31:31]),.I4(m_2[30:30]),.I5(reg3_1_1[30:30]),.O(N_1493));
defparam desc355.INIT=64'hFF0DFF01000C0000;
  LUT6 desc356(.I0(un3_reg3_s_25),.I1(inf_abs0_2[19:19]),.I2(inf_abs0_2[20:20]),.I3(inf_abs0_2[31:31]),.I4(m_2[28:28]),.I5(reg3_1_1[28:28]),.O(N_1363));
defparam desc356.INIT=64'hFFFBFF0B00F80008;
  LUT6 desc357(.I0(un3_reg3_s_24),.I1(inf_abs0_2[19:19]),.I2(inf_abs0_2[20:20]),.I3(inf_abs0_2[31:31]),.I4(m_2[27:27]),.I5(reg3_1_1[27:27]),.O(N_1362));
defparam desc357.INIT=64'hFFFBFF0B00F80008;
  LUT6 desc358(.I0(un3_reg3_s_23),.I1(inf_abs0_2[19:19]),.I2(inf_abs0_2[20:20]),.I3(inf_abs0_2[31:31]),.I4(m_2[26:26]),.I5(reg3_1_1[26:26]),.O(N_1361));
defparam desc358.INIT=64'hFFFBFF0B00F80008;
  LUT6 desc359(.I0(un3_reg3_s_16),.I1(inf_abs0_2[19:19]),.I2(inf_abs0_2[20:20]),.I3(inf_abs0_2[31:31]),.I4(m_2[19:19]),.I5(reg3_1_1[19:19]),.O(N_1354));
defparam desc359.INIT=64'hFFFBFF0B00F80008;
  LUT6 desc360(.I0(un3_reg3_s_15),.I1(inf_abs0_2[19:19]),.I2(inf_abs0_2[20:20]),.I3(inf_abs0_2[31:31]),.I4(m_2[18:18]),.I5(reg3_1_1[18:18]),.O(N_1353));
defparam desc360.INIT=64'hFFFBFF0B00F80008;
  LUT6 desc361(.I0(un3_reg3_s_14),.I1(inf_abs0_2[19:19]),.I2(inf_abs0_2[20:20]),.I3(inf_abs0_2[31:31]),.I4(m_2[17:17]),.I5(reg3_1_1[17:17]),.O(N_1352));
defparam desc361.INIT=64'hFFFBFF0B00F80008;
  LUT6 desc362(.I0(un3_reg3_s_13),.I1(inf_abs0_2[19:19]),.I2(inf_abs0_2[20:20]),.I3(inf_abs0_2[31:31]),.I4(m_2[16:16]),.I5(reg3_1_1[16:16]),.O(N_1351));
defparam desc362.INIT=64'hFFFBFF0B00F80008;
  LUT6 desc363(.I0(un3_reg3_s_12),.I1(inf_abs0_2[19:19]),.I2(inf_abs0_2[20:20]),.I3(inf_abs0_2[31:31]),.I4(m_2[15:15]),.I5(reg3_1_1[15:15]),.O(N_1350));
defparam desc363.INIT=64'hFFFBFF0B00F80008;
  LUT6 desc364(.I0(un3_reg3_s_11),.I1(inf_abs0_2[19:19]),.I2(inf_abs0_2[20:20]),.I3(inf_abs0_2[31:31]),.I4(m_2[14:14]),.I5(reg3_1_1[14:14]),.O(N_1349));
defparam desc364.INIT=64'hFFFBFF0B00F80008;
  LUT6 desc365(.I0(un3_reg3_s_10),.I1(inf_abs0_2[19:19]),.I2(inf_abs0_2[20:20]),.I3(inf_abs0_2[31:31]),.I4(m_2[13:13]),.I5(reg3_1_1[13:13]),.O(N_1348));
defparam desc365.INIT=64'hFFFBFF0B00F80008;
  LUT6 desc366(.I0(un3_reg3_s_9),.I1(inf_abs0_2[19:19]),.I2(inf_abs0_2[20:20]),.I3(inf_abs0_2[31:31]),.I4(m_2[12:12]),.I5(reg3_1_1[12:12]),.O(N_1347));
defparam desc366.INIT=64'hFFFBFF0B00F80008;
  LUT6 desc367(.I0(un3_reg3_s_8),.I1(inf_abs0_2[19:19]),.I2(inf_abs0_2[20:20]),.I3(inf_abs0_2[31:31]),.I4(m_2[11:11]),.I5(reg3_1_1[11:11]),.O(N_1346));
defparam desc367.INIT=64'hFFFBFF0B00F80008;
  LUT6 desc368(.I0(un3_reg3_s_7),.I1(inf_abs0_2[19:19]),.I2(inf_abs0_2[20:20]),.I3(inf_abs0_2[31:31]),.I4(m_2[10:10]),.I5(reg3_1_1[10:10]),.O(N_1345));
defparam desc368.INIT=64'hFFFBFF0B00F80008;
  LUT6 desc369(.I0(un3_reg3_s_6),.I1(inf_abs0_2[19:19]),.I2(inf_abs0_2[20:20]),.I3(inf_abs0_2[31:31]),.I4(m_2[9:9]),.I5(reg3_1_1[9:9]),.O(N_1344));
defparam desc369.INIT=64'hFFFBFF0B00F80008;
  LUT6 desc370(.I0(un3_reg3_s_5),.I1(inf_abs0_2[19:19]),.I2(inf_abs0_2[20:20]),.I3(inf_abs0_2[31:31]),.I4(m_2[8:8]),.I5(reg3_1_1[8:8]),.O(N_1343));
defparam desc370.INIT=64'hFFFBFF0B00F80008;
  LUT6 desc371(.I0(un3_reg3_s_4),.I1(inf_abs0_2[19:19]),.I2(inf_abs0_2[20:20]),.I3(inf_abs0_2[31:31]),.I4(m_2[7:7]),.I5(reg3_1_1[7:7]),.O(N_1342));
defparam desc371.INIT=64'hFFFBFF0B00F80008;
  LUT6 desc372(.I0(un3_reg3_s_3),.I1(inf_abs0_2[19:19]),.I2(inf_abs0_2[20:20]),.I3(inf_abs0_2[31:31]),.I4(m_2[6:6]),.I5(reg3_1_1[6:6]),.O(N_1341));
defparam desc372.INIT=64'hFFFBFF0B00F80008;
  LUT6 desc373(.I0(un3_reg3_s_2),.I1(inf_abs0_2[19:19]),.I2(inf_abs0_2[20:20]),.I3(inf_abs0_2[31:31]),.I4(m_2[5:5]),.I5(reg3_1_1[5:5]),.O(N_1340));
defparam desc373.INIT=64'hFFFBFF0B00F80008;
  LUT6 desc374(.I0(un3_reg3_s_1),.I1(inf_abs0_2[19:19]),.I2(inf_abs0_2[20:20]),.I3(inf_abs0_2[31:31]),.I4(m_2[4:4]),.I5(reg3_1_1[4:4]),.O(N_1339));
defparam desc374.INIT=64'hFFFBFF0B00F80008;
  LUT6 desc375(.I0(reg3[3:3]),.I1(inf_abs0_2[19:19]),.I2(inf_abs0_2[20:20]),.I3(inf_abs0_2[31:31]),.I4(m_2[3:3]),.I5(reg3_1_1[3:3]),.O(N_1338));
defparam desc375.INIT=64'hFFF7FF0700F40004;
  LUT6 desc376(.I0(reg3[2:2]),.I1(inf_abs0_2[19:19]),.I2(inf_abs0_2[20:20]),.I3(inf_abs0_2[31:31]),.I4(m_2[2:2]),.I5(reg3_1_1[2:2]),.O(N_1337));
defparam desc376.INIT=64'hFFFBFF0B00F80008;
  LUT6 desc377(.I0(reg3[1:1]),.I1(inf_abs0_2[19:19]),.I2(inf_abs0_2[20:20]),.I3(inf_abs0_2[31:31]),.I4(m_2[1:1]),.I5(reg3_1_1[1:1]),.O(N_1336));
defparam desc377.INIT=64'hFFFBFF0B00F80008;
  LUT6 desc378(.I0(un3_reg3_s_22),.I1(inf_abs0_2[19:19]),.I2(inf_abs0_2[31:31]),.I3(\d_cnst_sn.reg0_28_a0_1 [7:7]),.I4(\d_cnst_sn.reg2_16_0 [25:25]),.I5(reg3_1_1[25:25]),.O(\d_cnst_sn.reg2_16_1 [25:25]));
defparam desc378.INIT=64'hFBFF000008FF0000;
  LUT6 desc379(.I0(un3_reg3_s_21),.I1(inf_abs0_2[19:19]),.I2(inf_abs0_2[31:31]),.I3(\d_cnst_sn.reg0_28_a0_1 [7:7]),.I4(\d_cnst_sn.reg2_16_0 [24:24]),.I5(reg3_1_1[24:24]),.O(\d_cnst_sn.reg2_16_1 [24:24]));
defparam desc379.INIT=64'hFBFF000008FF0000;
  LUT6 desc380(.I0(un3_reg3_s_20),.I1(inf_abs0_2[19:19]),.I2(inf_abs0_2[31:31]),.I3(\d_cnst_sn.reg0_28_a0_1 [7:7]),.I4(\d_cnst_sn.reg2_16_0 [23:23]),.I5(reg3_1_1[23:23]),.O(\d_cnst_sn.reg2_16_1 [23:23]));
defparam desc380.INIT=64'hFBFF000008FF0000;
  LUT6 desc381(.I0(un3_reg3_s_19),.I1(inf_abs0_2[19:19]),.I2(inf_abs0_2[31:31]),.I3(\d_cnst_sn.reg0_28_a0_1 [7:7]),.I4(\d_cnst_sn.reg2_16_0 [22:22]),.I5(reg3_1_1[22:22]),.O(\d_cnst_sn.reg2_16_1 [22:22]));
defparam desc381.INIT=64'hFBFF000008FF0000;
  LUT6 desc382(.I0(un3_reg3_s_18),.I1(inf_abs0_2[19:19]),.I2(inf_abs0_2[31:31]),.I3(\d_cnst_sn.reg0_28_a0_1 [7:7]),.I4(reg3_1_1[21:21]),.I5(\d_cnst_sn.reg2_16_0 [21:21]),.O(\d_cnst_sn.reg2_16_1 [21:21]));
defparam desc382.INIT=64'hFBFF08FF00000000;
  LUT6 desc383(.I0(inf_abs0_2[21:21]),.I1(inf_abs0_2[31:31]),.I2(inf_abs0_2[28:28]),.I3(r_4[15:15]),.I4(reg3_1_1[16:16]),.I5(t_1[16:16]),.O(N_1083));
defparam desc383.INIT=64'hFDDD2000FFDF2202;
  LUT6 desc384(.I0(inf_abs0_2[21:21]),.I1(inf_abs0_2[31:31]),.I2(inf_abs0_2[28:28]),.I3(r_4[14:14]),.I4(reg3_1_1[15:15]),.I5(t_1[15:15]),.O(N_1082));
defparam desc384.INIT=64'hFDDD2000FFDF2202;
  LUT6 desc385(.I0(inf_abs0_2[21:21]),.I1(inf_abs0_2[31:31]),.I2(inf_abs0_2[28:28]),.I3(r_4[13:13]),.I4(reg3_1_1[14:14]),.I5(t_1[14:14]),.O(N_1081));
defparam desc385.INIT=64'hFDDD2000FFDF2202;
  LUT6 desc386(.I0(inf_abs0_2[21:21]),.I1(inf_abs0_2[31:31]),.I2(inf_abs0_2[28:28]),.I3(r_4[12:12]),.I4(reg3_1_1[13:13]),.I5(t_1[13:13]),.O(N_1080));
defparam desc386.INIT=64'hFDDD2000FFDF2202;
  LUT6 desc387(.I0(inf_abs0_2[21:21]),.I1(inf_abs0_2[31:31]),.I2(inf_abs0_2[28:28]),.I3(r_4[11:11]),.I4(reg3_1_1[12:12]),.I5(t_1[12:12]),.O(N_1079));
defparam desc387.INIT=64'hFDDD2000FFDF2202;
  LUT6 desc388(.I0(inf_abs0_2[21:21]),.I1(inf_abs0_2[31:31]),.I2(inf_abs0_2[28:28]),.I3(r_4[10:10]),.I4(reg3_1_1[11:11]),.I5(t_1[11:11]),.O(N_1078));
defparam desc388.INIT=64'hFDDD2000FFDF2202;
  LUT6 desc389(.I0(inf_abs0_2[21:21]),.I1(inf_abs0_2[31:31]),.I2(inf_abs0_2[28:28]),.I3(r_4[9:9]),.I4(reg3_1_1[10:10]),.I5(t_1[10:10]),.O(N_1077));
defparam desc389.INIT=64'hFDDD2000FFDF2202;
  LUT6 desc390(.I0(inf_abs0_2[21:21]),.I1(inf_abs0_2[31:31]),.I2(inf_abs0_2[28:28]),.I3(r_4[8:8]),.I4(reg3_1_1[9:9]),.I5(t_1[9:9]),.O(N_1076));
defparam desc390.INIT=64'hFDDD2000FFDF2202;
  LUT6_L desc391(.I0(inf_abs0_2[21:21]),.I1(inf_abs0_2[31:31]),.I2(inf_abs0_2[28:28]),.I3(reg3_1_1[2:2]),.I4(r_4[1:1]),.I5(t_1[2:2]),.LO(N_1069));
defparam desc391.INIT=64'hFD20DD00FF22DF02;
  LUT6 desc392(.I0(inf_abs0_2[21:21]),.I1(inf_abs0_2[31:31]),.I2(inf_abs0_2[28:28]),.I3(reg3_1_1[1:1]),.I4(r_4[0:0]),.I5(t_1[1:1]),.O(N_1068));
defparam desc392.INIT=64'hFD20DD00FF22DF02;
  LUT6 desc393(.I0(inf_abs0_2[20:20]),.I1(inf_abs0_2[21:21]),.I2(inf_abs0_2[22:22]),.I3(inf_abs0_2[31:31]),.I4(N_3568),.I5(reg3_1_1[30:30]),.O(\d_cnst_sn.reg0_28_14_0 ));
defparam desc393.INIT=64'hFFFFC101FFFF0000;
  LUT6 desc394(.I0(reg1[4:4]),.I1(un3_reg3_s_1),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[29:29]),.I4(inf_abs0_2[30:30]),.I5(N_919),.O(r_4[4:4]));
defparam desc394.INIT=64'hFCFFFAFF0C000A00;
  LUT6 desc395(.I0(reg1[4:4]),.I1(un3_reg3_s_1),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[29:29]),.I4(inf_abs0_2[30:30]),.I5(N_919),.O(un3_t_axb_4));
defparam desc395.INIT=64'h03000500F3FFF5FF;
  LUT6 desc396(.I0(reg1[1:1]),.I1(reg3[1:1]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[29:29]),.I4(inf_abs0_2[30:30]),.I5(N_916),.O(un3_t_axb_1));
defparam desc396.INIT=64'h03000500F3FFF5FF;
  LUT6 desc397(.I0(reg1[1:1]),.I1(reg3[1:1]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[29:29]),.I4(inf_abs0_2[30:30]),.I5(N_916),.O(r_4[1:1]));
defparam desc397.INIT=64'hFCFFFAFF0C000A00;
  LUT6 desc398(.I0(reg1[0:0]),.I1(reg3[0:0]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[29:29]),.I4(inf_abs0_2[30:30]),.I5(N_915),.O(r_4[0:0]));
defparam desc398.INIT=64'hFCFFFAFF0C000A00;
  LUT6 desc399(.I0(reg1[0:0]),.I1(reg3[0:0]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[29:29]),.I4(inf_abs0_2[30:30]),.I5(N_915),.O(un3_t_axb_0));
defparam desc399.INIT=64'h03000500F3FFF5FF;
  LUT6 desc400(.I0(reg1[24:24]),.I1(un3_reg3_s_21),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[29:29]),.I4(inf_abs0_2[30:30]),.I5(N_939),.O(r_4[24:24]));
defparam desc400.INIT=64'hFCFFFAFF0C000A00;
  LUT6 desc401(.I0(reg1[24:24]),.I1(un3_reg3_s_21),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[29:29]),.I4(inf_abs0_2[30:30]),.I5(N_939),.O(un3_t_axb_24));
defparam desc401.INIT=64'h03000500F3FFF5FF;
  LUT6 desc402(.I0(reg1[23:23]),.I1(un3_reg3_s_20),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[29:29]),.I4(inf_abs0_2[30:30]),.I5(N_938),.O(r_4[23:23]));
defparam desc402.INIT=64'hFCFFFAFF0C000A00;
  LUT6 desc403(.I0(reg1[23:23]),.I1(un3_reg3_s_20),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[29:29]),.I4(inf_abs0_2[30:30]),.I5(N_938),.O(un3_t_axb_23));
defparam desc403.INIT=64'h03000500F3FFF5FF;
  LUT6 desc404(.I0(reg1[27:27]),.I1(un3_reg3_s_24),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[29:29]),.I4(inf_abs0_2[30:30]),.I5(N_942),.O(r_4[27:27]));
defparam desc404.INIT=64'hFCFFFAFF0C000A00;
  LUT6 desc405(.I0(reg1[27:27]),.I1(un3_reg3_s_24),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[29:29]),.I4(inf_abs0_2[30:30]),.I5(N_942),.O(un3_t_axb_27));
defparam desc405.INIT=64'h03000500F3FFF5FF;
  LUT6 desc406(.I0(reg1[20:20]),.I1(un3_reg3_s_17),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[29:29]),.I4(inf_abs0_2[30:30]),.I5(N_935),.O(r_4[20:20]));
defparam desc406.INIT=64'hFCFFFAFF0C000A00;
  LUT6 desc407(.I0(reg1[20:20]),.I1(un3_reg3_s_17),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[29:29]),.I4(inf_abs0_2[30:30]),.I5(N_935),.O(un3_t_axb_20));
defparam desc407.INIT=64'h03000500F3FFF5FF;
  LUT6 desc408(.I0(reg0[25:25]),.I1(reg2[25:25]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[29:29]),.I4(inf_abs0_2[30:30]),.I5(N_972),.O(r_4[25:25]));
defparam desc408.INIT=64'hAFACAFAAA0ACA0AA;
  LUT6 desc409(.I0(reg0[25:25]),.I1(reg2[25:25]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[29:29]),.I4(inf_abs0_2[30:30]),.I5(N_972),.O(un3_t_axb_25));
defparam desc409.INIT=64'h505350555F535F55;
  LUT6 desc410(.I0(reg0[28:28]),.I1(reg2[28:28]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[29:29]),.I4(inf_abs0_2[30:30]),.I5(N_975),.O(r_4[28:28]));
defparam desc410.INIT=64'hAFACAFAAA0ACA0AA;
  LUT6 desc411(.I0(reg0[28:28]),.I1(reg2[28:28]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[29:29]),.I4(inf_abs0_2[30:30]),.I5(N_975),.O(un3_t_axb_28));
defparam desc411.INIT=64'h505350555F535F55;
  LUT6 desc412(.I0(reg0[26:26]),.I1(reg2[26:26]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[29:29]),.I4(inf_abs0_2[30:30]),.I5(N_973),.O(r_4[26:26]));
defparam desc412.INIT=64'hAFACAFAAA0ACA0AA;
  LUT6 desc413(.I0(reg0[26:26]),.I1(reg2[26:26]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[29:29]),.I4(inf_abs0_2[30:30]),.I5(N_973),.O(un3_t_axb_26));
defparam desc413.INIT=64'h505350555F535F55;
  LUT6 desc414(.I0(reg1[22:22]),.I1(un3_reg3_s_19),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[29:29]),.I4(inf_abs0_2[30:30]),.I5(N_937),.O(un3_t_axb_22));
defparam desc414.INIT=64'h03000500F3FFF5FF;
  LUT6 desc415(.I0(reg1[22:22]),.I1(un3_reg3_s_19),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[29:29]),.I4(inf_abs0_2[30:30]),.I5(N_937),.O(r_4[22:22]));
defparam desc415.INIT=64'hFCFFFAFF0C000A00;
  LUT6 desc416(.I0(reg1[3:3]),.I1(reg3[3:3]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[29:29]),.I4(inf_abs0_2[30:30]),.I5(N_918),.O(r_4[3:3]));
defparam desc416.INIT=64'hF3FFFAFF03000A00;
  LUT6 desc417(.I0(reg1[3:3]),.I1(reg3[3:3]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[29:29]),.I4(inf_abs0_2[30:30]),.I5(N_918),.O(un3_t_axb_3));
defparam desc417.INIT=64'h0C000500FCFFF5FF;
  LUT5 desc418(.I0(inf_abs0_2[31:31]),.I1(inf_abs0_2[28:28]),.I2(inf_abs0_2[29:29]),.I3(N_967),.I4(N_935),.O(\d_cnst_sn.reg3_17_a2_2_0 [21:21]));
defparam desc418.INIT=32'h44044000;
  LUT5 desc419(.I0(inf_abs0_2[31:31]),.I1(inf_abs0_2[28:28]),.I2(inf_abs0_2[29:29]),.I3(N_941),.I4(N_973),.O(\d_cnst_sn.reg3_17_4_a2_0 [27:27]));
defparam desc419.INIT=32'h44400400;
  LUT5 desc420(.I0(inf_abs0_2[31:31]),.I1(inf_abs0_2[28:28]),.I2(inf_abs0_2[29:29]),.I3(N_971),.I4(N_939),.O(\d_cnst_sn.reg3_17_4_a2_0 [25:25]));
defparam desc420.INIT=32'h44044000;
  LUT5 desc421(.I0(inf_abs0_2[31:31]),.I1(inf_abs0_2[28:28]),.I2(inf_abs0_2[29:29]),.I3(N_974),.I4(N_942),.O(\d_cnst_sn.reg3_17_4_a2_0 [28:28]));
defparam desc421.INIT=32'h44044000;
  LUT5 desc422(.I0(inf_abs0_2[31:31]),.I1(inf_abs0_2[28:28]),.I2(inf_abs0_2[29:29]),.I3(N_940),.I4(N_972),.O(\d_cnst_sn.reg3_17_4_a2_0 [26:26]));
defparam desc422.INIT=32'h44400400;
  LUT6 desc423(.I0(inf_abs0_2[21:21]),.I1(inf_abs0_2[31:31]),.I2(inf_abs0_2[29:29]),.I3(N_970),.I4(N_938),.I5(reg3_1_1[24:24]),.O(reg0_28_7_d[24:24]));
defparam desc423.INIT=64'hFFDFFDDD22022000;
  LUT6 desc424(.I0(datai[26:26]),.I1(inf_abs0_2[31:31]),.I2(inf_abs0_2[29:29]),.I3(N_941),.I4(N_973),.I5(m7),.O(un32_reg0_axb_26));
defparam desc424.INIT=64'h00CF30FFAA659A55;
  LUT6 desc425(.I0(datai[25:25]),.I1(inf_abs0_2[31:31]),.I2(inf_abs0_2[29:29]),.I3(N_940),.I4(N_972),.I5(m7),.O(un32_reg0_axb_25));
defparam desc425.INIT=64'h00CF30FFAA659A55;
  LUT6 desc426(.I0(datai[23:23]),.I1(inf_abs0_2[31:31]),.I2(inf_abs0_2[29:29]),.I3(N_970),.I4(N_938),.I5(m7),.O(un32_reg0_axb_23));
defparam desc426.INIT=64'h0030CFFFAA9A6555;
  LUT6 desc427(.I0(inf_abs0_2[31:31]),.I1(inf_abs0_2[29:29]),.I2(r_4_2_a0[1:1]),.I3(\d_cnst_sn.r_4_0_0 [1:1]),.I4(N_916),.I5(m_2[1:1]),.O(un32_reg0_axb_1));
defparam desc427.INIT=64'hBFBB04004044FBFF;
  LUT6 desc428(.I0(inf_abs0_2[31:31]),.I1(inf_abs0_2[29:29]),.I2(m_2_i[0:0]),.I3(r_4_2_a0[0:0]),.I4(\d_cnst_sn.r_4_0_0 [0:0]),.I5(N_915),.O(N_1035));
defparam desc428.INIT=64'h4B0F4B4BF0B4F0F0;
  LUT6 desc429(.I0(datai[28:28]),.I1(inf_abs0_2[31:31]),.I2(inf_abs0_2[29:29]),.I3(N_943),.I4(N_975),.I5(m7),.O(un32_reg0_axb_28));
defparam desc429.INIT=64'h00CF30FFAA659A55;
  LUT6 desc430(.I0(datai[27:27]),.I1(inf_abs0_2[31:31]),.I2(inf_abs0_2[29:29]),.I3(N_974),.I4(N_942),.I5(m7),.O(un32_reg0_axb_27));
defparam desc430.INIT=64'h0030CFFFAA9A6555;
  LUT6 desc431(.I0(datai[20:20]),.I1(inf_abs0_2[31:31]),.I2(inf_abs0_2[29:29]),.I3(N_967),.I4(N_935),.I5(m7),.O(un32_reg0_axb_20));
defparam desc431.INIT=64'h0030CFFFAA9A6555;
  LUT6 desc432(.I0(datai[24:24]),.I1(inf_abs0_2[31:31]),.I2(inf_abs0_2[29:29]),.I3(N_971),.I4(N_939),.I5(m7),.O(un32_reg0_axb_24));
defparam desc432.INIT=64'h0030CFFFAA9A6555;
  LUT6 desc433(.I0(datai[22:22]),.I1(inf_abs0_2[31:31]),.I2(inf_abs0_2[29:29]),.I3(N_969),.I4(N_937),.I5(m7),.O(un32_reg0_axb_22));
defparam desc433.INIT=64'h0030CFFFAA9A6555;
  LUT6 desc434(.I0(datai[21:21]),.I1(inf_abs0_2[31:31]),.I2(inf_abs0_2[29:29]),.I3(N_936),.I4(N_968),.I5(m7),.O(un32_reg0_axb_21));
defparam desc434.INIT=64'h00CF30FFAA659A55;
  LUT5 desc435(.I0(state),.I1(inf_abs0_2[23:23]),.I2(inf_abs0_2[31:31]),.I3(un1_df_1),.I4(un36_df),.O(dce));
defparam desc435.INIT=32'h000000A2;
  LUT6 desc436(.I0(state),.I1(inf_abs0_2[23:23]),.I2(inf_abs0_2[31:31]),.I3(N_1892),.I4(un36_df),.I5(N_1890),.O(\d_cnst_sn.un1_state_3_1 ));
defparam desc436.INIT=64'hFFFFFF5DFFFFFFFF;
  LUT4 desc437(.I0(inf_abs0_2[31:31]),.I1(inf_abs0_2[28:28]),.I2(N_28),.I3(t_1[3:3]),.O(t_6[3:3]));
defparam desc437.INIT=16'h40FB;
  LUT6 desc438(.I0(inf_abs0_2[21:21]),.I1(inf_abs0_2[22:22]),.I2(inf_abs0_2[31:31]),.I3(N_1033),.I4(un32_reg0_s_28),.I5(un11_reg0_s_28),.O(N_3614));
defparam desc438.INIT=64'h0606060000060000;
  LUT5 un11_reg0_axb_29_cZ(.I0(datai[29:29]),.I1(inf_abs0_2[31:31]),.I2(inf_abs0_2[27:27]),.I3(inf_abs0_2[28:28]),.I4(r_4[29:29]),.O(un11_reg0_axb_29));
defparam un11_reg0_axb_29_cZ.INIT=32'hDDDF2220;
  LUT6 desc439(.I0(reg0[19:19]),.I1(reg2[19:19]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[29:29]),.I4(inf_abs0_2[30:30]),.I5(N_2722),.O(r_4[19:19]));
defparam desc439.INIT=64'hAFACAFAAA0ACA0AA;
  LUT6 desc440(.I0(reg0[19:19]),.I1(reg2[19:19]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[29:29]),.I4(inf_abs0_2[30:30]),.I5(N_2722),.O(un3_t_axb_19));
defparam desc440.INIT=64'h505350555F535F55;
  LUT6 desc441(.I0(reg0[6:6]),.I1(reg2[6:6]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[29:29]),.I4(inf_abs0_2[30:30]),.I5(N_953),.O(r_4[6:6]));
defparam desc441.INIT=64'hAFACAFAAA0ACA0AA;
  LUT6 desc442(.I0(reg0[6:6]),.I1(reg2[6:6]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[29:29]),.I4(inf_abs0_2[30:30]),.I5(N_953),.O(un3_t_axb_6));
defparam desc442.INIT=64'h505350555F535F55;
  LUT6 desc443(.I0(reg0[12:12]),.I1(reg2[12:12]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[29:29]),.I4(inf_abs0_2[30:30]),.I5(N_959),.O(un3_t_axb_12));
defparam desc443.INIT=64'h505350555F535F55;
  LUT6 desc444(.I0(reg0[12:12]),.I1(reg2[12:12]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[29:29]),.I4(inf_abs0_2[30:30]),.I5(N_959),.O(r_4[12:12]));
defparam desc444.INIT=64'hAFACAFAAA0ACA0AA;
  LUT6 desc445(.I0(reg0[5:5]),.I1(reg2[5:5]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[29:29]),.I4(inf_abs0_2[30:30]),.I5(N_952),.O(r_4[5:5]));
defparam desc445.INIT=64'hAFACAFAAA0ACA0AA;
  LUT6 desc446(.I0(reg0[5:5]),.I1(reg2[5:5]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[29:29]),.I4(inf_abs0_2[30:30]),.I5(N_952),.O(un3_t_axb_5));
defparam desc446.INIT=64'h505350555F535F55;
  LUT6 desc447(.I0(reg0[17:17]),.I1(reg2[17:17]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[29:29]),.I4(inf_abs0_2[30:30]),.I5(N_964),.O(r_4[17:17]));
defparam desc447.INIT=64'hAFACAFAAA0ACA0AA;
  LUT6 desc448(.I0(reg0[17:17]),.I1(reg2[17:17]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[29:29]),.I4(inf_abs0_2[30:30]),.I5(N_964),.O(un3_t_axb_17));
defparam desc448.INIT=64'h505350555F535F55;
  LUT6 desc449(.I0(reg0[7:7]),.I1(reg2[7:7]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[29:29]),.I4(inf_abs0_2[30:30]),.I5(N_954),.O(r_4[7:7]));
defparam desc449.INIT=64'hAFACAFAAA0ACA0AA;
  LUT6 desc450(.I0(reg0[7:7]),.I1(reg2[7:7]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[29:29]),.I4(inf_abs0_2[30:30]),.I5(N_954),.O(un3_t_axb_7));
defparam desc450.INIT=64'h505350555F535F55;
  LUT6 desc451(.I0(reg0[9:9]),.I1(reg2[9:9]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[29:29]),.I4(inf_abs0_2[30:30]),.I5(N_956),.O(r_4[9:9]));
defparam desc451.INIT=64'hAFACAFAAA0ACA0AA;
  LUT6 desc452(.I0(reg0[9:9]),.I1(reg2[9:9]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[29:29]),.I4(inf_abs0_2[30:30]),.I5(N_956),.O(un3_t_axb_9));
defparam desc452.INIT=64'h505350555F535F55;
  LUT6 desc453(.I0(reg0[10:10]),.I1(reg2[10:10]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[29:29]),.I4(inf_abs0_2[30:30]),.I5(N_957),.O(r_4[10:10]));
defparam desc453.INIT=64'hAFACAFAAA0ACA0AA;
  LUT6 desc454(.I0(reg0[10:10]),.I1(reg2[10:10]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[29:29]),.I4(inf_abs0_2[30:30]),.I5(N_957),.O(un3_t_axb_10));
defparam desc454.INIT=64'h505350555F535F55;
  LUT6 desc455(.I0(reg0[14:14]),.I1(reg2[14:14]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[29:29]),.I4(inf_abs0_2[30:30]),.I5(N_961),.O(un3_t_axb_14));
defparam desc455.INIT=64'h505350555F535F55;
  LUT6 desc456(.I0(reg0[14:14]),.I1(reg2[14:14]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[29:29]),.I4(inf_abs0_2[30:30]),.I5(N_961),.O(r_4[14:14]));
defparam desc456.INIT=64'hAFACAFAAA0ACA0AA;
  LUT6 desc457(.I0(reg0[16:16]),.I1(reg2[16:16]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[29:29]),.I4(inf_abs0_2[30:30]),.I5(N_963),.O(r_4[16:16]));
defparam desc457.INIT=64'hAFACAFAAA0ACA0AA;
  LUT6 desc458(.I0(reg0[16:16]),.I1(reg2[16:16]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[29:29]),.I4(inf_abs0_2[30:30]),.I5(N_963),.O(un3_t_axb_16));
defparam desc458.INIT=64'h505350555F535F55;
  LUT6 desc459(.I0(reg0[13:13]),.I1(reg2[13:13]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[29:29]),.I4(inf_abs0_2[30:30]),.I5(N_960),.O(r_4[13:13]));
defparam desc459.INIT=64'hAFACAFAAA0ACA0AA;
  LUT6 desc460(.I0(reg0[13:13]),.I1(reg2[13:13]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[29:29]),.I4(inf_abs0_2[30:30]),.I5(N_960),.O(un3_t_axb_13));
defparam desc460.INIT=64'h505350555F535F55;
  LUT6 desc461(.I0(reg0[11:11]),.I1(reg2[11:11]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[29:29]),.I4(inf_abs0_2[30:30]),.I5(N_958),.O(r_4[11:11]));
defparam desc461.INIT=64'hAFACAFAAA0ACA0AA;
  LUT6 desc462(.I0(reg0[11:11]),.I1(reg2[11:11]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[29:29]),.I4(inf_abs0_2[30:30]),.I5(N_958),.O(un3_t_axb_11));
defparam desc462.INIT=64'h505350555F535F55;
  LUT6 desc463(.I0(reg1[4:4]),.I1(inf_abs0_2[30:30]),.I2(\d_cnst_sn.r_4_0_0 [4:4]),.I3(N_919),.I4(m_2[4:4]),.I5(N_13),.O(un32_reg0_axb_4));
defparam desc463.INIT=64'hFF0000FFE0E01F1F;
  LUT6 desc464(.I0(reg0[15:15]),.I1(reg2[15:15]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[29:29]),.I4(inf_abs0_2[30:30]),.I5(N_962),.O(r_4[15:15]));
defparam desc464.INIT=64'hAFACAFAAA0ACA0AA;
  LUT6 desc465(.I0(reg0[15:15]),.I1(reg2[15:15]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[29:29]),.I4(inf_abs0_2[30:30]),.I5(N_962),.O(un3_t_axb_15));
defparam desc465.INIT=64'h505350555F535F55;
  LUT6_L desc466(.I0(state),.I1(un1_inf_abs0_10[1:1]),.I2(inf_abs0_2[27:27]),.I3(inf_abs0_2[28:28]),.I4(\d_cnst_sn.addr_20_iv_8_627_i_1 ),.I5(N_2641),.LO(N_2315_i));
defparam desc466.INIT=64'h000000000000DFFF;
  LUT6 desc467(.I0(reg0[8:8]),.I1(reg2[8:8]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[29:29]),.I4(inf_abs0_2[30:30]),.I5(N_955),.O(r_4[8:8]));
defparam desc467.INIT=64'hAFACAFAAA0ACA0AA;
  LUT6 desc468(.I0(reg0[8:8]),.I1(reg2[8:8]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[29:29]),.I4(inf_abs0_2[30:30]),.I5(N_955),.O(un3_t_axb_8));
defparam desc468.INIT=64'h505350555F535F55;
  LUT6_L desc469(.I0(reg2[0:0]),.I1(inf_abs0_2[0:0]),.I2(inf_abs0_2[28:28]),.I3(\d_cnst_sn.addr_20_iv_7_654_i_1 ),.I4(N_2660_2),.I5(N_2641),.LO(N_2335_i));
defparam desc469.INIT=64'h00000000006F00FF;
  LUT6 desc470(.I0(reg1[3:3]),.I1(inf_abs0_2[30:30]),.I2(\d_cnst_sn.r_4_0_0 [3:3]),.I3(N_918),.I4(m_2[3:3]),.I5(N_13),.O(un32_reg0_axb_3));
defparam desc470.INIT=64'hFF0000FFE0E01F1F;
  LUT6 desc471(.I0(datai[2:2]),.I1(inf_abs0_2[2:2]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[27:27]),.I4(inf_abs0_2[28:28]),.I5(N_28),.O(un32_reg0_axb_2));
defparam desc471.INIT=64'hCACACACC35353533;
  LUT4 desc472(.I0(inf_abs0_2[20:20]),.I1(inf_abs0_2[31:31]),.I2(un32_reg0_s_22),.I3(un11_reg0_s_22),.O(N_1581));
defparam desc472.INIT=16'hFD20;
  LUT6 un11_r_df22_cZ(.I0(N_969),.I1(N_937),.I2(m_2[22:22]),.I3(m_2[23:23]),.I4(N_13),.I5(r_4[23:23]),.O(un11_r_df22));
defparam un11_r_df22_cZ.INIT=64'hC300A50000C300A5;
  LUT6 un11_r_lt22_cZ(.I0(N_969),.I1(N_937),.I2(m_2[22:22]),.I3(m_2[23:23]),.I4(N_13),.I5(r_4[23:23]),.O(un11_r_lt22));
defparam un11_r_lt22_cZ.INIT=64'h30005000FF30FF50;
  LUT6 un26_r_lt22_cZ(.I0(N_969),.I1(N_937),.I2(m_2[22:22]),.I3(m_2[23:23]),.I4(N_13),.I5(r_4[23:23]),.O(un26_r_lt22));
defparam un26_r_lt22_cZ.INIT=64'h30005000FF30FF50;
  LUT6 un26_r_df22_cZ(.I0(N_969),.I1(N_937),.I2(m_2[22:22]),.I3(m_2[23:23]),.I4(N_13),.I5(r_4[23:23]),.O(un26_r_df22));
defparam un26_r_df22_cZ.INIT=64'hC300A50000C300A5;
  LUT6 b18_df22_cZ(.I0(N_969),.I1(N_937),.I2(m_2[22:22]),.I3(m_2[23:23]),.I4(N_13),.I5(r_4[23:23]),.O(b18_df22));
defparam b18_df22_cZ.INIT=64'hC300A50000C300A5;
  LUT6 b18_lt22_cZ(.I0(N_969),.I1(N_937),.I2(m_2[22:22]),.I3(m_2[23:23]),.I4(N_13),.I5(r_4[23:23]),.O(b18_lt22));
defparam b18_lt22_cZ.INIT=64'h0CFF0AFF000C000A;
  LUT4 desc473(.I0(inf_abs0_2[19:19]),.I1(inf_abs0_2[31:31]),.I2(un32_reg0_s_8),.I3(un11_reg0_s_8),.O(N_1375));
defparam desc473.INIT=16'hFD20;
  LUT4 desc474(.I0(inf_abs0_2[20:20]),.I1(inf_abs0_2[31:31]),.I2(un32_reg0_s_23),.I3(un11_reg0_s_23),.O(N_1582));
defparam desc474.INIT=16'hFD20;
  LUT4_L desc475(.I0(inf_abs0_2[20:20]),.I1(inf_abs0_2[31:31]),.I2(b18),.I3(un26_r_cry[30:30]),.LO(N_895));
defparam desc475.INIT=16'h2F0D;
  LUT4 desc476(.I0(inf_abs0_2[20:20]),.I1(inf_abs0_2[31:31]),.I2(un32_reg0_s_21),.I3(un11_reg0_s_21),.O(N_1580));
defparam desc476.INIT=16'hFD20;
  LUT4 desc477(.I0(inf_abs0_2[20:20]),.I1(inf_abs0_2[31:31]),.I2(un32_reg0_s_16),.I3(un11_reg0_s_16),.O(N_1575));
defparam desc477.INIT=16'hFD20;
  LUT4 desc478(.I0(inf_abs0_2[19:19]),.I1(inf_abs0_2[31:31]),.I2(un32_reg0_s_14),.I3(un11_reg0_s_14),.O(N_1381));
defparam desc478.INIT=16'hFD20;
  LUT4 desc479(.I0(inf_abs0_2[20:20]),.I1(inf_abs0_2[31:31]),.I2(un32_reg0_s_24),.I3(un11_reg0_s_24),.O(N_1583));
defparam desc479.INIT=16'hFD20;
  LUT6_L desc480(.I0(r_4_2_a0[1:1]),.I1(\d_cnst_sn.r_4_0_0 [1:1]),.I2(N_916),.I3(N_527_i),.I4(N_13),.I5(t_1[2:2]),.LO(t_6[2:2]));
defparam desc480.INIT=64'hF0004400F0FF44FF;
  LUT4 desc481(.I0(inf_abs0_2[19:19]),.I1(inf_abs0_2[31:31]),.I2(un11_reg0_s_2),.I3(un32_reg0_s_2),.O(N_1369));
defparam desc481.INIT=16'hF2D0;
  LUT6_L desc482(.I0(r_4_2_a1_lut6_2_O5[3:3]),.I1(\d_cnst_sn.r_4_0_0 [4:4]),.I2(N_919),.I3(N_527_i),.I4(N_13),.I5(t_1[5:5]),.LO(t_6[5:5]));
defparam desc482.INIT=64'hF0004400F0FF44FF;
  LUT6_L desc483(.I0(r_4_2_a1_lut6_2_O5[3:3]),.I1(\d_cnst_sn.r_4_0_0 [4:4]),.I2(N_919),.I3(N_527_i),.I4(N_13),.I5(t_1[5:5]),.LO(r_4_2_a1_lut6_2_RNI5V8R3[3:3]));
defparam desc483.INIT=64'h0FFFBBFF0F00BB00;
  LUT6_L desc484(.I0(reg1[19:19]),.I1(reg0[19:19]),.I2(reg2[19:19]),.I3(un3_reg3_s_16),.I4(inf_abs0_2[29:29]),.I5(inf_abs0_2[30:30]),.LO(N_2724));
defparam desc484.INIT=64'hFF00F0F0AAAACCCC;
  LUT6_L desc485(.I0(r_4_2_a1_lut6_2_O6[3:3]),.I1(\d_cnst_sn.r_4_0_0 [3:3]),.I2(N_918),.I3(N_527_i),.I4(N_13),.I5(t_1[4:4]),.LO(t_6[4:4]));
defparam desc485.INIT=64'hF0004400F0FF44FF;
  LUT6_L desc486(.I0(r_4_2_a1_lut6_2_O6[3:3]),.I1(\d_cnst_sn.r_4_0_0 [3:3]),.I2(N_918),.I3(N_527_i),.I4(N_13),.I5(t_1[4:4]),.LO(r_4_2_a1_lut6_2_RNI2T8R3[3:3]));
defparam desc486.INIT=64'h0FFFBBFF0F00BB00;
  LUT6 desc487(.I0(inf_abs0_2[19:19]),.I1(inf_abs0_2[20:20]),.I2(inf_abs0_2[21:21]),.I3(inf_abs0_2[31:31]),.I4(un32_reg0_s_8),.I5(un11_reg0_s_8),.O(N_1043));
defparam desc487.INIT=64'hFFFFFF3500CA0000;
  LUT6 un11_r_df20_cZ(.I0(N_967),.I1(N_935),.I2(m_2[20:20]),.I3(m_2[21:21]),.I4(N_13),.I5(r_4[21:21]),.O(un11_r_df20));
defparam un11_r_df20_cZ.INIT=64'hC300A50000C300A5;
  LUT6 un11_r_lt20_cZ(.I0(N_967),.I1(N_935),.I2(m_2[20:20]),.I3(m_2[21:21]),.I4(N_13),.I5(r_4[21:21]),.O(un11_r_lt20));
defparam un11_r_lt20_cZ.INIT=64'h30005000FF30FF50;
  LUT6 un26_r_df20_cZ(.I0(N_967),.I1(N_935),.I2(m_2[20:20]),.I3(m_2[21:21]),.I4(N_13),.I5(r_4[21:21]),.O(un26_r_df20));
defparam un26_r_df20_cZ.INIT=64'hC300A50000C300A5;
  LUT6 un26_r_lt20_cZ(.I0(N_967),.I1(N_935),.I2(m_2[20:20]),.I3(m_2[21:21]),.I4(N_13),.I5(r_4[21:21]),.O(un26_r_lt20));
defparam un26_r_lt20_cZ.INIT=64'h30005000FF30FF50;
  LUT6 b18_df20_cZ(.I0(N_967),.I1(N_935),.I2(m_2[20:20]),.I3(m_2[21:21]),.I4(N_13),.I5(r_4[21:21]),.O(b18_df20));
defparam b18_df20_cZ.INIT=64'hC300A50000C300A5;
  LUT6 b18_lt20_cZ(.I0(N_967),.I1(N_935),.I2(m_2[20:20]),.I3(m_2[21:21]),.I4(N_13),.I5(r_4[21:21]),.O(b18_lt20));
defparam b18_lt20_cZ.INIT=64'h0CFF0AFF000C000A;
  LUT4 desc488(.I0(inf_abs0_2[19:19]),.I1(inf_abs0_2[31:31]),.I2(un32_reg0_s_12),.I3(un11_reg0_s_12),.O(N_1379));
defparam desc488.INIT=16'hFD20;
  LUT6_L desc489(.I0(N_513_i),.I1(m_2[0:0]),.I2(N_527_i),.I3(N_3916),.I4(N_1035),.I5(t_1[0:0]),.LO(reg1_16[0:0]));
defparam desc489.INIT=64'h0044FF44004EFF4E;
  LUT6_L desc490(.I0(N_513_i),.I1(m_2[0:0]),.I2(N_527_i),.I3(N_3916),.I4(N_1035),.I5(t_1[0:0]),.LO(reg0_28[0:0]));
defparam desc490.INIT=64'h0044FF44004EFF4E;
  LUT4 desc491(.I0(inf_abs0_2[20:20]),.I1(inf_abs0_2[31:31]),.I2(un32_reg0_s_15),.I3(un11_reg0_s_15),.O(N_1574));
defparam desc491.INIT=16'hFD20;
  LUT6 desc492(.I0(inf_abs0_2[19:19]),.I1(inf_abs0_2[20:20]),.I2(inf_abs0_2[21:21]),.I3(inf_abs0_2[31:31]),.I4(un32_reg0_s_7),.I5(un11_reg0_s_7),.O(N_1042));
defparam desc492.INIT=64'hFFFFFF3500CA0000;
  LUT6 desc493(.I0(inf_abs0_2[19:19]),.I1(inf_abs0_2[20:20]),.I2(inf_abs0_2[21:21]),.I3(inf_abs0_2[31:31]),.I4(un32_reg0_s_11),.I5(un11_reg0_s_11),.O(N_1046));
defparam desc493.INIT=64'hFFFFFF3500CA0000;
  LUT4 desc494(.I0(inf_abs0_2[19:19]),.I1(inf_abs0_2[31:31]),.I2(un32_reg0_s_13),.I3(un11_reg0_s_13),.O(N_1380));
defparam desc494.INIT=16'hFD20;
  LUT6 desc495(.I0(inf_abs0_2[19:19]),.I1(inf_abs0_2[20:20]),.I2(inf_abs0_2[21:21]),.I3(inf_abs0_2[31:31]),.I4(un32_reg0_s_13),.I5(un11_reg0_s_13),.O(N_1048));
defparam desc495.INIT=64'hFFFFFF3500CA0000;
  LUT4 desc496(.I0(inf_abs0_2[19:19]),.I1(inf_abs0_2[31:31]),.I2(un32_reg0_s_11),.I3(un11_reg0_s_11),.O(N_1378));
defparam desc496.INIT=16'hFD20;
  LUT4 desc497(.I0(inf_abs0_2[19:19]),.I1(inf_abs0_2[31:31]),.I2(un32_reg0_s_10),.I3(un11_reg0_s_10),.O(N_1377));
defparam desc497.INIT=16'hFD20;
  LUT4 desc498(.I0(inf_abs0_2[19:19]),.I1(inf_abs0_2[31:31]),.I2(un32_reg0_s_9),.I3(un11_reg0_s_9),.O(N_1376));
defparam desc498.INIT=16'hFD20;
  LUT4 desc499(.I0(inf_abs0_2[19:19]),.I1(inf_abs0_2[31:31]),.I2(un32_reg0_s_6),.I3(un11_reg0_s_6),.O(N_1373));
defparam desc499.INIT=16'hFD20;
  LUT4 desc500(.I0(inf_abs0_2[19:19]),.I1(inf_abs0_2[31:31]),.I2(un32_reg0_s_3),.I3(un11_reg0_s_3),.O(N_1370));
defparam desc500.INIT=16'hFD20;
  LUT4 desc501(.I0(inf_abs0_2[19:19]),.I1(inf_abs0_2[31:31]),.I2(un11_reg0_s_1),.I3(un32_reg0_s_1),.O(N_1368));
defparam desc501.INIT=16'hF2D0;
  LUT6 un11_r_df28_cZ(.I0(N_943),.I1(N_975),.I2(m_2[29:29]),.I3(m_2[28:28]),.I4(N_13),.I5(r_4[29:29]),.O(un11_r_df28));
defparam un11_r_df28_cZ.INIT=64'hA050C0300A050C03;
  LUT6 un11_r_lt28_cZ(.I0(N_943),.I1(N_975),.I2(m_2[29:29]),.I3(m_2[28:28]),.I4(N_13),.I5(r_4[29:29]),.O(un11_r_lt28));
defparam un11_r_lt28_cZ.INIT=64'h50003000F5F0F3F0;
  LUT6 un26_r_df28_cZ(.I0(N_943),.I1(N_975),.I2(m_2[29:29]),.I3(m_2[28:28]),.I4(N_13),.I5(r_4[29:29]),.O(un26_r_df28));
defparam un26_r_df28_cZ.INIT=64'hA050C0300A050C03;
  LUT6 un26_r_lt28_cZ(.I0(N_943),.I1(N_975),.I2(m_2[29:29]),.I3(m_2[28:28]),.I4(N_13),.I5(r_4[29:29]),.O(un26_r_lt28));
defparam un26_r_lt28_cZ.INIT=64'h50003000F5F0F3F0;
  LUT6 b18_df28_cZ(.I0(N_943),.I1(N_975),.I2(m_2[29:29]),.I3(m_2[28:28]),.I4(N_13),.I5(r_4[29:29]),.O(b18_df28));
defparam b18_df28_cZ.INIT=64'hA050C0300A050C03;
  LUT6 b18_lt28_cZ(.I0(N_943),.I1(N_975),.I2(m_2[29:29]),.I3(m_2[28:28]),.I4(N_13),.I5(r_4[29:29]),.O(b18_lt28));
defparam b18_lt28_cZ.INIT=64'h0FAF0FCF000A000C;
  LUT6 un11_r_df26_cZ(.I0(N_941),.I1(N_973),.I2(m_2[26:26]),.I3(m_2[27:27]),.I4(N_13),.I5(r_4[27:27]),.O(un11_r_df26));
defparam un11_r_df26_cZ.INIT=64'hA500C30000A500C3;
  LUT6 un11_r_lt26_cZ(.I0(N_941),.I1(N_973),.I2(m_2[26:26]),.I3(m_2[27:27]),.I4(N_13),.I5(r_4[27:27]),.O(un11_r_lt26));
defparam un11_r_lt26_cZ.INIT=64'h50003000FF50FF30;
  LUT6 b18_df26_cZ(.I0(N_941),.I1(N_973),.I2(m_2[26:26]),.I3(m_2[27:27]),.I4(N_13),.I5(r_4[27:27]),.O(b18_df26));
defparam b18_df26_cZ.INIT=64'hA500C30000A500C3;
  LUT6 un26_r_df26_cZ(.I0(N_941),.I1(N_973),.I2(m_2[26:26]),.I3(m_2[27:27]),.I4(N_13),.I5(r_4[27:27]),.O(un26_r_df26));
defparam un26_r_df26_cZ.INIT=64'hA500C30000A500C3;
  LUT6 un26_r_lt26_cZ(.I0(N_941),.I1(N_973),.I2(m_2[26:26]),.I3(m_2[27:27]),.I4(N_13),.I5(r_4[27:27]),.O(un26_r_lt26));
defparam un26_r_lt26_cZ.INIT=64'h50003000FF50FF30;
  LUT6 b18_lt26_cZ(.I0(N_941),.I1(N_973),.I2(m_2[26:26]),.I3(m_2[27:27]),.I4(N_13),.I5(r_4[27:27]),.O(b18_lt26));
defparam b18_lt26_cZ.INIT=64'h0AFF0CFF000A000C;
  LUT6 un11_r_lt24_cZ(.I0(N_940),.I1(N_972),.I2(m_2[24:24]),.I3(m_2[25:25]),.I4(N_13),.I5(r_4[24:24]),.O(un11_r_lt24));
defparam un11_r_lt24_cZ.INIT=64'h55003300F550F330;
  LUT6 un11_r_df24_cZ(.I0(N_940),.I1(N_972),.I2(m_2[24:24]),.I3(m_2[25:25]),.I4(N_13),.I5(r_4[24:24]),.O(un11_r_df24));
defparam un11_r_df24_cZ.INIT=64'hA050C0300A050C03;
  LUT6 b18_df24_cZ(.I0(N_940),.I1(N_972),.I2(m_2[24:24]),.I3(m_2[25:25]),.I4(N_13),.I5(r_4[24:24]),.O(b18_df24));
defparam b18_df24_cZ.INIT=64'hA050C0300A050C03;
  LUT6 b18_lt24_cZ(.I0(N_940),.I1(N_972),.I2(m_2[24:24]),.I3(m_2[25:25]),.I4(N_13),.I5(r_4[24:24]),.O(b18_lt24));
defparam b18_lt24_cZ.INIT=64'h0AAF0CCF00AA00CC;
  LUT6 un26_r_df24_cZ(.I0(N_940),.I1(N_972),.I2(m_2[24:24]),.I3(m_2[25:25]),.I4(N_13),.I5(r_4[24:24]),.O(un26_r_df24));
defparam un26_r_df24_cZ.INIT=64'hA050C0300A050C03;
  LUT6 un26_r_lt24_cZ(.I0(N_940),.I1(N_972),.I2(m_2[24:24]),.I3(m_2[25:25]),.I4(N_13),.I5(r_4[24:24]),.O(un26_r_lt24));
defparam un26_r_lt24_cZ.INIT=64'h55003300F550F330;
  LUT6_L desc502(.I0(r_4_2_a0[0:0]),.I1(\d_cnst_sn.r_4_0_0 [0:0]),.I2(N_915),.I3(N_527_i),.I4(N_13),.I5(t_1[1:1]),.LO(t_6[1:1]));
defparam desc502.INIT=64'hF0004400F0FF44FF;
  LUT6 desc503(.I0(inf_abs0_2[19:19]),.I1(inf_abs0_2[20:20]),.I2(inf_abs0_2[21:21]),.I3(inf_abs0_2[31:31]),.I4(un32_reg0_s_9),.I5(un11_reg0_s_9),.O(N_1044));
defparam desc503.INIT=64'hFFFFFF3500CA0000;
  LUT6 desc504(.I0(inf_abs0_2[19:19]),.I1(inf_abs0_2[20:20]),.I2(inf_abs0_2[21:21]),.I3(inf_abs0_2[31:31]),.I4(un11_reg0_s_1),.I5(un32_reg0_s_1),.O(N_1036));
defparam desc504.INIT=64'hFFFF00CAFF350000;
  LUT6 desc505(.I0(inf_abs0_2[19:19]),.I1(inf_abs0_2[20:20]),.I2(inf_abs0_2[21:21]),.I3(inf_abs0_2[31:31]),.I4(un11_reg0_s_2),.I5(un32_reg0_s_2),.O(N_1037));
defparam desc505.INIT=64'hFFFF00CAFF350000;
  LUT6 desc506(.I0(inf_abs0_2[19:19]),.I1(inf_abs0_2[20:20]),.I2(inf_abs0_2[21:21]),.I3(inf_abs0_2[31:31]),.I4(un32_reg0_s_6),.I5(un11_reg0_s_6),.O(N_1041));
defparam desc506.INIT=64'hFFFFFF3500CA0000;
  LUT6 desc507(.I0(inf_abs0_2[19:19]),.I1(inf_abs0_2[21:21]),.I2(inf_abs0_2[22:22]),.I3(inf_abs0_2[31:31]),.I4(un32_reg0_s_22),.I5(un11_reg0_s_22),.O(reg2_16_11_a4[22:22]));
defparam desc507.INIT=64'h0000002000100030;
  LUT6 desc508(.I0(inf_abs0_2[19:19]),.I1(inf_abs0_2[21:21]),.I2(inf_abs0_2[22:22]),.I3(inf_abs0_2[31:31]),.I4(un32_reg0_s_21),.I5(un11_reg0_s_21),.O(reg2_16_11_a4[21:21]));
defparam desc508.INIT=64'h0000002000100030;
  LUT6 desc509(.I0(inf_abs0_2[20:20]),.I1(inf_abs0_2[21:21]),.I2(inf_abs0_2[22:22]),.I3(inf_abs0_2[31:31]),.I4(un32_reg0_s_17),.I5(un11_reg0_s_17),.O(reg2_16_11_a2[17:17]));
defparam desc509.INIT=64'h000000080004000C;
  LUT6 desc510(.I0(inf_abs0_2[19:19]),.I1(inf_abs0_2[20:20]),.I2(inf_abs0_2[21:21]),.I3(inf_abs0_2[22:22]),.I4(inf_abs0_2[31:31]),.I5(un32_reg0_s_20),.O(\d_cnst_sn.reg2_16_1 [20:20]));
defparam desc510.INIT=64'hFFFFFFFFFFFFF53F;
  LUT4 desc511(.I0(inf_abs0_2[20:20]),.I1(inf_abs0_2[31:31]),.I2(un32_reg0_s_14),.I3(un11_reg0_s_14),.O(N_1573));
defparam desc511.INIT=16'hFD20;
  LUT4 desc512(.I0(inf_abs0_2[20:20]),.I1(inf_abs0_2[31:31]),.I2(un32_reg0_s_13),.I3(un11_reg0_s_13),.O(N_1572));
defparam desc512.INIT=16'hFD20;
  LUT4 desc513(.I0(inf_abs0_2[20:20]),.I1(inf_abs0_2[31:31]),.I2(un32_reg0_s_12),.I3(un11_reg0_s_12),.O(N_1571));
defparam desc513.INIT=16'hFD20;
  LUT4 desc514(.I0(inf_abs0_2[20:20]),.I1(inf_abs0_2[31:31]),.I2(un32_reg0_s_11),.I3(un11_reg0_s_11),.O(N_1570));
defparam desc514.INIT=16'hFD20;
  LUT4 desc515(.I0(inf_abs0_2[20:20]),.I1(inf_abs0_2[31:31]),.I2(un32_reg0_s_10),.I3(un11_reg0_s_10),.O(N_1569));
defparam desc515.INIT=16'hFD20;
  LUT5 desc516(.I0(state),.I1(inf_abs0_2[27:27]),.I2(inf_abs0_2[28:28]),.I3(un1_inf_abs0_10[7:7]),.I4(un1_inf_abs0_11[7:7]),.O(\d_cnst_sn.addr_20_iv_14_443_i_2 ));
defparam desc516.INIT=32'h008022A2;
  LUT4 desc517(.I0(inf_abs0_2[19:19]),.I1(inf_abs0_2[31:31]),.I2(un32_reg0_s_15),.I3(un11_reg0_s_15),.O(N_1382));
defparam desc517.INIT=16'hFD20;
  LUT6 desc518(.I0(inf_abs0_2[19:19]),.I1(inf_abs0_2[21:21]),.I2(inf_abs0_2[22:22]),.I3(inf_abs0_2[31:31]),.I4(un32_reg0_s_25),.I5(un11_reg0_s_25),.O(reg2_16_11_a4[25:25]));
defparam desc518.INIT=64'h0000002000100030;
  LUT4 desc519(.I0(inf_abs0_2[19:19]),.I1(inf_abs0_2[31:31]),.I2(un32_reg0_s_5),.I3(un11_reg0_s_5),.O(N_1372));
defparam desc519.INIT=16'hFD20;
  LUT6 desc520(.I0(inf_abs0_2[19:19]),.I1(inf_abs0_2[20:20]),.I2(inf_abs0_2[21:21]),.I3(inf_abs0_2[31:31]),.I4(un32_reg0_s_16),.I5(un11_reg0_s_16),.O(N_1051));
defparam desc520.INIT=64'hFFFFFF3500CA0000;
  LUT4 desc521(.I0(inf_abs0_2[19:19]),.I1(inf_abs0_2[31:31]),.I2(un32_reg0_s_4),.I3(un11_reg0_s_4),.O(N_1371));
defparam desc521.INIT=16'hFD20;
  LUT6 desc522(.I0(inf_abs0_2[19:19]),.I1(inf_abs0_2[20:20]),.I2(inf_abs0_2[21:21]),.I3(inf_abs0_2[31:31]),.I4(un32_reg0_s_15),.I5(un11_reg0_s_15),.O(N_1050));
defparam desc522.INIT=64'hFFFFFF3500CA0000;
  LUT6 desc523(.I0(inf_abs0_2[19:19]),.I1(inf_abs0_2[20:20]),.I2(inf_abs0_2[21:21]),.I3(inf_abs0_2[31:31]),.I4(un32_reg0_s_17),.I5(un11_reg0_s_17),.O(N_1052));
defparam desc523.INIT=64'hFFFFFF3500CA0000;
  LUT4 desc524(.I0(inf_abs0_2[19:19]),.I1(inf_abs0_2[31:31]),.I2(un32_reg0_s_16),.I3(un11_reg0_s_16),.O(N_1383));
defparam desc524.INIT=16'hFD20;
  LUT6 desc525(.I0(inf_abs0_2[19:19]),.I1(inf_abs0_2[21:21]),.I2(inf_abs0_2[22:22]),.I3(inf_abs0_2[31:31]),.I4(un32_reg0_s_29),.I5(un11_reg0_s_29),.O(reg2_16_11_a3[29:29]));
defparam desc525.INIT=64'h0030001000200000;
  LUT6 desc526(.I0(inf_abs0_2[19:19]),.I1(inf_abs0_2[21:21]),.I2(inf_abs0_2[22:22]),.I3(inf_abs0_2[31:31]),.I4(un32_reg0_s_24),.I5(un11_reg0_s_24),.O(reg2_16_11_a4[24:24]));
defparam desc526.INIT=64'h0000002000100030;
  LUT6 desc527(.I0(inf_abs0_2[20:20]),.I1(inf_abs0_2[21:21]),.I2(inf_abs0_2[22:22]),.I3(inf_abs0_2[31:31]),.I4(un32_reg0_s_18),.I5(un11_reg0_s_18),.O(reg2_16_11_a2[18:18]));
defparam desc527.INIT=64'h000000080004000C;
  LUT4 desc528(.I0(inf_abs0_2[20:20]),.I1(inf_abs0_2[31:31]),.I2(un32_reg0_s_5),.I3(un11_reg0_s_5),.O(N_1564));
defparam desc528.INIT=16'hFD20;
  LUT6 desc529(.I0(inf_abs0_2[19:19]),.I1(inf_abs0_2[20:20]),.I2(inf_abs0_2[21:21]),.I3(inf_abs0_2[31:31]),.I4(un32_reg0_s_10),.I5(un11_reg0_s_10),.O(N_1045));
defparam desc529.INIT=64'hFFFFFF3500CA0000;
  LUT6 desc530(.I0(inf_abs0_2[19:19]),.I1(inf_abs0_2[20:20]),.I2(inf_abs0_2[21:21]),.I3(inf_abs0_2[31:31]),.I4(un32_reg0_s_14),.I5(un11_reg0_s_14),.O(N_1049));
defparam desc530.INIT=64'hFFFFFF3500CA0000;
  LUT4 desc531(.I0(inf_abs0_2[20:20]),.I1(inf_abs0_2[31:31]),.I2(un32_reg0_s_9),.I3(un11_reg0_s_9),.O(N_1568));
defparam desc531.INIT=16'hFD20;
  LUT6 desc532(.I0(inf_abs0_2[20:20]),.I1(inf_abs0_2[21:21]),.I2(inf_abs0_2[22:22]),.I3(inf_abs0_2[31:31]),.I4(un32_reg0_s_19),.I5(un11_reg0_s_19),.O(reg2_16_11_a2[19:19]));
defparam desc532.INIT=64'h000000080004000C;
  LUT6 desc533(.I0(inf_abs0_2[19:19]),.I1(inf_abs0_2[20:20]),.I2(inf_abs0_2[21:21]),.I3(inf_abs0_2[31:31]),.I4(un32_reg0_s_4),.I5(un11_reg0_s_4),.O(N_1039));
defparam desc533.INIT=64'hFFFFFF3500CA0000;
  LUT6 desc534(.I0(inf_abs0_2[19:19]),.I1(inf_abs0_2[20:20]),.I2(inf_abs0_2[21:21]),.I3(inf_abs0_2[31:31]),.I4(un32_reg0_s_18),.I5(un11_reg0_s_18),.O(N_1053));
defparam desc534.INIT=64'hFFFFFF3500CA0000;
  LUT4 desc535(.I0(inf_abs0_2[20:20]),.I1(inf_abs0_2[31:31]),.I2(un32_reg0_s_6),.I3(un11_reg0_s_6),.O(N_1565));
defparam desc535.INIT=16'hFD20;
  LUT4 desc536(.I0(inf_abs0_2[19:19]),.I1(inf_abs0_2[31:31]),.I2(un32_reg0_s_7),.I3(un11_reg0_s_7),.O(N_1374));
defparam desc536.INIT=16'hFD20;
  LUT4 desc537(.I0(inf_abs0_2[20:20]),.I1(inf_abs0_2[31:31]),.I2(un32_reg0_s_8),.I3(un11_reg0_s_8),.O(N_1567));
defparam desc537.INIT=16'hFD20;
  LUT6 desc538(.I0(inf_abs0_2[19:19]),.I1(inf_abs0_2[21:21]),.I2(inf_abs0_2[22:22]),.I3(inf_abs0_2[31:31]),.I4(un32_reg0_s_23),.I5(un11_reg0_s_23),.O(reg2_16_11_a4[23:23]));
defparam desc538.INIT=64'h0000002000100030;
  LUT6 desc539(.I0(inf_abs0_2[19:19]),.I1(inf_abs0_2[20:20]),.I2(inf_abs0_2[21:21]),.I3(inf_abs0_2[31:31]),.I4(un32_reg0_s_5),.I5(un11_reg0_s_5),.O(N_1040));
defparam desc539.INIT=64'hFFFFFF3500CA0000;
  LUT6 desc540(.I0(inf_abs0_2[19:19]),.I1(inf_abs0_2[20:20]),.I2(inf_abs0_2[21:21]),.I3(inf_abs0_2[31:31]),.I4(un32_reg0_s_3),.I5(un11_reg0_s_3),.O(N_1038));
defparam desc540.INIT=64'hFFFFFF3500CA0000;
  LUT6 desc541(.I0(inf_abs0_2[19:19]),.I1(inf_abs0_2[20:20]),.I2(inf_abs0_2[21:21]),.I3(inf_abs0_2[31:31]),.I4(un32_reg0_s_12),.I5(un11_reg0_s_12),.O(N_1047));
defparam desc541.INIT=64'hFFFFFF3500CA0000;
  LUT4 desc542(.I0(inf_abs0_2[20:20]),.I1(inf_abs0_2[21:21]),.I2(inf_abs0_2[22:22]),.I3(reg3_1_1[27:27]),.O(\d_cnst_sn.reg0_28_11_2228_a6_1_1 ));
defparam desc542.INIT=16'h0100;
  LUT4 desc543(.I0(inf_abs0_2[20:20]),.I1(inf_abs0_2[31:31]),.I2(un11_reg0_s_2),.I3(un32_reg0_s_2),.O(N_1561));
defparam desc543.INIT=16'hF2D0;
  LUT4 desc544(.I0(inf_abs0_2[20:20]),.I1(inf_abs0_2[31:31]),.I2(un32_reg0_s_25),.I3(un11_reg0_s_25),.O(N_1584));
defparam desc544.INIT=16'hFD20;
  LUT4 desc545(.I0(inf_abs0_2[20:20]),.I1(inf_abs0_2[31:31]),.I2(un32_reg0_s_4),.I3(un11_reg0_s_4),.O(N_1563));
defparam desc545.INIT=16'hFD20;
  LUT4 desc546(.I0(inf_abs0_2[20:20]),.I1(inf_abs0_2[31:31]),.I2(un32_reg0_s_7),.I3(un11_reg0_s_7),.O(N_1566));
defparam desc546.INIT=16'hFD20;
  LUT4 desc547(.I0(inf_abs0_2[20:20]),.I1(inf_abs0_2[31:31]),.I2(un32_reg0_s_3),.I3(un11_reg0_s_3),.O(N_1562));
defparam desc547.INIT=16'hFD20;
  LUT6 desc548(.I0(datai[20:20]),.I1(un3_reg3_s_17),.I2(inf_abs0_2[20:20]),.I3(inf_abs0_2[31:31]),.I4(inf_abs0_2[27:27]),.I5(inf_abs0_2[28:28]),.O(reg2_16_2_d[20:20]));
defparam desc548.INIT=64'hCCACCCACCCACCC0C;
  LUT4 desc549(.I0(inf_abs0_2[20:20]),.I1(inf_abs0_2[31:31]),.I2(un11_reg0_s_1),.I3(un32_reg0_s_1),.O(N_1560));
defparam desc549.INIT=16'hF2D0;
  LUT6_L desc550(.I0(inf_abs0_2[31:31]),.I1(inf_abs0_2[28:28]),.I2(inf_abs0_2[29:29]),.I3(N_921),.I4(N_953),.I5(t_1[7:7]),.LO(t_6[7:7]));
defparam desc550.INIT=64'h44400400FFFBBFBB;
  LUT6_L desc551(.I0(inf_abs0_2[31:31]),.I1(inf_abs0_2[28:28]),.I2(inf_abs0_2[29:29]),.I3(N_920),.I4(N_952),.I5(t_1[6:6]),.LO(t_6[6:6]));
defparam desc551.INIT=64'h44400400FFFBBFBB;
  LUT6_L desc552(.I0(inf_abs0_2[31:31]),.I1(inf_abs0_2[28:28]),.I2(inf_abs0_2[29:29]),.I3(N_927),.I4(N_959),.I5(t_1[13:13]),.LO(t_6[13:13]));
defparam desc552.INIT=64'h44400400FFFBBFBB;
  LUT6_L desc553(.I0(inf_abs0_2[31:31]),.I1(inf_abs0_2[28:28]),.I2(inf_abs0_2[29:29]),.I3(N_929),.I4(N_961),.I5(t_1[15:15]),.LO(t_6[15:15]));
defparam desc553.INIT=64'h44400400FFFBBFBB;
  LUT6_L desc554(.I0(inf_abs0_2[31:31]),.I1(inf_abs0_2[28:28]),.I2(inf_abs0_2[29:29]),.I3(N_930),.I4(N_962),.I5(t_1[16:16]),.LO(t_6[16:16]));
defparam desc554.INIT=64'h44400400FFFBBFBB;
  LUT6_L desc555(.I0(inf_abs0_2[31:31]),.I1(inf_abs0_2[28:28]),.I2(inf_abs0_2[29:29]),.I3(N_928),.I4(N_960),.I5(t_1[14:14]),.LO(t_6[14:14]));
defparam desc555.INIT=64'h44400400FFFBBFBB;
  LUT5 desc556(.I0(inf_abs0_2[31:31]),.I1(inf_abs0_2[28:28]),.I2(inf_abs0_2[29:29]),.I3(N_934),.I4(N_2722),.O(\d_cnst_sn.reg3_17_4_a2_0 [20:20]));
defparam desc556.INIT=32'h44400400;
  LUT6_L desc557(.I0(N_513_i),.I1(N_514_i),.I2(N_527_i),.I3(N_1335),.I4(N_1035),.I5(t_1[0:0]),.LO(reg2_16[0:0]));
defparam desc557.INIT=64'h1100776619087F6E;
  LUT6_L desc558(.I0(inf_abs0_2[31:31]),.I1(inf_abs0_2[28:28]),.I2(inf_abs0_2[29:29]),.I3(N_923),.I4(N_955),.I5(t_1[9:9]),.LO(r_4_1_RNIIQ731[8:8]));
defparam desc558.INIT=64'hBBBFFBFF00044044;
  LUT6_L desc559(.I0(inf_abs0_2[31:31]),.I1(inf_abs0_2[28:28]),.I2(inf_abs0_2[29:29]),.I3(N_925),.I4(N_957),.I5(t_1[11:11]),.LO(t_6[11:11]));
defparam desc559.INIT=64'h44400400FFFBBFBB;
  LUT6_L desc560(.I0(inf_abs0_2[31:31]),.I1(inf_abs0_2[28:28]),.I2(inf_abs0_2[29:29]),.I3(N_926),.I4(N_958),.I5(t_1[12:12]),.LO(t_6[12:12]));
defparam desc560.INIT=64'h44400400FFFBBFBB;
  LUT6_L desc561(.I0(inf_abs0_2[31:31]),.I1(inf_abs0_2[28:28]),.I2(inf_abs0_2[29:29]),.I3(N_920),.I4(N_952),.I5(t_1[6:6]),.LO(r_4_1_RNI9K731[5:5]));
defparam desc561.INIT=64'hBBBFFBFF00044044;
  LUT6_L desc562(.I0(inf_abs0_2[31:31]),.I1(inf_abs0_2[28:28]),.I2(inf_abs0_2[29:29]),.I3(N_921),.I4(N_953),.I5(t_1[7:7]),.LO(r_4_1_RNICM731[6:6]));
defparam desc562.INIT=64'hBBBFFBFF00044044;
  LUT6_L desc563(.I0(inf_abs0_2[31:31]),.I1(inf_abs0_2[28:28]),.I2(inf_abs0_2[29:29]),.I3(N_925),.I4(N_957),.I5(t_1[11:11]),.LO(r_4_1_RNIDBOH1[10:10]));
defparam desc563.INIT=64'hBBBFFBFF00044044;
  LUT6_L desc564(.I0(inf_abs0_2[31:31]),.I1(inf_abs0_2[28:28]),.I2(inf_abs0_2[29:29]),.I3(N_924),.I4(N_956),.I5(t_1[10:10]),.LO(r_4_1_RNIS3K91[9:9]));
defparam desc564.INIT=64'hBBBFFBFF00044044;
  LUT6_L desc565(.I0(inf_abs0_2[31:31]),.I1(inf_abs0_2[28:28]),.I2(inf_abs0_2[29:29]),.I3(N_922),.I4(N_954),.I5(t_1[8:8]),.LO(r_4_1_RNIFO731[7:7]));
defparam desc565.INIT=64'hBBBFFBFF00044044;
  LUT6 desc566(.I0(inf_abs0_2[21:21]),.I1(inf_abs0_2[31:31]),.I2(inf_abs0_2[28:28]),.I3(inf_abs0_2[29:29]),.I4(N_931),.I5(N_963),.O(reg0_28_7_a1[17:17]));
defparam desc566.INIT=64'h0000002020002020;
  LUT6_L desc567(.I0(inf_abs0_2[31:31]),.I1(inf_abs0_2[28:28]),.I2(inf_abs0_2[29:29]),.I3(N_922),.I4(N_954),.I5(t_1[8:8]),.LO(t_6[8:8]));
defparam desc567.INIT=64'h44400400FFFBBFBB;
  LUT6_L desc568(.I0(inf_abs0_2[31:31]),.I1(inf_abs0_2[28:28]),.I2(inf_abs0_2[29:29]),.I3(N_923),.I4(N_955),.I5(t_1[9:9]),.LO(t_6[9:9]));
defparam desc568.INIT=64'h44400400FFFBBFBB;
  LUT6 desc569(.I0(inf_abs0_2[21:21]),.I1(inf_abs0_2[31:31]),.I2(inf_abs0_2[28:28]),.I3(inf_abs0_2[29:29]),.I4(N_932),.I5(N_964),.O(reg0_28_7_a1[18:18]));
defparam desc569.INIT=64'h0000002020002020;
  LUT6_L desc570(.I0(inf_abs0_2[31:31]),.I1(inf_abs0_2[28:28]),.I2(inf_abs0_2[29:29]),.I3(N_924),.I4(N_956),.I5(t_1[10:10]),.LO(t_6[10:10]));
defparam desc570.INIT=64'h44400400FFFBBFBB;
  LUT6_L desc571(.I0(N_7_i),.I1(un36_df),.I2(un1_b59),.I3(un87_df),.I4(un32_reg0_s_23),.I5(un11_reg0_s_23),.LO(N_1742));
defparam desc571.INIT=64'hFFFFEFFF10000000;
  LUT6_L desc572(.I0(N_7_i),.I1(un36_df),.I2(un1_b59),.I3(un87_df),.I4(un32_reg0_s_24),.I5(un11_reg0_s_24),.LO(N_1743));
defparam desc572.INIT=64'hFFFFEFFF10000000;
  LUT6_L desc573(.I0(inf_abs0_2[21:21]),.I1(inf_abs0_2[31:31]),.I2(inf_abs0_2[28:28]),.I3(r_4[17:17]),.I4(reg3_1_1[18:18]),.I5(t_1[18:18]),.LO(N_1085));
defparam desc573.INIT=64'hFDDD2000FFDF2202;
  LUT6 desc574(.I0(N_7_i),.I1(un36_df),.I2(un1_b59),.I3(un87_df),.I4(un32_reg0_s_13),.I5(un11_reg0_s_13),.O(N_1732));
defparam desc574.INIT=64'hFFFFEFFF10000000;
  LUT6_L desc575(.I0(inf_abs0_2[21:21]),.I1(inf_abs0_2[31:31]),.I2(inf_abs0_2[28:28]),.I3(r_4[16:16]),.I4(reg3_1_1[17:17]),.I5(t_1[17:17]),.LO(N_1084));
defparam desc575.INIT=64'hFDDD2000FFDF2202;
  LUT5 desc576(.I0(datai[0:0]),.I1(m_2[0:0]),.I2(N_1035),.I3(un1_cf),.I4(N_1810),.O(N_1812));
defparam desc576.INIT=32'hCCAA0F0F;
  LUT6_L desc577(.I0(N_7_i),.I1(un36_df),.I2(un1_b59),.I3(un87_df),.I4(un32_reg0_s_22),.I5(un11_reg0_s_22),.LO(N_1741));
defparam desc577.INIT=64'hFFFFEFFF10000000;
  LUT6_L desc578(.I0(N_7_i),.I1(un36_df),.I2(un1_b59),.I3(un87_df),.I4(un32_reg0_s_21),.I5(un11_reg0_s_21),.LO(N_1740));
defparam desc578.INIT=64'hFFFFEFFF10000000;
  MUXCY_L un3_t_cry_0_cy_cZ(.DI(GND),.CI(VCC),.S(r_4_3_ci[31:31]),.LO(un3_t_cry_0_cy));
  LUT6 desc579(.I0(reg0[31:31]),.I1(reg1[31:31]),.I2(reg2[31:31]),.I3(inf_abs0_2[31:31]),.I4(inf_abs0_2[29:29]),.I5(inf_abs0_2[30:30]),.O(r_4_3_ci[31:31]));
defparam desc579.INIT=64'hAA00AAF0AACCAAAA;
  MUXCY_L t_1_cry_0_cy_cZ(.DI(GND),.CI(VCC),.S(r_4_i[31:31]),.LO(t_1_cry_0_cy));
  LUT5 desc580(.I0(reg0[2:2]),.I1(reg2[2:2]),.I2(inf_abs0_2[31:31]),.I3(\d_cnst_sn.m19_0_1 ),.I4(\d_cnst_sn.m26_0_1 ),.O(N_28));
defparam desc580.INIT=32'hACA0AFAA;
  LUT5 un3_t_axb_2_cZ(.I0(reg0[2:2]),.I1(reg2[2:2]),.I2(inf_abs0_2[31:31]),.I3(\d_cnst_sn.m19_0_1 ),.I4(\d_cnst_sn.m26_0_1 ),.O(un3_t_axb_2));
defparam un3_t_axb_2_cZ.INIT=32'h535F5055;
  LUT5_L desc581(.I0(inf_abs0_2[31:31]),.I1(\d_cnst_sn.reg0_28_14_2135_1_a0_2 ),.I2(reg3_1_1[30:30]),.I3(\d_cnst_sn.reg0_28_14_0 ),.I4(t_1[30:30]),.LO(N_3550));
defparam desc581.INIT=32'hFFA0FFEC;
  LUT4 desc582(.I0(m_2[21:21]),.I1(\d_cnst_sn.reg3_17_a2_2_0 [21:21]),.I2(\d_cnst_sn.reg3_17_sn_m7_0 ),.I3(reg3_14_sqmuxa),.O(\d_cnst_sn.reg3_17_0_tz [21:21]));
defparam desc582.INIT=16'hC00A;
  LUT5_L desc583(.I0(N_3916),.I1(\d_cnst_sn.reg0_28_7_a0_0 [9:9]),.I2(\d_cnst_sn.reg0_0 [17:17]),.I3(t_1[17:17]),.I4(N_1052),.LO(reg0_28[17:17]));
defparam desc583.INIT=32'hB0F01050;
  LUT5_L desc584(.I0(N_3916),.I1(\d_cnst_sn.reg0_28_7_a0_0 [9:9]),.I2(\d_cnst_sn.reg1_0 [18:18]),.I3(t_1[18:18]),.I4(N_1053),.LO(reg1_16[18:18]));
defparam desc584.INIT=32'hB0F01050;
  LUT1_L desc585(.I0(state),.LO(state_i));
defparam desc585.INIT=2'h1;
  LUT2 un1_inf_abs0_0_s_19_RNO(.I0(reg1[19:19]),.I1(inf_abs0_2[19:19]),.O(un1_inf_abs0_0_axb_19));
defparam un1_inf_abs0_0_s_19_RNO.INIT=4'h6;
  LUT2 un1_inf_abs0_s_19_RNO(.I0(reg2[19:19]),.I1(inf_abs0_2[19:19]),.O(un1_inf_abs0_axb_19));
defparam un1_inf_abs0_s_19_RNO.INIT=4'h6;
  LUT2 desc586(.I0(inf_abs0_2[31:31]),.I1(inf_abs0_2[30:30]),.O(N_3_0));
defparam desc586.INIT=4'h4;
  LUT3_L desc587(.I0(datai[8:8]),.I1(state),.I2(inf_abs0_2[8:8]),.LO(ir_3[8:8]));
defparam desc587.INIT=8'hE2;
  LUT3_L desc588(.I0(datai[16:16]),.I1(state),.I2(inf_abs0_2[16:16]),.LO(ir_3[16:16]));
defparam desc588.INIT=8'hE2;
  LUT3_L desc589(.I0(datai[3:3]),.I1(state),.I2(inf_abs0_2[3:3]),.LO(ir_3[3:3]));
defparam desc589.INIT=8'hE2;
  LUT3_L desc590(.I0(datai[0:0]),.I1(state),.I2(inf_abs0_2[0:0]),.LO(ir_3[0:0]));
defparam desc590.INIT=8'hE2;
  LUT3_L desc591(.I0(datai[27:27]),.I1(state),.I2(inf_abs0_2[27:27]),.LO(ir_3[27:27]));
defparam desc591.INIT=8'hE2;
  LUT3_L desc592(.I0(datai[23:23]),.I1(state),.I2(inf_abs0_2[23:23]),.LO(ir_3[23:23]));
defparam desc592.INIT=8'hE2;
  LUT3_L desc593(.I0(datai[26:26]),.I1(state),.I2(inf_abs0_2[26:26]),.LO(ir_3[26:26]));
defparam desc593.INIT=8'hE2;
  LUT3_L desc594(.I0(datai[5:5]),.I1(state),.I2(inf_abs0_2[5:5]),.LO(ir_3[5:5]));
defparam desc594.INIT=8'hE2;
  LUT3_L desc595(.I0(datai[2:2]),.I1(state),.I2(inf_abs0_2[2:2]),.LO(ir_3[2:2]));
defparam desc595.INIT=8'hE2;
  LUT3_L desc596(.I0(datai[18:18]),.I1(state),.I2(inf_abs0_2[18:18]),.LO(ir_3[18:18]));
defparam desc596.INIT=8'hE2;
  LUT3_L desc597(.I0(datai[19:19]),.I1(state),.I2(inf_abs0_2[19:19]),.LO(ir_3[19:19]));
defparam desc597.INIT=8'hE2;
  LUT3_L desc598(.I0(datai[10:10]),.I1(state),.I2(inf_abs0_2[10:10]),.LO(ir_3[10:10]));
defparam desc598.INIT=8'hE2;
  LUT3_L desc599(.I0(datai[9:9]),.I1(state),.I2(inf_abs0_2[9:9]),.LO(ir_3[9:9]));
defparam desc599.INIT=8'hE2;
  LUT3_L desc600(.I0(datai[6:6]),.I1(state),.I2(inf_abs0_2[6:6]),.LO(ir_3[6:6]));
defparam desc600.INIT=8'hE2;
  LUT3_L desc601(.I0(datai[4:4]),.I1(state),.I2(inf_abs0_2[4:4]),.LO(ir_3[4:4]));
defparam desc601.INIT=8'hE2;
  LUT3_L desc602(.I0(datai[22:22]),.I1(state),.I2(inf_abs0_2[22:22]),.LO(ir_3[22:22]));
defparam desc602.INIT=8'hE2;
  LUT3 desc603(.I0(reg1[19:19]),.I1(un3_reg3_s_16),.I2(inf_abs0_2[30:30]),.O(N_2722));
defparam desc603.INIT=8'hCA;
  LUT3_L desc604(.I0(datai[21:21]),.I1(state),.I2(inf_abs0_2[21:21]),.LO(ir_3[21:21]));
defparam desc604.INIT=8'hE2;
  LUT3_L desc605(.I0(datai[1:1]),.I1(state),.I2(inf_abs0_2[1:1]),.LO(ir_3[1:1]));
defparam desc605.INIT=8'hE2;
  LUT3_L desc606(.I0(datai[7:7]),.I1(state),.I2(inf_abs0_2[7:7]),.LO(ir_3[7:7]));
defparam desc606.INIT=8'hE2;
  LUT3_L desc607(.I0(datai[25:25]),.I1(state),.I2(inf_abs0_2[25:25]),.LO(ir_3[25:25]));
defparam desc607.INIT=8'hE2;
  LUT3_L desc608(.I0(datai[24:24]),.I1(state),.I2(inf_abs0_2[24:24]),.LO(ir_3[24:24]));
defparam desc608.INIT=8'hE2;
  LUT3_L desc609(.I0(datai[29:29]),.I1(state),.I2(inf_abs0_2[29:29]),.LO(ir_3[29:29]));
defparam desc609.INIT=8'hE2;
  LUT3_L desc610(.I0(datai[11:11]),.I1(state),.I2(inf_abs0_2[11:11]),.LO(ir_3[11:11]));
defparam desc610.INIT=8'hE2;
  LUT3 desc611(.I0(reg3[0:0]),.I1(inf_abs0_2[31:31]),.I2(inf_abs0_2[30:30]),.O(r_4_2_a0[0:0]));
defparam desc611.INIT=8'h10;
  LUT3 desc612(.I0(reg3[1:1]),.I1(inf_abs0_2[31:31]),.I2(inf_abs0_2[30:30]),.O(r_4_2_a0[1:1]));
defparam desc612.INIT=8'h10;
  LUT3 desc613(.I0(reg1[0:0]),.I1(inf_abs0_2[31:31]),.I2(inf_abs0_2[30:30]),.O(\d_cnst_sn.r_4_0_0 [0:0]));
defparam desc613.INIT=8'hBA;
  LUT3 desc614(.I0(reg1[1:1]),.I1(inf_abs0_2[31:31]),.I2(inf_abs0_2[30:30]),.O(\d_cnst_sn.r_4_0_0 [1:1]));
defparam desc614.INIT=8'hBA;
  LUT3 desc615(.I0(inf_abs0_2[31:31]),.I1(inf_abs0_2[27:27]),.I2(inf_abs0_2[28:28]),.O(m7));
defparam desc615.INIT=8'hAB;
  LUT2 inf_abs0_2_axb_30_cZ(.I0(ir[30:30]),.I1(ir[31:31]),.O(inf_abs0_2_axb_30));
defparam inf_abs0_2_axb_30_cZ.INIT=4'h6;
  LUT2 desc616(.I0(inf_abs0_2[23:23]),.I1(inf_abs0_2[31:31]),.O(N_7_i));
defparam desc616.INIT=4'h2;
  LUT2 desc617(.I0(inf_abs0_2[31:31]),.I1(inf_abs0_2[29:29]),.O(N_13));
defparam desc617.INIT=4'hB;
  LUT2 desc618(.I0(inf_abs0_2[22:22]),.I1(inf_abs0_2[31:31]),.O(N_514_i));
defparam desc618.INIT=4'h2;
  LUT2 desc619(.I0(inf_abs0_2[21:21]),.I1(inf_abs0_2[31:31]),.O(N_513_i));
defparam desc619.INIT=4'h2;
  LUT4 desc620(.I0(reg0[11:11]),.I1(reg2[11:11]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[30:30]),.O(N_926));
defparam desc620.INIT=16'hACAA;
  LUT4 desc621(.I0(reg0[26:26]),.I1(reg2[26:26]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[30:30]),.O(N_941));
defparam desc621.INIT=16'hACAA;
  LUT4 desc622(.I0(reg1[11:11]),.I1(un3_reg3_s_8),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[30:30]),.O(N_958));
defparam desc622.INIT=16'hACAA;
  LUT4 desc623(.I0(reg1[26:26]),.I1(un3_reg3_s_23),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[30:30]),.O(N_973));
defparam desc623.INIT=16'hACAA;
  LUT4 desc624(.I0(reg0[28:28]),.I1(reg2[28:28]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[30:30]),.O(N_943));
defparam desc624.INIT=16'hACAA;
  LUT4 desc625(.I0(reg1[28:28]),.I1(un3_reg3_s_25),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[30:30]),.O(N_975));
defparam desc625.INIT=16'hACAA;
  LUT4 desc626(.I0(reg0[25:25]),.I1(reg2[25:25]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[30:30]),.O(N_940));
defparam desc626.INIT=16'hACAA;
  LUT4 desc627(.I0(reg1[25:25]),.I1(un3_reg3_s_22),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[30:30]),.O(N_972));
defparam desc627.INIT=16'hACAA;
  LUT4 desc628(.I0(reg0[13:13]),.I1(reg2[13:13]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[30:30]),.O(N_928));
defparam desc628.INIT=16'hACAA;
  LUT4 desc629(.I0(reg1[13:13]),.I1(un3_reg3_s_10),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[30:30]),.O(N_960));
defparam desc629.INIT=16'hACAA;
  LUT4 desc630(.I0(reg0[16:16]),.I1(reg2[16:16]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[30:30]),.O(N_931));
defparam desc630.INIT=16'hACAA;
  LUT4 desc631(.I0(reg1[16:16]),.I1(un3_reg3_s_13),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[30:30]),.O(N_963));
defparam desc631.INIT=16'hACAA;
  LUT4 desc632(.I0(reg0[14:14]),.I1(reg2[14:14]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[30:30]),.O(N_929));
defparam desc632.INIT=16'hACAA;
  LUT4 desc633(.I0(reg1[14:14]),.I1(un3_reg3_s_11),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[30:30]),.O(N_961));
defparam desc633.INIT=16'hACAA;
  LUT4 desc634(.I0(reg0[10:10]),.I1(reg2[10:10]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[30:30]),.O(N_925));
defparam desc634.INIT=16'hACAA;
  LUT4 desc635(.I0(reg1[10:10]),.I1(un3_reg3_s_7),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[30:30]),.O(N_957));
defparam desc635.INIT=16'hACAA;
  LUT4 desc636(.I0(reg0[9:9]),.I1(reg2[9:9]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[30:30]),.O(N_924));
defparam desc636.INIT=16'hACAA;
  LUT4 desc637(.I0(reg1[9:9]),.I1(un3_reg3_s_6),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[30:30]),.O(N_956));
defparam desc637.INIT=16'hACAA;
  LUT4 desc638(.I0(reg0[7:7]),.I1(reg2[7:7]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[30:30]),.O(N_922));
defparam desc638.INIT=16'hACAA;
  LUT4 desc639(.I0(reg0[8:8]),.I1(reg2[8:8]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[30:30]),.O(N_923));
defparam desc639.INIT=16'hACAA;
  LUT4 desc640(.I0(reg1[7:7]),.I1(un3_reg3_s_4),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[30:30]),.O(N_954));
defparam desc640.INIT=16'hACAA;
  LUT4 desc641(.I0(reg1[8:8]),.I1(un3_reg3_s_5),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[30:30]),.O(N_955));
defparam desc641.INIT=16'hACAA;
  LUT4 desc642(.I0(reg0[21:21]),.I1(reg2[21:21]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[30:30]),.O(N_936));
defparam desc642.INIT=16'hACAA;
  LUT4 desc643(.I0(reg1[21:21]),.I1(un3_reg3_s_18),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[30:30]),.O(N_968));
defparam desc643.INIT=16'hACAA;
  LUT4 desc644(.I0(reg0[20:20]),.I1(reg2[20:20]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[30:30]),.O(N_935));
defparam desc644.INIT=16'hACAA;
  LUT4 desc645(.I0(reg1[20:20]),.I1(un3_reg3_s_17),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[30:30]),.O(N_967));
defparam desc645.INIT=16'hACAA;
  LUT4 desc646(.I0(reg0[15:15]),.I1(reg2[15:15]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[30:30]),.O(N_930));
defparam desc646.INIT=16'hACAA;
  LUT4 desc647(.I0(reg0[17:17]),.I1(reg2[17:17]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[30:30]),.O(N_932));
defparam desc647.INIT=16'hACAA;
  LUT4 desc648(.I0(reg1[15:15]),.I1(un3_reg3_s_12),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[30:30]),.O(N_962));
defparam desc648.INIT=16'hACAA;
  LUT4 desc649(.I0(reg1[17:17]),.I1(un3_reg3_s_14),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[30:30]),.O(N_964));
defparam desc649.INIT=16'hACAA;
  LUT4 desc650(.I0(reg0[5:5]),.I1(reg2[5:5]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[30:30]),.O(N_920));
defparam desc650.INIT=16'hACAA;
  LUT4 desc651(.I0(reg1[5:5]),.I1(un3_reg3_s_2),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[30:30]),.O(N_952));
defparam desc651.INIT=16'hACAA;
  LUT4 desc652(.I0(reg0[27:27]),.I1(reg2[27:27]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[30:30]),.O(N_942));
defparam desc652.INIT=16'hACAA;
  LUT4 desc653(.I0(reg1[27:27]),.I1(un3_reg3_s_24),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[30:30]),.O(N_974));
defparam desc653.INIT=16'hACAA;
  LUT4 desc654(.I0(reg0[18:18]),.I1(reg2[18:18]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[30:30]),.O(N_933));
defparam desc654.INIT=16'hACAA;
  LUT4 desc655(.I0(reg1[18:18]),.I1(un3_reg3_s_15),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[30:30]),.O(N_965));
defparam desc655.INIT=16'hACAA;
  LUT4 desc656(.I0(reg0[22:22]),.I1(reg2[22:22]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[30:30]),.O(N_937));
defparam desc656.INIT=16'hACAA;
  LUT4 desc657(.I0(reg1[22:22]),.I1(un3_reg3_s_19),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[30:30]),.O(N_969));
defparam desc657.INIT=16'hACAA;
  LUT4 desc658(.I0(reg0[12:12]),.I1(reg2[12:12]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[30:30]),.O(N_927));
defparam desc658.INIT=16'hACAA;
  LUT4 desc659(.I0(reg1[12:12]),.I1(un3_reg3_s_9),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[30:30]),.O(N_959));
defparam desc659.INIT=16'hACAA;
  LUT4 desc660(.I0(reg0[6:6]),.I1(reg2[6:6]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[30:30]),.O(N_921));
defparam desc660.INIT=16'hACAA;
  LUT4 desc661(.I0(reg1[6:6]),.I1(un3_reg3_s_3),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[30:30]),.O(N_953));
defparam desc661.INIT=16'hACAA;
  LUT4 desc662(.I0(reg0[19:19]),.I1(reg2[19:19]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[30:30]),.O(N_934));
defparam desc662.INIT=16'hACAA;
  LUT4 desc663(.I0(reg1[23:23]),.I1(un3_reg3_s_20),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[30:30]),.O(N_970));
defparam desc663.INIT=16'hACAA;
  LUT4 desc664(.I0(reg0[23:23]),.I1(reg2[23:23]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[30:30]),.O(N_938));
defparam desc664.INIT=16'hACAA;
  LUT4 desc665(.I0(reg1[24:24]),.I1(un3_reg3_s_21),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[30:30]),.O(N_971));
defparam desc665.INIT=16'hACAA;
  LUT4 desc666(.I0(reg0[24:24]),.I1(reg2[24:24]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[30:30]),.O(N_939));
defparam desc666.INIT=16'hACAA;
  LUT4 desc667(.I0(reg1[2:2]),.I1(reg3[2:2]),.I2(inf_abs0_2[29:29]),.I3(inf_abs0_2[30:30]),.O(\d_cnst_sn.m19_0_1 ));
defparam desc667.INIT=16'hCFA0;
  LUT4 desc668(.I0(reg1[2:2]),.I1(reg3[2:2]),.I2(inf_abs0_2[29:29]),.I3(inf_abs0_2[30:30]),.O(\d_cnst_sn.m26_0_1 ));
defparam desc668.INIT=16'h3F50;
  LUT4 desc669(.I0(reg1[3:3]),.I1(reg3[3:3]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[30:30]),.O(\d_cnst_sn.r_4_0_0 [3:3]));
defparam desc669.INIT=16'hA3AF;
  LUT4 desc670(.I0(reg1[4:4]),.I1(un3_reg3_s_1),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[30:30]),.O(\d_cnst_sn.r_4_0_0 [4:4]));
defparam desc670.INIT=16'hACAF;
  LUT6 desc671(.I0(m_2[22:22]),.I1(m_2[23:23]),.I2(m_2[21:21]),.I3(r_4[21:21]),.I4(r_4[23:23]),.I5(r_4[22:22]),.O(un14_r_0_N_56));
defparam desc671.INIT=64'h8008200240041001;
  LUT5 desc672(.I0(state),.I1(inf_abs0_2[24:24]),.I2(inf_abs0_2[23:23]),.I3(inf_abs0_2[25:25]),.I4(inf_abs0_2[26:26]),.O(N_2641));
defparam desc672.INIT=32'h08000000;
  LUT6 desc673(.I0(m_2[24:24]),.I1(m_2[25:25]),.I2(m_2[26:26]),.I3(r_4[24:24]),.I4(r_4[25:25]),.I5(r_4[26:26]),.O(un14_r_0_N_35));
defparam desc673.INIT=64'h8040201008040201;
  LUT4 desc674(.I0(reg0[0:0]),.I1(reg2[0:0]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[30:30]),.O(N_915));
defparam desc674.INIT=16'hACAA;
  LUT4 desc675(.I0(reg0[1:1]),.I1(reg2[1:1]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[30:30]),.O(N_916));
defparam desc675.INIT=16'hACAA;
  LUT6_L desc676(.I0(reg0[29:29]),.I1(reg1[29:29]),.I2(reg2[29:29]),.I3(un3_reg3_cry_25),.I4(inf_abs0_2[29:29]),.I5(inf_abs0_2[30:30]),.LO(r_4_3_6_1508_i_m2));
defparam desc676.INIT=64'hFF00F0F0CCCCAAAA;
  LUT6_L desc677(.I0(reg1[28:28]),.I1(reg0[28:28]),.I2(reg2[28:28]),.I3(un3_reg3_s_25),.I4(inf_abs0_2[29:29]),.I5(inf_abs0_2[30:30]),.LO(r_4_3_5_1534_i_m2));
defparam desc677.INIT=64'hFF00F0F0AAAACCCC;
  LUT6_L desc678(.I0(reg0[24:24]),.I1(reg2[24:24]),.I2(reg1[24:24]),.I3(un3_reg3_s_21),.I4(inf_abs0_2[29:29]),.I5(inf_abs0_2[30:30]),.LO(r_4_3_1_1638_i_m2));
defparam desc678.INIT=64'hFF00CCCCF0F0AAAA;
  LUT6_L desc679(.I0(reg1[16:16]),.I1(reg0[16:16]),.I2(reg2[16:16]),.I3(un3_reg3_s_13),.I4(inf_abs0_2[29:29]),.I5(inf_abs0_2[30:30]),.LO(r_4_3_18_1208_i_m2));
defparam desc679.INIT=64'hFF00F0F0AAAACCCC;
  LUT6_L desc680(.I0(reg1[13:13]),.I1(reg0[13:13]),.I2(reg2[13:13]),.I3(un3_reg3_s_10),.I4(inf_abs0_2[29:29]),.I5(inf_abs0_2[30:30]),.LO(r_4_3_15_1286_i_m2));
defparam desc680.INIT=64'hFF00F0F0AAAACCCC;
  LUT6_L desc681(.I0(reg1[11:11]),.I1(reg0[11:11]),.I2(reg2[11:11]),.I3(un3_reg3_s_8),.I4(inf_abs0_2[29:29]),.I5(inf_abs0_2[30:30]),.LO(r_4_3_13_1338_i_m2));
defparam desc681.INIT=64'hFF00F0F0AAAACCCC;
  LUT6_L desc682(.I0(reg1[17:17]),.I1(reg0[17:17]),.I2(reg2[17:17]),.I3(un3_reg3_s_14),.I4(inf_abs0_2[29:29]),.I5(inf_abs0_2[30:30]),.LO(r_4_3_19_1182_i_m2));
defparam desc682.INIT=64'hFF00F0F0AAAACCCC;
  LUT6_L desc683(.I0(reg1[12:12]),.I1(reg0[12:12]),.I2(reg2[12:12]),.I3(un3_reg3_s_9),.I4(inf_abs0_2[29:29]),.I5(inf_abs0_2[30:30]),.LO(r_4_3_14_1312_i_m2));
defparam desc683.INIT=64'hFF00F0F0AAAACCCC;
  LUT6_L desc684(.I0(reg1[10:10]),.I1(reg0[10:10]),.I2(reg2[10:10]),.I3(un3_reg3_s_7),.I4(inf_abs0_2[29:29]),.I5(inf_abs0_2[30:30]),.LO(r_4_3_12_1364_i_m2));
defparam desc684.INIT=64'hFF00F0F0AAAACCCC;
  LUT6_L desc685(.I0(reg1[26:26]),.I1(reg0[26:26]),.I2(reg2[26:26]),.I3(un3_reg3_s_23),.I4(inf_abs0_2[29:29]),.I5(inf_abs0_2[30:30]),.LO(r_4_3_3_1586_i_m2));
defparam desc685.INIT=64'hFF00F0F0AAAACCCC;
  LUT6_L desc686(.I0(reg1[14:14]),.I1(reg0[14:14]),.I2(reg2[14:14]),.I3(un3_reg3_s_11),.I4(inf_abs0_2[29:29]),.I5(inf_abs0_2[30:30]),.LO(r_4_3_16_1260_i_m2));
defparam desc686.INIT=64'hFF00F0F0AAAACCCC;
  LUT6_L desc687(.I0(reg1[9:9]),.I1(reg0[9:9]),.I2(reg2[9:9]),.I3(un3_reg3_s_6),.I4(inf_abs0_2[29:29]),.I5(inf_abs0_2[30:30]),.LO(r_4_3_11_1390_i_m2));
defparam desc687.INIT=64'hFF00F0F0AAAACCCC;
  LUT6_L desc688(.I0(reg1[6:6]),.I1(reg0[6:6]),.I2(reg2[6:6]),.I3(un3_reg3_s_3),.I4(inf_abs0_2[29:29]),.I5(inf_abs0_2[30:30]),.LO(r_4_3_30_680_i_m2));
defparam desc688.INIT=64'hFF00F0F0AAAACCCC;
  LUT6_L desc689(.I0(reg1[8:8]),.I1(reg0[8:8]),.I2(reg2[8:8]),.I3(un3_reg3_s_5),.I4(inf_abs0_2[29:29]),.I5(inf_abs0_2[30:30]),.LO(r_4_3_10_1416_i_m2));
defparam desc689.INIT=64'hFF00F0F0AAAACCCC;
  LUT6_L desc690(.I0(reg1[7:7]),.I1(reg0[7:7]),.I2(reg2[7:7]),.I3(un3_reg3_s_4),.I4(inf_abs0_2[29:29]),.I5(inf_abs0_2[30:30]),.LO(r_4_3_9_1442_i_m2));
defparam desc690.INIT=64'hFF00F0F0AAAACCCC;
  LUT6_L desc691(.I0(reg0[23:23]),.I1(reg2[23:23]),.I2(reg1[23:23]),.I3(un3_reg3_s_20),.I4(inf_abs0_2[29:29]),.I5(inf_abs0_2[30:30]),.LO(r_4_3_0_1664_i_m2));
defparam desc691.INIT=64'hFF00CCCCF0F0AAAA;
  LUT6_L desc692(.I0(reg0[20:20]),.I1(reg2[20:20]),.I2(reg1[20:20]),.I3(un3_reg3_s_17),.I4(inf_abs0_2[29:29]),.I5(inf_abs0_2[30:30]),.LO(r_4_3_22_1104_i_m2));
defparam desc692.INIT=64'hFF00CCCCF0F0AAAA;
  LUT6_L desc693(.I0(reg0[1:1]),.I1(reg2[1:1]),.I2(reg1[1:1]),.I3(reg3[1:1]),.I4(inf_abs0_2[29:29]),.I5(inf_abs0_2[30:30]),.LO(r_4_3_25_810_i_m2));
defparam desc693.INIT=64'hFF00CCCCF0F0AAAA;
  LUT6_L desc694(.I0(reg1[15:15]),.I1(reg0[15:15]),.I2(reg2[15:15]),.I3(un3_reg3_s_12),.I4(inf_abs0_2[29:29]),.I5(inf_abs0_2[30:30]),.LO(r_4_3_17_1234_i_m2));
defparam desc694.INIT=64'hFF00F0F0AAAACCCC;
  LUT6_L desc695(.I0(reg1[5:5]),.I1(reg0[5:5]),.I2(reg2[5:5]),.I3(un3_reg3_s_2),.I4(inf_abs0_2[29:29]),.I5(inf_abs0_2[30:30]),.LO(r_4_3_29_706_i_m2));
defparam desc695.INIT=64'hFF00F0F0AAAACCCC;
  LUT6_L desc696(.I0(reg0[0:0]),.I1(reg2[0:0]),.I2(reg1[0:0]),.I3(reg3[0:0]),.I4(inf_abs0_2[29:29]),.I5(inf_abs0_2[30:30]),.LO(r_4_3_24_836_i_m2));
defparam desc696.INIT=64'hFF00CCCCF0F0AAAA;
  LUT6_L desc697(.I0(reg0[27:27]),.I1(reg2[27:27]),.I2(reg1[27:27]),.I3(un3_reg3_s_24),.I4(inf_abs0_2[29:29]),.I5(inf_abs0_2[30:30]),.LO(r_4_3_4_1560_i_m2));
defparam desc697.INIT=64'hFF00CCCCF0F0AAAA;
  LUT4 desc698(.I0(datai[29:29]),.I1(inf_abs0_2[31:31]),.I2(inf_abs0_2[27:27]),.I3(inf_abs0_2[28:28]),.O(m_2[29:29]));
defparam desc698.INIT=16'h2220;
  LUT6_L desc699(.I0(reg1[18:18]),.I1(reg0[18:18]),.I2(reg2[18:18]),.I3(un3_reg3_s_15),.I4(inf_abs0_2[29:29]),.I5(inf_abs0_2[30:30]),.LO(r_4_3_20_1156_i_m2));
defparam desc699.INIT=64'hFF00F0F0AAAACCCC;
  LUT6_L desc700(.I0(reg0[22:22]),.I1(reg2[22:22]),.I2(reg1[22:22]),.I3(un3_reg3_s_19),.I4(inf_abs0_2[29:29]),.I5(inf_abs0_2[30:30]),.LO(r_4_3_1690_i_m2));
defparam desc700.INIT=64'hFF00CCCCF0F0AAAA;
  LUT6_L desc701(.I0(reg0[4:4]),.I1(reg2[4:4]),.I2(reg1[4:4]),.I3(un3_reg3_s_1),.I4(inf_abs0_2[29:29]),.I5(inf_abs0_2[30:30]),.LO(r_4_3_28_732_i_m2));
defparam desc701.INIT=64'hFF00CCCCF0F0AAAA;
  LUT6_L desc702(.I0(reg1[25:25]),.I1(reg0[25:25]),.I2(reg2[25:25]),.I3(un3_reg3_s_22),.I4(inf_abs0_2[29:29]),.I5(inf_abs0_2[30:30]),.LO(r_4_3_2_1612_i_m2));
defparam desc702.INIT=64'hFF00F0F0AAAACCCC;
  LUT6_L desc703(.I0(reg1[21:21]),.I1(reg0[21:21]),.I2(reg2[21:21]),.I3(un3_reg3_s_18),.I4(inf_abs0_2[29:29]),.I5(inf_abs0_2[30:30]),.LO(r_4_3_23_1078_i_m2));
defparam desc703.INIT=64'hFF00F0F0AAAACCCC;
  LUT6_L desc704(.I0(reg0[3:3]),.I1(reg2[3:3]),.I2(reg1[3:3]),.I3(reg3[3:3]),.I4(inf_abs0_2[29:29]),.I5(inf_abs0_2[30:30]),.LO(r_4_3_27_758_i_m2));
defparam desc704.INIT=64'h00FFCCCCF0F0AAAA;
  LUT3 desc705(.I0(inf_abs0_2[19:19]),.I1(inf_abs0_2[20:20]),.I2(inf_abs0_2[31:31]),.O(N_1901));
defparam desc705.INIT=8'h0E;
  LUT5 desc706(.I0(datai[5:5]),.I1(inf_abs0_2[5:5]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[27:27]),.I4(inf_abs0_2[28:28]),.O(m_2[5:5]));
defparam desc706.INIT=32'hCACACACC;
  LUT5 desc707(.I0(datai[8:8]),.I1(inf_abs0_2[8:8]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[27:27]),.I4(inf_abs0_2[28:28]),.O(m_2[8:8]));
defparam desc707.INIT=32'hCACACACC;
  LUT5 desc708(.I0(datai[15:15]),.I1(inf_abs0_2[15:15]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[27:27]),.I4(inf_abs0_2[28:28]),.O(m_2[15:15]));
defparam desc708.INIT=32'hCACACACC;
  LUT5 desc709(.I0(datai[16:16]),.I1(inf_abs0_2[16:16]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[27:27]),.I4(inf_abs0_2[28:28]),.O(m_2[16:16]));
defparam desc709.INIT=32'hCACACACC;
  LUT5 desc710(.I0(datai[3:3]),.I1(inf_abs0_2[3:3]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[27:27]),.I4(inf_abs0_2[28:28]),.O(m_2[3:3]));
defparam desc710.INIT=32'hCACACACC;
  LUT5 desc711(.I0(datai[1:1]),.I1(inf_abs0_2[1:1]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[27:27]),.I4(inf_abs0_2[28:28]),.O(m_2[1:1]));
defparam desc711.INIT=32'hCACACACC;
  LUT5_L desc712(.I0(reg0[31:31]),.I1(reg1[31:31]),.I2(reg2[31:31]),.I3(inf_abs0_2[29:29]),.I4(inf_abs0_2[30:30]),.LO(r_4_3_8_1467));
defparam desc712.INIT=32'h00F0CCAA;
  LUT5 desc713(.I0(datai[13:13]),.I1(inf_abs0_2[13:13]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[27:27]),.I4(inf_abs0_2[28:28]),.O(m_2[13:13]));
defparam desc713.INIT=32'hCACACACC;
  LUT5 desc714(.I0(datai[19:19]),.I1(inf_abs0_2[19:19]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[27:27]),.I4(inf_abs0_2[28:28]),.O(m_2[19:19]));
defparam desc714.INIT=32'hCACACACC;
  LUT5 desc715(.I0(datai[14:14]),.I1(inf_abs0_2[14:14]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[27:27]),.I4(inf_abs0_2[28:28]),.O(m_2[14:14]));
defparam desc715.INIT=32'hCACACACC;
  LUT5 desc716(.I0(datai[18:18]),.I1(inf_abs0_2[18:18]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[27:27]),.I4(inf_abs0_2[28:28]),.O(m_2[18:18]));
defparam desc716.INIT=32'hCACACACC;
  LUT5 desc717(.I0(datai[12:12]),.I1(inf_abs0_2[12:12]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[27:27]),.I4(inf_abs0_2[28:28]),.O(m_2[12:12]));
defparam desc717.INIT=32'hCACACACC;
  LUT5 desc718(.I0(datai[17:17]),.I1(inf_abs0_2[17:17]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[27:27]),.I4(inf_abs0_2[28:28]),.O(m_2[17:17]));
defparam desc718.INIT=32'hCACACACC;
  LUT5 desc719(.I0(datai[10:10]),.I1(inf_abs0_2[10:10]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[27:27]),.I4(inf_abs0_2[28:28]),.O(m_2[10:10]));
defparam desc719.INIT=32'hCACACACC;
  LUT5 desc720(.I0(datai[11:11]),.I1(inf_abs0_2[11:11]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[27:27]),.I4(inf_abs0_2[28:28]),.O(m_2[11:11]));
defparam desc720.INIT=32'hCACACACC;
  LUT5 desc721(.I0(datai[9:9]),.I1(inf_abs0_2[9:9]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[27:27]),.I4(inf_abs0_2[28:28]),.O(m_2[9:9]));
defparam desc721.INIT=32'hCACACACC;
  LUT5 desc722(.I0(datai[2:2]),.I1(inf_abs0_2[2:2]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[27:27]),.I4(inf_abs0_2[28:28]),.O(m_2[2:2]));
defparam desc722.INIT=32'hCACACACC;
  LUT5 desc723(.I0(datai[6:6]),.I1(inf_abs0_2[6:6]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[27:27]),.I4(inf_abs0_2[28:28]),.O(m_2[6:6]));
defparam desc723.INIT=32'hCACACACC;
  LUT5 desc724(.I0(datai[7:7]),.I1(inf_abs0_2[7:7]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[27:27]),.I4(inf_abs0_2[28:28]),.O(m_2[7:7]));
defparam desc724.INIT=32'hCACACACC;
  LUT5 desc725(.I0(datai[4:4]),.I1(inf_abs0_2[4:4]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[27:27]),.I4(inf_abs0_2[28:28]),.O(m_2[4:4]));
defparam desc725.INIT=32'hCACACACC;
  LUT5_L desc726(.I0(reg3[11:11]),.I1(state),.I2(inf_abs0_2[11:11]),.I3(inf_abs0_2[28:28]),.I4(N_2641),.LO(\d_cnst_sn.addr_20_iv_18_335_i_1 ));
defparam desc726.INIT=32'hFFFF111D;
  LUT5_L desc727(.I0(reg3[6:6]),.I1(state),.I2(inf_abs0_2[6:6]),.I3(inf_abs0_2[28:28]),.I4(N_2641),.LO(\d_cnst_sn.addr_20_iv_13_470_i_1 ));
defparam desc727.INIT=32'hFFFF111D;
  LUT5_L desc728(.I0(reg3[10:10]),.I1(state),.I2(inf_abs0_2[10:10]),.I3(inf_abs0_2[28:28]),.I4(N_2641),.LO(\d_cnst_sn.addr_20_iv_17_362_i_1 ));
defparam desc728.INIT=32'hFFFF111D;
  LUT5_L desc729(.I0(reg3[8:8]),.I1(state),.I2(inf_abs0_2[8:8]),.I3(inf_abs0_2[28:28]),.I4(N_2641),.LO(\d_cnst_sn.addr_20_iv_15_416_i_1 ));
defparam desc729.INIT=32'hFFFF111D;
  LUT5_L desc730(.I0(reg3[3:3]),.I1(state),.I2(inf_abs0_2[3:3]),.I3(inf_abs0_2[28:28]),.I4(N_2641),.LO(\d_cnst_sn.addr_20_iv_10_562_i_1 ));
defparam desc730.INIT=32'hFFFF111D;
  LUT5_L desc731(.I0(reg3[5:5]),.I1(state),.I2(inf_abs0_2[5:5]),.I3(inf_abs0_2[28:28]),.I4(N_2641),.LO(\d_cnst_sn.addr_20_iv_12_497_i_1 ));
defparam desc731.INIT=32'hFFFF111D;
  LUT5_L desc732(.I0(reg3[9:9]),.I1(state),.I2(inf_abs0_2[9:9]),.I3(inf_abs0_2[28:28]),.I4(N_2641),.LO(\d_cnst_sn.addr_20_iv_16_389_i_1 ));
defparam desc732.INIT=32'hFFFF111D;
  LUT6 desc733(.I0(reg3[1:1]),.I1(state),.I2(inf_abs0_2[1:1]),.I3(un1_inf_abs0_11[1:1]),.I4(inf_abs0_2[27:27]),.I5(inf_abs0_2[28:28]),.O(\d_cnst_sn.addr_20_iv_8_627_i_1 ));
defparam desc733.INIT=64'h111111DD1D1D1DDD;
  LUT4 desc734(.I0(reg0[4:4]),.I1(reg2[4:4]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[30:30]),.O(N_919));
defparam desc734.INIT=16'hACAA;
  LUT4 desc735(.I0(reg0[3:3]),.I1(reg2[3:3]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[30:30]),.O(N_918));
defparam desc735.INIT=16'hACAA;
  LUT5 desc736(.I0(inf_abs0_2[19:19]),.I1(inf_abs0_2[20:20]),.I2(inf_abs0_2[21:21]),.I3(inf_abs0_2[22:22]),.I4(inf_abs0_2[31:31]),.O(N_1890));
defparam desc736.INIT=32'hFFFFFFFD;
  LUT4 desc737(.I0(inf_abs0_2[24:24]),.I1(inf_abs0_2[25:25]),.I2(inf_abs0_2[26:26]),.I3(inf_abs0_2[31:31]),.O(un36_df));
defparam desc737.INIT=16'h0080;
  LUT5 desc738(.I0(datai[0:0]),.I1(inf_abs0_2[0:0]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[27:27]),.I4(inf_abs0_2[28:28]),.O(m_2[0:0]));
defparam desc738.INIT=32'hCACACACC;
  LUT6 desc739(.I0(datai[30:30]),.I1(inf_abs0_2[20:20]),.I2(inf_abs0_2[21:21]),.I3(inf_abs0_2[22:22]),.I4(inf_abs0_2[31:31]),.I5(g0_2_0_i2_lut6_2_O6),.O(N_3568));
defparam desc739.INIT=64'h0000000000000008;
  LUT4 reg3_1_1_axb_31_cZ(.I0(datai[31:31]),.I1(inf_abs0_2[31:31]),.I2(inf_abs0_2[27:27]),.I3(inf_abs0_2[28:28]),.O(reg3_1_1_axb_31));
defparam reg3_1_1_axb_31_cZ.INIT=16'hDDDF;
  LUT6 desc740(.I0(reg0[29:29]),.I1(reg1[29:29]),.I2(reg2[29:29]),.I3(un3_reg3_cry_25),.I4(N_3_0),.I5(N_13),.O(r_4[29:29]));
defparam desc740.INIT=64'hF0F0AAAAFF00CCCC;
  LUT6_L desc741(.I0(reg0[2:2]),.I1(reg1[2:2]),.I2(reg2[2:2]),.I3(reg3[2:2]),.I4(inf_abs0_2[29:29]),.I5(inf_abs0_2[30:30]),.LO(N_36_i));
defparam desc741.INIT=64'hFF00F0F0CCCCAAAA;
  LUT6 un11_reg0_axb_19_cZ(.I0(datai[19:19]),.I1(inf_abs0_2[19:19]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[27:27]),.I4(inf_abs0_2[28:28]),.I5(r_4[19:19]),.O(un11_reg0_axb_19));
defparam un11_reg0_axb_19_cZ.INIT=64'h35353533CACACACC;
  LUT6 un11_reg0_axb_18_cZ(.I0(datai[18:18]),.I1(inf_abs0_2[18:18]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[27:27]),.I4(inf_abs0_2[28:28]),.I5(r_4[18:18]),.O(un11_reg0_axb_18));
defparam un11_reg0_axb_18_cZ.INIT=64'h35353533CACACACC;
  LUT6 un11_reg0_axb_17_cZ(.I0(datai[17:17]),.I1(inf_abs0_2[17:17]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[27:27]),.I4(inf_abs0_2[28:28]),.I5(r_4[17:17]),.O(un11_reg0_axb_17));
defparam un11_reg0_axb_17_cZ.INIT=64'h35353533CACACACC;
  LUT6 un11_reg0_axb_16_cZ(.I0(datai[16:16]),.I1(inf_abs0_2[16:16]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[27:27]),.I4(inf_abs0_2[28:28]),.I5(r_4[16:16]),.O(un11_reg0_axb_16));
defparam un11_reg0_axb_16_cZ.INIT=64'h35353533CACACACC;
  LUT6 un11_reg0_axb_15_cZ(.I0(datai[15:15]),.I1(inf_abs0_2[15:15]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[27:27]),.I4(inf_abs0_2[28:28]),.I5(r_4[15:15]),.O(un11_reg0_axb_15));
defparam un11_reg0_axb_15_cZ.INIT=64'h35353533CACACACC;
  LUT6 un11_reg0_axb_14_cZ(.I0(datai[14:14]),.I1(inf_abs0_2[14:14]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[27:27]),.I4(inf_abs0_2[28:28]),.I5(r_4[14:14]),.O(un11_reg0_axb_14));
defparam un11_reg0_axb_14_cZ.INIT=64'h35353533CACACACC;
  LUT6 un11_reg0_axb_13_cZ(.I0(datai[13:13]),.I1(inf_abs0_2[13:13]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[27:27]),.I4(inf_abs0_2[28:28]),.I5(r_4[13:13]),.O(un11_reg0_axb_13));
defparam un11_reg0_axb_13_cZ.INIT=64'h35353533CACACACC;
  LUT6 un11_reg0_axb_12_cZ(.I0(datai[12:12]),.I1(inf_abs0_2[12:12]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[27:27]),.I4(inf_abs0_2[28:28]),.I5(r_4[12:12]),.O(un11_reg0_axb_12));
defparam un11_reg0_axb_12_cZ.INIT=64'h35353533CACACACC;
  LUT6 un11_reg0_axb_11_cZ(.I0(datai[11:11]),.I1(inf_abs0_2[11:11]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[27:27]),.I4(inf_abs0_2[28:28]),.I5(r_4[11:11]),.O(un11_reg0_axb_11));
defparam un11_reg0_axb_11_cZ.INIT=64'h35353533CACACACC;
  LUT6 un11_reg0_axb_10_cZ(.I0(datai[10:10]),.I1(inf_abs0_2[10:10]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[27:27]),.I4(inf_abs0_2[28:28]),.I5(r_4[10:10]),.O(un11_reg0_axb_10));
defparam un11_reg0_axb_10_cZ.INIT=64'h35353533CACACACC;
  LUT6 un11_reg0_axb_9_cZ(.I0(datai[9:9]),.I1(inf_abs0_2[9:9]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[27:27]),.I4(inf_abs0_2[28:28]),.I5(r_4[9:9]),.O(un11_reg0_axb_9));
defparam un11_reg0_axb_9_cZ.INIT=64'h35353533CACACACC;
  LUT6 un11_reg0_axb_8_cZ(.I0(datai[8:8]),.I1(inf_abs0_2[8:8]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[27:27]),.I4(inf_abs0_2[28:28]),.I5(r_4[8:8]),.O(un11_reg0_axb_8));
defparam un11_reg0_axb_8_cZ.INIT=64'h35353533CACACACC;
  LUT6 un11_reg0_axb_7_cZ(.I0(datai[7:7]),.I1(inf_abs0_2[7:7]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[27:27]),.I4(inf_abs0_2[28:28]),.I5(r_4[7:7]),.O(un11_reg0_axb_7));
defparam un11_reg0_axb_7_cZ.INIT=64'h35353533CACACACC;
  LUT6 un11_reg0_axb_6_cZ(.I0(datai[6:6]),.I1(inf_abs0_2[6:6]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[27:27]),.I4(inf_abs0_2[28:28]),.I5(r_4[6:6]),.O(un11_reg0_axb_6));
defparam un11_reg0_axb_6_cZ.INIT=64'h35353533CACACACC;
  LUT6 un11_reg0_axb_5_cZ(.I0(datai[5:5]),.I1(inf_abs0_2[5:5]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[27:27]),.I4(inf_abs0_2[28:28]),.I5(r_4[5:5]),.O(un11_reg0_axb_5));
defparam un11_reg0_axb_5_cZ.INIT=64'h35353533CACACACC;
  LUT6 un11_reg0_axb_4_cZ(.I0(datai[4:4]),.I1(inf_abs0_2[4:4]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[27:27]),.I4(inf_abs0_2[28:28]),.I5(r_4[4:4]),.O(un11_reg0_axb_4));
defparam un11_reg0_axb_4_cZ.INIT=64'h35353533CACACACC;
  LUT6 un11_reg0_axb_3_cZ(.I0(datai[3:3]),.I1(inf_abs0_2[3:3]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[27:27]),.I4(inf_abs0_2[28:28]),.I5(r_4[3:3]),.O(un11_reg0_axb_3));
defparam un11_reg0_axb_3_cZ.INIT=64'h35353533CACACACC;
  LUT6 un11_reg0_axb_2_cZ(.I0(datai[2:2]),.I1(inf_abs0_2[2:2]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[27:27]),.I4(inf_abs0_2[28:28]),.I5(N_28),.O(un11_reg0_axb_2));
defparam un11_reg0_axb_2_cZ.INIT=64'h35353533CACACACC;
  LUT6 un11_reg0_axb_1_cZ(.I0(datai[1:1]),.I1(inf_abs0_2[1:1]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[27:27]),.I4(inf_abs0_2[28:28]),.I5(r_4[1:1]),.O(un11_reg0_axb_1));
defparam un11_reg0_axb_1_cZ.INIT=64'h35353533CACACACC;
  LUT5 reg3_1_1_axb_19_cZ(.I0(datai[19:19]),.I1(inf_abs0_2[19:19]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[27:27]),.I4(inf_abs0_2[28:28]),.O(reg3_1_1_axb_19));
defparam reg3_1_1_axb_19_cZ.INIT=32'h35353533;
  LUT5 reg3_1_1_axb_18_cZ(.I0(datai[18:18]),.I1(inf_abs0_2[18:18]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[27:27]),.I4(inf_abs0_2[28:28]),.O(reg3_1_1_axb_18));
defparam reg3_1_1_axb_18_cZ.INIT=32'h35353533;
  LUT5 reg3_1_1_axb_17_cZ(.I0(datai[17:17]),.I1(inf_abs0_2[17:17]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[27:27]),.I4(inf_abs0_2[28:28]),.O(reg3_1_1_axb_17));
defparam reg3_1_1_axb_17_cZ.INIT=32'h35353533;
  LUT5 reg3_1_1_axb_16_cZ(.I0(datai[16:16]),.I1(inf_abs0_2[16:16]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[27:27]),.I4(inf_abs0_2[28:28]),.O(reg3_1_1_axb_16));
defparam reg3_1_1_axb_16_cZ.INIT=32'h35353533;
  LUT5 reg3_1_1_axb_15_cZ(.I0(datai[15:15]),.I1(inf_abs0_2[15:15]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[27:27]),.I4(inf_abs0_2[28:28]),.O(reg3_1_1_axb_15));
defparam reg3_1_1_axb_15_cZ.INIT=32'h35353533;
  LUT5 reg3_1_1_axb_14_cZ(.I0(datai[14:14]),.I1(inf_abs0_2[14:14]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[27:27]),.I4(inf_abs0_2[28:28]),.O(reg3_1_1_axb_14));
defparam reg3_1_1_axb_14_cZ.INIT=32'h35353533;
  LUT5 reg3_1_1_axb_13_cZ(.I0(datai[13:13]),.I1(inf_abs0_2[13:13]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[27:27]),.I4(inf_abs0_2[28:28]),.O(reg3_1_1_axb_13));
defparam reg3_1_1_axb_13_cZ.INIT=32'h35353533;
  LUT5 reg3_1_1_axb_12_cZ(.I0(datai[12:12]),.I1(inf_abs0_2[12:12]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[27:27]),.I4(inf_abs0_2[28:28]),.O(reg3_1_1_axb_12));
defparam reg3_1_1_axb_12_cZ.INIT=32'h35353533;
  LUT5 reg3_1_1_axb_11_cZ(.I0(datai[11:11]),.I1(inf_abs0_2[11:11]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[27:27]),.I4(inf_abs0_2[28:28]),.O(reg3_1_1_axb_11));
defparam reg3_1_1_axb_11_cZ.INIT=32'h35353533;
  LUT5 reg3_1_1_axb_10_cZ(.I0(datai[10:10]),.I1(inf_abs0_2[10:10]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[27:27]),.I4(inf_abs0_2[28:28]),.O(reg3_1_1_axb_10));
defparam reg3_1_1_axb_10_cZ.INIT=32'h35353533;
  LUT5 reg3_1_1_axb_9_cZ(.I0(datai[9:9]),.I1(inf_abs0_2[9:9]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[27:27]),.I4(inf_abs0_2[28:28]),.O(reg3_1_1_axb_9));
defparam reg3_1_1_axb_9_cZ.INIT=32'h35353533;
  LUT5 reg3_1_1_axb_8_cZ(.I0(datai[8:8]),.I1(inf_abs0_2[8:8]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[27:27]),.I4(inf_abs0_2[28:28]),.O(reg3_1_1_axb_8));
defparam reg3_1_1_axb_8_cZ.INIT=32'h35353533;
  LUT5 reg3_1_1_axb_7_cZ(.I0(datai[7:7]),.I1(inf_abs0_2[7:7]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[27:27]),.I4(inf_abs0_2[28:28]),.O(reg3_1_1_axb_7));
defparam reg3_1_1_axb_7_cZ.INIT=32'h35353533;
  LUT5 reg3_1_1_axb_6_cZ(.I0(datai[6:6]),.I1(inf_abs0_2[6:6]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[27:27]),.I4(inf_abs0_2[28:28]),.O(reg3_1_1_axb_6));
defparam reg3_1_1_axb_6_cZ.INIT=32'h35353533;
  LUT5 reg3_1_1_axb_5_cZ(.I0(datai[5:5]),.I1(inf_abs0_2[5:5]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[27:27]),.I4(inf_abs0_2[28:28]),.O(reg3_1_1_axb_5));
defparam reg3_1_1_axb_5_cZ.INIT=32'h35353533;
  LUT5 reg3_1_1_axb_4_cZ(.I0(datai[4:4]),.I1(inf_abs0_2[4:4]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[27:27]),.I4(inf_abs0_2[28:28]),.O(reg3_1_1_axb_4));
defparam reg3_1_1_axb_4_cZ.INIT=32'h35353533;
  LUT5 reg3_1_1_axb_3_cZ(.I0(datai[3:3]),.I1(inf_abs0_2[3:3]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[27:27]),.I4(inf_abs0_2[28:28]),.O(reg3_1_1_axb_3));
defparam reg3_1_1_axb_3_cZ.INIT=32'h35353533;
  LUT5 reg3_1_1_axb_2_cZ(.I0(datai[2:2]),.I1(inf_abs0_2[2:2]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[27:27]),.I4(inf_abs0_2[28:28]),.O(reg3_1_1_axb_2));
defparam reg3_1_1_axb_2_cZ.INIT=32'h35353533;
  LUT5 reg3_1_1_axb_1_cZ(.I0(datai[1:1]),.I1(inf_abs0_2[1:1]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[27:27]),.I4(inf_abs0_2[28:28]),.O(reg3_1_1_axb_1));
defparam reg3_1_1_axb_1_cZ.INIT=32'h35353533;
  LUT6 desc742(.I0(reg0[31:31]),.I1(reg1[31:31]),.I2(reg2[31:31]),.I3(inf_abs0_2[31:31]),.I4(inf_abs0_2[29:29]),.I5(inf_abs0_2[30:30]),.O(r_4[31:31]));
defparam desc742.INIT=64'hAA00AAF0AACCAAAA;
  LUT4 desc743(.I0(inf_abs0_2[24:24]),.I1(inf_abs0_2[25:25]),.I2(inf_abs0_2[26:26]),.I3(inf_abs0_2[31:31]),.O(d_cnst_sm0));
defparam desc743.INIT=16'h00BC;
  LUT6 desc744(.I0(datai[19:19]),.I1(inf_abs0_2[19:19]),.I2(inf_abs0_2[20:20]),.I3(inf_abs0_2[31:31]),.I4(N_3873_2),.I5(g0_2_0_i2_lut6_2_O6),.O(\d_cnst_sn.reg0_28_3_2492_0 ));
defparam desc744.INIT=64'h00CC000000A00000;
  LUT6 desc745(.I0(reg1[0:0]),.I1(reg3[0:0]),.I2(state),.I3(inf_abs0_2[0:0]),.I4(inf_abs0_2[27:27]),.I5(inf_abs0_2[28:28]),.O(\d_cnst_sn.addr_20_iv_7_654_i_1 ));
defparam desc745.INIT=64'h0303A35303F3A3F3;
  LUT5 desc746(.I0(inf_abs0_2[24:24]),.I1(inf_abs0_2[25:25]),.I2(inf_abs0_2[26:26]),.I3(inf_abs0_2[22:22]),.I4(inf_abs0_2[31:31]),.O(\d_cnst_sn.reg3_5_sqmuxa_2_1 ));
defparam desc746.INIT=32'hFFFF007F;
  LUT5 desc747(.I0(inf_abs0_2[21:21]),.I1(inf_abs0_2[22:22]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[28:28]),.I4(r_4[28:28]),.O(reg2_16_11_a1[29:29]));
defparam desc747.INIT=32'h08000000;
  LUT6 desc748(.I0(N_3913),.I1(N_512_i),.I2(N_513_i),.I3(un11_r_cry[30:30]),.I4(un14_r_0_I_83),.I5(N_895),.O(N_3912));
defparam desc748.INIT=64'h5556595AA5A6A9AA;
  LUT6 un11_reg0_axb_0_cZ(.I0(datai[0:0]),.I1(inf_abs0_2[0:0]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[27:27]),.I4(inf_abs0_2[28:28]),.I5(r_4[0:0]),.O(un11_reg0_axb_0));
defparam un11_reg0_axb_0_cZ.INIT=64'h35353533CACACACC;
  LUT6 un3_t_axb_30_cZ(.I0(reg0[30:30]),.I1(reg1[30:30]),.I2(reg2[30:30]),.I3(inf_abs0_2[31:31]),.I4(inf_abs0_2[29:29]),.I5(inf_abs0_2[30:30]),.O(un3_t_axb_30));
defparam un3_t_axb_30_cZ.INIT=64'h55FF550F55335555;
  LUT6 un3_t_axb_29_cZ(.I0(reg0[29:29]),.I1(reg1[29:29]),.I2(reg2[29:29]),.I3(un3_reg3_cry_25),.I4(N_3_0),.I5(N_13),.O(un3_t_axb_29));
defparam un3_t_axb_29_cZ.INIT=64'h0F0F555500FF3333;
  LUT5 reg3_1_1_axb_0_cZ(.I0(datai[0:0]),.I1(inf_abs0_2[0:0]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[27:27]),.I4(inf_abs0_2[28:28]),.O(reg3_1_1_axb_0));
defparam reg3_1_1_axb_0_cZ.INIT=32'h35353533;
  LUT5 desc749(.I0(inf_abs0_2[24:24]),.I1(inf_abs0_2[23:23]),.I2(inf_abs0_2[25:25]),.I3(inf_abs0_2[26:26]),.I4(inf_abs0_2[31:31]),.O(addr_4_sqmuxa_1_1));
defparam desc749.INIT=32'h00002000;
  LUT6 desc750(.I0(reg0[31:31]),.I1(reg1[31:31]),.I2(reg2[31:31]),.I3(inf_abs0_2[31:31]),.I4(inf_abs0_2[29:29]),.I5(inf_abs0_2[30:30]),.O(r_4_i[31:31]));
defparam desc750.INIT=64'h55FF550F55335555;
  LUT6 un3_t_axb_31_cZ(.I0(reg0[31:31]),.I1(reg1[31:31]),.I2(reg2[31:31]),.I3(inf_abs0_2[31:31]),.I4(inf_abs0_2[29:29]),.I5(inf_abs0_2[30:30]),.O(un3_t_axb_31));
defparam un3_t_axb_31_cZ.INIT=64'h55FF550F55335555;
  LUT6 desc751(.I0(reg2[0:0]),.I1(reg1[0:0]),.I2(inf_abs0_2[0:0]),.I3(inf_abs0_2[31:31]),.I4(inf_abs0_2[27:27]),.I5(inf_abs0_2[28:28]),.O(N_2240_i));
defparam desc751.INIT=64'hF05AF03CF0F0F0F0;
  LUT6 desc752(.I0(b),.I1(inf_abs0_2[21:21]),.I2(inf_abs0_2[22:22]),.I3(inf_abs0_2[31:31]),.I4(inf_abs0_2[27:27]),.I5(inf_abs0_2[28:28]),.O(\d_cnst_sn.reg0_28_14_2135_1_a0_2 ));
defparam desc752.INIT=64'h00000000004000C0;
  LUT6 desc753(.I0(N_512_i),.I1(N_513_i),.I2(N_514_i),.I3(m_2[25:25]),.I4(N_527_i),.I5(r_4[24:24]),.O(\d_cnst_sn.reg2_16_0 [25:25]));
defparam desc753.INIT=64'hFFFDFFFD3F3DFFFD;
  LUT6 desc754(.I0(N_512_i),.I1(N_513_i),.I2(N_514_i),.I3(m_2[24:24]),.I4(N_527_i),.I5(r_4[23:23]),.O(\d_cnst_sn.reg2_16_0 [24:24]));
defparam desc754.INIT=64'hFFFDFFFD3F3DFFFD;
  LUT6 desc755(.I0(N_512_i),.I1(N_513_i),.I2(N_514_i),.I3(m_2[23:23]),.I4(N_527_i),.I5(r_4[22:22]),.O(\d_cnst_sn.reg2_16_0 [23:23]));
defparam desc755.INIT=64'hFFFDFFFD3F3DFFFD;
  LUT6 desc756(.I0(N_512_i),.I1(N_513_i),.I2(N_514_i),.I3(m_2[22:22]),.I4(N_527_i),.I5(r_4[21:21]),.O(\d_cnst_sn.reg2_16_0 [22:22]));
defparam desc756.INIT=64'hFFFDFFFD3F3DFFFD;
  LUT6_L desc757(.I0(N_512_i),.I1(N_513_i),.I2(N_514_i),.I3(m_2[21:21]),.I4(N_527_i),.I5(r_4[20:20]),.LO(\d_cnst_sn.reg2_16_0 [21:21]));
defparam desc757.INIT=64'hFFFDFFFD3F3DFFFD;
  LUT5 desc758(.I0(inf_abs0_2[19:19]),.I1(inf_abs0_2[20:20]),.I2(inf_abs0_2[21:21]),.I3(inf_abs0_2[22:22]),.I4(inf_abs0_2[31:31]),.O(un1_b59));
defparam desc758.INIT=32'h00000AC0;
  LUT5 desc759(.I0(inf_abs0_2[19:19]),.I1(inf_abs0_2[20:20]),.I2(inf_abs0_2[21:21]),.I3(inf_abs0_2[22:22]),.I4(inf_abs0_2[31:31]),.O(un1_b57));
defparam desc759.INIT=32'h00000530;
  LUT5 desc760(.I0(inf_abs0_2[21:21]),.I1(inf_abs0_2[22:22]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[28:28]),.I4(r_4[28:28]),.O(reg0_m9_i_a1));
defparam desc760.INIT=32'h08000000;
  LUT6 desc761(.I0(un3_reg3_cry_25),.I1(N_3913),.I2(N_512_i),.I3(\d_cnst_sn.reg1_16_a2_0 [5:5]),.I4(m_2[29:29]),.I5(reg3_1_1[29:29]),.O(reg2_16_11_a2[29:29]));
defparam desc761.INIT=64'hFE000E00F2000200;
  LUT6 desc762(.I0(state),.I1(inf_abs0_2[24:24]),.I2(inf_abs0_2[23:23]),.I3(inf_abs0_2[25:25]),.I4(inf_abs0_2[26:26]),.I5(inf_abs0_2[31:31]),.O(addr_4_sqmuxa_1));
defparam desc762.INIT=64'h0000000008000000;
  LUT4 desc763(.I0(inf_abs0_2[24:24]),.I1(inf_abs0_2[25:25]),.I2(inf_abs0_2[26:26]),.I3(inf_abs0_2[31:31]),.O(d_cnst));
defparam desc763.INIT=16'h00BA;
  LUT6_L desc764(.I0(inf_abs0_2[28:28]),.I1(un1_inf_abs0_10[10:10]),.I2(un1_inf_abs0_11[10:10]),.I3(N_2660_2),.I4(\d_cnst_sn.addr_20_iv_1052_i_a6_1_0 ),.I5(\d_cnst_sn.addr_20_iv_17_362_i_1 ),.LO(N_2119_i));
defparam desc764.INIT=64'h00000000D0F0DDFF;
  LUT6_L desc765(.I0(inf_abs0_2[28:28]),.I1(un1_inf_abs0_10[9:9]),.I2(un1_inf_abs0_11[9:9]),.I3(N_2660_2),.I4(\d_cnst_sn.addr_20_iv_1052_i_a6_1_0 ),.I5(\d_cnst_sn.addr_20_iv_16_389_i_1 ),.LO(N_2139_i));
defparam desc765.INIT=64'h00000000D0F0DDFF;
  LUT6_L desc766(.I0(state),.I1(inf_abs0_2[27:27]),.I2(inf_abs0_2[28:28]),.I3(un1_inf_abs0_10[8:8]),.I4(un1_inf_abs0_11[8:8]),.I5(\d_cnst_sn.addr_20_iv_15_416_i_1 ),.LO(N_2159_i));
defparam desc766.INIT=64'h00000000FF7FDD5D;
  LUT6_L desc767(.I0(reg3[7:7]),.I1(state),.I2(inf_abs0_2[7:7]),.I3(inf_abs0_2[28:28]),.I4(\d_cnst_sn.addr_20_iv_14_443_i_2 ),.I5(N_2641),.LO(N_2179_i));
defparam desc767.INIT=64'h000000000000EEE2;
  LUT6_L desc768(.I0(state),.I1(inf_abs0_2[27:27]),.I2(inf_abs0_2[28:28]),.I3(un1_inf_abs0_10[6:6]),.I4(un1_inf_abs0_11[6:6]),.I5(\d_cnst_sn.addr_20_iv_13_470_i_1 ),.LO(N_2199_i));
defparam desc768.INIT=64'h00000000FF7FDD5D;
  LUT6_L desc769(.I0(state),.I1(inf_abs0_2[27:27]),.I2(inf_abs0_2[28:28]),.I3(un1_inf_abs0_10[5:5]),.I4(un1_inf_abs0_11[5:5]),.I5(\d_cnst_sn.addr_20_iv_12_497_i_1 ),.LO(N_2219_i));
defparam desc769.INIT=64'h00000000FF7FDD5D;
  LUT6_L desc770(.I0(state),.I1(inf_abs0_2[27:27]),.I2(inf_abs0_2[28:28]),.I3(un1_inf_abs0_10[3:3]),.I4(un1_inf_abs0_11[3:3]),.I5(\d_cnst_sn.addr_20_iv_10_562_i_1 ),.LO(N_2267_i));
defparam desc770.INIT=64'h00000000FF7FDD5D;
  LUT6 desc771(.I0(\d_cnst_sn.reg2_N_3_mux ),.I1(reg2_16_2_d[20:20]),.I2(\d_cnst_sn.reg1_16_a2_0 [5:5]),.I3(\d_cnst_sn.reg0_28_a1_1 [4:4]),.I4(r_4[19:19]),.I5(reg3_1_1[20:20]),.O(\d_cnst_sn.reg2_16_0 [20:20]));
defparam desc771.INIT=64'hEFEF00EF4F4F004F;
  LUT6 desc772(.I0(m_2[2:2]),.I1(m_2[1:1]),.I2(m_2[0:0]),.I3(r_4[0:0]),.I4(r_4[1:1]),.I5(N_28),.O(un14_r_0_N_70));
defparam desc772.INIT=64'h8008200240041001;
  LUT6 desc773(.I0(m_2[15:15]),.I1(m_2[16:16]),.I2(m_2[17:17]),.I3(r_4[15:15]),.I4(r_4[16:16]),.I5(r_4[17:17]),.O(un14_r_0_N_42));
defparam desc773.INIT=64'h8040201008040201;
  LUT6 desc774(.I0(m_2[3:3]),.I1(m_2[4:4]),.I2(m_2[5:5]),.I3(r_4[3:3]),.I4(r_4[4:4]),.I5(r_4[5:5]),.O(un14_r_0_N_14));
defparam desc774.INIT=64'h8040201008040201;
  LUT6 desc775(.I0(m_2[19:19]),.I1(m_2[20:20]),.I2(m_2[18:18]),.I3(r_4[19:19]),.I4(r_4[18:18]),.I5(r_4[20:20]),.O(un14_r_0_N_49));
defparam desc775.INIT=64'h8040080420100201;
  LUT6 desc776(.I0(m_2[12:12]),.I1(m_2[13:13]),.I2(m_2[14:14]),.I3(r_4[12:12]),.I4(r_4[13:13]),.I5(r_4[14:14]),.O(un14_r_0_N_7));
defparam desc776.INIT=64'h8040201008040201;
  LUT6 desc777(.I0(m_2[9:9]),.I1(m_2[10:10]),.I2(m_2[11:11]),.I3(r_4[11:11]),.I4(r_4[9:9]),.I5(r_4[10:10]),.O(un14_r_0_N_28));
defparam desc777.INIT=64'h8008400420021001;
  LUT6 desc778(.I0(m_2[7:7]),.I1(m_2[6:6]),.I2(m_2[8:8]),.I3(r_4[6:6]),.I4(r_4[8:8]),.I5(r_4[7:7]),.O(un14_r_0_N_21));
defparam desc778.INIT=64'h8020080240100401;
  LUT6 desc779(.I0(reg0[30:30]),.I1(reg1[30:30]),.I2(reg2[30:30]),.I3(N_3_0),.I4(r_4[31:31]),.I5(N_13),.O(r_6[30:30]));
defparam desc779.INIT=64'hF0AA000000CC0000;
  LUT6 desc780(.I0(N_3910),.I1(\d_cnst_sn.reg0_28_a0_1 [7:7]),.I2(m_2[7:7]),.I3(\d_cnst_sn.reg0_28_a1_1 [4:4]),.I4(r_4[6:6]),.I5(reg3_1_1[7:7]),.O(\d_cnst_sn.reg0_1 [7:7]));
defparam desc780.INIT=64'hF5F500F531310031;
  LUT6 desc781(.I0(m_2[29:29]),.I1(m_2[27:27]),.I2(m_2[28:28]),.I3(r_4[27:27]),.I4(r_4[28:28]),.I5(r_4[29:29]),.O(un14_r_0_N_63));
defparam desc781.INIT=64'h8020080240100401;
  LUT6 desc782(.I0(N_526_i),.I1(N_1901),.I2(N_513_i),.I3(N_514_i),.I4(un36_df),.I5(N_527_i),.O(b_2_sqmuxa));
defparam desc782.INIT=64'h0000200000000000;
  LUT6_L desc783(.I0(state),.I1(inf_abs0_2[27:27]),.I2(inf_abs0_2[28:28]),.I3(un1_inf_abs0_10[11:11]),.I4(un1_inf_abs0_11[11:11]),.I5(\d_cnst_sn.addr_20_iv_18_335_i_1 ),.LO(N_2099_i));
defparam desc783.INIT=64'h00000000FF7FDD5D;
  LUT6_L desc784(.I0(\d_cnst_sn.addr_20_iv_6_863_i_0 ),.I1(un1_inf_abs0_10[19:19]),.I2(un1_inf_abs0_11[19:19]),.I3(\d_cnst_sn.addr_20_iv_1052_i_a6_1_0 ),.I4(\d_cnst_sn.addr_20_iv_1052_i_a6_2_0 ),.I5(N_2641),.LO(N_2516_i));
defparam desc784.INIT=64'h0000000040445055;
  LUT6_L desc785(.I0(\d_cnst_sn.addr_20_iv_5_890_i_0 ),.I1(un1_inf_abs0_10[18:18]),.I2(un1_inf_abs0_11[18:18]),.I3(\d_cnst_sn.addr_20_iv_1052_i_a6_1_0 ),.I4(\d_cnst_sn.addr_20_iv_1052_i_a6_2_0 ),.I5(N_2641),.LO(N_2536_i));
defparam desc785.INIT=64'h0000000040445055;
  LUT6_L desc786(.I0(\d_cnst_sn.addr_20_iv_4_917_i_0 ),.I1(un1_inf_abs0_10[17:17]),.I2(un1_inf_abs0_11[17:17]),.I3(\d_cnst_sn.addr_20_iv_1052_i_a6_1_0 ),.I4(\d_cnst_sn.addr_20_iv_1052_i_a6_2_0 ),.I5(N_2641),.LO(N_2556_i));
defparam desc786.INIT=64'h0000000040445055;
  LUT6_L desc787(.I0(\d_cnst_sn.addr_20_iv_3_944_i_0 ),.I1(un1_inf_abs0_10[16:16]),.I2(un1_inf_abs0_11[16:16]),.I3(\d_cnst_sn.addr_20_iv_1052_i_a6_1_0 ),.I4(\d_cnst_sn.addr_20_iv_1052_i_a6_2_0 ),.I5(N_2641),.LO(N_2576_i));
defparam desc787.INIT=64'h0000000040445055;
  LUT6_L desc788(.I0(\d_cnst_sn.addr_20_iv_2_971_i_0 ),.I1(un1_inf_abs0_10[15:15]),.I2(un1_inf_abs0_11[15:15]),.I3(\d_cnst_sn.addr_20_iv_1052_i_a6_1_0 ),.I4(\d_cnst_sn.addr_20_iv_1052_i_a6_2_0 ),.I5(N_2641),.LO(N_2596_i));
defparam desc788.INIT=64'h0000000040445055;
  LUT6_L desc789(.I0(\d_cnst_sn.addr_20_iv_1_998_i_0 ),.I1(un1_inf_abs0_10[14:14]),.I2(un1_inf_abs0_11[14:14]),.I3(\d_cnst_sn.addr_20_iv_1052_i_a6_1_0 ),.I4(\d_cnst_sn.addr_20_iv_1052_i_a6_2_0 ),.I5(N_2641),.LO(N_2616_i));
defparam desc789.INIT=64'h0000000040445055;
  LUT6_L desc790(.I0(\d_cnst_sn.addr_20_iv_0_1025_i_0 ),.I1(un1_inf_abs0_10[13:13]),.I2(un1_inf_abs0_11[13:13]),.I3(\d_cnst_sn.addr_20_iv_1052_i_a6_1_0 ),.I4(\d_cnst_sn.addr_20_iv_1052_i_a6_2_0 ),.I5(N_2641),.LO(N_2636_i));
defparam desc790.INIT=64'h0000000040445055;
  LUT6_L desc791(.I0(\d_cnst_sn.addr_20_iv_1052_i_0 ),.I1(un1_inf_abs0_10[12:12]),.I2(un1_inf_abs0_11[12:12]),.I3(\d_cnst_sn.addr_20_iv_1052_i_a6_1_0 ),.I4(\d_cnst_sn.addr_20_iv_1052_i_a6_2_0 ),.I5(N_2641),.LO(N_2656_i));
defparam desc791.INIT=64'h0000000040445055;
  LUT6 desc792(.I0(\d_cnst_sn.reg2_16_0_1_tz [28:28]),.I1(\d_cnst_sn.reg1_16_a2_0 [5:5]),.I2(\d_cnst_sn.reg0_28_a1_1 [4:4]),.I3(r_4[27:27]),.I4(N_1363),.I5(un32_reg0_s_28),.O(\d_cnst_sn.reg2_16_0_1_0 [28:28]));
defparam desc792.INIT=64'hFF0F3303AA0A2202;
  LUT6 desc793(.I0(\d_cnst_sn.reg2_16_0_1_tz [28:28]),.I1(\d_cnst_sn.reg1_16_a2_0 [5:5]),.I2(\d_cnst_sn.reg0_28_a1_1 [4:4]),.I3(r_4[26:26]),.I4(N_1362),.I5(un32_reg0_s_27),.O(\d_cnst_sn.reg2_16_0_1_0 [27:27]));
defparam desc793.INIT=64'hFF0F3303AA0A2202;
  LUT6 desc794(.I0(\d_cnst_sn.reg2_16_0_1_tz [28:28]),.I1(\d_cnst_sn.reg1_16_a2_0 [5:5]),.I2(\d_cnst_sn.reg0_28_a1_1 [4:4]),.I3(r_4[25:25]),.I4(N_1361),.I5(un32_reg0_s_26),.O(\d_cnst_sn.reg2_16_0_1_0 [26:26]));
defparam desc794.INIT=64'hFF0F3303AA0A2202;
  LUT6 desc795(.I0(N_3913),.I1(N_513_i),.I2(N_514_i),.I3(N_1352),.I4(un32_reg0_s_17),.I5(un11_reg0_s_17),.O(reg2_16_11_a3[17:17]));
defparam desc795.INIT=64'h0003101320233033;
  LUT6 desc796(.I0(N_3913),.I1(N_513_i),.I2(N_514_i),.I3(N_1354),.I4(un32_reg0_s_19),.I5(un11_reg0_s_19),.O(reg2_16_11_a3[19:19]));
defparam desc796.INIT=64'h0003101320233033;
  LUT6 desc797(.I0(N_3913),.I1(N_513_i),.I2(N_514_i),.I3(N_1353),.I4(un32_reg0_s_18),.I5(un11_reg0_s_18),.O(reg2_16_11_a3[18:18]));
defparam desc797.INIT=64'h0003101320233033;
  LUT6_L desc798(.I0(inf_abs0_2[22:22]),.I1(reg0_28_sn_m6_lut6_2_O5),.I2(N_513_i),.I3(N_527_i),.I4(N_1493),.I5(t_1[30:30]),.LO(reg2_16[30:30]));
defparam desc798.INIT=64'h0F0F00000F2F0020;
  LUT6 desc799(.I0(\d_cnst_sn.reg0_m9_i_a3_0 ),.I1(N_1033),.I2(\d_cnst_sn.reg0_28_9_2294_a6_3_0 ),.I3(m_2[27:27]),.I4(un32_reg0_s_27),.I5(un11_reg0_s_27),.O(\d_cnst_sn.reg1_16_8_1837_0 ));
defparam desc799.INIT=64'hFAAAF888F222F000;
  LUT6 desc800(.I0(\d_cnst_sn.reg0_m9_i_a3_0 ),.I1(N_1033),.I2(\d_cnst_sn.reg0_28_9_2294_a6_3_0 ),.I3(m_2[26:26]),.I4(un32_reg0_s_26),.I5(un11_reg0_s_26),.O(\d_cnst_sn.reg1_16_7_1870_0 ));
defparam desc800.INIT=64'hFAAAF888F222F000;
  LUT6 desc801(.I0(\d_cnst_sn.reg0_m9_i_a3_0 ),.I1(N_1033),.I2(\d_cnst_sn.reg0_28_9_2294_a6_3_0 ),.I3(m_2[25:25]),.I4(un32_reg0_s_25),.I5(un11_reg0_s_25),.O(\d_cnst_sn.reg0_28_9_2294_0 ));
defparam desc801.INIT=64'hFAAAF888F222F000;
  LUT6 desc802(.I0(\d_cnst_sn.reg0_m9_i_a3_0 ),.I1(N_1033),.I2(\d_cnst_sn.reg0_28_9_2294_a6_3_0 ),.I3(m_2[23:23]),.I4(un32_reg0_s_23),.I5(un11_reg0_s_23),.O(\d_cnst_sn.reg0_28_7_2360_0 ));
defparam desc802.INIT=64'hFAAAF888F222F000;
  LUT6 desc803(.I0(\d_cnst_sn.reg0_m9_i_a3_0 ),.I1(N_1033),.I2(\d_cnst_sn.reg0_28_9_2294_a6_3_0 ),.I3(m_2[22:22]),.I4(un32_reg0_s_22),.I5(un11_reg0_s_22),.O(\d_cnst_sn.reg0_28_6_2393_0 ));
defparam desc803.INIT=64'hFAAAF888F222F000;
  LUT6 desc804(.I0(\d_cnst_sn.reg0_m9_i_a3_0 ),.I1(N_1033),.I2(\d_cnst_sn.reg0_28_9_2294_a6_3_0 ),.I3(m_2[21:21]),.I4(un32_reg0_s_21),.I5(un11_reg0_s_21),.O(\d_cnst_sn.reg0_28_5_2426_0 ));
defparam desc804.INIT=64'hFAAAF888F222F000;
  LUT6 desc805(.I0(\d_cnst_sn.reg0_m9_i_a3_0 ),.I1(N_1033),.I2(\d_cnst_sn.reg0_28_9_2294_a6_3_0 ),.I3(m_2[24:24]),.I4(un32_reg0_s_24),.I5(un11_reg0_s_24),.O(\d_cnst_sn.reg0_28_8_2327_0 ));
defparam desc805.INIT=64'hFAAAF888F222F000;
  LUT6 desc806(.I0(\d_cnst_sn.reg0_m9_i_a3_0 ),.I1(N_1033),.I2(\d_cnst_sn.reg0_28_9_2294_a6_3_0 ),.I3(m_2[20:20]),.I4(un32_reg0_s_20),.I5(un11_reg0_s_20),.O(\d_cnst_sn.reg0_28_4_2459_0 ));
defparam desc806.INIT=64'hFAAAF888F222F000;
  LUT5 desc807(.I0(\d_cnst_sn.reg0_m9_i_a3_0 ),.I1(N_1033),.I2(\d_cnst_sn.reg0_28_3_2492_0 ),.I3(un32_reg0_s_19),.I4(un11_reg0_s_19),.O(\d_cnst_sn.reg0_28_3_2492_1 ));
defparam desc807.INIT=32'hFAF8F2F0;
  LUT6 desc808(.I0(N_512_i),.I1(\d_cnst_sn.b60_0 ),.I2(reg2_16_11_a1[29:29]),.I3(reg2_16_11_a2[29:29]),.I4(un32_reg0_s_29),.I5(un11_reg0_s_29),.O(\d_cnst_sn.reg2_16_1 [29:29]));
defparam desc808.INIT=64'hFFFCFFF4FFF8FFF0;
  LUT6_L desc809(.I0(N_513_i),.I1(N_514_i),.I2(N_1338),.I3(N_1370),.I4(N_1562),.I5(t_6[3:3]),.LO(reg2_16[3:3]));
defparam desc809.INIT=64'hFEBADC9876325410;
  LUT6_L desc810(.I0(N_513_i),.I1(N_514_i),.I2(N_1339),.I3(N_1371),.I4(N_1563),.I5(t_6[4:4]),.LO(reg2_16[4:4]));
defparam desc810.INIT=64'hFEBADC9876325410;
  LUT6_L desc811(.I0(N_513_i),.I1(N_514_i),.I2(N_1340),.I3(N_1372),.I4(N_1564),.I5(t_6[5:5]),.LO(reg2_16[5:5]));
defparam desc811.INIT=64'hFEBADC9876325410;
  LUT6_L desc812(.I0(N_513_i),.I1(N_514_i),.I2(N_1341),.I3(N_1373),.I4(N_1565),.I5(t_6[6:6]),.LO(reg2_16[6:6]));
defparam desc812.INIT=64'hFEBADC9876325410;
  LUT6_L desc813(.I0(N_513_i),.I1(N_514_i),.I2(N_1344),.I3(N_1376),.I4(N_1568),.I5(t_6[9:9]),.LO(reg2_16[9:9]));
defparam desc813.INIT=64'hFEBADC9876325410;
  LUT6_L desc814(.I0(N_513_i),.I1(N_514_i),.I2(N_1345),.I3(N_1377),.I4(N_1569),.I5(t_6[10:10]),.LO(reg2_16[10:10]));
defparam desc814.INIT=64'hFEBADC9876325410;
  LUT6_L desc815(.I0(N_513_i),.I1(N_514_i),.I2(N_1346),.I3(N_1378),.I4(N_1570),.I5(t_6[11:11]),.LO(reg2_16[11:11]));
defparam desc815.INIT=64'hFEBADC9876325410;
  LUT6_L desc816(.I0(N_513_i),.I1(N_514_i),.I2(N_1347),.I3(N_1379),.I4(N_1571),.I5(t_6[12:12]),.LO(reg2_16[12:12]));
defparam desc816.INIT=64'hFEBADC9876325410;
  LUT6_L desc817(.I0(N_513_i),.I1(N_514_i),.I2(N_1348),.I3(N_1380),.I4(N_1572),.I5(t_6[13:13]),.LO(reg2_16[13:13]));
defparam desc817.INIT=64'hFEBADC9876325410;
  LUT6_L desc818(.I0(N_513_i),.I1(N_514_i),.I2(N_1349),.I3(N_1381),.I4(N_1573),.I5(t_6[14:14]),.LO(reg2_16[14:14]));
defparam desc818.INIT=64'hFEBADC9876325410;
  LUT6_L desc819(.I0(N_513_i),.I1(N_514_i),.I2(N_1350),.I3(N_1382),.I4(N_1574),.I5(t_6[15:15]),.LO(reg2_16[15:15]));
defparam desc819.INIT=64'hFEBADC9876325410;
  LUT6_L desc820(.I0(N_513_i),.I1(N_514_i),.I2(N_1351),.I3(N_1383),.I4(N_1575),.I5(t_6[16:16]),.LO(reg2_16[16:16]));
defparam desc820.INIT=64'hFEBADC9876325410;
  LUT6_L desc821(.I0(state),.I1(N_7_i),.I2(N_513_i),.I3(N_514_i),.I4(un36_df),.I5(m7),.LO(rd_18));
defparam desc821.INIT=64'h55555555DDDDDFFF;
  LUT6_L desc822(.I0(N_513_i),.I1(N_514_i),.I2(N_1343),.I3(N_1375),.I4(N_1567),.I5(t_6[8:8]),.LO(reg2_16[8:8]));
defparam desc822.INIT=64'hFEBADC9876325410;
  LUT6_L desc823(.I0(N_513_i),.I1(N_514_i),.I2(N_1337),.I3(N_1369),.I4(N_1561),.I5(t_6[2:2]),.LO(reg2_16[2:2]));
defparam desc823.INIT=64'hFEBADC9876325410;
  LUT6_L desc824(.I0(N_513_i),.I1(N_514_i),.I2(N_1342),.I3(N_1374),.I4(N_1566),.I5(t_6[7:7]),.LO(reg2_16[7:7]));
defparam desc824.INIT=64'hFEBADC9876325410;
  LUT6 desc825(.I0(state),.I1(N_7_i),.I2(N_513_i),.I3(N_514_i),.I4(un36_df),.I5(m7),.O(addr_0_sqmuxa_1_i));
defparam desc825.INIT=64'h77775555FFFFDFFF;
  LUT6 desc826(.I0(\d_cnst_sn.reg0_28_12_2195_a6_1_2_0 ),.I1(\d_cnst_sn.reg0_m8_e_0 ),.I2(N_513_i),.I3(N_527_i),.I4(r_4[27:27]),.I5(reg3_1_1[28:28]),.O(\d_cnst_sn.reg1_16_9_1804_3_tz ));
defparam desc826.INIT=64'hBBBBABBBB0B0A0B0;
  LUT6_L desc827(.I0(\d_cnst_sn.reg0_28_a1_1 [4:4]),.I1(\d_cnst_sn.reg1_16_a0_1 [3:3]),.I2(r_4[16:16]),.I3(t_1[17:17]),.I4(reg2_16_11_a2[17:17]),.I5(reg2_16_11_a3[17:17]),.LO(reg2_16[17:17]));
defparam desc827.INIT=64'h00000000000031F5;
  LUT6_L desc828(.I0(\d_cnst_sn.reg0_28_a1_1 [4:4]),.I1(\d_cnst_sn.reg1_16_a0_1 [3:3]),.I2(r_4[18:18]),.I3(t_1[19:19]),.I4(reg2_16_11_a2[19:19]),.I5(reg2_16_11_a3[19:19]),.LO(reg2_16[19:19]));
defparam desc828.INIT=64'h00000000000031F5;
  LUT6_L desc829(.I0(\d_cnst_sn.reg0_28_a1_1 [4:4]),.I1(\d_cnst_sn.reg1_16_a0_1 [3:3]),.I2(r_4[17:17]),.I3(t_1[18:18]),.I4(reg2_16_11_a2[18:18]),.I5(reg2_16_11_a3[18:18]),.LO(reg2_16[18:18]));
defparam desc829.INIT=64'h00000000000031F5;
  LUT6_L desc830(.I0(\d_cnst_sn.reg2_16_11_1_tz [28:28]),.I1(\d_cnst_sn.reg1_16_a0_1 [3:3]),.I2(\d_cnst_sn.reg2_16_0 [20:20]),.I3(un11_reg0_s_20),.I4(\d_cnst_sn.reg2_16_1 [20:20]),.I5(t_1[20:20]),.LO(reg2_16[20:20]));
defparam desc830.INIT=64'h30200000F0A00000;
  LUT5_L desc831(.I0(\d_cnst_sn.reg2_16_11_1_tz [28:28]),.I1(\d_cnst_sn.reg1_16_a0_1 [3:3]),.I2(un11_reg0_s_28),.I3(\d_cnst_sn.reg2_16_0_1_0 [28:28]),.I4(t_1[28:28]),.LO(reg2_16[28:28]));
defparam desc831.INIT=32'h3200FA00;
  LUT5_L desc832(.I0(\d_cnst_sn.reg2_16_11_1_tz [28:28]),.I1(\d_cnst_sn.reg1_16_a0_1 [3:3]),.I2(un11_reg0_s_27),.I3(\d_cnst_sn.reg2_16_0_1_0 [27:27]),.I4(t_1[27:27]),.LO(reg2_16[27:27]));
defparam desc832.INIT=32'h3200FA00;
  LUT5_L desc833(.I0(\d_cnst_sn.reg2_16_11_1_tz [28:28]),.I1(\d_cnst_sn.reg1_16_a0_1 [3:3]),.I2(un11_reg0_s_26),.I3(\d_cnst_sn.reg2_16_0_1_0 [26:26]),.I4(t_1[26:26]),.LO(reg2_16[26:26]));
defparam desc833.INIT=32'h3200FA00;
  LUT5_L desc834(.I0(d[0:0]),.I1(d[1:1]),.I2(un1_df_1),.I3(d_cnst),.I4(d_cnst_sm0),.LO(un86_df));
defparam desc834.INIT=32'h404F4040;
  LUT6_L desc835(.I0(\d_cnst_sn.reg0_28_2526_a5_1_0 ),.I1(\d_cnst_sn.reg1_16_8_1837_2_tz ),.I2(\d_cnst_sn.reg0_28_7_a0_0 [9:9]),.I3(\d_cnst_sn.reg0_28_0 [20:20]),.I4(t_1[20:20]),.I5(\d_cnst_sn.reg0_28_4_2459_0 ),.LO(reg0_28_4_2459));
defparam desc835.INIT=64'hFFFFFFFF0E00EE00;
  LUT5_L desc836(.I0(\d_cnst_sn.reg0_28_7_a0_0 [9:9]),.I1(\d_cnst_sn.reg0_28_11_2228_a6_1_1 ),.I2(\d_cnst_sn.reg1_16_8_1837_3_1 ),.I3(t_1[27:27]),.I4(\d_cnst_sn.reg1_16_8_1837_0 ),.LO(reg1_16_8_1837));
defparam desc836.INIT=32'hFFFF54FC;
  LUT5_L desc837(.I0(\d_cnst_sn.reg0_28_7_a0_0 [9:9]),.I1(\d_cnst_sn.reg0_28_7_2360_3_1 ),.I2(\d_cnst_sn.reg0_28_7_2360_a6_1_1 ),.I3(t_1[23:23]),.I4(\d_cnst_sn.reg0_28_7_2360_0 ),.LO(reg0_28_7_2360));
defparam desc837.INIT=32'hFFFF54FC;
  LUT5_L desc838(.I0(\d_cnst_sn.reg0_28_7_a0_0 [9:9]),.I1(\d_cnst_sn.reg0_28_10_2261_a6_1_1 ),.I2(\d_cnst_sn.reg1_16_7_1870_3_1 ),.I3(t_1[26:26]),.I4(\d_cnst_sn.reg1_16_7_1870_0 ),.LO(reg1_16_7_1870));
defparam desc838.INIT=32'hFFFF54FC;
  LUT5_L desc839(.I0(\d_cnst_sn.reg0_28_7_a0_0 [9:9]),.I1(\d_cnst_sn.reg0_28_5_2426_3_1 ),.I2(\d_cnst_sn.reg0_28_5_2426_a6_1_1 ),.I3(t_1[21:21]),.I4(\d_cnst_sn.reg0_28_5_2426_0 ),.LO(reg0_28_5_2426));
defparam desc839.INIT=32'hFFFF54FC;
  LUT6_L desc840(.I0(\d_cnst_sn.reg0_28_2526_a5_1_0 ),.I1(\d_cnst_sn.reg1_16_8_1837_2_tz ),.I2(\d_cnst_sn.reg0_28_7_a0_0 [9:9]),.I3(\d_cnst_sn.reg0_28_0 [19:19]),.I4(t_1[19:19]),.I5(\d_cnst_sn.reg0_28_3_2492_1 ),.LO(reg0_28_3_2492));
defparam desc840.INIT=64'hFFFFFFFF0E00EE00;
  LUT5_L desc841(.I0(\d_cnst_sn.reg0_28_7_a0_0 [9:9]),.I1(\d_cnst_sn.reg0_28_6_2393_3_1 ),.I2(\d_cnst_sn.reg0_28_6_2393_a6_1_1 ),.I3(t_1[22:22]),.I4(\d_cnst_sn.reg0_28_6_2393_0 ),.LO(reg0_28_6_2393));
defparam desc841.INIT=32'hFFFF54FC;
  LUT5_L desc842(.I0(\d_cnst_sn.reg0_28_7_a0_0 [9:9]),.I1(\d_cnst_sn.reg0_28_9_2294_3_1 ),.I2(\d_cnst_sn.reg0_28_9_2294_a6_1_1 ),.I3(t_1[25:25]),.I4(\d_cnst_sn.reg0_28_9_2294_0 ),.LO(N_3673));
defparam desc842.INIT=32'hFFFF54FC;
  LUT6_L desc843(.I0(\d_cnst_sn.reg1_16_8_1837_2_tz ),.I1(\d_cnst_sn.reg0_28_7_a0_0 [9:9]),.I2(reg0_28_7_d[24:24]),.I3(\d_cnst_sn.reg0_28_8_2327_a6_1_1 ),.I4(t_1[24:24]),.I5(\d_cnst_sn.reg0_28_8_2327_0 ),.LO(reg0_28_8_2327));
defparam desc843.INIT=64'hFFFFFFFF3320FFA8;
  LUT6_L desc844(.I0(\d_cnst_sn.reg0_m9_i_a0_0 ),.I1(N_514_i),.I2(N_527_i),.I3(t_1[29:29]),.I4(reg2_16_11_a3[29:29]),.I5(\d_cnst_sn.reg2_16_1 [29:29]),.LO(reg2_16[29:29]));
defparam desc844.INIT=64'hFFFFFFFFFFFF0008;
  LUT6_L desc845(.I0(\d_cnst_sn.b64_0 ),.I1(\d_cnst_sn.b60_0 ),.I2(\d_cnst_sn.reg1_16_a0_1 [3:3]),.I3(\d_cnst_sn.reg0_1 [7:7]),.I4(t_1[7:7]),.I5(N_1042),.LO(reg0_28[7:7]));
defparam desc845.INIT=64'h0F00FF0001001100;
  LUT6_L desc846(.I0(\d_cnst_sn.b60_0 ),.I1(\d_cnst_sn.reg1_16_a0_1 [3:3]),.I2(\d_cnst_sn.reg2_16_1 [25:25]),.I3(t_1[25:25]),.I4(reg2_16_11_a4[25:25]),.I5(N_1584),.LO(reg2_16[25:25]));
defparam desc846.INIT=64'h000030F000001050;
  LUT6_L desc847(.I0(\d_cnst_sn.b60_0 ),.I1(\d_cnst_sn.reg1_16_a0_1 [3:3]),.I2(\d_cnst_sn.reg2_16_1 [24:24]),.I3(t_1[24:24]),.I4(reg2_16_11_a4[24:24]),.I5(N_1583),.LO(reg2_16[24:24]));
defparam desc847.INIT=64'h000030F000001050;
  LUT6_L desc848(.I0(\d_cnst_sn.b60_0 ),.I1(\d_cnst_sn.reg1_16_a0_1 [3:3]),.I2(\d_cnst_sn.reg2_16_1 [23:23]),.I3(t_1[23:23]),.I4(reg2_16_11_a4[23:23]),.I5(N_1582),.LO(reg2_16[23:23]));
defparam desc848.INIT=64'h000030F000001050;
  LUT6_L desc849(.I0(\d_cnst_sn.b60_0 ),.I1(\d_cnst_sn.reg1_16_a0_1 [3:3]),.I2(\d_cnst_sn.reg2_16_1 [22:22]),.I3(t_1[22:22]),.I4(reg2_16_11_a4[22:22]),.I5(N_1581),.LO(reg2_16[22:22]));
defparam desc849.INIT=64'h000030F000001050;
  LUT6_L desc850(.I0(\d_cnst_sn.b60_0 ),.I1(\d_cnst_sn.reg1_16_a0_1 [3:3]),.I2(\d_cnst_sn.reg2_16_1 [21:21]),.I3(t_1[21:21]),.I4(reg2_16_11_a4[21:21]),.I5(N_1580),.LO(reg2_16[21:21]));
defparam desc850.INIT=64'h000030F000001050;
  LUT6_L b_e(.I0(b),.I1(state),.I2(N_7_i),.I3(N_514_i),.I4(b_2_sqmuxa),.I5(N_3912),.LO(b_0));
defparam b_e.INIT=64'hA222AA2AE2E2EAEA;
  LUT6 desc851(.I0(d[0:0]),.I1(d[1:1]),.I2(un1_df_1),.I3(d_cnst),.I4(d_cnst_sm0),.I5(un36_df),.O(un1_df_17_2));
defparam desc851.INIT=64'h000000008F808080;
  LUT6_L desc852(.I0(inf_abs0_2[4:4]),.I1(inf_abs0_2[27:27]),.I2(inf_abs0_2[28:28]),.I3(un1_inf_abs0_10[4:4]),.I4(un1_inf_abs0_11[4:4]),.I5(addr_4_sqmuxa_1_1),.LO(N_54));
defparam desc852.INIT=64'hFFFFFFFF04C435F5;
  LUT6_L desc853(.I0(inf_abs0_2[2:2]),.I1(inf_abs0_2[27:27]),.I2(inf_abs0_2[28:28]),.I3(un1_inf_abs0_10[2:2]),.I4(un1_inf_abs0_11[2:2]),.I5(addr_4_sqmuxa_1_1),.LO(N_45));
defparam desc853.INIT=64'hFFFFFFFF04C435F5;
  LUT6 desc854(.I0(d[0:0]),.I1(d[1:1]),.I2(un1_df_1),.I3(N_3910),.I4(d_cnst),.I5(d_cnst_sm0),.O(N_1132));
defparam desc854.INIT=64'h1000100010001F00;
  LUT6 desc855(.I0(d[0:0]),.I1(d[1:1]),.I2(un1_df_1),.I3(N_3910),.I4(d_cnst),.I5(d_cnst_sm0),.O(N_1270));
defparam desc855.INIT=64'h200020002F002000;
  LUT6_L desc856(.I0(\d_cnst_sn.reg0_28_9_2294_a6_3_0 ),.I1(m_2[28:28]),.I2(\d_cnst_sn.reg0_28_7_a0_0 [9:9]),.I3(\d_cnst_sn.reg1_16_9_1804_3_tz ),.I4(t_1[28:28]),.I5(N_3614),.LO(reg1_16_9));
defparam desc856.INIT=64'hFFFFFFFF8F88FF88;
  LUT6 desc857(.I0(N_7_i),.I1(N_1901),.I2(N_513_i),.I3(N_514_i),.I4(un36_df),.I5(un87_df),.O(reg3_1_sqmuxa));
defparam desc857.INIT=64'h0000000100000000;
  LUT6 desc858(.I0(N_7_i),.I1(N_1901),.I2(N_513_i),.I3(N_514_i),.I4(un36_df),.I5(un87_df),.O(reg3_14_sqmuxa));
defparam desc858.INIT=64'h0000100000000000;
  LUT6 desc859(.I0(d[0:0]),.I1(d[1:1]),.I2(un1_df_1),.I3(d_cnst),.I4(d_cnst_sm0),.I5(\d_cnst_sn.un1_state_3_1 ),.O(un1_state_3_i));
defparam desc859.INIT=64'h0000000020202F20;
  LUT6 desc860(.I0(d[0:0]),.I1(d[1:1]),.I2(un1_df_1),.I3(d_cnst),.I4(d_cnst_sm0),.I5(\d_cnst_sn.un1_state_3_1 ),.O(un1_state_4_i));
defparam desc860.INIT=64'h000000001010101F;
  LUT5_L desc861(.I0(m_2[15:15]),.I1(N_3916),.I2(N_1132),.I3(N_1050),.I4(N_1082),.LO(reg0_28[15:15]));
defparam desc861.INIT=32'hAFA3ACA0;
  LUT5_L desc862(.I0(m_2[15:15]),.I1(N_3916),.I2(N_1270),.I3(N_1050),.I4(N_1082),.LO(reg1_16[15:15]));
defparam desc862.INIT=32'hAFA3ACA0;
  LUT5_L desc863(.I0(m_2[1:1]),.I1(N_3916),.I2(N_1132),.I3(N_1036),.I4(N_1068),.LO(reg0_28[1:1]));
defparam desc863.INIT=32'hAFA3ACA0;
  LUT5_L desc864(.I0(m_2[16:16]),.I1(N_3916),.I2(N_1132),.I3(N_1051),.I4(N_1083),.LO(reg0_28[16:16]));
defparam desc864.INIT=32'hAFA3ACA0;
  LUT5_L desc865(.I0(m_2[18:18]),.I1(N_3916),.I2(N_1132),.I3(N_1053),.I4(N_1085),.LO(reg0_28[18:18]));
defparam desc865.INIT=32'hAFA3ACA0;
  LUT5_L desc866(.I0(m_2[1:1]),.I1(N_3916),.I2(N_1270),.I3(N_1036),.I4(N_1068),.LO(reg1_16[1:1]));
defparam desc866.INIT=32'hAFA3ACA0;
  LUT5_L desc867(.I0(m_2[16:16]),.I1(N_3916),.I2(N_1270),.I3(N_1051),.I4(N_1083),.LO(reg1_16[16:16]));
defparam desc867.INIT=32'hAFA3ACA0;
  LUT5_L desc868(.I0(m_2[13:13]),.I1(N_3916),.I2(N_1132),.I3(N_1048),.I4(N_1080),.LO(reg0_28[13:13]));
defparam desc868.INIT=32'hAFA3ACA0;
  LUT5_L desc869(.I0(m_2[13:13]),.I1(N_3916),.I2(N_1270),.I3(N_1048),.I4(N_1080),.LO(reg1_16[13:13]));
defparam desc869.INIT=32'hAFA3ACA0;
  LUT5_L desc870(.I0(m_2[9:9]),.I1(N_3916),.I2(N_1132),.I3(N_1044),.I4(N_1076),.LO(reg0_28[9:9]));
defparam desc870.INIT=32'hAFA3ACA0;
  LUT5_L desc871(.I0(m_2[10:10]),.I1(N_3916),.I2(N_1132),.I3(N_1045),.I4(N_1077),.LO(reg0_28[10:10]));
defparam desc871.INIT=32'hAFA3ACA0;
  LUT5_L desc872(.I0(m_2[11:11]),.I1(N_3916),.I2(N_1132),.I3(N_1046),.I4(N_1078),.LO(reg0_28[11:11]));
defparam desc872.INIT=32'hAFA3ACA0;
  LUT5_L desc873(.I0(m_2[12:12]),.I1(N_3916),.I2(N_1132),.I3(N_1047),.I4(N_1079),.LO(reg0_28[12:12]));
defparam desc873.INIT=32'hAFA3ACA0;
  LUT5_L desc874(.I0(m_2[14:14]),.I1(N_3916),.I2(N_1132),.I3(N_1049),.I4(N_1081),.LO(reg0_28[14:14]));
defparam desc874.INIT=32'hAFA3ACA0;
  LUT5_L desc875(.I0(m_2[2:2]),.I1(N_3916),.I2(N_1270),.I3(N_1037),.I4(N_1069),.LO(reg1_16[2:2]));
defparam desc875.INIT=32'hAFA3ACA0;
  LUT5_L desc876(.I0(m_2[9:9]),.I1(N_3916),.I2(N_1270),.I3(N_1044),.I4(N_1076),.LO(reg1_16[9:9]));
defparam desc876.INIT=32'hAFA3ACA0;
  LUT5_L desc877(.I0(m_2[10:10]),.I1(N_3916),.I2(N_1270),.I3(N_1045),.I4(N_1077),.LO(reg1_16[10:10]));
defparam desc877.INIT=32'hAFA3ACA0;
  LUT5_L desc878(.I0(m_2[11:11]),.I1(N_3916),.I2(N_1270),.I3(N_1046),.I4(N_1078),.LO(reg1_16[11:11]));
defparam desc878.INIT=32'hAFA3ACA0;
  LUT5_L desc879(.I0(m_2[12:12]),.I1(N_3916),.I2(N_1270),.I3(N_1047),.I4(N_1079),.LO(reg1_16[12:12]));
defparam desc879.INIT=32'hAFA3ACA0;
  LUT5_L desc880(.I0(m_2[14:14]),.I1(N_3916),.I2(N_1270),.I3(N_1049),.I4(N_1081),.LO(reg1_16[14:14]));
defparam desc880.INIT=32'hAFA3ACA0;
  LUT5_L desc881(.I0(m_2[17:17]),.I1(N_3916),.I2(N_1270),.I3(N_1052),.I4(N_1084),.LO(reg1_16[17:17]));
defparam desc881.INIT=32'hAFA3ACA0;
  LUT6 desc882(.I0(N_7_i),.I1(N_1901),.I2(N_513_i),.I3(N_514_i),.I4(un1_df_17_2),.I5(rd_4_sqmuxa),.O(reg3_17_sn_N_5));
defparam desc882.INIT=64'h00000000EFFFFFFF;
  LUT6 desc883(.I0(state),.I1(N_7_i),.I2(N_1892),.I3(un36_df),.I4(N_1890),.I5(un86_df),.O(un1_state_1_0_i));
defparam desc883.INIT=64'h0002000200000002;
  LUT3 desc884(.I0(reg3[1:1]),.I1(reg3_1_1[1:1]),.I2(reg3_1_sqmuxa),.O(N_1689));
defparam desc884.INIT=8'hCA;
  LUT3 desc885(.I0(reg3[2:2]),.I1(reg3_1_1[2:2]),.I2(reg3_1_sqmuxa),.O(N_1690));
defparam desc885.INIT=8'hCA;
  LUT3 desc886(.I0(reg3[0:0]),.I1(m_2[0:0]),.I2(reg3_1_sqmuxa),.O(N_1688));
defparam desc886.INIT=8'hCA;
  LUT6 desc887(.I0(N_513_i),.I1(m_2[18:18]),.I2(N_3916),.I3(reg0_28_7_a1[18:18]),.I4(N_1270),.I5(reg3_1_1[18:18]),.O(\d_cnst_sn.reg1_0 [18:18]));
defparam desc887.INIT=64'hCCCCF0FFCCCCF0FA;
  LUT6 desc888(.I0(N_513_i),.I1(m_2[17:17]),.I2(N_3916),.I3(reg0_28_7_a1[17:17]),.I4(N_1132),.I5(reg3_1_1[17:17]),.O(\d_cnst_sn.reg0_0 [17:17]));
defparam desc888.INIT=64'hCCCCF0FFCCCCF0FA;
  LUT6 desc889(.I0(\d_cnst_sn.reg1_16_a2_0 [5:5]),.I1(m_2[8:8]),.I2(\d_cnst_sn.reg0_28_a1_1 [4:4]),.I3(r_4[7:7]),.I4(reg3_1_1[8:8]),.I5(N_1132),.O(\d_cnst_sn.reg0_1 [8:8]));
defparam desc889.INIT=64'hCCCCCCCCFF0F5505;
  LUT6 desc890(.I0(\d_cnst_sn.reg1_16_a2_0 [5:5]),.I1(m_2[8:8]),.I2(\d_cnst_sn.reg0_28_a1_1 [4:4]),.I3(r_4[7:7]),.I4(reg3_1_1[8:8]),.I5(N_1270),.O(\d_cnst_sn.reg1_1 [8:8]));
defparam desc890.INIT=64'hCCCCCCCCFF0F5505;
  LUT6 desc891(.I0(\d_cnst_sn.reg1_16_a2_0 [5:5]),.I1(m_2[6:6]),.I2(\d_cnst_sn.reg0_28_a1_1 [4:4]),.I3(r_4[5:5]),.I4(reg3_1_1[6:6]),.I5(N_1132),.O(\d_cnst_sn.reg0_1 [6:6]));
defparam desc891.INIT=64'hCCCCCCCCFF0F5505;
  LUT6 desc892(.I0(\d_cnst_sn.reg1_16_a2_0 [5:5]),.I1(m_2[6:6]),.I2(\d_cnst_sn.reg0_28_a1_1 [4:4]),.I3(r_4[5:5]),.I4(reg3_1_1[6:6]),.I5(N_1270),.O(\d_cnst_sn.reg1_1 [6:6]));
defparam desc892.INIT=64'hCCCCCCCCFF0F5505;
  LUT6 desc893(.I0(\d_cnst_sn.reg1_16_a2_0 [5:5]),.I1(m_2[5:5]),.I2(\d_cnst_sn.reg0_28_a1_1 [4:4]),.I3(r_4[4:4]),.I4(reg3_1_1[5:5]),.I5(N_1132),.O(\d_cnst_sn.reg0_1 [5:5]));
defparam desc893.INIT=64'hCCCCCCCCFF0F5505;
  LUT6 desc894(.I0(\d_cnst_sn.reg1_16_a2_0 [5:5]),.I1(m_2[5:5]),.I2(\d_cnst_sn.reg0_28_a1_1 [4:4]),.I3(r_4[4:4]),.I4(reg3_1_1[5:5]),.I5(N_1270),.O(\d_cnst_sn.reg1_1 [5:5]));
defparam desc894.INIT=64'hCCCCCCCCFF0F5505;
  LUT6 desc895(.I0(\d_cnst_sn.reg1_16_a2_0 [5:5]),.I1(m_2[4:4]),.I2(\d_cnst_sn.reg0_28_a1_1 [4:4]),.I3(r_4[3:3]),.I4(reg3_1_1[4:4]),.I5(N_1270),.O(\d_cnst_sn.reg1_1 [4:4]));
defparam desc895.INIT=64'hCCCCCCCCFF0F5505;
  LUT6 desc896(.I0(\d_cnst_sn.reg1_16_a2_0 [5:5]),.I1(m_2[4:4]),.I2(\d_cnst_sn.reg0_28_a1_1 [4:4]),.I3(r_4[3:3]),.I4(reg3_1_1[4:4]),.I5(N_1132),.O(\d_cnst_sn.reg0_1 [4:4]));
defparam desc896.INIT=64'hCCCCCCCCFF0F5505;
  LUT6 desc897(.I0(\d_cnst_sn.reg1_16_a2_0 [5:5]),.I1(m_2[3:3]),.I2(\d_cnst_sn.reg0_28_a1_1 [4:4]),.I3(reg3_1_1[3:3]),.I4(N_28),.I5(N_1270),.O(\d_cnst_sn.reg1_1 [3:3]));
defparam desc897.INIT=64'hCCCCCCCCFF550F05;
  LUT6 desc898(.I0(\d_cnst_sn.reg1_16_a2_0 [5:5]),.I1(m_2[3:3]),.I2(\d_cnst_sn.reg0_28_a1_1 [4:4]),.I3(reg3_1_1[3:3]),.I4(N_28),.I5(N_1132),.O(\d_cnst_sn.reg0_1 [3:3]));
defparam desc898.INIT=64'hCCCCCCCCFF550F05;
  LUT6 desc899(.I0(\d_cnst_sn.reg1_16_a2_0 [5:5]),.I1(m_2[2:2]),.I2(\d_cnst_sn.reg0_28_a1_1 [4:4]),.I3(reg3_1_1[2:2]),.I4(r_4[1:1]),.I5(N_1132),.O(\d_cnst_sn.reg0_1 [2:2]));
defparam desc899.INIT=64'hCCCCCCCCFF550F05;
  LUT6_L desc900(.I0(reg3[4:4]),.I1(state),.I2(inf_abs0_2[31:31]),.I3(N_2240_i),.I4(addr_4_sqmuxa_1_1),.I5(N_54),.LO(N_56_i));
defparam desc900.INIT=64'hEE22E222EEEEEEEE;
  LUT6_L desc901(.I0(reg3[2:2]),.I1(state),.I2(inf_abs0_2[31:31]),.I3(N_2240_i),.I4(addr_4_sqmuxa_1_1),.I5(N_45),.LO(N_47_i));
defparam desc901.INIT=64'hEE22E222EEEEEEEE;
  LUT5 desc902(.I0(reg3[3:3]),.I1(inf_abs0_2[3:3]),.I2(reg3_1_1[3:3]),.I3(rd_4_sqmuxa),.I4(reg3_1_sqmuxa),.O(reg3_N_7_i_RNO));
defparam desc902.INIT=32'h330F33AA;
  LUT5 desc903(.I0(un3_reg3_s_1),.I1(inf_abs0_2[4:4]),.I2(reg3_1_1[4:4]),.I3(rd_4_sqmuxa),.I4(reg3_1_sqmuxa),.O(reg3_1_sqmuxa_RNIEMUH1));
defparam desc903.INIT=32'h330F3355;
  LUT5 desc904(.I0(un3_reg3_s_2),.I1(inf_abs0_2[5:5]),.I2(reg3_1_1[5:5]),.I3(rd_4_sqmuxa),.I4(reg3_1_sqmuxa),.O(reg3_1_sqmuxa_RNIHMUH1));
defparam desc904.INIT=32'h330F3355;
  LUT5 desc905(.I0(un3_reg3_s_4),.I1(inf_abs0_2[7:7]),.I2(reg3_1_1[7:7]),.I3(rd_4_sqmuxa),.I4(reg3_1_sqmuxa),.O(reg3_1_sqmuxa_RNINMUH1));
defparam desc905.INIT=32'h330F3355;
  LUT5 desc906(.I0(un3_reg3_s_3),.I1(inf_abs0_2[6:6]),.I2(reg3_1_1[6:6]),.I3(rd_4_sqmuxa),.I4(reg3_1_sqmuxa),.O(reg3_1_sqmuxa_RNIKMUH1));
defparam desc906.INIT=32'h330F3355;
  LUT5 desc907(.I0(un3_reg3_s_6),.I1(inf_abs0_2[9:9]),.I2(reg3_1_1[9:9]),.I3(rd_4_sqmuxa),.I4(reg3_1_sqmuxa),.O(reg3_1_sqmuxa_RNITMUH1));
defparam desc907.INIT=32'h330F3355;
  LUT5 desc908(.I0(un3_reg3_s_5),.I1(inf_abs0_2[8:8]),.I2(reg3_1_1[8:8]),.I3(rd_4_sqmuxa),.I4(reg3_1_sqmuxa),.O(reg3_1_sqmuxa_RNIQMUH1));
defparam desc908.INIT=32'h330F3355;
  LUT5 desc909(.I0(un3_reg3_s_7),.I1(inf_abs0_2[10:10]),.I2(reg3_1_1[10:10]),.I3(rd_4_sqmuxa),.I4(reg3_1_sqmuxa),.O(reg3_1_sqmuxa_RNIE1DM1));
defparam desc909.INIT=32'h330F3355;
  LUT5 desc910(.I0(un3_reg3_s_8),.I1(inf_abs0_2[11:11]),.I2(reg3_1_1[11:11]),.I3(rd_4_sqmuxa),.I4(reg3_1_sqmuxa),.O(reg3_1_sqmuxa_RNIH1DM1));
defparam desc910.INIT=32'h330F3355;
  LUT5_L desc911(.I0(un1_df_16),.I1(N_1810),.I2(un11_reg0_s_1),.I3(un32_reg0_s_1),.I4(N_1658),.LO(N_1813));
defparam desc911.INIT=32'hFEDC3210;
  LUT5_L desc912(.I0(un1_df_16),.I1(N_1810),.I2(N_1684),.I3(un32_reg0_s_27),.I4(un11_reg0_s_27),.LO(N_1839));
defparam desc912.INIT=32'hF3D1E2C0;
  LUT5_L desc913(.I0(un1_df_16),.I1(N_1810),.I2(N_1685),.I3(un32_reg0_s_28),.I4(un11_reg0_s_28),.LO(N_1840));
defparam desc913.INIT=32'hF3D1E2C0;
  LUT5_L desc914(.I0(un1_df_16),.I1(N_1810),.I2(N_1673),.I3(un32_reg0_s_16),.I4(un11_reg0_s_16),.LO(N_1828));
defparam desc914.INIT=32'hF3D1E2C0;
  LUT5 desc915(.I0(un1_df_16),.I1(N_1810),.I2(N_1666),.I3(un32_reg0_s_9),.I4(un11_reg0_s_9),.O(N_1821));
defparam desc915.INIT=32'hF3D1E2C0;
  LUT5_L desc916(.I0(un1_df_16),.I1(N_1810),.I2(N_1676),.I3(un32_reg0_s_19),.I4(un11_reg0_s_19),.LO(N_1831));
defparam desc916.INIT=32'hF3D1E2C0;
  LUT5_L desc917(.I0(un1_df_16),.I1(N_1810),.I2(N_1677),.I3(un32_reg0_s_20),.I4(un11_reg0_s_20),.LO(N_1832));
defparam desc917.INIT=32'hF3D1E2C0;
  LUT5_L desc918(.I0(un1_df_16),.I1(N_1810),.I2(N_1671),.I3(un32_reg0_s_14),.I4(un11_reg0_s_14),.LO(N_1826));
defparam desc918.INIT=32'hF3D1E2C0;
  LUT5_L desc919(.I0(un1_df_16),.I1(N_1810),.I2(N_1675),.I3(un32_reg0_s_18),.I4(un11_reg0_s_18),.LO(N_1830));
defparam desc919.INIT=32'hF3D1E2C0;
  LUT5 desc920(.I0(un1_df_16),.I1(N_1810),.I2(N_1662),.I3(un32_reg0_s_5),.I4(un11_reg0_s_5),.O(N_1817));
defparam desc920.INIT=32'hF3D1E2C0;
  LUT5_L desc921(.I0(un1_df_16),.I1(N_1810),.I2(N_1669),.I3(un32_reg0_s_12),.I4(un11_reg0_s_12),.LO(N_1824));
defparam desc921.INIT=32'hF3D1E2C0;
  LUT5_L desc922(.I0(un1_df_16),.I1(N_1810),.I2(N_1674),.I3(un32_reg0_s_17),.I4(un11_reg0_s_17),.LO(N_1829));
defparam desc922.INIT=32'hF3D1E2C0;
  LUT5 desc923(.I0(un1_df_16),.I1(N_1810),.I2(N_1667),.I3(un32_reg0_s_10),.I4(un11_reg0_s_10),.O(N_1822));
defparam desc923.INIT=32'hF3D1E2C0;
  LUT5 desc924(.I0(un1_df_16),.I1(N_1810),.I2(N_1668),.I3(un32_reg0_s_11),.I4(un11_reg0_s_11),.O(N_1823));
defparam desc924.INIT=32'hF3D1E2C0;
  LUT5_L desc925(.I0(un1_df_16),.I1(N_1810),.I2(un11_reg0_s_2),.I3(un32_reg0_s_2),.I4(N_1659),.LO(N_1814));
defparam desc925.INIT=32'hFEDC3210;
  LUT5 desc926(.I0(un1_df_16),.I1(N_1810),.I2(N_1663),.I3(un32_reg0_s_6),.I4(un11_reg0_s_6),.O(N_1818));
defparam desc926.INIT=32'hF3D1E2C0;
  LUT5 desc927(.I0(un1_df_16),.I1(N_1810),.I2(N_1665),.I3(un32_reg0_s_8),.I4(un11_reg0_s_8),.O(N_1820));
defparam desc927.INIT=32'hF3D1E2C0;
  LUT5 desc928(.I0(un1_df_16),.I1(N_1810),.I2(un32_reg0_s_3),.I3(un11_reg0_s_3),.I4(N_1660),.O(N_1815));
defparam desc928.INIT=32'hFDEC3120;
  LUT5_L desc929(.I0(un1_df_16),.I1(N_1810),.I2(N_1672),.I3(un32_reg0_s_15),.I4(un11_reg0_s_15),.LO(N_1827));
defparam desc929.INIT=32'hF3D1E2C0;
  LUT5_L desc930(.I0(un1_df_16),.I1(N_1810),.I2(N_1683),.I3(un32_reg0_s_26),.I4(un11_reg0_s_26),.LO(N_1838));
defparam desc930.INIT=32'hF3D1E2C0;
  LUT5_L desc931(.I0(un1_df_16),.I1(N_1810),.I2(N_1682),.I3(un32_reg0_s_25),.I4(un11_reg0_s_25),.LO(N_1837));
defparam desc931.INIT=32'hF3D1E2C0;
  LUT5 desc932(.I0(un1_df_16),.I1(N_1810),.I2(N_1664),.I3(un32_reg0_s_7),.I4(un11_reg0_s_7),.O(N_1819));
defparam desc932.INIT=32'hF3D1E2C0;
  LUT5 desc933(.I0(un1_df_16),.I1(N_1810),.I2(N_1661),.I3(un32_reg0_s_4),.I4(un11_reg0_s_4),.O(N_1816));
defparam desc933.INIT=32'hF3D1E2C0;
  LUT6 desc934(.I0(un3_reg3_s_25),.I1(\d_cnst_sn.reg3_17_4_a2_0 [28:28]),.I2(rd_4_sqmuxa),.I3(reg3_1_1[28:28]),.I4(reg3_1_sqmuxa),.I5(reg3_14_sqmuxa),.O(\d_cnst_sn.reg3_17_6_0 [28:28]));
defparam desc934.INIT=64'hCCCCCCCC0F000A0A;
  LUT6 desc935(.I0(un3_reg3_s_24),.I1(\d_cnst_sn.reg3_17_4_a2_0 [27:27]),.I2(rd_4_sqmuxa),.I3(reg3_1_1[27:27]),.I4(reg3_1_sqmuxa),.I5(reg3_14_sqmuxa),.O(\d_cnst_sn.reg3_17_6_0 [27:27]));
defparam desc935.INIT=64'hCCCCCCCC0F000A0A;
  LUT6 desc936(.I0(un3_reg3_s_15),.I1(reg3_1_1[18:18]),.I2(rd_4_sqmuxa),.I3(reg3_1_sqmuxa),.I4(reg3_14_sqmuxa),.I5(\d_cnst_sn.reg3_17_6_0 [18:18]),.O(\d_cnst_sn.reg3_17_6_1 [18:18]));
defparam desc936.INIT=64'hFFFFFCFA00000000;
  LUT6 desc937(.I0(un3_reg3_s_16),.I1(reg3_1_1[19:19]),.I2(rd_4_sqmuxa),.I3(reg3_1_sqmuxa),.I4(reg3_14_sqmuxa),.I5(\d_cnst_sn.reg3_17_6_0 [19:19]),.O(\d_cnst_sn.reg3_17_6_1 [19:19]));
defparam desc937.INIT=64'hFFFFFCFA00000000;
  LUT6 desc938(.I0(un3_reg3_s_23),.I1(\d_cnst_sn.reg3_17_4_a2_0 [26:26]),.I2(rd_4_sqmuxa),.I3(reg3_1_1[26:26]),.I4(reg3_1_sqmuxa),.I5(reg3_14_sqmuxa),.O(\d_cnst_sn.reg3_17_6_0 [26:26]));
defparam desc938.INIT=64'hCCCCCCCC0F000A0A;
  LUT6 desc939(.I0(un3_reg3_s_14),.I1(reg3_1_1[17:17]),.I2(rd_4_sqmuxa),.I3(reg3_1_sqmuxa),.I4(reg3_14_sqmuxa),.I5(\d_cnst_sn.reg3_17_6_0 [17:17]),.O(\d_cnst_sn.reg3_17_6_1 [17:17]));
defparam desc939.INIT=64'hFFFFFCFA00000000;
  LUT6 desc940(.I0(un3_reg3_s_22),.I1(\d_cnst_sn.reg3_17_4_a2_0 [25:25]),.I2(rd_4_sqmuxa),.I3(reg3_1_1[25:25]),.I4(reg3_1_sqmuxa),.I5(reg3_14_sqmuxa),.O(\d_cnst_sn.reg3_17_6_0 [25:25]));
defparam desc940.INIT=64'hCCCCCCCC0F000A0A;
  LUT6 desc941(.I0(un3_reg3_s_13),.I1(reg3_1_1[16:16]),.I2(rd_4_sqmuxa),.I3(reg3_1_sqmuxa),.I4(reg3_14_sqmuxa),.I5(\d_cnst_sn.reg3_17_6_0 [16:16]),.O(\d_cnst_sn.reg3_17_6_1 [16:16]));
defparam desc941.INIT=64'hFFFFFCFA00000000;
  LUT6 desc942(.I0(un3_reg3_s_12),.I1(reg3_1_1[15:15]),.I2(rd_4_sqmuxa),.I3(reg3_1_sqmuxa),.I4(reg3_14_sqmuxa),.I5(\d_cnst_sn.reg3_17_6_0 [15:15]),.O(\d_cnst_sn.reg3_17_6_1 [15:15]));
defparam desc942.INIT=64'hFFFFFCFA00000000;
  LUT6 desc943(.I0(un3_reg3_s_11),.I1(reg3_1_1[14:14]),.I2(rd_4_sqmuxa),.I3(reg3_1_sqmuxa),.I4(reg3_14_sqmuxa),.I5(\d_cnst_sn.reg3_17_6_0 [14:14]),.O(\d_cnst_sn.reg3_17_6_1 [14:14]));
defparam desc943.INIT=64'hFFFFFCFA00000000;
  LUT6 desc944(.I0(un3_reg3_s_10),.I1(reg3_1_1[13:13]),.I2(rd_4_sqmuxa),.I3(reg3_1_sqmuxa),.I4(reg3_14_sqmuxa),.I5(\d_cnst_sn.reg3_17_6_0 [13:13]),.O(\d_cnst_sn.reg3_17_6_1 [13:13]));
defparam desc944.INIT=64'hFFFFFCFA00000000;
  LUT6 desc945(.I0(un3_reg3_s_17),.I1(\d_cnst_sn.reg3_17_4_a2_0 [20:20]),.I2(reg3_1_1[20:20]),.I3(rd_4_sqmuxa),.I4(reg3_1_sqmuxa),.I5(reg3_14_sqmuxa),.O(\d_cnst_sn.reg3_17_6_0 [20:20]));
defparam desc945.INIT=64'hCCCCCCCC00F000AA;
  LUT6 desc946(.I0(un3_reg3_s_9),.I1(reg3_1_1[12:12]),.I2(rd_4_sqmuxa),.I3(reg3_1_sqmuxa),.I4(reg3_14_sqmuxa),.I5(\d_cnst_sn.reg3_17_6_0 [12:12]),.O(\d_cnst_sn.reg3_17_6_1 [12:12]));
defparam desc946.INIT=64'hFFFFFCFA00000000;
  LUT6 desc947(.I0(un3_reg3_s_21),.I1(reg3_1_1[24:24]),.I2(N_1810),.I3(\d_cnst_sn.reg3_17_sn_m7_0 ),.I4(reg3_1_sqmuxa),.I5(reg3_17_sn_N_5),.O(reg3_17_a0[24:24]));
defparam desc947.INIT=64'hC000A00000000000;
  LUT6 desc948(.I0(un3_reg3_s_20),.I1(reg3_1_1[23:23]),.I2(N_1810),.I3(\d_cnst_sn.reg3_17_sn_m7_0 ),.I4(reg3_1_sqmuxa),.I5(reg3_17_sn_N_5),.O(reg3_17_a0[23:23]));
defparam desc948.INIT=64'hC000A00000000000;
  LUT6 desc949(.I0(un3_reg3_s_19),.I1(reg3_1_1[22:22]),.I2(N_1810),.I3(\d_cnst_sn.reg3_17_sn_m7_0 ),.I4(reg3_1_sqmuxa),.I5(reg3_17_sn_N_5),.O(reg3_17_a0[22:22]));
defparam desc949.INIT=64'hC000A00000000000;
  LUT6 desc950(.I0(un3_reg3_s_18),.I1(reg3_1_1[21:21]),.I2(N_1810),.I3(\d_cnst_sn.reg3_17_sn_m7_0 ),.I4(reg3_1_sqmuxa),.I5(reg3_17_sn_N_5),.O(reg3_17_a0[21:21]));
defparam desc950.INIT=64'hC000A00000000000;
  LUT6_L desc951(.I0(N_1810),.I1(\d_cnst_sn.reg3_17_sn_m7_0 ),.I2(reg3_17_sn_N_5),.I3(N_1689),.I4(N_1751),.I5(N_1813),.LO(reg3_17[1:1]));
defparam desc951.INIT=64'hFF7FF77788088000;
  LUT5_L desc952(.I0(reg3_17_sn_N_5),.I1(N_1690),.I2(N_1841),.I3(N_1752),.I4(N_1814),.LO(reg3_17[2:2]));
defparam desc952.INIT=32'hDF8FD080;
  LUT6_L desc953(.I0(N_1810),.I1(\d_cnst_sn.reg3_17_sn_m7_0 ),.I2(reg3_17_sn_N_5),.I3(N_1812),.I4(N_1688),.I5(N_1750),.LO(reg3_17[0:0]));
defparam desc953.INIT=64'hFF887F08F7807700;
  LUT6_L desc954(.I0(\d_cnst_sn.b64_0 ),.I1(\d_cnst_sn.b60_0 ),.I2(\d_cnst_sn.reg1_16_a0_1 [3:3]),.I3(\d_cnst_sn.reg0_1 [3:3]),.I4(t_1[3:3]),.I5(N_1038),.LO(reg0_28[3:3]));
defparam desc954.INIT=64'h0F00FF0001001100;
  LUT6_L desc955(.I0(\d_cnst_sn.b64_0 ),.I1(\d_cnst_sn.b60_0 ),.I2(\d_cnst_sn.reg1_16_a0_1 [3:3]),.I3(\d_cnst_sn.reg0_1 [2:2]),.I4(t_1[2:2]),.I5(N_1037),.LO(reg0_28[2:2]));
defparam desc955.INIT=64'h0F00FF0001001100;
  LUT6_L desc956(.I0(\d_cnst_sn.b64_0 ),.I1(\d_cnst_sn.b60_0 ),.I2(\d_cnst_sn.reg1_16_a0_1 [3:3]),.I3(\d_cnst_sn.reg1_1 [3:3]),.I4(t_1[3:3]),.I5(N_1038),.LO(reg1_16[3:3]));
defparam desc956.INIT=64'h0F00FF0001001100;
  LUT6_L desc957(.I0(\d_cnst_sn.b64_0 ),.I1(\d_cnst_sn.b60_0 ),.I2(\d_cnst_sn.reg1_16_a0_1 [3:3]),.I3(\d_cnst_sn.reg0_1 [8:8]),.I4(t_1[8:8]),.I5(N_1043),.LO(reg0_28[8:8]));
defparam desc957.INIT=64'h0F00FF0001001100;
  LUT6_L desc958(.I0(\d_cnst_sn.b64_0 ),.I1(\d_cnst_sn.b60_0 ),.I2(\d_cnst_sn.reg1_16_a0_1 [3:3]),.I3(\d_cnst_sn.reg1_1 [8:8]),.I4(t_1[8:8]),.I5(N_1043),.LO(reg1_16[8:8]));
defparam desc958.INIT=64'h0F00FF0001001100;
  LUT6_L desc959(.I0(\d_cnst_sn.b64_0 ),.I1(\d_cnst_sn.b60_0 ),.I2(\d_cnst_sn.reg1_16_a0_1 [3:3]),.I3(\d_cnst_sn.reg1_1 [6:6]),.I4(t_1[6:6]),.I5(N_1041),.LO(reg1_16[6:6]));
defparam desc959.INIT=64'h0F00FF0001001100;
  LUT6_L desc960(.I0(\d_cnst_sn.b64_0 ),.I1(\d_cnst_sn.b60_0 ),.I2(\d_cnst_sn.reg1_16_a0_1 [3:3]),.I3(\d_cnst_sn.reg0_1 [5:5]),.I4(t_1[5:5]),.I5(N_1040),.LO(reg0_28[5:5]));
defparam desc960.INIT=64'h0F00FF0001001100;
  LUT6_L desc961(.I0(\d_cnst_sn.b64_0 ),.I1(\d_cnst_sn.b60_0 ),.I2(\d_cnst_sn.reg1_16_a0_1 [3:3]),.I3(\d_cnst_sn.reg0_1 [6:6]),.I4(t_1[6:6]),.I5(N_1041),.LO(reg0_28[6:6]));
defparam desc961.INIT=64'h0F00FF0001001100;
  LUT6_L desc962(.I0(\d_cnst_sn.b64_0 ),.I1(\d_cnst_sn.b60_0 ),.I2(\d_cnst_sn.reg1_16_a0_1 [3:3]),.I3(\d_cnst_sn.reg1_1 [4:4]),.I4(t_1[4:4]),.I5(N_1039),.LO(reg1_16[4:4]));
defparam desc962.INIT=64'h0F00FF0001001100;
  LUT6_L desc963(.I0(\d_cnst_sn.b64_0 ),.I1(\d_cnst_sn.b60_0 ),.I2(\d_cnst_sn.reg1_16_a0_1 [3:3]),.I3(\d_cnst_sn.reg1_1 [5:5]),.I4(t_1[5:5]),.I5(N_1040),.LO(reg1_16[5:5]));
defparam desc963.INIT=64'h0F00FF0001001100;
  LUT6_L desc964(.I0(\d_cnst_sn.b64_0 ),.I1(\d_cnst_sn.b60_0 ),.I2(\d_cnst_sn.reg1_16_a0_1 [3:3]),.I3(\d_cnst_sn.reg0_1 [4:4]),.I4(t_1[4:4]),.I5(N_1039),.LO(reg0_28[4:4]));
defparam desc964.INIT=64'h0F00FF0001001100;
  LUT6_L desc965(.I0(N_1810),.I1(\d_cnst_sn.reg3_17_sn_m7_0 ),.I2(reg3_14_sqmuxa),.I3(reg3_1_sqmuxa_RNIEMUH1),.I4(N_1816),.I5(r_4_2_a1_lut6_2_RNI2T8R3[3:3]),.LO(reg3_17[4:4]));
defparam desc965.INIT=64'h777F0008F7FF8088;
  LUT6_L desc966(.I0(N_1810),.I1(\d_cnst_sn.reg3_17_sn_m7_0 ),.I2(reg3_14_sqmuxa),.I3(reg3_1_sqmuxa_RNIHMUH1),.I4(N_1817),.I5(r_4_2_a1_lut6_2_RNI5V8R3[3:3]),.LO(reg3_17[5:5]));
defparam desc966.INIT=64'h777F0008F7FF8088;
  LUT6_L desc967(.I0(N_1810),.I1(\d_cnst_sn.reg3_17_sn_m7_0 ),.I2(reg3_14_sqmuxa),.I3(reg3_1_sqmuxa_RNINMUH1),.I4(N_1819),.I5(r_4_1_RNICM731[6:6]),.LO(reg3_17[7:7]));
defparam desc967.INIT=64'h777F0008F7FF8088;
  LUT6_L desc968(.I0(N_1810),.I1(\d_cnst_sn.reg3_17_sn_m7_0 ),.I2(reg3_14_sqmuxa),.I3(reg3_1_sqmuxa_RNIKMUH1),.I4(N_1818),.I5(r_4_1_RNI9K731[5:5]),.LO(reg3_17[6:6]));
defparam desc968.INIT=64'h777F0008F7FF8088;
  LUT6_L desc969(.I0(N_1810),.I1(\d_cnst_sn.reg3_17_sn_m7_0 ),.I2(reg3_14_sqmuxa),.I3(reg3_1_sqmuxa_RNITMUH1),.I4(N_1821),.I5(r_4_1_RNIIQ731[8:8]),.LO(reg3_17[9:9]));
defparam desc969.INIT=64'h777F0008F7FF8088;
  LUT6_L desc970(.I0(N_1810),.I1(\d_cnst_sn.reg3_17_sn_m7_0 ),.I2(reg3_14_sqmuxa),.I3(reg3_1_sqmuxa_RNIQMUH1),.I4(N_1820),.I5(r_4_1_RNIFO731[7:7]),.LO(reg3_17[8:8]));
defparam desc970.INIT=64'h777F0008F7FF8088;
  LUT6_L desc971(.I0(N_1810),.I1(\d_cnst_sn.reg3_17_sn_m7_0 ),.I2(reg3_14_sqmuxa),.I3(reg3_1_sqmuxa_RNIE1DM1),.I4(N_1822),.I5(r_4_1_RNIS3K91[9:9]),.LO(reg3_17[10:10]));
defparam desc971.INIT=64'h777F0008F7FF8088;
  LUT6_L desc972(.I0(N_1810),.I1(\d_cnst_sn.reg3_17_sn_m7_0 ),.I2(reg3_14_sqmuxa),.I3(reg3_1_sqmuxa_RNIH1DM1),.I4(N_1823),.I5(r_4_1_RNIDBOH1[10:10]),.LO(reg3_17[11:11]));
defparam desc972.INIT=64'h777F0008F7FF8088;
  LUT6_L desc973(.I0(N_1810),.I1(\d_cnst_sn.reg3_17_sn_m7_0 ),.I2(N_1670),.I3(\d_cnst_sn.reg3_17_6_1 [13:13]),.I4(N_1732),.I5(reg3_17_4_a2[13:13]),.LO(reg3_17[13:13]));
defparam desc973.INIT=64'h75752020FD75A820;
  LUT6_L desc974(.I0(N_527_i),.I1(reg3_14_sqmuxa),.I2(\d_cnst_sn.reg3_17_6_0 [27:27]),.I3(N_1841),.I4(t_1[27:27]),.I5(N_1839),.LO(reg3_17[27:27]));
defparam desc974.INIT=64'hF0FFF4FFF000F400;
  LUT6_L desc975(.I0(N_527_i),.I1(reg3_14_sqmuxa),.I2(\d_cnst_sn.reg3_17_6_0 [28:28]),.I3(N_1841),.I4(t_1[28:28]),.I5(N_1840),.LO(reg3_17[28:28]));
defparam desc975.INIT=64'hF0FFF4FFF000F400;
  LUT6_L desc976(.I0(N_527_i),.I1(reg3_14_sqmuxa),.I2(N_1841),.I3(\d_cnst_sn.reg3_17_6_1 [16:16]),.I4(t_1[16:16]),.I5(N_1828),.LO(reg3_17[16:16]));
defparam desc976.INIT=64'hBF0FFF0FB000F000;
  LUT6_L desc977(.I0(N_527_i),.I1(reg3_14_sqmuxa),.I2(N_1841),.I3(\d_cnst_sn.reg3_17_6_1 [19:19]),.I4(t_1[19:19]),.I5(N_1831),.LO(reg3_17[19:19]));
defparam desc977.INIT=64'hBF0FFF0FB000F000;
  LUT6_L desc978(.I0(N_527_i),.I1(reg3_14_sqmuxa),.I2(\d_cnst_sn.reg3_17_6_0 [20:20]),.I3(N_1841),.I4(t_1[20:20]),.I5(N_1832),.LO(reg3_17[20:20]));
defparam desc978.INIT=64'hF0FFF4FFF000F400;
  LUT6_L desc979(.I0(N_527_i),.I1(reg3_14_sqmuxa),.I2(t_1[14:14]),.I3(N_1841),.I4(\d_cnst_sn.reg3_17_6_1 [14:14]),.I5(N_1826),.LO(reg3_17[14:14]));
defparam desc979.INIT=64'hBFFF00FFBF000000;
  LUT6_L desc980(.I0(N_527_i),.I1(reg3_14_sqmuxa),.I2(N_1841),.I3(\d_cnst_sn.reg3_17_6_1 [18:18]),.I4(t_1[18:18]),.I5(N_1830),.LO(reg3_17[18:18]));
defparam desc980.INIT=64'hBF0FFF0FB000F000;
  LUT6_L desc981(.I0(N_527_i),.I1(reg3_14_sqmuxa),.I2(t_1[12:12]),.I3(N_1841),.I4(\d_cnst_sn.reg3_17_6_1 [12:12]),.I5(N_1824),.LO(reg3_17[12:12]));
defparam desc981.INIT=64'hBFFF00FFBF000000;
  LUT6_L desc982(.I0(N_527_i),.I1(reg3_14_sqmuxa),.I2(N_1841),.I3(\d_cnst_sn.reg3_17_6_1 [17:17]),.I4(t_1[17:17]),.I5(N_1829),.LO(reg3_17[17:17]));
defparam desc982.INIT=64'hBF0FFF0FB000F000;
  LUT6_L desc983(.I0(N_527_i),.I1(reg3_14_sqmuxa),.I2(N_1841),.I3(\d_cnst_sn.reg3_17_6_1 [15:15]),.I4(t_1[15:15]),.I5(N_1827),.LO(reg3_17[15:15]));
defparam desc983.INIT=64'hBF0FFF0FB000F000;
  LUT6_L desc984(.I0(N_527_i),.I1(reg3_14_sqmuxa),.I2(\d_cnst_sn.reg3_17_6_0 [26:26]),.I3(N_1841),.I4(t_1[26:26]),.I5(N_1838),.LO(reg3_17[26:26]));
defparam desc984.INIT=64'hF0FFF4FFF000F400;
  LUT6_L desc985(.I0(N_527_i),.I1(reg3_14_sqmuxa),.I2(\d_cnst_sn.reg3_17_6_0 [25:25]),.I3(N_1841),.I4(t_1[25:25]),.I5(N_1837),.LO(reg3_17[25:25]));
defparam desc985.INIT=64'hF0FFF4FFF000F400;
  LUT6_L desc986(.I0(N_1810),.I1(reg3_17_a0[24:24]),.I2(\d_cnst_sn.reg3_17_a1_2 [24:24]),.I3(\d_cnst_sn.reg3_17_0_tz [24:24]),.I4(t_1[24:24]),.I5(N_1743),.LO(reg3_17[24:24]));
defparam desc986.INIT=64'hFFDDFFFDEECCFEFC;
  LUT6_L desc987(.I0(N_1810),.I1(reg3_17_a0[23:23]),.I2(\d_cnst_sn.reg3_17_a1_2 [24:24]),.I3(\d_cnst_sn.reg3_17_0_tz [23:23]),.I4(t_1[23:23]),.I5(N_1742),.LO(reg3_17[23:23]));
defparam desc987.INIT=64'hFFDDFFFDEECCFEFC;
  LUT6_L desc988(.I0(N_1810),.I1(reg3_17_a0[22:22]),.I2(\d_cnst_sn.reg3_17_a1_2 [24:24]),.I3(\d_cnst_sn.reg3_17_0_tz [22:22]),.I4(t_1[22:22]),.I5(N_1741),.LO(reg3_17[22:22]));
defparam desc988.INIT=64'hFFDDFFFDEECCFEFC;
  LUT6_L desc989(.I0(N_1810),.I1(\d_cnst_sn.reg3_17_0_tz [21:21]),.I2(reg3_17_a0[21:21]),.I3(\d_cnst_sn.reg3_17_a1_2 [24:24]),.I4(t_1[21:21]),.I5(N_1740),.LO(reg3_17[21:21]));
defparam desc989.INIT=64'hFDFDFFFDF8F8FFF8;
  LUT6_L desc990(.I0(N_1810),.I1(\d_cnst_sn.reg3_17_sn_m7_0 ),.I2(reg3_14_sqmuxa),.I3(reg3_N_7_i_RNO),.I4(N_1815),.I5(t_6[3:3]),.LO(\d_cnst_sn.reg3_N_7_i ));
defparam desc990.INIT=64'hF7FF8088777F0008;
  LUT5 desc991(.I0(datai[20:20]),.I1(inf_abs0_2[31:31]),.I2(inf_abs0_2[27:27]),.I3(inf_abs0_2[28:28]),.I4(r_4[20:20]),.O(un11_reg0_axb_20));
defparam desc991.INIT=32'hDDDF2220;
  LUT4 desc992(.I0(datai[20:20]),.I1(inf_abs0_2[31:31]),.I2(inf_abs0_2[27:27]),.I3(inf_abs0_2[28:28]),.O(m_2[20:20]));
defparam desc992.INIT=16'h2220;
  LUT5 desc993(.I0(datai[21:21]),.I1(inf_abs0_2[31:31]),.I2(inf_abs0_2[27:27]),.I3(inf_abs0_2[28:28]),.I4(r_4[21:21]),.O(un11_reg0_axb_21));
defparam desc993.INIT=32'hDDDF2220;
  LUT4 desc994(.I0(datai[21:21]),.I1(inf_abs0_2[31:31]),.I2(inf_abs0_2[27:27]),.I3(inf_abs0_2[28:28]),.O(m_2[21:21]));
defparam desc994.INIT=16'h2220;
  LUT5 desc995(.I0(datai[22:22]),.I1(inf_abs0_2[31:31]),.I2(inf_abs0_2[27:27]),.I3(inf_abs0_2[28:28]),.I4(r_4[22:22]),.O(un11_reg0_axb_22));
defparam desc995.INIT=32'hDDDF2220;
  LUT4 desc996(.I0(datai[22:22]),.I1(inf_abs0_2[31:31]),.I2(inf_abs0_2[27:27]),.I3(inf_abs0_2[28:28]),.O(m_2[22:22]));
defparam desc996.INIT=16'h2220;
  LUT5 desc997(.I0(datai[23:23]),.I1(inf_abs0_2[31:31]),.I2(inf_abs0_2[27:27]),.I3(inf_abs0_2[28:28]),.I4(r_4[23:23]),.O(un11_reg0_axb_23));
defparam desc997.INIT=32'hDDDF2220;
  LUT4 desc998(.I0(datai[23:23]),.I1(inf_abs0_2[31:31]),.I2(inf_abs0_2[27:27]),.I3(inf_abs0_2[28:28]),.O(m_2[23:23]));
defparam desc998.INIT=16'h2220;
  LUT5 desc999(.I0(datai[24:24]),.I1(inf_abs0_2[31:31]),.I2(inf_abs0_2[27:27]),.I3(inf_abs0_2[28:28]),.I4(r_4[24:24]),.O(un11_reg0_axb_24));
defparam desc999.INIT=32'hDDDF2220;
  LUT4 desc1000(.I0(datai[24:24]),.I1(inf_abs0_2[31:31]),.I2(inf_abs0_2[27:27]),.I3(inf_abs0_2[28:28]),.O(m_2[24:24]));
defparam desc1000.INIT=16'h2220;
  LUT5 desc1001(.I0(datai[25:25]),.I1(inf_abs0_2[31:31]),.I2(inf_abs0_2[27:27]),.I3(inf_abs0_2[28:28]),.I4(r_4[25:25]),.O(un11_reg0_axb_25));
defparam desc1001.INIT=32'hDDDF2220;
  LUT4 desc1002(.I0(datai[25:25]),.I1(inf_abs0_2[31:31]),.I2(inf_abs0_2[27:27]),.I3(inf_abs0_2[28:28]),.O(m_2[25:25]));
defparam desc1002.INIT=16'h2220;
  LUT5 desc1003(.I0(datai[26:26]),.I1(inf_abs0_2[31:31]),.I2(inf_abs0_2[27:27]),.I3(inf_abs0_2[28:28]),.I4(r_4[26:26]),.O(un11_reg0_axb_26));
defparam desc1003.INIT=32'hDDDF2220;
  LUT4 desc1004(.I0(datai[26:26]),.I1(inf_abs0_2[31:31]),.I2(inf_abs0_2[27:27]),.I3(inf_abs0_2[28:28]),.O(m_2[26:26]));
defparam desc1004.INIT=16'h2220;
  LUT5 desc1005(.I0(datai[27:27]),.I1(inf_abs0_2[31:31]),.I2(inf_abs0_2[27:27]),.I3(inf_abs0_2[28:28]),.I4(r_4[27:27]),.O(un11_reg0_axb_27));
defparam desc1005.INIT=32'hDDDF2220;
  LUT4 desc1006(.I0(datai[27:27]),.I1(inf_abs0_2[31:31]),.I2(inf_abs0_2[27:27]),.I3(inf_abs0_2[28:28]),.O(m_2[27:27]));
defparam desc1006.INIT=16'h2220;
  LUT5 desc1007(.I0(datai[28:28]),.I1(inf_abs0_2[31:31]),.I2(inf_abs0_2[27:27]),.I3(inf_abs0_2[28:28]),.I4(r_4[28:28]),.O(un11_reg0_axb_28));
defparam desc1007.INIT=32'hDDDF2220;
  LUT4 desc1008(.I0(datai[28:28]),.I1(inf_abs0_2[31:31]),.I2(inf_abs0_2[27:27]),.I3(inf_abs0_2[28:28]),.O(m_2[28:28]));
defparam desc1008.INIT=16'h2220;
  LUT5 desc1009(.I0(inf_abs0_2[31:31]),.I1(inf_abs0_2[29:29]),.I2(N_920),.I3(N_952),.I4(m_2[5:5]),.O(un32_reg0_axb_5));
defparam desc1009.INIT=32'hF4B00B4F;
  LUT5 desc1010(.I0(inf_abs0_2[31:31]),.I1(inf_abs0_2[29:29]),.I2(N_921),.I3(N_953),.I4(m_2[6:6]),.O(un32_reg0_axb_6));
defparam desc1010.INIT=32'hF4B00B4F;
  LUT5 desc1011(.I0(inf_abs0_2[31:31]),.I1(inf_abs0_2[29:29]),.I2(N_922),.I3(N_954),.I4(m_2[7:7]),.O(un32_reg0_axb_7));
defparam desc1011.INIT=32'hF4B00B4F;
  LUT5 desc1012(.I0(inf_abs0_2[31:31]),.I1(inf_abs0_2[29:29]),.I2(N_923),.I3(N_955),.I4(m_2[8:8]),.O(un32_reg0_axb_8));
defparam desc1012.INIT=32'hF4B00B4F;
  LUT5 desc1013(.I0(inf_abs0_2[31:31]),.I1(inf_abs0_2[29:29]),.I2(N_924),.I3(N_956),.I4(m_2[9:9]),.O(un32_reg0_axb_9));
defparam desc1013.INIT=32'hF4B00B4F;
  LUT5 desc1014(.I0(inf_abs0_2[31:31]),.I1(inf_abs0_2[29:29]),.I2(N_925),.I3(N_957),.I4(m_2[10:10]),.O(un32_reg0_axb_10));
defparam desc1014.INIT=32'hF4B00B4F;
  LUT5 desc1015(.I0(inf_abs0_2[31:31]),.I1(inf_abs0_2[29:29]),.I2(N_926),.I3(N_958),.I4(m_2[11:11]),.O(un32_reg0_axb_11));
defparam desc1015.INIT=32'hF4B00B4F;
  LUT5 desc1016(.I0(inf_abs0_2[31:31]),.I1(inf_abs0_2[29:29]),.I2(N_927),.I3(N_959),.I4(m_2[12:12]),.O(un32_reg0_axb_12));
defparam desc1016.INIT=32'hF4B00B4F;
  LUT5 desc1017(.I0(inf_abs0_2[31:31]),.I1(inf_abs0_2[29:29]),.I2(N_928),.I3(N_960),.I4(m_2[13:13]),.O(un32_reg0_axb_13));
defparam desc1017.INIT=32'hF4B00B4F;
  LUT5 desc1018(.I0(inf_abs0_2[31:31]),.I1(inf_abs0_2[29:29]),.I2(N_929),.I3(N_961),.I4(m_2[14:14]),.O(un32_reg0_axb_14));
defparam desc1018.INIT=32'hF4B00B4F;
  LUT5 desc1019(.I0(inf_abs0_2[31:31]),.I1(inf_abs0_2[29:29]),.I2(N_930),.I3(N_962),.I4(m_2[15:15]),.O(un32_reg0_axb_15));
defparam desc1019.INIT=32'hF4B00B4F;
  LUT5 desc1020(.I0(inf_abs0_2[31:31]),.I1(inf_abs0_2[29:29]),.I2(N_931),.I3(N_963),.I4(m_2[16:16]),.O(un32_reg0_axb_16));
defparam desc1020.INIT=32'hF4B00B4F;
  LUT5 desc1021(.I0(inf_abs0_2[31:31]),.I1(inf_abs0_2[29:29]),.I2(N_932),.I3(N_964),.I4(m_2[17:17]),.O(un32_reg0_axb_17));
defparam desc1021.INIT=32'hF4B00B4F;
  LUT5 desc1022(.I0(inf_abs0_2[31:31]),.I1(inf_abs0_2[29:29]),.I2(N_933),.I3(N_965),.I4(m_2[18:18]),.O(un32_reg0_axb_18));
defparam desc1022.INIT=32'hF4B00B4F;
  LUT5 desc1023(.I0(inf_abs0_2[31:31]),.I1(inf_abs0_2[29:29]),.I2(N_934),.I3(N_2722),.I4(m_2[19:19]),.O(un32_reg0_axb_19));
defparam desc1023.INIT=32'hF4B00B4F;
  XORCY t_1_s_31(.LI(r_4[31:31]),.CI(t_1_cry_30),.O(t_1[31:31]));
  XORCY t_1_s_30(.LI(N_4571_i),.CI(t_1_cry_29),.O(t_1[30:30]));
  MUXCY_L t_1_cry_30_cZ(.DI(VCC),.CI(t_1_cry_29),.S(N_4571_i),.LO(t_1_cry_30));
  XORCY t_1_s_29(.LI(N_4570_i),.CI(t_1_cry_28),.O(t_1[29:29]));
  MUXCY_L t_1_cry_29_cZ(.DI(VCC),.CI(t_1_cry_28),.S(N_4570_i),.LO(t_1_cry_29));
  XORCY t_1_s_28(.LI(N_4569_i),.CI(t_1_cry_27),.O(t_1[28:28]));
  MUXCY_L t_1_cry_28_cZ(.DI(VCC),.CI(t_1_cry_27),.S(N_4569_i),.LO(t_1_cry_28));
  XORCY t_1_s_27(.LI(N_4568_i),.CI(t_1_cry_26),.O(t_1[27:27]));
  MUXCY_L t_1_cry_27_cZ(.DI(VCC),.CI(t_1_cry_26),.S(N_4568_i),.LO(t_1_cry_27));
  XORCY t_1_s_26(.LI(N_4567_i),.CI(t_1_cry_25),.O(t_1[26:26]));
  MUXCY_L t_1_cry_26_cZ(.DI(VCC),.CI(t_1_cry_25),.S(N_4567_i),.LO(t_1_cry_26));
  XORCY t_1_s_25(.LI(N_4566_i),.CI(t_1_cry_24),.O(t_1[25:25]));
  MUXCY_L t_1_cry_25_cZ(.DI(VCC),.CI(t_1_cry_24),.S(N_4566_i),.LO(t_1_cry_25));
  XORCY t_1_s_24(.LI(N_4565_i),.CI(t_1_cry_23),.O(t_1[24:24]));
  MUXCY_L t_1_cry_24_cZ(.DI(VCC),.CI(t_1_cry_23),.S(N_4565_i),.LO(t_1_cry_24));
  XORCY t_1_s_23(.LI(N_4564_i),.CI(t_1_cry_22),.O(t_1[23:23]));
  MUXCY_L t_1_cry_23_cZ(.DI(VCC),.CI(t_1_cry_22),.S(N_4564_i),.LO(t_1_cry_23));
  XORCY t_1_s_22(.LI(N_4563_i),.CI(t_1_cry_21),.O(t_1[22:22]));
  MUXCY_L t_1_cry_22_cZ(.DI(VCC),.CI(t_1_cry_21),.S(N_4563_i),.LO(t_1_cry_22));
  XORCY t_1_s_21(.LI(N_4562_i),.CI(t_1_cry_20),.O(t_1[21:21]));
  MUXCY_L t_1_cry_21_cZ(.DI(VCC),.CI(t_1_cry_20),.S(N_4562_i),.LO(t_1_cry_21));
  XORCY t_1_s_20(.LI(N_4561_i),.CI(t_1_cry_19),.O(t_1[20:20]));
  MUXCY_L t_1_cry_20_cZ(.DI(VCC),.CI(t_1_cry_19),.S(N_4561_i),.LO(t_1_cry_20));
  XORCY t_1_s_19(.LI(N_4560_i),.CI(t_1_cry_18),.O(t_1[19:19]));
  MUXCY_L t_1_cry_19_cZ(.DI(VCC),.CI(t_1_cry_18),.S(N_4560_i),.LO(t_1_cry_19));
  XORCY t_1_s_18(.LI(N_4559_i),.CI(t_1_cry_17),.O(t_1[18:18]));
  MUXCY_L t_1_cry_18_cZ(.DI(VCC),.CI(t_1_cry_17),.S(N_4559_i),.LO(t_1_cry_18));
  XORCY t_1_s_17(.LI(N_4558_i),.CI(t_1_cry_16),.O(t_1[17:17]));
  MUXCY_L t_1_cry_17_cZ(.DI(VCC),.CI(t_1_cry_16),.S(N_4558_i),.LO(t_1_cry_17));
  XORCY t_1_s_16(.LI(N_4557_i),.CI(t_1_cry_15),.O(t_1[16:16]));
  MUXCY_L t_1_cry_16_cZ(.DI(VCC),.CI(t_1_cry_15),.S(N_4557_i),.LO(t_1_cry_16));
  XORCY t_1_s_15(.LI(N_4556_i),.CI(t_1_cry_14),.O(t_1[15:15]));
  MUXCY_L t_1_cry_15_cZ(.DI(VCC),.CI(t_1_cry_14),.S(N_4556_i),.LO(t_1_cry_15));
  XORCY t_1_s_14(.LI(N_4555_i),.CI(t_1_cry_13),.O(t_1[14:14]));
  MUXCY_L t_1_cry_14_cZ(.DI(VCC),.CI(t_1_cry_13),.S(N_4555_i),.LO(t_1_cry_14));
  XORCY t_1_s_13(.LI(N_4554_i),.CI(t_1_cry_12),.O(t_1[13:13]));
  MUXCY_L t_1_cry_13_cZ(.DI(VCC),.CI(t_1_cry_12),.S(N_4554_i),.LO(t_1_cry_13));
  XORCY t_1_s_12(.LI(N_4553_i),.CI(t_1_cry_11),.O(t_1[12:12]));
  MUXCY_L t_1_cry_12_cZ(.DI(VCC),.CI(t_1_cry_11),.S(N_4553_i),.LO(t_1_cry_12));
  XORCY t_1_s_11(.LI(N_4552_i),.CI(t_1_cry_10),.O(t_1[11:11]));
  MUXCY_L t_1_cry_11_cZ(.DI(VCC),.CI(t_1_cry_10),.S(N_4552_i),.LO(t_1_cry_11));
  XORCY t_1_s_10(.LI(N_4551_i),.CI(t_1_cry_9),.O(t_1[10:10]));
  MUXCY_L t_1_cry_10_cZ(.DI(VCC),.CI(t_1_cry_9),.S(N_4551_i),.LO(t_1_cry_10));
  XORCY t_1_s_9(.LI(N_4550_i),.CI(t_1_cry_8),.O(t_1[9:9]));
  MUXCY_L t_1_cry_9_cZ(.DI(VCC),.CI(t_1_cry_8),.S(N_4550_i),.LO(t_1_cry_9));
  XORCY t_1_s_8(.LI(N_4549_i),.CI(t_1_cry_7),.O(t_1[8:8]));
  MUXCY_L t_1_cry_8_cZ(.DI(VCC),.CI(t_1_cry_7),.S(N_4549_i),.LO(t_1_cry_8));
  XORCY t_1_s_7(.LI(N_4548_i),.CI(t_1_cry_6),.O(t_1[7:7]));
  MUXCY_L t_1_cry_7_cZ(.DI(VCC),.CI(t_1_cry_6),.S(N_4548_i),.LO(t_1_cry_7));
  XORCY t_1_s_6(.LI(N_4547_i),.CI(t_1_cry_5),.O(t_1[6:6]));
  MUXCY_L t_1_cry_6_cZ(.DI(VCC),.CI(t_1_cry_5),.S(N_4547_i),.LO(t_1_cry_6));
  XORCY t_1_s_5(.LI(N_4546_i),.CI(t_1_cry_4),.O(t_1[5:5]));
  MUXCY_L t_1_cry_5_cZ(.DI(VCC),.CI(t_1_cry_4),.S(N_4546_i),.LO(t_1_cry_5));
  XORCY t_1_s_4(.LI(N_4545_i),.CI(t_1_cry_3),.O(t_1[4:4]));
  MUXCY_L t_1_cry_4_cZ(.DI(VCC),.CI(t_1_cry_3),.S(N_4545_i),.LO(t_1_cry_4));
  XORCY t_1_s_3(.LI(N_4544_i),.CI(t_1_cry_2),.O(t_1[3:3]));
  MUXCY_L t_1_cry_3_cZ(.DI(VCC),.CI(t_1_cry_2),.S(N_4544_i),.LO(t_1_cry_3));
  XORCY t_1_s_2(.LI(N_4543_i),.CI(t_1_cry_1),.O(t_1[2:2]));
  MUXCY_L t_1_cry_2_cZ(.DI(VCC),.CI(t_1_cry_1),.S(N_4543_i),.LO(t_1_cry_2));
  XORCY t_1_s_1(.LI(N_4542_i),.CI(t_1_cry_0),.O(t_1[1:1]));
  MUXCY_L t_1_cry_1_cZ(.DI(VCC),.CI(t_1_cry_0),.S(N_4542_i),.LO(t_1_cry_1));
  XORCY t_1_s_0(.LI(N_4541_i),.CI(t_1_cry_0_cy),.O(t_1[0:0]));
  MUXCY_L t_1_cry_0_cZ(.DI(VCC),.CI(t_1_cry_0_cy),.S(N_4541_i),.LO(t_1_cry_0));
  XORCY un3_reg3_s_25_cZ(.LI(un3_reg3_axb_25),.CI(un3_reg3_cry_24),.O(un3_reg3_s_25));
  MUXCY un3_reg3_cry_25_cZ(.DI(GND),.CI(un3_reg3_cry_24),.S(un3_reg3_axb_25),.O(un3_reg3_cry_25_0));
  XORCY un3_reg3_s_24_cZ(.LI(un3_reg3_axb_24),.CI(un3_reg3_cry_23),.O(un3_reg3_s_24));
  MUXCY_L un3_reg3_cry_24_cZ(.DI(GND),.CI(un3_reg3_cry_23),.S(un3_reg3_axb_24),.LO(un3_reg3_cry_24));
  XORCY un3_reg3_s_23_cZ(.LI(un3_reg3_axb_23),.CI(un3_reg3_cry_22),.O(un3_reg3_s_23));
  MUXCY_L un3_reg3_cry_23_cZ(.DI(GND),.CI(un3_reg3_cry_22),.S(un3_reg3_axb_23),.LO(un3_reg3_cry_23));
  XORCY un3_reg3_s_22_cZ(.LI(un3_reg3_axb_22),.CI(un3_reg3_cry_21),.O(un3_reg3_s_22));
  MUXCY_L un3_reg3_cry_22_cZ(.DI(GND),.CI(un3_reg3_cry_21),.S(un3_reg3_axb_22),.LO(un3_reg3_cry_22));
  XORCY un3_reg3_s_21_cZ(.LI(un3_reg3_axb_21),.CI(un3_reg3_cry_20),.O(un3_reg3_s_21));
  MUXCY_L un3_reg3_cry_21_cZ(.DI(GND),.CI(un3_reg3_cry_20),.S(un3_reg3_axb_21),.LO(un3_reg3_cry_21));
  XORCY un3_reg3_s_20_cZ(.LI(un3_reg3_axb_20),.CI(un3_reg3_cry_19),.O(un3_reg3_s_20));
  MUXCY_L un3_reg3_cry_20_cZ(.DI(GND),.CI(un3_reg3_cry_19),.S(un3_reg3_axb_20),.LO(un3_reg3_cry_20));
  XORCY un3_reg3_s_19_cZ(.LI(un3_reg3_axb_19),.CI(un3_reg3_cry_18),.O(un3_reg3_s_19));
  MUXCY_L un3_reg3_cry_19_cZ(.DI(GND),.CI(un3_reg3_cry_18),.S(un3_reg3_axb_19),.LO(un3_reg3_cry_19));
  XORCY un3_reg3_s_18_cZ(.LI(un3_reg3_axb_18),.CI(un3_reg3_cry_17),.O(un3_reg3_s_18));
  MUXCY_L un3_reg3_cry_18_cZ(.DI(GND),.CI(un3_reg3_cry_17),.S(un3_reg3_axb_18),.LO(un3_reg3_cry_18));
  XORCY un3_reg3_s_17_cZ(.LI(un3_reg3_axb_17),.CI(un3_reg3_cry_16),.O(un3_reg3_s_17));
  MUXCY_L un3_reg3_cry_17_cZ(.DI(GND),.CI(un3_reg3_cry_16),.S(un3_reg3_axb_17),.LO(un3_reg3_cry_17));
  XORCY un3_reg3_s_16_cZ(.LI(un3_reg3_axb_16),.CI(un3_reg3_cry_15),.O(un3_reg3_s_16));
  MUXCY_L un3_reg3_cry_16_cZ(.DI(GND),.CI(un3_reg3_cry_15),.S(un3_reg3_axb_16),.LO(un3_reg3_cry_16));
  XORCY un3_reg3_s_15_cZ(.LI(un3_reg3_axb_15),.CI(un3_reg3_cry_14),.O(un3_reg3_s_15));
  MUXCY_L un3_reg3_cry_15_cZ(.DI(GND),.CI(un3_reg3_cry_14),.S(un3_reg3_axb_15),.LO(un3_reg3_cry_15));
  XORCY un3_reg3_s_14_cZ(.LI(un3_reg3_axb_14),.CI(un3_reg3_cry_13),.O(un3_reg3_s_14));
  MUXCY_L un3_reg3_cry_14_cZ(.DI(GND),.CI(un3_reg3_cry_13),.S(un3_reg3_axb_14),.LO(un3_reg3_cry_14));
  XORCY un3_reg3_s_13_cZ(.LI(un3_reg3_axb_13),.CI(un3_reg3_cry_12),.O(un3_reg3_s_13));
  MUXCY_L un3_reg3_cry_13_cZ(.DI(GND),.CI(un3_reg3_cry_12),.S(un3_reg3_axb_13),.LO(un3_reg3_cry_13));
  XORCY un3_reg3_s_12_cZ(.LI(un3_reg3_axb_12),.CI(un3_reg3_cry_11),.O(un3_reg3_s_12));
  MUXCY_L un3_reg3_cry_12_cZ(.DI(GND),.CI(un3_reg3_cry_11),.S(un3_reg3_axb_12),.LO(un3_reg3_cry_12));
  XORCY un3_reg3_s_11_cZ(.LI(un3_reg3_axb_11),.CI(un3_reg3_cry_10),.O(un3_reg3_s_11));
  MUXCY_L un3_reg3_cry_11_cZ(.DI(GND),.CI(un3_reg3_cry_10),.S(un3_reg3_axb_11),.LO(un3_reg3_cry_11));
  XORCY un3_reg3_s_10_cZ(.LI(un3_reg3_axb_10),.CI(un3_reg3_cry_9),.O(un3_reg3_s_10));
  MUXCY_L un3_reg3_cry_10_cZ(.DI(GND),.CI(un3_reg3_cry_9),.S(un3_reg3_axb_10),.LO(un3_reg3_cry_10));
  XORCY un3_reg3_s_9_cZ(.LI(un3_reg3_axb_9),.CI(un3_reg3_cry_8),.O(un3_reg3_s_9));
  MUXCY_L un3_reg3_cry_9_cZ(.DI(GND),.CI(un3_reg3_cry_8),.S(un3_reg3_axb_9),.LO(un3_reg3_cry_9));
  XORCY un3_reg3_s_8_cZ(.LI(un3_reg3_axb_8),.CI(un3_reg3_cry_7),.O(un3_reg3_s_8));
  MUXCY_L un3_reg3_cry_8_cZ(.DI(GND),.CI(un3_reg3_cry_7),.S(un3_reg3_axb_8),.LO(un3_reg3_cry_8));
  XORCY un3_reg3_s_7_cZ(.LI(un3_reg3_axb_7),.CI(un3_reg3_cry_6),.O(un3_reg3_s_7));
  MUXCY_L un3_reg3_cry_7_cZ(.DI(GND),.CI(un3_reg3_cry_6),.S(un3_reg3_axb_7),.LO(un3_reg3_cry_7));
  XORCY un3_reg3_s_6_cZ(.LI(un3_reg3_axb_6),.CI(un3_reg3_cry_5),.O(un3_reg3_s_6));
  MUXCY_L un3_reg3_cry_6_cZ(.DI(GND),.CI(un3_reg3_cry_5),.S(un3_reg3_axb_6),.LO(un3_reg3_cry_6));
  XORCY un3_reg3_s_5_cZ(.LI(un3_reg3_axb_5),.CI(un3_reg3_cry_4),.O(un3_reg3_s_5));
  MUXCY_L un3_reg3_cry_5_cZ(.DI(GND),.CI(un3_reg3_cry_4),.S(un3_reg3_axb_5),.LO(un3_reg3_cry_5));
  XORCY un3_reg3_s_4_cZ(.LI(un3_reg3_axb_4),.CI(un3_reg3_cry_3),.O(un3_reg3_s_4));
  MUXCY_L un3_reg3_cry_4_cZ(.DI(GND),.CI(un3_reg3_cry_3),.S(un3_reg3_axb_4),.LO(un3_reg3_cry_4));
  XORCY un3_reg3_s_3_cZ(.LI(un3_reg3_axb_3),.CI(un3_reg3_cry_2),.O(un3_reg3_s_3));
  MUXCY_L un3_reg3_cry_3_cZ(.DI(GND),.CI(un3_reg3_cry_2),.S(un3_reg3_axb_3),.LO(un3_reg3_cry_3));
  XORCY un3_reg3_s_2_cZ(.LI(un3_reg3_axb_2),.CI(un3_reg3_cry_1),.O(un3_reg3_s_2));
  MUXCY_L un3_reg3_cry_2_cZ(.DI(GND),.CI(un3_reg3_cry_1),.S(un3_reg3_axb_2),.LO(un3_reg3_cry_2));
  XORCY un3_reg3_s_1_cZ(.LI(un3_reg3_axb_1),.CI(reg3[3:3]),.O(un3_reg3_s_1));
  MUXCY_L un3_reg3_cry_1_cZ(.DI(GND),.CI(reg3[3:3]),.S(un3_reg3_axb_1),.LO(un3_reg3_cry_1));
  XORCY un1_inf_abs0_0_s_19(.LI(un1_inf_abs0_0_axb_19),.CI(un1_inf_abs0_0_cry_18),.O(un1_inf_abs0_11[19:19]));
  XORCY un1_inf_abs0_0_s_18(.LI(un1_inf_abs0_0_axb_18),.CI(un1_inf_abs0_0_cry_17),.O(un1_inf_abs0_11[18:18]));
  MUXCY_L un1_inf_abs0_0_cry_18_cZ(.DI(inf_abs0_2[18:18]),.CI(un1_inf_abs0_0_cry_17),.S(un1_inf_abs0_0_axb_18),.LO(un1_inf_abs0_0_cry_18));
  XORCY un1_inf_abs0_0_s_17(.LI(un1_inf_abs0_0_axb_17),.CI(un1_inf_abs0_0_cry_16),.O(un1_inf_abs0_11[17:17]));
  MUXCY_L un1_inf_abs0_0_cry_17_cZ(.DI(inf_abs0_2[17:17]),.CI(un1_inf_abs0_0_cry_16),.S(un1_inf_abs0_0_axb_17),.LO(un1_inf_abs0_0_cry_17));
  XORCY un1_inf_abs0_0_s_16(.LI(un1_inf_abs0_0_axb_16),.CI(un1_inf_abs0_0_cry_15),.O(un1_inf_abs0_11[16:16]));
  MUXCY_L un1_inf_abs0_0_cry_16_cZ(.DI(inf_abs0_2[16:16]),.CI(un1_inf_abs0_0_cry_15),.S(un1_inf_abs0_0_axb_16),.LO(un1_inf_abs0_0_cry_16));
  XORCY un1_inf_abs0_0_s_15(.LI(un1_inf_abs0_0_axb_15),.CI(un1_inf_abs0_0_cry_14),.O(un1_inf_abs0_11[15:15]));
  MUXCY_L un1_inf_abs0_0_cry_15_cZ(.DI(inf_abs0_2[15:15]),.CI(un1_inf_abs0_0_cry_14),.S(un1_inf_abs0_0_axb_15),.LO(un1_inf_abs0_0_cry_15));
  XORCY un1_inf_abs0_0_s_14(.LI(un1_inf_abs0_0_axb_14),.CI(un1_inf_abs0_0_cry_13),.O(un1_inf_abs0_11[14:14]));
  MUXCY_L un1_inf_abs0_0_cry_14_cZ(.DI(inf_abs0_2[14:14]),.CI(un1_inf_abs0_0_cry_13),.S(un1_inf_abs0_0_axb_14),.LO(un1_inf_abs0_0_cry_14));
  XORCY un1_inf_abs0_0_s_13(.LI(un1_inf_abs0_0_axb_13),.CI(un1_inf_abs0_0_cry_12),.O(un1_inf_abs0_11[13:13]));
  MUXCY_L un1_inf_abs0_0_cry_13_cZ(.DI(inf_abs0_2[13:13]),.CI(un1_inf_abs0_0_cry_12),.S(un1_inf_abs0_0_axb_13),.LO(un1_inf_abs0_0_cry_13));
  XORCY un1_inf_abs0_0_s_12(.LI(un1_inf_abs0_0_axb_12),.CI(un1_inf_abs0_0_cry_11),.O(un1_inf_abs0_11[12:12]));
  MUXCY_L un1_inf_abs0_0_cry_12_cZ(.DI(inf_abs0_2[12:12]),.CI(un1_inf_abs0_0_cry_11),.S(un1_inf_abs0_0_axb_12),.LO(un1_inf_abs0_0_cry_12));
  XORCY un1_inf_abs0_0_s_11(.LI(un1_inf_abs0_0_axb_11),.CI(un1_inf_abs0_0_cry_10),.O(un1_inf_abs0_11[11:11]));
  MUXCY_L un1_inf_abs0_0_cry_11_cZ(.DI(inf_abs0_2[11:11]),.CI(un1_inf_abs0_0_cry_10),.S(un1_inf_abs0_0_axb_11),.LO(un1_inf_abs0_0_cry_11));
  XORCY un1_inf_abs0_0_s_10(.LI(un1_inf_abs0_0_axb_10),.CI(un1_inf_abs0_0_cry_9),.O(un1_inf_abs0_11[10:10]));
  MUXCY_L un1_inf_abs0_0_cry_10_cZ(.DI(inf_abs0_2[10:10]),.CI(un1_inf_abs0_0_cry_9),.S(un1_inf_abs0_0_axb_10),.LO(un1_inf_abs0_0_cry_10));
  XORCY un1_inf_abs0_0_s_9(.LI(un1_inf_abs0_0_axb_9),.CI(un1_inf_abs0_0_cry_8),.O(un1_inf_abs0_11[9:9]));
  MUXCY_L un1_inf_abs0_0_cry_9_cZ(.DI(inf_abs0_2[9:9]),.CI(un1_inf_abs0_0_cry_8),.S(un1_inf_abs0_0_axb_9),.LO(un1_inf_abs0_0_cry_9));
  XORCY un1_inf_abs0_0_s_8(.LI(un1_inf_abs0_0_axb_8),.CI(un1_inf_abs0_0_cry_7),.O(un1_inf_abs0_11[8:8]));
  MUXCY_L un1_inf_abs0_0_cry_8_cZ(.DI(inf_abs0_2[8:8]),.CI(un1_inf_abs0_0_cry_7),.S(un1_inf_abs0_0_axb_8),.LO(un1_inf_abs0_0_cry_8));
  XORCY un1_inf_abs0_0_s_7(.LI(un1_inf_abs0_0_axb_7),.CI(un1_inf_abs0_0_cry_6),.O(un1_inf_abs0_11[7:7]));
  MUXCY_L un1_inf_abs0_0_cry_7_cZ(.DI(inf_abs0_2[7:7]),.CI(un1_inf_abs0_0_cry_6),.S(un1_inf_abs0_0_axb_7),.LO(un1_inf_abs0_0_cry_7));
  XORCY un1_inf_abs0_0_s_6(.LI(un1_inf_abs0_0_axb_6),.CI(un1_inf_abs0_0_cry_5),.O(un1_inf_abs0_11[6:6]));
  MUXCY_L un1_inf_abs0_0_cry_6_cZ(.DI(inf_abs0_2[6:6]),.CI(un1_inf_abs0_0_cry_5),.S(un1_inf_abs0_0_axb_6),.LO(un1_inf_abs0_0_cry_6));
  XORCY un1_inf_abs0_0_s_5(.LI(un1_inf_abs0_0_axb_5),.CI(un1_inf_abs0_0_cry_4),.O(un1_inf_abs0_11[5:5]));
  MUXCY_L un1_inf_abs0_0_cry_5_cZ(.DI(inf_abs0_2[5:5]),.CI(un1_inf_abs0_0_cry_4),.S(un1_inf_abs0_0_axb_5),.LO(un1_inf_abs0_0_cry_5));
  XORCY un1_inf_abs0_0_s_4(.LI(un1_inf_abs0_0_axb_4),.CI(un1_inf_abs0_0_cry_3),.O(un1_inf_abs0_11[4:4]));
  MUXCY_L un1_inf_abs0_0_cry_4_cZ(.DI(inf_abs0_2[4:4]),.CI(un1_inf_abs0_0_cry_3),.S(un1_inf_abs0_0_axb_4),.LO(un1_inf_abs0_0_cry_4));
  XORCY un1_inf_abs0_0_s_3(.LI(un1_inf_abs0_0_axb_3),.CI(un1_inf_abs0_0_cry_2),.O(un1_inf_abs0_11[3:3]));
  MUXCY_L un1_inf_abs0_0_cry_3_cZ(.DI(inf_abs0_2[3:3]),.CI(un1_inf_abs0_0_cry_2),.S(un1_inf_abs0_0_axb_3),.LO(un1_inf_abs0_0_cry_3));
  XORCY un1_inf_abs0_0_s_2(.LI(un1_inf_abs0_0_axb_2),.CI(un1_inf_abs0_0_cry_1),.O(un1_inf_abs0_11[2:2]));
  MUXCY_L un1_inf_abs0_0_cry_2_cZ(.DI(inf_abs0_2[2:2]),.CI(un1_inf_abs0_0_cry_1),.S(un1_inf_abs0_0_axb_2),.LO(un1_inf_abs0_0_cry_2));
  XORCY un1_inf_abs0_0_s_1(.LI(un1_inf_abs0_0_axb_1),.CI(un1_inf_abs0_0_cry_0),.O(un1_inf_abs0_11[1:1]));
  MUXCY_L un1_inf_abs0_0_cry_1_cZ(.DI(inf_abs0_2[1:1]),.CI(un1_inf_abs0_0_cry_0),.S(un1_inf_abs0_0_axb_1),.LO(un1_inf_abs0_0_cry_1));
  MUXCY_L un1_inf_abs0_0_cry_0_cZ(.DI(inf_abs0_2[0:0]),.CI(GND),.S(un1_inf_abs0_11[0:0]),.LO(un1_inf_abs0_0_cry_0));
  XORCY un1_inf_abs0_s_19(.LI(un1_inf_abs0_axb_19),.CI(un1_inf_abs0_cry_18),.O(un1_inf_abs0_10[19:19]));
  XORCY un1_inf_abs0_s_18(.LI(un1_inf_abs0_axb_18),.CI(un1_inf_abs0_cry_17),.O(un1_inf_abs0_10[18:18]));
  MUXCY_L un1_inf_abs0_cry_18_cZ(.DI(inf_abs0_2[18:18]),.CI(un1_inf_abs0_cry_17),.S(un1_inf_abs0_axb_18),.LO(un1_inf_abs0_cry_18));
  XORCY un1_inf_abs0_s_17(.LI(un1_inf_abs0_axb_17),.CI(un1_inf_abs0_cry_16),.O(un1_inf_abs0_10[17:17]));
  MUXCY_L un1_inf_abs0_cry_17_cZ(.DI(inf_abs0_2[17:17]),.CI(un1_inf_abs0_cry_16),.S(un1_inf_abs0_axb_17),.LO(un1_inf_abs0_cry_17));
  XORCY un1_inf_abs0_s_16(.LI(un1_inf_abs0_axb_16),.CI(un1_inf_abs0_cry_15),.O(un1_inf_abs0_10[16:16]));
  MUXCY_L un1_inf_abs0_cry_16_cZ(.DI(inf_abs0_2[16:16]),.CI(un1_inf_abs0_cry_15),.S(un1_inf_abs0_axb_16),.LO(un1_inf_abs0_cry_16));
  XORCY un1_inf_abs0_s_15(.LI(un1_inf_abs0_axb_15),.CI(un1_inf_abs0_cry_14),.O(un1_inf_abs0_10[15:15]));
  MUXCY_L un1_inf_abs0_cry_15_cZ(.DI(inf_abs0_2[15:15]),.CI(un1_inf_abs0_cry_14),.S(un1_inf_abs0_axb_15),.LO(un1_inf_abs0_cry_15));
  XORCY un1_inf_abs0_s_14(.LI(un1_inf_abs0_axb_14),.CI(un1_inf_abs0_cry_13),.O(un1_inf_abs0_10[14:14]));
  MUXCY_L un1_inf_abs0_cry_14_cZ(.DI(inf_abs0_2[14:14]),.CI(un1_inf_abs0_cry_13),.S(un1_inf_abs0_axb_14),.LO(un1_inf_abs0_cry_14));
  XORCY un1_inf_abs0_s_13(.LI(un1_inf_abs0_axb_13),.CI(un1_inf_abs0_cry_12),.O(un1_inf_abs0_10[13:13]));
  MUXCY_L un1_inf_abs0_cry_13_cZ(.DI(inf_abs0_2[13:13]),.CI(un1_inf_abs0_cry_12),.S(un1_inf_abs0_axb_13),.LO(un1_inf_abs0_cry_13));
  XORCY un1_inf_abs0_s_12(.LI(un1_inf_abs0_axb_12),.CI(un1_inf_abs0_cry_11),.O(un1_inf_abs0_10[12:12]));
  MUXCY_L un1_inf_abs0_cry_12_cZ(.DI(inf_abs0_2[12:12]),.CI(un1_inf_abs0_cry_11),.S(un1_inf_abs0_axb_12),.LO(un1_inf_abs0_cry_12));
  XORCY un1_inf_abs0_s_11(.LI(un1_inf_abs0_axb_11),.CI(un1_inf_abs0_cry_10),.O(un1_inf_abs0_10[11:11]));
  MUXCY_L un1_inf_abs0_cry_11_cZ(.DI(inf_abs0_2[11:11]),.CI(un1_inf_abs0_cry_10),.S(un1_inf_abs0_axb_11),.LO(un1_inf_abs0_cry_11));
  XORCY un1_inf_abs0_s_10(.LI(un1_inf_abs0_axb_10),.CI(un1_inf_abs0_cry_9),.O(un1_inf_abs0_10[10:10]));
  MUXCY_L un1_inf_abs0_cry_10_cZ(.DI(inf_abs0_2[10:10]),.CI(un1_inf_abs0_cry_9),.S(un1_inf_abs0_axb_10),.LO(un1_inf_abs0_cry_10));
  XORCY un1_inf_abs0_s_9(.LI(un1_inf_abs0_axb_9),.CI(un1_inf_abs0_cry_8),.O(un1_inf_abs0_10[9:9]));
  MUXCY_L un1_inf_abs0_cry_9_cZ(.DI(inf_abs0_2[9:9]),.CI(un1_inf_abs0_cry_8),.S(un1_inf_abs0_axb_9),.LO(un1_inf_abs0_cry_9));
  XORCY un1_inf_abs0_s_8(.LI(un1_inf_abs0_axb_8),.CI(un1_inf_abs0_cry_7),.O(un1_inf_abs0_10[8:8]));
  MUXCY_L un1_inf_abs0_cry_8_cZ(.DI(inf_abs0_2[8:8]),.CI(un1_inf_abs0_cry_7),.S(un1_inf_abs0_axb_8),.LO(un1_inf_abs0_cry_8));
  XORCY un1_inf_abs0_s_7(.LI(un1_inf_abs0_axb_7),.CI(un1_inf_abs0_cry_6),.O(un1_inf_abs0_10[7:7]));
  MUXCY_L un1_inf_abs0_cry_7_cZ(.DI(inf_abs0_2[7:7]),.CI(un1_inf_abs0_cry_6),.S(un1_inf_abs0_axb_7),.LO(un1_inf_abs0_cry_7));
  XORCY un1_inf_abs0_s_6(.LI(un1_inf_abs0_axb_6),.CI(un1_inf_abs0_cry_5),.O(un1_inf_abs0_10[6:6]));
  MUXCY_L un1_inf_abs0_cry_6_cZ(.DI(inf_abs0_2[6:6]),.CI(un1_inf_abs0_cry_5),.S(un1_inf_abs0_axb_6),.LO(un1_inf_abs0_cry_6));
  XORCY un1_inf_abs0_s_5(.LI(un1_inf_abs0_axb_5),.CI(un1_inf_abs0_cry_4),.O(un1_inf_abs0_10[5:5]));
  MUXCY_L un1_inf_abs0_cry_5_cZ(.DI(inf_abs0_2[5:5]),.CI(un1_inf_abs0_cry_4),.S(un1_inf_abs0_axb_5),.LO(un1_inf_abs0_cry_5));
  XORCY un1_inf_abs0_s_4(.LI(un1_inf_abs0_axb_4),.CI(un1_inf_abs0_cry_3),.O(un1_inf_abs0_10[4:4]));
  MUXCY_L un1_inf_abs0_cry_4_cZ(.DI(inf_abs0_2[4:4]),.CI(un1_inf_abs0_cry_3),.S(un1_inf_abs0_axb_4),.LO(un1_inf_abs0_cry_4));
  XORCY un1_inf_abs0_s_3(.LI(un1_inf_abs0_axb_3),.CI(un1_inf_abs0_cry_2),.O(un1_inf_abs0_10[3:3]));
  MUXCY_L un1_inf_abs0_cry_3_cZ(.DI(inf_abs0_2[3:3]),.CI(un1_inf_abs0_cry_2),.S(un1_inf_abs0_axb_3),.LO(un1_inf_abs0_cry_3));
  XORCY un1_inf_abs0_s_2(.LI(un1_inf_abs0_axb_2),.CI(un1_inf_abs0_cry_1),.O(un1_inf_abs0_10[2:2]));
  MUXCY_L un1_inf_abs0_cry_2_cZ(.DI(inf_abs0_2[2:2]),.CI(un1_inf_abs0_cry_1),.S(un1_inf_abs0_axb_2),.LO(un1_inf_abs0_cry_2));
  XORCY un1_inf_abs0_s_1(.LI(un1_inf_abs0_axb_1),.CI(un1_inf_abs0_cry_0),.O(un1_inf_abs0_10[1:1]));
  MUXCY_L un1_inf_abs0_cry_1_cZ(.DI(inf_abs0_2[1:1]),.CI(un1_inf_abs0_cry_0),.S(un1_inf_abs0_axb_1),.LO(un1_inf_abs0_cry_1));
  MUXCY_L un1_inf_abs0_cry_0_cZ(.DI(inf_abs0_2[0:0]),.CI(GND),.S(un1_inf_abs0_10[0:0]),.LO(un1_inf_abs0_cry_0));
  XORCY un32_reg0_s_29_cZ(.LI(un32_reg0_axb_29),.CI(un32_reg0_cry_28),.O(un32_reg0_s_29));
  XORCY un32_reg0_s_28_cZ(.LI(un32_reg0_axb_28),.CI(un32_reg0_cry_27),.O(un32_reg0_s_28));
  MUXCY_L un32_reg0_cry_28_cZ(.DI(r_4[28:28]),.CI(un32_reg0_cry_27),.S(un32_reg0_axb_28),.LO(un32_reg0_cry_28));
  XORCY un32_reg0_s_27_cZ(.LI(un32_reg0_axb_27),.CI(un32_reg0_cry_26),.O(un32_reg0_s_27));
  MUXCY_L un32_reg0_cry_27_cZ(.DI(r_4[27:27]),.CI(un32_reg0_cry_26),.S(un32_reg0_axb_27),.LO(un32_reg0_cry_27));
  XORCY un32_reg0_s_26_cZ(.LI(un32_reg0_axb_26),.CI(un32_reg0_cry_25),.O(un32_reg0_s_26));
  MUXCY_L un32_reg0_cry_26_cZ(.DI(r_4[26:26]),.CI(un32_reg0_cry_25),.S(un32_reg0_axb_26),.LO(un32_reg0_cry_26));
  XORCY un32_reg0_s_25_cZ(.LI(un32_reg0_axb_25),.CI(un32_reg0_cry_24),.O(un32_reg0_s_25));
  MUXCY_L un32_reg0_cry_25_cZ(.DI(r_4[25:25]),.CI(un32_reg0_cry_24),.S(un32_reg0_axb_25),.LO(un32_reg0_cry_25));
  XORCY un32_reg0_s_24_cZ(.LI(un32_reg0_axb_24),.CI(un32_reg0_cry_23),.O(un32_reg0_s_24));
  MUXCY_L un32_reg0_cry_24_cZ(.DI(r_4[24:24]),.CI(un32_reg0_cry_23),.S(un32_reg0_axb_24),.LO(un32_reg0_cry_24));
  XORCY un32_reg0_s_23_cZ(.LI(un32_reg0_axb_23),.CI(un32_reg0_cry_22),.O(un32_reg0_s_23));
  MUXCY_L un32_reg0_cry_23_cZ(.DI(r_4[23:23]),.CI(un32_reg0_cry_22),.S(un32_reg0_axb_23),.LO(un32_reg0_cry_23));
  XORCY un32_reg0_s_22_cZ(.LI(un32_reg0_axb_22),.CI(un32_reg0_cry_21),.O(un32_reg0_s_22));
  MUXCY_L un32_reg0_cry_22_cZ(.DI(r_4[22:22]),.CI(un32_reg0_cry_21),.S(un32_reg0_axb_22),.LO(un32_reg0_cry_22));
  XORCY un32_reg0_s_21_cZ(.LI(un32_reg0_axb_21),.CI(un32_reg0_cry_20),.O(un32_reg0_s_21));
  MUXCY_L un32_reg0_cry_21_cZ(.DI(r_4[21:21]),.CI(un32_reg0_cry_20),.S(un32_reg0_axb_21),.LO(un32_reg0_cry_21));
  XORCY un32_reg0_s_20_cZ(.LI(un32_reg0_axb_20),.CI(un32_reg0_cry_19),.O(un32_reg0_s_20));
  MUXCY_L un32_reg0_cry_20_cZ(.DI(r_4[20:20]),.CI(un32_reg0_cry_19),.S(un32_reg0_axb_20),.LO(un32_reg0_cry_20));
  XORCY un32_reg0_s_19_cZ(.LI(un32_reg0_axb_19),.CI(un32_reg0_cry_18),.O(un32_reg0_s_19));
  MUXCY_L un32_reg0_cry_19_cZ(.DI(r_4[19:19]),.CI(un32_reg0_cry_18),.S(un32_reg0_axb_19),.LO(un32_reg0_cry_19));
  XORCY un32_reg0_s_18_cZ(.LI(un32_reg0_axb_18),.CI(un32_reg0_cry_17),.O(un32_reg0_s_18));
  MUXCY_L un32_reg0_cry_18_cZ(.DI(r_4[18:18]),.CI(un32_reg0_cry_17),.S(un32_reg0_axb_18),.LO(un32_reg0_cry_18));
  XORCY un32_reg0_s_17_cZ(.LI(un32_reg0_axb_17),.CI(un32_reg0_cry_16),.O(un32_reg0_s_17));
  MUXCY_L un32_reg0_cry_17_cZ(.DI(r_4[17:17]),.CI(un32_reg0_cry_16),.S(un32_reg0_axb_17),.LO(un32_reg0_cry_17));
  XORCY un32_reg0_s_16_cZ(.LI(un32_reg0_axb_16),.CI(un32_reg0_cry_15),.O(un32_reg0_s_16));
  MUXCY_L un32_reg0_cry_16_cZ(.DI(r_4[16:16]),.CI(un32_reg0_cry_15),.S(un32_reg0_axb_16),.LO(un32_reg0_cry_16));
  XORCY un32_reg0_s_15_cZ(.LI(un32_reg0_axb_15),.CI(un32_reg0_cry_14),.O(un32_reg0_s_15));
  MUXCY_L un32_reg0_cry_15_cZ(.DI(r_4[15:15]),.CI(un32_reg0_cry_14),.S(un32_reg0_axb_15),.LO(un32_reg0_cry_15));
  XORCY un32_reg0_s_14_cZ(.LI(un32_reg0_axb_14),.CI(un32_reg0_cry_13),.O(un32_reg0_s_14));
  MUXCY_L un32_reg0_cry_14_cZ(.DI(r_4[14:14]),.CI(un32_reg0_cry_13),.S(un32_reg0_axb_14),.LO(un32_reg0_cry_14));
  XORCY un32_reg0_s_13_cZ(.LI(un32_reg0_axb_13),.CI(un32_reg0_cry_12),.O(un32_reg0_s_13));
  MUXCY_L un32_reg0_cry_13_cZ(.DI(r_4[13:13]),.CI(un32_reg0_cry_12),.S(un32_reg0_axb_13),.LO(un32_reg0_cry_13));
  XORCY un32_reg0_s_12_cZ(.LI(un32_reg0_axb_12),.CI(un32_reg0_cry_11),.O(un32_reg0_s_12));
  MUXCY_L un32_reg0_cry_12_cZ(.DI(r_4[12:12]),.CI(un32_reg0_cry_11),.S(un32_reg0_axb_12),.LO(un32_reg0_cry_12));
  XORCY un32_reg0_s_11_cZ(.LI(un32_reg0_axb_11),.CI(un32_reg0_cry_10),.O(un32_reg0_s_11));
  MUXCY_L un32_reg0_cry_11_cZ(.DI(r_4[11:11]),.CI(un32_reg0_cry_10),.S(un32_reg0_axb_11),.LO(un32_reg0_cry_11));
  XORCY un32_reg0_s_10_cZ(.LI(un32_reg0_axb_10),.CI(un32_reg0_cry_9),.O(un32_reg0_s_10));
  MUXCY_L un32_reg0_cry_10_cZ(.DI(r_4[10:10]),.CI(un32_reg0_cry_9),.S(un32_reg0_axb_10),.LO(un32_reg0_cry_10));
  XORCY un32_reg0_s_9_cZ(.LI(un32_reg0_axb_9),.CI(un32_reg0_cry_8),.O(un32_reg0_s_9));
  MUXCY_L un32_reg0_cry_9_cZ(.DI(r_4[9:9]),.CI(un32_reg0_cry_8),.S(un32_reg0_axb_9),.LO(un32_reg0_cry_9));
  XORCY un32_reg0_s_8_cZ(.LI(un32_reg0_axb_8),.CI(un32_reg0_cry_7),.O(un32_reg0_s_8));
  MUXCY_L un32_reg0_cry_8_cZ(.DI(r_4[8:8]),.CI(un32_reg0_cry_7),.S(un32_reg0_axb_8),.LO(un32_reg0_cry_8));
  XORCY un32_reg0_s_7_cZ(.LI(un32_reg0_axb_7),.CI(un32_reg0_cry_6),.O(un32_reg0_s_7));
  MUXCY_L un32_reg0_cry_7_cZ(.DI(r_4[7:7]),.CI(un32_reg0_cry_6),.S(un32_reg0_axb_7),.LO(un32_reg0_cry_7));
  XORCY un32_reg0_s_6_cZ(.LI(un32_reg0_axb_6),.CI(un32_reg0_cry_5),.O(un32_reg0_s_6));
  MUXCY_L un32_reg0_cry_6_cZ(.DI(r_4[6:6]),.CI(un32_reg0_cry_5),.S(un32_reg0_axb_6),.LO(un32_reg0_cry_6));
  XORCY un32_reg0_s_5_cZ(.LI(un32_reg0_axb_5),.CI(un32_reg0_cry_4),.O(un32_reg0_s_5));
  MUXCY_L un32_reg0_cry_5_cZ(.DI(r_4[5:5]),.CI(un32_reg0_cry_4),.S(un32_reg0_axb_5),.LO(un32_reg0_cry_5));
  XORCY un32_reg0_s_4_cZ(.LI(un32_reg0_axb_4),.CI(un32_reg0_cry_3),.O(un32_reg0_s_4));
  MUXCY_L un32_reg0_cry_4_cZ(.DI(r_4[4:4]),.CI(un32_reg0_cry_3),.S(un32_reg0_axb_4),.LO(un32_reg0_cry_4));
  XORCY un32_reg0_s_3_cZ(.LI(un32_reg0_axb_3),.CI(un32_reg0_cry_2),.O(un32_reg0_s_3));
  MUXCY_L un32_reg0_cry_3_cZ(.DI(r_4[3:3]),.CI(un32_reg0_cry_2),.S(un32_reg0_axb_3),.LO(un32_reg0_cry_3));
  XORCY un32_reg0_s_2_cZ(.LI(un32_reg0_axb_2),.CI(un32_reg0_cry_1),.O(un32_reg0_s_2));
  MUXCY_L un32_reg0_cry_2_cZ(.DI(N_28),.CI(un32_reg0_cry_1),.S(un32_reg0_axb_2),.LO(un32_reg0_cry_2));
  XORCY un32_reg0_s_1_cZ(.LI(un32_reg0_axb_1),.CI(un32_reg0_cry_0),.O(un32_reg0_s_1));
  MUXCY_L un32_reg0_cry_1_cZ(.DI(r_4[1:1]),.CI(un32_reg0_cry_0),.S(un32_reg0_axb_1),.LO(un32_reg0_cry_1));
  MUXCY_L un32_reg0_cry_0_cZ(.DI(r_4[0:0]),.CI(VCC),.S(N_1035),.LO(un32_reg0_cry_0));
  XORCY un11_reg0_s_29_cZ(.LI(un11_reg0_axb_29),.CI(un11_reg0_cry_28),.O(un11_reg0_s_29));
  XORCY un11_reg0_s_28_cZ(.LI(un11_reg0_axb_28),.CI(un11_reg0_cry_27),.O(un11_reg0_s_28));
  MUXCY_L un11_reg0_cry_28_cZ(.DI(m_2[28:28]),.CI(un11_reg0_cry_27),.S(un11_reg0_axb_28),.LO(un11_reg0_cry_28));
  XORCY un11_reg0_s_27_cZ(.LI(un11_reg0_axb_27),.CI(un11_reg0_cry_26),.O(un11_reg0_s_27));
  MUXCY_L un11_reg0_cry_27_cZ(.DI(m_2[27:27]),.CI(un11_reg0_cry_26),.S(un11_reg0_axb_27),.LO(un11_reg0_cry_27));
  XORCY un11_reg0_s_26_cZ(.LI(un11_reg0_axb_26),.CI(un11_reg0_cry_25),.O(un11_reg0_s_26));
  MUXCY_L un11_reg0_cry_26_cZ(.DI(m_2[26:26]),.CI(un11_reg0_cry_25),.S(un11_reg0_axb_26),.LO(un11_reg0_cry_26));
  XORCY un11_reg0_s_25_cZ(.LI(un11_reg0_axb_25),.CI(un11_reg0_cry_24),.O(un11_reg0_s_25));
  MUXCY_L un11_reg0_cry_25_cZ(.DI(m_2[25:25]),.CI(un11_reg0_cry_24),.S(un11_reg0_axb_25),.LO(un11_reg0_cry_25));
  XORCY un11_reg0_s_24_cZ(.LI(un11_reg0_axb_24),.CI(un11_reg0_cry_23),.O(un11_reg0_s_24));
  MUXCY_L un11_reg0_cry_24_cZ(.DI(m_2[24:24]),.CI(un11_reg0_cry_23),.S(un11_reg0_axb_24),.LO(un11_reg0_cry_24));
  XORCY un11_reg0_s_23_cZ(.LI(un11_reg0_axb_23),.CI(un11_reg0_cry_22),.O(un11_reg0_s_23));
  MUXCY_L un11_reg0_cry_23_cZ(.DI(m_2[23:23]),.CI(un11_reg0_cry_22),.S(un11_reg0_axb_23),.LO(un11_reg0_cry_23));
  XORCY un11_reg0_s_22_cZ(.LI(un11_reg0_axb_22),.CI(un11_reg0_cry_21),.O(un11_reg0_s_22));
  MUXCY_L un11_reg0_cry_22_cZ(.DI(m_2[22:22]),.CI(un11_reg0_cry_21),.S(un11_reg0_axb_22),.LO(un11_reg0_cry_22));
  XORCY un11_reg0_s_21_cZ(.LI(un11_reg0_axb_21),.CI(un11_reg0_cry_20),.O(un11_reg0_s_21));
  MUXCY_L un11_reg0_cry_21_cZ(.DI(m_2[21:21]),.CI(un11_reg0_cry_20),.S(un11_reg0_axb_21),.LO(un11_reg0_cry_21));
  XORCY un11_reg0_s_20_cZ(.LI(un11_reg0_axb_20),.CI(un11_reg0_cry_19),.O(un11_reg0_s_20));
  MUXCY_L un11_reg0_cry_20_cZ(.DI(m_2[20:20]),.CI(un11_reg0_cry_19),.S(un11_reg0_axb_20),.LO(un11_reg0_cry_20));
  XORCY un11_reg0_s_19_cZ(.LI(un11_reg0_axb_19),.CI(un11_reg0_cry_18),.O(un11_reg0_s_19));
  MUXCY_L un11_reg0_cry_19_cZ(.DI(r_4[19:19]),.CI(un11_reg0_cry_18),.S(un11_reg0_axb_19),.LO(un11_reg0_cry_19));
  XORCY un11_reg0_s_18_cZ(.LI(un11_reg0_axb_18),.CI(un11_reg0_cry_17),.O(un11_reg0_s_18));
  MUXCY_L un11_reg0_cry_18_cZ(.DI(r_4[18:18]),.CI(un11_reg0_cry_17),.S(un11_reg0_axb_18),.LO(un11_reg0_cry_18));
  XORCY un11_reg0_s_17_cZ(.LI(un11_reg0_axb_17),.CI(un11_reg0_cry_16),.O(un11_reg0_s_17));
  MUXCY_L un11_reg0_cry_17_cZ(.DI(r_4[17:17]),.CI(un11_reg0_cry_16),.S(un11_reg0_axb_17),.LO(un11_reg0_cry_17));
  XORCY un11_reg0_s_16_cZ(.LI(un11_reg0_axb_16),.CI(un11_reg0_cry_15),.O(un11_reg0_s_16));
  MUXCY_L un11_reg0_cry_16_cZ(.DI(r_4[16:16]),.CI(un11_reg0_cry_15),.S(un11_reg0_axb_16),.LO(un11_reg0_cry_16));
  XORCY un11_reg0_s_15_cZ(.LI(un11_reg0_axb_15),.CI(un11_reg0_cry_14),.O(un11_reg0_s_15));
  MUXCY_L un11_reg0_cry_15_cZ(.DI(r_4[15:15]),.CI(un11_reg0_cry_14),.S(un11_reg0_axb_15),.LO(un11_reg0_cry_15));
  XORCY un11_reg0_s_14_cZ(.LI(un11_reg0_axb_14),.CI(un11_reg0_cry_13),.O(un11_reg0_s_14));
  MUXCY_L un11_reg0_cry_14_cZ(.DI(r_4[14:14]),.CI(un11_reg0_cry_13),.S(un11_reg0_axb_14),.LO(un11_reg0_cry_14));
  XORCY un11_reg0_s_13_cZ(.LI(un11_reg0_axb_13),.CI(un11_reg0_cry_12),.O(un11_reg0_s_13));
  MUXCY_L un11_reg0_cry_13_cZ(.DI(r_4[13:13]),.CI(un11_reg0_cry_12),.S(un11_reg0_axb_13),.LO(un11_reg0_cry_13));
  XORCY un11_reg0_s_12_cZ(.LI(un11_reg0_axb_12),.CI(un11_reg0_cry_11),.O(un11_reg0_s_12));
  MUXCY_L un11_reg0_cry_12_cZ(.DI(r_4[12:12]),.CI(un11_reg0_cry_11),.S(un11_reg0_axb_12),.LO(un11_reg0_cry_12));
  XORCY un11_reg0_s_11_cZ(.LI(un11_reg0_axb_11),.CI(un11_reg0_cry_10),.O(un11_reg0_s_11));
  MUXCY_L un11_reg0_cry_11_cZ(.DI(r_4[11:11]),.CI(un11_reg0_cry_10),.S(un11_reg0_axb_11),.LO(un11_reg0_cry_11));
  XORCY un11_reg0_s_10_cZ(.LI(un11_reg0_axb_10),.CI(un11_reg0_cry_9),.O(un11_reg0_s_10));
  MUXCY_L un11_reg0_cry_10_cZ(.DI(r_4[10:10]),.CI(un11_reg0_cry_9),.S(un11_reg0_axb_10),.LO(un11_reg0_cry_10));
  XORCY un11_reg0_s_9_cZ(.LI(un11_reg0_axb_9),.CI(un11_reg0_cry_8),.O(un11_reg0_s_9));
  MUXCY_L un11_reg0_cry_9_cZ(.DI(r_4[9:9]),.CI(un11_reg0_cry_8),.S(un11_reg0_axb_9),.LO(un11_reg0_cry_9));
  XORCY un11_reg0_s_8_cZ(.LI(un11_reg0_axb_8),.CI(un11_reg0_cry_7),.O(un11_reg0_s_8));
  MUXCY_L un11_reg0_cry_8_cZ(.DI(r_4[8:8]),.CI(un11_reg0_cry_7),.S(un11_reg0_axb_8),.LO(un11_reg0_cry_8));
  XORCY un11_reg0_s_7_cZ(.LI(un11_reg0_axb_7),.CI(un11_reg0_cry_6),.O(un11_reg0_s_7));
  MUXCY_L un11_reg0_cry_7_cZ(.DI(r_4[7:7]),.CI(un11_reg0_cry_6),.S(un11_reg0_axb_7),.LO(un11_reg0_cry_7));
  XORCY un11_reg0_s_6_cZ(.LI(un11_reg0_axb_6),.CI(un11_reg0_cry_5),.O(un11_reg0_s_6));
  MUXCY_L un11_reg0_cry_6_cZ(.DI(r_4[6:6]),.CI(un11_reg0_cry_5),.S(un11_reg0_axb_6),.LO(un11_reg0_cry_6));
  XORCY un11_reg0_s_5_cZ(.LI(un11_reg0_axb_5),.CI(un11_reg0_cry_4),.O(un11_reg0_s_5));
  MUXCY_L un11_reg0_cry_5_cZ(.DI(r_4[5:5]),.CI(un11_reg0_cry_4),.S(un11_reg0_axb_5),.LO(un11_reg0_cry_5));
  XORCY un11_reg0_s_4_cZ(.LI(un11_reg0_axb_4),.CI(un11_reg0_cry_3),.O(un11_reg0_s_4));
  MUXCY_L un11_reg0_cry_4_cZ(.DI(r_4[4:4]),.CI(un11_reg0_cry_3),.S(un11_reg0_axb_4),.LO(un11_reg0_cry_4));
  XORCY un11_reg0_s_3_cZ(.LI(un11_reg0_axb_3),.CI(un11_reg0_cry_2),.O(un11_reg0_s_3));
  MUXCY_L un11_reg0_cry_3_cZ(.DI(r_4[3:3]),.CI(un11_reg0_cry_2),.S(un11_reg0_axb_3),.LO(un11_reg0_cry_3));
  XORCY un11_reg0_s_2_cZ(.LI(un11_reg0_axb_2),.CI(un11_reg0_cry_1),.O(un11_reg0_s_2));
  MUXCY_L un11_reg0_cry_2_cZ(.DI(N_28),.CI(un11_reg0_cry_1),.S(un11_reg0_axb_2),.LO(un11_reg0_cry_2));
  XORCY un11_reg0_s_1_cZ(.LI(un11_reg0_axb_1),.CI(un11_reg0_cry_0),.O(un11_reg0_s_1));
  MUXCY_L un11_reg0_cry_1_cZ(.DI(r_4[1:1]),.CI(un11_reg0_cry_0),.S(un11_reg0_axb_1),.LO(un11_reg0_cry_1));
  MUXCY_L un11_reg0_cry_0_cZ(.DI(r_4[0:0]),.CI(GND),.S(un11_reg0_axb_0),.LO(un11_reg0_cry_0));
  XORCY un3_t_s_31_cZ(.LI(un3_t_axb_31),.CI(un3_t_cry_30),.O(un3_t_s_31));
  XORCY un3_t_s_30_cZ(.LI(un3_t_axb_30),.CI(un3_t_cry_29),.O(un3_t_s_30));
  MUXCY_L un3_t_cry_30_cZ(.DI(GND),.CI(un3_t_cry_29),.S(un3_t_axb_30),.LO(un3_t_cry_30));
  XORCY un3_t_s_29_cZ(.LI(un3_t_axb_29),.CI(un3_t_cry_28),.O(un3_t_s_29));
  MUXCY_L un3_t_cry_29_cZ(.DI(GND),.CI(un3_t_cry_28),.S(un3_t_axb_29),.LO(un3_t_cry_29));
  XORCY un3_t_s_28_cZ(.LI(un3_t_axb_28),.CI(un3_t_cry_27),.O(un3_t_s_28));
  MUXCY_L un3_t_cry_28_cZ(.DI(GND),.CI(un3_t_cry_27),.S(un3_t_axb_28),.LO(un3_t_cry_28));
  XORCY un3_t_s_27_cZ(.LI(un3_t_axb_27),.CI(un3_t_cry_26),.O(un3_t_s_27));
  MUXCY_L un3_t_cry_27_cZ(.DI(GND),.CI(un3_t_cry_26),.S(un3_t_axb_27),.LO(un3_t_cry_27));
  XORCY un3_t_s_26_cZ(.LI(un3_t_axb_26),.CI(un3_t_cry_25),.O(un3_t_s_26));
  MUXCY_L un3_t_cry_26_cZ(.DI(GND),.CI(un3_t_cry_25),.S(un3_t_axb_26),.LO(un3_t_cry_26));
  XORCY un3_t_s_25_cZ(.LI(un3_t_axb_25),.CI(un3_t_cry_24),.O(un3_t_s_25));
  MUXCY_L un3_t_cry_25_cZ(.DI(GND),.CI(un3_t_cry_24),.S(un3_t_axb_25),.LO(un3_t_cry_25));
  XORCY un3_t_s_24_cZ(.LI(un3_t_axb_24),.CI(un3_t_cry_23),.O(un3_t_s_24));
  MUXCY_L un3_t_cry_24_cZ(.DI(GND),.CI(un3_t_cry_23),.S(un3_t_axb_24),.LO(un3_t_cry_24));
  XORCY un3_t_s_23_cZ(.LI(un3_t_axb_23),.CI(un3_t_cry_22),.O(un3_t_s_23));
  MUXCY_L un3_t_cry_23_cZ(.DI(GND),.CI(un3_t_cry_22),.S(un3_t_axb_23),.LO(un3_t_cry_23));
  XORCY un3_t_s_22_cZ(.LI(un3_t_axb_22),.CI(un3_t_cry_21),.O(un3_t_s_22));
  MUXCY_L un3_t_cry_22_cZ(.DI(GND),.CI(un3_t_cry_21),.S(un3_t_axb_22),.LO(un3_t_cry_22));
  XORCY un3_t_s_21_cZ(.LI(un3_t_axb_21),.CI(un3_t_cry_20),.O(un3_t_s_21));
  MUXCY_L un3_t_cry_21_cZ(.DI(GND),.CI(un3_t_cry_20),.S(un3_t_axb_21),.LO(un3_t_cry_21));
  XORCY un3_t_s_20_cZ(.LI(un3_t_axb_20),.CI(un3_t_cry_19),.O(un3_t_s_20));
  MUXCY_L un3_t_cry_20_cZ(.DI(GND),.CI(un3_t_cry_19),.S(un3_t_axb_20),.LO(un3_t_cry_20));
  XORCY un3_t_s_19_cZ(.LI(un3_t_axb_19),.CI(un3_t_cry_18),.O(un3_t_s_19));
  MUXCY_L un3_t_cry_19_cZ(.DI(GND),.CI(un3_t_cry_18),.S(un3_t_axb_19),.LO(un3_t_cry_19));
  XORCY un3_t_s_18_cZ(.LI(un3_t_axb_18),.CI(un3_t_cry_17),.O(un3_t_s_18));
  MUXCY_L un3_t_cry_18_cZ(.DI(GND),.CI(un3_t_cry_17),.S(un3_t_axb_18),.LO(un3_t_cry_18));
  XORCY un3_t_s_17_cZ(.LI(un3_t_axb_17),.CI(un3_t_cry_16),.O(un3_t_s_17));
  MUXCY_L un3_t_cry_17_cZ(.DI(GND),.CI(un3_t_cry_16),.S(un3_t_axb_17),.LO(un3_t_cry_17));
  XORCY un3_t_s_16_cZ(.LI(un3_t_axb_16),.CI(un3_t_cry_15),.O(un3_t_s_16));
  MUXCY_L un3_t_cry_16_cZ(.DI(GND),.CI(un3_t_cry_15),.S(un3_t_axb_16),.LO(un3_t_cry_16));
  XORCY un3_t_s_15_cZ(.LI(un3_t_axb_15),.CI(un3_t_cry_14),.O(un3_t_s_15));
  MUXCY_L un3_t_cry_15_cZ(.DI(GND),.CI(un3_t_cry_14),.S(un3_t_axb_15),.LO(un3_t_cry_15));
  XORCY un3_t_s_14_cZ(.LI(un3_t_axb_14),.CI(un3_t_cry_13),.O(un3_t_s_14));
  MUXCY_L un3_t_cry_14_cZ(.DI(GND),.CI(un3_t_cry_13),.S(un3_t_axb_14),.LO(un3_t_cry_14));
  XORCY un3_t_s_13_cZ(.LI(un3_t_axb_13),.CI(un3_t_cry_12),.O(un3_t_s_13));
  MUXCY_L un3_t_cry_13_cZ(.DI(GND),.CI(un3_t_cry_12),.S(un3_t_axb_13),.LO(un3_t_cry_13));
  XORCY un3_t_s_12_cZ(.LI(un3_t_axb_12),.CI(un3_t_cry_11),.O(un3_t_s_12));
  MUXCY_L un3_t_cry_12_cZ(.DI(GND),.CI(un3_t_cry_11),.S(un3_t_axb_12),.LO(un3_t_cry_12));
  XORCY un3_t_s_11_cZ(.LI(un3_t_axb_11),.CI(un3_t_cry_10),.O(un3_t_s_11));
  MUXCY_L un3_t_cry_11_cZ(.DI(GND),.CI(un3_t_cry_10),.S(un3_t_axb_11),.LO(un3_t_cry_11));
  XORCY un3_t_s_10_cZ(.LI(un3_t_axb_10),.CI(un3_t_cry_9),.O(un3_t_s_10));
  MUXCY_L un3_t_cry_10_cZ(.DI(GND),.CI(un3_t_cry_9),.S(un3_t_axb_10),.LO(un3_t_cry_10));
  XORCY un3_t_s_9_cZ(.LI(un3_t_axb_9),.CI(un3_t_cry_8),.O(un3_t_s_9));
  MUXCY_L un3_t_cry_9_cZ(.DI(GND),.CI(un3_t_cry_8),.S(un3_t_axb_9),.LO(un3_t_cry_9));
  XORCY un3_t_s_8_cZ(.LI(un3_t_axb_8),.CI(un3_t_cry_7),.O(un3_t_s_8));
  MUXCY_L un3_t_cry_8_cZ(.DI(GND),.CI(un3_t_cry_7),.S(un3_t_axb_8),.LO(un3_t_cry_8));
  XORCY un3_t_s_7_cZ(.LI(un3_t_axb_7),.CI(un3_t_cry_6),.O(un3_t_s_7));
  MUXCY_L un3_t_cry_7_cZ(.DI(GND),.CI(un3_t_cry_6),.S(un3_t_axb_7),.LO(un3_t_cry_7));
  XORCY un3_t_s_6_cZ(.LI(un3_t_axb_6),.CI(un3_t_cry_5),.O(un3_t_s_6));
  MUXCY_L un3_t_cry_6_cZ(.DI(GND),.CI(un3_t_cry_5),.S(un3_t_axb_6),.LO(un3_t_cry_6));
  XORCY un3_t_s_5_cZ(.LI(un3_t_axb_5),.CI(un3_t_cry_4),.O(un3_t_s_5));
  MUXCY_L un3_t_cry_5_cZ(.DI(GND),.CI(un3_t_cry_4),.S(un3_t_axb_5),.LO(un3_t_cry_5));
  XORCY un3_t_s_4_cZ(.LI(un3_t_axb_4),.CI(un3_t_cry_3),.O(un3_t_s_4));
  MUXCY_L un3_t_cry_4_cZ(.DI(GND),.CI(un3_t_cry_3),.S(un3_t_axb_4),.LO(un3_t_cry_4));
  XORCY un3_t_s_3_cZ(.LI(un3_t_axb_3),.CI(un3_t_cry_2),.O(un3_t_s_3));
  MUXCY_L un3_t_cry_3_cZ(.DI(GND),.CI(un3_t_cry_2),.S(un3_t_axb_3),.LO(un3_t_cry_3));
  XORCY un3_t_s_2_cZ(.LI(un3_t_axb_2),.CI(un3_t_cry_1),.O(un3_t_s_2));
  MUXCY_L un3_t_cry_2_cZ(.DI(GND),.CI(un3_t_cry_1),.S(un3_t_axb_2),.LO(un3_t_cry_2));
  XORCY un3_t_s_1_cZ(.LI(un3_t_axb_1),.CI(un3_t_cry_0),.O(un3_t_s_1));
  MUXCY_L un3_t_cry_1_cZ(.DI(GND),.CI(un3_t_cry_0),.S(un3_t_axb_1),.LO(un3_t_cry_1));
  MUXCY_L un3_t_cry_0_cZ(.DI(GND),.CI(un3_t_cry_0_cy),.S(un3_t_axb_0),.LO(un3_t_cry_0));
  XORCY reg3_1_1_s_31(.LI(reg3_1_1_axb_31),.CI(reg3_1_1_cry_30),.O(reg3_1_1[31:31]));
  XORCY reg3_1_1_s_30(.LI(reg3_1_1_axb_30),.CI(reg3_1_1_cry_29),.O(reg3_1_1[30:30]));
  MUXCY_L reg3_1_1_cry_30_cZ(.DI(GND),.CI(reg3_1_1_cry_29),.S(reg3_1_1_axb_30),.LO(reg3_1_1_cry_30));
  XORCY reg3_1_1_s_29(.LI(reg3_1_1_axb_29),.CI(reg3_1_1_cry_28),.O(reg3_1_1[29:29]));
  MUXCY_L reg3_1_1_cry_29_cZ(.DI(GND),.CI(reg3_1_1_cry_28),.S(reg3_1_1_axb_29),.LO(reg3_1_1_cry_29));
  XORCY reg3_1_1_s_28(.LI(reg3_1_1_axb_28),.CI(reg3_1_1_cry_27),.O(reg3_1_1[28:28]));
  MUXCY_L reg3_1_1_cry_28_cZ(.DI(GND),.CI(reg3_1_1_cry_27),.S(reg3_1_1_axb_28),.LO(reg3_1_1_cry_28));
  XORCY reg3_1_1_s_27(.LI(reg3_1_1_axb_27),.CI(reg3_1_1_cry_26),.O(reg3_1_1[27:27]));
  MUXCY_L reg3_1_1_cry_27_cZ(.DI(GND),.CI(reg3_1_1_cry_26),.S(reg3_1_1_axb_27),.LO(reg3_1_1_cry_27));
  XORCY reg3_1_1_s_26(.LI(reg3_1_1_axb_26),.CI(reg3_1_1_cry_25),.O(reg3_1_1[26:26]));
  MUXCY_L reg3_1_1_cry_26_cZ(.DI(GND),.CI(reg3_1_1_cry_25),.S(reg3_1_1_axb_26),.LO(reg3_1_1_cry_26));
  XORCY reg3_1_1_s_25(.LI(reg3_1_1_axb_25),.CI(reg3_1_1_cry_24),.O(reg3_1_1[25:25]));
  MUXCY_L reg3_1_1_cry_25_cZ(.DI(GND),.CI(reg3_1_1_cry_24),.S(reg3_1_1_axb_25),.LO(reg3_1_1_cry_25));
  XORCY reg3_1_1_s_24(.LI(reg3_1_1_axb_24),.CI(reg3_1_1_cry_23),.O(reg3_1_1[24:24]));
  MUXCY_L reg3_1_1_cry_24_cZ(.DI(GND),.CI(reg3_1_1_cry_23),.S(reg3_1_1_axb_24),.LO(reg3_1_1_cry_24));
  XORCY reg3_1_1_s_23(.LI(reg3_1_1_axb_23),.CI(reg3_1_1_cry_22),.O(reg3_1_1[23:23]));
  MUXCY_L reg3_1_1_cry_23_cZ(.DI(GND),.CI(reg3_1_1_cry_22),.S(reg3_1_1_axb_23),.LO(reg3_1_1_cry_23));
  XORCY reg3_1_1_s_22(.LI(reg3_1_1_axb_22),.CI(reg3_1_1_cry_21),.O(reg3_1_1[22:22]));
  MUXCY_L reg3_1_1_cry_22_cZ(.DI(GND),.CI(reg3_1_1_cry_21),.S(reg3_1_1_axb_22),.LO(reg3_1_1_cry_22));
  XORCY reg3_1_1_s_21(.LI(reg3_1_1_axb_21),.CI(reg3_1_1_cry_20),.O(reg3_1_1[21:21]));
  MUXCY_L reg3_1_1_cry_21_cZ(.DI(GND),.CI(reg3_1_1_cry_20),.S(reg3_1_1_axb_21),.LO(reg3_1_1_cry_21));
  XORCY reg3_1_1_s_20(.LI(reg3_1_1_axb_20),.CI(reg3_1_1_cry_19),.O(reg3_1_1[20:20]));
  MUXCY_L reg3_1_1_cry_20_cZ(.DI(GND),.CI(reg3_1_1_cry_19),.S(reg3_1_1_axb_20),.LO(reg3_1_1_cry_20));
  XORCY reg3_1_1_s_19(.LI(reg3_1_1_axb_19),.CI(reg3_1_1_cry_18),.O(reg3_1_1[19:19]));
  MUXCY_L reg3_1_1_cry_19_cZ(.DI(GND),.CI(reg3_1_1_cry_18),.S(reg3_1_1_axb_19),.LO(reg3_1_1_cry_19));
  XORCY reg3_1_1_s_18(.LI(reg3_1_1_axb_18),.CI(reg3_1_1_cry_17),.O(reg3_1_1[18:18]));
  MUXCY_L reg3_1_1_cry_18_cZ(.DI(GND),.CI(reg3_1_1_cry_17),.S(reg3_1_1_axb_18),.LO(reg3_1_1_cry_18));
  XORCY reg3_1_1_s_17(.LI(reg3_1_1_axb_17),.CI(reg3_1_1_cry_16),.O(reg3_1_1[17:17]));
  MUXCY_L reg3_1_1_cry_17_cZ(.DI(GND),.CI(reg3_1_1_cry_16),.S(reg3_1_1_axb_17),.LO(reg3_1_1_cry_17));
  XORCY reg3_1_1_s_16(.LI(reg3_1_1_axb_16),.CI(reg3_1_1_cry_15),.O(reg3_1_1[16:16]));
  MUXCY_L reg3_1_1_cry_16_cZ(.DI(GND),.CI(reg3_1_1_cry_15),.S(reg3_1_1_axb_16),.LO(reg3_1_1_cry_16));
  XORCY reg3_1_1_s_15(.LI(reg3_1_1_axb_15),.CI(reg3_1_1_cry_14),.O(reg3_1_1[15:15]));
  MUXCY_L reg3_1_1_cry_15_cZ(.DI(GND),.CI(reg3_1_1_cry_14),.S(reg3_1_1_axb_15),.LO(reg3_1_1_cry_15));
  XORCY reg3_1_1_s_14(.LI(reg3_1_1_axb_14),.CI(reg3_1_1_cry_13),.O(reg3_1_1[14:14]));
  MUXCY_L reg3_1_1_cry_14_cZ(.DI(GND),.CI(reg3_1_1_cry_13),.S(reg3_1_1_axb_14),.LO(reg3_1_1_cry_14));
  XORCY reg3_1_1_s_13(.LI(reg3_1_1_axb_13),.CI(reg3_1_1_cry_12),.O(reg3_1_1[13:13]));
  MUXCY_L reg3_1_1_cry_13_cZ(.DI(GND),.CI(reg3_1_1_cry_12),.S(reg3_1_1_axb_13),.LO(reg3_1_1_cry_13));
  XORCY reg3_1_1_s_12(.LI(reg3_1_1_axb_12),.CI(reg3_1_1_cry_11),.O(reg3_1_1[12:12]));
  MUXCY_L reg3_1_1_cry_12_cZ(.DI(GND),.CI(reg3_1_1_cry_11),.S(reg3_1_1_axb_12),.LO(reg3_1_1_cry_12));
  XORCY reg3_1_1_s_11(.LI(reg3_1_1_axb_11),.CI(reg3_1_1_cry_10),.O(reg3_1_1[11:11]));
  MUXCY_L reg3_1_1_cry_11_cZ(.DI(GND),.CI(reg3_1_1_cry_10),.S(reg3_1_1_axb_11),.LO(reg3_1_1_cry_11));
  XORCY reg3_1_1_s_10(.LI(reg3_1_1_axb_10),.CI(reg3_1_1_cry_9),.O(reg3_1_1[10:10]));
  MUXCY_L reg3_1_1_cry_10_cZ(.DI(GND),.CI(reg3_1_1_cry_9),.S(reg3_1_1_axb_10),.LO(reg3_1_1_cry_10));
  XORCY reg3_1_1_s_9(.LI(reg3_1_1_axb_9),.CI(reg3_1_1_cry_8),.O(reg3_1_1[9:9]));
  MUXCY_L reg3_1_1_cry_9_cZ(.DI(GND),.CI(reg3_1_1_cry_8),.S(reg3_1_1_axb_9),.LO(reg3_1_1_cry_9));
  XORCY reg3_1_1_s_8(.LI(reg3_1_1_axb_8),.CI(reg3_1_1_cry_7),.O(reg3_1_1[8:8]));
  MUXCY_L reg3_1_1_cry_8_cZ(.DI(GND),.CI(reg3_1_1_cry_7),.S(reg3_1_1_axb_8),.LO(reg3_1_1_cry_8));
  XORCY reg3_1_1_s_7(.LI(reg3_1_1_axb_7),.CI(reg3_1_1_cry_6),.O(reg3_1_1[7:7]));
  MUXCY_L reg3_1_1_cry_7_cZ(.DI(GND),.CI(reg3_1_1_cry_6),.S(reg3_1_1_axb_7),.LO(reg3_1_1_cry_7));
  XORCY reg3_1_1_s_6(.LI(reg3_1_1_axb_6),.CI(reg3_1_1_cry_5),.O(reg3_1_1[6:6]));
  MUXCY_L reg3_1_1_cry_6_cZ(.DI(GND),.CI(reg3_1_1_cry_5),.S(reg3_1_1_axb_6),.LO(reg3_1_1_cry_6));
  XORCY reg3_1_1_s_5(.LI(reg3_1_1_axb_5),.CI(reg3_1_1_cry_4),.O(reg3_1_1[5:5]));
  MUXCY_L reg3_1_1_cry_5_cZ(.DI(GND),.CI(reg3_1_1_cry_4),.S(reg3_1_1_axb_5),.LO(reg3_1_1_cry_5));
  XORCY reg3_1_1_s_4(.LI(reg3_1_1_axb_4),.CI(reg3_1_1_cry_3),.O(reg3_1_1[4:4]));
  MUXCY_L reg3_1_1_cry_4_cZ(.DI(GND),.CI(reg3_1_1_cry_3),.S(reg3_1_1_axb_4),.LO(reg3_1_1_cry_4));
  XORCY reg3_1_1_s_3(.LI(reg3_1_1_axb_3),.CI(reg3_1_1_cry_2),.O(reg3_1_1[3:3]));
  MUXCY_L reg3_1_1_cry_3_cZ(.DI(GND),.CI(reg3_1_1_cry_2),.S(reg3_1_1_axb_3),.LO(reg3_1_1_cry_3));
  XORCY reg3_1_1_s_2(.LI(reg3_1_1_axb_2),.CI(reg3_1_1_cry_1),.O(reg3_1_1[2:2]));
  MUXCY_L reg3_1_1_cry_2_cZ(.DI(GND),.CI(reg3_1_1_cry_1),.S(reg3_1_1_axb_2),.LO(reg3_1_1_cry_2));
  XORCY reg3_1_1_s_1(.LI(reg3_1_1_axb_1),.CI(reg3_1_1_cry_0),.O(reg3_1_1[1:1]));
  MUXCY_L reg3_1_1_cry_1_cZ(.DI(GND),.CI(reg3_1_1_cry_0),.S(reg3_1_1_axb_1),.LO(reg3_1_1_cry_1));
  MUXCY_L reg3_1_1_cry_0_cZ(.DI(GND),.CI(VCC),.S(reg3_1_1_axb_0),.LO(reg3_1_1_cry_0));
  XORCY inf_abs0_2_s_30(.LI(inf_abs0_2_axb_30),.CI(inf_abs0_2_cry_29),.O(inf_abs0_2[30:30]));
  MUXCY inf_abs0_2_cry_30(.DI(GND),.CI(inf_abs0_2_cry_29),.S(inf_abs0_2_axb_30),.O(inf_abs0_2_0[31:31]));
  XORCY inf_abs0_2_s_29(.LI(inf_abs0_2_axb_29),.CI(inf_abs0_2_cry_28),.O(inf_abs0_2[29:29]));
  XORCY inf_abs0_2_s_28(.LI(inf_abs0_2_axb_28),.CI(inf_abs0_2_cry_27),.O(inf_abs0_2[28:28]));
  MUXCY_L inf_abs0_2_cry_28_cZ(.DI(GND),.CI(inf_abs0_2_cry_27),.S(inf_abs0_2_axb_28),.LO(inf_abs0_2_cry_28));
  XORCY inf_abs0_2_s_27(.LI(inf_abs0_2_axb_27),.CI(inf_abs0_2_cry_26),.O(inf_abs0_2[27:27]));
  MUXCY_L inf_abs0_2_cry_27_cZ(.DI(GND),.CI(inf_abs0_2_cry_26),.S(inf_abs0_2_axb_27),.LO(inf_abs0_2_cry_27));
  XORCY inf_abs0_2_s_26(.LI(inf_abs0_2_axb_26),.CI(inf_abs0_2_cry_25),.O(inf_abs0_2[26:26]));
  MUXCY_L inf_abs0_2_cry_26_cZ(.DI(GND),.CI(inf_abs0_2_cry_25),.S(inf_abs0_2_axb_26),.LO(inf_abs0_2_cry_26));
  XORCY inf_abs0_2_s_25(.LI(inf_abs0_2_axb_25),.CI(inf_abs0_2_cry_24),.O(inf_abs0_2[25:25]));
  MUXCY_L inf_abs0_2_cry_25_cZ(.DI(GND),.CI(inf_abs0_2_cry_24),.S(inf_abs0_2_axb_25),.LO(inf_abs0_2_cry_25));
  XORCY inf_abs0_2_s_24(.LI(inf_abs0_2_axb_24),.CI(inf_abs0_2_cry_23),.O(inf_abs0_2[24:24]));
  MUXCY_L inf_abs0_2_cry_24_cZ(.DI(GND),.CI(inf_abs0_2_cry_23),.S(inf_abs0_2_axb_24),.LO(inf_abs0_2_cry_24));
  XORCY inf_abs0_2_s_23(.LI(inf_abs0_2_axb_23),.CI(inf_abs0_2_cry_22),.O(inf_abs0_2[23:23]));
  MUXCY_L inf_abs0_2_cry_23_cZ(.DI(GND),.CI(inf_abs0_2_cry_22),.S(inf_abs0_2_axb_23),.LO(inf_abs0_2_cry_23));
  XORCY inf_abs0_2_s_22(.LI(inf_abs0_2_axb_22),.CI(inf_abs0_2_cry_21),.O(inf_abs0_2[22:22]));
  MUXCY_L inf_abs0_2_cry_22_cZ(.DI(GND),.CI(inf_abs0_2_cry_21),.S(inf_abs0_2_axb_22),.LO(inf_abs0_2_cry_22));
  XORCY inf_abs0_2_s_21(.LI(inf_abs0_2_axb_21),.CI(inf_abs0_2_cry_20),.O(inf_abs0_2[21:21]));
  MUXCY_L inf_abs0_2_cry_21_cZ(.DI(GND),.CI(inf_abs0_2_cry_20),.S(inf_abs0_2_axb_21),.LO(inf_abs0_2_cry_21));
  XORCY inf_abs0_2_s_20(.LI(inf_abs0_2_axb_20),.CI(inf_abs0_2_cry_19),.O(inf_abs0_2[20:20]));
  MUXCY_L inf_abs0_2_cry_20_cZ(.DI(GND),.CI(inf_abs0_2_cry_19),.S(inf_abs0_2_axb_20),.LO(inf_abs0_2_cry_20));
  XORCY inf_abs0_2_s_19(.LI(inf_abs0_2_axb_19),.CI(inf_abs0_2_cry_18),.O(inf_abs0_2[19:19]));
  MUXCY_L inf_abs0_2_cry_19_cZ(.DI(GND),.CI(inf_abs0_2_cry_18),.S(inf_abs0_2_axb_19),.LO(inf_abs0_2_cry_19));
  XORCY inf_abs0_2_s_18(.LI(inf_abs0_2_axb_18),.CI(inf_abs0_2_cry_17),.O(inf_abs0_2[18:18]));
  MUXCY_L inf_abs0_2_cry_18_cZ(.DI(GND),.CI(inf_abs0_2_cry_17),.S(inf_abs0_2_axb_18),.LO(inf_abs0_2_cry_18));
  XORCY inf_abs0_2_s_17(.LI(inf_abs0_2_axb_17),.CI(inf_abs0_2_cry_16),.O(inf_abs0_2[17:17]));
  MUXCY_L inf_abs0_2_cry_17_cZ(.DI(GND),.CI(inf_abs0_2_cry_16),.S(inf_abs0_2_axb_17),.LO(inf_abs0_2_cry_17));
  XORCY inf_abs0_2_s_16(.LI(inf_abs0_2_axb_16),.CI(inf_abs0_2_cry_15),.O(inf_abs0_2[16:16]));
  MUXCY_L inf_abs0_2_cry_16_cZ(.DI(GND),.CI(inf_abs0_2_cry_15),.S(inf_abs0_2_axb_16),.LO(inf_abs0_2_cry_16));
  XORCY inf_abs0_2_s_15(.LI(inf_abs0_2_axb_15),.CI(inf_abs0_2_cry_14),.O(inf_abs0_2[15:15]));
  MUXCY_L inf_abs0_2_cry_15_cZ(.DI(GND),.CI(inf_abs0_2_cry_14),.S(inf_abs0_2_axb_15),.LO(inf_abs0_2_cry_15));
  XORCY inf_abs0_2_s_14(.LI(inf_abs0_2_axb_14),.CI(inf_abs0_2_cry_13),.O(inf_abs0_2[14:14]));
  MUXCY_L inf_abs0_2_cry_14_cZ(.DI(GND),.CI(inf_abs0_2_cry_13),.S(inf_abs0_2_axb_14),.LO(inf_abs0_2_cry_14));
  XORCY inf_abs0_2_s_13(.LI(inf_abs0_2_axb_13),.CI(inf_abs0_2_cry_12),.O(inf_abs0_2[13:13]));
  MUXCY_L inf_abs0_2_cry_13_cZ(.DI(GND),.CI(inf_abs0_2_cry_12),.S(inf_abs0_2_axb_13),.LO(inf_abs0_2_cry_13));
  XORCY inf_abs0_2_s_12(.LI(inf_abs0_2_axb_12),.CI(inf_abs0_2_cry_11),.O(inf_abs0_2[12:12]));
  MUXCY_L inf_abs0_2_cry_12_cZ(.DI(GND),.CI(inf_abs0_2_cry_11),.S(inf_abs0_2_axb_12),.LO(inf_abs0_2_cry_12));
  XORCY inf_abs0_2_s_11(.LI(inf_abs0_2_axb_11),.CI(inf_abs0_2_cry_10),.O(inf_abs0_2[11:11]));
  MUXCY_L inf_abs0_2_cry_11_cZ(.DI(GND),.CI(inf_abs0_2_cry_10),.S(inf_abs0_2_axb_11),.LO(inf_abs0_2_cry_11));
  XORCY inf_abs0_2_s_10(.LI(inf_abs0_2_axb_10),.CI(inf_abs0_2_cry_9),.O(inf_abs0_2[10:10]));
  MUXCY_L inf_abs0_2_cry_10_cZ(.DI(GND),.CI(inf_abs0_2_cry_9),.S(inf_abs0_2_axb_10),.LO(inf_abs0_2_cry_10));
  XORCY inf_abs0_2_s_9(.LI(inf_abs0_2_axb_9),.CI(inf_abs0_2_cry_8),.O(inf_abs0_2[9:9]));
  MUXCY_L inf_abs0_2_cry_9_cZ(.DI(GND),.CI(inf_abs0_2_cry_8),.S(inf_abs0_2_axb_9),.LO(inf_abs0_2_cry_9));
  XORCY inf_abs0_2_s_8(.LI(inf_abs0_2_axb_8),.CI(inf_abs0_2_cry_7),.O(inf_abs0_2[8:8]));
  MUXCY_L inf_abs0_2_cry_8_cZ(.DI(GND),.CI(inf_abs0_2_cry_7),.S(inf_abs0_2_axb_8),.LO(inf_abs0_2_cry_8));
  XORCY inf_abs0_2_s_7(.LI(inf_abs0_2_axb_7),.CI(inf_abs0_2_cry_6),.O(inf_abs0_2[7:7]));
  MUXCY_L inf_abs0_2_cry_7_cZ(.DI(GND),.CI(inf_abs0_2_cry_6),.S(inf_abs0_2_axb_7),.LO(inf_abs0_2_cry_7));
  XORCY inf_abs0_2_s_6(.LI(inf_abs0_2_axb_6),.CI(inf_abs0_2_cry_5),.O(inf_abs0_2[6:6]));
  MUXCY_L inf_abs0_2_cry_6_cZ(.DI(GND),.CI(inf_abs0_2_cry_5),.S(inf_abs0_2_axb_6),.LO(inf_abs0_2_cry_6));
  XORCY inf_abs0_2_s_5(.LI(inf_abs0_2_axb_5),.CI(inf_abs0_2_cry_4),.O(inf_abs0_2[5:5]));
  MUXCY_L inf_abs0_2_cry_5_cZ(.DI(GND),.CI(inf_abs0_2_cry_4),.S(inf_abs0_2_axb_5),.LO(inf_abs0_2_cry_5));
  XORCY inf_abs0_2_s_4(.LI(inf_abs0_2_axb_4),.CI(inf_abs0_2_cry_3),.O(inf_abs0_2[4:4]));
  MUXCY_L inf_abs0_2_cry_4_cZ(.DI(GND),.CI(inf_abs0_2_cry_3),.S(inf_abs0_2_axb_4),.LO(inf_abs0_2_cry_4));
  XORCY inf_abs0_2_s_3(.LI(inf_abs0_2_axb_3),.CI(inf_abs0_2_cry_2),.O(inf_abs0_2[3:3]));
  MUXCY_L inf_abs0_2_cry_3_cZ(.DI(GND),.CI(inf_abs0_2_cry_2),.S(inf_abs0_2_axb_3),.LO(inf_abs0_2_cry_3));
  XORCY inf_abs0_2_s_2(.LI(inf_abs0_2_axb_2),.CI(inf_abs0_2_cry_1),.O(inf_abs0_2[2:2]));
  MUXCY_L inf_abs0_2_cry_2_cZ(.DI(GND),.CI(inf_abs0_2_cry_1),.S(inf_abs0_2_axb_2),.LO(inf_abs0_2_cry_2));
  XORCY inf_abs0_2_s_1(.LI(inf_abs0_2_axb_1),.CI(inf_abs0_2_cry_0),.O(inf_abs0_2[1:1]));
  MUXCY_L inf_abs0_2_cry_1_cZ(.DI(GND),.CI(inf_abs0_2_cry_0),.S(inf_abs0_2_axb_1),.LO(inf_abs0_2_cry_1));
  XORCY inf_abs0_2_s_0(.LI(inf_abs0_2_axb_0),.CI(ir_fast[31:31]),.O(inf_abs0_2[0:0]));
  MUXCY_L inf_abs0_2_cry_0_cZ(.DI(GND),.CI(ir_fast[31:31]),.S(inf_abs0_2_axb_0),.LO(inf_abs0_2_cry_0));
  LUT4 un26_r_lt30_cZ(.I0(m_2_i[31:31]),.I1(m_2[30:30]),.I2(r_4_i[31:31]),.I3(r_6[30:30]),.O(un26_r_lt30));
defparam un26_r_lt30_cZ.INIT=16'h0A8E;
  MUXCY_L desc1024(.DI(un26_r_lt28),.CI(un26_r_cry[26:26]),.S(un26_r_df28),.LO(un26_r_cry[28:28]));
  MUXCY_L desc1025(.DI(un26_r_lt26),.CI(un26_r_cry[24:24]),.S(un26_r_df26),.LO(un26_r_cry[26:26]));
  MUXCY_L desc1026(.DI(un26_r_lt24),.CI(un26_r_cry[22:22]),.S(un26_r_df24),.LO(un26_r_cry[24:24]));
  MUXCY_L desc1027(.DI(un26_r_lt22),.CI(un26_r_cry[20:20]),.S(un26_r_df22),.LO(un26_r_cry[22:22]));
  MUXCY_L desc1028(.DI(un26_r_lt20),.CI(un26_r_cry[18:18]),.S(un26_r_df20),.LO(un26_r_cry[20:20]));
  MUXCY_L desc1029(.DI(un26_r_lt18),.CI(un26_r_cry[16:16]),.S(un26_r_df18),.LO(un26_r_cry[18:18]));
  LUT4 un26_r_lt18_cZ(.I0(m_2[19:19]),.I1(m_2[18:18]),.I2(r_4[19:19]),.I3(r_4[18:18]),.O(un26_r_lt18));
defparam un26_r_lt18_cZ.INIT=16'h0A8E;
  MUXCY_L desc1030(.DI(un26_r_lt16),.CI(un26_r_cry[14:14]),.S(un26_r_df16),.LO(un26_r_cry[16:16]));
  LUT4 un26_r_lt16_cZ(.I0(m_2[16:16]),.I1(m_2[17:17]),.I2(r_4[16:16]),.I3(r_4[17:17]),.O(un26_r_lt16));
defparam un26_r_lt16_cZ.INIT=16'h08CE;
  MUXCY_L desc1031(.DI(un26_r_lt14),.CI(un26_r_cry[12:12]),.S(un26_r_df14),.LO(un26_r_cry[14:14]));
  LUT4 un26_r_lt14_cZ(.I0(m_2[14:14]),.I1(m_2[15:15]),.I2(r_4[14:14]),.I3(r_4[15:15]),.O(un26_r_lt14));
defparam un26_r_lt14_cZ.INIT=16'h08CE;
  MUXCY_L desc1032(.DI(un26_r_lt12),.CI(un26_r_cry[10:10]),.S(un26_r_df12),.LO(un26_r_cry[12:12]));
  LUT4 un26_r_lt12_cZ(.I0(m_2[12:12]),.I1(m_2[13:13]),.I2(r_4[12:12]),.I3(r_4[13:13]),.O(un26_r_lt12));
defparam un26_r_lt12_cZ.INIT=16'h08CE;
  MUXCY_L desc1033(.DI(un26_r_lt10),.CI(un26_r_cry[8:8]),.S(un26_r_df10),.LO(un26_r_cry[10:10]));
  LUT4 un26_r_lt10_cZ(.I0(m_2[10:10]),.I1(m_2[11:11]),.I2(r_4[11:11]),.I3(r_4[10:10]),.O(un26_r_lt10));
defparam un26_r_lt10_cZ.INIT=16'h0C8E;
  MUXCY_L desc1034(.DI(un26_r_lt8),.CI(un26_r_cry[6:6]),.S(un26_r_df8),.LO(un26_r_cry[8:8]));
  LUT4 un26_r_lt8_cZ(.I0(m_2[8:8]),.I1(m_2[9:9]),.I2(r_4[8:8]),.I3(r_4[9:9]),.O(un26_r_lt8));
defparam un26_r_lt8_cZ.INIT=16'h08CE;
  MUXCY_L desc1035(.DI(un26_r_lt6),.CI(un26_r_cry[4:4]),.S(un26_r_df6),.LO(un26_r_cry[6:6]));
  LUT4 un26_r_lt6_cZ(.I0(m_2[7:7]),.I1(m_2[6:6]),.I2(r_4[6:6]),.I3(r_4[7:7]),.O(un26_r_lt6));
defparam un26_r_lt6_cZ.INIT=16'h08AE;
  MUXCY_L desc1036(.DI(un26_r_lt4),.CI(un26_r_cry[2:2]),.S(un26_r_df4),.LO(un26_r_cry[4:4]));
  LUT4 un26_r_lt4_cZ(.I0(m_2[4:4]),.I1(m_2[5:5]),.I2(r_4[4:4]),.I3(r_4[5:5]),.O(un26_r_lt4));
defparam un26_r_lt4_cZ.INIT=16'h08CE;
  MUXCY_L desc1037(.DI(un26_r_lt2),.CI(un26_r_cry[0:0]),.S(un26_r_df2),.LO(un26_r_cry[2:2]));
  LUT4 un26_r_lt2_cZ(.I0(m_2[2:2]),.I1(m_2[3:3]),.I2(r_4[3:3]),.I3(N_28),.O(un26_r_lt2));
defparam un26_r_lt2_cZ.INIT=16'h0C8E;
  MUXCY_L desc1038(.DI(un26_r_lt0),.CI(GND),.S(un26_r_df0),.LO(un26_r_cry[0:0]));
  LUT4 un26_r_lt0_cZ(.I0(m_2[1:1]),.I1(m_2[0:0]),.I2(r_4[0:0]),.I3(r_4[1:1]),.O(un26_r_lt0));
defparam un26_r_lt0_cZ.INIT=16'h08AE;
  MUXCY_L desc1039(.DI(b18_lt28),.CI(b18_cry[26:26]),.S(b18_df28),.LO(b18_cry[28:28]));
  MUXCY_L desc1040(.DI(b18_lt26),.CI(b18_cry[24:24]),.S(b18_df26),.LO(b18_cry[26:26]));
  MUXCY_L desc1041(.DI(b18_lt24),.CI(b18_cry[22:22]),.S(b18_df24),.LO(b18_cry[24:24]));
  MUXCY_L desc1042(.DI(b18_lt22),.CI(b18_cry[20:20]),.S(b18_df22),.LO(b18_cry[22:22]));
  MUXCY_L desc1043(.DI(b18_lt20),.CI(b18_cry[18:18]),.S(b18_df20),.LO(b18_cry[20:20]));
  MUXCY_L desc1044(.DI(b18_lt18),.CI(b18_cry[16:16]),.S(b18_df18),.LO(b18_cry[18:18]));
  LUT4 b18_lt18_cZ(.I0(m_2[19:19]),.I1(m_2[18:18]),.I2(r_4[19:19]),.I3(r_4[18:18]),.O(b18_lt18));
defparam b18_lt18_cZ.INIT=16'h7150;
  MUXCY_L desc1045(.DI(b18_lt16),.CI(b18_cry[14:14]),.S(b18_df16),.LO(b18_cry[16:16]));
  LUT4 b18_lt16_cZ(.I0(m_2[16:16]),.I1(m_2[17:17]),.I2(r_4[16:16]),.I3(r_4[17:17]),.O(b18_lt16));
defparam b18_lt16_cZ.INIT=16'h7310;
  MUXCY_L desc1046(.DI(b18_lt14),.CI(b18_cry[12:12]),.S(b18_df14),.LO(b18_cry[14:14]));
  LUT4 b18_lt14_cZ(.I0(m_2[14:14]),.I1(m_2[15:15]),.I2(r_4[14:14]),.I3(r_4[15:15]),.O(b18_lt14));
defparam b18_lt14_cZ.INIT=16'h7310;
  MUXCY_L desc1047(.DI(b18_lt12),.CI(b18_cry[10:10]),.S(b18_df12),.LO(b18_cry[12:12]));
  LUT4 b18_lt12_cZ(.I0(m_2[12:12]),.I1(m_2[13:13]),.I2(r_4[12:12]),.I3(r_4[13:13]),.O(b18_lt12));
defparam b18_lt12_cZ.INIT=16'h7310;
  MUXCY_L desc1048(.DI(b18_lt10),.CI(b18_cry[8:8]),.S(b18_df10),.LO(b18_cry[10:10]));
  LUT4 b18_lt10_cZ(.I0(m_2[10:10]),.I1(m_2[11:11]),.I2(r_4[11:11]),.I3(r_4[10:10]),.O(b18_lt10));
defparam b18_lt10_cZ.INIT=16'h7130;
  MUXCY_L desc1049(.DI(b18_lt8),.CI(b18_cry[6:6]),.S(b18_df8),.LO(b18_cry[8:8]));
  LUT4 b18_lt8_cZ(.I0(m_2[8:8]),.I1(m_2[9:9]),.I2(r_4[8:8]),.I3(r_4[9:9]),.O(b18_lt8));
defparam b18_lt8_cZ.INIT=16'h7310;
  MUXCY_L desc1050(.DI(b18_lt6),.CI(b18_cry[4:4]),.S(b18_df6),.LO(b18_cry[6:6]));
  LUT4 b18_lt6_cZ(.I0(m_2[7:7]),.I1(m_2[6:6]),.I2(r_4[6:6]),.I3(r_4[7:7]),.O(b18_lt6));
defparam b18_lt6_cZ.INIT=16'h7510;
  MUXCY_L desc1051(.DI(b18_lt4),.CI(b18_cry[2:2]),.S(b18_df4),.LO(b18_cry[4:4]));
  LUT4 b18_lt4_cZ(.I0(m_2[4:4]),.I1(m_2[5:5]),.I2(r_4[4:4]),.I3(r_4[5:5]),.O(b18_lt4));
defparam b18_lt4_cZ.INIT=16'h7310;
  MUXCY_L desc1052(.DI(b18_lt2),.CI(b18_cry[0:0]),.S(b18_df2),.LO(b18_cry[2:2]));
  LUT4 b18_lt2_cZ(.I0(m_2[2:2]),.I1(m_2[3:3]),.I2(r_4[3:3]),.I3(N_28),.O(b18_lt2));
defparam b18_lt2_cZ.INIT=16'h7130;
  MUXCY_L desc1053(.DI(b18_lt0),.CI(GND),.S(b18_df0),.LO(b18_cry[0:0]));
  LUT4 b18_lt0_cZ(.I0(m_2[1:1]),.I1(m_2[0:0]),.I2(r_4[0:0]),.I3(r_4[1:1]),.O(b18_lt0));
defparam b18_lt0_cZ.INIT=16'h7510;
  MUXCY_L desc1054(.DI(un11_r_lt28),.CI(un11_r_cry[26:26]),.S(un11_r_df28),.LO(un11_r_cry[28:28]));
  MUXCY_L desc1055(.DI(un11_r_lt26),.CI(un11_r_cry[24:24]),.S(un11_r_df26),.LO(un11_r_cry[26:26]));
  MUXCY_L desc1056(.DI(un11_r_lt24),.CI(un11_r_cry[22:22]),.S(un11_r_df24),.LO(un11_r_cry[24:24]));
  MUXCY_L desc1057(.DI(un11_r_lt22),.CI(un11_r_cry[20:20]),.S(un11_r_df22),.LO(un11_r_cry[22:22]));
  MUXCY_L desc1058(.DI(un11_r_lt20),.CI(un11_r_cry[18:18]),.S(un11_r_df20),.LO(un11_r_cry[20:20]));
  MUXCY_L desc1059(.DI(un11_r_lt18),.CI(un11_r_cry[16:16]),.S(un11_r_df18),.LO(un11_r_cry[18:18]));
  LUT4 un11_r_lt18_cZ(.I0(m_2[19:19]),.I1(m_2[18:18]),.I2(r_4[19:19]),.I3(r_4[18:18]),.O(un11_r_lt18));
defparam un11_r_lt18_cZ.INIT=16'h0A8E;
  MUXCY_L desc1060(.DI(un11_r_lt16),.CI(un11_r_cry[14:14]),.S(un11_r_df16),.LO(un11_r_cry[16:16]));
  LUT4 un11_r_lt16_cZ(.I0(m_2[16:16]),.I1(m_2[17:17]),.I2(r_4[16:16]),.I3(r_4[17:17]),.O(un11_r_lt16));
defparam un11_r_lt16_cZ.INIT=16'h08CE;
  MUXCY_L desc1061(.DI(un11_r_lt14),.CI(un11_r_cry[12:12]),.S(un11_r_df14),.LO(un11_r_cry[14:14]));
  LUT4 un11_r_lt14_cZ(.I0(m_2[14:14]),.I1(m_2[15:15]),.I2(r_4[14:14]),.I3(r_4[15:15]),.O(un11_r_lt14));
defparam un11_r_lt14_cZ.INIT=16'h08CE;
  MUXCY_L desc1062(.DI(un11_r_lt12),.CI(un11_r_cry[10:10]),.S(un11_r_df12),.LO(un11_r_cry[12:12]));
  LUT4 un11_r_lt12_cZ(.I0(m_2[12:12]),.I1(m_2[13:13]),.I2(r_4[12:12]),.I3(r_4[13:13]),.O(un11_r_lt12));
defparam un11_r_lt12_cZ.INIT=16'h08CE;
  MUXCY_L desc1063(.DI(un11_r_lt10),.CI(un11_r_cry[8:8]),.S(un11_r_df10),.LO(un11_r_cry[10:10]));
  LUT4 un11_r_lt10_cZ(.I0(m_2[10:10]),.I1(m_2[11:11]),.I2(r_4[11:11]),.I3(r_4[10:10]),.O(un11_r_lt10));
defparam un11_r_lt10_cZ.INIT=16'h0C8E;
  MUXCY_L desc1064(.DI(un11_r_lt8),.CI(un11_r_cry[6:6]),.S(un11_r_df8),.LO(un11_r_cry[8:8]));
  LUT4 un11_r_lt8_cZ(.I0(m_2[8:8]),.I1(m_2[9:9]),.I2(r_4[8:8]),.I3(r_4[9:9]),.O(un11_r_lt8));
defparam un11_r_lt8_cZ.INIT=16'h08CE;
  MUXCY_L desc1065(.DI(un11_r_lt6),.CI(un11_r_cry[4:4]),.S(un11_r_df6),.LO(un11_r_cry[6:6]));
  LUT4 un11_r_lt6_cZ(.I0(m_2[7:7]),.I1(m_2[6:6]),.I2(r_4[6:6]),.I3(r_4[7:7]),.O(un11_r_lt6));
defparam un11_r_lt6_cZ.INIT=16'h08AE;
  MUXCY_L desc1066(.DI(un11_r_lt4),.CI(un11_r_cry[2:2]),.S(un11_r_df4),.LO(un11_r_cry[4:4]));
  LUT4 un11_r_lt4_cZ(.I0(m_2[4:4]),.I1(m_2[5:5]),.I2(r_4[4:4]),.I3(r_4[5:5]),.O(un11_r_lt4));
defparam un11_r_lt4_cZ.INIT=16'h08CE;
  MUXCY_L desc1067(.DI(un11_r_lt2),.CI(un11_r_cry[0:0]),.S(un11_r_df2),.LO(un11_r_cry[2:2]));
  LUT4 un11_r_lt2_cZ(.I0(m_2[2:2]),.I1(m_2[3:3]),.I2(r_4[3:3]),.I3(N_28),.O(un11_r_lt2));
defparam un11_r_lt2_cZ.INIT=16'h0C8E;
  MUXCY_L desc1068(.DI(un11_r_lt0),.CI(GND),.S(un11_r_df0),.LO(un11_r_cry[0:0]));
  LUT4 un11_r_lt0_cZ(.I0(m_2[1:1]),.I1(m_2[0:0]),.I2(r_4[0:0]),.I3(r_4[1:1]),.O(un11_r_lt0));
defparam un11_r_lt0_cZ.INIT=16'h08AE;
  MUXCY_L un14_r_0_I_75(.DI(GND),.CI(un14_r_0_data_tmp[3:3]),.S(un14_r_0_N_7),.LO(un14_r_0_data_tmp[4:4]));
  MUXCY_L un14_r_0_I_67(.DI(GND),.CI(un14_r_0_data_tmp[0:0]),.S(un14_r_0_N_14),.LO(un14_r_0_data_tmp[1:1]));
  MUXCY_L un14_r_0_I_59(.DI(GND),.CI(un14_r_0_data_tmp[1:1]),.S(un14_r_0_N_21),.LO(un14_r_0_data_tmp[2:2]));
  MUXCY_L un14_r_0_I_51(.DI(GND),.CI(un14_r_0_data_tmp[2:2]),.S(un14_r_0_N_28),.LO(un14_r_0_data_tmp[3:3]));
  MUXCY_L un14_r_0_I_43(.DI(GND),.CI(un14_r_0_data_tmp[7:7]),.S(un14_r_0_N_35),.LO(un14_r_0_data_tmp[8:8]));
  MUXCY_L un14_r_0_I_35(.DI(GND),.CI(un14_r_0_data_tmp[4:4]),.S(un14_r_0_N_42),.LO(un14_r_0_data_tmp[5:5]));
  MUXCY_L un14_r_0_I_27(.DI(GND),.CI(un14_r_0_data_tmp[5:5]),.S(un14_r_0_N_49),.LO(un14_r_0_data_tmp[6:6]));
  MUXCY_L un14_r_0_I_19(.DI(GND),.CI(un14_r_0_data_tmp[6:6]),.S(un14_r_0_N_56),.LO(un14_r_0_data_tmp[7:7]));
  MUXCY_L un14_r_0_I_11(.DI(GND),.CI(un14_r_0_data_tmp[8:8]),.S(un14_r_0_N_63),.LO(un14_r_0_data_tmp[9:9]));
  MUXCY_L un14_r_0_I_1(.DI(GND),.CI(VCC),.S(un14_r_0_N_70),.LO(un14_r_0_data_tmp[0:0]));
  LUT4 desc1069(.I0(inf_abs0_2[20:20]),.I1(inf_abs0_2[21:21]),.I2(inf_abs0_2[22:22]),.I3(reg3_1_1[21:21]),.O(\d_cnst_sn.reg0_28_5_2426_a6_1_1 ));
defparam desc1069.INIT=16'h0100;
  LUT3 desc1070(.I0(inf_abs0_2[20:20]),.I1(inf_abs0_2[21:21]),.I2(inf_abs0_2[22:22]),.O(\d_cnst_sn.reg0_28_12_2195_a6_1_2_0 ));
defparam desc1070.INIT=8'h01;
  LUT4 desc1071(.I0(inf_abs0_2[20:20]),.I1(inf_abs0_2[21:21]),.I2(inf_abs0_2[22:22]),.I3(reg3_1_1[25:25]),.O(\d_cnst_sn.reg0_28_9_2294_a6_1_1 ));
defparam desc1071.INIT=16'h0100;
  LUT4 desc1072(.I0(inf_abs0_2[20:20]),.I1(inf_abs0_2[21:21]),.I2(inf_abs0_2[22:22]),.I3(reg3_1_1[26:26]),.O(\d_cnst_sn.reg0_28_10_2261_a6_1_1 ));
defparam desc1072.INIT=16'h0100;
  LUT2 desc1073(.I0(reg1[3:3]),.I1(inf_abs0_2[30:30]),.O(r_4_2_a1_lut6_2_O6[3:3]));
defparam desc1073.INIT=4'h1;
  LUT2 desc1074(.I0(reg1[4:4]),.I1(inf_abs0_2[30:30]),.O(r_4_2_a1_lut6_2_O5[3:3]));
defparam desc1074.INIT=4'h1;
  LUT4 desc1075(.I0(inf_abs0_2[20:20]),.I1(inf_abs0_2[21:21]),.I2(inf_abs0_2[22:22]),.I3(reg3_1_1[23:23]),.O(\d_cnst_sn.reg0_28_7_2360_a6_1_1 ));
defparam desc1075.INIT=16'h0100;
  LUT2 desc1076(.I0(inf_abs0_2[21:21]),.I1(inf_abs0_2[22:22]),.O(N_3873_2));
defparam desc1076.INIT=4'h1;
  LUT2 desc1077(.I0(datai[31:31]),.I1(inf_abs0_2[20:20]),.O(\d_cnst_sn.g0_0_0_a5_0_0 ));
defparam desc1077.INIT=4'h8;
  LUT3 desc1078(.I0(datai[20:20]),.I1(state),.I2(inf_abs0_2[20:20]),.O(ir_3[20:20]));
defparam desc1078.INIT=8'hE2;
  LUT3 desc1079(.I0(state),.I1(inf_abs0_2[27:27]),.I2(inf_abs0_2[28:28]),.O(\d_cnst_sn.addr_20_iv_1052_i_a6_2_0 ));
defparam desc1079.INIT=8'h80;
  LUT3 desc1080(.I0(datai[30:30]),.I1(state),.I2(inf_abs0_2[30:30]),.O(ir_3[30:30]));
defparam desc1080.INIT=8'hE2;
  LUT2 desc1081(.I0(state),.I1(inf_abs0_2[27:27]),.O(\d_cnst_sn.addr_20_iv_1052_i_a6_1_0 ));
defparam desc1081.INIT=4'h2;
  LUT3 desc1082(.I0(datai[31:31]),.I1(state),.I2(inf_abs0_2[31:31]),.O(ir_3[31:31]));
defparam desc1082.INIT=8'hE2;
  LUT3 desc1083(.I0(inf_abs0_2[20:20]),.I1(inf_abs0_2[21:21]),.I2(inf_abs0_2[22:22]),.O(\d_cnst_sn.reg0_28_2526_a5_1_0 ));
defparam desc1083.INIT=8'h01;
  LUT4 desc1084(.I0(inf_abs0_2[21:21]),.I1(inf_abs0_2[22:22]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[28:28]),.O(\d_cnst_sn.g0_0_0_a5_2 ));
defparam desc1084.INIT=16'h0008;
  LUT4 desc1085(.I0(inf_abs0_2[20:20]),.I1(inf_abs0_2[21:21]),.I2(inf_abs0_2[22:22]),.I3(inf_abs0_2[31:31]),.O(\d_cnst_sn.reg0_N_13_0 ));
defparam desc1085.INIT=16'h003E;
  LUT3 desc1086(.I0(inf_abs0_2[21:21]),.I1(inf_abs0_2[22:22]),.I2(inf_abs0_2[31:31]),.O(\d_cnst_sn.reg0_m8_e_0 ));
defparam desc1086.INIT=8'h07;
  LUT4 desc1087(.I0(inf_abs0_2[20:20]),.I1(inf_abs0_2[21:21]),.I2(inf_abs0_2[22:22]),.I3(reg3_1_1[24:24]),.O(\d_cnst_sn.reg0_28_8_2327_a6_1_1 ));
defparam desc1087.INIT=16'h0100;
  LUT3 desc1088(.I0(inf_abs0_2[21:21]),.I1(inf_abs0_2[22:22]),.I2(inf_abs0_2[31:31]),.O(\d_cnst_sn.reg1_16_8_1837_2_tz ));
defparam desc1088.INIT=8'hF8;
  LUT2 desc1089(.I0(inf_abs0_2[31:31]),.I1(inf_abs0_2[28:28]),.O(N_527_i));
defparam desc1089.INIT=4'h4;
  LUT5 desc1090(.I0(inf_abs0_2[21:21]),.I1(inf_abs0_2[31:31]),.I2(inf_abs0_2[28:28]),.I3(r_4[18:18]),.I4(reg3_1_1[19:19]),.O(\d_cnst_sn.reg0_28_0 [19:19]));
defparam desc1090.INIT=32'hFFDF2202;
  LUT4 desc1091(.I0(reg3[19:19]),.I1(state),.I2(inf_abs0_2[19:19]),.I3(inf_abs0_2[28:28]),.O(\d_cnst_sn.addr_20_iv_6_863_i_0 ));
defparam desc1091.INIT=16'h111D;
  LUT3 desc1092(.I0(datai[28:28]),.I1(state),.I2(inf_abs0_2[28:28]),.O(ir_3[28:28]));
defparam desc1092.INIT=8'hE2;
  LUT2 desc1093(.I0(inf_abs0_2[27:27]),.I1(inf_abs0_2[28:28]),.O(g0_2_0_i2_lut6_2_O6));
defparam desc1093.INIT=4'h1;
  LUT4 desc1094(.I0(reg3[18:18]),.I1(state),.I2(inf_abs0_2[18:18]),.I3(inf_abs0_2[28:28]),.O(\d_cnst_sn.addr_20_iv_5_890_i_0 ));
defparam desc1094.INIT=16'h111D;
  LUT4 desc1095(.I0(reg3[17:17]),.I1(state),.I2(inf_abs0_2[17:17]),.I3(inf_abs0_2[28:28]),.O(\d_cnst_sn.addr_20_iv_4_917_i_0 ));
defparam desc1095.INIT=16'h111D;
  LUT3 desc1096(.I0(datai[17:17]),.I1(state),.I2(inf_abs0_2[17:17]),.O(ir_3[17:17]));
defparam desc1096.INIT=8'hE2;
  LUT2 desc1097(.I0(inf_abs0_2[27:27]),.I1(inf_abs0_2[28:28]),.O(N_7));
defparam desc1097.INIT=4'hE;
  LUT4 desc1098(.I0(reg3[16:16]),.I1(state),.I2(inf_abs0_2[16:16]),.I3(inf_abs0_2[28:28]),.O(\d_cnst_sn.addr_20_iv_3_944_i_0 ));
defparam desc1098.INIT=16'h111D;
  LUT4 desc1099(.I0(reg3[13:13]),.I1(state),.I2(inf_abs0_2[13:13]),.I3(inf_abs0_2[28:28]),.O(\d_cnst_sn.addr_20_iv_0_1025_i_0 ));
defparam desc1099.INIT=16'h111D;
  LUT3 desc1100(.I0(datai[13:13]),.I1(state),.I2(inf_abs0_2[13:13]),.O(ir_3[13:13]));
defparam desc1100.INIT=8'hE2;
  LUT4 desc1101(.I0(reg3[12:12]),.I1(state),.I2(inf_abs0_2[12:12]),.I3(inf_abs0_2[28:28]),.O(\d_cnst_sn.addr_20_iv_1052_i_0 ));
defparam desc1101.INIT=16'h111D;
  LUT3 desc1102(.I0(datai[12:12]),.I1(state),.I2(inf_abs0_2[12:12]),.O(ir_3[12:12]));
defparam desc1102.INIT=8'hE2;
  LUT4 desc1103(.I0(reg3[14:14]),.I1(state),.I2(inf_abs0_2[14:14]),.I3(inf_abs0_2[28:28]),.O(\d_cnst_sn.addr_20_iv_1_998_i_0 ));
defparam desc1103.INIT=16'h111D;
  LUT3 desc1104(.I0(datai[14:14]),.I1(state),.I2(inf_abs0_2[14:14]),.O(ir_3[14:14]));
defparam desc1104.INIT=8'hE2;
  LUT4 desc1105(.I0(reg3[15:15]),.I1(state),.I2(inf_abs0_2[15:15]),.I3(inf_abs0_2[28:28]),.O(\d_cnst_sn.addr_20_iv_2_971_i_0 ));
defparam desc1105.INIT=16'h111D;
  LUT3 desc1106(.I0(datai[15:15]),.I1(state),.I2(inf_abs0_2[15:15]),.O(ir_3[15:15]));
defparam desc1106.INIT=8'hE2;
  LUT4 desc1107(.I0(inf_abs0_2[20:20]),.I1(inf_abs0_2[21:21]),.I2(inf_abs0_2[22:22]),.I3(reg3_1_1[22:22]),.O(\d_cnst_sn.reg0_28_6_2393_a6_1_1 ));
defparam desc1107.INIT=16'h0100;
  LUT3 desc1108(.I0(inf_abs0_2[21:21]),.I1(inf_abs0_2[22:22]),.I2(inf_abs0_2[31:31]),.O(\d_cnst_sn.b60_0 ));
defparam desc1108.INIT=8'h02;
  LUT2 desc1109(.I0(inf_abs0_2[20:20]),.I1(inf_abs0_2[31:31]),.O(N_512_i));
defparam desc1109.INIT=4'h2;
  LUT3 desc1110(.I0(inf_abs0_2[21:21]),.I1(inf_abs0_2[22:22]),.I2(inf_abs0_2[31:31]),.O(\d_cnst_sn.reg0_m9_i_a3_0 ));
defparam desc1110.INIT=8'h06;
  LUT5 desc1111(.I0(inf_abs0_2[21:21]),.I1(inf_abs0_2[31:31]),.I2(inf_abs0_2[28:28]),.I3(r_4[19:19]),.I4(reg3_1_1[20:20]),.O(\d_cnst_sn.reg0_28_0 [20:20]));
defparam desc1111.INIT=32'hFFDF2202;
  LUT3 desc1112(.I0(inf_abs0_2[21:21]),.I1(inf_abs0_2[31:31]),.I2(inf_abs0_2[28:28]),.O(\d_cnst_sn.reg0_28_7_a0_0 [9:9]));
defparam desc1112.INIT=8'h02;
  LUT3 desc1113(.I0(inf_abs0_2[21:21]),.I1(inf_abs0_2[22:22]),.I2(inf_abs0_2[31:31]),.O(\d_cnst_sn.reg1_16_a2_0 [5:5]));
defparam desc1113.INIT=8'hF1;
  LUT2 desc1114(.I0(inf_abs0_2[19:19]),.I1(inf_abs0_2[31:31]),.O(N_3913));
defparam desc1114.INIT=4'hD;
  LUT3 desc1115(.I0(inf_abs0_2[19:19]),.I1(inf_abs0_2[20:20]),.I2(inf_abs0_2[31:31]),.O(\d_cnst_sn.reg2_N_3_mux ));
defparam desc1115.INIT=8'hF1;
  LUT5 desc1116(.I0(reg3[0:0]),.I1(inf_abs0_2[19:19]),.I2(inf_abs0_2[20:20]),.I3(inf_abs0_2[31:31]),.I4(m_2[0:0]),.O(N_1335));
defparam desc1116.INIT=32'hFFFB0008;
  LUT3 desc1117(.I0(inf_abs0_2[21:21]),.I1(inf_abs0_2[22:22]),.I2(inf_abs0_2[31:31]),.O(\d_cnst_sn.b64_0 ));
defparam desc1117.INIT=8'h04;
  LUT2 desc1118(.I0(inf_abs0_2[31:31]),.I1(inf_abs0_2[27:27]),.O(N_526_i));
defparam desc1118.INIT=4'h4;
  LUT4 desc1119(.I0(datai[30:30]),.I1(inf_abs0_2[31:31]),.I2(inf_abs0_2[27:27]),.I3(inf_abs0_2[28:28]),.O(m_2[30:30]));
defparam desc1119.INIT=16'h2220;
  LUT4 desc1120(.I0(datai[31:31]),.I1(inf_abs0_2[31:31]),.I2(inf_abs0_2[27:27]),.I3(inf_abs0_2[28:28]),.O(m_2[31:31]));
defparam desc1120.INIT=16'h2220;
  LUT3 desc1121(.I0(inf_abs0_2[21:21]),.I1(inf_abs0_2[22:22]),.I2(inf_abs0_2[31:31]),.O(N_3916));
defparam desc1121.INIT=8'h06;
  LUT3 desc1122(.I0(b),.I1(inf_abs0_2[31:31]),.I2(inf_abs0_2[27:27]),.O(reg0_28_sn_m6_lut6_2_O5));
defparam desc1122.INIT=8'h20;
  LUT4 desc1123(.I0(b),.I1(inf_abs0_2[21:21]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[27:27]),.O(\d_cnst_sn.reg0_m9_i_a0_0 ));
defparam desc1123.INIT=16'h040C;
  LUT2 desc1124(.I0(state),.I1(inf_abs0_2[27:27]),.O(N_2660_2));
defparam desc1124.INIT=4'h8;
  LUT4 desc1125(.I0(inf_abs0_2[20:20]),.I1(inf_abs0_2[21:21]),.I2(inf_abs0_2[22:22]),.I3(inf_abs0_2[31:31]),.O(N_3910));
defparam desc1125.INIT=16'h0002;
  LUT4 desc1126(.I0(inf_abs0_2[21:21]),.I1(inf_abs0_2[22:22]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[28:28]),.O(\d_cnst_sn.g0_3_a2_2 ));
defparam desc1126.INIT=16'h0008;
  LUT4 desc1127(.I0(inf_abs0_2[21:21]),.I1(inf_abs0_2[22:22]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[28:28]),.O(\d_cnst_sn.reg0_28_a1_1 [4:4]));
defparam desc1127.INIT=16'h0800;
  LUT4 desc1128(.I0(inf_abs0_2[20:20]),.I1(inf_abs0_2[21:21]),.I2(inf_abs0_2[22:22]),.I3(inf_abs0_2[31:31]),.O(\d_cnst_sn.reg0_28_9_2294_a6_3_0 ));
defparam desc1128.INIT=16'h0002;
  LUT4 desc1129(.I0(inf_abs0_2[20:20]),.I1(inf_abs0_2[21:21]),.I2(inf_abs0_2[22:22]),.I3(inf_abs0_2[31:31]),.O(\d_cnst_sn.reg0_28_a0_1 [7:7]));
defparam desc1129.INIT=16'hFF01;
  LUT4 desc1130(.I0(inf_abs0_2[21:21]),.I1(inf_abs0_2[22:22]),.I2(inf_abs0_2[31:31]),.I3(inf_abs0_2[28:28]),.O(\d_cnst_sn.reg1_16_a0_1 [3:3]));
defparam desc1130.INIT=16'h0008;
  LUT4 desc1131(.I0(datai[31:31]),.I1(inf_abs0_2[31:31]),.I2(inf_abs0_2[27:27]),.I3(inf_abs0_2[28:28]),.O(m_2_i[31:31]));
defparam desc1131.INIT=16'hDDDF;
  LUT3 desc1132(.I0(datai[31:31]),.I1(state),.I2(inf_abs0_2[31:31]),.O(ir_3_fast[31:31]));
defparam desc1132.INIT=8'hE2;
  LUT4 desc1133(.I0(inf_abs0_2[19:19]),.I1(inf_abs0_2[20:20]),.I2(inf_abs0_2[21:21]),.I3(inf_abs0_2[31:31]),.O(N_1033));
defparam desc1133.INIT=16'hFF35;
  LUT5 desc1134(.I0(inf_abs0_2[19:19]),.I1(inf_abs0_2[20:20]),.I2(inf_abs0_2[21:21]),.I3(inf_abs0_2[22:22]),.I4(inf_abs0_2[31:31]),.O(\d_cnst_sn.reg2_16_11_1_tz [28:28]));
defparam desc1134.INIT=32'hFFFFFACF;
  LUT5 desc1135(.I0(inf_abs0_2[19:19]),.I1(inf_abs0_2[20:20]),.I2(inf_abs0_2[21:21]),.I3(inf_abs0_2[22:22]),.I4(inf_abs0_2[31:31]),.O(N_1892));
defparam desc1135.INIT=32'h0000E000;
  LUT5 desc1136(.I0(inf_abs0_2[19:19]),.I1(inf_abs0_2[20:20]),.I2(inf_abs0_2[21:21]),.I3(inf_abs0_2[22:22]),.I4(inf_abs0_2[31:31]),.O(\d_cnst_sn.reg2_16_0_1_tz [28:28]));
defparam desc1136.INIT=32'hFFFFF53F;
  LUT4 b18_df30_lut6_2_o6(.I0(m_2_i[31:31]),.I1(r_4[30:30]),.I2(m_2[30:30]),.I3(r_4_i[31:31]),.O(b18_df30));
defparam b18_df30_lut6_2_o6.INIT=16'h8241;
  LUT4 b18_df30_lut6_2_o5(.I0(m_2_i[31:31]),.I1(r_4[30:30]),.I2(m_2[30:30]),.I3(r_4_i[31:31]),.O(b18_lt30));
defparam b18_df30_lut6_2_o5.INIT=16'h5D04;
  LUT4 un11_r_df30_lut6_2_o6(.I0(m_2_i[31:31]),.I1(r_4[30:30]),.I2(m_2[30:30]),.I3(r_4_i[31:31]),.O(un11_r_df30));
defparam un11_r_df30_lut6_2_o6.INIT=16'h8241;
  LUT4 un11_r_df30_lut6_2_o5(.I0(m_2_i[31:31]),.I1(r_4[30:30]),.I2(m_2[30:30]),.I3(r_4_i[31:31]),.O(un11_r_lt30));
defparam un11_r_df30_lut6_2_o5.INIT=16'h20BA;
endmodule