module \$__ABC9_LUT5 (input SEL, D, C, B, A, output Z);
	specify
		(SEL => Z) = 171;
		(D => Z) = 303;
		(C => Z) = 311;
		(B => Z) = 309;
		(A => Z) = 306;
	endspecify
endmodule