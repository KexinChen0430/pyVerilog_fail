module imp_test_mod2;
   import imp_test_pkg::*;
   word_t some_word;
endmodule