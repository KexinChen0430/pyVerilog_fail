module fir_inj (x_in,clk,y,p_desc0_p_O_FD,p_desc1_p_O_FD,p_desc2_p_O_FD,p_desc3_p_O_FD,p_desc4_p_O_FD,p_desc5_p_O_FD,p_desc6_p_O_FD,p_desc7_p_O_FD,p_desc8_p_O_FD,p_desc9_p_O_FD,p_desc10_p_O_FD,p_desc11_p_O_FD,p_desc12_p_O_FD,p_desc13_p_O_FD,p_desc14_p_O_FD,p_desc15_p_O_FD,p_desc16_p_O_FD,p_desc17_p_O_FD,p_desc18_p_O_FD,p_desc19_p_O_FD,p_desc20_p_O_FD,p_desc21_p_O_FD,p_desc22_p_O_FD,p_desc23_p_O_FD,p_desc24_p_O_FD,p_desc25_p_O_FD,p_desc26_p_O_FD,p_desc27_p_O_FD,p_desc28_p_O_FD,p_desc29_p_O_FD,p_desc30_p_O_FD,p_desc31_p_O_FD,p_desc32_p_O_FD,p_x_14_pipe_0_Z_p_O_FD,p_x_14_pipe_9_Z_p_O_FD,p_x_14_pipe_10_Z_p_O_FD,p_x_14_pipe_11_Z_p_O_FD,p_x_14_pipe_12_Z_p_O_FD,p_x_14_pipe_13_Z_p_O_FD,p_x_14_pipe_14_Z_p_O_FD,p_x_14_pipe_15_Z_p_O_FD,p_x_14_pipe_16_Z_p_O_FD,p_x_14_pipe_17_Z_p_O_FD,p_x_9_pipe_1_Z_p_O_FD,p_x_9_pipe_2_Z_p_O_FD,p_x_9_pipe_3_Z_p_O_FD,p_x_9_pipe_4_Z_p_O_FD,p_x_9_pipe_5_Z_p_O_FD,p_x_9_pipe_6_Z_p_O_FD,p_x_9_pipe_7_Z_p_O_FD,p_x_9_pipe_8_Z_p_O_FD,p_x_15_pipe_0_0_15_Z_p_O_FD,p_x_15_pipe_0_0_16_Z_p_O_FD,p_x_15_pipe_0_0_17_Z_p_O_FD,p_x_15_pipe_0_0_18_Z_p_O_FD,p_x_15_pipe_0_0_19_Z_p_O_FD,p_x_15_pipe_0_0_20_Z_p_O_FD,p_x_15_pipe_0_0_21_Z_p_O_FD,p_x_15_pipe_0_0_22_Z_p_O_FD,p_x_15_pipe_0_0_23_Z_p_O_FD,p_x_15_pipe_0_0_24_Z_p_O_FD,p_x_15_pipe_0_0_25_Z_p_O_FD,p_x_15_pipe_0_0_26_Z_p_O_FD,p_x_15_pipe_0_0_27_Z_p_O_FD,p_x_15_pipe_0_0_28_Z_p_O_FD,p_x_15_pipe_0_0_29_Z_p_O_FD,p_x_16_pipe_0_0_0_Z_p_O_FD,p_x_16_pipe_0_0_1_Z_p_O_FD,p_x_16_pipe_0_0_2_Z_p_O_FD,p_x_16_pipe_0_0_3_Z_p_O_FD,p_x_16_pipe_0_0_4_Z_p_O_FD,p_x_16_pipe_0_0_5_Z_p_O_FD,p_x_16_pipe_0_0_6_Z_p_O_FD,p_x_16_pipe_0_0_7_Z_p_O_FD,p_x_16_pipe_0_0_8_Z_p_O_FD,p_x_16_pipe_0_0_9_Z_p_O_FD,p_x_16_pipe_0_0_10_Z_p_O_FD,p_x_16_pipe_0_0_11_Z_p_O_FD,p_x_16_pipe_0_0_12_Z_p_O_FD,p_x_16_pipe_0_0_13_Z_p_O_FD,p_x_16_pipe_0_0_14_Z_p_O_FD,p_desc33_p_O_FD,p_desc34_p_O_FD,p_desc35_p_O_FD,p_desc36_p_O_FD,p_desc37_p_O_FD,p_desc38_p_O_FD,p_desc39_p_O_FD,p_desc40_p_O_FD,p_desc41_p_O_FD,p_desc42_p_O_FD,p_desc43_p_O_FD,p_desc44_p_O_FD,p_desc45_p_O_FD,p_desc46_p_O_FD,p_desc47_p_O_FD,p_desc48_p_O_FD,p_desc49_p_O_FD,p_desc50_p_O_FD,p_desc51_p_O_FD,p_desc52_p_O_FD,p_desc53_p_O_FD,p_desc54_p_O_FD,p_desc55_p_O_FD,p_desc56_p_O_FD);
input [7:0] x_in ;
input clk ;
output [7:0] y ;
wire clk ;
wire [7:0] x_0 ;
wire [15:4] un1_x_1 ;
wire [15:5] un1_x_2 ;
wire [15:4] un1_x_3 ;
wire [7:0] x_4 ;
wire [15:2] un1_x_4 ;
wire [14:0] un84_sop_0_0_0_0_5 ;
wire [7:0] x_7 ;
wire [7:0] x_8 ;
wire x_9 ;
wire [7:0] x_12 ;
wire [7:0] x_13 ;
wire [9:0] un84_sop_0_0_0_0_0 ;
wire [9:0] un84_sop_0_0_0_0_1 ;
wire [15:4] un1_x_14_0_0 ;
wire [15:5] un1_x_13_0_0 ;
wire [15:4] un1_x_12_0_0 ;
wire [14:7] un1_x_11_0_0 ;
wire [14:0] un84_sop_0_0_0_10_0 ;
wire [15:8] un1_x_10_0_0 ;
wire [15:5] un1_x_9_0 ;
wire [15:4] un1_x_8_0 ;
wire [15:2] un1_x_7_0 ;
wire [15:1] un1_x_6_0 ;
wire [14:0] un84_sop_0_0_0_5_0 ;
wire [47:11] P_uc ;
wire [29:0] ACOUT ;
wire [3:0] CARRYOUT ;
wire [47:0] PCOUT ;
wire [47:11] P_uc_0 ;
wire [29:0] ACOUT_0 ;
wire [3:0] CARRYOUT_0 ;
wire [47:0] PCOUT_0 ;
wire [47:11] P_uc_1 ;
wire [29:0] ACOUT_1 ;
wire [17:0] BCOUT_1 ;
wire [3:0] CARRYOUT_1 ;
wire [47:0] PCOUT_1 ;
wire [47:12] P_uc_2 ;
wire [29:0] ACOUT_2 ;
wire [3:0] CARRYOUT_2 ;
wire [47:0] PCOUT_2 ;
wire [47:12] P_uc_3 ;
wire [29:0] ACOUT_3 ;
wire [3:0] CARRYOUT_3 ;
wire [47:0] PCOUT_3 ;
wire [47:12] P_uc_4 ;
wire [29:0] ACOUT_4 ;
wire [3:0] CARRYOUT_4 ;
wire [47:0] PCOUT_4 ;
wire [47:12] P_uc_5 ;
wire [29:0] ACOUT_5 ;
wire [3:0] CARRYOUT_5 ;
wire [47:0] PCOUT_5 ;
wire [47:12] P_uc_6 ;
wire [29:0] ACOUT_6 ;
wire [3:0] CARRYOUT_6 ;
wire [47:0] PCOUT_6 ;
wire [47:14] P_uc_7 ;
wire [29:0] ACOUT_7 ;
wire [3:0] CARRYOUT_7 ;
wire [47:0] PCOUT_7 ;
wire [47:14] P_uc_8 ;
wire [29:0] ACOUT_8 ;
wire [3:0] CARRYOUT_8 ;
wire [47:0] PCOUT_8 ;
wire [47:15] P_uc_9 ;
wire [29:0] ACOUT_9 ;
wire [17:0] BCOUT_9 ;
wire [3:0] CARRYOUT_9 ;
wire [47:0] PCOUT_9 ;
wire [7:0] x_10_0 ;
wire [7:7] x_10_1 ;
wire [7:7] x_10_2 ;
wire [7:7] x_10_3 ;
wire [7:7] x_10_4 ;
wire [7:7] x_10_5 ;
wire [7:7] x_10_6 ;
wire [7:7] x_10_7 ;
wire [7:7] x_10_8 ;
wire [7:7] x_10_9 ;
wire [7:7] x_10_10 ;
wire [7:0] x_9_0 ;
wire [7:7] x_9_1 ;
wire [7:7] x_9_2 ;
wire [7:7] x_9_3 ;
wire [7:7] x_9_4 ;
wire [7:7] x_9_5 ;
wire [7:7] x_9_6 ;
wire [7:7] x_9_7 ;
wire [7:7] x_9_8 ;
wire [7:7] x_9_9 ;
wire [7:7] x_9_10 ;
wire [7:0] x_6_0 ;
wire [7:7] x_6_1 ;
wire [7:7] x_6_2 ;
wire [7:7] x_6_3 ;
wire [7:7] x_6_4 ;
wire [7:7] x_6_5 ;
wire [7:7] x_6_6 ;
wire [7:7] x_6_7 ;
wire [7:7] x_6_8 ;
wire [7:7] x_6_9 ;
wire [7:7] x_6_10 ;
wire [7:0] x_5_0 ;
wire [7:7] x_5_1 ;
wire [7:7] x_5_2 ;
wire [7:7] x_5_3 ;
wire [7:7] x_5_4 ;
wire [7:7] x_5_5 ;
wire [7:7] x_5_6 ;
wire [7:7] x_5_7 ;
wire [7:7] x_5_8 ;
wire [7:7] x_5_9 ;
wire [7:7] x_5_10 ;
wire [7:0] x_4_0 ;
wire [7:7] x_4_1 ;
wire [7:7] x_4_2 ;
wire [7:7] x_4_3 ;
wire [7:7] x_4_4 ;
wire [7:7] x_4_5 ;
wire [7:7] x_4_6 ;
wire [7:7] x_4_7 ;
wire [7:7] x_4_8 ;
wire [7:7] x_4_9 ;
wire [7:7] x_4_10 ;
wire [7:0] x_3_0 ;
wire [7:7] x_3_1 ;
wire [7:7] x_3_2 ;
wire [7:7] x_3_3 ;
wire [7:7] x_3_4 ;
wire [7:7] x_3_5 ;
wire [7:7] x_3_6 ;
wire [7:7] x_3_7 ;
wire [7:7] x_3_8 ;
wire [7:7] x_3_9 ;
wire [7:7] x_3_10 ;
wire [7:0] x_2_0 ;
wire [7:7] x_2_1 ;
wire [7:7] x_2_2 ;
wire [7:7] x_2_3 ;
wire [7:7] x_2_4 ;
wire [7:7] x_2_5 ;
wire [7:7] x_2_6 ;
wire [7:7] x_2_7 ;
wire [7:7] x_2_8 ;
wire [7:7] x_2_9 ;
wire [7:7] x_2_10 ;
wire [7:0] x_1_0 ;
wire [7:7] x_1_1 ;
wire [7:7] x_1_2 ;
wire [7:7] x_1_3 ;
wire [7:7] x_1_4 ;
wire [7:7] x_1_5 ;
wire [7:7] x_1_6 ;
wire [7:7] x_1_7 ;
wire [7:7] x_1_8 ;
wire [7:7] x_1_9 ;
wire [7:7] x_1_10 ;
wire [7:0] x_0_0 ;
wire [7:7] x_0_1 ;
wire [7:7] x_0_2 ;
wire [7:7] x_0_3 ;
wire [7:7] x_0_4 ;
wire [7:7] x_0_5 ;
wire [7:7] x_0_6 ;
wire [7:7] x_0_7 ;
wire [7:7] x_0_8 ;
wire [7:7] x_0_9 ;
wire [7:7] x_0_10 ;
wire [14:3] un84_sop_0_0_0_1_6_8 ;
wire [14:0] un84_sop_1_7 ;
wire [14:0] un84_sop_0_0_0_0_11_7 ;
wire [14:0] un84_sop_1_4 ;
wire [10:2] un1_x_10_4 ;
wire [14:0] un84_sop_0_0_0_1_6_4 ;
wire [14:0] un84_sop_0_0_0_0_11_6 ;
wire [14:0] un84_sop_0_0_0_0_8 ;
wire [14:0] un84_sop_0_0_0_1_6_6 ;
wire [14:0] un84_sop_1_6 ;
wire [14:7] un1_x_15_0_0_0 ;
wire [14:7] un1_x_11_0_0_0 ;
wire [14:7] un1_x_16_0_0_0 ;
wire x_12_6_tmp_d_array_0 ;
wire x_12_5_tmp_d_array_0 ;
wire x_12_4_tmp_d_array_0 ;
wire x_12_3_tmp_d_array_0 ;
wire x_12_2_tmp_d_array_0 ;
wire x_12_1_tmp_d_array_0 ;
wire x_12_0_tmp_d_array_0 ;
wire x_12_tmp_d_array_0 ;
wire x_7_6_tmp_d_array_0 ;
wire x_7_5_tmp_d_array_0 ;
wire x_7_4_tmp_d_array_0 ;
wire x_7_3_tmp_d_array_0 ;
wire x_7_2_tmp_d_array_0 ;
wire x_7_1_tmp_d_array_0 ;
wire x_7_0_tmp_d_array_0 ;
wire x_7_tmp_d_array_0 ;
wire x_4_6_tmp_d_array_0 ;
wire x_4_5_tmp_d_array_0 ;
wire x_4_4_tmp_d_array_0 ;
wire x_4_3_tmp_d_array_0 ;
wire x_4_2_tmp_d_array_0 ;
wire x_4_1_tmp_d_array_0 ;
wire x_4_0_tmp_d_array_0 ;
wire x_4_tmp_d_array_0 ;
wire [4:4] un1_x_14_0_0_0 ;
wire [5:5] un1_x_9_0_0 ;
wire [4:4] un1_x_3_0 ;
wire VCC ;
wire GND ;
wire un84_sop_1_s_7 ;
wire un84_sop_1_s_8 ;
wire un84_sop_1_s_9 ;
wire un84_sop_1_s_10 ;
wire un84_sop_1_s_11 ;
wire un84_sop_1_s_12 ;
wire un84_sop_1_s_13 ;
wire un84_sop_1_s_14 ;
wire un1_x_10_s_2_sf ;
wire un1_x_10_axb_3 ;
wire CARRYCASCOUT ;
wire OVERFLOW ;
wire MULTSIGNOUT ;
wire PATTERNBDETECT ;
wire PATTERNDETECT ;
wire UNDERFLOW ;
wire CARRYCASCOUT_0 ;
wire OVERFLOW_0 ;
wire MULTSIGNOUT_0 ;
wire PATTERNBDETECT_0 ;
wire PATTERNDETECT_0 ;
wire UNDERFLOW_0 ;
wire CARRYCASCOUT_1 ;
wire OVERFLOW_1 ;
wire MULTSIGNOUT_1 ;
wire PATTERNBDETECT_1 ;
wire PATTERNDETECT_1 ;
wire UNDERFLOW_1 ;
wire CARRYCASCOUT_2 ;
wire OVERFLOW_2 ;
wire MULTSIGNOUT_2 ;
wire PATTERNBDETECT_2 ;
wire PATTERNDETECT_2 ;
wire UNDERFLOW_2 ;
wire CARRYCASCOUT_3 ;
wire OVERFLOW_3 ;
wire MULTSIGNOUT_3 ;
wire PATTERNBDETECT_3 ;
wire PATTERNDETECT_3 ;
wire UNDERFLOW_3 ;
wire CARRYCASCOUT_4 ;
wire OVERFLOW_4 ;
wire MULTSIGNOUT_4 ;
wire PATTERNBDETECT_4 ;
wire PATTERNDETECT_4 ;
wire UNDERFLOW_4 ;
wire CARRYCASCOUT_5 ;
wire OVERFLOW_5 ;
wire MULTSIGNOUT_5 ;
wire PATTERNBDETECT_5 ;
wire PATTERNDETECT_5 ;
wire UNDERFLOW_5 ;
wire CARRYCASCOUT_6 ;
wire OVERFLOW_6 ;
wire MULTSIGNOUT_6 ;
wire PATTERNBDETECT_6 ;
wire PATTERNDETECT_6 ;
wire UNDERFLOW_6 ;
wire CARRYCASCOUT_7 ;
wire OVERFLOW_7 ;
wire MULTSIGNOUT_7 ;
wire PATTERNBDETECT_7 ;
wire PATTERNDETECT_7 ;
wire UNDERFLOW_7 ;
wire CARRYCASCOUT_8 ;
wire OVERFLOW_8 ;
wire MULTSIGNOUT_8 ;
wire PATTERNBDETECT_8 ;
wire PATTERNDETECT_8 ;
wire UNDERFLOW_8 ;
wire CARRYCASCOUT_9 ;
wire OVERFLOW_9 ;
wire MULTSIGNOUT_9 ;
wire PATTERNBDETECT_9 ;
wire PATTERNDETECT_9 ;
wire UNDERFLOW_9 ;
wire un84_sop_1_6_0_axb_1_lut6_2_O5 ;
wire un84_sop_1_6_0_o5_2 ;
wire un84_sop_1_6_0_o5_3 ;
wire un84_sop_1_6_0_o5_4 ;
wire un84_sop_1_6_0_o5_5 ;
wire un84_sop_1_6_0_o5_6 ;
wire un84_sop_1_6_0_o5_7 ;
wire un84_sop_1_6_0_o5_8 ;
wire un84_sop_1_6_0_o5_9 ;
wire un84_sop_1_6_0_o5_10 ;
wire un84_sop_1_6_0_o5_11 ;
wire un84_sop_0_0_0_1_6_8_axb_2_lut6_2_O5 ;
wire un84_sop_0_0_0_1_6_8_o5_3 ;
wire un84_sop_0_0_0_1_6_8_o5_4 ;
wire un84_sop_0_0_0_1_6_8_o5_5 ;
wire un84_sop_0_0_0_1_6_8_o5_6 ;
wire un84_sop_0_0_0_1_6_8_o5_7 ;
wire un84_sop_0_0_0_6_6_0_axb_1_lut6_2_O5 ;
wire un84_sop_0_0_0_6_6_0_o5_2 ;
wire un84_sop_0_0_0_6_6_0_o5_3 ;
wire un84_sop_0_0_0_6_6_0_o5_4 ;
wire un84_sop_0_0_0_6_6_0_o5_5 ;
wire un84_sop_0_0_0_6_6_0_o5_6 ;
wire un84_sop_0_0_0_6_6_0_o5_7 ;
wire un84_sop_0_0_0_6_6_0_o5_8 ;
wire un84_sop_0_0_0_6_6_0_o5_9 ;
wire un84_sop_0_0_0_6_6_0_o5_10 ;
wire un84_sop_0_0_0_6_6_0_o5_11 ;
wire un84_sop_0_0_0_6_6_0_o5_12 ;
wire un84_sop_0_0_0_11_0_o5_2 ;
wire un84_sop_0_0_0_11_0_o5_3 ;
wire un84_sop_0_0_0_11_0_o5_4 ;
wire un84_sop_0_0_0_11_0_o5_5 ;
wire un84_sop_0_0_0_11_0_o5_6 ;
wire un84_sop_0_0_0_11_0_o5_7 ;
wire un84_sop_0_0_0_11_0_o5_8 ;
wire un84_sop_0_0_0_11_0_o5_9 ;
wire un84_sop_0_0_0_11_0_o5_10 ;
wire un84_sop_0_0_0_11_0_o5_11 ;
wire un84_sop_0_0_0_11_0_o5_12 ;
wire un84_sop_0_0_0_11_6_0_axb_1_lut6_2_O5 ;
wire un84_sop_0_0_0_11_6_0_o5_2 ;
wire un84_sop_0_0_0_11_6_0_o5_3 ;
wire un84_sop_0_0_0_11_6_0_o5_4 ;
wire un84_sop_0_0_0_11_6_0_o5_5 ;
wire un84_sop_0_0_0_11_6_0_o5_6 ;
wire un84_sop_0_0_0_11_6_0_o5_7 ;
wire un84_sop_0_0_0_11_6_0_o5_8 ;
wire un84_sop_0_0_0_11_6_0_o5_9 ;
wire un84_sop_0_0_0_11_6_0_o5_10 ;
wire un84_sop_0_0_0_11_6_0_o5_11 ;
wire un84_sop_0_0_0_11_6_0_cry_0 ;
wire un84_sop_0_0_0_11_6_0_axb_1 ;
wire un84_sop_0_0_0_11_6_0_cry_1 ;
wire un84_sop_0_0_0_11_6_0_axb_2 ;
wire un84_sop_0_0_0_11_6_0_cry_2 ;
wire un84_sop_0_0_0_11_6_0_axb_3 ;
wire un84_sop_0_0_0_11_6_0_cry_3 ;
wire un84_sop_0_0_0_11_6_0_axb_4 ;
wire un84_sop_0_0_0_11_6_0_cry_4 ;
wire un84_sop_0_0_0_11_6_0_axb_5 ;
wire un84_sop_0_0_0_11_6_0_cry_5 ;
wire un84_sop_0_0_0_11_6_0_axb_6 ;
wire un84_sop_0_0_0_11_6_0_cry_6 ;
wire un84_sop_0_0_0_11_6_0_axb_7 ;
wire un84_sop_0_0_0_11_6_0_cry_7 ;
wire un84_sop_0_0_0_11_6_0_axb_8 ;
wire un84_sop_0_0_0_11_6_0_cry_8 ;
wire un84_sop_0_0_0_11_6_0_axb_9 ;
wire un84_sop_0_0_0_11_6_0_cry_9 ;
wire un84_sop_0_0_0_11_6_0_axb_10 ;
wire un84_sop_0_0_0_11_6_0_cry_10 ;
wire un84_sop_0_0_0_11_6_0_axb_11 ;
wire un84_sop_0_0_0_11_6_0_cry_11 ;
wire un84_sop_0_0_0_11_6_0_axb_12 ;
wire un84_sop_0_0_0_11_6_0_cry_12 ;
wire un84_sop_0_0_0_11_6_0_axb_13 ;
wire un84_sop_0_0_0_11_0_axb_0 ;
wire un84_sop_0_0_0_11_0_cry_0 ;
wire un84_sop_0_0_0_11_0_axb_1 ;
wire un84_sop_0_0_0_11_0_cry_1 ;
wire un84_sop_0_0_0_11_0_cry_2_RNO ;
wire un84_sop_0_0_0_11_0_axb_2 ;
wire un84_sop_0_0_0_11_0_cry_2 ;
wire un84_sop_0_0_0_11_0_axb_3 ;
wire un84_sop_0_0_0_11_0_cry_3 ;
wire un84_sop_0_0_0_11_0_axb_4 ;
wire un84_sop_0_0_0_11_0_cry_4 ;
wire un84_sop_0_0_0_11_0_axb_5 ;
wire un84_sop_0_0_0_11_0_cry_5 ;
wire un84_sop_0_0_0_11_0_axb_6 ;
wire un84_sop_0_0_0_11_0_cry_6 ;
wire un84_sop_0_0_0_11_0_axb_7 ;
wire un84_sop_0_0_0_11_0_cry_7 ;
wire un84_sop_0_0_0_11_0_axb_8 ;
wire un84_sop_0_0_0_11_0_cry_8 ;
wire un84_sop_0_0_0_11_0_axb_9 ;
wire un84_sop_0_0_0_11_0_cry_9 ;
wire un84_sop_0_0_0_11_0_axb_10 ;
wire un84_sop_0_0_0_11_0_cry_10 ;
wire un84_sop_0_0_0_11_0_axb_11 ;
wire un84_sop_0_0_0_11_0_cry_11 ;
wire un84_sop_0_0_0_11_0_axb_12 ;
wire un84_sop_0_0_0_11_0_cry_12 ;
wire un84_sop_0_0_0_11_0_axb_13 ;
wire un84_sop_0_0_0_11_0_cry_13 ;
wire un84_sop_0_0_0_11_0_axb_14 ;
wire un84_sop_0_0_0_6_6_0_cry_0 ;
wire un84_sop_0_0_0_6_6_0_axb_1 ;
wire un84_sop_0_0_0_6_6_0_cry_1 ;
wire un84_sop_0_0_0_6_6_0_axb_2 ;
wire un84_sop_0_0_0_6_6_0_cry_2 ;
wire un84_sop_0_0_0_6_6_0_axb_3 ;
wire un84_sop_0_0_0_6_6_0_cry_3 ;
wire un84_sop_0_0_0_6_6_0_axb_4 ;
wire un84_sop_0_0_0_6_6_0_cry_4 ;
wire un84_sop_0_0_0_6_6_0_axb_5 ;
wire un84_sop_0_0_0_6_6_0_cry_5 ;
wire un84_sop_0_0_0_6_6_0_axb_6 ;
wire un84_sop_0_0_0_6_6_0_cry_6 ;
wire un84_sop_0_0_0_6_6_0_axb_7 ;
wire un84_sop_0_0_0_6_6_0_cry_7 ;
wire un84_sop_0_0_0_6_6_0_axb_8 ;
wire un84_sop_0_0_0_6_6_0_cry_8 ;
wire un84_sop_0_0_0_6_6_0_axb_9 ;
wire un84_sop_0_0_0_6_6_0_cry_9 ;
wire un84_sop_0_0_0_6_6_0_axb_10 ;
wire un84_sop_0_0_0_6_6_0_cry_10 ;
wire un84_sop_0_0_0_6_6_0_axb_11 ;
wire un84_sop_0_0_0_6_6_0_cry_11 ;
wire un84_sop_0_0_0_6_6_0_axb_12 ;
wire un84_sop_0_0_0_6_6_0_cry_12 ;
wire un84_sop_0_0_0_6_6_0_axb_13 ;
wire un84_sop_0_0_0_6_6_0_cry_13 ;
wire un84_sop_0_0_0_6_6_0_axb_14 ;
wire un84_sop_0_0_0_1_6_8_cry_0 ;
wire un84_sop_0_0_0_1_6_8_axb_1 ;
wire un84_sop_0_0_0_1_6_8_cry_1 ;
wire un84_sop_0_0_0_1_6_8_axb_2 ;
wire un84_sop_0_0_0_1_6_8_cry_2 ;
wire un84_sop_0_0_0_1_6_8_axb_3 ;
wire un84_sop_0_0_0_1_6_8_cry_3 ;
wire un84_sop_0_0_0_1_6_8_axb_4 ;
wire un84_sop_0_0_0_1_6_8_cry_4 ;
wire un84_sop_0_0_0_1_6_8_axb_5 ;
wire un84_sop_0_0_0_1_6_8_cry_5 ;
wire un84_sop_0_0_0_1_6_8_axb_6 ;
wire un84_sop_0_0_0_1_6_8_cry_6 ;
wire un84_sop_0_0_0_1_6_8_axb_7 ;
wire un84_sop_0_0_0_1_6_8_cry_7 ;
wire un84_sop_0_0_0_1_6_8_axb_8 ;
wire un84_sop_0_0_0_1_6_8_cry_8 ;
wire un84_sop_0_0_0_1_6_8_axb_9 ;
wire un84_sop_0_0_0_1_6_8_cry_9 ;
wire un84_sop_0_0_0_1_6_8_axb_10 ;
wire un84_sop_0_0_0_1_6_8_cry_10 ;
wire un84_sop_0_0_0_1_6_8_axb_11 ;
wire un84_sop_1_6_0_cry_0 ;
wire un84_sop_1_6_0_axb_1 ;
wire un84_sop_1_6_0_cry_1 ;
wire un84_sop_1_6_0_axb_2 ;
wire un84_sop_1_6_0_cry_2 ;
wire un84_sop_1_6_0_axb_3 ;
wire un84_sop_1_6_0_cry_3 ;
wire un84_sop_1_6_0_axb_4 ;
wire un84_sop_1_6_0_cry_4 ;
wire un84_sop_1_6_0_axb_5 ;
wire un84_sop_1_6_0_cry_5 ;
wire un84_sop_1_6_0_axb_6 ;
wire un84_sop_1_6_0_cry_6 ;
wire un84_sop_1_6_0_axb_7 ;
wire un84_sop_1_6_0_cry_7 ;
wire un84_sop_1_6_0_axb_8 ;
wire un84_sop_1_6_0_cry_8 ;
wire un84_sop_1_6_0_axb_9 ;
wire un84_sop_1_6_0_cry_9 ;
wire un84_sop_1_6_0_axb_10 ;
wire un84_sop_1_6_0_cry_10 ;
wire un84_sop_1_6_0_axb_11 ;
wire un84_sop_1_6_0_cry_11 ;
wire un84_sop_1_6_0_axb_12 ;
wire un84_sop_1_6_0_cry_12 ;
wire un84_sop_1_6_0_axb_13 ;
wire un1_x_10_cry_3 ;
wire un1_x_10_axb_4 ;
wire un1_x_10_cry_4 ;
wire un1_x_10_axb_5 ;
wire un1_x_10_cry_5 ;
wire un1_x_10_axb_6 ;
wire un1_x_10_cry_6 ;
wire un1_x_10_axb_7 ;
wire un1_x_10_cry_7 ;
wire un1_x_10_axb_8 ;
wire un1_x_10_cry_8 ;
wire un1_x_10_axb_9 ;
wire un1_x_10_cry_9 ;
wire un1_x_10_axb_10 ;
wire un1_x_10_cry_10 ;
wire un1_x_10_axb_11 ;
wire un84_sop_0_0_0_1_6_4_cry_0 ;
wire un84_sop_0_0_0_1_6_4_axb_1 ;
wire un84_sop_0_0_0_1_6_4_cry_1 ;
wire un84_sop_0_0_0_1_6_4_axb_2 ;
wire un84_sop_0_0_0_1_6_4_cry_2 ;
wire un84_sop_0_0_0_1_6_4_axb_3 ;
wire un84_sop_0_0_0_1_6_4_cry_3 ;
wire un84_sop_0_0_0_1_6_4_axb_4 ;
wire un84_sop_0_0_0_1_6_4_cry_4 ;
wire un84_sop_0_0_0_1_6_4_axb_5 ;
wire un84_sop_0_0_0_1_6_4_cry_5 ;
wire un84_sop_0_0_0_1_6_4_axb_6 ;
wire un84_sop_0_0_0_1_6_4_cry_6 ;
wire un84_sop_0_0_0_1_6_4_axb_7 ;
wire un84_sop_0_0_0_1_6_4_cry_7 ;
wire un84_sop_0_0_0_1_6_4_axb_8 ;
wire un84_sop_0_0_0_1_6_4_cry_8 ;
wire un84_sop_0_0_0_1_6_4_axb_9 ;
wire un84_sop_0_0_0_1_6_4_cry_9 ;
wire un84_sop_0_0_0_1_6_4_axb_10 ;
wire un84_sop_0_0_0_1_6_4_cry_10 ;
wire un84_sop_0_0_0_1_6_4_axb_11 ;
wire un84_sop_0_0_0_1_6_4_cry_11 ;
wire un84_sop_0_0_0_1_6_4_axb_12 ;
wire un84_sop_0_0_0_1_6_4_cry_12 ;
wire un84_sop_0_0_0_1_6_4_axb_13 ;
wire un84_sop_0_0_0_1_6_4_cry_13 ;
wire un84_sop_0_0_0_1_6_4_axb_14 ;
wire un84_sop_0_0_0_1_6_cry_0 ;
wire un84_sop_0_0_0_1_6_axb_1 ;
wire un84_sop_0_0_0_1_6_cry_1 ;
wire un84_sop_0_0_0_1_6_axb_2 ;
wire un84_sop_0_0_0_1_6_cry_2 ;
wire un84_sop_0_0_0_1_6_axb_3 ;
wire un84_sop_0_0_0_1_6_cry_3 ;
wire un84_sop_0_0_0_1_6_axb_4 ;
wire un84_sop_0_0_0_1_6_cry_4 ;
wire un84_sop_0_0_0_1_6_axb_5 ;
wire un84_sop_0_0_0_1_6_cry_5 ;
wire un84_sop_0_0_0_1_6_axb_6 ;
wire un84_sop_0_0_0_1_6_cry_6 ;
wire un84_sop_0_0_0_1_6_axb_7 ;
wire un84_sop_0_0_0_1_6_cry_7 ;
wire un84_sop_0_0_0_1_6_axb_8 ;
wire un84_sop_0_0_0_1_6_cry_8 ;
wire un84_sop_0_0_0_1_6_axb_9 ;
wire un84_sop_0_0_0_1_6_cry_9 ;
wire un84_sop_0_0_0_1_6_axb_10 ;
wire un84_sop_0_0_0_1_6_cry_10 ;
wire un84_sop_0_0_0_1_6_axb_11 ;
wire un84_sop_0_0_0_1_6_cry_11 ;
wire un84_sop_0_0_0_1_6_axb_12 ;
wire un84_sop_0_0_0_1_6_cry_12 ;
wire un84_sop_0_0_0_1_6_axb_13 ;
wire un84_sop_0_0_0_1_6_cry_13 ;
wire un84_sop_0_0_0_1_6_axb_14 ;
wire un1_x_0_0_c4 ;
wire un1_x_10_5_c5 ;
wire un84_sop_1_7_cry_0 ;
wire un84_sop_1_7_axb_1 ;
wire un84_sop_1_7_cry_1 ;
wire un84_sop_1_7_axb_2 ;
wire un84_sop_1_7_cry_2 ;
wire un84_sop_1_7_axb_3 ;
wire un84_sop_1_7_cry_3 ;
wire un84_sop_1_7_axb_4 ;
wire un84_sop_1_7_cry_4 ;
wire un84_sop_1_7_axb_5 ;
wire un84_sop_1_7_cry_5 ;
wire un84_sop_1_7_axb_6 ;
wire un84_sop_1_7_cry_6 ;
wire un84_sop_1_7_axb_7 ;
wire un84_sop_1_7_cry_7 ;
wire un84_sop_1_7_axb_8 ;
wire un84_sop_1_7_cry_8 ;
wire un84_sop_1_7_axb_9 ;
wire un84_sop_1_7_cry_9 ;
wire un84_sop_1_7_axb_10 ;
wire un84_sop_1_7_cry_10 ;
wire un84_sop_1_7_axb_11 ;
wire un84_sop_1_7_cry_11 ;
wire un84_sop_1_7_axb_12 ;
wire un84_sop_1_7_cry_12 ;
wire un84_sop_1_7_axb_13 ;
wire un84_sop_1_7_cry_13 ;
wire un84_sop_1_7_axb_14 ;
wire un84_sop_0_0_0_0_11_7_cry_0 ;
wire un84_sop_0_0_0_0_11_7_axb_1 ;
wire un84_sop_0_0_0_0_11_7_cry_1 ;
wire un84_sop_0_0_0_0_11_7_axb_2 ;
wire un84_sop_0_0_0_0_11_7_cry_2 ;
wire un84_sop_0_0_0_0_11_7_axb_3 ;
wire un84_sop_0_0_0_0_11_7_cry_3 ;
wire un84_sop_0_0_0_0_11_7_axb_4 ;
wire un84_sop_0_0_0_0_11_7_cry_4 ;
wire un84_sop_0_0_0_0_11_7_axb_5 ;
wire un84_sop_0_0_0_0_11_7_cry_5 ;
wire un84_sop_0_0_0_0_11_7_axb_6 ;
wire un84_sop_0_0_0_0_11_7_cry_6 ;
wire un84_sop_0_0_0_0_11_7_axb_7 ;
wire un84_sop_0_0_0_0_11_7_cry_7 ;
wire un84_sop_0_0_0_0_11_7_axb_8 ;
wire un84_sop_0_0_0_0_11_7_cry_8 ;
wire un84_sop_0_0_0_0_11_7_axb_9 ;
wire un84_sop_0_0_0_0_11_7_cry_9 ;
wire un84_sop_0_0_0_0_11_7_axb_10 ;
wire un84_sop_1_4_cry_0 ;
wire un84_sop_1_4_axb_1 ;
wire un84_sop_1_4_cry_1 ;
wire un84_sop_1_4_axb_2 ;
wire un84_sop_1_4_cry_2 ;
wire un84_sop_1_4_axb_3 ;
wire un84_sop_1_4_cry_3 ;
wire un84_sop_1_4_axb_4 ;
wire un84_sop_1_4_cry_4 ;
wire un84_sop_1_4_axb_5 ;
wire un84_sop_1_4_cry_5 ;
wire un84_sop_1_4_axb_6 ;
wire un84_sop_1_4_cry_6 ;
wire un84_sop_1_4_axb_7 ;
wire un84_sop_1_4_cry_7 ;
wire un84_sop_1_4_axb_8 ;
wire un84_sop_1_4_cry_8 ;
wire un84_sop_1_4_axb_9 ;
wire un84_sop_1_4_cry_9 ;
wire un84_sop_1_4_axb_10 ;
wire un84_sop_1_4_cry_10 ;
wire un84_sop_1_4_axb_11 ;
wire un84_sop_1_4_cry_11 ;
wire un84_sop_1_4_axb_12 ;
wire un84_sop_1_4_cry_12 ;
wire un84_sop_1_4_axb_13 ;
wire un84_sop_1_4_cry_13 ;
wire un84_sop_1_4_axb_14 ;
wire un84_sop_1_axb_0 ;
wire un84_sop_1_cry_0 ;
wire un84_sop_1_axb_1 ;
wire un84_sop_1_cry_1 ;
wire un84_sop_1_axb_2 ;
wire un84_sop_1_cry_2 ;
wire un84_sop_1_axb_3 ;
wire un84_sop_1_cry_3 ;
wire un84_sop_1_axb_4 ;
wire un84_sop_1_cry_4 ;
wire un84_sop_1_axb_5 ;
wire un84_sop_1_cry_5 ;
wire un84_sop_1_axb_6 ;
wire un84_sop_1_cry_6 ;
wire un84_sop_1_axb_7 ;
wire un84_sop_1_cry_7 ;
wire un84_sop_1_axb_8 ;
wire un84_sop_1_cry_8 ;
wire un84_sop_1_axb_9 ;
wire un84_sop_1_cry_9 ;
wire un84_sop_1_axb_10 ;
wire un84_sop_1_cry_10 ;
wire un84_sop_1_axb_11 ;
wire un84_sop_1_cry_11 ;
wire un84_sop_1_axb_12 ;
wire un84_sop_1_cry_12 ;
wire un84_sop_1_axb_13 ;
wire un84_sop_1_cry_13 ;
wire un84_sop_1_axb_14 ;
wire un1_x_10_4_cry_1 ;
wire un1_x_10_4_axb_2 ;
wire un1_x_10_4_cry_2 ;
wire un1_x_10_4_axb_3 ;
wire un1_x_10_4_cry_3 ;
wire un1_x_10_4_axb_4 ;
wire un1_x_10_4_cry_4 ;
wire un1_x_10_4_axb_5 ;
wire un1_x_10_4_cry_5 ;
wire un1_x_10_4_axb_6 ;
wire un1_x_10_4_cry_6 ;
wire un1_x_10_4_axb_7 ;
wire un1_x_10_4_cry_7 ;
wire un1_x_15_0_axb_0 ;
wire un1_x_15_0_cry_0 ;
wire un1_x_15_0_axb_1 ;
wire un1_x_15_0_cry_1 ;
wire un1_x_15_0_axb_2 ;
wire un1_x_15_0_cry_2 ;
wire un1_x_15_0_axb_3 ;
wire un1_x_15_0_cry_3 ;
wire un1_x_15_0_axb_4 ;
wire un1_x_15_0_cry_4 ;
wire un1_x_15_0_axb_5 ;
wire un1_x_15_0_cry_5 ;
wire un1_x_15_0_axb_6 ;
wire un1_x_15_0_cry_6 ;
wire un1_x_15_0_axb_7 ;
wire un1_x_15_0_cry_7 ;
wire un1_x_15_0_axb_8 ;
wire un1_x_11_0_axb_0 ;
wire un1_x_11_0_cry_0 ;
wire un1_x_11_0_axb_1 ;
wire un1_x_11_0_cry_1 ;
wire un1_x_11_0_axb_2 ;
wire un1_x_11_0_cry_2 ;
wire un1_x_11_0_axb_3 ;
wire un1_x_11_0_cry_3 ;
wire un1_x_11_0_axb_4 ;
wire un1_x_11_0_cry_4 ;
wire un1_x_11_0_axb_5 ;
wire un1_x_11_0_cry_5 ;
wire un1_x_11_0_axb_6 ;
wire un1_x_11_0_cry_6 ;
wire un1_x_11_0_axb_7 ;
wire un1_x_11_0_cry_7 ;
wire un1_x_11_0_axb_8 ;
wire un1_x_16_0_axb_0 ;
wire un1_x_16_0_cry_0 ;
wire un1_x_16_0_axb_1 ;
wire un1_x_16_0_cry_1 ;
wire un1_x_16_0_axb_2 ;
wire un1_x_16_0_cry_2 ;
wire un1_x_16_0_axb_3 ;
wire un1_x_16_0_cry_3 ;
wire un1_x_16_0_axb_4 ;
wire un1_x_16_0_cry_4 ;
wire un1_x_16_0_axb_5 ;
wire un1_x_16_0_cry_5 ;
wire un1_x_16_0_axb_6 ;
wire un1_x_16_0_cry_6 ;
wire un1_x_16_0_axb_7 ;
wire un1_x_16_0_cry_7 ;
wire un1_x_16_0_axb_8 ;
wire un84_sop_0_0_0_1_cry_0 ;
wire un84_sop_0_0_0_1_axb_1 ;
wire un84_sop_0_0_0_1_cry_1 ;
wire un84_sop_0_0_0_1_axb_2 ;
wire un84_sop_0_0_0_1_cry_2 ;
wire un84_sop_0_0_0_1_axb_3 ;
wire un84_sop_0_0_0_1_cry_3 ;
wire un84_sop_0_0_0_1_axb_4 ;
wire un84_sop_0_0_0_1_cry_4 ;
wire un84_sop_0_0_0_1_axb_5 ;
wire un84_sop_0_0_0_1_cry_5 ;
wire un84_sop_0_0_0_1_axb_6 ;
wire un84_sop_0_0_0_1_cry_6 ;
wire un84_sop_0_0_0_1_axb_7 ;
wire un84_sop_0_0_0_1_cry_7 ;
wire un84_sop_0_0_0_1_axb_8 ;
wire un84_sop_0_0_0_1_cry_8 ;
wire un84_sop_0_0_0_1_axb_9 ;
wire un1_x_10_4_cry_1_sf ;
wire un84_sop_0_0_0_0_11_7_axb_0_ci ;
wire un84_sop_0_0_0_11_0_cry_0_cy ;
wire un84_sop_0_0_0_11_6_0_cry_0_cy ;
wire un84_sop_0_0_0_6_6_0_cry_0_cy ;
wire un84_sop_1_6_0_cry_0_cy ;
wire un84_sop_0_0_0_6_0_axb_0_0 ;
wire un84_sop_0_0_0_6_0_axb_0_1 ;
wire un84_sop_1_6_0_axb_0_0 ;
wire un1_x_10_4_s_8_false ;
wire x_4_x_4_1Q_Q31 ;
wire x_4_0_x_4_1Q_Q31 ;
wire x_4_1_x_4_1Q_Q31 ;
wire x_4_2_x_4_1Q_Q31 ;
wire x_4_3_x_4_1Q_Q31 ;
wire x_4_4_x_4_1Q_Q31 ;
wire x_4_5_x_4_1Q_Q31 ;
wire x_4_6_x_4_1Q_Q31 ;
wire x_7_x_7_1Q_Q31 ;
wire x_7_0_x_7_1Q_Q31 ;
wire x_7_1_x_7_1Q_Q31 ;
wire x_7_2_x_7_1Q_Q31 ;
wire x_7_3_x_7_1Q_Q31 ;
wire x_7_4_x_7_1Q_Q31 ;
wire x_7_5_x_7_1Q_Q31 ;
wire x_7_6_x_7_1Q_Q31 ;
wire x_12_x_4_1Q_Q31 ;
wire x_12_0_x_4_1Q_Q31 ;
wire x_12_1_x_4_1Q_Q31 ;
wire x_12_2_x_4_1Q_Q31 ;
wire x_12_3_x_4_1Q_Q31 ;
wire x_12_4_x_4_1Q_Q31 ;
wire x_12_5_x_4_1Q_Q31 ;
wire x_12_6_x_7_1Q_Q31 ;
input p_desc0_p_O_FD ;
input p_desc1_p_O_FD ;
input p_desc2_p_O_FD ;
input p_desc3_p_O_FD ;
input p_desc4_p_O_FD ;
input p_desc5_p_O_FD ;
input p_desc6_p_O_FD ;
input p_desc7_p_O_FD ;
input p_desc8_p_O_FD ;
input p_desc9_p_O_FD ;
input p_desc10_p_O_FD ;
input p_desc11_p_O_FD ;
input p_desc12_p_O_FD ;
input p_desc13_p_O_FD ;
input p_desc14_p_O_FD ;
input p_desc15_p_O_FD ;
input p_desc16_p_O_FD ;
input p_desc17_p_O_FD ;
input p_desc18_p_O_FD ;
input p_desc19_p_O_FD ;
input p_desc20_p_O_FD ;
input p_desc21_p_O_FD ;
input p_desc22_p_O_FD ;
input p_desc23_p_O_FD ;
input p_desc24_p_O_FD ;
input p_desc25_p_O_FD ;
input p_desc26_p_O_FD ;
input p_desc27_p_O_FD ;
input p_desc28_p_O_FD ;
input p_desc29_p_O_FD ;
input p_desc30_p_O_FD ;
input p_desc31_p_O_FD ;
input p_desc32_p_O_FD ;
input p_x_14_pipe_0_Z_p_O_FD ;
input p_x_14_pipe_9_Z_p_O_FD ;
input p_x_14_pipe_10_Z_p_O_FD ;
input p_x_14_pipe_11_Z_p_O_FD ;
input p_x_14_pipe_12_Z_p_O_FD ;
input p_x_14_pipe_13_Z_p_O_FD ;
input p_x_14_pipe_14_Z_p_O_FD ;
input p_x_14_pipe_15_Z_p_O_FD ;
input p_x_14_pipe_16_Z_p_O_FD ;
input p_x_14_pipe_17_Z_p_O_FD ;
input p_x_9_pipe_1_Z_p_O_FD ;
input p_x_9_pipe_2_Z_p_O_FD ;
input p_x_9_pipe_3_Z_p_O_FD ;
input p_x_9_pipe_4_Z_p_O_FD ;
input p_x_9_pipe_5_Z_p_O_FD ;
input p_x_9_pipe_6_Z_p_O_FD ;
input p_x_9_pipe_7_Z_p_O_FD ;
input p_x_9_pipe_8_Z_p_O_FD ;
input p_x_15_pipe_0_0_15_Z_p_O_FD ;
input p_x_15_pipe_0_0_16_Z_p_O_FD ;
input p_x_15_pipe_0_0_17_Z_p_O_FD ;
input p_x_15_pipe_0_0_18_Z_p_O_FD ;
input p_x_15_pipe_0_0_19_Z_p_O_FD ;
input p_x_15_pipe_0_0_20_Z_p_O_FD ;
input p_x_15_pipe_0_0_21_Z_p_O_FD ;
input p_x_15_pipe_0_0_22_Z_p_O_FD ;
input p_x_15_pipe_0_0_23_Z_p_O_FD ;
input p_x_15_pipe_0_0_24_Z_p_O_FD ;
input p_x_15_pipe_0_0_25_Z_p_O_FD ;
input p_x_15_pipe_0_0_26_Z_p_O_FD ;
input p_x_15_pipe_0_0_27_Z_p_O_FD ;
input p_x_15_pipe_0_0_28_Z_p_O_FD ;
input p_x_15_pipe_0_0_29_Z_p_O_FD ;
input p_x_16_pipe_0_0_0_Z_p_O_FD ;
input p_x_16_pipe_0_0_1_Z_p_O_FD ;
input p_x_16_pipe_0_0_2_Z_p_O_FD ;
input p_x_16_pipe_0_0_3_Z_p_O_FD ;
input p_x_16_pipe_0_0_4_Z_p_O_FD ;
input p_x_16_pipe_0_0_5_Z_p_O_FD ;
input p_x_16_pipe_0_0_6_Z_p_O_FD ;
input p_x_16_pipe_0_0_7_Z_p_O_FD ;
input p_x_16_pipe_0_0_8_Z_p_O_FD ;
input p_x_16_pipe_0_0_9_Z_p_O_FD ;
input p_x_16_pipe_0_0_10_Z_p_O_FD ;
input p_x_16_pipe_0_0_11_Z_p_O_FD ;
input p_x_16_pipe_0_0_12_Z_p_O_FD ;
input p_x_16_pipe_0_0_13_Z_p_O_FD ;
input p_x_16_pipe_0_0_14_Z_p_O_FD ;
input p_desc33_p_O_FD ;
input p_desc34_p_O_FD ;
input p_desc35_p_O_FD ;
input p_desc36_p_O_FD ;
input p_desc37_p_O_FD ;
input p_desc38_p_O_FD ;
input p_desc39_p_O_FD ;
input p_desc40_p_O_FD ;
input p_desc41_p_O_FD ;
input p_desc42_p_O_FD ;
input p_desc43_p_O_FD ;
input p_desc44_p_O_FD ;
input p_desc45_p_O_FD ;
input p_desc46_p_O_FD ;
input p_desc47_p_O_FD ;
input p_desc48_p_O_FD ;
input p_desc49_p_O_FD ;
input p_desc50_p_O_FD ;
input p_desc51_p_O_FD ;
input p_desc52_p_O_FD ;
input p_desc53_p_O_FD ;
input p_desc54_p_O_FD ;
input p_desc55_p_O_FD ;
input p_desc56_p_O_FD ;
// instances
  GND GND_cZ(.G(GND));
  VCC VCC_cZ(.P(VCC));
  SRLC32E x_12_6_x_7_1Q(.Q(x_12_6_tmp_d_array_0),.Q31(x_12_6_x_7_1Q_Q31),.A({GND,GND,GND,GND,VCC}),.D(x_9),.CLK(clk),.CE(VCC));
  SRLC32E x_12_5_x_4_1Q(.Q(x_12_5_tmp_d_array_0),.Q31(x_12_5_x_4_1Q_Q31),.A({GND,GND,GND,VCC,GND}),.D(x_8[1:1]),.CLK(clk),.CE(VCC));
  SRLC32E x_12_4_x_4_1Q(.Q(x_12_4_tmp_d_array_0),.Q31(x_12_4_x_4_1Q_Q31),.A({GND,GND,GND,VCC,GND}),.D(x_8[2:2]),.CLK(clk),.CE(VCC));
  SRLC32E x_12_3_x_4_1Q(.Q(x_12_3_tmp_d_array_0),.Q31(x_12_3_x_4_1Q_Q31),.A({GND,GND,GND,VCC,GND}),.D(x_8[3:3]),.CLK(clk),.CE(VCC));
  SRLC32E x_12_2_x_4_1Q(.Q(x_12_2_tmp_d_array_0),.Q31(x_12_2_x_4_1Q_Q31),.A({GND,GND,GND,VCC,GND}),.D(x_8[4:4]),.CLK(clk),.CE(VCC));
  SRLC32E x_12_1_x_4_1Q(.Q(x_12_1_tmp_d_array_0),.Q31(x_12_1_x_4_1Q_Q31),.A({GND,GND,GND,VCC,GND}),.D(x_8[5:5]),.CLK(clk),.CE(VCC));
  SRLC32E x_12_0_x_4_1Q(.Q(x_12_0_tmp_d_array_0),.Q31(x_12_0_x_4_1Q_Q31),.A({GND,GND,GND,VCC,GND}),.D(x_8[6:6]),.CLK(clk),.CE(VCC));
  SRLC32E x_12_x_4_1Q(.Q(x_12_tmp_d_array_0),.Q31(x_12_x_4_1Q_Q31),.A({GND,GND,GND,VCC,GND}),.D(x_8[7:7]),.CLK(clk),.CE(VCC));
  SRLC32E x_7_6_x_7_1Q(.Q(x_7_6_tmp_d_array_0),.Q31(x_7_6_x_7_1Q_Q31),.A({GND,GND,GND,GND,VCC}),.D(x_4[0:0]),.CLK(clk),.CE(VCC));
  SRLC32E x_7_5_x_7_1Q(.Q(x_7_5_tmp_d_array_0),.Q31(x_7_5_x_7_1Q_Q31),.A({GND,GND,GND,GND,VCC}),.D(x_4[1:1]),.CLK(clk),.CE(VCC));
  SRLC32E x_7_4_x_7_1Q(.Q(x_7_4_tmp_d_array_0),.Q31(x_7_4_x_7_1Q_Q31),.A({GND,GND,GND,GND,VCC}),.D(x_4[2:2]),.CLK(clk),.CE(VCC));
  SRLC32E x_7_3_x_7_1Q(.Q(x_7_3_tmp_d_array_0),.Q31(x_7_3_x_7_1Q_Q31),.A({GND,GND,GND,GND,VCC}),.D(x_4[3:3]),.CLK(clk),.CE(VCC));
  SRLC32E x_7_2_x_7_1Q(.Q(x_7_2_tmp_d_array_0),.Q31(x_7_2_x_7_1Q_Q31),.A({GND,GND,GND,GND,VCC}),.D(x_4[4:4]),.CLK(clk),.CE(VCC));
  SRLC32E x_7_1_x_7_1Q(.Q(x_7_1_tmp_d_array_0),.Q31(x_7_1_x_7_1Q_Q31),.A({GND,GND,GND,GND,VCC}),.D(x_4[5:5]),.CLK(clk),.CE(VCC));
  SRLC32E x_7_0_x_7_1Q(.Q(x_7_0_tmp_d_array_0),.Q31(x_7_0_x_7_1Q_Q31),.A({GND,GND,GND,GND,VCC}),.D(x_4[6:6]),.CLK(clk),.CE(VCC));
  SRLC32E x_7_x_7_1Q(.Q(x_7_tmp_d_array_0),.Q31(x_7_x_7_1Q_Q31),.A({GND,GND,GND,GND,VCC}),.D(x_4[7:7]),.CLK(clk),.CE(VCC));
  SRLC32E x_4_6_x_4_1Q(.Q(x_4_6_tmp_d_array_0),.Q31(x_4_6_x_4_1Q_Q31),.A({GND,GND,GND,VCC,GND}),.D(x_0[0:0]),.CLK(clk),.CE(VCC));
  SRLC32E x_4_5_x_4_1Q(.Q(x_4_5_tmp_d_array_0),.Q31(x_4_5_x_4_1Q_Q31),.A({GND,GND,GND,VCC,GND}),.D(x_0[1:1]),.CLK(clk),.CE(VCC));
  SRLC32E x_4_4_x_4_1Q(.Q(x_4_4_tmp_d_array_0),.Q31(x_4_4_x_4_1Q_Q31),.A({GND,GND,GND,VCC,GND}),.D(x_0[2:2]),.CLK(clk),.CE(VCC));
  SRLC32E x_4_3_x_4_1Q(.Q(x_4_3_tmp_d_array_0),.Q31(x_4_3_x_4_1Q_Q31),.A({GND,GND,GND,VCC,GND}),.D(x_0[3:3]),.CLK(clk),.CE(VCC));
  SRLC32E x_4_2_x_4_1Q(.Q(x_4_2_tmp_d_array_0),.Q31(x_4_2_x_4_1Q_Q31),.A({GND,GND,GND,VCC,GND}),.D(x_0[4:4]),.CLK(clk),.CE(VCC));
  SRLC32E x_4_1_x_4_1Q(.Q(x_4_1_tmp_d_array_0),.Q31(x_4_1_x_4_1Q_Q31),.A({GND,GND,GND,VCC,GND}),.D(x_0[5:5]),.CLK(clk),.CE(VCC));
  SRLC32E x_4_0_x_4_1Q(.Q(x_4_0_tmp_d_array_0),.Q31(x_4_0_x_4_1Q_Q31),.A({GND,GND,GND,VCC,GND}),.D(x_0[6:6]),.CLK(clk),.CE(VCC));
  SRLC32E x_4_x_4_1Q(.Q(x_4_tmp_d_array_0),.Q31(x_4_x_4_1Q_Q31),.A({GND,GND,GND,VCC,GND}),.D(x_0[7:7]),.CLK(clk),.CE(VCC));
  LUT1 un1_x_10_4_s_8_false_cZ(.I0(GND),.O(un1_x_10_4_s_8_false));
defparam un1_x_10_4_s_8_false_cZ.INIT=2'h0;
  LUT3 un84_sop_1_6_0_s_0_lut(.I0(un1_x_1[4:4]),.I1(un1_x_2[5:5]),.I2(un1_x_3[4:4]),.O(un84_sop_1_6[0:0]));
defparam un84_sop_1_6_0_s_0_lut.INIT=8'h96;
  LUT3 un84_sop_0_0_0_11_6_0_s_0_lut(.I0(un1_x_12_0_0[4:4]),.I1(un1_x_13_0_0[5:5]),.I2(un1_x_14_0_0[4:4]),.O(un84_sop_0_0_0_0_11_6[0:0]));
defparam un84_sop_0_0_0_11_6_0_s_0_lut.INIT=8'h96;
  LUT3 un84_sop_0_0_0_6_6_0_s_0_lut(.I0(un1_x_7_0[2:2]),.I1(un1_x_8_0[4:4]),.I2(un1_x_9_0[5:5]),.O(un84_sop_0_0_0_1_6_6[0:0]));
defparam un84_sop_0_0_0_6_6_0_s_0_lut.INIT=8'h96;
  LUT2 un84_sop_0_0_0_6_0_axb_0_0_cZ(.I0(un1_x_12_0_0[4:4]),.I1(un1_x_13_0_0[5:5]),.O(un84_sop_0_0_0_6_0_axb_0_0));
defparam un84_sop_0_0_0_6_0_axb_0_0_cZ.INIT=4'h6;
  LUT3 un84_sop_0_0_0_11_6_0_axb_12_cZ(.I0(un1_x_12_0_0[15:15]),.I1(un1_x_13_0_0[15:15]),.I2(un1_x_14_0_0[15:15]),.O(un84_sop_0_0_0_11_6_0_axb_12));
defparam un84_sop_0_0_0_11_6_0_axb_12_cZ.INIT=8'h7E;
  LUT2 un84_sop_0_0_0_6_0_axb_0_1_cZ(.I0(un1_x_7_0[2:2]),.I1(un1_x_8_0[4:4]),.O(un84_sop_0_0_0_6_0_axb_0_1));
defparam un84_sop_0_0_0_6_0_axb_0_1_cZ.INIT=4'h6;
  LUT4 un84_sop_0_0_0_6_6_0_axb_12_cZ(.I0(un1_x_7_0[13:13]),.I1(un1_x_7_0[14:14]),.I2(un1_x_8_0[15:15]),.I3(un1_x_9_0[15:15]),.O(un84_sop_0_0_0_6_6_0_axb_12));
defparam un84_sop_0_0_0_6_6_0_axb_12_cZ.INIT=16'h399C;
  LUT4 un84_sop_0_0_0_6_6_0_axb_13_cZ(.I0(un1_x_7_0[14:14]),.I1(un1_x_7_0[15:15]),.I2(un1_x_8_0[15:15]),.I3(un1_x_9_0[15:15]),.O(un84_sop_0_0_0_6_6_0_axb_13));
defparam un84_sop_0_0_0_6_6_0_axb_13_cZ.INIT=16'h399C;
  LUT2 un84_sop_0_0_0_1_6_8_axb_0(.I0(un84_sop_0_0_0_10_0[3:3]),.I1(x_4[0:0]),.O(un84_sop_0_0_0_1_6_8[3:3]));
defparam un84_sop_0_0_0_1_6_8_axb_0.INIT=4'h6;
  LUT2 un84_sop_0_0_0_1_6_8_axb_1_cZ(.I0(un84_sop_0_0_0_10_0[4:4]),.I1(x_4[1:1]),.O(un84_sop_0_0_0_1_6_8_axb_1));
defparam un84_sop_0_0_0_1_6_8_axb_1_cZ.INIT=4'h6;
  LUT4 un84_sop_0_0_0_1_6_8_axb_9_cZ(.I0(un84_sop_0_0_0_10_0[11:11]),.I1(un84_sop_0_0_0_10_0[12:12]),.I2(x_4[6:6]),.I3(x_4[7:7]),.O(un84_sop_0_0_0_1_6_8_axb_9));
defparam un84_sop_0_0_0_1_6_8_axb_9_cZ.INIT=16'h366C;
  LUT2 un84_sop_0_0_0_1_6_8_axb_10_cZ(.I0(un84_sop_0_0_0_10_0[13:13]),.I1(x_4[7:7]),.O(un84_sop_0_0_0_1_6_8_axb_10));
defparam un84_sop_0_0_0_1_6_8_axb_10_cZ.INIT=4'h6;
  LUT2 un84_sop_1_6_0_axb_0_0_cZ(.I0(un1_x_1[4:4]),.I1(un1_x_2[5:5]),.O(un84_sop_1_6_0_axb_0_0));
defparam un84_sop_1_6_0_axb_0_0_cZ.INIT=4'h6;
  LUT3 un84_sop_1_6_0_axb_12_cZ(.I0(un1_x_1[15:15]),.I1(un1_x_2[15:15]),.I2(un1_x_3[15:15]),.O(un84_sop_1_6_0_axb_12));
defparam un84_sop_1_6_0_axb_12_cZ.INIT=8'h7E;
  LUT3 un1_x_10_axb_4_cZ(.I0(un1_x_10_4[4:4]),.I1(x_8[0:0]),.I2(x_8[1:1]),.O(un1_x_10_axb_4));
defparam un1_x_10_axb_4_cZ.INIT=8'h96;
  LUT4 un1_x_10_axb_5_cZ(.I0(un1_x_10_4[5:5]),.I1(x_8[0:0]),.I2(x_8[1:1]),.I3(x_8[2:2]),.O(un1_x_10_axb_5));
defparam un1_x_10_axb_5_cZ.INIT=16'hA956;
  LUT3 un1_x_10_axb_8_cZ(.I0(un1_x_10_4[8:8]),.I1(un1_x_10_5_c5),.I2(x_8[5:5]),.O(un1_x_10_axb_8));
defparam un1_x_10_axb_8_cZ.INIT=8'h69;
  LUT4 un1_x_10_axb_9_cZ(.I0(un1_x_10_5_c5),.I1(x_8[5:5]),.I2(x_8[6:6]),.I3(x_8[7:7]),.O(un1_x_10_axb_9));
defparam un1_x_10_axb_9_cZ.INIT=16'hD22D;
  LUT3 un1_x_10_axb_10_cZ(.I0(un1_x_10_5_c5),.I1(x_8[5:5]),.I2(x_8[6:6]),.O(un1_x_10_axb_10));
defparam un1_x_10_axb_10_cZ.INIT=8'hFD;
  LUT2 un84_sop_0_0_0_1_6_4_axb_0(.I0(un1_x_6_0[1:1]),.I1(un84_sop_0_0_0_10_0[0:0]),.O(un84_sop_0_0_0_1_6_4[0:0]));
defparam un84_sop_0_0_0_1_6_4_axb_0.INIT=4'h6;
  LUT2 un84_sop_0_0_0_1_6_4_axb_1_cZ(.I0(un1_x_6_0[2:2]),.I1(un84_sop_0_0_0_10_0[1:1]),.O(un84_sop_0_0_0_1_6_4_axb_1));
defparam un84_sop_0_0_0_1_6_4_axb_1_cZ.INIT=4'h6;
  LUT2 un84_sop_0_0_0_1_6_4_axb_2_cZ(.I0(un1_x_6_0[3:3]),.I1(un84_sop_0_0_0_10_0[2:2]),.O(un84_sop_0_0_0_1_6_4_axb_2));
defparam un84_sop_0_0_0_1_6_4_axb_2_cZ.INIT=4'h6;
  LUT3 un84_sop_0_0_0_1_6_4_axb_3_cZ(.I0(un1_x_6_0[4:4]),.I1(un84_sop_0_0_0_10_0[3:3]),.I2(x_4[0:0]),.O(un84_sop_0_0_0_1_6_4_axb_3));
defparam un84_sop_0_0_0_1_6_4_axb_3_cZ.INIT=8'h96;
  LUT2 un84_sop_0_0_0_1_6_4_axb_4_cZ(.I0(un1_x_6_0[5:5]),.I1(un84_sop_0_0_0_1_6_8[4:4]),.O(un84_sop_0_0_0_1_6_4_axb_4));
defparam un84_sop_0_0_0_1_6_4_axb_4_cZ.INIT=4'h6;
  LUT2 un84_sop_0_0_0_1_6_4_axb_5_cZ(.I0(un1_x_6_0[6:6]),.I1(un84_sop_0_0_0_1_6_8[5:5]),.O(un84_sop_0_0_0_1_6_4_axb_5));
defparam un84_sop_0_0_0_1_6_4_axb_5_cZ.INIT=4'h6;
  LUT2 un84_sop_0_0_0_1_6_4_axb_6_cZ(.I0(un1_x_6_0[7:7]),.I1(un84_sop_0_0_0_1_6_8[6:6]),.O(un84_sop_0_0_0_1_6_4_axb_6));
defparam un84_sop_0_0_0_1_6_4_axb_6_cZ.INIT=4'h6;
  LUT2 un84_sop_0_0_0_1_6_4_axb_7_cZ(.I0(un1_x_6_0[8:8]),.I1(un84_sop_0_0_0_1_6_8[7:7]),.O(un84_sop_0_0_0_1_6_4_axb_7));
defparam un84_sop_0_0_0_1_6_4_axb_7_cZ.INIT=4'h6;
  LUT2 un84_sop_0_0_0_1_6_4_axb_8_cZ(.I0(un1_x_6_0[9:9]),.I1(un84_sop_0_0_0_1_6_8[8:8]),.O(un84_sop_0_0_0_1_6_4_axb_8));
defparam un84_sop_0_0_0_1_6_4_axb_8_cZ.INIT=4'h6;
  LUT2 un84_sop_0_0_0_1_6_4_axb_9_cZ(.I0(un1_x_6_0[10:10]),.I1(un84_sop_0_0_0_1_6_8[9:9]),.O(un84_sop_0_0_0_1_6_4_axb_9));
defparam un84_sop_0_0_0_1_6_4_axb_9_cZ.INIT=4'h6;
  LUT2 un84_sop_0_0_0_1_6_4_axb_10_cZ(.I0(un1_x_6_0[11:11]),.I1(un84_sop_0_0_0_1_6_8[10:10]),.O(un84_sop_0_0_0_1_6_4_axb_10));
defparam un84_sop_0_0_0_1_6_4_axb_10_cZ.INIT=4'h6;
  LUT2 un84_sop_0_0_0_1_6_4_axb_11_cZ(.I0(un1_x_6_0[12:12]),.I1(un84_sop_0_0_0_1_6_8[11:11]),.O(un84_sop_0_0_0_1_6_4_axb_11));
defparam un84_sop_0_0_0_1_6_4_axb_11_cZ.INIT=4'h6;
  LUT2 un84_sop_0_0_0_1_6_4_axb_12_cZ(.I0(un1_x_6_0[13:13]),.I1(un84_sop_0_0_0_1_6_8[12:12]),.O(un84_sop_0_0_0_1_6_4_axb_12));
defparam un84_sop_0_0_0_1_6_4_axb_12_cZ.INIT=4'h6;
  LUT2 un84_sop_0_0_0_1_6_4_axb_13_cZ(.I0(un1_x_6_0[14:14]),.I1(un84_sop_0_0_0_1_6_8[13:13]),.O(un84_sop_0_0_0_1_6_4_axb_13));
defparam un84_sop_0_0_0_1_6_4_axb_13_cZ.INIT=4'h6;
  LUT2 un84_sop_1_7_axb_1_cZ(.I0(un1_x_4[3:3]),.I1(un84_sop_0_0_0_0_5[1:1]),.O(un84_sop_1_7_axb_1));
defparam un84_sop_1_7_axb_1_cZ.INIT=4'h6;
  LUT2 un84_sop_1_7_axb_2_cZ(.I0(un1_x_4[4:4]),.I1(un84_sop_0_0_0_0_5[2:2]),.O(un84_sop_1_7_axb_2));
defparam un84_sop_1_7_axb_2_cZ.INIT=4'h6;
  LUT2 un84_sop_1_7_axb_3_cZ(.I0(un1_x_4[5:5]),.I1(un84_sop_0_0_0_0_5[3:3]),.O(un84_sop_1_7_axb_3));
defparam un84_sop_1_7_axb_3_cZ.INIT=4'h6;
  LUT2 un84_sop_1_7_axb_4_cZ(.I0(un1_x_4[6:6]),.I1(un84_sop_0_0_0_0_5[4:4]),.O(un84_sop_1_7_axb_4));
defparam un84_sop_1_7_axb_4_cZ.INIT=4'h6;
  LUT2 un84_sop_1_7_axb_5_cZ(.I0(un1_x_4[7:7]),.I1(un84_sop_0_0_0_0_5[5:5]),.O(un84_sop_1_7_axb_5));
defparam un84_sop_1_7_axb_5_cZ.INIT=4'h6;
  LUT2 un84_sop_1_7_axb_6_cZ(.I0(un1_x_4[8:8]),.I1(un84_sop_0_0_0_0_5[6:6]),.O(un84_sop_1_7_axb_6));
defparam un84_sop_1_7_axb_6_cZ.INIT=4'h6;
  LUT2 un84_sop_1_7_axb_7_cZ(.I0(un1_x_4[9:9]),.I1(un84_sop_0_0_0_0_5[7:7]),.O(un84_sop_1_7_axb_7));
defparam un84_sop_1_7_axb_7_cZ.INIT=4'h6;
  LUT2 un84_sop_1_7_axb_8_cZ(.I0(un1_x_4[10:10]),.I1(un84_sop_0_0_0_0_5[8:8]),.O(un84_sop_1_7_axb_8));
defparam un84_sop_1_7_axb_8_cZ.INIT=4'h6;
  LUT2 un84_sop_1_7_axb_9_cZ(.I0(un1_x_4[11:11]),.I1(un84_sop_0_0_0_0_5[9:9]),.O(un84_sop_1_7_axb_9));
defparam un84_sop_1_7_axb_9_cZ.INIT=4'h6;
  LUT2 un84_sop_1_7_axb_10_cZ(.I0(un1_x_4[12:12]),.I1(un84_sop_0_0_0_0_5[10:10]),.O(un84_sop_1_7_axb_10));
defparam un84_sop_1_7_axb_10_cZ.INIT=4'h6;
  LUT2 un84_sop_1_7_axb_11_cZ(.I0(un1_x_4[13:13]),.I1(un84_sop_0_0_0_0_5[11:11]),.O(un84_sop_1_7_axb_11));
defparam un84_sop_1_7_axb_11_cZ.INIT=4'h6;
  LUT2 un84_sop_1_7_axb_12_cZ(.I0(un1_x_4[14:14]),.I1(un84_sop_0_0_0_0_5[12:12]),.O(un84_sop_1_7_axb_12));
defparam un84_sop_1_7_axb_12_cZ.INIT=4'h6;
  LUT2 un84_sop_1_7_axb_13_cZ(.I0(un1_x_4[15:15]),.I1(un84_sop_0_0_0_0_5[13:13]),.O(un84_sop_1_7_axb_13));
defparam un84_sop_1_7_axb_13_cZ.INIT=4'h6;
  LUT2 un84_sop_0_0_0_0_11_7_axb_0(.I0(un84_sop_0_0_0_0_0[0:0]),.I1(x_9),.O(un84_sop_0_0_0_0_11_7[0:0]));
defparam un84_sop_0_0_0_0_11_7_axb_0.INIT=4'h6;
  LUT2 un84_sop_0_0_0_0_11_7_axb_1_cZ(.I0(un1_x_11_0_0[7:7]),.I1(un84_sop_0_0_0_0_0[1:1]),.O(un84_sop_0_0_0_0_11_7_axb_1));
defparam un84_sop_0_0_0_0_11_7_axb_1_cZ.INIT=4'h6;
  LUT2 un84_sop_0_0_0_0_11_7_axb_2_cZ(.I0(un1_x_11_0_0[8:8]),.I1(un84_sop_0_0_0_0_0[2:2]),.O(un84_sop_0_0_0_0_11_7_axb_2));
defparam un84_sop_0_0_0_0_11_7_axb_2_cZ.INIT=4'h6;
  LUT2 un84_sop_0_0_0_0_11_7_axb_3_cZ(.I0(un1_x_11_0_0[9:9]),.I1(un84_sop_0_0_0_0_0[3:3]),.O(un84_sop_0_0_0_0_11_7_axb_3));
defparam un84_sop_0_0_0_0_11_7_axb_3_cZ.INIT=4'h6;
  LUT2 un84_sop_0_0_0_0_11_7_axb_4_cZ(.I0(un1_x_11_0_0[10:10]),.I1(un84_sop_0_0_0_0_0[4:4]),.O(un84_sop_0_0_0_0_11_7_axb_4));
defparam un84_sop_0_0_0_0_11_7_axb_4_cZ.INIT=4'h6;
  LUT2 un84_sop_0_0_0_0_11_7_axb_5_cZ(.I0(un1_x_11_0_0[11:11]),.I1(un84_sop_0_0_0_0_0[5:5]),.O(un84_sop_0_0_0_0_11_7_axb_5));
defparam un84_sop_0_0_0_0_11_7_axb_5_cZ.INIT=4'h6;
  LUT2 un84_sop_0_0_0_0_11_7_axb_6_cZ(.I0(un1_x_11_0_0[12:12]),.I1(un84_sop_0_0_0_0_0[6:6]),.O(un84_sop_0_0_0_0_11_7_axb_6));
defparam un84_sop_0_0_0_0_11_7_axb_6_cZ.INIT=4'h6;
  LUT2 un84_sop_0_0_0_0_11_7_axb_7_cZ(.I0(un1_x_11_0_0[13:13]),.I1(un84_sop_0_0_0_0_0[7:7]),.O(un84_sop_0_0_0_0_11_7_axb_7));
defparam un84_sop_0_0_0_0_11_7_axb_7_cZ.INIT=4'h6;
  LUT2 un84_sop_0_0_0_0_11_7_axb_8_cZ(.I0(un1_x_11_0_0[14:14]),.I1(un84_sop_0_0_0_0_0[8:8]),.O(un84_sop_0_0_0_0_11_7_axb_8));
defparam un84_sop_0_0_0_0_11_7_axb_8_cZ.INIT=4'h6;
  LUT2 un84_sop_0_0_0_0_11_7_axb_9_cZ(.I0(un1_x_11_0_0[14:14]),.I1(un84_sop_0_0_0_0_0[9:9]),.O(un84_sop_0_0_0_0_11_7_axb_9));
defparam un84_sop_0_0_0_0_11_7_axb_9_cZ.INIT=4'h6;
  LUT3 un84_sop_1_4_cry_0_RNO(.I0(un1_x_4[2:2]),.I1(un84_sop_0_0_0_0_5[0:0]),.I2(x_0[0:0]),.O(un84_sop_1_4[0:0]));
defparam un84_sop_1_4_cry_0_RNO.INIT=8'h96;
  LUT3 un84_sop_1_4_axb_1_cZ(.I0(un84_sop_1_7[1:1]),.I1(x_0[0:0]),.I2(x_0[1:1]),.O(un84_sop_1_4_axb_1));
defparam un84_sop_1_4_axb_1_cZ.INIT=8'h96;
  LUT4 un84_sop_1_4_axb_2_cZ(.I0(un84_sop_1_7[2:2]),.I1(x_0[0:0]),.I2(x_0[1:1]),.I3(x_0[2:2]),.O(un84_sop_1_4_axb_2));
defparam un84_sop_1_4_axb_2_cZ.INIT=16'hA956;
  LUT4 un84_sop_1_4_axb_5_cZ(.I0(un1_x_0_0_c4),.I1(un84_sop_1_7[5:5]),.I2(x_0[4:4]),.I3(x_0[5:5]),.O(un84_sop_1_4_axb_5));
defparam un84_sop_1_4_axb_5_cZ.INIT=16'hC639;
  LUT4 un84_sop_1_axb_0_cZ(.I0(un1_x_4[2:2]),.I1(un84_sop_0_0_0_0_5[0:0]),.I2(un84_sop_1_6[0:0]),.I3(x_0[0:0]),.O(un84_sop_1_axb_0));
defparam un84_sop_1_axb_0_cZ.INIT=16'h6996;
  LUT2 un84_sop_1_axb_1_cZ(.I0(un84_sop_1_4[1:1]),.I1(un84_sop_1_6[1:1]),.O(un84_sop_1_axb_1));
defparam un84_sop_1_axb_1_cZ.INIT=4'h6;
  LUT2 un84_sop_1_axb_2_cZ(.I0(un84_sop_1_4[2:2]),.I1(un84_sop_1_6[2:2]),.O(un84_sop_1_axb_2));
defparam un84_sop_1_axb_2_cZ.INIT=4'h6;
  LUT2 un84_sop_1_axb_3_cZ(.I0(un84_sop_1_4[3:3]),.I1(un84_sop_1_6[3:3]),.O(un84_sop_1_axb_3));
defparam un84_sop_1_axb_3_cZ.INIT=4'h6;
  LUT2 un84_sop_1_axb_4_cZ(.I0(un84_sop_1_4[4:4]),.I1(un84_sop_1_6[4:4]),.O(un84_sop_1_axb_4));
defparam un84_sop_1_axb_4_cZ.INIT=4'h6;
  LUT2 un84_sop_1_axb_5_cZ(.I0(un84_sop_1_4[5:5]),.I1(un84_sop_1_6[5:5]),.O(un84_sop_1_axb_5));
defparam un84_sop_1_axb_5_cZ.INIT=4'h6;
  LUT2 un84_sop_1_axb_6_cZ(.I0(un84_sop_1_4[6:6]),.I1(un84_sop_1_6[6:6]),.O(un84_sop_1_axb_6));
defparam un84_sop_1_axb_6_cZ.INIT=4'h6;
  LUT2 un1_x_10_4_cry_1_RNO(.I0(x_8[0:0]),.I1(x_8[1:1]),.O(un1_x_10_4_cry_1_sf));
defparam un1_x_10_4_cry_1_RNO.INIT=4'h6;
  LUT2 un1_x_10_4_axb_2_cZ(.I0(x_8[1:1]),.I1(x_8[2:2]),.O(un1_x_10_4_axb_2));
defparam un1_x_10_4_axb_2_cZ.INIT=4'h6;
  LUT2 un1_x_10_4_axb_3_cZ(.I0(x_8[2:2]),.I1(x_8[3:3]),.O(un1_x_10_4_axb_3));
defparam un1_x_10_4_axb_3_cZ.INIT=4'h6;
  LUT2 un1_x_10_4_axb_4_cZ(.I0(x_8[3:3]),.I1(x_8[4:4]),.O(un1_x_10_4_axb_4));
defparam un1_x_10_4_axb_4_cZ.INIT=4'h6;
  LUT2 un1_x_10_4_axb_5_cZ(.I0(x_8[4:4]),.I1(x_8[5:5]),.O(un1_x_10_4_axb_5));
defparam un1_x_10_4_axb_5_cZ.INIT=4'h6;
  LUT2 un1_x_10_4_axb_6_cZ(.I0(x_8[5:5]),.I1(x_8[6:6]),.O(un1_x_10_4_axb_6));
defparam un1_x_10_4_axb_6_cZ.INIT=4'h6;
  LUT2 un1_x_10_4_axb_7_cZ(.I0(x_8[6:6]),.I1(x_8[7:7]),.O(un1_x_10_4_axb_7));
defparam un1_x_10_4_axb_7_cZ.INIT=4'h6;
  LUT1 un1_x_15_0_axb_0_cZ(.I0(x_12[0:0]),.O(un1_x_15_0_axb_0));
defparam un1_x_15_0_axb_0_cZ.INIT=2'h1;
  LUT1 un1_x_15_0_axb_1_cZ(.I0(x_12[1:1]),.O(un1_x_15_0_axb_1));
defparam un1_x_15_0_axb_1_cZ.INIT=2'h1;
  LUT1 un1_x_15_0_axb_2_cZ(.I0(x_12[2:2]),.O(un1_x_15_0_axb_2));
defparam un1_x_15_0_axb_2_cZ.INIT=2'h1;
  LUT1 un1_x_15_0_axb_3_cZ(.I0(x_12[3:3]),.O(un1_x_15_0_axb_3));
defparam un1_x_15_0_axb_3_cZ.INIT=2'h1;
  LUT1 un1_x_15_0_axb_4_cZ(.I0(x_12[4:4]),.O(un1_x_15_0_axb_4));
defparam un1_x_15_0_axb_4_cZ.INIT=2'h1;
  LUT1 un1_x_15_0_axb_5_cZ(.I0(x_12[5:5]),.O(un1_x_15_0_axb_5));
defparam un1_x_15_0_axb_5_cZ.INIT=2'h1;
  LUT1 un1_x_15_0_axb_6_cZ(.I0(x_12[6:6]),.O(un1_x_15_0_axb_6));
defparam un1_x_15_0_axb_6_cZ.INIT=2'h1;
  LUT1 un1_x_15_0_axb_7_cZ(.I0(x_12[7:7]),.O(un1_x_15_0_axb_7));
defparam un1_x_15_0_axb_7_cZ.INIT=2'h1;
  LUT1 un1_x_11_0_axb_0_cZ(.I0(x_8[0:0]),.O(un1_x_11_0_axb_0));
defparam un1_x_11_0_axb_0_cZ.INIT=2'h1;
  LUT1 un1_x_16_0_axb_0_cZ(.I0(x_13[0:0]),.O(un1_x_16_0_axb_0));
defparam un1_x_16_0_axb_0_cZ.INIT=2'h1;
  LUT1 un1_x_16_0_axb_1_cZ(.I0(x_13[1:1]),.O(un1_x_16_0_axb_1));
defparam un1_x_16_0_axb_1_cZ.INIT=2'h1;
  LUT1 un1_x_16_0_axb_2_cZ(.I0(x_13[2:2]),.O(un1_x_16_0_axb_2));
defparam un1_x_16_0_axb_2_cZ.INIT=2'h1;
  LUT1 un1_x_16_0_axb_3_cZ(.I0(x_13[3:3]),.O(un1_x_16_0_axb_3));
defparam un1_x_16_0_axb_3_cZ.INIT=2'h1;
  LUT1 un1_x_16_0_axb_4_cZ(.I0(x_13[4:4]),.O(un1_x_16_0_axb_4));
defparam un1_x_16_0_axb_4_cZ.INIT=2'h1;
  LUT1 un1_x_16_0_axb_5_cZ(.I0(x_13[5:5]),.O(un1_x_16_0_axb_5));
defparam un1_x_16_0_axb_5_cZ.INIT=2'h1;
  LUT1 un1_x_16_0_axb_6_cZ(.I0(x_13[6:6]),.O(un1_x_16_0_axb_6));
defparam un1_x_16_0_axb_6_cZ.INIT=2'h1;
  LUT1 un1_x_16_0_axb_7_cZ(.I0(x_13[7:7]),.O(un1_x_16_0_axb_7));
defparam un1_x_16_0_axb_7_cZ.INIT=2'h1;
  LUT2 un84_sop_0_0_0_0_11_7_axb_0_ci_cZ(.I0(un84_sop_0_0_0_0_0[0:0]),.I1(x_9),.O(un84_sop_0_0_0_0_11_7_axb_0_ci));
defparam un84_sop_0_0_0_0_11_7_axb_0_ci_cZ.INIT=4'h6;
  LUT1 un84_sop_0_0_0_11_6_0_cry_0_thru(.I0(un1_x_14_0_0[4:4]),.O(un1_x_14_0_0_0[4:4]));
defparam un84_sop_0_0_0_11_6_0_cry_0_thru.INIT=2'h2;
  LUT1 un84_sop_0_0_0_6_6_0_cry_0_thru(.I0(un1_x_9_0[5:5]),.O(un1_x_9_0_0[5:5]));
defparam un84_sop_0_0_0_6_6_0_cry_0_thru.INIT=2'h2;
  LUT1 un84_sop_1_6_0_cry_0_thru(.I0(un1_x_3[4:4]),.O(un1_x_3_0[4:4]));
defparam un84_sop_1_6_0_cry_0_thru.INIT=2'h2;
  p_O_FD desc0(.Q(x_0[0:0]),.D(x_in[0:0]),.C(clk),.E(p_desc0_p_O_FD));
  p_O_FD desc1(.Q(x_0[1:1]),.D(x_in[1:1]),.C(clk),.E(p_desc1_p_O_FD));
  p_O_FD desc2(.Q(x_0[2:2]),.D(x_in[2:2]),.C(clk),.E(p_desc2_p_O_FD));
  p_O_FD desc3(.Q(x_0[3:3]),.D(x_in[3:3]),.C(clk),.E(p_desc3_p_O_FD));
  p_O_FD desc4(.Q(x_0[4:4]),.D(x_in[4:4]),.C(clk),.E(p_desc4_p_O_FD));
  p_O_FD desc5(.Q(x_0[5:5]),.D(x_in[5:5]),.C(clk),.E(p_desc5_p_O_FD));
  p_O_FD desc6(.Q(x_0[6:6]),.D(x_in[6:6]),.C(clk),.E(p_desc6_p_O_FD));
  p_O_FD desc7(.Q(x_0[7:7]),.D(x_in[7:7]),.C(clk),.E(p_desc7_p_O_FD));
  p_O_FD desc8(.Q(y[7:7]),.D(un84_sop_1_s_14),.C(clk),.E(p_desc8_p_O_FD));
  p_O_FD desc9(.Q(y[0:0]),.D(un84_sop_1_s_7),.C(clk),.E(p_desc9_p_O_FD));
  p_O_FD desc10(.Q(y[1:1]),.D(un84_sop_1_s_8),.C(clk),.E(p_desc10_p_O_FD));
  p_O_FD desc11(.Q(y[2:2]),.D(un84_sop_1_s_9),.C(clk),.E(p_desc11_p_O_FD));
  p_O_FD desc12(.Q(y[3:3]),.D(un84_sop_1_s_10),.C(clk),.E(p_desc12_p_O_FD));
  p_O_FD desc13(.Q(y[4:4]),.D(un84_sop_1_s_11),.C(clk),.E(p_desc13_p_O_FD));
  p_O_FD desc14(.Q(y[5:5]),.D(un84_sop_1_s_12),.C(clk),.E(p_desc14_p_O_FD));
  p_O_FD desc15(.Q(y[6:6]),.D(un84_sop_1_s_13),.C(clk),.E(p_desc15_p_O_FD));
  p_O_FD desc16(.Q(x_8[7:7]),.D(x_7[7:7]),.C(clk),.E(p_desc16_p_O_FD));
  p_O_FD desc17(.Q(x_8[6:6]),.D(x_7[6:6]),.C(clk),.E(p_desc17_p_O_FD));
  p_O_FD desc18(.Q(x_8[5:5]),.D(x_7[5:5]),.C(clk),.E(p_desc18_p_O_FD));
  p_O_FD desc19(.Q(x_8[4:4]),.D(x_7[4:4]),.C(clk),.E(p_desc19_p_O_FD));
  p_O_FD desc20(.Q(x_8[3:3]),.D(x_7[3:3]),.C(clk),.E(p_desc20_p_O_FD));
  p_O_FD desc21(.Q(x_8[2:2]),.D(x_7[2:2]),.C(clk),.E(p_desc21_p_O_FD));
  p_O_FD desc22(.Q(x_8[1:1]),.D(x_7[1:1]),.C(clk),.E(p_desc22_p_O_FD));
  p_O_FD desc23(.Q(x_8[0:0]),.D(x_7[0:0]),.C(clk),.E(p_desc23_p_O_FD));
  p_O_FD desc24(.Q(x_9),.D(x_8[0:0]),.C(clk),.E(p_desc24_p_O_FD));
  p_O_FD desc25(.Q(x_13[7:7]),.D(x_12[7:7]),.C(clk),.E(p_desc25_p_O_FD));
  p_O_FD desc26(.Q(x_13[6:6]),.D(x_12[6:6]),.C(clk),.E(p_desc26_p_O_FD));
  p_O_FD desc27(.Q(x_13[5:5]),.D(x_12[5:5]),.C(clk),.E(p_desc27_p_O_FD));
  p_O_FD desc28(.Q(x_13[4:4]),.D(x_12[4:4]),.C(clk),.E(p_desc28_p_O_FD));
  p_O_FD desc29(.Q(x_13[3:3]),.D(x_12[3:3]),.C(clk),.E(p_desc29_p_O_FD));
  p_O_FD desc30(.Q(x_13[2:2]),.D(x_12[2:2]),.C(clk),.E(p_desc30_p_O_FD));
  p_O_FD desc31(.Q(x_13[1:1]),.D(x_12[1:1]),.C(clk),.E(p_desc31_p_O_FD));
  p_O_FD desc32(.Q(x_13[0:0]),.D(x_12[0:0]),.C(clk),.E(p_desc32_p_O_FD));
  p_O_FD x_14_pipe_0_Z(.Q(un84_sop_0_0_0_0_0[0:0]),.D(un84_sop_0_0_0_0_1[0:0]),.C(clk),.E(p_x_14_pipe_0_Z_p_O_FD));
  p_O_FD x_14_pipe_9_Z(.Q(un84_sop_0_0_0_0_0[1:1]),.D(un84_sop_0_0_0_0_1[1:1]),.C(clk),.E(p_x_14_pipe_9_Z_p_O_FD));
  p_O_FD x_14_pipe_10_Z(.Q(un84_sop_0_0_0_0_0[2:2]),.D(un84_sop_0_0_0_0_1[2:2]),.C(clk),.E(p_x_14_pipe_10_Z_p_O_FD));
  p_O_FD x_14_pipe_11_Z(.Q(un84_sop_0_0_0_0_0[3:3]),.D(un84_sop_0_0_0_0_1[3:3]),.C(clk),.E(p_x_14_pipe_11_Z_p_O_FD));
  p_O_FD x_14_pipe_12_Z(.Q(un84_sop_0_0_0_0_0[4:4]),.D(un84_sop_0_0_0_0_1[4:4]),.C(clk),.E(p_x_14_pipe_12_Z_p_O_FD));
  p_O_FD x_14_pipe_13_Z(.Q(un84_sop_0_0_0_0_0[5:5]),.D(un84_sop_0_0_0_0_1[5:5]),.C(clk),.E(p_x_14_pipe_13_Z_p_O_FD));
  p_O_FD x_14_pipe_14_Z(.Q(un84_sop_0_0_0_0_0[6:6]),.D(un84_sop_0_0_0_0_1[6:6]),.C(clk),.E(p_x_14_pipe_14_Z_p_O_FD));
  p_O_FD x_14_pipe_15_Z(.Q(un84_sop_0_0_0_0_0[7:7]),.D(un84_sop_0_0_0_0_1[7:7]),.C(clk),.E(p_x_14_pipe_15_Z_p_O_FD));
  p_O_FD x_14_pipe_16_Z(.Q(un84_sop_0_0_0_0_0[8:8]),.D(un84_sop_0_0_0_0_1[8:8]),.C(clk),.E(p_x_14_pipe_16_Z_p_O_FD));
  p_O_FD x_14_pipe_17_Z(.Q(un84_sop_0_0_0_0_0[9:9]),.D(un84_sop_0_0_0_0_1[9:9]),.C(clk),.E(p_x_14_pipe_17_Z_p_O_FD));
  p_O_FD x_9_pipe_1_Z(.Q(un1_x_11_0_0[7:7]),.D(un1_x_11_0_0_0[7:7]),.C(clk),.E(p_x_9_pipe_1_Z_p_O_FD));
  p_O_FD x_9_pipe_2_Z(.Q(un1_x_11_0_0[8:8]),.D(un1_x_11_0_0_0[8:8]),.C(clk),.E(p_x_9_pipe_2_Z_p_O_FD));
  p_O_FD x_9_pipe_3_Z(.Q(un1_x_11_0_0[9:9]),.D(un1_x_11_0_0_0[9:9]),.C(clk),.E(p_x_9_pipe_3_Z_p_O_FD));
  p_O_FD x_9_pipe_4_Z(.Q(un1_x_11_0_0[10:10]),.D(un1_x_11_0_0_0[10:10]),.C(clk),.E(p_x_9_pipe_4_Z_p_O_FD));
  p_O_FD x_9_pipe_5_Z(.Q(un1_x_11_0_0[11:11]),.D(un1_x_11_0_0_0[11:11]),.C(clk),.E(p_x_9_pipe_5_Z_p_O_FD));
  p_O_FD x_9_pipe_6_Z(.Q(un1_x_11_0_0[12:12]),.D(un1_x_11_0_0_0[12:12]),.C(clk),.E(p_x_9_pipe_6_Z_p_O_FD));
  p_O_FD x_9_pipe_7_Z(.Q(un1_x_11_0_0[13:13]),.D(un1_x_11_0_0_0[13:13]),.C(clk),.E(p_x_9_pipe_7_Z_p_O_FD));
  p_O_FD x_9_pipe_8_Z(.Q(un1_x_11_0_0[14:14]),.D(un1_x_11_0_0_0[14:14]),.C(clk),.E(p_x_9_pipe_8_Z_p_O_FD));
  p_O_FD x_15_pipe_0_0_15_Z(.Q(un84_sop_0_0_0_10_0[0:0]),.D(un84_sop_0_0_0_0_8[0:0]),.C(clk),.E(p_x_15_pipe_0_0_15_Z_p_O_FD));
  p_O_FD x_15_pipe_0_0_16_Z(.Q(un84_sop_0_0_0_10_0[1:1]),.D(un84_sop_0_0_0_0_8[1:1]),.C(clk),.E(p_x_15_pipe_0_0_16_Z_p_O_FD));
  p_O_FD x_15_pipe_0_0_17_Z(.Q(un84_sop_0_0_0_10_0[2:2]),.D(un84_sop_0_0_0_0_8[2:2]),.C(clk),.E(p_x_15_pipe_0_0_17_Z_p_O_FD));
  p_O_FD x_15_pipe_0_0_18_Z(.Q(un84_sop_0_0_0_10_0[3:3]),.D(un84_sop_0_0_0_0_8[3:3]),.C(clk),.E(p_x_15_pipe_0_0_18_Z_p_O_FD));
  p_O_FD x_15_pipe_0_0_19_Z(.Q(un84_sop_0_0_0_10_0[4:4]),.D(un84_sop_0_0_0_0_8[4:4]),.C(clk),.E(p_x_15_pipe_0_0_19_Z_p_O_FD));
  p_O_FD x_15_pipe_0_0_20_Z(.Q(un84_sop_0_0_0_10_0[5:5]),.D(un84_sop_0_0_0_0_8[5:5]),.C(clk),.E(p_x_15_pipe_0_0_20_Z_p_O_FD));
  p_O_FD x_15_pipe_0_0_21_Z(.Q(un84_sop_0_0_0_10_0[6:6]),.D(un84_sop_0_0_0_0_8[6:6]),.C(clk),.E(p_x_15_pipe_0_0_21_Z_p_O_FD));
  p_O_FD x_15_pipe_0_0_22_Z(.Q(un84_sop_0_0_0_10_0[7:7]),.D(un84_sop_0_0_0_0_8[7:7]),.C(clk),.E(p_x_15_pipe_0_0_22_Z_p_O_FD));
  p_O_FD x_15_pipe_0_0_23_Z(.Q(un84_sop_0_0_0_10_0[8:8]),.D(un84_sop_0_0_0_0_8[8:8]),.C(clk),.E(p_x_15_pipe_0_0_23_Z_p_O_FD));
  p_O_FD x_15_pipe_0_0_24_Z(.Q(un84_sop_0_0_0_10_0[9:9]),.D(un84_sop_0_0_0_0_8[9:9]),.C(clk),.E(p_x_15_pipe_0_0_24_Z_p_O_FD));
  p_O_FD x_15_pipe_0_0_25_Z(.Q(un84_sop_0_0_0_10_0[10:10]),.D(un84_sop_0_0_0_0_8[10:10]),.C(clk),.E(p_x_15_pipe_0_0_25_Z_p_O_FD));
  p_O_FD x_15_pipe_0_0_26_Z(.Q(un84_sop_0_0_0_10_0[11:11]),.D(un84_sop_0_0_0_0_8[11:11]),.C(clk),.E(p_x_15_pipe_0_0_26_Z_p_O_FD));
  p_O_FD x_15_pipe_0_0_27_Z(.Q(un84_sop_0_0_0_10_0[12:12]),.D(un84_sop_0_0_0_0_8[12:12]),.C(clk),.E(p_x_15_pipe_0_0_27_Z_p_O_FD));
  p_O_FD x_15_pipe_0_0_28_Z(.Q(un84_sop_0_0_0_10_0[13:13]),.D(un84_sop_0_0_0_0_8[13:13]),.C(clk),.E(p_x_15_pipe_0_0_28_Z_p_O_FD));
  p_O_FD x_15_pipe_0_0_29_Z(.Q(un84_sop_0_0_0_10_0[14:14]),.D(un84_sop_0_0_0_0_8[14:14]),.C(clk),.E(p_x_15_pipe_0_0_29_Z_p_O_FD));
  p_O_FD x_16_pipe_0_0_0_Z(.Q(un84_sop_0_0_0_0_5[0:0]),.D(un84_sop_0_0_0_5_0[0:0]),.C(clk),.E(p_x_16_pipe_0_0_0_Z_p_O_FD));
  p_O_FD x_16_pipe_0_0_1_Z(.Q(un84_sop_0_0_0_0_5[1:1]),.D(un84_sop_0_0_0_5_0[1:1]),.C(clk),.E(p_x_16_pipe_0_0_1_Z_p_O_FD));
  p_O_FD x_16_pipe_0_0_2_Z(.Q(un84_sop_0_0_0_0_5[2:2]),.D(un84_sop_0_0_0_5_0[2:2]),.C(clk),.E(p_x_16_pipe_0_0_2_Z_p_O_FD));
  p_O_FD x_16_pipe_0_0_3_Z(.Q(un84_sop_0_0_0_0_5[3:3]),.D(un84_sop_0_0_0_5_0[3:3]),.C(clk),.E(p_x_16_pipe_0_0_3_Z_p_O_FD));
  p_O_FD x_16_pipe_0_0_4_Z(.Q(un84_sop_0_0_0_0_5[4:4]),.D(un84_sop_0_0_0_5_0[4:4]),.C(clk),.E(p_x_16_pipe_0_0_4_Z_p_O_FD));
  p_O_FD x_16_pipe_0_0_5_Z(.Q(un84_sop_0_0_0_0_5[5:5]),.D(un84_sop_0_0_0_5_0[5:5]),.C(clk),.E(p_x_16_pipe_0_0_5_Z_p_O_FD));
  p_O_FD x_16_pipe_0_0_6_Z(.Q(un84_sop_0_0_0_0_5[6:6]),.D(un84_sop_0_0_0_5_0[6:6]),.C(clk),.E(p_x_16_pipe_0_0_6_Z_p_O_FD));
  p_O_FD x_16_pipe_0_0_7_Z(.Q(un84_sop_0_0_0_0_5[7:7]),.D(un84_sop_0_0_0_5_0[7:7]),.C(clk),.E(p_x_16_pipe_0_0_7_Z_p_O_FD));
  p_O_FD x_16_pipe_0_0_8_Z(.Q(un84_sop_0_0_0_0_5[8:8]),.D(un84_sop_0_0_0_5_0[8:8]),.C(clk),.E(p_x_16_pipe_0_0_8_Z_p_O_FD));
  p_O_FD x_16_pipe_0_0_9_Z(.Q(un84_sop_0_0_0_0_5[9:9]),.D(un84_sop_0_0_0_5_0[9:9]),.C(clk),.E(p_x_16_pipe_0_0_9_Z_p_O_FD));
  p_O_FD x_16_pipe_0_0_10_Z(.Q(un84_sop_0_0_0_0_5[10:10]),.D(un84_sop_0_0_0_5_0[10:10]),.C(clk),.E(p_x_16_pipe_0_0_10_Z_p_O_FD));
  p_O_FD x_16_pipe_0_0_11_Z(.Q(un84_sop_0_0_0_0_5[11:11]),.D(un84_sop_0_0_0_5_0[11:11]),.C(clk),.E(p_x_16_pipe_0_0_11_Z_p_O_FD));
  p_O_FD x_16_pipe_0_0_12_Z(.Q(un84_sop_0_0_0_0_5[12:12]),.D(un84_sop_0_0_0_5_0[12:12]),.C(clk),.E(p_x_16_pipe_0_0_12_Z_p_O_FD));
  p_O_FD x_16_pipe_0_0_13_Z(.Q(un84_sop_0_0_0_0_5[13:13]),.D(un84_sop_0_0_0_5_0[13:13]),.C(clk),.E(p_x_16_pipe_0_0_13_Z_p_O_FD));
  p_O_FD x_16_pipe_0_0_14_Z(.Q(un84_sop_0_0_0_0_5[14:14]),.D(un84_sop_0_0_0_5_0[14:14]),.C(clk),.E(p_x_16_pipe_0_0_14_Z_p_O_FD));
  p_O_FD desc33(.Q(x_4[7:7]),.D(x_4_tmp_d_array_0),.C(clk),.E(p_desc33_p_O_FD));
  p_O_FD desc34(.Q(x_4[6:6]),.D(x_4_0_tmp_d_array_0),.C(clk),.E(p_desc34_p_O_FD));
  p_O_FD desc35(.Q(x_4[5:5]),.D(x_4_1_tmp_d_array_0),.C(clk),.E(p_desc35_p_O_FD));
  p_O_FD desc36(.Q(x_4[4:4]),.D(x_4_2_tmp_d_array_0),.C(clk),.E(p_desc36_p_O_FD));
  p_O_FD desc37(.Q(x_4[3:3]),.D(x_4_3_tmp_d_array_0),.C(clk),.E(p_desc37_p_O_FD));
  p_O_FD desc38(.Q(x_4[2:2]),.D(x_4_4_tmp_d_array_0),.C(clk),.E(p_desc38_p_O_FD));
  p_O_FD desc39(.Q(x_4[1:1]),.D(x_4_5_tmp_d_array_0),.C(clk),.E(p_desc39_p_O_FD));
  p_O_FD desc40(.Q(x_4[0:0]),.D(x_4_6_tmp_d_array_0),.C(clk),.E(p_desc40_p_O_FD));
  p_O_FD desc41(.Q(x_7[7:7]),.D(x_7_tmp_d_array_0),.C(clk),.E(p_desc41_p_O_FD));
  p_O_FD desc42(.Q(x_7[6:6]),.D(x_7_0_tmp_d_array_0),.C(clk),.E(p_desc42_p_O_FD));
  p_O_FD desc43(.Q(x_7[5:5]),.D(x_7_1_tmp_d_array_0),.C(clk),.E(p_desc43_p_O_FD));
  p_O_FD desc44(.Q(x_7[4:4]),.D(x_7_2_tmp_d_array_0),.C(clk),.E(p_desc44_p_O_FD));
  p_O_FD desc45(.Q(x_7[3:3]),.D(x_7_3_tmp_d_array_0),.C(clk),.E(p_desc45_p_O_FD));
  p_O_FD desc46(.Q(x_7[2:2]),.D(x_7_4_tmp_d_array_0),.C(clk),.E(p_desc46_p_O_FD));
  p_O_FD desc47(.Q(x_7[1:1]),.D(x_7_5_tmp_d_array_0),.C(clk),.E(p_desc47_p_O_FD));
  p_O_FD desc48(.Q(x_7[0:0]),.D(x_7_6_tmp_d_array_0),.C(clk),.E(p_desc48_p_O_FD));
  p_O_FD desc49(.Q(x_12[7:7]),.D(x_12_tmp_d_array_0),.C(clk),.E(p_desc49_p_O_FD));
  p_O_FD desc50(.Q(x_12[6:6]),.D(x_12_0_tmp_d_array_0),.C(clk),.E(p_desc50_p_O_FD));
  p_O_FD desc51(.Q(x_12[5:5]),.D(x_12_1_tmp_d_array_0),.C(clk),.E(p_desc51_p_O_FD));
  p_O_FD desc52(.Q(x_12[4:4]),.D(x_12_2_tmp_d_array_0),.C(clk),.E(p_desc52_p_O_FD));
  p_O_FD desc53(.Q(x_12[3:3]),.D(x_12_3_tmp_d_array_0),.C(clk),.E(p_desc53_p_O_FD));
  p_O_FD desc54(.Q(x_12[2:2]),.D(x_12_4_tmp_d_array_0),.C(clk),.E(p_desc54_p_O_FD));
  p_O_FD desc55(.Q(x_12[1:1]),.D(x_12_5_tmp_d_array_0),.C(clk),.E(p_desc55_p_O_FD));
  p_O_FD desc56(.Q(x_12[0:0]),.D(x_12_6_tmp_d_array_0),.C(clk),.E(p_desc56_p_O_FD));
  MUXCY_L un84_sop_1_6_0_cry_0_cy_cZ(.DI(GND),.CI(VCC),.S(un1_x_3_0[4:4]),.LO(un84_sop_1_6_0_cry_0_cy));
  MUXCY_L un84_sop_0_0_0_6_6_0_cry_0_cy_cZ(.DI(GND),.CI(VCC),.S(un1_x_9_0_0[5:5]),.LO(un84_sop_0_0_0_6_6_0_cry_0_cy));
  MUXCY_L un84_sop_0_0_0_11_6_0_cry_0_cy_cZ(.DI(GND),.CI(VCC),.S(un1_x_14_0_0_0[4:4]),.LO(un84_sop_0_0_0_11_6_0_cry_0_cy));
  LUT3 un84_sop_0_0_0_11_0_cry_2_RNO_cZ(.I0(x_8[1:1]),.I1(x_8[0:0]),.I2(un84_sop_0_0_0_0_11_7[1:1]),.O(un84_sop_0_0_0_11_0_cry_2_RNO));
defparam un84_sop_0_0_0_11_0_cry_2_RNO_cZ.INIT=8'h60;
  LUT6 un84_sop_0_0_0_11_6_0_axb_8_cZ(.I0(un1_x_12_0_0[11:11]),.I1(un1_x_12_0_0[12:12]),.I2(un1_x_13_0_0[12:12]),.I3(un1_x_13_0_0[13:13]),.I4(un1_x_14_0_0[11:11]),.I5(un1_x_14_0_0[12:12]),.O(un84_sop_0_0_0_11_6_0_axb_8));
defparam un84_sop_0_0_0_11_6_0_axb_8_cZ.INIT=64'h36C96C93C936936C;
  LUT6 un84_sop_0_0_0_11_6_0_axb_3_cZ(.I0(un1_x_12_0_0[6:6]),.I1(un1_x_12_0_0[7:7]),.I2(un1_x_13_0_0[7:7]),.I3(un1_x_13_0_0[8:8]),.I4(un1_x_14_0_0[6:6]),.I5(un1_x_14_0_0[7:7]),.O(un84_sop_0_0_0_11_6_0_axb_3));
defparam un84_sop_0_0_0_11_6_0_axb_3_cZ.INIT=64'h36C96C93C936936C;
  LUT6 un84_sop_0_0_0_11_6_0_axb_4_cZ(.I0(un1_x_12_0_0[7:7]),.I1(un1_x_12_0_0[8:8]),.I2(un1_x_13_0_0[8:8]),.I3(un1_x_13_0_0[9:9]),.I4(un1_x_14_0_0[7:7]),.I5(un1_x_14_0_0[8:8]),.O(un84_sop_0_0_0_11_6_0_axb_4));
defparam un84_sop_0_0_0_11_6_0_axb_4_cZ.INIT=64'h36C96C93C936936C;
  LUT6 un84_sop_0_0_0_11_6_0_axb_9_cZ(.I0(un1_x_12_0_0[12:12]),.I1(un1_x_12_0_0[13:13]),.I2(un1_x_13_0_0[13:13]),.I3(un1_x_13_0_0[14:14]),.I4(un1_x_14_0_0[12:12]),.I5(un1_x_14_0_0[13:13]),.O(un84_sop_0_0_0_11_6_0_axb_9));
defparam un84_sop_0_0_0_11_6_0_axb_9_cZ.INIT=64'h36C96C93C936936C;
  LUT5 un84_sop_0_0_0_11_6_0_axb_11_cZ(.I0(un1_x_12_0_0[14:14]),.I1(un1_x_14_0_0[14:14]),.I2(un1_x_12_0_0[15:15]),.I3(un1_x_14_0_0[15:15]),.I4(un1_x_13_0_0[15:15]),.O(un84_sop_0_0_0_11_6_0_axb_11));
defparam un84_sop_0_0_0_11_6_0_axb_11_cZ.INIT=32'h1EE18778;
  LUT6 un84_sop_1_6_0_axb_4_cZ(.I0(un1_x_1[7:7]),.I1(un1_x_1[8:8]),.I2(un1_x_2[8:8]),.I3(un1_x_2[9:9]),.I4(un1_x_3[7:7]),.I5(un1_x_3[8:8]),.O(un84_sop_1_6_0_axb_4));
defparam un84_sop_1_6_0_axb_4_cZ.INIT=64'h36C96C93C936936C;
  LUT6 un84_sop_0_0_0_11_6_0_axb_10_cZ(.I0(un1_x_12_0_0[13:13]),.I1(un1_x_12_0_0[14:14]),.I2(un1_x_13_0_0[14:14]),.I3(un1_x_14_0_0[13:13]),.I4(un1_x_14_0_0[14:14]),.I5(un1_x_13_0_0[15:15]),.O(un84_sop_0_0_0_11_6_0_axb_10));
defparam un84_sop_0_0_0_11_6_0_axb_10_cZ.INIT=64'h366CC993C993366C;
  LUT6 un84_sop_0_0_0_11_6_0_axb_2_cZ(.I0(un1_x_12_0_0[5:5]),.I1(un1_x_12_0_0[6:6]),.I2(un1_x_13_0_0[6:6]),.I3(un1_x_13_0_0[7:7]),.I4(un1_x_14_0_0[5:5]),.I5(un1_x_14_0_0[6:6]),.O(un84_sop_0_0_0_11_6_0_axb_2));
defparam un84_sop_0_0_0_11_6_0_axb_2_cZ.INIT=64'h36C96C93C936936C;
  LUT6_L un84_sop_0_0_0_11_0_axb_5_cZ(.I0(un84_sop_0_0_0_0_11_7[4:4]),.I1(un84_sop_0_0_0_0_11_7[5:5]),.I2(un84_sop_0_0_0_0_11_6[4:4]),.I3(un84_sop_0_0_0_0_11_6[5:5]),.I4(un1_x_10_0_0[8:8]),.I5(un1_x_10_0_0[9:9]),.LO(un84_sop_0_0_0_11_0_axb_5));
defparam un84_sop_0_0_0_11_0_axb_5_cZ.INIT=64'h36C96C93C936936C;
  LUT6_L un84_sop_0_0_0_11_0_axb_6_cZ(.I0(un84_sop_0_0_0_0_11_7[5:5]),.I1(un84_sop_0_0_0_0_11_7[6:6]),.I2(un84_sop_0_0_0_0_11_6[5:5]),.I3(un84_sop_0_0_0_0_11_6[6:6]),.I4(un1_x_10_0_0[9:9]),.I5(un1_x_10_0_0[10:10]),.LO(un84_sop_0_0_0_11_0_axb_6));
defparam un84_sop_0_0_0_11_0_axb_6_cZ.INIT=64'h36C96C93C936936C;
  LUT6 un84_sop_0_0_0_11_6_0_axb_6_cZ(.I0(un1_x_12_0_0[9:9]),.I1(un1_x_12_0_0[10:10]),.I2(un1_x_13_0_0[10:10]),.I3(un1_x_13_0_0[11:11]),.I4(un1_x_14_0_0[9:9]),.I5(un1_x_14_0_0[10:10]),.O(un84_sop_0_0_0_11_6_0_axb_6));
defparam un84_sop_0_0_0_11_6_0_axb_6_cZ.INIT=64'h36C96C93C936936C;
  LUT6 un84_sop_0_0_0_11_6_0_axb_7_cZ(.I0(un1_x_12_0_0[10:10]),.I1(un1_x_12_0_0[11:11]),.I2(un1_x_13_0_0[11:11]),.I3(un1_x_13_0_0[12:12]),.I4(un1_x_14_0_0[10:10]),.I5(un1_x_14_0_0[11:11]),.O(un84_sop_0_0_0_11_6_0_axb_7));
defparam un84_sop_0_0_0_11_6_0_axb_7_cZ.INIT=64'h36C96C93C936936C;
  LUT6_L un84_sop_0_0_0_11_0_axb_10_cZ(.I0(un84_sop_0_0_0_0_11_7[9:9]),.I1(un84_sop_0_0_0_0_11_7[14:14]),.I2(un84_sop_0_0_0_0_11_6[9:9]),.I3(un84_sop_0_0_0_0_11_6[10:10]),.I4(un1_x_10_0_0[13:13]),.I5(un1_x_10_0_0[14:14]),.LO(un84_sop_0_0_0_11_0_axb_10));
defparam un84_sop_0_0_0_11_0_axb_10_cZ.INIT=64'h36C96C93C936936C;
  LUT4_L un84_sop_0_0_0_11_0_axb_12_cZ(.I0(un84_sop_0_0_0_0_11_7[14:14]),.I1(un84_sop_0_0_0_0_11_6[11:11]),.I2(un84_sop_0_0_0_0_11_6[12:12]),.I3(un1_x_10_0_0[15:15]),.LO(un84_sop_0_0_0_11_0_axb_12));
defparam un84_sop_0_0_0_11_0_axb_12_cZ.INIT=16'h4BD2;
  LUT4_L un84_sop_0_0_0_11_0_axb_13_cZ(.I0(un84_sop_0_0_0_0_11_7[14:14]),.I1(un84_sop_0_0_0_0_11_6[14:14]),.I2(un84_sop_0_0_0_0_11_6[12:12]),.I3(un1_x_10_0_0[15:15]),.LO(un84_sop_0_0_0_11_0_axb_13));
defparam un84_sop_0_0_0_11_0_axb_13_cZ.INIT=16'h63C6;
  LUT3 un84_sop_0_0_0_11_6_0_axb_13_cZ(.I0(un1_x_12_0_0[15:15]),.I1(un1_x_14_0_0[15:15]),.I2(un1_x_13_0_0[15:15]),.O(un84_sop_0_0_0_11_6_0_axb_13));
defparam un84_sop_0_0_0_11_6_0_axb_13_cZ.INIT=8'h7E;
  LUT6_L un84_sop_0_0_0_11_0_axb_3_cZ(.I0(un84_sop_0_0_0_0_11_7[2:2]),.I1(un84_sop_0_0_0_0_11_7[3:3]),.I2(un84_sop_0_0_0_0_11_6[2:2]),.I3(un1_x_10_s_2_sf),.I4(un1_x_10_axb_3),.I5(un84_sop_0_0_0_0_11_6[3:3]),.LO(un84_sop_0_0_0_11_0_axb_3));
defparam un84_sop_0_0_0_11_0_axb_3_cZ.INIT=64'h366CC993C993366C;
  LUT6_L un84_sop_0_0_0_11_0_axb_4_cZ(.I0(un84_sop_0_0_0_0_11_7[3:3]),.I1(un84_sop_0_0_0_0_11_7[4:4]),.I2(un1_x_10_axb_3),.I3(un84_sop_0_0_0_0_11_6[3:3]),.I4(un84_sop_0_0_0_0_11_6[4:4]),.I5(un1_x_10_0_0[8:8]),.LO(un84_sop_0_0_0_11_0_axb_4));
defparam un84_sop_0_0_0_11_0_axb_4_cZ.INIT=64'h366CC993C993366C;
  LUT6 un84_sop_0_0_0_6_6_0_axb_5_cZ(.I0(un1_x_7_0[6:6]),.I1(un1_x_7_0[7:7]),.I2(un1_x_8_0[8:8]),.I3(un1_x_8_0[9:9]),.I4(un1_x_9_0[9:9]),.I5(un1_x_9_0[10:10]),.O(un84_sop_0_0_0_6_6_0_axb_5));
defparam un84_sop_0_0_0_6_6_0_axb_5_cZ.INIT=64'h36C96C93C936936C;
  LUT6 un84_sop_0_0_0_6_6_0_axb_6_cZ(.I0(un1_x_7_0[7:7]),.I1(un1_x_7_0[8:8]),.I2(un1_x_8_0[9:9]),.I3(un1_x_8_0[10:10]),.I4(un1_x_9_0[10:10]),.I5(un1_x_9_0[11:11]),.O(un84_sop_0_0_0_6_6_0_axb_6));
defparam un84_sop_0_0_0_6_6_0_axb_6_cZ.INIT=64'h36C96C93C936936C;
  LUT6 un84_sop_0_0_0_6_6_0_axb_10_cZ(.I0(un1_x_7_0[11:11]),.I1(un1_x_7_0[12:12]),.I2(un1_x_8_0[13:13]),.I3(un1_x_8_0[14:14]),.I4(un1_x_9_0[14:14]),.I5(un1_x_9_0[15:15]),.O(un84_sop_0_0_0_6_6_0_axb_10));
defparam un84_sop_0_0_0_6_6_0_axb_10_cZ.INIT=64'h36C96C93C936936C;
  LUT5 un84_sop_0_0_0_6_6_0_axb_11_cZ(.I0(un1_x_7_0[12:12]),.I1(un1_x_7_0[13:13]),.I2(un1_x_8_0[14:14]),.I3(un1_x_8_0[15:15]),.I4(un1_x_9_0[15:15]),.O(un84_sop_0_0_0_6_6_0_axb_11));
defparam un84_sop_0_0_0_6_6_0_axb_11_cZ.INIT=32'h36C9936C;
  LUT6 un84_sop_0_0_0_1_6_8_axb_3_cZ(.I0(un84_sop_0_0_0_10_0[5:5]),.I1(un84_sop_0_0_0_10_0[6:6]),.I2(x_4[1:1]),.I3(x_4[0:0]),.I4(x_4[2:2]),.I5(x_4[3:3]),.O(un84_sop_0_0_0_1_6_8_axb_3));
defparam un84_sop_0_0_0_1_6_8_axb_3_cZ.INIT=64'h3C6969C3C396963C;
  LUT6 un84_sop_0_0_0_1_6_8_axb_4_cZ(.I0(un84_sop_0_0_0_10_0[6:6]),.I1(un84_sop_0_0_0_10_0[7:7]),.I2(x_4[1:1]),.I3(x_4[2:2]),.I4(x_4[3:3]),.I5(x_4[4:4]),.O(un84_sop_0_0_0_1_6_8_axb_4));
defparam un84_sop_0_0_0_1_6_8_axb_4_cZ.INIT=64'h36C96C93C936936C;
  LUT6 un84_sop_0_0_0_1_6_8_axb_5_cZ(.I0(un84_sop_0_0_0_10_0[7:7]),.I1(un84_sop_0_0_0_10_0[8:8]),.I2(x_4[2:2]),.I3(x_4[3:3]),.I4(x_4[4:4]),.I5(x_4[5:5]),.O(un84_sop_0_0_0_1_6_8_axb_5));
defparam un84_sop_0_0_0_1_6_8_axb_5_cZ.INIT=64'h36C96C93C936936C;
  LUT6 un84_sop_0_0_0_1_6_8_axb_6_cZ(.I0(un84_sop_0_0_0_10_0[8:8]),.I1(un84_sop_0_0_0_10_0[9:9]),.I2(x_4[6:6]),.I3(x_4[3:3]),.I4(x_4[4:4]),.I5(x_4[5:5]),.O(un84_sop_0_0_0_1_6_8_axb_6));
defparam un84_sop_0_0_0_1_6_8_axb_6_cZ.INIT=64'h3C69C39669C3963C;
  LUT6 un84_sop_0_0_0_1_6_8_axb_7_cZ(.I0(un84_sop_0_0_0_10_0[9:9]),.I1(un84_sop_0_0_0_10_0[10:10]),.I2(x_4[6:6]),.I3(x_4[4:4]),.I4(x_4[5:5]),.I5(x_4[7:7]),.O(un84_sop_0_0_0_1_6_8_axb_7));
defparam un84_sop_0_0_0_1_6_8_axb_7_cZ.INIT=64'h366CC993C993366C;
  LUT5 un84_sop_0_0_0_1_6_8_axb_8_cZ(.I0(un84_sop_0_0_0_10_0[11:11]),.I1(un84_sop_0_0_0_10_0[10:10]),.I2(x_4[6:6]),.I3(x_4[5:5]),.I4(x_4[7:7]),.O(un84_sop_0_0_0_1_6_8_axb_8));
defparam un84_sop_0_0_0_1_6_8_axb_8_cZ.INIT=32'h5A69965A;
  LUT6 un84_sop_0_0_0_11_6_0_axb_5_cZ(.I0(un1_x_12_0_0[8:8]),.I1(un1_x_12_0_0[9:9]),.I2(un1_x_13_0_0[9:9]),.I3(un1_x_13_0_0[10:10]),.I4(un1_x_14_0_0[8:8]),.I5(un1_x_14_0_0[9:9]),.O(un84_sop_0_0_0_11_6_0_axb_5));
defparam un84_sop_0_0_0_11_6_0_axb_5_cZ.INIT=64'h36C96C93C936936C;
  LUT6 un84_sop_1_6_0_axb_2_cZ(.I0(un1_x_1[5:5]),.I1(un1_x_1[6:6]),.I2(un1_x_2[6:6]),.I3(un1_x_2[7:7]),.I4(un1_x_3[5:5]),.I5(un1_x_3[6:6]),.O(un84_sop_1_6_0_axb_2));
defparam un84_sop_1_6_0_axb_2_cZ.INIT=64'h36C96C93C936936C;
  LUT6 un84_sop_1_6_0_axb_3_cZ(.I0(un1_x_1[6:6]),.I1(un1_x_1[7:7]),.I2(un1_x_2[7:7]),.I3(un1_x_2[8:8]),.I4(un1_x_3[6:6]),.I5(un1_x_3[7:7]),.O(un84_sop_1_6_0_axb_3));
defparam un84_sop_1_6_0_axb_3_cZ.INIT=64'h36C96C93C936936C;
  LUT6 un84_sop_1_6_0_axb_5_cZ(.I0(un1_x_1[8:8]),.I1(un1_x_1[9:9]),.I2(un1_x_2[9:9]),.I3(un1_x_2[10:10]),.I4(un1_x_3[8:8]),.I5(un1_x_3[9:9]),.O(un84_sop_1_6_0_axb_5));
defparam un84_sop_1_6_0_axb_5_cZ.INIT=64'h36C96C93C936936C;
  LUT6 un84_sop_1_6_0_axb_6_cZ(.I0(un1_x_1[9:9]),.I1(un1_x_1[10:10]),.I2(un1_x_2[10:10]),.I3(un1_x_2[11:11]),.I4(un1_x_3[9:9]),.I5(un1_x_3[10:10]),.O(un84_sop_1_6_0_axb_6));
defparam un84_sop_1_6_0_axb_6_cZ.INIT=64'h36C96C93C936936C;
  LUT6 un84_sop_1_6_0_axb_7_cZ(.I0(un1_x_1[10:10]),.I1(un1_x_1[11:11]),.I2(un1_x_2[11:11]),.I3(un1_x_2[12:12]),.I4(un1_x_3[10:10]),.I5(un1_x_3[11:11]),.O(un84_sop_1_6_0_axb_7));
defparam un84_sop_1_6_0_axb_7_cZ.INIT=64'h36C96C93C936936C;
  LUT6 un84_sop_1_6_0_axb_8_cZ(.I0(un1_x_1[11:11]),.I1(un1_x_1[12:12]),.I2(un1_x_2[12:12]),.I3(un1_x_2[13:13]),.I4(un1_x_3[11:11]),.I5(un1_x_3[12:12]),.O(un84_sop_1_6_0_axb_8));
defparam un84_sop_1_6_0_axb_8_cZ.INIT=64'h36C96C93C936936C;
  LUT6 un84_sop_1_6_0_axb_9_cZ(.I0(un1_x_1[12:12]),.I1(un1_x_1[13:13]),.I2(un1_x_2[13:13]),.I3(un1_x_2[14:14]),.I4(un1_x_3[12:12]),.I5(un1_x_3[13:13]),.O(un84_sop_1_6_0_axb_9));
defparam un84_sop_1_6_0_axb_9_cZ.INIT=64'h36C96C93C936936C;
  LUT6 un84_sop_1_6_0_axb_10_cZ(.I0(un1_x_1[13:13]),.I1(un1_x_1[14:14]),.I2(un1_x_2[14:14]),.I3(un1_x_3[13:13]),.I4(un1_x_3[14:14]),.I5(un1_x_2[15:15]),.O(un84_sop_1_6_0_axb_10));
defparam un84_sop_1_6_0_axb_10_cZ.INIT=64'h366CC993C993366C;
  LUT5 un84_sop_1_6_0_axb_11_cZ(.I0(un1_x_1[14:14]),.I1(un1_x_3[14:14]),.I2(un1_x_1[15:15]),.I3(un1_x_3[15:15]),.I4(un1_x_2[15:15]),.O(un84_sop_1_6_0_axb_11));
defparam un84_sop_1_6_0_axb_11_cZ.INIT=32'h1EE18778;
  LUT3 un84_sop_1_6_0_axb_13_cZ(.I0(un1_x_1[15:15]),.I1(un1_x_3[15:15]),.I2(un1_x_2[15:15]),.O(un84_sop_1_6_0_axb_13));
defparam un84_sop_1_6_0_axb_13_cZ.INIT=8'h7E;
  LUT6_L un84_sop_0_0_0_11_0_axb_7_cZ(.I0(un84_sop_0_0_0_0_11_7[6:6]),.I1(un84_sop_0_0_0_0_11_7[7:7]),.I2(un84_sop_0_0_0_0_11_6[6:6]),.I3(un84_sop_0_0_0_0_11_6[7:7]),.I4(un1_x_10_0_0[10:10]),.I5(un1_x_10_0_0[11:11]),.LO(un84_sop_0_0_0_11_0_axb_7));
defparam un84_sop_0_0_0_11_0_axb_7_cZ.INIT=64'h36C96C93C936936C;
  LUT6_L un84_sop_0_0_0_11_0_axb_8_cZ(.I0(un84_sop_0_0_0_0_11_7[7:7]),.I1(un84_sop_0_0_0_0_11_7[8:8]),.I2(un84_sop_0_0_0_0_11_6[7:7]),.I3(un84_sop_0_0_0_0_11_6[8:8]),.I4(un1_x_10_0_0[11:11]),.I5(un1_x_10_0_0[12:12]),.LO(un84_sop_0_0_0_11_0_axb_8));
defparam un84_sop_0_0_0_11_0_axb_8_cZ.INIT=64'h36C96C93C936936C;
  LUT6_L un84_sop_0_0_0_11_0_axb_9_cZ(.I0(un84_sop_0_0_0_0_11_7[8:8]),.I1(un84_sop_0_0_0_0_11_7[9:9]),.I2(un84_sop_0_0_0_0_11_6[8:8]),.I3(un84_sop_0_0_0_0_11_6[9:9]),.I4(un1_x_10_0_0[12:12]),.I5(un1_x_10_0_0[13:13]),.LO(un84_sop_0_0_0_11_0_axb_9));
defparam un84_sop_0_0_0_11_0_axb_9_cZ.INIT=64'h36C96C93C936936C;
  LUT4_L un84_sop_0_0_0_11_0_axb_1_cZ(.I0(x_8[1:1]),.I1(x_8[0:0]),.I2(un84_sop_0_0_0_0_11_7[1:1]),.I3(un84_sop_0_0_0_0_11_6[1:1]),.LO(un84_sop_0_0_0_11_0_axb_1));
defparam un84_sop_0_0_0_11_0_axb_1_cZ.INIT=16'h6996;
  LUT5_L un84_sop_0_0_0_11_0_axb_11_cZ(.I0(un84_sop_0_0_0_0_11_7[14:14]),.I1(un84_sop_0_0_0_0_11_6[10:10]),.I2(un84_sop_0_0_0_0_11_6[11:11]),.I3(un1_x_10_0_0[14:14]),.I4(un1_x_10_0_0[15:15]),.LO(un84_sop_0_0_0_11_0_axb_11));
defparam un84_sop_0_0_0_11_0_axb_11_cZ.INIT=32'h4B2DB4D2;
  LUT3 un84_sop_0_0_0_1_6_axb_0(.I0(un84_sop_0_0_0_10_0[0:0]),.I1(un1_x_6_0[1:1]),.I2(un84_sop_0_0_0_1_6_6[0:0]),.O(un84_sop_0_0_0_5_0[0:0]));
defparam un84_sop_0_0_0_1_6_axb_0.INIT=8'h96;
  LUT6 un84_sop_1_4_axb_4_cZ(.I0(x_0[3:3]),.I1(x_0[2:2]),.I2(x_0[1:1]),.I3(x_0[0:0]),.I4(x_0[4:4]),.I5(un84_sop_1_7[4:4]),.O(un84_sop_1_4_axb_4));
defparam un84_sop_1_4_axb_4_cZ.INIT=64'hFFFE00010001FFFE;
  LUT6 un84_sop_0_0_0_6_6_0_axb_2_cZ(.I0(un1_x_7_0[3:3]),.I1(un1_x_7_0[4:4]),.I2(un1_x_8_0[5:5]),.I3(un1_x_8_0[6:6]),.I4(un1_x_9_0[6:6]),.I5(un1_x_9_0[7:7]),.O(un84_sop_0_0_0_6_6_0_axb_2));
defparam un84_sop_0_0_0_6_6_0_axb_2_cZ.INIT=64'h36C96C93C936936C;
  LUT6 un84_sop_0_0_0_6_6_0_axb_3_cZ(.I0(un1_x_7_0[4:4]),.I1(un1_x_7_0[5:5]),.I2(un1_x_8_0[6:6]),.I3(un1_x_8_0[7:7]),.I4(un1_x_9_0[7:7]),.I5(un1_x_9_0[8:8]),.O(un84_sop_0_0_0_6_6_0_axb_3));
defparam un84_sop_0_0_0_6_6_0_axb_3_cZ.INIT=64'h36C96C93C936936C;
  LUT6 un84_sop_0_0_0_6_6_0_axb_4_cZ(.I0(un1_x_7_0[5:5]),.I1(un1_x_7_0[6:6]),.I2(un1_x_8_0[7:7]),.I3(un1_x_8_0[8:8]),.I4(un1_x_9_0[8:8]),.I5(un1_x_9_0[9:9]),.O(un84_sop_0_0_0_6_6_0_axb_4));
defparam un84_sop_0_0_0_6_6_0_axb_4_cZ.INIT=64'h36C96C93C936936C;
  LUT6_L un84_sop_0_0_0_11_6_0_s_2_RNIGK751(.I0(x_8[1:1]),.I1(x_8[0:0]),.I2(un84_sop_0_0_0_0_11_7[1:1]),.I3(un84_sop_0_0_0_0_11_7[2:2]),.I4(un84_sop_0_0_0_0_11_6[2:2]),.I5(un1_x_10_s_2_sf),.LO(un84_sop_0_0_0_11_0_axb_2));
defparam un84_sop_0_0_0_11_6_0_s_2_RNIGK751.INIT=64'h9F60609F609F9F60;
  LUT6 un84_sop_0_0_0_6_6_0_axb_7_cZ(.I0(un1_x_7_0[8:8]),.I1(un1_x_7_0[9:9]),.I2(un1_x_8_0[10:10]),.I3(un1_x_8_0[11:11]),.I4(un1_x_9_0[11:11]),.I5(un1_x_9_0[12:12]),.O(un84_sop_0_0_0_6_6_0_axb_7));
defparam un84_sop_0_0_0_6_6_0_axb_7_cZ.INIT=64'h36C96C93C936936C;
  LUT6 un84_sop_0_0_0_6_6_0_axb_8_cZ(.I0(un1_x_7_0[9:9]),.I1(un1_x_7_0[10:10]),.I2(un1_x_8_0[11:11]),.I3(un1_x_8_0[12:12]),.I4(un1_x_9_0[12:12]),.I5(un1_x_9_0[13:13]),.O(un84_sop_0_0_0_6_6_0_axb_8));
defparam un84_sop_0_0_0_6_6_0_axb_8_cZ.INIT=64'h36C96C93C936936C;
  LUT6 un84_sop_0_0_0_6_6_0_axb_9_cZ(.I0(un1_x_7_0[10:10]),.I1(un1_x_7_0[11:11]),.I2(un1_x_8_0[12:12]),.I3(un1_x_8_0[13:13]),.I4(un1_x_9_0[13:13]),.I5(un1_x_9_0[14:14]),.O(un84_sop_0_0_0_6_6_0_axb_9));
defparam un84_sop_0_0_0_6_6_0_axb_9_cZ.INIT=64'h36C96C93C936936C;
  LUT4 un1_x_10_axb_11_cZ(.I0(x_8[6:6]),.I1(x_8[7:7]),.I2(x_8[5:5]),.I3(un1_x_10_5_c5),.O(un1_x_10_axb_11));
defparam un1_x_10_axb_11_cZ.INIT=16'hFEFF;
  LUT3_L un84_sop_0_0_0_11_0_axb_14_cZ(.I0(un84_sop_0_0_0_0_11_7[14:14]),.I1(un84_sop_0_0_0_0_11_6[14:14]),.I2(un1_x_10_0_0[15:15]),.LO(un84_sop_0_0_0_11_0_axb_14));
defparam un84_sop_0_0_0_11_0_axb_14_cZ.INIT=8'h7E;
  LUT3 un84_sop_0_0_0_6_6_0_axb_14_cZ(.I0(un1_x_7_0[15:15]),.I1(un1_x_8_0[15:15]),.I2(un1_x_9_0[15:15]),.O(un84_sop_0_0_0_6_6_0_axb_14));
defparam un84_sop_0_0_0_6_6_0_axb_14_cZ.INIT=8'h7E;
  MUXCY_L un84_sop_0_0_0_11_0_cry_0_cy_cZ(.DI(GND),.CI(VCC),.S(un84_sop_0_0_0_0_11_7_axb_0_ci),.LO(un84_sop_0_0_0_11_0_cry_0_cy));
  LUT1 un1_x_10_4_s_2_RNI13H1(.I0(un1_x_10_4[2:2]),.O(un1_x_10_s_2_sf));
defparam un1_x_10_4_s_2_RNI13H1.INIT=2'h2;
  LUT2_L un84_sop_0_0_0_1_axb_9_cZ(.I0(un1_x_16_0_0_0[14:14]),.I1(un1_x_15_0_0_0[14:14]),.LO(un84_sop_0_0_0_1_axb_9));
defparam un84_sop_0_0_0_1_axb_9_cZ.INIT=4'h6;
  LUT2_L un84_sop_0_0_0_1_axb_8_cZ(.I0(un1_x_16_0_0_0[14:14]),.I1(un1_x_15_0_0_0[14:14]),.LO(un84_sop_0_0_0_1_axb_8));
defparam un84_sop_0_0_0_1_axb_8_cZ.INIT=4'h6;
  LUT2_L un84_sop_0_0_0_1_axb_7_cZ(.I0(un1_x_16_0_0_0[13:13]),.I1(un1_x_15_0_0_0[13:13]),.LO(un84_sop_0_0_0_1_axb_7));
defparam un84_sop_0_0_0_1_axb_7_cZ.INIT=4'h6;
  LUT2_L un84_sop_0_0_0_1_axb_6_cZ(.I0(un1_x_16_0_0_0[12:12]),.I1(un1_x_15_0_0_0[12:12]),.LO(un84_sop_0_0_0_1_axb_6));
defparam un84_sop_0_0_0_1_axb_6_cZ.INIT=4'h6;
  LUT2_L un84_sop_0_0_0_1_axb_5_cZ(.I0(un1_x_16_0_0_0[11:11]),.I1(un1_x_15_0_0_0[11:11]),.LO(un84_sop_0_0_0_1_axb_5));
defparam un84_sop_0_0_0_1_axb_5_cZ.INIT=4'h6;
  LUT2_L un84_sop_0_0_0_1_axb_4_cZ(.I0(un1_x_16_0_0_0[10:10]),.I1(un1_x_15_0_0_0[10:10]),.LO(un84_sop_0_0_0_1_axb_4));
defparam un84_sop_0_0_0_1_axb_4_cZ.INIT=4'h6;
  LUT2_L un84_sop_0_0_0_1_axb_3_cZ(.I0(un1_x_16_0_0_0[9:9]),.I1(un1_x_15_0_0_0[9:9]),.LO(un84_sop_0_0_0_1_axb_3));
defparam un84_sop_0_0_0_1_axb_3_cZ.INIT=4'h6;
  LUT2_L un84_sop_0_0_0_1_axb_2_cZ(.I0(un1_x_16_0_0_0[8:8]),.I1(un1_x_15_0_0_0[8:8]),.LO(un84_sop_0_0_0_1_axb_2));
defparam un84_sop_0_0_0_1_axb_2_cZ.INIT=4'h6;
  LUT2_L un84_sop_0_0_0_1_axb_1_cZ(.I0(un1_x_16_0_0_0[7:7]),.I1(un1_x_15_0_0_0[7:7]),.LO(un84_sop_0_0_0_1_axb_1));
defparam un84_sop_0_0_0_1_axb_1_cZ.INIT=4'h6;
  LUT2 un84_sop_0_0_0_1_axb_0(.I0(x_12[0:0]),.I1(x_13[0:0]),.O(un84_sop_0_0_0_0_1[0:0]));
defparam un84_sop_0_0_0_1_axb_0.INIT=4'h6;
  LUT1 un1_x_16_0_axb_8_cZ(.I0(x_13[7:7]),.O(un1_x_16_0_axb_8));
defparam un1_x_16_0_axb_8_cZ.INIT=2'h1;
  LUT1_L un1_x_11_0_axb_8_cZ(.I0(x_8[7:7]),.LO(un1_x_11_0_axb_8));
defparam un1_x_11_0_axb_8_cZ.INIT=2'h1;
  LUT1_L un1_x_11_0_axb_7_cZ(.I0(x_8[7:7]),.LO(un1_x_11_0_axb_7));
defparam un1_x_11_0_axb_7_cZ.INIT=2'h1;
  LUT1_L un1_x_11_0_axb_6_cZ(.I0(x_8[6:6]),.LO(un1_x_11_0_axb_6));
defparam un1_x_11_0_axb_6_cZ.INIT=2'h1;
  LUT1_L un1_x_11_0_axb_5_cZ(.I0(x_8[5:5]),.LO(un1_x_11_0_axb_5));
defparam un1_x_11_0_axb_5_cZ.INIT=2'h1;
  LUT1_L un1_x_11_0_axb_4_cZ(.I0(x_8[4:4]),.LO(un1_x_11_0_axb_4));
defparam un1_x_11_0_axb_4_cZ.INIT=2'h1;
  LUT1_L un1_x_11_0_axb_3_cZ(.I0(x_8[3:3]),.LO(un1_x_11_0_axb_3));
defparam un1_x_11_0_axb_3_cZ.INIT=2'h1;
  LUT1_L un1_x_11_0_axb_2_cZ(.I0(x_8[2:2]),.LO(un1_x_11_0_axb_2));
defparam un1_x_11_0_axb_2_cZ.INIT=2'h1;
  LUT1_L un1_x_11_0_axb_1_cZ(.I0(x_8[1:1]),.LO(un1_x_11_0_axb_1));
defparam un1_x_11_0_axb_1_cZ.INIT=2'h1;
  LUT1 un1_x_15_0_axb_8_cZ(.I0(x_12[7:7]),.O(un1_x_15_0_axb_8));
defparam un1_x_15_0_axb_8_cZ.INIT=2'h1;
  LUT1 un1_x_10_4_axb_10(.I0(x_8[7:7]),.O(un1_x_10_4[10:10]));
defparam un1_x_10_4_axb_10.INIT=2'h2;
  LUT1 un1_x_10_4_axb_9(.I0(x_8[7:7]),.O(un1_x_10_4[9:9]));
defparam un1_x_10_4_axb_9.INIT=2'h2;
  LUT2_L un84_sop_1_axb_14_cZ(.I0(un84_sop_1_6[14:14]),.I1(un84_sop_1_4[14:14]),.LO(un84_sop_1_axb_14));
defparam un84_sop_1_axb_14_cZ.INIT=4'h6;
  LUT2_L un84_sop_1_axb_13_cZ(.I0(un84_sop_1_6[14:14]),.I1(un84_sop_1_4[13:13]),.LO(un84_sop_1_axb_13));
defparam un84_sop_1_axb_13_cZ.INIT=4'h6;
  LUT2_L un84_sop_1_axb_12_cZ(.I0(un84_sop_1_6[12:12]),.I1(un84_sop_1_4[12:12]),.LO(un84_sop_1_axb_12));
defparam un84_sop_1_axb_12_cZ.INIT=4'h6;
  LUT2_L un84_sop_1_axb_11_cZ(.I0(un84_sop_1_6[11:11]),.I1(un84_sop_1_4[11:11]),.LO(un84_sop_1_axb_11));
defparam un84_sop_1_axb_11_cZ.INIT=4'h6;
  LUT2_L un84_sop_1_axb_10_cZ(.I0(un84_sop_1_6[10:10]),.I1(un84_sop_1_4[10:10]),.LO(un84_sop_1_axb_10));
defparam un84_sop_1_axb_10_cZ.INIT=4'h6;
  LUT2_L un84_sop_1_axb_9_cZ(.I0(un84_sop_1_6[9:9]),.I1(un84_sop_1_4[9:9]),.LO(un84_sop_1_axb_9));
defparam un84_sop_1_axb_9_cZ.INIT=4'h6;
  LUT2_L un84_sop_1_axb_8_cZ(.I0(un84_sop_1_6[8:8]),.I1(un84_sop_1_4[8:8]),.LO(un84_sop_1_axb_8));
defparam un84_sop_1_axb_8_cZ.INIT=4'h6;
  LUT2_L un84_sop_1_axb_7_cZ(.I0(un84_sop_1_6[7:7]),.I1(un84_sop_1_4[7:7]),.LO(un84_sop_1_axb_7));
defparam un84_sop_1_axb_7_cZ.INIT=4'h6;
  LUT2 un84_sop_0_0_0_0_11_7_axb_10_cZ(.I0(un1_x_11_0_0[14:14]),.I1(un84_sop_0_0_0_0_0[9:9]),.O(un84_sop_0_0_0_0_11_7_axb_10));
defparam un84_sop_0_0_0_0_11_7_axb_10_cZ.INIT=4'h6;
  LUT2 un84_sop_1_7_axb_14_cZ(.I0(un84_sop_0_0_0_0_5[14:14]),.I1(un1_x_4[15:15]),.O(un84_sop_1_7_axb_14));
defparam un84_sop_1_7_axb_14_cZ.INIT=4'h6;
  LUT2_L un84_sop_0_0_0_1_6_axb_14_cZ(.I0(un84_sop_0_0_0_1_6_6[14:14]),.I1(un84_sop_0_0_0_1_6_4[14:14]),.LO(un84_sop_0_0_0_1_6_axb_14));
defparam un84_sop_0_0_0_1_6_axb_14_cZ.INIT=4'h6;
  LUT2_L un84_sop_0_0_0_1_6_axb_13_cZ(.I0(un84_sop_0_0_0_1_6_6[13:13]),.I1(un84_sop_0_0_0_1_6_4[13:13]),.LO(un84_sop_0_0_0_1_6_axb_13));
defparam un84_sop_0_0_0_1_6_axb_13_cZ.INIT=4'h6;
  LUT2_L un84_sop_0_0_0_1_6_axb_12_cZ(.I0(un84_sop_0_0_0_1_6_6[12:12]),.I1(un84_sop_0_0_0_1_6_4[12:12]),.LO(un84_sop_0_0_0_1_6_axb_12));
defparam un84_sop_0_0_0_1_6_axb_12_cZ.INIT=4'h6;
  LUT2_L un84_sop_0_0_0_1_6_axb_11_cZ(.I0(un84_sop_0_0_0_1_6_6[11:11]),.I1(un84_sop_0_0_0_1_6_4[11:11]),.LO(un84_sop_0_0_0_1_6_axb_11));
defparam un84_sop_0_0_0_1_6_axb_11_cZ.INIT=4'h6;
  LUT2_L un84_sop_0_0_0_1_6_axb_10_cZ(.I0(un84_sop_0_0_0_1_6_6[10:10]),.I1(un84_sop_0_0_0_1_6_4[10:10]),.LO(un84_sop_0_0_0_1_6_axb_10));
defparam un84_sop_0_0_0_1_6_axb_10_cZ.INIT=4'h6;
  LUT2_L un84_sop_0_0_0_1_6_axb_9_cZ(.I0(un84_sop_0_0_0_1_6_6[9:9]),.I1(un84_sop_0_0_0_1_6_4[9:9]),.LO(un84_sop_0_0_0_1_6_axb_9));
defparam un84_sop_0_0_0_1_6_axb_9_cZ.INIT=4'h6;
  LUT2_L un84_sop_0_0_0_1_6_axb_8_cZ(.I0(un84_sop_0_0_0_1_6_6[8:8]),.I1(un84_sop_0_0_0_1_6_4[8:8]),.LO(un84_sop_0_0_0_1_6_axb_8));
defparam un84_sop_0_0_0_1_6_axb_8_cZ.INIT=4'h6;
  LUT2_L un84_sop_0_0_0_1_6_axb_7_cZ(.I0(un84_sop_0_0_0_1_6_6[7:7]),.I1(un84_sop_0_0_0_1_6_4[7:7]),.LO(un84_sop_0_0_0_1_6_axb_7));
defparam un84_sop_0_0_0_1_6_axb_7_cZ.INIT=4'h6;
  LUT2_L un84_sop_0_0_0_1_6_axb_6_cZ(.I0(un84_sop_0_0_0_1_6_6[6:6]),.I1(un84_sop_0_0_0_1_6_4[6:6]),.LO(un84_sop_0_0_0_1_6_axb_6));
defparam un84_sop_0_0_0_1_6_axb_6_cZ.INIT=4'h6;
  LUT2_L un84_sop_0_0_0_1_6_axb_5_cZ(.I0(un84_sop_0_0_0_1_6_6[5:5]),.I1(un84_sop_0_0_0_1_6_4[5:5]),.LO(un84_sop_0_0_0_1_6_axb_5));
defparam un84_sop_0_0_0_1_6_axb_5_cZ.INIT=4'h6;
  LUT2_L un84_sop_0_0_0_1_6_axb_4_cZ(.I0(un84_sop_0_0_0_1_6_6[4:4]),.I1(un84_sop_0_0_0_1_6_4[4:4]),.LO(un84_sop_0_0_0_1_6_axb_4));
defparam un84_sop_0_0_0_1_6_axb_4_cZ.INIT=4'h6;
  LUT2_L un84_sop_0_0_0_1_6_axb_3_cZ(.I0(un84_sop_0_0_0_1_6_4[3:3]),.I1(un84_sop_0_0_0_1_6_6[3:3]),.LO(un84_sop_0_0_0_1_6_axb_3));
defparam un84_sop_0_0_0_1_6_axb_3_cZ.INIT=4'h6;
  LUT2_L un84_sop_0_0_0_1_6_axb_2_cZ(.I0(un84_sop_0_0_0_1_6_4[2:2]),.I1(un84_sop_0_0_0_1_6_6[2:2]),.LO(un84_sop_0_0_0_1_6_axb_2));
defparam un84_sop_0_0_0_1_6_axb_2_cZ.INIT=4'h6;
  LUT2_L un84_sop_0_0_0_1_6_axb_1_cZ(.I0(un84_sop_0_0_0_1_6_4[1:1]),.I1(un84_sop_0_0_0_1_6_6[1:1]),.LO(un84_sop_0_0_0_1_6_axb_1));
defparam un84_sop_0_0_0_1_6_axb_1_cZ.INIT=4'h6;
  LUT2 un84_sop_0_0_0_1_6_4_axb_14_cZ(.I0(un1_x_6_0[15:15]),.I1(un84_sop_0_0_0_1_6_8[14:14]),.O(un84_sop_0_0_0_1_6_4_axb_14));
defparam un84_sop_0_0_0_1_6_4_axb_14_cZ.INIT=4'h6;
  LUT2 un1_x_10_axb_3_cZ(.I0(x_8[0:0]),.I1(un1_x_10_4[3:3]),.O(un1_x_10_axb_3));
defparam un1_x_10_axb_3_cZ.INIT=4'h6;
  LUT2 un84_sop_0_0_0_1_6_8_axb_11_cZ(.I0(un84_sop_0_0_0_10_0[14:14]),.I1(x_4[7:7]),.O(un84_sop_0_0_0_1_6_8_axb_11));
defparam un84_sop_0_0_0_1_6_8_axb_11_cZ.INIT=4'h6;
  LUT2_L un84_sop_0_0_0_11_0_axb_0_cZ(.I0(x_8[0:0]),.I1(un84_sop_0_0_0_0_11_6[0:0]),.LO(un84_sop_0_0_0_11_0_axb_0));
defparam un84_sop_0_0_0_11_0_axb_0_cZ.INIT=4'h6;
  LUT4 un1_x_0_0_ac0_5(.I0(x_0[3:3]),.I1(x_0[2:2]),.I2(x_0[1:1]),.I3(x_0[0:0]),.O(un1_x_0_0_c4));
defparam un1_x_0_0_ac0_5.INIT=16'h0001;
  LUT3 un84_sop_0_0_0_11_6_0_o5_11_cZ(.I0(un1_x_12_0_0[15:15]),.I1(un1_x_14_0_0[15:15]),.I2(un1_x_13_0_0[15:15]),.O(un84_sop_0_0_0_11_6_0_o5_11));
defparam un84_sop_0_0_0_11_6_0_o5_11_cZ.INIT=8'hE8;
  LUT3 un84_sop_0_0_0_11_6_0_o5_10_cZ(.I0(un1_x_12_0_0[14:14]),.I1(un1_x_14_0_0[14:14]),.I2(un1_x_13_0_0[15:15]),.O(un84_sop_0_0_0_11_6_0_o5_10));
defparam un84_sop_0_0_0_11_6_0_o5_10_cZ.INIT=8'hE8;
  LUT3 un84_sop_0_0_0_11_6_0_o5_9_cZ(.I0(un1_x_12_0_0[13:13]),.I1(un1_x_13_0_0[14:14]),.I2(un1_x_14_0_0[13:13]),.O(un84_sop_0_0_0_11_6_0_o5_9));
defparam un84_sop_0_0_0_11_6_0_o5_9_cZ.INIT=8'hE8;
  LUT3 un84_sop_0_0_0_11_6_0_o5_8_cZ(.I0(un1_x_12_0_0[12:12]),.I1(un1_x_13_0_0[13:13]),.I2(un1_x_14_0_0[12:12]),.O(un84_sop_0_0_0_11_6_0_o5_8));
defparam un84_sop_0_0_0_11_6_0_o5_8_cZ.INIT=8'hE8;
  LUT3 un84_sop_0_0_0_11_6_0_o5_7_cZ(.I0(un1_x_12_0_0[11:11]),.I1(un1_x_13_0_0[12:12]),.I2(un1_x_14_0_0[11:11]),.O(un84_sop_0_0_0_11_6_0_o5_7));
defparam un84_sop_0_0_0_11_6_0_o5_7_cZ.INIT=8'hE8;
  LUT3 un84_sop_0_0_0_11_6_0_o5_6_cZ(.I0(un1_x_12_0_0[10:10]),.I1(un1_x_13_0_0[11:11]),.I2(un1_x_14_0_0[10:10]),.O(un84_sop_0_0_0_11_6_0_o5_6));
defparam un84_sop_0_0_0_11_6_0_o5_6_cZ.INIT=8'hE8;
  LUT3 un84_sop_0_0_0_11_6_0_o5_5_cZ(.I0(un1_x_12_0_0[9:9]),.I1(un1_x_13_0_0[10:10]),.I2(un1_x_14_0_0[9:9]),.O(un84_sop_0_0_0_11_6_0_o5_5));
defparam un84_sop_0_0_0_11_6_0_o5_5_cZ.INIT=8'hE8;
  LUT3 un84_sop_0_0_0_11_6_0_o5_4_cZ(.I0(un1_x_12_0_0[8:8]),.I1(un1_x_13_0_0[9:9]),.I2(un1_x_14_0_0[8:8]),.O(un84_sop_0_0_0_11_6_0_o5_4));
defparam un84_sop_0_0_0_11_6_0_o5_4_cZ.INIT=8'hE8;
  LUT3 un84_sop_0_0_0_11_6_0_o5_3_cZ(.I0(un1_x_12_0_0[7:7]),.I1(un1_x_13_0_0[8:8]),.I2(un1_x_14_0_0[7:7]),.O(un84_sop_0_0_0_11_6_0_o5_3));
defparam un84_sop_0_0_0_11_6_0_o5_3_cZ.INIT=8'hE8;
  LUT3 un84_sop_0_0_0_11_6_0_o5_2_cZ(.I0(un1_x_12_0_0[6:6]),.I1(un1_x_13_0_0[7:7]),.I2(un1_x_14_0_0[6:6]),.O(un84_sop_0_0_0_11_6_0_o5_2));
defparam un84_sop_0_0_0_11_6_0_o5_2_cZ.INIT=8'hE8;
  LUT3 un84_sop_0_0_0_11_0_o5_12_cZ(.I0(un84_sop_0_0_0_0_11_7[14:14]),.I1(un84_sop_0_0_0_0_11_6[12:12]),.I2(un1_x_10_0_0[15:15]),.O(un84_sop_0_0_0_11_0_o5_12));
defparam un84_sop_0_0_0_11_0_o5_12_cZ.INIT=8'hE8;
  LUT3 un84_sop_0_0_0_11_0_o5_11_cZ(.I0(un84_sop_0_0_0_0_11_7[14:14]),.I1(un84_sop_0_0_0_0_11_6[11:11]),.I2(un1_x_10_0_0[15:15]),.O(un84_sop_0_0_0_11_0_o5_11));
defparam un84_sop_0_0_0_11_0_o5_11_cZ.INIT=8'hE8;
  LUT3 un84_sop_0_0_0_11_0_o5_10_cZ(.I0(un84_sop_0_0_0_0_11_7[14:14]),.I1(un84_sop_0_0_0_0_11_6[10:10]),.I2(un1_x_10_0_0[14:14]),.O(un84_sop_0_0_0_11_0_o5_10));
defparam un84_sop_0_0_0_11_0_o5_10_cZ.INIT=8'hE8;
  LUT3 un84_sop_0_0_0_11_0_o5_9_cZ(.I0(un84_sop_0_0_0_0_11_7[9:9]),.I1(un84_sop_0_0_0_0_11_6[9:9]),.I2(un1_x_10_0_0[13:13]),.O(un84_sop_0_0_0_11_0_o5_9));
defparam un84_sop_0_0_0_11_0_o5_9_cZ.INIT=8'hE8;
  LUT3 un84_sop_0_0_0_11_0_o5_8_cZ(.I0(un84_sop_0_0_0_0_11_7[8:8]),.I1(un84_sop_0_0_0_0_11_6[8:8]),.I2(un1_x_10_0_0[12:12]),.O(un84_sop_0_0_0_11_0_o5_8));
defparam un84_sop_0_0_0_11_0_o5_8_cZ.INIT=8'hE8;
  LUT3 un84_sop_0_0_0_11_0_o5_7_cZ(.I0(un84_sop_0_0_0_0_11_7[7:7]),.I1(un84_sop_0_0_0_0_11_6[7:7]),.I2(un1_x_10_0_0[11:11]),.O(un84_sop_0_0_0_11_0_o5_7));
defparam un84_sop_0_0_0_11_0_o5_7_cZ.INIT=8'hE8;
  LUT3 un84_sop_0_0_0_11_0_o5_6_cZ(.I0(un84_sop_0_0_0_0_11_7[6:6]),.I1(un84_sop_0_0_0_0_11_6[6:6]),.I2(un1_x_10_0_0[10:10]),.O(un84_sop_0_0_0_11_0_o5_6));
defparam un84_sop_0_0_0_11_0_o5_6_cZ.INIT=8'hE8;
  LUT3 un84_sop_0_0_0_11_0_o5_5_cZ(.I0(un84_sop_0_0_0_0_11_7[5:5]),.I1(un84_sop_0_0_0_0_11_6[5:5]),.I2(un1_x_10_0_0[9:9]),.O(un84_sop_0_0_0_11_0_o5_5));
defparam un84_sop_0_0_0_11_0_o5_5_cZ.INIT=8'hE8;
  LUT3 un84_sop_0_0_0_11_0_o5_4_cZ(.I0(un84_sop_0_0_0_0_11_7[4:4]),.I1(un84_sop_0_0_0_0_11_6[4:4]),.I2(un1_x_10_0_0[8:8]),.O(un84_sop_0_0_0_11_0_o5_4));
defparam un84_sop_0_0_0_11_0_o5_4_cZ.INIT=8'hE8;
  LUT3 un84_sop_0_0_0_11_0_o5_3_cZ(.I0(un84_sop_0_0_0_0_11_7[3:3]),.I1(un1_x_10_axb_3),.I2(un84_sop_0_0_0_0_11_6[3:3]),.O(un84_sop_0_0_0_11_0_o5_3));
defparam un84_sop_0_0_0_11_0_o5_3_cZ.INIT=8'hE8;
  LUT3 un84_sop_0_0_0_11_0_o5_2_cZ(.I0(un84_sop_0_0_0_0_11_7[2:2]),.I1(un84_sop_0_0_0_0_11_6[2:2]),.I2(un1_x_10_s_2_sf),.O(un84_sop_0_0_0_11_0_o5_2));
defparam un84_sop_0_0_0_11_0_o5_2_cZ.INIT=8'hE8;
  LUT3 un84_sop_0_0_0_6_6_0_o5_12_cZ(.I0(un1_x_7_0[14:14]),.I1(un1_x_8_0[15:15]),.I2(un1_x_9_0[15:15]),.O(un84_sop_0_0_0_6_6_0_o5_12));
defparam un84_sop_0_0_0_6_6_0_o5_12_cZ.INIT=8'hE8;
  LUT3 un84_sop_0_0_0_6_6_0_o5_11_cZ(.I0(un1_x_7_0[13:13]),.I1(un1_x_8_0[15:15]),.I2(un1_x_9_0[15:15]),.O(un84_sop_0_0_0_6_6_0_o5_11));
defparam un84_sop_0_0_0_6_6_0_o5_11_cZ.INIT=8'hE8;
  LUT3 un84_sop_0_0_0_6_6_0_o5_10_cZ(.I0(un1_x_7_0[12:12]),.I1(un1_x_8_0[14:14]),.I2(un1_x_9_0[15:15]),.O(un84_sop_0_0_0_6_6_0_o5_10));
defparam un84_sop_0_0_0_6_6_0_o5_10_cZ.INIT=8'hE8;
  LUT3 un84_sop_0_0_0_6_6_0_o5_9_cZ(.I0(un1_x_7_0[11:11]),.I1(un1_x_8_0[13:13]),.I2(un1_x_9_0[14:14]),.O(un84_sop_0_0_0_6_6_0_o5_9));
defparam un84_sop_0_0_0_6_6_0_o5_9_cZ.INIT=8'hE8;
  LUT3 un84_sop_0_0_0_6_6_0_o5_8_cZ(.I0(un1_x_7_0[10:10]),.I1(un1_x_8_0[12:12]),.I2(un1_x_9_0[13:13]),.O(un84_sop_0_0_0_6_6_0_o5_8));
defparam un84_sop_0_0_0_6_6_0_o5_8_cZ.INIT=8'hE8;
  LUT3 un84_sop_0_0_0_6_6_0_o5_7_cZ(.I0(un1_x_7_0[9:9]),.I1(un1_x_8_0[11:11]),.I2(un1_x_9_0[12:12]),.O(un84_sop_0_0_0_6_6_0_o5_7));
defparam un84_sop_0_0_0_6_6_0_o5_7_cZ.INIT=8'hE8;
  LUT3 un84_sop_0_0_0_6_6_0_o5_6_cZ(.I0(un1_x_7_0[8:8]),.I1(un1_x_8_0[10:10]),.I2(un1_x_9_0[11:11]),.O(un84_sop_0_0_0_6_6_0_o5_6));
defparam un84_sop_0_0_0_6_6_0_o5_6_cZ.INIT=8'hE8;
  LUT3 un84_sop_0_0_0_6_6_0_o5_5_cZ(.I0(un1_x_7_0[7:7]),.I1(un1_x_8_0[9:9]),.I2(un1_x_9_0[10:10]),.O(un84_sop_0_0_0_6_6_0_o5_5));
defparam un84_sop_0_0_0_6_6_0_o5_5_cZ.INIT=8'hE8;
  LUT3 un84_sop_0_0_0_6_6_0_o5_4_cZ(.I0(un1_x_7_0[6:6]),.I1(un1_x_8_0[8:8]),.I2(un1_x_9_0[9:9]),.O(un84_sop_0_0_0_6_6_0_o5_4));
defparam un84_sop_0_0_0_6_6_0_o5_4_cZ.INIT=8'hE8;
  LUT3 un84_sop_0_0_0_6_6_0_o5_3_cZ(.I0(un1_x_7_0[5:5]),.I1(un1_x_8_0[7:7]),.I2(un1_x_9_0[8:8]),.O(un84_sop_0_0_0_6_6_0_o5_3));
defparam un84_sop_0_0_0_6_6_0_o5_3_cZ.INIT=8'hE8;
  LUT3 un84_sop_0_0_0_6_6_0_o5_2_cZ(.I0(un1_x_7_0[4:4]),.I1(un1_x_8_0[6:6]),.I2(un1_x_9_0[7:7]),.O(un84_sop_0_0_0_6_6_0_o5_2));
defparam un84_sop_0_0_0_6_6_0_o5_2_cZ.INIT=8'hE8;
  LUT3 un84_sop_0_0_0_1_6_8_o5_7_cZ(.I0(un84_sop_0_0_0_10_0[10:10]),.I1(x_4[5:5]),.I2(x_4[7:7]),.O(un84_sop_0_0_0_1_6_8_o5_7));
defparam un84_sop_0_0_0_1_6_8_o5_7_cZ.INIT=8'hE8;
  LUT3 un84_sop_0_0_0_1_6_8_o5_6_cZ(.I0(un84_sop_0_0_0_10_0[9:9]),.I1(x_4[6:6]),.I2(x_4[4:4]),.O(un84_sop_0_0_0_1_6_8_o5_6));
defparam un84_sop_0_0_0_1_6_8_o5_6_cZ.INIT=8'hE8;
  LUT3 un84_sop_0_0_0_1_6_8_o5_5_cZ(.I0(un84_sop_0_0_0_10_0[8:8]),.I1(x_4[3:3]),.I2(x_4[5:5]),.O(un84_sop_0_0_0_1_6_8_o5_5));
defparam un84_sop_0_0_0_1_6_8_o5_5_cZ.INIT=8'hE8;
  LUT3 un84_sop_0_0_0_1_6_8_o5_4_cZ(.I0(un84_sop_0_0_0_10_0[7:7]),.I1(x_4[2:2]),.I2(x_4[4:4]),.O(un84_sop_0_0_0_1_6_8_o5_4));
defparam un84_sop_0_0_0_1_6_8_o5_4_cZ.INIT=8'hE8;
  LUT3 un84_sop_0_0_0_1_6_8_o5_3_cZ(.I0(un84_sop_0_0_0_10_0[6:6]),.I1(x_4[1:1]),.I2(x_4[3:3]),.O(un84_sop_0_0_0_1_6_8_o5_3));
defparam un84_sop_0_0_0_1_6_8_o5_3_cZ.INIT=8'hE8;
  LUT3 un84_sop_1_6_0_o5_11_cZ(.I0(un1_x_1[15:15]),.I1(un1_x_3[15:15]),.I2(un1_x_2[15:15]),.O(un84_sop_1_6_0_o5_11));
defparam un84_sop_1_6_0_o5_11_cZ.INIT=8'hE8;
  LUT3 un84_sop_1_6_0_o5_10_cZ(.I0(un1_x_1[14:14]),.I1(un1_x_3[14:14]),.I2(un1_x_2[15:15]),.O(un84_sop_1_6_0_o5_10));
defparam un84_sop_1_6_0_o5_10_cZ.INIT=8'hE8;
  LUT3 un84_sop_1_6_0_o5_9_cZ(.I0(un1_x_1[13:13]),.I1(un1_x_2[14:14]),.I2(un1_x_3[13:13]),.O(un84_sop_1_6_0_o5_9));
defparam un84_sop_1_6_0_o5_9_cZ.INIT=8'hE8;
  LUT3 un84_sop_1_6_0_o5_8_cZ(.I0(un1_x_1[12:12]),.I1(un1_x_2[13:13]),.I2(un1_x_3[12:12]),.O(un84_sop_1_6_0_o5_8));
defparam un84_sop_1_6_0_o5_8_cZ.INIT=8'hE8;
  LUT3 un84_sop_1_6_0_o5_7_cZ(.I0(un1_x_1[11:11]),.I1(un1_x_2[12:12]),.I2(un1_x_3[11:11]),.O(un84_sop_1_6_0_o5_7));
defparam un84_sop_1_6_0_o5_7_cZ.INIT=8'hE8;
  LUT3 un84_sop_1_6_0_o5_6_cZ(.I0(un1_x_1[10:10]),.I1(un1_x_2[11:11]),.I2(un1_x_3[10:10]),.O(un84_sop_1_6_0_o5_6));
defparam un84_sop_1_6_0_o5_6_cZ.INIT=8'hE8;
  LUT3 un84_sop_1_6_0_o5_5_cZ(.I0(un1_x_1[9:9]),.I1(un1_x_2[10:10]),.I2(un1_x_3[9:9]),.O(un84_sop_1_6_0_o5_5));
defparam un84_sop_1_6_0_o5_5_cZ.INIT=8'hE8;
  LUT3 un84_sop_1_6_0_o5_4_cZ(.I0(un1_x_1[8:8]),.I1(un1_x_2[9:9]),.I2(un1_x_3[8:8]),.O(un84_sop_1_6_0_o5_4));
defparam un84_sop_1_6_0_o5_4_cZ.INIT=8'hE8;
  LUT3 un84_sop_1_6_0_o5_3_cZ(.I0(un1_x_1[7:7]),.I1(un1_x_2[8:8]),.I2(un1_x_3[7:7]),.O(un84_sop_1_6_0_o5_3));
defparam un84_sop_1_6_0_o5_3_cZ.INIT=8'hE8;
  LUT3 un84_sop_1_6_0_o5_2_cZ(.I0(un1_x_1[6:6]),.I1(un1_x_2[7:7]),.I2(un1_x_3[6:6]),.O(un84_sop_1_6_0_o5_2));
defparam un84_sop_1_6_0_o5_2_cZ.INIT=8'hE8;
  LUT5 un84_sop_1_4_axb_3_cZ(.I0(x_0[3:3]),.I1(x_0[2:2]),.I2(x_0[1:1]),.I3(x_0[0:0]),.I4(un84_sop_1_7[3:3]),.O(un84_sop_1_4_axb_3));
defparam un84_sop_1_4_axb_3_cZ.INIT=32'hAAA95556;
  LUT5 un1_x_10_5_ac0_7(.I0(x_8[4:4]),.I1(x_8[3:3]),.I2(x_8[2:2]),.I3(x_8[1:1]),.I4(x_8[0:0]),.O(un1_x_10_5_c5));
defparam un1_x_10_5_ac0_7.INIT=32'h00000001;
  LUT5 un1_x_10_axb_6_cZ(.I0(x_8[3:3]),.I1(x_8[2:2]),.I2(x_8[1:1]),.I3(x_8[0:0]),.I4(un1_x_10_4[6:6]),.O(un1_x_10_axb_6));
defparam un1_x_10_axb_6_cZ.INIT=32'hAAA95556;
  LUT6 un1_x_10_axb_7_cZ(.I0(x_8[4:4]),.I1(x_8[3:3]),.I2(x_8[2:2]),.I3(x_8[1:1]),.I4(x_8[0:0]),.I5(un1_x_10_4[7:7]),.O(un1_x_10_axb_7));
defparam un1_x_10_axb_7_cZ.INIT=64'hAAAAAAA955555556;
  LUT5 un84_sop_1_4_axb_6_cZ(.I0(x_0[6:6]),.I1(x_0[5:5]),.I2(x_0[4:4]),.I3(un1_x_0_0_c4),.I4(un84_sop_1_7[6:6]),.O(un84_sop_1_4_axb_6));
defparam un84_sop_1_4_axb_6_cZ.INIT=32'hA9AA5655;
  LUT6 un84_sop_1_4_axb_7_cZ(.I0(x_0[7:7]),.I1(x_0[6:6]),.I2(x_0[5:5]),.I3(x_0[4:4]),.I4(un1_x_0_0_c4),.I5(un84_sop_1_7[7:7]),.O(un84_sop_1_4_axb_7));
defparam un84_sop_1_4_axb_7_cZ.INIT=64'hAAA9AAAA55565555;
  LUT6 un84_sop_1_4_axb_14_cZ(.I0(x_0[7:7]),.I1(x_0[6:6]),.I2(x_0[5:5]),.I3(x_0[4:4]),.I4(un1_x_0_0_c4),.I5(un84_sop_1_7[14:14]),.O(un84_sop_1_4_axb_14));
defparam un84_sop_1_4_axb_14_cZ.INIT=64'hAAABAAAA55545555;
  LUT6 un84_sop_1_4_axb_13_cZ(.I0(x_0[7:7]),.I1(x_0[6:6]),.I2(x_0[5:5]),.I3(x_0[4:4]),.I4(un1_x_0_0_c4),.I5(un84_sop_1_7[13:13]),.O(un84_sop_1_4_axb_13));
defparam un84_sop_1_4_axb_13_cZ.INIT=64'hAAABAAAA55545555;
  LUT6 un84_sop_1_4_axb_12_cZ(.I0(x_0[7:7]),.I1(x_0[6:6]),.I2(x_0[5:5]),.I3(x_0[4:4]),.I4(un1_x_0_0_c4),.I5(un84_sop_1_7[12:12]),.O(un84_sop_1_4_axb_12));
defparam un84_sop_1_4_axb_12_cZ.INIT=64'hAAABAAAA55545555;
  LUT6 un84_sop_1_4_axb_11_cZ(.I0(x_0[7:7]),.I1(x_0[6:6]),.I2(x_0[5:5]),.I3(x_0[4:4]),.I4(un1_x_0_0_c4),.I5(un84_sop_1_7[11:11]),.O(un84_sop_1_4_axb_11));
defparam un84_sop_1_4_axb_11_cZ.INIT=64'hAAABAAAA55545555;
  LUT6 un84_sop_1_4_axb_10_cZ(.I0(x_0[7:7]),.I1(x_0[6:6]),.I2(x_0[5:5]),.I3(x_0[4:4]),.I4(un1_x_0_0_c4),.I5(un84_sop_1_7[10:10]),.O(un84_sop_1_4_axb_10));
defparam un84_sop_1_4_axb_10_cZ.INIT=64'hAAABAAAA55545555;
  LUT6 un84_sop_1_4_axb_9_cZ(.I0(x_0[7:7]),.I1(x_0[6:6]),.I2(x_0[5:5]),.I3(x_0[4:4]),.I4(un1_x_0_0_c4),.I5(un84_sop_1_7[9:9]),.O(un84_sop_1_4_axb_9));
defparam un84_sop_1_4_axb_9_cZ.INIT=64'hAAABAAAA55545555;
  LUT6 un84_sop_1_4_axb_8_cZ(.I0(x_0[7:7]),.I1(x_0[6:6]),.I2(x_0[5:5]),.I3(x_0[4:4]),.I4(un1_x_0_0_c4),.I5(un84_sop_1_7[8:8]),.O(un84_sop_1_4_axb_8));
defparam un84_sop_1_4_axb_8_cZ.INIT=64'hAAABAAAA55545555;
  LUT2 x_16_pipe_0_0_0_RNI0KBH(.I0(un84_sop_0_0_0_0_5[0:0]),.I1(un1_x_4[2:2]),.O(un84_sop_1_7[0:0]));
defparam x_16_pipe_0_0_0_RNI0KBH.INIT=4'h6;
  XORCY un84_sop_0_0_0_1_s_9(.LI(un84_sop_0_0_0_1_axb_9),.CI(un84_sop_0_0_0_1_cry_8),.O(un84_sop_0_0_0_0_1[9:9]));
  XORCY un84_sop_0_0_0_1_s_8(.LI(un84_sop_0_0_0_1_axb_8),.CI(un84_sop_0_0_0_1_cry_7),.O(un84_sop_0_0_0_0_1[8:8]));
  MUXCY_L un84_sop_0_0_0_1_cry_8_cZ(.DI(un1_x_15_0_0_0[14:14]),.CI(un84_sop_0_0_0_1_cry_7),.S(un84_sop_0_0_0_1_axb_8),.LO(un84_sop_0_0_0_1_cry_8));
  XORCY un84_sop_0_0_0_1_s_7(.LI(un84_sop_0_0_0_1_axb_7),.CI(un84_sop_0_0_0_1_cry_6),.O(un84_sop_0_0_0_0_1[7:7]));
  MUXCY_L un84_sop_0_0_0_1_cry_7_cZ(.DI(un1_x_15_0_0_0[13:13]),.CI(un84_sop_0_0_0_1_cry_6),.S(un84_sop_0_0_0_1_axb_7),.LO(un84_sop_0_0_0_1_cry_7));
  XORCY un84_sop_0_0_0_1_s_6(.LI(un84_sop_0_0_0_1_axb_6),.CI(un84_sop_0_0_0_1_cry_5),.O(un84_sop_0_0_0_0_1[6:6]));
  MUXCY_L un84_sop_0_0_0_1_cry_6_cZ(.DI(un1_x_15_0_0_0[12:12]),.CI(un84_sop_0_0_0_1_cry_5),.S(un84_sop_0_0_0_1_axb_6),.LO(un84_sop_0_0_0_1_cry_6));
  XORCY un84_sop_0_0_0_1_s_5(.LI(un84_sop_0_0_0_1_axb_5),.CI(un84_sop_0_0_0_1_cry_4),.O(un84_sop_0_0_0_0_1[5:5]));
  MUXCY_L un84_sop_0_0_0_1_cry_5_cZ(.DI(un1_x_15_0_0_0[11:11]),.CI(un84_sop_0_0_0_1_cry_4),.S(un84_sop_0_0_0_1_axb_5),.LO(un84_sop_0_0_0_1_cry_5));
  XORCY un84_sop_0_0_0_1_s_4(.LI(un84_sop_0_0_0_1_axb_4),.CI(un84_sop_0_0_0_1_cry_3),.O(un84_sop_0_0_0_0_1[4:4]));
  MUXCY_L un84_sop_0_0_0_1_cry_4_cZ(.DI(un1_x_15_0_0_0[10:10]),.CI(un84_sop_0_0_0_1_cry_3),.S(un84_sop_0_0_0_1_axb_4),.LO(un84_sop_0_0_0_1_cry_4));
  XORCY un84_sop_0_0_0_1_s_3(.LI(un84_sop_0_0_0_1_axb_3),.CI(un84_sop_0_0_0_1_cry_2),.O(un84_sop_0_0_0_0_1[3:3]));
  MUXCY_L un84_sop_0_0_0_1_cry_3_cZ(.DI(un1_x_15_0_0_0[9:9]),.CI(un84_sop_0_0_0_1_cry_2),.S(un84_sop_0_0_0_1_axb_3),.LO(un84_sop_0_0_0_1_cry_3));
  XORCY un84_sop_0_0_0_1_s_2(.LI(un84_sop_0_0_0_1_axb_2),.CI(un84_sop_0_0_0_1_cry_1),.O(un84_sop_0_0_0_0_1[2:2]));
  MUXCY_L un84_sop_0_0_0_1_cry_2_cZ(.DI(un1_x_15_0_0_0[8:8]),.CI(un84_sop_0_0_0_1_cry_1),.S(un84_sop_0_0_0_1_axb_2),.LO(un84_sop_0_0_0_1_cry_2));
  XORCY un84_sop_0_0_0_1_s_1(.LI(un84_sop_0_0_0_1_axb_1),.CI(un84_sop_0_0_0_1_cry_0),.O(un84_sop_0_0_0_0_1[1:1]));
  MUXCY_L un84_sop_0_0_0_1_cry_1_cZ(.DI(un1_x_15_0_0_0[7:7]),.CI(un84_sop_0_0_0_1_cry_0),.S(un84_sop_0_0_0_1_axb_1),.LO(un84_sop_0_0_0_1_cry_1));
  MUXCY_L un84_sop_0_0_0_1_cry_0_cZ(.DI(x_13[0:0]),.CI(GND),.S(un84_sop_0_0_0_0_1[0:0]),.LO(un84_sop_0_0_0_1_cry_0));
  XORCY un1_x_16_0_s_8(.LI(un1_x_16_0_axb_8),.CI(un1_x_16_0_cry_7),.O(un1_x_16_0_0_0[14:14]));
  XORCY un1_x_16_0_s_7(.LI(un1_x_16_0_axb_7),.CI(un1_x_16_0_cry_6),.O(un1_x_16_0_0_0[13:13]));
  MUXCY_L un1_x_16_0_cry_7_cZ(.DI(GND),.CI(un1_x_16_0_cry_6),.S(un1_x_16_0_axb_7),.LO(un1_x_16_0_cry_7));
  XORCY un1_x_16_0_s_6(.LI(un1_x_16_0_axb_6),.CI(un1_x_16_0_cry_5),.O(un1_x_16_0_0_0[12:12]));
  MUXCY_L un1_x_16_0_cry_6_cZ(.DI(GND),.CI(un1_x_16_0_cry_5),.S(un1_x_16_0_axb_6),.LO(un1_x_16_0_cry_6));
  XORCY un1_x_16_0_s_5(.LI(un1_x_16_0_axb_5),.CI(un1_x_16_0_cry_4),.O(un1_x_16_0_0_0[11:11]));
  MUXCY_L un1_x_16_0_cry_5_cZ(.DI(GND),.CI(un1_x_16_0_cry_4),.S(un1_x_16_0_axb_5),.LO(un1_x_16_0_cry_5));
  XORCY un1_x_16_0_s_4(.LI(un1_x_16_0_axb_4),.CI(un1_x_16_0_cry_3),.O(un1_x_16_0_0_0[10:10]));
  MUXCY_L un1_x_16_0_cry_4_cZ(.DI(GND),.CI(un1_x_16_0_cry_3),.S(un1_x_16_0_axb_4),.LO(un1_x_16_0_cry_4));
  XORCY un1_x_16_0_s_3(.LI(un1_x_16_0_axb_3),.CI(un1_x_16_0_cry_2),.O(un1_x_16_0_0_0[9:9]));
  MUXCY_L un1_x_16_0_cry_3_cZ(.DI(GND),.CI(un1_x_16_0_cry_2),.S(un1_x_16_0_axb_3),.LO(un1_x_16_0_cry_3));
  XORCY un1_x_16_0_s_2(.LI(un1_x_16_0_axb_2),.CI(un1_x_16_0_cry_1),.O(un1_x_16_0_0_0[8:8]));
  MUXCY_L un1_x_16_0_cry_2_cZ(.DI(GND),.CI(un1_x_16_0_cry_1),.S(un1_x_16_0_axb_2),.LO(un1_x_16_0_cry_2));
  XORCY un1_x_16_0_s_1(.LI(un1_x_16_0_axb_1),.CI(un1_x_16_0_cry_0),.O(un1_x_16_0_0_0[7:7]));
  MUXCY_L un1_x_16_0_cry_1_cZ(.DI(GND),.CI(un1_x_16_0_cry_0),.S(un1_x_16_0_axb_1),.LO(un1_x_16_0_cry_1));
  MUXCY_L un1_x_16_0_cry_0_cZ(.DI(GND),.CI(VCC),.S(un1_x_16_0_axb_0),.LO(un1_x_16_0_cry_0));
  XORCY un1_x_11_0_s_8(.LI(un1_x_11_0_axb_8),.CI(un1_x_11_0_cry_7),.O(un1_x_11_0_0_0[14:14]));
  XORCY un1_x_11_0_s_7(.LI(un1_x_11_0_axb_7),.CI(un1_x_11_0_cry_6),.O(un1_x_11_0_0_0[13:13]));
  MUXCY_L un1_x_11_0_cry_7_cZ(.DI(GND),.CI(un1_x_11_0_cry_6),.S(un1_x_11_0_axb_7),.LO(un1_x_11_0_cry_7));
  XORCY un1_x_11_0_s_6(.LI(un1_x_11_0_axb_6),.CI(un1_x_11_0_cry_5),.O(un1_x_11_0_0_0[12:12]));
  MUXCY_L un1_x_11_0_cry_6_cZ(.DI(GND),.CI(un1_x_11_0_cry_5),.S(un1_x_11_0_axb_6),.LO(un1_x_11_0_cry_6));
  XORCY un1_x_11_0_s_5(.LI(un1_x_11_0_axb_5),.CI(un1_x_11_0_cry_4),.O(un1_x_11_0_0_0[11:11]));
  MUXCY_L un1_x_11_0_cry_5_cZ(.DI(GND),.CI(un1_x_11_0_cry_4),.S(un1_x_11_0_axb_5),.LO(un1_x_11_0_cry_5));
  XORCY un1_x_11_0_s_4(.LI(un1_x_11_0_axb_4),.CI(un1_x_11_0_cry_3),.O(un1_x_11_0_0_0[10:10]));
  MUXCY_L un1_x_11_0_cry_4_cZ(.DI(GND),.CI(un1_x_11_0_cry_3),.S(un1_x_11_0_axb_4),.LO(un1_x_11_0_cry_4));
  XORCY un1_x_11_0_s_3(.LI(un1_x_11_0_axb_3),.CI(un1_x_11_0_cry_2),.O(un1_x_11_0_0_0[9:9]));
  MUXCY_L un1_x_11_0_cry_3_cZ(.DI(GND),.CI(un1_x_11_0_cry_2),.S(un1_x_11_0_axb_3),.LO(un1_x_11_0_cry_3));
  XORCY un1_x_11_0_s_2(.LI(un1_x_11_0_axb_2),.CI(un1_x_11_0_cry_1),.O(un1_x_11_0_0_0[8:8]));
  MUXCY_L un1_x_11_0_cry_2_cZ(.DI(GND),.CI(un1_x_11_0_cry_1),.S(un1_x_11_0_axb_2),.LO(un1_x_11_0_cry_2));
  XORCY un1_x_11_0_s_1(.LI(un1_x_11_0_axb_1),.CI(un1_x_11_0_cry_0),.O(un1_x_11_0_0_0[7:7]));
  MUXCY_L un1_x_11_0_cry_1_cZ(.DI(GND),.CI(un1_x_11_0_cry_0),.S(un1_x_11_0_axb_1),.LO(un1_x_11_0_cry_1));
  MUXCY_L un1_x_11_0_cry_0_cZ(.DI(GND),.CI(VCC),.S(un1_x_11_0_axb_0),.LO(un1_x_11_0_cry_0));
  XORCY un1_x_15_0_s_8(.LI(un1_x_15_0_axb_8),.CI(un1_x_15_0_cry_7),.O(un1_x_15_0_0_0[14:14]));
  XORCY un1_x_15_0_s_7(.LI(un1_x_15_0_axb_7),.CI(un1_x_15_0_cry_6),.O(un1_x_15_0_0_0[13:13]));
  MUXCY_L un1_x_15_0_cry_7_cZ(.DI(GND),.CI(un1_x_15_0_cry_6),.S(un1_x_15_0_axb_7),.LO(un1_x_15_0_cry_7));
  XORCY un1_x_15_0_s_6(.LI(un1_x_15_0_axb_6),.CI(un1_x_15_0_cry_5),.O(un1_x_15_0_0_0[12:12]));
  MUXCY_L un1_x_15_0_cry_6_cZ(.DI(GND),.CI(un1_x_15_0_cry_5),.S(un1_x_15_0_axb_6),.LO(un1_x_15_0_cry_6));
  XORCY un1_x_15_0_s_5(.LI(un1_x_15_0_axb_5),.CI(un1_x_15_0_cry_4),.O(un1_x_15_0_0_0[11:11]));
  MUXCY_L un1_x_15_0_cry_5_cZ(.DI(GND),.CI(un1_x_15_0_cry_4),.S(un1_x_15_0_axb_5),.LO(un1_x_15_0_cry_5));
  XORCY un1_x_15_0_s_4(.LI(un1_x_15_0_axb_4),.CI(un1_x_15_0_cry_3),.O(un1_x_15_0_0_0[10:10]));
  MUXCY_L un1_x_15_0_cry_4_cZ(.DI(GND),.CI(un1_x_15_0_cry_3),.S(un1_x_15_0_axb_4),.LO(un1_x_15_0_cry_4));
  XORCY un1_x_15_0_s_3(.LI(un1_x_15_0_axb_3),.CI(un1_x_15_0_cry_2),.O(un1_x_15_0_0_0[9:9]));
  MUXCY_L un1_x_15_0_cry_3_cZ(.DI(GND),.CI(un1_x_15_0_cry_2),.S(un1_x_15_0_axb_3),.LO(un1_x_15_0_cry_3));
  XORCY un1_x_15_0_s_2(.LI(un1_x_15_0_axb_2),.CI(un1_x_15_0_cry_1),.O(un1_x_15_0_0_0[8:8]));
  MUXCY_L un1_x_15_0_cry_2_cZ(.DI(GND),.CI(un1_x_15_0_cry_1),.S(un1_x_15_0_axb_2),.LO(un1_x_15_0_cry_2));
  XORCY un1_x_15_0_s_1(.LI(un1_x_15_0_axb_1),.CI(un1_x_15_0_cry_0),.O(un1_x_15_0_0_0[7:7]));
  MUXCY_L un1_x_15_0_cry_1_cZ(.DI(GND),.CI(un1_x_15_0_cry_0),.S(un1_x_15_0_axb_1),.LO(un1_x_15_0_cry_1));
  MUXCY_L un1_x_15_0_cry_0_cZ(.DI(GND),.CI(VCC),.S(un1_x_15_0_axb_0),.LO(un1_x_15_0_cry_0));
  XORCY un1_x_10_4_s_8(.LI(un1_x_10_4_s_8_false),.CI(un1_x_10_4_cry_7),.O(un1_x_10_4[8:8]));
  XORCY un1_x_10_4_s_7(.LI(un1_x_10_4_axb_7),.CI(un1_x_10_4_cry_6),.O(un1_x_10_4[7:7]));
  MUXCY_L un1_x_10_4_cry_7_cZ(.DI(x_8[6:6]),.CI(un1_x_10_4_cry_6),.S(un1_x_10_4_axb_7),.LO(un1_x_10_4_cry_7));
  XORCY un1_x_10_4_s_6(.LI(un1_x_10_4_axb_6),.CI(un1_x_10_4_cry_5),.O(un1_x_10_4[6:6]));
  MUXCY_L un1_x_10_4_cry_6_cZ(.DI(x_8[5:5]),.CI(un1_x_10_4_cry_5),.S(un1_x_10_4_axb_6),.LO(un1_x_10_4_cry_6));
  XORCY un1_x_10_4_s_5(.LI(un1_x_10_4_axb_5),.CI(un1_x_10_4_cry_4),.O(un1_x_10_4[5:5]));
  MUXCY_L un1_x_10_4_cry_5_cZ(.DI(x_8[4:4]),.CI(un1_x_10_4_cry_4),.S(un1_x_10_4_axb_5),.LO(un1_x_10_4_cry_5));
  XORCY un1_x_10_4_s_4(.LI(un1_x_10_4_axb_4),.CI(un1_x_10_4_cry_3),.O(un1_x_10_4[4:4]));
  MUXCY_L un1_x_10_4_cry_4_cZ(.DI(x_8[3:3]),.CI(un1_x_10_4_cry_3),.S(un1_x_10_4_axb_4),.LO(un1_x_10_4_cry_4));
  XORCY un1_x_10_4_s_3(.LI(un1_x_10_4_axb_3),.CI(un1_x_10_4_cry_2),.O(un1_x_10_4[3:3]));
  MUXCY_L un1_x_10_4_cry_3_cZ(.DI(x_8[2:2]),.CI(un1_x_10_4_cry_2),.S(un1_x_10_4_axb_3),.LO(un1_x_10_4_cry_3));
  XORCY un1_x_10_4_s_2(.LI(un1_x_10_4_axb_2),.CI(un1_x_10_4_cry_1),.O(un1_x_10_4[2:2]));
  MUXCY_L un1_x_10_4_cry_2_cZ(.DI(x_8[1:1]),.CI(un1_x_10_4_cry_1),.S(un1_x_10_4_axb_2),.LO(un1_x_10_4_cry_2));
  MUXCY_L un1_x_10_4_cry_1_cZ(.DI(x_8[0:0]),.CI(GND),.S(un1_x_10_4_cry_1_sf),.LO(un1_x_10_4_cry_1));
  XORCY un84_sop_1_s_14_cZ(.LI(un84_sop_1_axb_14),.CI(un84_sop_1_cry_13),.O(un84_sop_1_s_14));
  XORCY un84_sop_1_s_13_cZ(.LI(un84_sop_1_axb_13),.CI(un84_sop_1_cry_12),.O(un84_sop_1_s_13));
  MUXCY_L un84_sop_1_cry_13_cZ(.DI(un84_sop_1_4[13:13]),.CI(un84_sop_1_cry_12),.S(un84_sop_1_axb_13),.LO(un84_sop_1_cry_13));
  XORCY un84_sop_1_s_12_cZ(.LI(un84_sop_1_axb_12),.CI(un84_sop_1_cry_11),.O(un84_sop_1_s_12));
  MUXCY_L un84_sop_1_cry_12_cZ(.DI(un84_sop_1_4[12:12]),.CI(un84_sop_1_cry_11),.S(un84_sop_1_axb_12),.LO(un84_sop_1_cry_12));
  XORCY un84_sop_1_s_11_cZ(.LI(un84_sop_1_axb_11),.CI(un84_sop_1_cry_10),.O(un84_sop_1_s_11));
  MUXCY_L un84_sop_1_cry_11_cZ(.DI(un84_sop_1_4[11:11]),.CI(un84_sop_1_cry_10),.S(un84_sop_1_axb_11),.LO(un84_sop_1_cry_11));
  XORCY un84_sop_1_s_10_cZ(.LI(un84_sop_1_axb_10),.CI(un84_sop_1_cry_9),.O(un84_sop_1_s_10));
  MUXCY_L un84_sop_1_cry_10_cZ(.DI(un84_sop_1_4[10:10]),.CI(un84_sop_1_cry_9),.S(un84_sop_1_axb_10),.LO(un84_sop_1_cry_10));
  XORCY un84_sop_1_s_9_cZ(.LI(un84_sop_1_axb_9),.CI(un84_sop_1_cry_8),.O(un84_sop_1_s_9));
  MUXCY_L un84_sop_1_cry_9_cZ(.DI(un84_sop_1_4[9:9]),.CI(un84_sop_1_cry_8),.S(un84_sop_1_axb_9),.LO(un84_sop_1_cry_9));
  XORCY un84_sop_1_s_8_cZ(.LI(un84_sop_1_axb_8),.CI(un84_sop_1_cry_7),.O(un84_sop_1_s_8));
  MUXCY_L un84_sop_1_cry_8_cZ(.DI(un84_sop_1_4[8:8]),.CI(un84_sop_1_cry_7),.S(un84_sop_1_axb_8),.LO(un84_sop_1_cry_8));
  XORCY un84_sop_1_s_7_cZ(.LI(un84_sop_1_axb_7),.CI(un84_sop_1_cry_6),.O(un84_sop_1_s_7));
  MUXCY_L un84_sop_1_cry_7_cZ(.DI(un84_sop_1_4[7:7]),.CI(un84_sop_1_cry_6),.S(un84_sop_1_axb_7),.LO(un84_sop_1_cry_7));
  MUXCY_L un84_sop_1_cry_6_cZ(.DI(un84_sop_1_4[6:6]),.CI(un84_sop_1_cry_5),.S(un84_sop_1_axb_6),.LO(un84_sop_1_cry_6));
  MUXCY_L un84_sop_1_cry_5_cZ(.DI(un84_sop_1_4[5:5]),.CI(un84_sop_1_cry_4),.S(un84_sop_1_axb_5),.LO(un84_sop_1_cry_5));
  MUXCY_L un84_sop_1_cry_4_cZ(.DI(un84_sop_1_4[4:4]),.CI(un84_sop_1_cry_3),.S(un84_sop_1_axb_4),.LO(un84_sop_1_cry_4));
  MUXCY_L un84_sop_1_cry_3_cZ(.DI(un84_sop_1_4[3:3]),.CI(un84_sop_1_cry_2),.S(un84_sop_1_axb_3),.LO(un84_sop_1_cry_3));
  MUXCY_L un84_sop_1_cry_2_cZ(.DI(un84_sop_1_4[2:2]),.CI(un84_sop_1_cry_1),.S(un84_sop_1_axb_2),.LO(un84_sop_1_cry_2));
  MUXCY_L un84_sop_1_cry_1_cZ(.DI(un84_sop_1_4[1:1]),.CI(un84_sop_1_cry_0),.S(un84_sop_1_axb_1),.LO(un84_sop_1_cry_1));
  MUXCY_L un84_sop_1_cry_0_cZ(.DI(un84_sop_1_6[0:0]),.CI(GND),.S(un84_sop_1_axb_0),.LO(un84_sop_1_cry_0));
  XORCY un84_sop_1_4_s_14(.LI(un84_sop_1_4_axb_14),.CI(un84_sop_1_4_cry_13),.O(un84_sop_1_4[14:14]));
  XORCY un84_sop_1_4_s_13(.LI(un84_sop_1_4_axb_13),.CI(un84_sop_1_4_cry_12),.O(un84_sop_1_4[13:13]));
  MUXCY_L un84_sop_1_4_cry_13_cZ(.DI(un84_sop_1_7[13:13]),.CI(un84_sop_1_4_cry_12),.S(un84_sop_1_4_axb_13),.LO(un84_sop_1_4_cry_13));
  XORCY un84_sop_1_4_s_12(.LI(un84_sop_1_4_axb_12),.CI(un84_sop_1_4_cry_11),.O(un84_sop_1_4[12:12]));
  MUXCY_L un84_sop_1_4_cry_12_cZ(.DI(un84_sop_1_7[12:12]),.CI(un84_sop_1_4_cry_11),.S(un84_sop_1_4_axb_12),.LO(un84_sop_1_4_cry_12));
  XORCY un84_sop_1_4_s_11(.LI(un84_sop_1_4_axb_11),.CI(un84_sop_1_4_cry_10),.O(un84_sop_1_4[11:11]));
  MUXCY_L un84_sop_1_4_cry_11_cZ(.DI(un84_sop_1_7[11:11]),.CI(un84_sop_1_4_cry_10),.S(un84_sop_1_4_axb_11),.LO(un84_sop_1_4_cry_11));
  XORCY un84_sop_1_4_s_10(.LI(un84_sop_1_4_axb_10),.CI(un84_sop_1_4_cry_9),.O(un84_sop_1_4[10:10]));
  MUXCY_L un84_sop_1_4_cry_10_cZ(.DI(un84_sop_1_7[10:10]),.CI(un84_sop_1_4_cry_9),.S(un84_sop_1_4_axb_10),.LO(un84_sop_1_4_cry_10));
  XORCY un84_sop_1_4_s_9(.LI(un84_sop_1_4_axb_9),.CI(un84_sop_1_4_cry_8),.O(un84_sop_1_4[9:9]));
  MUXCY_L un84_sop_1_4_cry_9_cZ(.DI(un84_sop_1_7[9:9]),.CI(un84_sop_1_4_cry_8),.S(un84_sop_1_4_axb_9),.LO(un84_sop_1_4_cry_9));
  XORCY un84_sop_1_4_s_8(.LI(un84_sop_1_4_axb_8),.CI(un84_sop_1_4_cry_7),.O(un84_sop_1_4[8:8]));
  MUXCY_L un84_sop_1_4_cry_8_cZ(.DI(un84_sop_1_7[8:8]),.CI(un84_sop_1_4_cry_7),.S(un84_sop_1_4_axb_8),.LO(un84_sop_1_4_cry_8));
  XORCY un84_sop_1_4_s_7(.LI(un84_sop_1_4_axb_7),.CI(un84_sop_1_4_cry_6),.O(un84_sop_1_4[7:7]));
  MUXCY_L un84_sop_1_4_cry_7_cZ(.DI(un84_sop_1_7[7:7]),.CI(un84_sop_1_4_cry_6),.S(un84_sop_1_4_axb_7),.LO(un84_sop_1_4_cry_7));
  XORCY un84_sop_1_4_s_6(.LI(un84_sop_1_4_axb_6),.CI(un84_sop_1_4_cry_5),.O(un84_sop_1_4[6:6]));
  MUXCY_L un84_sop_1_4_cry_6_cZ(.DI(un84_sop_1_7[6:6]),.CI(un84_sop_1_4_cry_5),.S(un84_sop_1_4_axb_6),.LO(un84_sop_1_4_cry_6));
  XORCY un84_sop_1_4_s_5(.LI(un84_sop_1_4_axb_5),.CI(un84_sop_1_4_cry_4),.O(un84_sop_1_4[5:5]));
  MUXCY_L un84_sop_1_4_cry_5_cZ(.DI(un84_sop_1_7[5:5]),.CI(un84_sop_1_4_cry_4),.S(un84_sop_1_4_axb_5),.LO(un84_sop_1_4_cry_5));
  XORCY un84_sop_1_4_s_4(.LI(un84_sop_1_4_axb_4),.CI(un84_sop_1_4_cry_3),.O(un84_sop_1_4[4:4]));
  MUXCY_L un84_sop_1_4_cry_4_cZ(.DI(un84_sop_1_7[4:4]),.CI(un84_sop_1_4_cry_3),.S(un84_sop_1_4_axb_4),.LO(un84_sop_1_4_cry_4));
  XORCY un84_sop_1_4_s_3(.LI(un84_sop_1_4_axb_3),.CI(un84_sop_1_4_cry_2),.O(un84_sop_1_4[3:3]));
  MUXCY_L un84_sop_1_4_cry_3_cZ(.DI(un84_sop_1_7[3:3]),.CI(un84_sop_1_4_cry_2),.S(un84_sop_1_4_axb_3),.LO(un84_sop_1_4_cry_3));
  XORCY un84_sop_1_4_s_2(.LI(un84_sop_1_4_axb_2),.CI(un84_sop_1_4_cry_1),.O(un84_sop_1_4[2:2]));
  MUXCY_L un84_sop_1_4_cry_2_cZ(.DI(un84_sop_1_7[2:2]),.CI(un84_sop_1_4_cry_1),.S(un84_sop_1_4_axb_2),.LO(un84_sop_1_4_cry_2));
  XORCY un84_sop_1_4_s_1(.LI(un84_sop_1_4_axb_1),.CI(un84_sop_1_4_cry_0),.O(un84_sop_1_4[1:1]));
  MUXCY_L un84_sop_1_4_cry_1_cZ(.DI(un84_sop_1_7[1:1]),.CI(un84_sop_1_4_cry_0),.S(un84_sop_1_4_axb_1),.LO(un84_sop_1_4_cry_1));
  MUXCY_L un84_sop_1_4_cry_0_cZ(.DI(un84_sop_1_7[0:0]),.CI(GND),.S(un84_sop_1_4[0:0]),.LO(un84_sop_1_4_cry_0));
  XORCY un84_sop_0_0_0_0_11_7_s_10(.LI(un84_sop_0_0_0_0_11_7_axb_10),.CI(un84_sop_0_0_0_0_11_7_cry_9),.O(un84_sop_0_0_0_0_11_7[14:14]));
  XORCY un84_sop_0_0_0_0_11_7_s_9(.LI(un84_sop_0_0_0_0_11_7_axb_9),.CI(un84_sop_0_0_0_0_11_7_cry_8),.O(un84_sop_0_0_0_0_11_7[9:9]));
  MUXCY_L un84_sop_0_0_0_0_11_7_cry_9_cZ(.DI(un84_sop_0_0_0_0_0[9:9]),.CI(un84_sop_0_0_0_0_11_7_cry_8),.S(un84_sop_0_0_0_0_11_7_axb_9),.LO(un84_sop_0_0_0_0_11_7_cry_9));
  XORCY un84_sop_0_0_0_0_11_7_s_8(.LI(un84_sop_0_0_0_0_11_7_axb_8),.CI(un84_sop_0_0_0_0_11_7_cry_7),.O(un84_sop_0_0_0_0_11_7[8:8]));
  MUXCY_L un84_sop_0_0_0_0_11_7_cry_8_cZ(.DI(un84_sop_0_0_0_0_0[8:8]),.CI(un84_sop_0_0_0_0_11_7_cry_7),.S(un84_sop_0_0_0_0_11_7_axb_8),.LO(un84_sop_0_0_0_0_11_7_cry_8));
  XORCY un84_sop_0_0_0_0_11_7_s_7(.LI(un84_sop_0_0_0_0_11_7_axb_7),.CI(un84_sop_0_0_0_0_11_7_cry_6),.O(un84_sop_0_0_0_0_11_7[7:7]));
  MUXCY_L un84_sop_0_0_0_0_11_7_cry_7_cZ(.DI(un84_sop_0_0_0_0_0[7:7]),.CI(un84_sop_0_0_0_0_11_7_cry_6),.S(un84_sop_0_0_0_0_11_7_axb_7),.LO(un84_sop_0_0_0_0_11_7_cry_7));
  XORCY un84_sop_0_0_0_0_11_7_s_6(.LI(un84_sop_0_0_0_0_11_7_axb_6),.CI(un84_sop_0_0_0_0_11_7_cry_5),.O(un84_sop_0_0_0_0_11_7[6:6]));
  MUXCY_L un84_sop_0_0_0_0_11_7_cry_6_cZ(.DI(un84_sop_0_0_0_0_0[6:6]),.CI(un84_sop_0_0_0_0_11_7_cry_5),.S(un84_sop_0_0_0_0_11_7_axb_6),.LO(un84_sop_0_0_0_0_11_7_cry_6));
  XORCY un84_sop_0_0_0_0_11_7_s_5(.LI(un84_sop_0_0_0_0_11_7_axb_5),.CI(un84_sop_0_0_0_0_11_7_cry_4),.O(un84_sop_0_0_0_0_11_7[5:5]));
  MUXCY_L un84_sop_0_0_0_0_11_7_cry_5_cZ(.DI(un84_sop_0_0_0_0_0[5:5]),.CI(un84_sop_0_0_0_0_11_7_cry_4),.S(un84_sop_0_0_0_0_11_7_axb_5),.LO(un84_sop_0_0_0_0_11_7_cry_5));
  XORCY un84_sop_0_0_0_0_11_7_s_4(.LI(un84_sop_0_0_0_0_11_7_axb_4),.CI(un84_sop_0_0_0_0_11_7_cry_3),.O(un84_sop_0_0_0_0_11_7[4:4]));
  MUXCY_L un84_sop_0_0_0_0_11_7_cry_4_cZ(.DI(un84_sop_0_0_0_0_0[4:4]),.CI(un84_sop_0_0_0_0_11_7_cry_3),.S(un84_sop_0_0_0_0_11_7_axb_4),.LO(un84_sop_0_0_0_0_11_7_cry_4));
  XORCY un84_sop_0_0_0_0_11_7_s_3(.LI(un84_sop_0_0_0_0_11_7_axb_3),.CI(un84_sop_0_0_0_0_11_7_cry_2),.O(un84_sop_0_0_0_0_11_7[3:3]));
  MUXCY_L un84_sop_0_0_0_0_11_7_cry_3_cZ(.DI(un84_sop_0_0_0_0_0[3:3]),.CI(un84_sop_0_0_0_0_11_7_cry_2),.S(un84_sop_0_0_0_0_11_7_axb_3),.LO(un84_sop_0_0_0_0_11_7_cry_3));
  XORCY un84_sop_0_0_0_0_11_7_s_2(.LI(un84_sop_0_0_0_0_11_7_axb_2),.CI(un84_sop_0_0_0_0_11_7_cry_1),.O(un84_sop_0_0_0_0_11_7[2:2]));
  MUXCY_L un84_sop_0_0_0_0_11_7_cry_2_cZ(.DI(un84_sop_0_0_0_0_0[2:2]),.CI(un84_sop_0_0_0_0_11_7_cry_1),.S(un84_sop_0_0_0_0_11_7_axb_2),.LO(un84_sop_0_0_0_0_11_7_cry_2));
  XORCY un84_sop_0_0_0_0_11_7_s_1(.LI(un84_sop_0_0_0_0_11_7_axb_1),.CI(un84_sop_0_0_0_0_11_7_cry_0),.O(un84_sop_0_0_0_0_11_7[1:1]));
  MUXCY_L un84_sop_0_0_0_0_11_7_cry_1_cZ(.DI(un84_sop_0_0_0_0_0[1:1]),.CI(un84_sop_0_0_0_0_11_7_cry_0),.S(un84_sop_0_0_0_0_11_7_axb_1),.LO(un84_sop_0_0_0_0_11_7_cry_1));
  MUXCY_L un84_sop_0_0_0_0_11_7_cry_0_cZ(.DI(un84_sop_0_0_0_0_0[0:0]),.CI(GND),.S(un84_sop_0_0_0_0_11_7[0:0]),.LO(un84_sop_0_0_0_0_11_7_cry_0));
  XORCY un84_sop_1_7_s_14(.LI(un84_sop_1_7_axb_14),.CI(un84_sop_1_7_cry_13),.O(un84_sop_1_7[14:14]));
  XORCY un84_sop_1_7_s_13(.LI(un84_sop_1_7_axb_13),.CI(un84_sop_1_7_cry_12),.O(un84_sop_1_7[13:13]));
  MUXCY_L un84_sop_1_7_cry_13_cZ(.DI(un84_sop_0_0_0_0_5[13:13]),.CI(un84_sop_1_7_cry_12),.S(un84_sop_1_7_axb_13),.LO(un84_sop_1_7_cry_13));
  XORCY un84_sop_1_7_s_12(.LI(un84_sop_1_7_axb_12),.CI(un84_sop_1_7_cry_11),.O(un84_sop_1_7[12:12]));
  MUXCY_L un84_sop_1_7_cry_12_cZ(.DI(un84_sop_0_0_0_0_5[12:12]),.CI(un84_sop_1_7_cry_11),.S(un84_sop_1_7_axb_12),.LO(un84_sop_1_7_cry_12));
  XORCY un84_sop_1_7_s_11(.LI(un84_sop_1_7_axb_11),.CI(un84_sop_1_7_cry_10),.O(un84_sop_1_7[11:11]));
  MUXCY_L un84_sop_1_7_cry_11_cZ(.DI(un84_sop_0_0_0_0_5[11:11]),.CI(un84_sop_1_7_cry_10),.S(un84_sop_1_7_axb_11),.LO(un84_sop_1_7_cry_11));
  XORCY un84_sop_1_7_s_10(.LI(un84_sop_1_7_axb_10),.CI(un84_sop_1_7_cry_9),.O(un84_sop_1_7[10:10]));
  MUXCY_L un84_sop_1_7_cry_10_cZ(.DI(un84_sop_0_0_0_0_5[10:10]),.CI(un84_sop_1_7_cry_9),.S(un84_sop_1_7_axb_10),.LO(un84_sop_1_7_cry_10));
  XORCY un84_sop_1_7_s_9(.LI(un84_sop_1_7_axb_9),.CI(un84_sop_1_7_cry_8),.O(un84_sop_1_7[9:9]));
  MUXCY_L un84_sop_1_7_cry_9_cZ(.DI(un84_sop_0_0_0_0_5[9:9]),.CI(un84_sop_1_7_cry_8),.S(un84_sop_1_7_axb_9),.LO(un84_sop_1_7_cry_9));
  XORCY un84_sop_1_7_s_8(.LI(un84_sop_1_7_axb_8),.CI(un84_sop_1_7_cry_7),.O(un84_sop_1_7[8:8]));
  MUXCY_L un84_sop_1_7_cry_8_cZ(.DI(un84_sop_0_0_0_0_5[8:8]),.CI(un84_sop_1_7_cry_7),.S(un84_sop_1_7_axb_8),.LO(un84_sop_1_7_cry_8));
  XORCY un84_sop_1_7_s_7(.LI(un84_sop_1_7_axb_7),.CI(un84_sop_1_7_cry_6),.O(un84_sop_1_7[7:7]));
  MUXCY_L un84_sop_1_7_cry_7_cZ(.DI(un84_sop_0_0_0_0_5[7:7]),.CI(un84_sop_1_7_cry_6),.S(un84_sop_1_7_axb_7),.LO(un84_sop_1_7_cry_7));
  XORCY un84_sop_1_7_s_6(.LI(un84_sop_1_7_axb_6),.CI(un84_sop_1_7_cry_5),.O(un84_sop_1_7[6:6]));
  MUXCY_L un84_sop_1_7_cry_6_cZ(.DI(un84_sop_0_0_0_0_5[6:6]),.CI(un84_sop_1_7_cry_5),.S(un84_sop_1_7_axb_6),.LO(un84_sop_1_7_cry_6));
  XORCY un84_sop_1_7_s_5(.LI(un84_sop_1_7_axb_5),.CI(un84_sop_1_7_cry_4),.O(un84_sop_1_7[5:5]));
  MUXCY_L un84_sop_1_7_cry_5_cZ(.DI(un84_sop_0_0_0_0_5[5:5]),.CI(un84_sop_1_7_cry_4),.S(un84_sop_1_7_axb_5),.LO(un84_sop_1_7_cry_5));
  XORCY un84_sop_1_7_s_4(.LI(un84_sop_1_7_axb_4),.CI(un84_sop_1_7_cry_3),.O(un84_sop_1_7[4:4]));
  MUXCY_L un84_sop_1_7_cry_4_cZ(.DI(un84_sop_0_0_0_0_5[4:4]),.CI(un84_sop_1_7_cry_3),.S(un84_sop_1_7_axb_4),.LO(un84_sop_1_7_cry_4));
  XORCY un84_sop_1_7_s_3(.LI(un84_sop_1_7_axb_3),.CI(un84_sop_1_7_cry_2),.O(un84_sop_1_7[3:3]));
  MUXCY_L un84_sop_1_7_cry_3_cZ(.DI(un84_sop_0_0_0_0_5[3:3]),.CI(un84_sop_1_7_cry_2),.S(un84_sop_1_7_axb_3),.LO(un84_sop_1_7_cry_3));
  XORCY un84_sop_1_7_s_2(.LI(un84_sop_1_7_axb_2),.CI(un84_sop_1_7_cry_1),.O(un84_sop_1_7[2:2]));
  MUXCY_L un84_sop_1_7_cry_2_cZ(.DI(un84_sop_0_0_0_0_5[2:2]),.CI(un84_sop_1_7_cry_1),.S(un84_sop_1_7_axb_2),.LO(un84_sop_1_7_cry_2));
  XORCY un84_sop_1_7_s_1(.LI(un84_sop_1_7_axb_1),.CI(un84_sop_1_7_cry_0),.O(un84_sop_1_7[1:1]));
  MUXCY_L un84_sop_1_7_cry_1_cZ(.DI(un84_sop_0_0_0_0_5[1:1]),.CI(un84_sop_1_7_cry_0),.S(un84_sop_1_7_axb_1),.LO(un84_sop_1_7_cry_1));
  MUXCY_L un84_sop_1_7_cry_0_cZ(.DI(un84_sop_0_0_0_0_5[0:0]),.CI(GND),.S(un84_sop_1_7[0:0]),.LO(un84_sop_1_7_cry_0));
  XORCY un84_sop_0_0_0_1_6_s_14(.LI(un84_sop_0_0_0_1_6_axb_14),.CI(un84_sop_0_0_0_1_6_cry_13),.O(un84_sop_0_0_0_5_0[14:14]));
  XORCY un84_sop_0_0_0_1_6_s_13(.LI(un84_sop_0_0_0_1_6_axb_13),.CI(un84_sop_0_0_0_1_6_cry_12),.O(un84_sop_0_0_0_5_0[13:13]));
  MUXCY_L un84_sop_0_0_0_1_6_cry_13_cZ(.DI(un84_sop_0_0_0_1_6_4[13:13]),.CI(un84_sop_0_0_0_1_6_cry_12),.S(un84_sop_0_0_0_1_6_axb_13),.LO(un84_sop_0_0_0_1_6_cry_13));
  XORCY un84_sop_0_0_0_1_6_s_12(.LI(un84_sop_0_0_0_1_6_axb_12),.CI(un84_sop_0_0_0_1_6_cry_11),.O(un84_sop_0_0_0_5_0[12:12]));
  MUXCY_L un84_sop_0_0_0_1_6_cry_12_cZ(.DI(un84_sop_0_0_0_1_6_4[12:12]),.CI(un84_sop_0_0_0_1_6_cry_11),.S(un84_sop_0_0_0_1_6_axb_12),.LO(un84_sop_0_0_0_1_6_cry_12));
  XORCY un84_sop_0_0_0_1_6_s_11(.LI(un84_sop_0_0_0_1_6_axb_11),.CI(un84_sop_0_0_0_1_6_cry_10),.O(un84_sop_0_0_0_5_0[11:11]));
  MUXCY_L un84_sop_0_0_0_1_6_cry_11_cZ(.DI(un84_sop_0_0_0_1_6_4[11:11]),.CI(un84_sop_0_0_0_1_6_cry_10),.S(un84_sop_0_0_0_1_6_axb_11),.LO(un84_sop_0_0_0_1_6_cry_11));
  XORCY un84_sop_0_0_0_1_6_s_10(.LI(un84_sop_0_0_0_1_6_axb_10),.CI(un84_sop_0_0_0_1_6_cry_9),.O(un84_sop_0_0_0_5_0[10:10]));
  MUXCY_L un84_sop_0_0_0_1_6_cry_10_cZ(.DI(un84_sop_0_0_0_1_6_4[10:10]),.CI(un84_sop_0_0_0_1_6_cry_9),.S(un84_sop_0_0_0_1_6_axb_10),.LO(un84_sop_0_0_0_1_6_cry_10));
  XORCY un84_sop_0_0_0_1_6_s_9(.LI(un84_sop_0_0_0_1_6_axb_9),.CI(un84_sop_0_0_0_1_6_cry_8),.O(un84_sop_0_0_0_5_0[9:9]));
  MUXCY_L un84_sop_0_0_0_1_6_cry_9_cZ(.DI(un84_sop_0_0_0_1_6_4[9:9]),.CI(un84_sop_0_0_0_1_6_cry_8),.S(un84_sop_0_0_0_1_6_axb_9),.LO(un84_sop_0_0_0_1_6_cry_9));
  XORCY un84_sop_0_0_0_1_6_s_8(.LI(un84_sop_0_0_0_1_6_axb_8),.CI(un84_sop_0_0_0_1_6_cry_7),.O(un84_sop_0_0_0_5_0[8:8]));
  MUXCY_L un84_sop_0_0_0_1_6_cry_8_cZ(.DI(un84_sop_0_0_0_1_6_4[8:8]),.CI(un84_sop_0_0_0_1_6_cry_7),.S(un84_sop_0_0_0_1_6_axb_8),.LO(un84_sop_0_0_0_1_6_cry_8));
  XORCY un84_sop_0_0_0_1_6_s_7(.LI(un84_sop_0_0_0_1_6_axb_7),.CI(un84_sop_0_0_0_1_6_cry_6),.O(un84_sop_0_0_0_5_0[7:7]));
  MUXCY_L un84_sop_0_0_0_1_6_cry_7_cZ(.DI(un84_sop_0_0_0_1_6_4[7:7]),.CI(un84_sop_0_0_0_1_6_cry_6),.S(un84_sop_0_0_0_1_6_axb_7),.LO(un84_sop_0_0_0_1_6_cry_7));
  XORCY un84_sop_0_0_0_1_6_s_6(.LI(un84_sop_0_0_0_1_6_axb_6),.CI(un84_sop_0_0_0_1_6_cry_5),.O(un84_sop_0_0_0_5_0[6:6]));
  MUXCY_L un84_sop_0_0_0_1_6_cry_6_cZ(.DI(un84_sop_0_0_0_1_6_4[6:6]),.CI(un84_sop_0_0_0_1_6_cry_5),.S(un84_sop_0_0_0_1_6_axb_6),.LO(un84_sop_0_0_0_1_6_cry_6));
  XORCY un84_sop_0_0_0_1_6_s_5(.LI(un84_sop_0_0_0_1_6_axb_5),.CI(un84_sop_0_0_0_1_6_cry_4),.O(un84_sop_0_0_0_5_0[5:5]));
  MUXCY_L un84_sop_0_0_0_1_6_cry_5_cZ(.DI(un84_sop_0_0_0_1_6_4[5:5]),.CI(un84_sop_0_0_0_1_6_cry_4),.S(un84_sop_0_0_0_1_6_axb_5),.LO(un84_sop_0_0_0_1_6_cry_5));
  XORCY un84_sop_0_0_0_1_6_s_4(.LI(un84_sop_0_0_0_1_6_axb_4),.CI(un84_sop_0_0_0_1_6_cry_3),.O(un84_sop_0_0_0_5_0[4:4]));
  MUXCY_L un84_sop_0_0_0_1_6_cry_4_cZ(.DI(un84_sop_0_0_0_1_6_4[4:4]),.CI(un84_sop_0_0_0_1_6_cry_3),.S(un84_sop_0_0_0_1_6_axb_4),.LO(un84_sop_0_0_0_1_6_cry_4));
  XORCY un84_sop_0_0_0_1_6_s_3(.LI(un84_sop_0_0_0_1_6_axb_3),.CI(un84_sop_0_0_0_1_6_cry_2),.O(un84_sop_0_0_0_5_0[3:3]));
  MUXCY_L un84_sop_0_0_0_1_6_cry_3_cZ(.DI(un84_sop_0_0_0_1_6_4[3:3]),.CI(un84_sop_0_0_0_1_6_cry_2),.S(un84_sop_0_0_0_1_6_axb_3),.LO(un84_sop_0_0_0_1_6_cry_3));
  XORCY un84_sop_0_0_0_1_6_s_2(.LI(un84_sop_0_0_0_1_6_axb_2),.CI(un84_sop_0_0_0_1_6_cry_1),.O(un84_sop_0_0_0_5_0[2:2]));
  MUXCY_L un84_sop_0_0_0_1_6_cry_2_cZ(.DI(un84_sop_0_0_0_1_6_4[2:2]),.CI(un84_sop_0_0_0_1_6_cry_1),.S(un84_sop_0_0_0_1_6_axb_2),.LO(un84_sop_0_0_0_1_6_cry_2));
  XORCY un84_sop_0_0_0_1_6_s_1(.LI(un84_sop_0_0_0_1_6_axb_1),.CI(un84_sop_0_0_0_1_6_cry_0),.O(un84_sop_0_0_0_5_0[1:1]));
  MUXCY_L un84_sop_0_0_0_1_6_cry_1_cZ(.DI(un84_sop_0_0_0_1_6_4[1:1]),.CI(un84_sop_0_0_0_1_6_cry_0),.S(un84_sop_0_0_0_1_6_axb_1),.LO(un84_sop_0_0_0_1_6_cry_1));
  MUXCY_L un84_sop_0_0_0_1_6_cry_0_cZ(.DI(un84_sop_0_0_0_1_6_6[0:0]),.CI(GND),.S(un84_sop_0_0_0_5_0[0:0]),.LO(un84_sop_0_0_0_1_6_cry_0));
  XORCY un84_sop_0_0_0_1_6_4_s_14(.LI(un84_sop_0_0_0_1_6_4_axb_14),.CI(un84_sop_0_0_0_1_6_4_cry_13),.O(un84_sop_0_0_0_1_6_4[14:14]));
  XORCY un84_sop_0_0_0_1_6_4_s_13(.LI(un84_sop_0_0_0_1_6_4_axb_13),.CI(un84_sop_0_0_0_1_6_4_cry_12),.O(un84_sop_0_0_0_1_6_4[13:13]));
  MUXCY_L un84_sop_0_0_0_1_6_4_cry_13_cZ(.DI(un84_sop_0_0_0_1_6_8[13:13]),.CI(un84_sop_0_0_0_1_6_4_cry_12),.S(un84_sop_0_0_0_1_6_4_axb_13),.LO(un84_sop_0_0_0_1_6_4_cry_13));
  XORCY un84_sop_0_0_0_1_6_4_s_12(.LI(un84_sop_0_0_0_1_6_4_axb_12),.CI(un84_sop_0_0_0_1_6_4_cry_11),.O(un84_sop_0_0_0_1_6_4[12:12]));
  MUXCY_L un84_sop_0_0_0_1_6_4_cry_12_cZ(.DI(un84_sop_0_0_0_1_6_8[12:12]),.CI(un84_sop_0_0_0_1_6_4_cry_11),.S(un84_sop_0_0_0_1_6_4_axb_12),.LO(un84_sop_0_0_0_1_6_4_cry_12));
  XORCY un84_sop_0_0_0_1_6_4_s_11(.LI(un84_sop_0_0_0_1_6_4_axb_11),.CI(un84_sop_0_0_0_1_6_4_cry_10),.O(un84_sop_0_0_0_1_6_4[11:11]));
  MUXCY_L un84_sop_0_0_0_1_6_4_cry_11_cZ(.DI(un84_sop_0_0_0_1_6_8[11:11]),.CI(un84_sop_0_0_0_1_6_4_cry_10),.S(un84_sop_0_0_0_1_6_4_axb_11),.LO(un84_sop_0_0_0_1_6_4_cry_11));
  XORCY un84_sop_0_0_0_1_6_4_s_10(.LI(un84_sop_0_0_0_1_6_4_axb_10),.CI(un84_sop_0_0_0_1_6_4_cry_9),.O(un84_sop_0_0_0_1_6_4[10:10]));
  MUXCY_L un84_sop_0_0_0_1_6_4_cry_10_cZ(.DI(un84_sop_0_0_0_1_6_8[10:10]),.CI(un84_sop_0_0_0_1_6_4_cry_9),.S(un84_sop_0_0_0_1_6_4_axb_10),.LO(un84_sop_0_0_0_1_6_4_cry_10));
  XORCY un84_sop_0_0_0_1_6_4_s_9(.LI(un84_sop_0_0_0_1_6_4_axb_9),.CI(un84_sop_0_0_0_1_6_4_cry_8),.O(un84_sop_0_0_0_1_6_4[9:9]));
  MUXCY_L un84_sop_0_0_0_1_6_4_cry_9_cZ(.DI(un84_sop_0_0_0_1_6_8[9:9]),.CI(un84_sop_0_0_0_1_6_4_cry_8),.S(un84_sop_0_0_0_1_6_4_axb_9),.LO(un84_sop_0_0_0_1_6_4_cry_9));
  XORCY un84_sop_0_0_0_1_6_4_s_8(.LI(un84_sop_0_0_0_1_6_4_axb_8),.CI(un84_sop_0_0_0_1_6_4_cry_7),.O(un84_sop_0_0_0_1_6_4[8:8]));
  MUXCY_L un84_sop_0_0_0_1_6_4_cry_8_cZ(.DI(un84_sop_0_0_0_1_6_8[8:8]),.CI(un84_sop_0_0_0_1_6_4_cry_7),.S(un84_sop_0_0_0_1_6_4_axb_8),.LO(un84_sop_0_0_0_1_6_4_cry_8));
  XORCY un84_sop_0_0_0_1_6_4_s_7(.LI(un84_sop_0_0_0_1_6_4_axb_7),.CI(un84_sop_0_0_0_1_6_4_cry_6),.O(un84_sop_0_0_0_1_6_4[7:7]));
  MUXCY_L un84_sop_0_0_0_1_6_4_cry_7_cZ(.DI(un84_sop_0_0_0_1_6_8[7:7]),.CI(un84_sop_0_0_0_1_6_4_cry_6),.S(un84_sop_0_0_0_1_6_4_axb_7),.LO(un84_sop_0_0_0_1_6_4_cry_7));
  XORCY un84_sop_0_0_0_1_6_4_s_6(.LI(un84_sop_0_0_0_1_6_4_axb_6),.CI(un84_sop_0_0_0_1_6_4_cry_5),.O(un84_sop_0_0_0_1_6_4[6:6]));
  MUXCY_L un84_sop_0_0_0_1_6_4_cry_6_cZ(.DI(un84_sop_0_0_0_1_6_8[6:6]),.CI(un84_sop_0_0_0_1_6_4_cry_5),.S(un84_sop_0_0_0_1_6_4_axb_6),.LO(un84_sop_0_0_0_1_6_4_cry_6));
  XORCY un84_sop_0_0_0_1_6_4_s_5(.LI(un84_sop_0_0_0_1_6_4_axb_5),.CI(un84_sop_0_0_0_1_6_4_cry_4),.O(un84_sop_0_0_0_1_6_4[5:5]));
  MUXCY_L un84_sop_0_0_0_1_6_4_cry_5_cZ(.DI(un84_sop_0_0_0_1_6_8[5:5]),.CI(un84_sop_0_0_0_1_6_4_cry_4),.S(un84_sop_0_0_0_1_6_4_axb_5),.LO(un84_sop_0_0_0_1_6_4_cry_5));
  XORCY un84_sop_0_0_0_1_6_4_s_4(.LI(un84_sop_0_0_0_1_6_4_axb_4),.CI(un84_sop_0_0_0_1_6_4_cry_3),.O(un84_sop_0_0_0_1_6_4[4:4]));
  MUXCY_L un84_sop_0_0_0_1_6_4_cry_4_cZ(.DI(un84_sop_0_0_0_1_6_8[4:4]),.CI(un84_sop_0_0_0_1_6_4_cry_3),.S(un84_sop_0_0_0_1_6_4_axb_4),.LO(un84_sop_0_0_0_1_6_4_cry_4));
  XORCY un84_sop_0_0_0_1_6_4_s_3(.LI(un84_sop_0_0_0_1_6_4_axb_3),.CI(un84_sop_0_0_0_1_6_4_cry_2),.O(un84_sop_0_0_0_1_6_4[3:3]));
  MUXCY_L un84_sop_0_0_0_1_6_4_cry_3_cZ(.DI(un1_x_6_0[4:4]),.CI(un84_sop_0_0_0_1_6_4_cry_2),.S(un84_sop_0_0_0_1_6_4_axb_3),.LO(un84_sop_0_0_0_1_6_4_cry_3));
  XORCY un84_sop_0_0_0_1_6_4_s_2(.LI(un84_sop_0_0_0_1_6_4_axb_2),.CI(un84_sop_0_0_0_1_6_4_cry_1),.O(un84_sop_0_0_0_1_6_4[2:2]));
  MUXCY_L un84_sop_0_0_0_1_6_4_cry_2_cZ(.DI(un1_x_6_0[3:3]),.CI(un84_sop_0_0_0_1_6_4_cry_1),.S(un84_sop_0_0_0_1_6_4_axb_2),.LO(un84_sop_0_0_0_1_6_4_cry_2));
  XORCY un84_sop_0_0_0_1_6_4_s_1(.LI(un84_sop_0_0_0_1_6_4_axb_1),.CI(un84_sop_0_0_0_1_6_4_cry_0),.O(un84_sop_0_0_0_1_6_4[1:1]));
  MUXCY_L un84_sop_0_0_0_1_6_4_cry_1_cZ(.DI(un1_x_6_0[2:2]),.CI(un84_sop_0_0_0_1_6_4_cry_0),.S(un84_sop_0_0_0_1_6_4_axb_1),.LO(un84_sop_0_0_0_1_6_4_cry_1));
  MUXCY_L un84_sop_0_0_0_1_6_4_cry_0_cZ(.DI(un1_x_6_0[1:1]),.CI(GND),.S(un84_sop_0_0_0_1_6_4[0:0]),.LO(un84_sop_0_0_0_1_6_4_cry_0));
  XORCY un1_x_10_s_11(.LI(un1_x_10_axb_11),.CI(un1_x_10_cry_10),.O(un1_x_10_0_0[15:15]));
  XORCY un1_x_10_s_10(.LI(un1_x_10_axb_10),.CI(un1_x_10_cry_9),.O(un1_x_10_0_0[14:14]));
  MUXCY_L un1_x_10_cry_10_cZ(.DI(un1_x_10_4[10:10]),.CI(un1_x_10_cry_9),.S(un1_x_10_axb_10),.LO(un1_x_10_cry_10));
  XORCY un1_x_10_s_9(.LI(un1_x_10_axb_9),.CI(un1_x_10_cry_8),.O(un1_x_10_0_0[13:13]));
  MUXCY_L un1_x_10_cry_9_cZ(.DI(un1_x_10_4[9:9]),.CI(un1_x_10_cry_8),.S(un1_x_10_axb_9),.LO(un1_x_10_cry_9));
  XORCY un1_x_10_s_8(.LI(un1_x_10_axb_8),.CI(un1_x_10_cry_7),.O(un1_x_10_0_0[12:12]));
  MUXCY_L un1_x_10_cry_8_cZ(.DI(un1_x_10_4[8:8]),.CI(un1_x_10_cry_7),.S(un1_x_10_axb_8),.LO(un1_x_10_cry_8));
  XORCY un1_x_10_s_7(.LI(un1_x_10_axb_7),.CI(un1_x_10_cry_6),.O(un1_x_10_0_0[11:11]));
  MUXCY_L un1_x_10_cry_7_cZ(.DI(un1_x_10_4[7:7]),.CI(un1_x_10_cry_6),.S(un1_x_10_axb_7),.LO(un1_x_10_cry_7));
  XORCY un1_x_10_s_6(.LI(un1_x_10_axb_6),.CI(un1_x_10_cry_5),.O(un1_x_10_0_0[10:10]));
  MUXCY_L un1_x_10_cry_6_cZ(.DI(un1_x_10_4[6:6]),.CI(un1_x_10_cry_5),.S(un1_x_10_axb_6),.LO(un1_x_10_cry_6));
  XORCY un1_x_10_s_5(.LI(un1_x_10_axb_5),.CI(un1_x_10_cry_4),.O(un1_x_10_0_0[9:9]));
  MUXCY_L un1_x_10_cry_5_cZ(.DI(un1_x_10_4[5:5]),.CI(un1_x_10_cry_4),.S(un1_x_10_axb_5),.LO(un1_x_10_cry_5));
  XORCY un1_x_10_s_4(.LI(un1_x_10_axb_4),.CI(un1_x_10_cry_3),.O(un1_x_10_0_0[8:8]));
  MUXCY_L un1_x_10_cry_4_cZ(.DI(un1_x_10_4[4:4]),.CI(un1_x_10_cry_3),.S(un1_x_10_axb_4),.LO(un1_x_10_cry_4));
  MUXCY_L un1_x_10_cry_3_cZ(.DI(un1_x_10_4[3:3]),.CI(GND),.S(un1_x_10_axb_3),.LO(un1_x_10_cry_3));
  XORCY un84_sop_1_6_0_s_13(.LI(un84_sop_1_6_0_axb_13),.CI(un84_sop_1_6_0_cry_12),.O(un84_sop_1_6[14:14]));
  XORCY un84_sop_1_6_0_s_12(.LI(un84_sop_1_6_0_axb_12),.CI(un84_sop_1_6_0_cry_11),.O(un84_sop_1_6[12:12]));
  MUXCY_L un84_sop_1_6_0_cry_12_cZ(.DI(un84_sop_1_6_0_o5_11),.CI(un84_sop_1_6_0_cry_11),.S(un84_sop_1_6_0_axb_12),.LO(un84_sop_1_6_0_cry_12));
  XORCY un84_sop_1_6_0_s_11(.LI(un84_sop_1_6_0_axb_11),.CI(un84_sop_1_6_0_cry_10),.O(un84_sop_1_6[11:11]));
  MUXCY_L un84_sop_1_6_0_cry_11_cZ(.DI(un84_sop_1_6_0_o5_10),.CI(un84_sop_1_6_0_cry_10),.S(un84_sop_1_6_0_axb_11),.LO(un84_sop_1_6_0_cry_11));
  XORCY un84_sop_1_6_0_s_10(.LI(un84_sop_1_6_0_axb_10),.CI(un84_sop_1_6_0_cry_9),.O(un84_sop_1_6[10:10]));
  MUXCY_L un84_sop_1_6_0_cry_10_cZ(.DI(un84_sop_1_6_0_o5_9),.CI(un84_sop_1_6_0_cry_9),.S(un84_sop_1_6_0_axb_10),.LO(un84_sop_1_6_0_cry_10));
  XORCY un84_sop_1_6_0_s_9(.LI(un84_sop_1_6_0_axb_9),.CI(un84_sop_1_6_0_cry_8),.O(un84_sop_1_6[9:9]));
  MUXCY_L un84_sop_1_6_0_cry_9_cZ(.DI(un84_sop_1_6_0_o5_8),.CI(un84_sop_1_6_0_cry_8),.S(un84_sop_1_6_0_axb_9),.LO(un84_sop_1_6_0_cry_9));
  XORCY un84_sop_1_6_0_s_8(.LI(un84_sop_1_6_0_axb_8),.CI(un84_sop_1_6_0_cry_7),.O(un84_sop_1_6[8:8]));
  MUXCY_L un84_sop_1_6_0_cry_8_cZ(.DI(un84_sop_1_6_0_o5_7),.CI(un84_sop_1_6_0_cry_7),.S(un84_sop_1_6_0_axb_8),.LO(un84_sop_1_6_0_cry_8));
  XORCY un84_sop_1_6_0_s_7(.LI(un84_sop_1_6_0_axb_7),.CI(un84_sop_1_6_0_cry_6),.O(un84_sop_1_6[7:7]));
  MUXCY_L un84_sop_1_6_0_cry_7_cZ(.DI(un84_sop_1_6_0_o5_6),.CI(un84_sop_1_6_0_cry_6),.S(un84_sop_1_6_0_axb_7),.LO(un84_sop_1_6_0_cry_7));
  XORCY un84_sop_1_6_0_s_6(.LI(un84_sop_1_6_0_axb_6),.CI(un84_sop_1_6_0_cry_5),.O(un84_sop_1_6[6:6]));
  MUXCY_L un84_sop_1_6_0_cry_6_cZ(.DI(un84_sop_1_6_0_o5_5),.CI(un84_sop_1_6_0_cry_5),.S(un84_sop_1_6_0_axb_6),.LO(un84_sop_1_6_0_cry_6));
  XORCY un84_sop_1_6_0_s_5(.LI(un84_sop_1_6_0_axb_5),.CI(un84_sop_1_6_0_cry_4),.O(un84_sop_1_6[5:5]));
  MUXCY_L un84_sop_1_6_0_cry_5_cZ(.DI(un84_sop_1_6_0_o5_4),.CI(un84_sop_1_6_0_cry_4),.S(un84_sop_1_6_0_axb_5),.LO(un84_sop_1_6_0_cry_5));
  XORCY un84_sop_1_6_0_s_4(.LI(un84_sop_1_6_0_axb_4),.CI(un84_sop_1_6_0_cry_3),.O(un84_sop_1_6[4:4]));
  MUXCY_L un84_sop_1_6_0_cry_4_cZ(.DI(un84_sop_1_6_0_o5_3),.CI(un84_sop_1_6_0_cry_3),.S(un84_sop_1_6_0_axb_4),.LO(un84_sop_1_6_0_cry_4));
  XORCY un84_sop_1_6_0_s_3(.LI(un84_sop_1_6_0_axb_3),.CI(un84_sop_1_6_0_cry_2),.O(un84_sop_1_6[3:3]));
  MUXCY_L un84_sop_1_6_0_cry_3_cZ(.DI(un84_sop_1_6_0_o5_2),.CI(un84_sop_1_6_0_cry_2),.S(un84_sop_1_6_0_axb_3),.LO(un84_sop_1_6_0_cry_3));
  XORCY un84_sop_1_6_0_s_2(.LI(un84_sop_1_6_0_axb_2),.CI(un84_sop_1_6_0_cry_1),.O(un84_sop_1_6[2:2]));
  MUXCY_L un84_sop_1_6_0_cry_2_cZ(.DI(un84_sop_1_6_0_axb_1_lut6_2_O5),.CI(un84_sop_1_6_0_cry_1),.S(un84_sop_1_6_0_axb_2),.LO(un84_sop_1_6_0_cry_2));
  XORCY un84_sop_1_6_0_s_1(.LI(un84_sop_1_6_0_axb_1),.CI(un84_sop_1_6_0_cry_0),.O(un84_sop_1_6[1:1]));
  MUXCY_L un84_sop_1_6_0_cry_1_cZ(.DI(GND),.CI(un84_sop_1_6_0_cry_0),.S(un84_sop_1_6_0_axb_1),.LO(un84_sop_1_6_0_cry_1));
  MUXCY_L un84_sop_1_6_0_cry_0_cZ(.DI(un1_x_2[5:5]),.CI(un84_sop_1_6_0_cry_0_cy),.S(un84_sop_1_6_0_axb_0_0),.LO(un84_sop_1_6_0_cry_0));
  XORCY un84_sop_0_0_0_1_6_8_s_11(.LI(un84_sop_0_0_0_1_6_8_axb_11),.CI(un84_sop_0_0_0_1_6_8_cry_10),.O(un84_sop_0_0_0_1_6_8[14:14]));
  XORCY un84_sop_0_0_0_1_6_8_s_10(.LI(un84_sop_0_0_0_1_6_8_axb_10),.CI(un84_sop_0_0_0_1_6_8_cry_9),.O(un84_sop_0_0_0_1_6_8[13:13]));
  MUXCY_L un84_sop_0_0_0_1_6_8_cry_10_cZ(.DI(un84_sop_0_0_0_10_0[13:13]),.CI(un84_sop_0_0_0_1_6_8_cry_9),.S(un84_sop_0_0_0_1_6_8_axb_10),.LO(un84_sop_0_0_0_1_6_8_cry_10));
  XORCY un84_sop_0_0_0_1_6_8_s_9(.LI(un84_sop_0_0_0_1_6_8_axb_9),.CI(un84_sop_0_0_0_1_6_8_cry_8),.O(un84_sop_0_0_0_1_6_8[12:12]));
  MUXCY_L un84_sop_0_0_0_1_6_8_cry_9_cZ(.DI(un84_sop_0_0_0_10_0[12:12]),.CI(un84_sop_0_0_0_1_6_8_cry_8),.S(un84_sop_0_0_0_1_6_8_axb_9),.LO(un84_sop_0_0_0_1_6_8_cry_9));
  XORCY un84_sop_0_0_0_1_6_8_s_8(.LI(un84_sop_0_0_0_1_6_8_axb_8),.CI(un84_sop_0_0_0_1_6_8_cry_7),.O(un84_sop_0_0_0_1_6_8[11:11]));
  MUXCY_L un84_sop_0_0_0_1_6_8_cry_8_cZ(.DI(un84_sop_0_0_0_1_6_8_o5_7),.CI(un84_sop_0_0_0_1_6_8_cry_7),.S(un84_sop_0_0_0_1_6_8_axb_8),.LO(un84_sop_0_0_0_1_6_8_cry_8));
  XORCY un84_sop_0_0_0_1_6_8_s_7(.LI(un84_sop_0_0_0_1_6_8_axb_7),.CI(un84_sop_0_0_0_1_6_8_cry_6),.O(un84_sop_0_0_0_1_6_8[10:10]));
  MUXCY_L un84_sop_0_0_0_1_6_8_cry_7_cZ(.DI(un84_sop_0_0_0_1_6_8_o5_6),.CI(un84_sop_0_0_0_1_6_8_cry_6),.S(un84_sop_0_0_0_1_6_8_axb_7),.LO(un84_sop_0_0_0_1_6_8_cry_7));
  XORCY un84_sop_0_0_0_1_6_8_s_6(.LI(un84_sop_0_0_0_1_6_8_axb_6),.CI(un84_sop_0_0_0_1_6_8_cry_5),.O(un84_sop_0_0_0_1_6_8[9:9]));
  MUXCY_L un84_sop_0_0_0_1_6_8_cry_6_cZ(.DI(un84_sop_0_0_0_1_6_8_o5_5),.CI(un84_sop_0_0_0_1_6_8_cry_5),.S(un84_sop_0_0_0_1_6_8_axb_6),.LO(un84_sop_0_0_0_1_6_8_cry_6));
  XORCY un84_sop_0_0_0_1_6_8_s_5(.LI(un84_sop_0_0_0_1_6_8_axb_5),.CI(un84_sop_0_0_0_1_6_8_cry_4),.O(un84_sop_0_0_0_1_6_8[8:8]));
  MUXCY_L un84_sop_0_0_0_1_6_8_cry_5_cZ(.DI(un84_sop_0_0_0_1_6_8_o5_4),.CI(un84_sop_0_0_0_1_6_8_cry_4),.S(un84_sop_0_0_0_1_6_8_axb_5),.LO(un84_sop_0_0_0_1_6_8_cry_5));
  XORCY un84_sop_0_0_0_1_6_8_s_4(.LI(un84_sop_0_0_0_1_6_8_axb_4),.CI(un84_sop_0_0_0_1_6_8_cry_3),.O(un84_sop_0_0_0_1_6_8[7:7]));
  MUXCY_L un84_sop_0_0_0_1_6_8_cry_4_cZ(.DI(un84_sop_0_0_0_1_6_8_o5_3),.CI(un84_sop_0_0_0_1_6_8_cry_3),.S(un84_sop_0_0_0_1_6_8_axb_4),.LO(un84_sop_0_0_0_1_6_8_cry_4));
  XORCY un84_sop_0_0_0_1_6_8_s_3(.LI(un84_sop_0_0_0_1_6_8_axb_3),.CI(un84_sop_0_0_0_1_6_8_cry_2),.O(un84_sop_0_0_0_1_6_8[6:6]));
  MUXCY_L un84_sop_0_0_0_1_6_8_cry_3_cZ(.DI(un84_sop_0_0_0_1_6_8_axb_2_lut6_2_O5),.CI(un84_sop_0_0_0_1_6_8_cry_2),.S(un84_sop_0_0_0_1_6_8_axb_3),.LO(un84_sop_0_0_0_1_6_8_cry_3));
  XORCY un84_sop_0_0_0_1_6_8_s_2(.LI(un84_sop_0_0_0_1_6_8_axb_2),.CI(un84_sop_0_0_0_1_6_8_cry_1),.O(un84_sop_0_0_0_1_6_8[5:5]));
  MUXCY_L un84_sop_0_0_0_1_6_8_cry_2_cZ(.DI(GND),.CI(un84_sop_0_0_0_1_6_8_cry_1),.S(un84_sop_0_0_0_1_6_8_axb_2),.LO(un84_sop_0_0_0_1_6_8_cry_2));
  XORCY un84_sop_0_0_0_1_6_8_s_1(.LI(un84_sop_0_0_0_1_6_8_axb_1),.CI(un84_sop_0_0_0_1_6_8_cry_0),.O(un84_sop_0_0_0_1_6_8[4:4]));
  MUXCY_L un84_sop_0_0_0_1_6_8_cry_1_cZ(.DI(un84_sop_0_0_0_10_0[4:4]),.CI(un84_sop_0_0_0_1_6_8_cry_0),.S(un84_sop_0_0_0_1_6_8_axb_1),.LO(un84_sop_0_0_0_1_6_8_cry_1));
  MUXCY_L un84_sop_0_0_0_1_6_8_cry_0_cZ(.DI(un84_sop_0_0_0_10_0[3:3]),.CI(GND),.S(un84_sop_0_0_0_1_6_8[3:3]),.LO(un84_sop_0_0_0_1_6_8_cry_0));
  XORCY un84_sop_0_0_0_6_6_0_s_14(.LI(un84_sop_0_0_0_6_6_0_axb_14),.CI(un84_sop_0_0_0_6_6_0_cry_13),.O(un84_sop_0_0_0_1_6_6[14:14]));
  XORCY un84_sop_0_0_0_6_6_0_s_13(.LI(un84_sop_0_0_0_6_6_0_axb_13),.CI(un84_sop_0_0_0_6_6_0_cry_12),.O(un84_sop_0_0_0_1_6_6[13:13]));
  MUXCY_L un84_sop_0_0_0_6_6_0_cry_13_cZ(.DI(un84_sop_0_0_0_6_6_0_o5_12),.CI(un84_sop_0_0_0_6_6_0_cry_12),.S(un84_sop_0_0_0_6_6_0_axb_13),.LO(un84_sop_0_0_0_6_6_0_cry_13));
  XORCY un84_sop_0_0_0_6_6_0_s_12(.LI(un84_sop_0_0_0_6_6_0_axb_12),.CI(un84_sop_0_0_0_6_6_0_cry_11),.O(un84_sop_0_0_0_1_6_6[12:12]));
  MUXCY_L un84_sop_0_0_0_6_6_0_cry_12_cZ(.DI(un84_sop_0_0_0_6_6_0_o5_11),.CI(un84_sop_0_0_0_6_6_0_cry_11),.S(un84_sop_0_0_0_6_6_0_axb_12),.LO(un84_sop_0_0_0_6_6_0_cry_12));
  XORCY un84_sop_0_0_0_6_6_0_s_11(.LI(un84_sop_0_0_0_6_6_0_axb_11),.CI(un84_sop_0_0_0_6_6_0_cry_10),.O(un84_sop_0_0_0_1_6_6[11:11]));
  MUXCY_L un84_sop_0_0_0_6_6_0_cry_11_cZ(.DI(un84_sop_0_0_0_6_6_0_o5_10),.CI(un84_sop_0_0_0_6_6_0_cry_10),.S(un84_sop_0_0_0_6_6_0_axb_11),.LO(un84_sop_0_0_0_6_6_0_cry_11));
  XORCY un84_sop_0_0_0_6_6_0_s_10(.LI(un84_sop_0_0_0_6_6_0_axb_10),.CI(un84_sop_0_0_0_6_6_0_cry_9),.O(un84_sop_0_0_0_1_6_6[10:10]));
  MUXCY_L un84_sop_0_0_0_6_6_0_cry_10_cZ(.DI(un84_sop_0_0_0_6_6_0_o5_9),.CI(un84_sop_0_0_0_6_6_0_cry_9),.S(un84_sop_0_0_0_6_6_0_axb_10),.LO(un84_sop_0_0_0_6_6_0_cry_10));
  XORCY un84_sop_0_0_0_6_6_0_s_9(.LI(un84_sop_0_0_0_6_6_0_axb_9),.CI(un84_sop_0_0_0_6_6_0_cry_8),.O(un84_sop_0_0_0_1_6_6[9:9]));
  MUXCY_L un84_sop_0_0_0_6_6_0_cry_9_cZ(.DI(un84_sop_0_0_0_6_6_0_o5_8),.CI(un84_sop_0_0_0_6_6_0_cry_8),.S(un84_sop_0_0_0_6_6_0_axb_9),.LO(un84_sop_0_0_0_6_6_0_cry_9));
  XORCY un84_sop_0_0_0_6_6_0_s_8(.LI(un84_sop_0_0_0_6_6_0_axb_8),.CI(un84_sop_0_0_0_6_6_0_cry_7),.O(un84_sop_0_0_0_1_6_6[8:8]));
  MUXCY_L un84_sop_0_0_0_6_6_0_cry_8_cZ(.DI(un84_sop_0_0_0_6_6_0_o5_7),.CI(un84_sop_0_0_0_6_6_0_cry_7),.S(un84_sop_0_0_0_6_6_0_axb_8),.LO(un84_sop_0_0_0_6_6_0_cry_8));
  XORCY un84_sop_0_0_0_6_6_0_s_7(.LI(un84_sop_0_0_0_6_6_0_axb_7),.CI(un84_sop_0_0_0_6_6_0_cry_6),.O(un84_sop_0_0_0_1_6_6[7:7]));
  MUXCY_L un84_sop_0_0_0_6_6_0_cry_7_cZ(.DI(un84_sop_0_0_0_6_6_0_o5_6),.CI(un84_sop_0_0_0_6_6_0_cry_6),.S(un84_sop_0_0_0_6_6_0_axb_7),.LO(un84_sop_0_0_0_6_6_0_cry_7));
  XORCY un84_sop_0_0_0_6_6_0_s_6(.LI(un84_sop_0_0_0_6_6_0_axb_6),.CI(un84_sop_0_0_0_6_6_0_cry_5),.O(un84_sop_0_0_0_1_6_6[6:6]));
  MUXCY_L un84_sop_0_0_0_6_6_0_cry_6_cZ(.DI(un84_sop_0_0_0_6_6_0_o5_5),.CI(un84_sop_0_0_0_6_6_0_cry_5),.S(un84_sop_0_0_0_6_6_0_axb_6),.LO(un84_sop_0_0_0_6_6_0_cry_6));
  XORCY un84_sop_0_0_0_6_6_0_s_5(.LI(un84_sop_0_0_0_6_6_0_axb_5),.CI(un84_sop_0_0_0_6_6_0_cry_4),.O(un84_sop_0_0_0_1_6_6[5:5]));
  MUXCY_L un84_sop_0_0_0_6_6_0_cry_5_cZ(.DI(un84_sop_0_0_0_6_6_0_o5_4),.CI(un84_sop_0_0_0_6_6_0_cry_4),.S(un84_sop_0_0_0_6_6_0_axb_5),.LO(un84_sop_0_0_0_6_6_0_cry_5));
  XORCY un84_sop_0_0_0_6_6_0_s_4(.LI(un84_sop_0_0_0_6_6_0_axb_4),.CI(un84_sop_0_0_0_6_6_0_cry_3),.O(un84_sop_0_0_0_1_6_6[4:4]));
  MUXCY_L un84_sop_0_0_0_6_6_0_cry_4_cZ(.DI(un84_sop_0_0_0_6_6_0_o5_3),.CI(un84_sop_0_0_0_6_6_0_cry_3),.S(un84_sop_0_0_0_6_6_0_axb_4),.LO(un84_sop_0_0_0_6_6_0_cry_4));
  XORCY un84_sop_0_0_0_6_6_0_s_3(.LI(un84_sop_0_0_0_6_6_0_axb_3),.CI(un84_sop_0_0_0_6_6_0_cry_2),.O(un84_sop_0_0_0_1_6_6[3:3]));
  MUXCY_L un84_sop_0_0_0_6_6_0_cry_3_cZ(.DI(un84_sop_0_0_0_6_6_0_o5_2),.CI(un84_sop_0_0_0_6_6_0_cry_2),.S(un84_sop_0_0_0_6_6_0_axb_3),.LO(un84_sop_0_0_0_6_6_0_cry_3));
  XORCY un84_sop_0_0_0_6_6_0_s_2(.LI(un84_sop_0_0_0_6_6_0_axb_2),.CI(un84_sop_0_0_0_6_6_0_cry_1),.O(un84_sop_0_0_0_1_6_6[2:2]));
  MUXCY_L un84_sop_0_0_0_6_6_0_cry_2_cZ(.DI(un84_sop_0_0_0_6_6_0_axb_1_lut6_2_O5),.CI(un84_sop_0_0_0_6_6_0_cry_1),.S(un84_sop_0_0_0_6_6_0_axb_2),.LO(un84_sop_0_0_0_6_6_0_cry_2));
  XORCY un84_sop_0_0_0_6_6_0_s_1(.LI(un84_sop_0_0_0_6_6_0_axb_1),.CI(un84_sop_0_0_0_6_6_0_cry_0),.O(un84_sop_0_0_0_1_6_6[1:1]));
  MUXCY_L un84_sop_0_0_0_6_6_0_cry_1_cZ(.DI(GND),.CI(un84_sop_0_0_0_6_6_0_cry_0),.S(un84_sop_0_0_0_6_6_0_axb_1),.LO(un84_sop_0_0_0_6_6_0_cry_1));
  MUXCY_L un84_sop_0_0_0_6_6_0_cry_0_cZ(.DI(un1_x_8_0[4:4]),.CI(un84_sop_0_0_0_6_6_0_cry_0_cy),.S(un84_sop_0_0_0_6_0_axb_0_1),.LO(un84_sop_0_0_0_6_6_0_cry_0));
  XORCY un84_sop_0_0_0_11_0_s_14(.LI(un84_sop_0_0_0_11_0_axb_14),.CI(un84_sop_0_0_0_11_0_cry_13),.O(un84_sop_0_0_0_0_8[14:14]));
  XORCY un84_sop_0_0_0_11_0_s_13(.LI(un84_sop_0_0_0_11_0_axb_13),.CI(un84_sop_0_0_0_11_0_cry_12),.O(un84_sop_0_0_0_0_8[13:13]));
  MUXCY_L un84_sop_0_0_0_11_0_cry_13_cZ(.DI(un84_sop_0_0_0_11_0_o5_12),.CI(un84_sop_0_0_0_11_0_cry_12),.S(un84_sop_0_0_0_11_0_axb_13),.LO(un84_sop_0_0_0_11_0_cry_13));
  XORCY un84_sop_0_0_0_11_0_s_12(.LI(un84_sop_0_0_0_11_0_axb_12),.CI(un84_sop_0_0_0_11_0_cry_11),.O(un84_sop_0_0_0_0_8[12:12]));
  MUXCY_L un84_sop_0_0_0_11_0_cry_12_cZ(.DI(un84_sop_0_0_0_11_0_o5_11),.CI(un84_sop_0_0_0_11_0_cry_11),.S(un84_sop_0_0_0_11_0_axb_12),.LO(un84_sop_0_0_0_11_0_cry_12));
  XORCY un84_sop_0_0_0_11_0_s_11(.LI(un84_sop_0_0_0_11_0_axb_11),.CI(un84_sop_0_0_0_11_0_cry_10),.O(un84_sop_0_0_0_0_8[11:11]));
  MUXCY_L un84_sop_0_0_0_11_0_cry_11_cZ(.DI(un84_sop_0_0_0_11_0_o5_10),.CI(un84_sop_0_0_0_11_0_cry_10),.S(un84_sop_0_0_0_11_0_axb_11),.LO(un84_sop_0_0_0_11_0_cry_11));
  XORCY un84_sop_0_0_0_11_0_s_10(.LI(un84_sop_0_0_0_11_0_axb_10),.CI(un84_sop_0_0_0_11_0_cry_9),.O(un84_sop_0_0_0_0_8[10:10]));
  MUXCY_L un84_sop_0_0_0_11_0_cry_10_cZ(.DI(un84_sop_0_0_0_11_0_o5_9),.CI(un84_sop_0_0_0_11_0_cry_9),.S(un84_sop_0_0_0_11_0_axb_10),.LO(un84_sop_0_0_0_11_0_cry_10));
  XORCY un84_sop_0_0_0_11_0_s_9(.LI(un84_sop_0_0_0_11_0_axb_9),.CI(un84_sop_0_0_0_11_0_cry_8),.O(un84_sop_0_0_0_0_8[9:9]));
  MUXCY_L un84_sop_0_0_0_11_0_cry_9_cZ(.DI(un84_sop_0_0_0_11_0_o5_8),.CI(un84_sop_0_0_0_11_0_cry_8),.S(un84_sop_0_0_0_11_0_axb_9),.LO(un84_sop_0_0_0_11_0_cry_9));
  XORCY un84_sop_0_0_0_11_0_s_8(.LI(un84_sop_0_0_0_11_0_axb_8),.CI(un84_sop_0_0_0_11_0_cry_7),.O(un84_sop_0_0_0_0_8[8:8]));
  MUXCY_L un84_sop_0_0_0_11_0_cry_8_cZ(.DI(un84_sop_0_0_0_11_0_o5_7),.CI(un84_sop_0_0_0_11_0_cry_7),.S(un84_sop_0_0_0_11_0_axb_8),.LO(un84_sop_0_0_0_11_0_cry_8));
  XORCY un84_sop_0_0_0_11_0_s_7(.LI(un84_sop_0_0_0_11_0_axb_7),.CI(un84_sop_0_0_0_11_0_cry_6),.O(un84_sop_0_0_0_0_8[7:7]));
  MUXCY_L un84_sop_0_0_0_11_0_cry_7_cZ(.DI(un84_sop_0_0_0_11_0_o5_6),.CI(un84_sop_0_0_0_11_0_cry_6),.S(un84_sop_0_0_0_11_0_axb_7),.LO(un84_sop_0_0_0_11_0_cry_7));
  XORCY un84_sop_0_0_0_11_0_s_6(.LI(un84_sop_0_0_0_11_0_axb_6),.CI(un84_sop_0_0_0_11_0_cry_5),.O(un84_sop_0_0_0_0_8[6:6]));
  MUXCY_L un84_sop_0_0_0_11_0_cry_6_cZ(.DI(un84_sop_0_0_0_11_0_o5_5),.CI(un84_sop_0_0_0_11_0_cry_5),.S(un84_sop_0_0_0_11_0_axb_6),.LO(un84_sop_0_0_0_11_0_cry_6));
  XORCY un84_sop_0_0_0_11_0_s_5(.LI(un84_sop_0_0_0_11_0_axb_5),.CI(un84_sop_0_0_0_11_0_cry_4),.O(un84_sop_0_0_0_0_8[5:5]));
  MUXCY_L un84_sop_0_0_0_11_0_cry_5_cZ(.DI(un84_sop_0_0_0_11_0_o5_4),.CI(un84_sop_0_0_0_11_0_cry_4),.S(un84_sop_0_0_0_11_0_axb_5),.LO(un84_sop_0_0_0_11_0_cry_5));
  XORCY un84_sop_0_0_0_11_0_s_4(.LI(un84_sop_0_0_0_11_0_axb_4),.CI(un84_sop_0_0_0_11_0_cry_3),.O(un84_sop_0_0_0_0_8[4:4]));
  MUXCY_L un84_sop_0_0_0_11_0_cry_4_cZ(.DI(un84_sop_0_0_0_11_0_o5_3),.CI(un84_sop_0_0_0_11_0_cry_3),.S(un84_sop_0_0_0_11_0_axb_4),.LO(un84_sop_0_0_0_11_0_cry_4));
  XORCY un84_sop_0_0_0_11_0_s_3(.LI(un84_sop_0_0_0_11_0_axb_3),.CI(un84_sop_0_0_0_11_0_cry_2),.O(un84_sop_0_0_0_0_8[3:3]));
  MUXCY_L un84_sop_0_0_0_11_0_cry_3_cZ(.DI(un84_sop_0_0_0_11_0_o5_2),.CI(un84_sop_0_0_0_11_0_cry_2),.S(un84_sop_0_0_0_11_0_axb_3),.LO(un84_sop_0_0_0_11_0_cry_3));
  XORCY un84_sop_0_0_0_11_0_s_2(.LI(un84_sop_0_0_0_11_0_axb_2),.CI(un84_sop_0_0_0_11_0_cry_1),.O(un84_sop_0_0_0_0_8[2:2]));
  MUXCY_L un84_sop_0_0_0_11_0_cry_2_cZ(.DI(un84_sop_0_0_0_11_0_cry_2_RNO),.CI(un84_sop_0_0_0_11_0_cry_1),.S(un84_sop_0_0_0_11_0_axb_2),.LO(un84_sop_0_0_0_11_0_cry_2));
  XORCY un84_sop_0_0_0_11_0_s_1(.LI(un84_sop_0_0_0_11_0_axb_1),.CI(un84_sop_0_0_0_11_0_cry_0),.O(un84_sop_0_0_0_0_8[1:1]));
  MUXCY_L un84_sop_0_0_0_11_0_cry_1_cZ(.DI(un84_sop_0_0_0_0_11_6[1:1]),.CI(un84_sop_0_0_0_11_0_cry_0),.S(un84_sop_0_0_0_11_0_axb_1),.LO(un84_sop_0_0_0_11_0_cry_1));
  XORCY un84_sop_0_0_0_11_0_s_0(.LI(un84_sop_0_0_0_11_0_axb_0),.CI(un84_sop_0_0_0_11_0_cry_0_cy),.O(un84_sop_0_0_0_0_8[0:0]));
  MUXCY_L un84_sop_0_0_0_11_0_cry_0_cZ(.DI(un84_sop_0_0_0_0_11_6[0:0]),.CI(un84_sop_0_0_0_11_0_cry_0_cy),.S(un84_sop_0_0_0_11_0_axb_0),.LO(un84_sop_0_0_0_11_0_cry_0));
  XORCY un84_sop_0_0_0_11_6_0_s_13(.LI(un84_sop_0_0_0_11_6_0_axb_13),.CI(un84_sop_0_0_0_11_6_0_cry_12),.O(un84_sop_0_0_0_0_11_6[14:14]));
  XORCY un84_sop_0_0_0_11_6_0_s_12(.LI(un84_sop_0_0_0_11_6_0_axb_12),.CI(un84_sop_0_0_0_11_6_0_cry_11),.O(un84_sop_0_0_0_0_11_6[12:12]));
  MUXCY_L un84_sop_0_0_0_11_6_0_cry_12_cZ(.DI(un84_sop_0_0_0_11_6_0_o5_11),.CI(un84_sop_0_0_0_11_6_0_cry_11),.S(un84_sop_0_0_0_11_6_0_axb_12),.LO(un84_sop_0_0_0_11_6_0_cry_12));
  XORCY un84_sop_0_0_0_11_6_0_s_11(.LI(un84_sop_0_0_0_11_6_0_axb_11),.CI(un84_sop_0_0_0_11_6_0_cry_10),.O(un84_sop_0_0_0_0_11_6[11:11]));
  MUXCY_L un84_sop_0_0_0_11_6_0_cry_11_cZ(.DI(un84_sop_0_0_0_11_6_0_o5_10),.CI(un84_sop_0_0_0_11_6_0_cry_10),.S(un84_sop_0_0_0_11_6_0_axb_11),.LO(un84_sop_0_0_0_11_6_0_cry_11));
  XORCY un84_sop_0_0_0_11_6_0_s_10(.LI(un84_sop_0_0_0_11_6_0_axb_10),.CI(un84_sop_0_0_0_11_6_0_cry_9),.O(un84_sop_0_0_0_0_11_6[10:10]));
  MUXCY_L un84_sop_0_0_0_11_6_0_cry_10_cZ(.DI(un84_sop_0_0_0_11_6_0_o5_9),.CI(un84_sop_0_0_0_11_6_0_cry_9),.S(un84_sop_0_0_0_11_6_0_axb_10),.LO(un84_sop_0_0_0_11_6_0_cry_10));
  XORCY un84_sop_0_0_0_11_6_0_s_9(.LI(un84_sop_0_0_0_11_6_0_axb_9),.CI(un84_sop_0_0_0_11_6_0_cry_8),.O(un84_sop_0_0_0_0_11_6[9:9]));
  MUXCY_L un84_sop_0_0_0_11_6_0_cry_9_cZ(.DI(un84_sop_0_0_0_11_6_0_o5_8),.CI(un84_sop_0_0_0_11_6_0_cry_8),.S(un84_sop_0_0_0_11_6_0_axb_9),.LO(un84_sop_0_0_0_11_6_0_cry_9));
  XORCY un84_sop_0_0_0_11_6_0_s_8(.LI(un84_sop_0_0_0_11_6_0_axb_8),.CI(un84_sop_0_0_0_11_6_0_cry_7),.O(un84_sop_0_0_0_0_11_6[8:8]));
  MUXCY_L un84_sop_0_0_0_11_6_0_cry_8_cZ(.DI(un84_sop_0_0_0_11_6_0_o5_7),.CI(un84_sop_0_0_0_11_6_0_cry_7),.S(un84_sop_0_0_0_11_6_0_axb_8),.LO(un84_sop_0_0_0_11_6_0_cry_8));
  XORCY un84_sop_0_0_0_11_6_0_s_7(.LI(un84_sop_0_0_0_11_6_0_axb_7),.CI(un84_sop_0_0_0_11_6_0_cry_6),.O(un84_sop_0_0_0_0_11_6[7:7]));
  MUXCY_L un84_sop_0_0_0_11_6_0_cry_7_cZ(.DI(un84_sop_0_0_0_11_6_0_o5_6),.CI(un84_sop_0_0_0_11_6_0_cry_6),.S(un84_sop_0_0_0_11_6_0_axb_7),.LO(un84_sop_0_0_0_11_6_0_cry_7));
  XORCY un84_sop_0_0_0_11_6_0_s_6(.LI(un84_sop_0_0_0_11_6_0_axb_6),.CI(un84_sop_0_0_0_11_6_0_cry_5),.O(un84_sop_0_0_0_0_11_6[6:6]));
  MUXCY_L un84_sop_0_0_0_11_6_0_cry_6_cZ(.DI(un84_sop_0_0_0_11_6_0_o5_5),.CI(un84_sop_0_0_0_11_6_0_cry_5),.S(un84_sop_0_0_0_11_6_0_axb_6),.LO(un84_sop_0_0_0_11_6_0_cry_6));
  XORCY un84_sop_0_0_0_11_6_0_s_5(.LI(un84_sop_0_0_0_11_6_0_axb_5),.CI(un84_sop_0_0_0_11_6_0_cry_4),.O(un84_sop_0_0_0_0_11_6[5:5]));
  MUXCY_L un84_sop_0_0_0_11_6_0_cry_5_cZ(.DI(un84_sop_0_0_0_11_6_0_o5_4),.CI(un84_sop_0_0_0_11_6_0_cry_4),.S(un84_sop_0_0_0_11_6_0_axb_5),.LO(un84_sop_0_0_0_11_6_0_cry_5));
  XORCY un84_sop_0_0_0_11_6_0_s_4(.LI(un84_sop_0_0_0_11_6_0_axb_4),.CI(un84_sop_0_0_0_11_6_0_cry_3),.O(un84_sop_0_0_0_0_11_6[4:4]));
  MUXCY_L un84_sop_0_0_0_11_6_0_cry_4_cZ(.DI(un84_sop_0_0_0_11_6_0_o5_3),.CI(un84_sop_0_0_0_11_6_0_cry_3),.S(un84_sop_0_0_0_11_6_0_axb_4),.LO(un84_sop_0_0_0_11_6_0_cry_4));
  XORCY un84_sop_0_0_0_11_6_0_s_3(.LI(un84_sop_0_0_0_11_6_0_axb_3),.CI(un84_sop_0_0_0_11_6_0_cry_2),.O(un84_sop_0_0_0_0_11_6[3:3]));
  MUXCY_L un84_sop_0_0_0_11_6_0_cry_3_cZ(.DI(un84_sop_0_0_0_11_6_0_o5_2),.CI(un84_sop_0_0_0_11_6_0_cry_2),.S(un84_sop_0_0_0_11_6_0_axb_3),.LO(un84_sop_0_0_0_11_6_0_cry_3));
  XORCY un84_sop_0_0_0_11_6_0_s_2(.LI(un84_sop_0_0_0_11_6_0_axb_2),.CI(un84_sop_0_0_0_11_6_0_cry_1),.O(un84_sop_0_0_0_0_11_6[2:2]));
  MUXCY_L un84_sop_0_0_0_11_6_0_cry_2_cZ(.DI(un84_sop_0_0_0_11_6_0_axb_1_lut6_2_O5),.CI(un84_sop_0_0_0_11_6_0_cry_1),.S(un84_sop_0_0_0_11_6_0_axb_2),.LO(un84_sop_0_0_0_11_6_0_cry_2));
  XORCY un84_sop_0_0_0_11_6_0_s_1(.LI(un84_sop_0_0_0_11_6_0_axb_1),.CI(un84_sop_0_0_0_11_6_0_cry_0),.O(un84_sop_0_0_0_0_11_6[1:1]));
  MUXCY_L un84_sop_0_0_0_11_6_0_cry_1_cZ(.DI(GND),.CI(un84_sop_0_0_0_11_6_0_cry_0),.S(un84_sop_0_0_0_11_6_0_axb_1),.LO(un84_sop_0_0_0_11_6_0_cry_1));
  MUXCY_L un84_sop_0_0_0_11_6_0_cry_0_cZ(.DI(un1_x_13_0_0[5:5]),.CI(un84_sop_0_0_0_11_6_0_cry_0_cy),.S(un84_sop_0_0_0_6_0_axb_0_0),.LO(un84_sop_0_0_0_11_6_0_cry_0));
  DSP48E1 desc57(.ACOUT(ACOUT[29:0]),.BCOUT({x_0_10[7:7],x_0_9[7:7],x_0_8[7:7],x_0_7[7:7],x_0_6[7:7],x_0_5[7:7],x_0_4[7:7],x_0_3[7:7],x_0_2[7:7],x_0_1[7:7],x_0_0[7:0]}),.CARRYCASCOUT(CARRYCASCOUT),.CARRYOUT(CARRYOUT[3:0]),.MULTSIGNOUT(MULTSIGNOUT),.OVERFLOW(OVERFLOW),.P({P_uc[47:12],un1_x_1[15:4]}),.PATTERNBDETECT(PATTERNBDETECT),.PATTERNDETECT(PATTERNDETECT),.PCOUT(PCOUT[47:0]),.UNDERFLOW(UNDERFLOW),.A({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,GND,VCC,VCC}),.ACIN({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.ALUMODE({GND,GND,GND,GND}),.B({x_in[7:7],x_in[7:7],x_in[7:7],x_in[7:7],x_in[7:7],x_in[7:7],x_in[7:7],x_in[7:7],x_in[7:7],x_in[7:7],x_in[7:0]}),.BCIN({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.C({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.CARRYCASCIN(GND),.CARRYIN(GND),.CARRYINSEL({GND,GND,GND}),.CEA1(GND),.CEA2(GND),.CEAD(GND),.CEALUMODE(GND),.CEB1(GND),.CEB2(VCC),.CEC(GND),.CECARRYIN(GND),.CECTRL(GND),.CED(GND),.CEINMODE(GND),.CEM(GND),.CEP(VCC),.CLK(clk),.D({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND}),.INMODE({GND,GND,GND,GND,GND}),.MULTSIGNIN(GND),.OPMODE({GND,GND,GND,GND,VCC,GND,VCC}),.PCIN({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND}),.RSTA(GND),.RSTALLCARRYIN(GND),.RSTALUMODE(GND),.RSTB(GND),.RSTC(GND),.RSTCTRL(GND),.RSTD(GND),.RSTINMODE(GND),.RSTM(GND),.RSTP(GND));
defparam desc57.ACASCREG=0;
defparam desc57.ADREG=0;
defparam desc57.ALUMODEREG=0;
defparam desc57.AREG=0;
defparam desc57.AUTORESET_PATDET="NO_RESET";
defparam desc57.A_INPUT="DIRECT";
defparam desc57.BCASCREG=1;
defparam desc57.BREG=1;
defparam desc57.B_INPUT="DIRECT";
defparam desc57.CARRYINREG=0;
defparam desc57.CARRYINSELREG=0;
defparam desc57.CREG=1;
defparam desc57.DREG=0;
defparam desc57.INMODEREG=0;
defparam desc57.MREG=0;
defparam desc57.OPMODEREG=0;
defparam desc57.PREG=1;
defparam desc57.USE_DPORT="FALSE";
defparam desc57.USE_MULT="MULTIPLY";
defparam desc57.USE_SIMD="ONE48";
  DSP48E1 desc58(.ACOUT(ACOUT_0[29:0]),.BCOUT({x_9_10[7:7],x_9_9[7:7],x_9_8[7:7],x_9_7[7:7],x_9_6[7:7],x_9_5[7:7],x_9_4[7:7],x_9_3[7:7],x_9_2[7:7],x_9_1[7:7],x_9_0[7:0]}),.CARRYCASCOUT(CARRYCASCOUT_0),.CARRYOUT(CARRYOUT_0[3:0]),.MULTSIGNOUT(MULTSIGNOUT_0),.OVERFLOW(OVERFLOW_0),.P({P_uc_0[47:12],un1_x_12_0_0[15:4]}),.PATTERNBDETECT(PATTERNBDETECT_0),.PATTERNDETECT(PATTERNDETECT_0),.PCOUT(PCOUT_0[47:0]),.UNDERFLOW(UNDERFLOW_0),.A({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,VCC,VCC,VCC}),.ACIN({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.ALUMODE({GND,GND,GND,GND}),.B({x_7[7:7],x_7[7:7],x_7[7:7],x_7[7:7],x_7[7:7],x_7[7:7],x_7[7:7],x_7[7:7],x_7[7:7],x_7[7:7],x_7[7:0]}),.BCIN({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.C({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.CARRYCASCIN(GND),.CARRYIN(GND),.CARRYINSEL({GND,GND,GND}),.CEA1(VCC),.CEA2(VCC),.CEAD(GND),.CEALUMODE(GND),.CEB1(VCC),.CEB2(VCC),.CEC(GND),.CECARRYIN(GND),.CECTRL(GND),.CED(GND),.CEINMODE(GND),.CEM(GND),.CEP(VCC),.CLK(clk),.D({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND}),.INMODE({GND,GND,GND,GND,GND}),.MULTSIGNIN(GND),.OPMODE({GND,GND,GND,GND,VCC,GND,VCC}),.PCIN({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND}),.RSTA(GND),.RSTALLCARRYIN(GND),.RSTALUMODE(GND),.RSTB(GND),.RSTC(GND),.RSTCTRL(GND),.RSTD(GND),.RSTINMODE(GND),.RSTM(GND),.RSTP(GND));
defparam desc58.ACASCREG=2;
defparam desc58.ADREG=0;
defparam desc58.ALUMODEREG=0;
defparam desc58.AREG=2;
defparam desc58.AUTORESET_PATDET="NO_RESET";
defparam desc58.A_INPUT="DIRECT";
defparam desc58.BCASCREG=2;
defparam desc58.BREG=2;
defparam desc58.B_INPUT="DIRECT";
defparam desc58.CARRYINREG=0;
defparam desc58.CARRYINSELREG=0;
defparam desc58.CREG=1;
defparam desc58.DREG=0;
defparam desc58.INMODEREG=0;
defparam desc58.MREG=0;
defparam desc58.OPMODEREG=0;
defparam desc58.PREG=1;
defparam desc58.USE_DPORT="FALSE";
defparam desc58.USE_MULT="MULTIPLY";
defparam desc58.USE_SIMD="ONE48";
  DSP48E1 desc59(.ACOUT(ACOUT_1[29:0]),.BCOUT(BCOUT_1[17:0]),.CARRYCASCOUT(CARRYCASCOUT_1),.CARRYOUT(CARRYOUT_1[3:0]),.MULTSIGNOUT(MULTSIGNOUT_1),.OVERFLOW(OVERFLOW_1),.P({P_uc_1[47:12],un1_x_14_0_0[15:4]}),.PATTERNBDETECT(PATTERNBDETECT_1),.PATTERNDETECT(PATTERNDETECT_1),.PCOUT(PCOUT_1[47:0]),.UNDERFLOW(UNDERFLOW_1),.A({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,GND,VCC,VCC}),.ACIN({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.ALUMODE({GND,GND,GND,GND}),.B({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.BCIN({x_10_10[7:7],x_10_9[7:7],x_10_8[7:7],x_10_7[7:7],x_10_6[7:7],x_10_5[7:7],x_10_4[7:7],x_10_3[7:7],x_10_2[7:7],x_10_1[7:7],x_10_0[7:0]}),.C({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.CARRYCASCIN(GND),.CARRYIN(GND),.CARRYINSEL({GND,GND,GND}),.CEA1(GND),.CEA2(GND),.CEAD(GND),.CEALUMODE(GND),.CEB1(GND),.CEB2(VCC),.CEC(GND),.CECARRYIN(GND),.CECTRL(GND),.CED(GND),.CEINMODE(GND),.CEM(GND),.CEP(VCC),.CLK(clk),.D({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND}),.INMODE({GND,GND,GND,GND,GND}),.MULTSIGNIN(GND),.OPMODE({GND,GND,GND,GND,VCC,GND,VCC}),.PCIN({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND}),.RSTA(GND),.RSTALLCARRYIN(GND),.RSTALUMODE(GND),.RSTB(GND),.RSTC(GND),.RSTCTRL(GND),.RSTD(GND),.RSTINMODE(GND),.RSTM(GND),.RSTP(GND));
defparam desc59.ACASCREG=0;
defparam desc59.ADREG=0;
defparam desc59.ALUMODEREG=0;
defparam desc59.AREG=0;
defparam desc59.AUTORESET_PATDET="NO_RESET";
defparam desc59.A_INPUT="DIRECT";
defparam desc59.BCASCREG=1;
defparam desc59.BREG=1;
defparam desc59.B_INPUT="CASCADE";
defparam desc59.CARRYINREG=0;
defparam desc59.CARRYINSELREG=0;
defparam desc59.CREG=1;
defparam desc59.DREG=0;
defparam desc59.INMODEREG=0;
defparam desc59.MREG=0;
defparam desc59.OPMODEREG=0;
defparam desc59.PREG=1;
defparam desc59.USE_DPORT="FALSE";
defparam desc59.USE_MULT="MULTIPLY";
defparam desc59.USE_SIMD="ONE48";
  DSP48E1 desc60(.ACOUT(ACOUT_2[29:0]),.BCOUT({x_2_10[7:7],x_2_9[7:7],x_2_8[7:7],x_2_7[7:7],x_2_6[7:7],x_2_5[7:7],x_2_4[7:7],x_2_3[7:7],x_2_2[7:7],x_2_1[7:7],x_2_0[7:0]}),.CARRYCASCOUT(CARRYCASCOUT_2),.CARRYOUT(CARRYOUT_2[3:0]),.MULTSIGNOUT(MULTSIGNOUT_2),.OVERFLOW(OVERFLOW_2),.P({P_uc_2[47:12],un1_x_3[15:4]}),.PATTERNBDETECT(PATTERNBDETECT_2),.PATTERNDETECT(PATTERNDETECT_2),.PCOUT(PCOUT_2[47:0]),.UNDERFLOW(UNDERFLOW_2),.A({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,VCC,VCC,VCC}),.ACIN({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.ALUMODE({GND,GND,GND,GND}),.B({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.BCIN({x_1_10[7:7],x_1_9[7:7],x_1_8[7:7],x_1_7[7:7],x_1_6[7:7],x_1_5[7:7],x_1_4[7:7],x_1_3[7:7],x_1_2[7:7],x_1_1[7:7],x_1_0[7:0]}),.C({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.CARRYCASCIN(GND),.CARRYIN(GND),.CARRYINSEL({GND,GND,GND}),.CEA1(GND),.CEA2(GND),.CEAD(GND),.CEALUMODE(GND),.CEB1(GND),.CEB2(VCC),.CEC(GND),.CECARRYIN(GND),.CECTRL(GND),.CED(GND),.CEINMODE(GND),.CEM(GND),.CEP(VCC),.CLK(clk),.D({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND}),.INMODE({GND,GND,GND,GND,GND}),.MULTSIGNIN(GND),.OPMODE({GND,GND,GND,GND,VCC,GND,VCC}),.PCIN({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND}),.RSTA(GND),.RSTALLCARRYIN(GND),.RSTALUMODE(GND),.RSTB(GND),.RSTC(GND),.RSTCTRL(GND),.RSTD(GND),.RSTINMODE(GND),.RSTM(GND),.RSTP(GND));
defparam desc60.ACASCREG=0;
defparam desc60.ADREG=0;
defparam desc60.ALUMODEREG=0;
defparam desc60.AREG=0;
defparam desc60.AUTORESET_PATDET="NO_RESET";
defparam desc60.A_INPUT="DIRECT";
defparam desc60.BCASCREG=1;
defparam desc60.BREG=1;
defparam desc60.B_INPUT="CASCADE";
defparam desc60.CARRYINREG=0;
defparam desc60.CARRYINSELREG=0;
defparam desc60.CREG=1;
defparam desc60.DREG=0;
defparam desc60.INMODEREG=0;
defparam desc60.MREG=0;
defparam desc60.OPMODEREG=0;
defparam desc60.PREG=1;
defparam desc60.USE_DPORT="FALSE";
defparam desc60.USE_MULT="MULTIPLY";
defparam desc60.USE_SIMD="ONE48";
  DSP48E1 desc61(.ACOUT(ACOUT_3[29:0]),.BCOUT({x_6_10[7:7],x_6_9[7:7],x_6_8[7:7],x_6_7[7:7],x_6_6[7:7],x_6_5[7:7],x_6_4[7:7],x_6_3[7:7],x_6_2[7:7],x_6_1[7:7],x_6_0[7:0]}),.CARRYCASCOUT(CARRYCASCOUT_3),.CARRYOUT(CARRYOUT_3[3:0]),.MULTSIGNOUT(MULTSIGNOUT_3),.OVERFLOW(OVERFLOW_3),.P({P_uc_3[47:12],un1_x_8_0[15:4]}),.PATTERNBDETECT(PATTERNBDETECT_3),.PATTERNDETECT(PATTERNDETECT_3),.PCOUT(PCOUT_3[47:0]),.UNDERFLOW(UNDERFLOW_3),.A({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,VCC,VCC,VCC}),.ACIN({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.ALUMODE({GND,GND,GND,GND}),.B({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.BCIN({x_5_10[7:7],x_5_9[7:7],x_5_8[7:7],x_5_7[7:7],x_5_6[7:7],x_5_5[7:7],x_5_4[7:7],x_5_3[7:7],x_5_2[7:7],x_5_1[7:7],x_5_0[7:0]}),.C({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.CARRYCASCIN(GND),.CARRYIN(GND),.CARRYINSEL({GND,GND,GND}),.CEA1(GND),.CEA2(GND),.CEAD(GND),.CEALUMODE(GND),.CEB1(GND),.CEB2(VCC),.CEC(GND),.CECARRYIN(GND),.CECTRL(GND),.CED(GND),.CEINMODE(GND),.CEM(GND),.CEP(VCC),.CLK(clk),.D({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND}),.INMODE({GND,GND,GND,GND,GND}),.MULTSIGNIN(GND),.OPMODE({GND,GND,GND,GND,VCC,GND,VCC}),.PCIN({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND}),.RSTA(GND),.RSTALLCARRYIN(GND),.RSTALUMODE(GND),.RSTB(GND),.RSTC(GND),.RSTCTRL(GND),.RSTD(GND),.RSTINMODE(GND),.RSTM(GND),.RSTP(GND));
defparam desc61.ACASCREG=0;
defparam desc61.ADREG=0;
defparam desc61.ALUMODEREG=0;
defparam desc61.AREG=0;
defparam desc61.AUTORESET_PATDET="NO_RESET";
defparam desc61.A_INPUT="DIRECT";
defparam desc61.BCASCREG=1;
defparam desc61.BREG=1;
defparam desc61.B_INPUT="CASCADE";
defparam desc61.CARRYINREG=0;
defparam desc61.CARRYINSELREG=0;
defparam desc61.CREG=1;
defparam desc61.DREG=0;
defparam desc61.INMODEREG=0;
defparam desc61.MREG=0;
defparam desc61.OPMODEREG=0;
defparam desc61.PREG=1;
defparam desc61.USE_DPORT="FALSE";
defparam desc61.USE_MULT="MULTIPLY";
defparam desc61.USE_SIMD="ONE48";
  DSP48E1 desc62(.ACOUT(ACOUT_4[29:0]),.BCOUT({x_4_10[7:7],x_4_9[7:7],x_4_8[7:7],x_4_7[7:7],x_4_6[7:7],x_4_5[7:7],x_4_4[7:7],x_4_3[7:7],x_4_2[7:7],x_4_1[7:7],x_4_0[7:0]}),.CARRYCASCOUT(CARRYCASCOUT_4),.CARRYOUT(CARRYOUT_4[3:0]),.MULTSIGNOUT(MULTSIGNOUT_4),.OVERFLOW(OVERFLOW_4),.P({P_uc_4[47:15],un1_x_6_0[15:1]}),.PATTERNBDETECT(PATTERNBDETECT_4),.PATTERNDETECT(PATTERNDETECT_4),.PCOUT(PCOUT_4[47:0]),.UNDERFLOW(UNDERFLOW_4),.A({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,VCC,GND,VCC,GND,GND,GND}),.ACIN({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.ALUMODE({GND,GND,GND,GND}),.B({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.BCIN({x_3_10[7:7],x_3_9[7:7],x_3_8[7:7],x_3_7[7:7],x_3_6[7:7],x_3_5[7:7],x_3_4[7:7],x_3_3[7:7],x_3_2[7:7],x_3_1[7:7],x_3_0[7:0]}),.C({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.CARRYCASCIN(GND),.CARRYIN(GND),.CARRYINSEL({GND,GND,GND}),.CEA1(GND),.CEA2(GND),.CEAD(GND),.CEALUMODE(GND),.CEB1(GND),.CEB2(VCC),.CEC(GND),.CECARRYIN(GND),.CECTRL(GND),.CED(GND),.CEINMODE(GND),.CEM(GND),.CEP(VCC),.CLK(clk),.D({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND}),.INMODE({GND,GND,GND,GND,GND}),.MULTSIGNIN(GND),.OPMODE({GND,GND,GND,GND,VCC,GND,VCC}),.PCIN({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND}),.RSTA(GND),.RSTALLCARRYIN(GND),.RSTALUMODE(GND),.RSTB(GND),.RSTC(GND),.RSTCTRL(GND),.RSTD(GND),.RSTINMODE(GND),.RSTM(GND),.RSTP(GND));
defparam desc62.ACASCREG=0;
defparam desc62.ADREG=0;
defparam desc62.ALUMODEREG=0;
defparam desc62.AREG=0;
defparam desc62.AUTORESET_PATDET="NO_RESET";
defparam desc62.A_INPUT="DIRECT";
defparam desc62.BCASCREG=1;
defparam desc62.BREG=1;
defparam desc62.B_INPUT="CASCADE";
defparam desc62.CARRYINREG=0;
defparam desc62.CARRYINSELREG=0;
defparam desc62.CREG=1;
defparam desc62.DREG=0;
defparam desc62.INMODEREG=0;
defparam desc62.MREG=0;
defparam desc62.OPMODEREG=0;
defparam desc62.PREG=1;
defparam desc62.USE_DPORT="FALSE";
defparam desc62.USE_MULT="MULTIPLY";
defparam desc62.USE_SIMD="ONE48";
  DSP48E1 desc63(.ACOUT(ACOUT_5[29:0]),.BCOUT({x_3_10[7:7],x_3_9[7:7],x_3_8[7:7],x_3_7[7:7],x_3_6[7:7],x_3_5[7:7],x_3_4[7:7],x_3_3[7:7],x_3_2[7:7],x_3_1[7:7],x_3_0[7:0]}),.CARRYCASCOUT(CARRYCASCOUT_5),.CARRYOUT(CARRYOUT_5[3:0]),.MULTSIGNOUT(MULTSIGNOUT_5),.OVERFLOW(OVERFLOW_5),.P({P_uc_5[47:15],P_uc_4[14:14],un1_x_4[15:2]}),.PATTERNBDETECT(PATTERNBDETECT_5),.PATTERNDETECT(PATTERNDETECT_5),.PCOUT(PCOUT_5[47:0]),.UNDERFLOW(UNDERFLOW_5),.A({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,VCC,VCC,GND,GND,VCC}),.ACIN({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.ALUMODE({GND,GND,GND,GND}),.B({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.BCIN({x_2_10[7:7],x_2_9[7:7],x_2_8[7:7],x_2_7[7:7],x_2_6[7:7],x_2_5[7:7],x_2_4[7:7],x_2_3[7:7],x_2_2[7:7],x_2_1[7:7],x_2_0[7:0]}),.C({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.CARRYCASCIN(GND),.CARRYIN(GND),.CARRYINSEL({GND,GND,GND}),.CEA1(GND),.CEA2(GND),.CEAD(GND),.CEALUMODE(GND),.CEB1(GND),.CEB2(VCC),.CEC(GND),.CECARRYIN(GND),.CECTRL(GND),.CED(GND),.CEINMODE(GND),.CEM(GND),.CEP(VCC),.CLK(clk),.D({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND}),.INMODE({GND,GND,GND,GND,GND}),.MULTSIGNIN(GND),.OPMODE({GND,GND,GND,GND,VCC,GND,VCC}),.PCIN({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND}),.RSTA(GND),.RSTALLCARRYIN(GND),.RSTALUMODE(GND),.RSTB(GND),.RSTC(GND),.RSTCTRL(GND),.RSTD(GND),.RSTINMODE(GND),.RSTM(GND),.RSTP(GND));
defparam desc63.ACASCREG=0;
defparam desc63.ADREG=0;
defparam desc63.ALUMODEREG=0;
defparam desc63.AREG=0;
defparam desc63.AUTORESET_PATDET="NO_RESET";
defparam desc63.A_INPUT="DIRECT";
defparam desc63.BCASCREG=1;
defparam desc63.BREG=1;
defparam desc63.B_INPUT="CASCADE";
defparam desc63.CARRYINREG=0;
defparam desc63.CARRYINSELREG=0;
defparam desc63.CREG=1;
defparam desc63.DREG=0;
defparam desc63.INMODEREG=0;
defparam desc63.MREG=0;
defparam desc63.OPMODEREG=0;
defparam desc63.PREG=1;
defparam desc63.USE_DPORT="FALSE";
defparam desc63.USE_MULT="MULTIPLY";
defparam desc63.USE_SIMD="ONE48";
  DSP48E1 desc64(.ACOUT(ACOUT_6[29:0]),.BCOUT({x_5_10[7:7],x_5_9[7:7],x_5_8[7:7],x_5_7[7:7],x_5_6[7:7],x_5_5[7:7],x_5_4[7:7],x_5_3[7:7],x_5_2[7:7],x_5_1[7:7],x_5_0[7:0]}),.CARRYCASCOUT(CARRYCASCOUT_6),.CARRYOUT(CARRYOUT_6[3:0]),.MULTSIGNOUT(MULTSIGNOUT_6),.OVERFLOW(OVERFLOW_6),.P({P_uc_6[47:15],P_uc_5[14:14],un1_x_7_0[15:2]}),.PATTERNBDETECT(PATTERNBDETECT_6),.PATTERNDETECT(PATTERNDETECT_6),.PCOUT(PCOUT_6[47:0]),.UNDERFLOW(UNDERFLOW_6),.A({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,VCC,VCC,GND,GND,VCC}),.ACIN({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.ALUMODE({GND,GND,GND,GND}),.B({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.BCIN({x_4_10[7:7],x_4_9[7:7],x_4_8[7:7],x_4_7[7:7],x_4_6[7:7],x_4_5[7:7],x_4_4[7:7],x_4_3[7:7],x_4_2[7:7],x_4_1[7:7],x_4_0[7:0]}),.C({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.CARRYCASCIN(GND),.CARRYIN(GND),.CARRYINSEL({GND,GND,GND}),.CEA1(GND),.CEA2(GND),.CEAD(GND),.CEALUMODE(GND),.CEB1(GND),.CEB2(VCC),.CEC(GND),.CECARRYIN(GND),.CECTRL(GND),.CED(GND),.CEINMODE(GND),.CEM(GND),.CEP(VCC),.CLK(clk),.D({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND}),.INMODE({GND,GND,GND,GND,GND}),.MULTSIGNIN(GND),.OPMODE({GND,GND,GND,GND,VCC,GND,VCC}),.PCIN({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND}),.RSTA(GND),.RSTALLCARRYIN(GND),.RSTALUMODE(GND),.RSTB(GND),.RSTC(GND),.RSTCTRL(GND),.RSTD(GND),.RSTINMODE(GND),.RSTM(GND),.RSTP(GND));
defparam desc64.ACASCREG=0;
defparam desc64.ADREG=0;
defparam desc64.ALUMODEREG=0;
defparam desc64.AREG=0;
defparam desc64.AUTORESET_PATDET="NO_RESET";
defparam desc64.A_INPUT="DIRECT";
defparam desc64.BCASCREG=1;
defparam desc64.BREG=1;
defparam desc64.B_INPUT="CASCADE";
defparam desc64.CARRYINREG=0;
defparam desc64.CARRYINSELREG=0;
defparam desc64.CREG=1;
defparam desc64.DREG=0;
defparam desc64.INMODEREG=0;
defparam desc64.MREG=0;
defparam desc64.OPMODEREG=0;
defparam desc64.PREG=1;
defparam desc64.USE_DPORT="FALSE";
defparam desc64.USE_MULT="MULTIPLY";
defparam desc64.USE_SIMD="ONE48";
  DSP48E1 desc65(.ACOUT(ACOUT_7[29:0]),.BCOUT({x_10_10[7:7],x_10_9[7:7],x_10_8[7:7],x_10_7[7:7],x_10_6[7:7],x_10_5[7:7],x_10_4[7:7],x_10_3[7:7],x_10_2[7:7],x_10_1[7:7],x_10_0[7:0]}),.CARRYCASCOUT(CARRYCASCOUT_7),.CARRYOUT(CARRYOUT_7[3:0]),.MULTSIGNOUT(MULTSIGNOUT_7),.OVERFLOW(OVERFLOW_7),.P({P_uc_7[47:15],P_uc_6[14:14],P_uc_4[13:12],P_uc[11:11],un1_x_13_0_0[15:5]}),.PATTERNBDETECT(PATTERNBDETECT_7),.PATTERNDETECT(PATTERNDETECT_7),.PCOUT(PCOUT_7[47:0]),.UNDERFLOW(UNDERFLOW_7),.A({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,GND,VCC}),.ACIN({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.ALUMODE({GND,GND,GND,GND}),.B({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.BCIN({x_9_10[7:7],x_9_9[7:7],x_9_8[7:7],x_9_7[7:7],x_9_6[7:7],x_9_5[7:7],x_9_4[7:7],x_9_3[7:7],x_9_2[7:7],x_9_1[7:7],x_9_0[7:0]}),.C({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.CARRYCASCIN(GND),.CARRYIN(GND),.CARRYINSEL({GND,GND,GND}),.CEA1(GND),.CEA2(GND),.CEAD(GND),.CEALUMODE(GND),.CEB1(GND),.CEB2(VCC),.CEC(GND),.CECARRYIN(GND),.CECTRL(GND),.CED(GND),.CEINMODE(GND),.CEM(GND),.CEP(VCC),.CLK(clk),.D({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND}),.INMODE({GND,GND,GND,GND,GND}),.MULTSIGNIN(GND),.OPMODE({GND,GND,GND,GND,VCC,GND,VCC}),.PCIN({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND}),.RSTA(GND),.RSTALLCARRYIN(GND),.RSTALUMODE(GND),.RSTB(GND),.RSTC(GND),.RSTCTRL(GND),.RSTD(GND),.RSTINMODE(GND),.RSTM(GND),.RSTP(GND));
defparam desc65.ACASCREG=0;
defparam desc65.ADREG=0;
defparam desc65.ALUMODEREG=0;
defparam desc65.AREG=0;
defparam desc65.AUTORESET_PATDET="NO_RESET";
defparam desc65.A_INPUT="DIRECT";
defparam desc65.BCASCREG=1;
defparam desc65.BREG=1;
defparam desc65.B_INPUT="CASCADE";
defparam desc65.CARRYINREG=0;
defparam desc65.CARRYINSELREG=0;
defparam desc65.CREG=1;
defparam desc65.DREG=0;
defparam desc65.INMODEREG=0;
defparam desc65.MREG=0;
defparam desc65.OPMODEREG=0;
defparam desc65.PREG=1;
defparam desc65.USE_DPORT="FALSE";
defparam desc65.USE_MULT="MULTIPLY";
defparam desc65.USE_SIMD="ONE48";
  DSP48E1 desc66(.ACOUT(ACOUT_8[29:0]),.BCOUT({x_1_10[7:7],x_1_9[7:7],x_1_8[7:7],x_1_7[7:7],x_1_6[7:7],x_1_5[7:7],x_1_4[7:7],x_1_3[7:7],x_1_2[7:7],x_1_1[7:7],x_1_0[7:0]}),.CARRYCASCOUT(CARRYCASCOUT_8),.CARRYOUT(CARRYOUT_8[3:0]),.MULTSIGNOUT(MULTSIGNOUT_8),.OVERFLOW(OVERFLOW_8),.P({P_uc_8[47:15],P_uc_7[14:14],P_uc_5[13:12],P_uc_0[11:11],un1_x_2[15:5]}),.PATTERNBDETECT(PATTERNBDETECT_8),.PATTERNDETECT(PATTERNDETECT_8),.PCOUT(PCOUT_8[47:0]),.UNDERFLOW(UNDERFLOW_8),.A({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,GND,VCC}),.ACIN({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.ALUMODE({GND,GND,GND,GND}),.B({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.BCIN({x_0_10[7:7],x_0_9[7:7],x_0_8[7:7],x_0_7[7:7],x_0_6[7:7],x_0_5[7:7],x_0_4[7:7],x_0_3[7:7],x_0_2[7:7],x_0_1[7:7],x_0_0[7:0]}),.C({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.CARRYCASCIN(GND),.CARRYIN(GND),.CARRYINSEL({GND,GND,GND}),.CEA1(GND),.CEA2(GND),.CEAD(GND),.CEALUMODE(GND),.CEB1(GND),.CEB2(VCC),.CEC(GND),.CECARRYIN(GND),.CECTRL(GND),.CED(GND),.CEINMODE(GND),.CEM(GND),.CEP(VCC),.CLK(clk),.D({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND}),.INMODE({GND,GND,GND,GND,GND}),.MULTSIGNIN(GND),.OPMODE({GND,GND,GND,GND,VCC,GND,VCC}),.PCIN({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND}),.RSTA(GND),.RSTALLCARRYIN(GND),.RSTALUMODE(GND),.RSTB(GND),.RSTC(GND),.RSTCTRL(GND),.RSTD(GND),.RSTINMODE(GND),.RSTM(GND),.RSTP(GND));
defparam desc66.ACASCREG=0;
defparam desc66.ADREG=0;
defparam desc66.ALUMODEREG=0;
defparam desc66.AREG=0;
defparam desc66.AUTORESET_PATDET="NO_RESET";
defparam desc66.A_INPUT="DIRECT";
defparam desc66.BCASCREG=1;
defparam desc66.BREG=1;
defparam desc66.B_INPUT="CASCADE";
defparam desc66.CARRYINREG=0;
defparam desc66.CARRYINSELREG=0;
defparam desc66.CREG=1;
defparam desc66.DREG=0;
defparam desc66.INMODEREG=0;
defparam desc66.MREG=0;
defparam desc66.OPMODEREG=0;
defparam desc66.PREG=1;
defparam desc66.USE_DPORT="FALSE";
defparam desc66.USE_MULT="MULTIPLY";
defparam desc66.USE_SIMD="ONE48";
  DSP48E1 desc67(.ACOUT(ACOUT_9[29:0]),.BCOUT(BCOUT_9[17:0]),.CARRYCASCOUT(CARRYCASCOUT_9),.CARRYOUT(CARRYOUT_9[3:0]),.MULTSIGNOUT(MULTSIGNOUT_9),.OVERFLOW(OVERFLOW_9),.P({P_uc_9[47:15],P_uc_8[14:14],P_uc_6[13:12],P_uc_1[11:11],un1_x_9_0[15:5]}),.PATTERNBDETECT(PATTERNBDETECT_9),.PATTERNDETECT(PATTERNDETECT_9),.PCOUT(PCOUT_9[47:0]),.UNDERFLOW(UNDERFLOW_9),.A({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,GND,VCC}),.ACIN({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.ALUMODE({GND,GND,GND,GND}),.B({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.BCIN({x_6_10[7:7],x_6_9[7:7],x_6_8[7:7],x_6_7[7:7],x_6_6[7:7],x_6_5[7:7],x_6_4[7:7],x_6_3[7:7],x_6_2[7:7],x_6_1[7:7],x_6_0[7:0]}),.C({VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC,VCC}),.CARRYCASCIN(GND),.CARRYIN(GND),.CARRYINSEL({GND,GND,GND}),.CEA1(GND),.CEA2(GND),.CEAD(GND),.CEALUMODE(GND),.CEB1(GND),.CEB2(VCC),.CEC(GND),.CECARRYIN(GND),.CECTRL(GND),.CED(GND),.CEINMODE(GND),.CEM(GND),.CEP(VCC),.CLK(clk),.D({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND}),.INMODE({GND,GND,GND,GND,GND}),.MULTSIGNIN(GND),.OPMODE({GND,GND,GND,GND,VCC,GND,VCC}),.PCIN({GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND,GND}),.RSTA(GND),.RSTALLCARRYIN(GND),.RSTALUMODE(GND),.RSTB(GND),.RSTC(GND),.RSTCTRL(GND),.RSTD(GND),.RSTINMODE(GND),.RSTM(GND),.RSTP(GND));
defparam desc67.ACASCREG=0;
defparam desc67.ADREG=0;
defparam desc67.ALUMODEREG=0;
defparam desc67.AREG=0;
defparam desc67.AUTORESET_PATDET="NO_RESET";
defparam desc67.A_INPUT="DIRECT";
defparam desc67.BCASCREG=1;
defparam desc67.BREG=1;
defparam desc67.B_INPUT="CASCADE";
defparam desc67.CARRYINREG=0;
defparam desc67.CARRYINSELREG=0;
defparam desc67.CREG=1;
defparam desc67.DREG=0;
defparam desc67.INMODEREG=0;
defparam desc67.MREG=0;
defparam desc67.OPMODEREG=0;
defparam desc67.PREG=1;
defparam desc67.USE_DPORT="FALSE";
defparam desc67.USE_MULT="MULTIPLY";
defparam desc67.USE_SIMD="ONE48";
  LUT3 un84_sop_0_0_0_11_6_0_axb_1_lut6_2_o6(.I0(un1_x_12_0_0[5:5]),.I1(un1_x_13_0_0[6:6]),.I2(un1_x_14_0_0[5:5]),.O(un84_sop_0_0_0_11_6_0_axb_1));
defparam un84_sop_0_0_0_11_6_0_axb_1_lut6_2_o6.INIT=8'h96;
  LUT3 un84_sop_0_0_0_11_6_0_axb_1_lut6_2_o5(.I0(un1_x_12_0_0[5:5]),.I1(un1_x_13_0_0[6:6]),.I2(un1_x_14_0_0[5:5]),.O(un84_sop_0_0_0_11_6_0_axb_1_lut6_2_O5));
defparam un84_sop_0_0_0_11_6_0_axb_1_lut6_2_o5.INIT=8'hE8;
  LUT3 un84_sop_0_0_0_6_6_0_axb_1_lut6_2_o6(.I0(un1_x_7_0[3:3]),.I1(un1_x_8_0[5:5]),.I2(un1_x_9_0[6:6]),.O(un84_sop_0_0_0_6_6_0_axb_1));
defparam un84_sop_0_0_0_6_6_0_axb_1_lut6_2_o6.INIT=8'h96;
  LUT3 un84_sop_0_0_0_6_6_0_axb_1_lut6_2_o5(.I0(un1_x_7_0[3:3]),.I1(un1_x_8_0[5:5]),.I2(un1_x_9_0[6:6]),.O(un84_sop_0_0_0_6_6_0_axb_1_lut6_2_O5));
defparam un84_sop_0_0_0_6_6_0_axb_1_lut6_2_o5.INIT=8'hE8;
  LUT3 un84_sop_0_0_0_1_6_8_axb_2_lut6_2_o6(.I0(un84_sop_0_0_0_10_0[5:5]),.I1(x_4[0:0]),.I2(x_4[2:2]),.O(un84_sop_0_0_0_1_6_8_axb_2));
defparam un84_sop_0_0_0_1_6_8_axb_2_lut6_2_o6.INIT=8'h96;
  LUT3 un84_sop_0_0_0_1_6_8_axb_2_lut6_2_o5(.I0(un84_sop_0_0_0_10_0[5:5]),.I1(x_4[0:0]),.I2(x_4[2:2]),.O(un84_sop_0_0_0_1_6_8_axb_2_lut6_2_O5));
defparam un84_sop_0_0_0_1_6_8_axb_2_lut6_2_o5.INIT=8'hE8;
  LUT3 un84_sop_1_6_0_axb_1_lut6_2_o6(.I0(un1_x_1[5:5]),.I1(un1_x_2[6:6]),.I2(un1_x_3[5:5]),.O(un84_sop_1_6_0_axb_1));
defparam un84_sop_1_6_0_axb_1_lut6_2_o6.INIT=8'h96;
  LUT3 un84_sop_1_6_0_axb_1_lut6_2_o5(.I0(un1_x_1[5:5]),.I1(un1_x_2[6:6]),.I2(un1_x_3[5:5]),.O(un84_sop_1_6_0_axb_1_lut6_2_O5));
defparam un84_sop_1_6_0_axb_1_lut6_2_o5.INIT=8'hE8;
endmodule