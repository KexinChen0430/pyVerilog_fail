module header
	// Internal signals
	// Generated Signal List
	// End of Generated Signal List
	// %COMPILER_OPTS%
	// Generated Signal Assignments
	// Generated Instances and Port Mappings
		// Generated Instance Port Map for inst_eca
		inst_eca_e inst_eca (
		);
		// End of Generated Instance Port Map for inst_eca
		// Generated Instance Port Map for inst_ecb
		inst_ecb_e inst_ecb (
		);
		// End of Generated Instance Port Map for inst_ecb
		// Generated Instance Port Map for inst_ecc
		inst_ecc_e inst_ecc (
		);
		// End of Generated Instance Port Map for inst_ecc
endmodule