module main;
   test tt();
   defparam foo = 3; /* This should generate an error. */
endmodule