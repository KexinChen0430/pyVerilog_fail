module mig_7series_v1_9_infrastructure #
  (
   parameter SIMULATION      = "FALSE",  // Should be TRUE during design simulations and
                                         // FALSE during implementations
   parameter TCQ             = 100,      // clk->out delay (sim only)
   parameter CLKIN_PERIOD    = 3000,     // Memory clock period
   parameter nCK_PER_CLK     = 2,        // Fabric clk period:Memory clk period
   parameter SYSCLK_TYPE     = "DIFFERENTIAL",
                                         // input clock type
                                         // "DIFFERENTIAL","SINGLE_ENDED"
   parameter UI_EXTRA_CLOCKS = "FALSE",
                                         // Generates extra clocks as
                                         // 1/2, 1/4 and 1/8 of fabrick clock.
                                         // Valid for DDR2/DDR3 AXI interfaces
                                         // based on GUI selection
   parameter CLKFBOUT_MULT   = 4,        // write PLL VCO multiplier
   parameter DIVCLK_DIVIDE   = 1,        // write PLL VCO divisor
   parameter CLKOUT0_PHASE   = 45.0,     // VCO output divisor for clkout0
   parameter CLKOUT0_DIVIDE   = 16,      // VCO output divisor for PLL clkout0
   parameter CLKOUT1_DIVIDE   = 4,       // VCO output divisor for PLL clkout1
   parameter CLKOUT2_DIVIDE   = 64,      // VCO output divisor for PLL clkout2
   parameter CLKOUT3_DIVIDE   = 16,      // VCO output divisor for PLL clkout3
   parameter MMCM_CLKOUT0_EN       = "FALSE",  // Enabled (or) Disable MMCM clkout0
   parameter MMCM_CLKOUT1_EN       = "FALSE",  // Enabled (or) Disable MMCM clkout1
   parameter MMCM_CLKOUT2_EN       = "FALSE",  // Enabled (or) Disable MMCM clkout2
   parameter MMCM_CLKOUT3_EN       = "FALSE",  // Enabled (or) Disable MMCM clkout3
   parameter MMCM_CLKOUT4_EN       = "FALSE",  // Enabled (or) Disable MMCM clkout4
   parameter MMCM_CLKOUT0_DIVIDE   = 1,  // VCO output divisor for MMCM clkout0
   parameter MMCM_CLKOUT1_DIVIDE   = 1,  // VCO output divisor for MMCM clkout1
   parameter MMCM_CLKOUT2_DIVIDE   = 1,  // VCO output divisor for MMCM clkout2
   parameter MMCM_CLKOUT3_DIVIDE   = 1,  // VCO output divisor for MMCM clkout3
   parameter MMCM_CLKOUT4_DIVIDE   = 1,  // VCO output divisor for MMCM clkout4
   parameter RST_ACT_LOW  = 1
   )
  (
   // Clock inputs
   input  mmcm_clk,           // System clock diff input
   // System reset input
   input  sys_rst,            // core reset from user application
   // PLLE2/IDELAYCTRL Lock status
   input  iodelay_ctrl_rdy,   // IDELAYCTRL lock status
   // Clock outputs
   output clk,                // fabric clock freq ; either  half rate or quarter rate and is
                              // determined by  PLL parameters settings.
   output mem_refclk,         // equal to  memory clock
   output freq_refclk,        // freq above 400 MHz:  set freq_refclk = mem_refclk
                              // freq below 400 MHz:  set freq_refclk = 2* mem_refclk or 4* mem_refclk;
                              // to hard PHY for phaser
   output sync_pulse,         // exactly 1/16 of mem_refclk and the sync pulse is exactly 1 memref_clk wide
   output auxout_clk,         // IO clk used to clock out Aux_Out ports
   output ui_addn_clk_0,      // MMCM out0 clk
   output ui_addn_clk_1,      // MMCM out1 clk
   output ui_addn_clk_2,      // MMCM out2 clk
   output ui_addn_clk_3,      // MMCM out3 clk
   output ui_addn_clk_4,      // MMCM out4 clk
   output pll_locked,         // locked output from PLLE2_ADV
   output mmcm_locked,        // locked output from MMCME2_ADV
   // Reset outputs
   output rstdiv0             // Reset CLK and CLKDIV logic (incl I/O),
   ,output rst_phaser_ref
   ,input  ref_dll_lock
	,output	ref_clk
	,input rst_tmp_idelay,
	input rst_ref
   );
  // # of clock cycles to delay deassertion of reset. Needs to be a fairly
  // high number not so much for metastability protection, but to give time
  // for reset (i.e. stable clock cycles) to propagate through all state
  // machines and to all control signals (i.e. not all control signals have
  // resets, instead they rely on base state logic being reset, and the effect
  // of that reset propagating through the logic). Need this because we may not
  // be getting stable clock cycles while reset asserted (i.e. since reset
  // depends on DCM lock status)
  localparam RST_SYNC_NUM = 25;
  // Round up for clk reset delay to ensure that CLKDIV reset deassertion
  // occurs at same time or after CLK reset deassertion (still need to
  // consider route delay - add one or two extra cycles to be sure!)
  localparam RST_DIV_SYNC_NUM = (RST_SYNC_NUM+1)/2;
  // Input clock is assumed to be equal to the memory clock frequency
  // User should change the parameter as necessary if a different input
  // clock frequency is used
  localparam real CLKIN1_PERIOD_NS = CLKIN_PERIOD / 1000.0;
  localparam CLKOUT4_DIVIDE = 2 * CLKOUT1_DIVIDE;
  localparam integer VCO_PERIOD
             = (CLKIN1_PERIOD_NS * DIVCLK_DIVIDE * 1000) / CLKFBOUT_MULT;
  localparam CLKOUT0_PERIOD = VCO_PERIOD * CLKOUT0_DIVIDE;
  localparam CLKOUT1_PERIOD = VCO_PERIOD * CLKOUT1_DIVIDE;
  localparam CLKOUT2_PERIOD = VCO_PERIOD * CLKOUT2_DIVIDE;
  localparam CLKOUT3_PERIOD = VCO_PERIOD * CLKOUT3_DIVIDE;
  localparam CLKOUT4_PERIOD = VCO_PERIOD * CLKOUT4_DIVIDE;
  localparam CLKOUT4_PHASE  = (SIMULATION == "TRUE") ? 22.5 : 168.75;
  localparam real CLKOUT3_PERIOD_NS = CLKOUT3_PERIOD / 1000.0;
  localparam real CLKOUT4_PERIOD_NS = CLKOUT4_PERIOD / 1000.0;
  localparam CLKOUT5_DIVIDE   = 4;
  localparam CLKOUT5_PHASE   = 0.000;
  //synthesis translate_off
  initial begin
    $display("############# Write Clocks PLLE2_ADV Parameters #############\n");
    $display("nCK_PER_CLK      = %7d",   nCK_PER_CLK     );
    $display("CLK_PERIOD       = %7d",   CLKIN_PERIOD    );
    $display("CLKIN1_PERIOD    = %7.3f", CLKIN1_PERIOD_NS);
    $display("DIVCLK_DIVIDE    = %7d",   DIVCLK_DIVIDE   );
    $display("CLKFBOUT_MULT    = %7d",   CLKFBOUT_MULT );
    $display("VCO_PERIOD       = %7d",   VCO_PERIOD      );
    $display("CLKOUT0_DIVIDE_F = %7d",   CLKOUT0_DIVIDE  );
    $display("CLKOUT1_DIVIDE   = %7d",   CLKOUT1_DIVIDE  );
    $display("CLKOUT2_DIVIDE   = %7d",   CLKOUT2_DIVIDE  );
    $display("CLKOUT3_DIVIDE   = %7d",   CLKOUT3_DIVIDE  );
    $display("CLKOUT0_PERIOD   = %7d",   CLKOUT0_PERIOD  );
    $display("CLKOUT1_PERIOD   = %7d",   CLKOUT1_PERIOD  );
    $display("CLKOUT2_PERIOD   = %7d",   CLKOUT2_PERIOD  );
    $display("CLKOUT3_PERIOD   = %7d",   CLKOUT3_PERIOD  );
    $display("CLKOUT4_PERIOD   = %7d",   CLKOUT4_PERIOD  );
    $display("############################################################\n");
  end
  //synthesis translate_on
  wire                       clk_bufg;
  wire                       clk_pll;
  wire                       clkfbout_pll;
  wire                       mmcm_clkfbout;
  (* keep = "true", max_fanout = 10 *) wire                       pll_locked_i
                             /* synthesis syn_maxfan = 10 */;
  reg [RST_DIV_SYNC_NUM-2:0] rstdiv0_sync_r;
  wire                       rst_tmp;
  (* keep = "true", max_fanout = 10 *) reg rstdiv0_sync_r1
                             /* synthesis syn_maxfan = 10 */;
  wire                       sys_rst_act_hi;
  wire                       rst_tmp_phaser_ref;
  (* keep = "true", max_fanout = 10 *) reg [RST_DIV_SYNC_NUM-1:0] rst_phaser_ref_sync_r
                             /* synthesis syn_maxfan = 10 */;
  // Instantiation of the MMCM primitive
  wire        clkfbout;
  wire        MMCM_Locked_i;
  wire        mmcm_clkout0;
  wire        mmcm_clkout1;
  wire        mmcm_clkout2;
  wire        mmcm_clkout3;
  wire        mmcm_clkout4;
  wire        ref_clk_mmcm_bufg;
  assign sys_rst_act_hi = RST_ACT_LOW ? ~sys_rst: sys_rst;
  // Assign global clocks:
  //   2. clk     : Half rate / Quarter rate(used for majority of internal logic)
  assign clk        = clk_bufg;
  assign pll_locked = pll_locked_i & MMCM_Locked_i;
  assign mmcm_locked = MMCM_Locked_i;
  assign	ref_clk = ref_clk_mmcm_bufg;
  // Global base clock generation and distribution
  // NOTES ON CALCULTING PROPER VCO FREQUENCY
  //  1. VCO frequency =
  //     1/((DIVCLK_DIVIDE * CLKIN_PERIOD)/(CLKFBOUT_MULT * nCK_PER_CLK))
  //  2. VCO frequency must be in the range [TBD, TBD]
  PLLE2_ADV #
    (
     .BANDWIDTH          ("OPTIMIZED"),
     .COMPENSATION       ("INTERNAL"),
     .STARTUP_WAIT       ("FALSE"),
     .CLKOUT0_DIVIDE     (CLKOUT0_DIVIDE),  // 4 freq_ref
     .CLKOUT1_DIVIDE     (CLKOUT1_DIVIDE),  // 4 mem_ref
     .CLKOUT2_DIVIDE     (CLKOUT2_DIVIDE),  // 16 sync
     .CLKOUT3_DIVIDE     (CLKOUT3_DIVIDE),  // 16 sysclk
     .CLKOUT4_DIVIDE     (CLKOUT4_DIVIDE),
     .CLKOUT5_DIVIDE     (CLKOUT5_DIVIDE),
     .DIVCLK_DIVIDE      (DIVCLK_DIVIDE),
     .CLKFBOUT_MULT      (CLKFBOUT_MULT),
     .CLKFBOUT_PHASE     (0.000),
     .CLKIN1_PERIOD      (CLKIN1_PERIOD_NS),
     .CLKIN2_PERIOD      (),
     .CLKOUT0_DUTY_CYCLE (0.500),
     .CLKOUT0_PHASE      (CLKOUT0_PHASE),
     .CLKOUT1_DUTY_CYCLE (0.500),
     .CLKOUT1_PHASE      (0.000),
     .CLKOUT2_DUTY_CYCLE (1.0/16.0),
     .CLKOUT2_PHASE      (9.84375),     // PHASE shift is required for sync pulse generation.
     .CLKOUT3_DUTY_CYCLE (0.500),
     .CLKOUT3_PHASE      (0.000),
     .CLKOUT4_DUTY_CYCLE (0.500),
     .CLKOUT4_PHASE      (CLKOUT4_PHASE),
     .CLKOUT5_DUTY_CYCLE (0.500),
     .CLKOUT5_PHASE      (CLKOUT5_PHASE),
     .REF_JITTER1        (0.010),
     .REF_JITTER2        (0.010)
     )
    plle2_i
      (
       .CLKFBOUT (pll_clkfbout),
       .CLKOUT0  (freq_refclk),
       .CLKOUT1  (mem_refclk),
       .CLKOUT2  (sync_pulse),  // always 1/16 of mem_ref_clk
       .CLKOUT3  (pll_clk3),
       .CLKOUT4  (auxout_clk_i),
       .CLKOUT5  (ref_clk_mmcm),
       .DO       (),
       .DRDY     (),
       .LOCKED   (pll_locked_i),
       .CLKFBIN  (pll_clkfbout),
       .CLKIN1   (mmcm_clk),
       .CLKIN2   (),
       .CLKINSEL (1'b1),
       .DADDR    (7'b0),
       .DCLK     (1'b0),
       .DEN      (1'b0),
       .DI       (16'b0),
       .DWE      (1'b0),
       .PWRDWN   (1'b0),
       .RST      ( sys_rst_act_hi)
       );
  BUFH u_bufh_auxout_clk
    (
     .O (auxout_clk),
     .I (auxout_clk_i)
     );
  BUFG u_bufg_clkdiv0
    (
     .O (clk_bufg),
     .I (clk_pll_i)
     );
	BUFG u_bufg_refclk
	(
		.O(ref_clk_mmcm_bufg),
		.I(ref_clk_mmcm)
		);
  localparam  integer MMCM_VCO_MIN_FREQ     = 600;
  localparam  integer MMCM_VCO_MAX_FREQ     = 1200; // This is the maximum VCO frequency for a -1 part
  localparam  real    MMCM_VCO_MIN_PERIOD   = 1000000.0/MMCM_VCO_MAX_FREQ;
  localparam  real    MMCM_VCO_MAX_PERIOD   = 1000000.0/MMCM_VCO_MIN_FREQ;
  localparam  real    MMCM_MULT_F_MID       = CLKOUT3_PERIOD/(MMCM_VCO_MAX_PERIOD*0.75);
  localparam  real    MMCM_EXPECTED_PERIOD  = CLKOUT3_PERIOD / MMCM_MULT_F_MID;
  localparam  real    MMCM_MULT_F           = ((MMCM_EXPECTED_PERIOD > MMCM_VCO_MAX_PERIOD) ? MMCM_MULT_F_MID + 1.0 : MMCM_MULT_F_MID);
  localparam  real    MMCM_VCO_FREQ         = MMCM_MULT_F / (1 * CLKOUT3_PERIOD_NS);
  localparam  real    MMCM_VCO_PERIOD       = (CLKOUT3_PERIOD_NS * 1000) / MMCM_MULT_F;
  //synthesis translate_off
  initial begin
    $display("############# MMCME2_ADV Parameters #############\n");
    $display("MMCM_VCO_MIN_PERIOD   = %7.3f", MMCM_VCO_MIN_PERIOD);
    $display("MMCM_VCO_MAX_PERIOD   = %7.3f", MMCM_VCO_MAX_PERIOD);
    $display("MMCM_MULT_F_MID       = %7.3f", MMCM_MULT_F_MID);
    $display("MMCM_EXPECTED_PERIOD  = %7.3f", MMCM_EXPECTED_PERIOD);
    $display("MMCM_MULT_F           = %7.3f", MMCM_MULT_F);
    $display("CLKOUT3_PERIOD_NS     = %7.3f", CLKOUT3_PERIOD_NS);
    $display("MMCM_VCO_FREQ (MHz)   = %7.3f", MMCM_VCO_FREQ*1000.0);
    $display("MMCM_VCO_PERIOD       = %7.3f", MMCM_VCO_PERIOD);
    $display("#################################################\n");
  end
  //synthesis translate_on
  generate
    if (UI_EXTRA_CLOCKS == "TRUE") begin: gen_ui_extra_clocks
      localparam MMCM_CLKOUT0_DIVIDE_CAL = (MMCM_CLKOUT0_EN == "TRUE") ? MMCM_CLKOUT0_DIVIDE : MMCM_MULT_F;
      localparam MMCM_CLKOUT1_DIVIDE_CAL = (MMCM_CLKOUT1_EN == "TRUE") ? MMCM_CLKOUT1_DIVIDE : MMCM_MULT_F;
      localparam MMCM_CLKOUT2_DIVIDE_CAL = (MMCM_CLKOUT2_EN == "TRUE") ? MMCM_CLKOUT2_DIVIDE : MMCM_MULT_F;
      localparam MMCM_CLKOUT3_DIVIDE_CAL = (MMCM_CLKOUT3_EN == "TRUE") ? MMCM_CLKOUT3_DIVIDE : MMCM_MULT_F;
      localparam MMCM_CLKOUT4_DIVIDE_CAL = (MMCM_CLKOUT4_EN == "TRUE") ? MMCM_CLKOUT4_DIVIDE : MMCM_MULT_F;
      MMCME2_ADV
      #(.BANDWIDTH            ("HIGH"),
        .CLKOUT4_CASCADE      ("FALSE"),
        .COMPENSATION         ("BUF_IN"),
        .STARTUP_WAIT         ("FALSE"),
        .DIVCLK_DIVIDE        (1),
        .CLKFBOUT_MULT_F      (MMCM_MULT_F),
        .CLKFBOUT_PHASE       (0.000),
        .CLKFBOUT_USE_FINE_PS ("FALSE"),
        .CLKOUT0_DIVIDE_F     (MMCM_CLKOUT0_DIVIDE_CAL),
        .CLKOUT0_PHASE        (0.000),
        .CLKOUT0_DUTY_CYCLE   (0.500),
        .CLKOUT0_USE_FINE_PS  ("FALSE"),
        .CLKOUT1_DIVIDE       (MMCM_CLKOUT1_DIVIDE_CAL),
        .CLKOUT1_PHASE        (0.000),
        .CLKOUT1_DUTY_CYCLE   (0.500),
        .CLKOUT1_USE_FINE_PS  ("FALSE"),
        .CLKOUT2_DIVIDE       (MMCM_CLKOUT2_DIVIDE_CAL),
        .CLKOUT2_PHASE        (0.000),
        .CLKOUT2_DUTY_CYCLE   (0.500),
        .CLKOUT2_USE_FINE_PS  ("FALSE"),
        .CLKOUT3_DIVIDE       (MMCM_CLKOUT3_DIVIDE_CAL),
        .CLKOUT3_PHASE        (0.000),
        .CLKOUT3_DUTY_CYCLE   (0.500),
        .CLKOUT3_USE_FINE_PS  ("FALSE"),
        .CLKOUT4_DIVIDE       (MMCM_CLKOUT4_DIVIDE_CAL),
        .CLKOUT4_PHASE        (0.000),
        .CLKOUT4_DUTY_CYCLE   (0.500),
        .CLKOUT4_USE_FINE_PS  ("FALSE"),
        .CLKIN1_PERIOD        (CLKOUT3_PERIOD_NS),
        .REF_JITTER1          (0.000))
      mmcm_i
        // Output clocks
       (.CLKFBOUT            (clk_pll_i),
        .CLKFBOUTB           (),
        .CLKOUT0             (mmcm_clkout0),
        .CLKOUT0B            (),
        .CLKOUT1             (mmcm_clkout1),
        .CLKOUT1B            (),
        .CLKOUT2             (mmcm_clkout2),
        .CLKOUT2B            (),
        .CLKOUT3             (mmcm_clkout3),
        .CLKOUT3B            (),
        .CLKOUT4             (mmcm_clkout4),
        .CLKOUT5             (),
        .CLKOUT6             (),
         // Input clock control
        .CLKFBIN             (clk_bufg),      // From BUFH network
        .CLKIN1              (pll_clk3),      // From PLL
        .CLKIN2              (1'b0),
         // Tied to always select the primary input clock
        .CLKINSEL            (1'b1),
        // Ports for dynamic reconfiguration
        .DADDR               (7'h0),
        .DCLK                (1'b0),
        .DEN                 (1'b0),
        .DI                  (16'h0),
        .DO                  (),
        .DRDY                (),
        .DWE                 (1'b0),
        // Ports for dynamic phase shift
        .PSCLK               (1'b0),
        .PSEN                (1'b0),
        .PSINCDEC            (1'b0),
        .PSDONE              (),
        // Other control and status signals
        .LOCKED              (MMCM_Locked_i),
        .CLKINSTOPPED        (),
        .CLKFBSTOPPED        (),
        .PWRDWN              (1'b0),
        .RST                 (~pll_locked_i));
      BUFG u_bufg_ui_addn_clk_0
        (
         .O (ui_addn_clk_0),
         .I (mmcm_clkout0)
         );
      BUFG u_bufg_ui_addn_clk_1
        (
         .O (ui_addn_clk_1),
         .I (mmcm_clkout1)
         );
      BUFG u_bufg_ui_addn_clk_2
        (
         .O (ui_addn_clk_2),
         .I (mmcm_clkout2)
         );
      BUFG u_bufg_ui_addn_clk_3
        (
         .O (ui_addn_clk_3),
         .I (mmcm_clkout3)
         );
      BUFG u_bufg_ui_addn_clk_4
        (
         .O (ui_addn_clk_4),
         .I (mmcm_clkout4)
         );
    end else begin: gen_mmcm
      MMCME2_ADV
      #(.BANDWIDTH            ("HIGH"),
        .CLKOUT4_CASCADE      ("FALSE"),
        .COMPENSATION         ("BUF_IN"),
        .STARTUP_WAIT         ("FALSE"),
        .DIVCLK_DIVIDE        (1),
        .CLKFBOUT_MULT_F      (MMCM_MULT_F),
        .CLKFBOUT_PHASE       (0.000),
        .CLKFBOUT_USE_FINE_PS ("FALSE"),
        .CLKOUT0_DIVIDE_F     (MMCM_MULT_F),
        .CLKOUT0_PHASE        (0.000),
        .CLKOUT0_DUTY_CYCLE   (0.500),
        .CLKOUT0_USE_FINE_PS  ("FALSE"),
        .CLKOUT1_DIVIDE       (),
        .CLKOUT1_PHASE        (0.000),
        .CLKOUT1_DUTY_CYCLE   (0.500),
        .CLKOUT1_USE_FINE_PS  ("FALSE"),
        .CLKIN1_PERIOD        (CLKOUT3_PERIOD_NS),
        .REF_JITTER1          (0.000))
      mmcm_i
        // Output clocks
       (.CLKFBOUT            (clk_pll_i),
        .CLKFBOUTB           (),
        .CLKOUT0             (),
        .CLKOUT0B            (),
        .CLKOUT1             (),
        .CLKOUT1B            (),
        .CLKOUT2             (),
        .CLKOUT2B            (),
        .CLKOUT3             (),
        .CLKOUT3B            (),
        .CLKOUT4             (),
        .CLKOUT5             (),
        .CLKOUT6             (),
         // Input clock control
        .CLKFBIN             (clk_bufg),      // From BUFH network
        .CLKIN1              (pll_clk3),      // From PLL
        .CLKIN2              (1'b0),
         // Tied to always select the primary input clock
        .CLKINSEL            (1'b1),
        // Ports for dynamic reconfiguration
        .DADDR               (7'h0),
        .DCLK                (1'b0),
        .DEN                 (1'b0),
        .DI                  (16'h0),
        .DO                  (),
        .DRDY                (),
        .DWE                 (1'b0),
        // Ports for dynamic phase shift
        .PSCLK               (1'b0),
        .PSEN                (1'b0),
        .PSINCDEC            (1'b0),
        .PSDONE              (),
        // Other control and status signals
        .LOCKED              (MMCM_Locked_i),
        .CLKINSTOPPED        (),
        .CLKFBSTOPPED        (),
        .PWRDWN              (1'b0),
        .RST                 (~pll_locked_i));
   end
  endgenerate
  // RESET SYNCHRONIZATION DESCRIPTION:
  //  Various resets are generated to ensure that:
  //   1. All resets are synchronously deasserted with respect to the clock
  //      domain they are interfacing to. There are several different clock
  //      domains - each one will receive a synchronized reset.
  //   2. The reset deassertion order starts with deassertion of SYS_RST,
  //      followed by deassertion of resets for various parts of the design
  //      (see "RESET ORDER" below) based on the lock status of PLLE2s.
  // RESET ORDER:
  //   1. User deasserts SYS_RST
  //   2. Reset PLLE2 and IDELAYCTRL
  //   3. Wait for PLLE2 and IDELAYCTRL to lock
  //   4. Release reset for all I/O primitives and internal logic
  // OTHER NOTES:
  //   1. Asynchronously assert reset. This way we can assert reset even if
  //      there is no clock (needed for things like 3-stating output buffers
  //      to prevent initial bus contention). Reset deassertion is synchronous.
  // CLKDIV logic reset
  // Wait for PLLE2 and IDELAYCTRL to lock before releasing reset
  // current O,25.0 unisim phaser_ref never locks.  Need to find out why .
  assign rst_tmp = sys_rst_act_hi | ~iodelay_ctrl_rdy |
                   ~ref_dll_lock | ~MMCM_Locked_i;
  always @(posedge clk_bufg or posedge rst_tmp) begin
    if (rst_tmp) begin
      rstdiv0_sync_r  <= #TCQ {RST_DIV_SYNC_NUM-1{1'b1}};
      rstdiv0_sync_r1 <= #TCQ 1'b1 ;
    end else begin
      rstdiv0_sync_r  <= #TCQ rstdiv0_sync_r << 1;
      rstdiv0_sync_r1 <= #TCQ rstdiv0_sync_r[RST_DIV_SYNC_NUM-2];
    end
  end
  assign rstdiv0 = rstdiv0_sync_r1 ;
  assign rst_tmp_phaser_ref = sys_rst_act_hi | ~pll_locked_i | ~iodelay_ctrl_rdy;
  always @(posedge clk_bufg or posedge rst_tmp_phaser_ref)
    if (rst_tmp_phaser_ref)
      rst_phaser_ref_sync_r <= #TCQ {RST_DIV_SYNC_NUM{1'b1}};
    else
      rst_phaser_ref_sync_r <= #TCQ rst_phaser_ref_sync_r << 1;
  assign rst_phaser_ref = rst_phaser_ref_sync_r[RST_DIV_SYNC_NUM-1];
endmodule