module sky130_fd_sc_hs__dlxtp (
    //# {{data|Data Signals}}
    input  D   ,
    output Q   ,
    //# {{clocks|Clocking}}
    input  GATE
);
    // Voltage supply signals
    supply1 VPWR;
    supply0 VGND;
endmodule