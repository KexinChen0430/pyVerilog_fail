module ne576ee
   (
    sys_clk,
    rst_n,
    fnddca9,
    ho79420,
    cm72a72,
    qv95390,
    ksa9c85,
    mtb4ec3,
    yk78c4c,
    shc6261,
    yz8514c,
    nt28a64,
    xj45326,
    ep29936,
    ay4c9b4,
    ld64da1,
    cb26d0e,
    mt36875,
    sjb43ac,
    oha1d64,
    bn2d5a3,
    ip6ad1f,
    mgac915,
    pf648a8,
    ohd0c6,
    me68634,
    qgef2ad,
    ep18d09,
    uvc684c,
    zx55a12,
    qg431a1,
    fa7944d,
    rgca26a,
    qt51353,
    ls89a9d,
    tu4d4eb,
    cz6a75a,
    tj9905,
    ec34264,
    zkeb509,
    gda1320,
    god4257,
    ba20bcf,
    bn22886,
    qvb47e9,
    rge1dc0,
    gbf8072,
    vka761d,
    rt64179,
    ea4c82f,
    th61a18,
    fp91fdb,
    yz8fede
    );
`ifdef LW1
parameter LANE_WIDTH = 1 ;
`else
`ifdef LW2
parameter LANE_WIDTH = 2 ;
`else
`ifdef LW4
parameter LANE_WIDTH = 4 ;
`else
parameter LANE_WIDTH = 1 ;
`endif
`endif
`endif
parameter D_WIDTH = 16 ;
parameter K27_7 = 8'hFB ;
parameter K28_0 = 8'h1C ;
parameter K28_2 = 8'h5C ;
parameter K28_3 = 8'h7C ;
parameter K28_5 = 8'hBC ;
parameter K29_7 = 8'hFD ;
parameter K30_7 = 8'hFE ;
parameter K23_7 = 8'hF7 ;
parameter K28_1 = 8'h3C ;
parameter D5_2  = 8'h45 ;
parameter D10_2 = 8'h4A ;
parameter D21_5 = 8'hB5 ;
parameter D26_5 = 8'hBA ;
parameter COM = K28_5 ;
parameter STP = K27_7 ;
parameter SDP = K28_2 ;
parameter END = K29_7 ;
parameter EDB = K30_7 ;
parameter SKP = K28_0 ;
parameter IDL = K28_3 ;
parameter PAD = K23_7 ;
parameter FTS = K28_1 ;
parameter OS_WIDTH      = 4 ;
parameter OS_T1_LIP_LAP = 4'd0 ;
parameter OS_T2_LIP_LAP = 4'd1 ;
parameter OS_COMPLI     = 4'd2 ;
parameter OS_T1         = 4'd3 ;
parameter OS_T2         = 4'd4 ;
parameter OS_IDLE       = 4'd5 ;
parameter OS_EIDLE      = 4'd6 ;
parameter OS_NFTS       = 4'd7 ;
parameter OS_BEACON     = 4'd8 ;
parameter DSM_WIDTH    = 2 ;
parameter PSM_WIDTH    = 2 ;
parameter RSM_WIDTH    = 2 ;
parameter L0SM_WIDTH   = 2 ;
parameter L0sTSM_WIDTH = 2 ;
parameter L0sRSM_WIDTH = 2 ;
parameter L1SM_WIDTH   = 1 ;
parameter L2SM_WIDTH   = 1 ;
parameter DISM_WIDTH   = 2 ;
parameter LBSM_WIDTH   = 2 ;
parameter HRSM_WIDTH   = 1 ;
parameter CFGSM_WIDTH  = 2 ;
parameter MSM_WIDTH    = 3 ;
parameter DETECT    = 4'd0 ;
parameter POLLING   = 4'd1 ;
parameter CONFIG    = 4'd2 ;
parameter L0        = 4'd3 ;
parameter L0s       = 4'd4 ;
parameter L1        = 4'd5 ;
parameter L2        = 4'd6 ;
parameter RECOVERY  = 4'd7 ;
parameter LOOPBACK  = 4'd8 ;
parameter HOTRST    = 4'd9 ;
parameter DISABLED  = 4'd10 ;
`ifdef VC1
parameter FADDR = 3 ;
`else
`ifdef VC2
parameter FADDR = 3 ;
`else
`ifdef VC3
parameter FADDR = 5 ;
`else
`ifdef VC4
parameter FADDR = 5 ;
`else
parameter FADDR = 6 ;
`endif
`endif
`endif
`endif
input                     sys_clk;
input                     rst_n;
input                     fnddca9;
input                     ho79420;
input                     cm72a72;
input   [15:0]            qv95390;
input   [1:0]             ksa9c85;
input                     mtb4ec3;
input                     yk78c4c;
input                     shc6261;
input                     nt28a64;
input                     yz8514c;
input   [7:0]             xj45326;
input                     ep29936;
input                     ay4c9b4;
input                     ld64da1;
input   [7:0]             cb26d0e;
input   [7:0]             mt36875;
output                    sjb43ac;
output  [7:0]             oha1d64;
output                    bn2d5a3;
output                    ip6ad1f;
output                    mgac915;
output                    pf648a8;
output                    ohd0c6;
output                    me68634;
output                    qgef2ad;
output                    ep18d09;
output                    uvc684c;
output                    zx55a12;
output                    qg431a1;
output                    fa7944d;
output                    tj9905;
output                    ec34264;
output                    tu4d4eb;
output                    cz6a75a;
output                    rgca26a;
output                    qt51353;
output                    ls89a9d;
output                    zkeb509;
output                    gda1320;
output                    god4257;
output                    ba20bcf;
output                    bn22886;
output                    qvb47e9;
output                    rge1dc0;
output                    gbf8072;
output                    vka761d;
output                    rt64179;
output                    ea4c82f;
output                    th61a18;
output                    fp91fdb;
output  [7:0]             yz8fede;
reg                      bn2d5a3;
reg                      ip6ad1f;
reg                      mgac915;
reg                      pf648a8;
reg                      jcd0a1a;
reg                      ep850d2;
reg                      jr28694;
reg                      su434a7;
reg                      sw1a539;
reg                      dzd29c8;
reg                      nt94e47;
reg                      jea723e;
reg                      mt391f2;
reg                      xjc8f94;
reg                      lq47ca7;
reg                      ks3e53a;
reg                      kdf29d1;
reg                      db94e8c;
reg                      hqa7466;
reg                      vk3a332;
reg                      sud1993;
reg                      god4257;
reg                      lq664c3;
reg                      bn22886;
reg                      qvb47e9;
reg                      rge1dc0;
reg                      qtc35d1;
reg                      co1ae8d;
reg                      jpd7469;
reg                      fpba34e;
reg                      uid1a77;
reg                      mg8d3b8;
reg  [7:0]               yz8fede;
reg  [15:0]              yx4ee02;
reg  [15:0]              os77014;
reg  [15:0]              lsb80a1;
reg  [1:0]               nec050a;
reg  [1:0]               cb2852;
reg  [1:0]               ri14294;
reg                      uxa14a3;
reg                      yma51d;
reg                      tu528e9;
reg                      lf9474b;
reg                      wya3a5f;
reg                      qv1d2f9;
reg   [2:0]              rte97cd;
reg   [1:0]              gb4be6f;
reg   [3:0]              dz5f37c;
reg   [1:0]              nrf9be6;
reg   [1:0]              jpcdf37;
reg   [1:0]              en6f9bf;
reg   [1:0]              fa7cdfd;
reg   [3:0]              xje6feb;
reg   [3:0]              zz37f5f;
reg   [1:0]              tjbfafe;
reg   [3:0]              alfd7f6;
reg   [3:0]              dmebfb4;
reg   [1:0]              zx5fda3;
reg   [3:0]              jcfed1f;
reg   [3:0]              zxf68fa;
reg   [1:0]              sjb47d6;
reg   [1:0]              mga3eb4;
reg   [1:0]              mg1f5a1;
reg   [1:0]              eafad08;
reg   [1:0]              kdd6840;
reg   [3:0]              qvb4205;
reg                      yza102c;
reg                      sjb43ac;
reg                      dz40b2c;
wire                     co5967;
wire                     wl2cb39;
wire                     qt659cc;
wire  [7:0]              qv2ce64;
wire  [7:0]              su67324;
wire  [7:0]              gd39920;
wire  [7:0]              encc905;
wire                     rt6482d;
wire                     wy2416e;
wire                     pu20b71 ;
wire                     gq5b8a ;
wire                     db2dc51 ;
wire                     vv6e28e;
wire                     jp71476;
`ifdef GEN2
`else
`endif
`ifdef GEN2
reg ux8a3b6 ;
`else
`endif
reg of51db5;
reg qt54e55;
reg by76d66;
reg [15 : 0] gqb6b32;
reg [1 : 0] xlb5990;
reg nt28480;
reg osffa9c;
reg uiea704;
reg mt90e17;
reg aa870bc;
reg [7 : 0] hd385e1;
reg jpc2f0e;
reg wl17876;
reg gqbc3b5;
reg [7 : 0] zke1da8;
reg [7 : 0] jeed42;
reg zk76a12;
reg tjb5092;
reg vka8496;
reg lq424b3;
reg qv1259b;
reg gq92cdc;
reg je966e1;
reg cob370a;
reg vx9b851;
reg endc28f;
reg xwe147d;
reg wya3eb;
reg en51f59;
reg qv8facc;
reg cm7d664;
reg tueb320;
reg qg59902;
reg mrcc810;
reg dz64085;
reg tw2042f;
reg sj217b;
reg sw10bdd;
reg yz85ee8;
reg pu2f745;
reg [15 : 0] nr7ba2a;
reg [15 : 0] fndd156;
reg [15 : 0] gbe8ab7;
reg [1 : 0] th455bc;
reg [1 : 0] xy2ade6;
reg [1 : 0] ay56f33;
reg ngb7999;
reg ymbccca;
reg the6651;
reg oh3328e;
reg ls99475;
reg byca3ab;
reg [2 : 0] sh51d5b;
reg [1 : 0] zz8eadc;
reg [3 : 0] yx756e6;
reg [1 : 0] kfab734;
reg [1 : 0] yx5b9a4;
reg [1 : 0] czdcd25;
reg [1 : 0] fne692c;
reg [3 : 0] ie34967;
reg [3 : 0] qva4b39;
reg [1 : 0] pu259cc;
reg [3 : 0] ir2ce62;
reg [3 : 0] go67314;
reg [1 : 0] oh398a0;
reg [3 : 0] qtcc505;
reg [3 : 0] cm6282c;
reg [1 : 0] ls14161;
reg [1 : 0] zza0b0b;
reg [1 : 0] ie585e;
reg [1 : 0] sj2c2f1;
reg [1 : 0] pf6178d;
reg [3 : 0] lsbc6f;
reg qt5e37a;
reg lqf1bd4;
reg mg8dea3;
reg cz6f519;
reg mr7a8cc;
reg [7 : 0] uid4664;
reg [7 : 0] qia3321;
reg [7 : 0] rv19908;
reg [7 : 0] uvcc846;
reg pf64235;
reg ks211af;
reg yz8d79;
reg su46bcd;
reg pu35e68;
reg vxaf343;
reg ho79a1e;
reg [2047:0] necf6c2;
wire [88:0] ld7b613;
`ifdef LW1
`else
`ifdef LW2
`else
`ifdef LW4
`else
`endif
`endif
`endif
`ifdef VC1
`else
`ifdef VC2
`else
`ifdef VC3
`else
`ifdef VC4
`else
`endif
`endif
`endif
`endif
`ifdef GEN2
`else
`endif
`ifdef GEN2
`else
`endif
localparam qgdb09f = 89,nrd84f8 = 32'hfdfff10b;
localparam [31:0] thc27c7 = nrd84f8;
localparam mt9f1ff = nrd84f8 & 4'hf;
localparam [11:0] fnc7fe5 = 'h7ff;
wire  [(1 << mt9f1ff)  -1:0] suff972;
reg    [qgdb09f-1:0] cme5c87;
reg [mt9f1ff-1:0] qg721c0 [0:1];
reg [mt9f1ff-1:0] ym8700c;
reg rv38061;
integer jcc030e;
integer vk1872;
`ifdef LW1
`else
`ifdef LW2
`else
`ifdef LW4
`else
`endif
`endif
`endif
`ifdef VC1
`else
`ifdef VC2
`else
`ifdef VC3
`else
`ifdef VC4
`else
`endif
`endif
`endif
`endif
`ifdef GEN2
`else
`endif
`ifdef GEN2
`else
`endif
`ifdef LW1
`else
`ifdef LW2
`else
`ifdef LW4
`else
`endif
`endif
`endif
`ifdef VC1
`else
`ifdef VC2
`else
`ifdef VC3
`else
`ifdef VC4
`else
`endif
`endif
`endif
`endif
always @(posedge sys_clk or negedge rst_n) begin   if (!rst_n) begin      yx4ee02 <= 0;      os77014 <= 0;      lsb80a1 <= 0;
      nec050a  <= 0;      cb2852  <= 0;      ri14294  <= 0;      uxa14a3 <= 0;      yma51d <= 0;      tu528e9 <= 0;   end   else begin                  yx4ee02 <= (by76d66) ? gqb6b32 : 15'hFF;      os77014 <= nr7ba2a;      lsb80a1 <= fndd156;      nec050a  <= (by76d66) ? xlb5990 : 0;      cb2852  <= th455bc;      ri14294  <= xy2ade6;            uxa14a3 <= qt54e55;      yma51d <= ngb7999;      tu528e9 <= ymbccca;   end
end
ir1d094 ene84a5 (        .sys_clk          ( sys_clk ),    .rst_n            ( rst_n ),
    .xl2d776           ( nr7ba2a ),    .xw5ddbf            ( th455bc ),
        .ps76fd3        ( co5967 ),    .rvbf4d2        ( wl2cb39 ),    .ald34b9      ( qt659cc ),    .rtd2e64        ( qv2ce64 ),    .wyb9938  ( rt6482d ),    .bl64e0d        ( su67324 ),    .bn38376  ( wy2416e ),    .irddb1        ( gd39920 ),    .by76c6f        ( encc905 )   ) ;
assign oha1d64 = uid4664;
always @(posedge sys_clk or negedge rst_n) begin   if (!rst_n) begin      lf9474b <= 1'b0;   end   else begin      lf9474b <= (((gbe8ab7[7:0] == K28_5) & (ay56f33[0] == 1'b1) &               (fndd156 == {IDL, IDL}) & (xy2ade6[1:0] == 2'b11)) |                      ((gbe8ab7[15:8] == K28_5) & (ay56f33[1] == 1'b1) &       ({gbe8ab7[7:0], fndd156[15:8]} == {IDL, IDL}) & ay56f33[0] & xy2ade6[1])             );   end
end
always @(posedge sys_clk or negedge rst_n) begin   if (!rst_n) begin      wya3a5f  <= 1'b0;   end   else  begin      wya3a5f <= (((fndd156 == {K28_5, SKP}) & (xy2ade6[1:0] == 2'b11)) |                    (({gbe8ab7[7:0],fndd156[15:8]}  == {K28_5, SKP}) & ay56f33[0] & xy2ade6[1]));   end
end
always @(posedge sys_clk or negedge rst_n) begin   if (!rst_n) begin      qv1d2f9  <= 1'b0;   end   else begin      qv1d2f9 <= ((({gbe8ab7, fndd156}  == {K28_5, FTS, FTS, FTS}) &                     ({ay56f33, xy2ade6} == 4'b1111)) |                    (({gbe8ab7[7:0], fndd156, nr7ba2a[15:8] }  == {K28_5, FTS, FTS, FTS}) &                     ({ay56f33[0], xy2ade6, th455bc[1]} == 4'b1111)));   end
end
always @(posedge sys_clk or negedge rst_n) begin   if (!rst_n) begin      yza102c <= 1'b0;   end   else begin      yza102c <= oh3328e || byca3ab;   end
end
assign pu20b71      = ((fndd156[7:0]  ==  8'h00) && (xy2ade6[0] == 1'b0)) ;
assign gq5b8a      = ((fndd156[15:8] ==  8'h00) && (xy2ade6[1] == 1'b0)) ;
assign db2dc51 = ((gbe8ab7[7:0]  ==  8'h00) && (ay56f33[0] == 1'b0)) ;
always @(posedge sys_clk or negedge rst_n) begin   if (!rst_n) begin      qvb4205 <= 0;   end   else begin      if (aa870bc) begin         qvb4205 <= 0;      end                  else if (((lsbc6f < 'd8) && ~of51db5) ||               ((lsbc6f < 'd3) &&  of51db5)) begin         case({su46bcd,yz8d79})            2'b00: qvb4205 <= 0;            2'b01: qvb4205 <= 4'd1;            2'b11: qvb4205 <= (pu35e68) ? (lsbc6f +4'd2) : 4'd2;            2'b10: qvb4205 <= (pu35e68) ? (lsbc6f +4'd1) : 0;         endcase      end   end
end
assign  vv6e28e  = (pf64235 == 1'b0) & (uid4664 == zke1da8);
assign  jp71476  = (ks211af == 1'b0) & (qia3321 == jeed42);
always @(posedge sys_clk or negedge rst_n) begin   if (!rst_n) begin      gb4be6f   <= 0;      dz5f37c  <= 0;      nrf9be6   <= 0;      jpcdf37    <= 0;      en6f9bf      <= 0;      fa7cdfd    <= 0;      xje6feb  <= 0;      zz37f5f  <= 0;      tjbfafe   <= 0;      alfd7f6  <= 0;      dmebfb4 <= 0;      zx5fda3          <= 0;      jcfed1f   <= 0;      zxf68fa   <= 0;      sjb47d6     <= 0;      mga3eb4      <= 0;      mg1f5a1      <= 0;      eafad08     <= 0;      kdd6840     <= 0;      rte97cd         <= 0;   end   else begin            if (qt5e37a | aa870bc) begin         gb4be6f <= 0;      end            else if (!zz8eadc[1]) begin         if (mg8dea3 && {uid4664,qia3321}== {PAD,PAD} && {pf64235,ks211af} == 2'b11) begin            gb4be6f <= zz8eadc + 1;         end         else if (mg8dea3 || cz6f519) begin            gb4be6f <= 0;         end      end            if (qt5e37a | aa870bc) begin         dz5f37c <= 0;      end      else if (!yx756e6[3]) begin
`ifdef GEN2
            if (({uid4664,qia3321}== {PAD,PAD}) &&        ({pf64235,ks211af} == 2'b11) &&        ((uvcc846[4] == 1'b0 && mg8dea3) ||                 (uvcc846[2] == 1'b1 && mg8dea3) ||                 (cz6f519)        )       ) begin               dz5f37c <= yx756e6 + 1;            end
`else
            if ((mg8dea3 || cz6f519) && {uid4664,qia3321}== {PAD,PAD} && {pf64235,ks211af} == 2'b11) begin               dz5f37c <= yx756e6 + 1;            end
`endif
         else if (mg8dea3 || cz6f519) begin            dz5f37c <= 0;         end      end            if (qt5e37a | aa870bc) begin         nrf9be6 <= 0;      end            else if (!kfab734[1]) begin         if (mg8dea3 && {uid4664,qia3321}== {zke1da8,PAD} && {pf64235,ks211af} == 2'b01) begin            nrf9be6 <= kfab734 + 1;         end         else if (mg8dea3 || cz6f519) begin            nrf9be6 <= 0;         end      end
             if (qt5e37a | aa870bc) begin         jpcdf37 <= 0;      end            else if (!yx5b9a4[1]) begin         if (mg8dea3 && {qia3321}== {PAD} && {pf64235,ks211af} == 2'b01) begin            jpcdf37 <= yx5b9a4 + 1;         end         else if (mg8dea3 || cz6f519) begin            jpcdf37 <= 0;         end      end             if (qt5e37a | aa870bc) begin         en6f9bf <= 0;      end            else if (!czdcd25[1]) begin         if (mg8dea3 && {qia3321}== {PAD} && ks211af == 1'b1) begin            en6f9bf <= czdcd25 + 1;         end         else if (mg8dea3 || cz6f519) begin            en6f9bf <= 0;         end      end            if (qt5e37a | aa870bc) begin         fa7cdfd <= 0;      end            else if (!fne692c[1]) begin         if (mg8dea3 && {uid4664}== {zke1da8} && {pf64235,ks211af} == 2'b00) begin            fa7cdfd <= fne692c + 1;         end         else if (mg8dea3 || cz6f519) begin            fa7cdfd <= 0;         end      end            if (qt5e37a | aa870bc) begin         xje6feb <= 0;      end            else if (!ie34967[3]) begin                  if (mg8dea3 && vxaf343 && !ho79a1e) begin            xje6feb <= ie34967 + 1;         end         else if (mg8dea3 || cz6f519) begin            xje6feb <= 0;         end      end             if (qt5e37a | aa870bc) begin         zz37f5f <= 0;      end            else if (!qva4b39[3]) begin                  if (mg8dea3 && !vxaf343 && ho79a1e) begin            zz37f5f <= qva4b39 + 1;         end         else if (mg8dea3 || cz6f519) begin            zz37f5f <= 0;         end      end
            if (qt5e37a | aa870bc) begin         tjbfafe <= 0;      end            else if (!pu259cc[1]) begin         if (mg8dea3 && {uid4664,qia3321}== {zke1da8,jeed42} && {pf64235,ks211af} == 2'b00) begin            tjbfafe <= pu259cc + 1;         end         else if (mg8dea3 || cz6f519) begin            tjbfafe <= 0;         end      end
            if (qt5e37a | aa870bc) begin         alfd7f6 <= 0;      end            else if (!ir2ce62[3]) begin         if ((mg8dea3 || cz6f519) && {uid4664,qia3321}== {zke1da8,jeed42} && {pf64235,ks211af} == 2'b00) begin            alfd7f6 <= ir2ce62 + 1;         end         else if (mg8dea3 || cz6f519) begin            alfd7f6 <= 0;         end      end             if (qt5e37a | aa870bc) begin         dmebfb4 <= 0;      end            else if (!go67314[3]) begin                  if (mg8dea3 && !vxaf343 && !ho79a1e) begin            dmebfb4 <= go67314 + 1;         end         else if (mg8dea3 || cz6f519) begin            dmebfb4 <= 0;         end      end             if (qt5e37a | aa870bc) begin         rte97cd <= 0;      end            else if (!sh51d5b[2]) begin         if (mg8dea3 || cz6f519) begin            rte97cd <= sh51d5b + 1;         end      end
            if (qt5e37a | aa870bc) begin         zx5fda3 <= 0;      end            else if (!oh398a0[1]) begin         if (cz6f519) begin            zx5fda3 <= oh398a0 + 1;         end         else if (mg8dea3) begin            zx5fda3 <= 0;         end      end            if (qt5e37a | aa870bc) begin         jcfed1f <= 0;      end            else if (!qtcc505[3]) begin         if (cz6f519 && {uid4664,qia3321}== {PAD,PAD} && {pf64235,ks211af} == 2'b11) begin            jcfed1f <= qtcc505 + 1;         end         else if (mg8dea3 || cz6f519) begin            jcfed1f <= 0;         end      end
            if (qt5e37a | aa870bc) begin         zxf68fa <= 0;      end            else if (!cm6282c[3]) begin         if (cz6f519 && {uid4664,qia3321}== {zke1da8,jeed42} && {pf64235,ks211af} == 2'b00) begin            zxf68fa <= cm6282c + 1;         end         else if (mg8dea3 || cz6f519) begin            zxf68fa <= 0;         end      end            if (qt5e37a | aa870bc) begin         sjb47d6 <= 0;      end            else if (!ls14161[1]) begin         if (mg8dea3 && uvcc846[0] == 1'b1 && vxaf343 && ho79a1e) begin            sjb47d6 <= ls14161 + 1;         end         else if (mg8dea3 || cz6f519) begin            sjb47d6 <= 0;         end      end            if (qt5e37a | aa870bc) begin         mga3eb4 <= 0;      end            else if (!zza0b0b[1]) begin         if (mg8dea3 && uvcc846[1] == 1'b1) begin            mga3eb4 <= zza0b0b + 1;         end         else if (mg8dea3 || cz6f519) begin            mga3eb4 <= 0;         end      end
             if (qt5e37a | aa870bc) begin         mg1f5a1 <= 0;      end            else if (!ie585e[1]) begin         if (mg8dea3 && uvcc846[2] == 1'b1) begin            mg1f5a1 <= ie585e + 1;         end         else if (mg8dea3 || cz6f519) begin            mg1f5a1 <= 0;         end      end             if (qt5e37a | aa870bc) begin         eafad08 <= 0;      end            else if (!sj2c2f1[1]) begin         if (mg8dea3 && uvcc846[2] == 1'b1 && {uid4664,qia3321} == {zke1da8,jeed42} &&            {pf64235,ks211af} == 2'b00 && rv19908 == hd385e1 ) begin            eafad08 <= sj2c2f1 + 1;         end         else if (mg8dea3 || cz6f519) begin            eafad08 <= 0;         end      end
             if (qt5e37a | aa870bc) begin         kdd6840 <= 0;      end            else if (!pf6178d[1]) begin         if (cz6f519 && uvcc846[3] == 1'b1) begin            kdd6840 <= pf6178d + 1;         end         else if (mg8dea3 || cz6f519) begin            kdd6840 <= 0;         end      end   end
end
always @(posedge sys_clk or negedge rst_n) begin   if (!rst_n) begin      mgac915    <= 1'b0;      pf648a8    <= 1'b0;      bn2d5a3           <= 1'b0;      ip6ad1f           <= 1'b0;      god4257         <= 1'b0;      bn22886        <= 1'b0;      rge1dc0          <= 1'b0;      yz8fede         <= 0;   end   else begin
      if (mg8dea3 && {uid4664,qia3321}== {zke1da8,jeed42} && {pf64235,ks211af}== 2'b00)         mgac915 <= 1'b1;      else         mgac915 <= 1'b0;      if (cz6f519 && {uid4664,qia3321}== {zke1da8,jeed42} && {pf64235,ks211af}== 2'b00)         pf648a8 <= 1'b1;      else         pf648a8 <= 1'b0;      bn2d5a3           <= mg8dea3;      ip6ad1f           <= cz6f519;      if (of51db5)      god4257         <= (lsbc6f >= 4'd3) ? 1'b1 : 1'b0;      else      god4257         <= (lsbc6f >= 4'd4) ? 1'b1 : 1'b0;
      bn22886        <= oh3328e;      rge1dc0          <= ls99475;      yz8fede         <= rv19908;   end
end
`ifdef GEN2
   always @(posedge sys_clk or negedge rst_n) begin      if (!rst_n)         ux8a3b6 <= 1'b0;      else if (ls99475)         ux8a3b6 <= 1'b1;      else if (gqbc3b5)         ux8a3b6  <= 1'b0;   end   always @(posedge sys_clk or negedge rst_n) begin      if (!rst_n)         qvb47e9 <= 1'b0;      else         qvb47e9 <= ((~the6651 & ymbccca & ~oh3328e) |                             (gqbc3b5 && ~ux8a3b6)) ? 1'b1 : 1'b0;   end
`else
   always @(posedge sys_clk or negedge rst_n) begin      if (!rst_n) begin         qvb47e9 <= 1'b0;      end      else begin         qvb47e9 <= (~the6651 & ymbccca & ~oh3328e) ? 1'b1 : 1'b0;      end   end
`endif
always @(posedge sys_clk or negedge rst_n) begin   if (!rst_n) begin      jcd0a1a         <= 1'b0;      ep850d2   <= 1'b0;      jr28694   <= 1'b0;      su434a7    <= 1'b0;      sw1a539  <= 1'b0;      dzd29c8   <= 1'b0;      nt94e47    <= 1'b0;      jea723e      <= 1'b0;      kdf29d1 <= 1'b0;      db94e8c  <= 1'b0;      hqa7466  <= 1'b0;      lq47ca7  <= 1'b0;      ks3e53a  <= 1'b0;      mt391f2          <= 1'b0;      xjc8f94   <= 1'b0;      vk3a332   <= 1'b0;      sud1993   <= 1'b0;      lq664c3        <= 1'b0;      qtc35d1      <= 1'b0;      co1ae8d     <= 1'b0;      jpd7469     <= 1'b0;      fpba34e      <= 1'b0;      uid1a77      <= 1'b0;      mg8d3b8     <= 1'b0;   end   else if (aa870bc) begin      jcd0a1a         <= 1'b0;      ep850d2   <= 1'b0;      jr28694   <= 1'b0;      su434a7    <= 1'b0;      sw1a539  <= 1'b0;      dzd29c8   <= 1'b0;      nt94e47    <= 1'b0;      jea723e      <= 1'b0;      kdf29d1 <= 1'b0;      db94e8c  <= 1'b0;      hqa7466  <= 1'b0;      lq47ca7  <= 1'b0;      ks3e53a  <= 1'b0;      mt391f2          <= 1'b0;      xjc8f94   <= 1'b0;      vk3a332   <= 1'b0;      sud1993   <= 1'b0;      lq664c3        <= 1'b0;      qtc35d1      <= 1'b0;      co1ae8d     <= 1'b0;      jpd7469     <= 1'b0;      fpba34e      <= 1'b0;      uid1a77      <= 1'b0;      mg8d3b8     <= 1'b0;   end   else begin      jcd0a1a         <= sh51d5b[2];                           ep850d2   <= zz8eadc[1];                     lq47ca7  <= yx756e6[3];                    jr28694   <= kfab734[1];                     su434a7    <= fne692c[1];                      sw1a539  <= (|ie34967[3:1]);               dzd29c8   <= pu259cc[1];                     ks3e53a  <= ir2ce62[3];                    nt94e47    <= yx5b9a4[1];                      jea723e      <= czdcd25[1];                        kdf29d1 <= go67314[3];                   db94e8c  <= qva4b39[3];                    hqa7466  <= ie34967[3];                    mt391f2          <= oh398a0[1];                            xjc8f94   <= (|cm6282c[3:1]);                vk3a332   <= qtcc505[3];                     sud1993   <= cm6282c[3];                     if (of51db5)      lq664c3        <= lsbc6f >= 'd3;                      else      lq664c3        <= lsbc6f[3];                          qtc35d1      <= sj2c2f1[1];                       co1ae8d     <= ls14161[1];                       jpd7469     <= pf6178d[1];                       fpba34e      <= (ie585e[1] || uiea704);        uid1a77      <= (zza0b0b[1] || osffa9c);        mg8d3b8     <= (ls14161[1]|| nt28480);    end
end
assign  ohd0c6         = zk76a12;
assign  me68634   = tjb5092;
assign  qgef2ad   = vka8496;
assign  ep18d09    = lq424b3;
assign  uvc684c  = qv1259b;
assign  zx55a12   = gq92cdc;
assign  qg431a1    = je966e1;
assign  fa7944d      = cob370a;
assign  rgca26a = en51f59;
assign  qt51353  = qv8facc;
assign  ls89a9d  = cm7d664;
assign  tu4d4eb  = xwe147d;
assign  cz6a75a  = wya3eb;
assign  tj9905          = vx9b851;
assign  ec34264   = endc28f;
assign  zkeb509   = tueb320;
assign  gda1320   = qg59902;
assign  ba20bcf        = mrcc810;
assign  gbf8072      = dz64085;
assign  vka761d     = tw2042f;
assign  rt64179     = sj217b;
assign  ea4c82f      = sw10bdd;
assign  th61a18      = yz85ee8;
assign  fp91fdb     = pu2f745;
always @(posedge sys_clk or negedge rst_n) begin   if (!rst_n) begin      dz40b2c     <= 1'b0;      sjb43ac      <= 1'b0;   end   else begin                  if (jpc2f0e == 1'b0) begin         dz40b2c <= 1'b0;      end      else if (mr7a8cc) begin         dz40b2c <= 1'b1;      end                  if (wl17876 == 1'b1) begin         sjb43ac <= 1'b0 ;      end      else if (mt90e17) begin         sjb43ac <= lqf1bd4;      end   end
end
always@* begin of51db5<=ld7b613[0];qt54e55<=ld7b613[1];by76d66<=ld7b613[2];gqb6b32<={qv95390>>1,ld7b613[3]};xlb5990<={ksa9c85>>1,ld7b613[4]};nt28480<=ld7b613[5];osffa9c<=ld7b613[6];uiea704<=ld7b613[7];mt90e17<=ld7b613[8];aa870bc<=ld7b613[9];hd385e1<={xj45326>>1,ld7b613[10]};jpc2f0e<=ld7b613[11];wl17876<=ld7b613[12];gqbc3b5<=ld7b613[13];zke1da8<={cb26d0e>>1,ld7b613[14]};jeed42<={mt36875>>1,ld7b613[15]};zk76a12<=ld7b613[16];tjb5092<=ld7b613[17];vka8496<=ld7b613[18];lq424b3<=ld7b613[19];qv1259b<=ld7b613[20];gq92cdc<=ld7b613[21];je966e1<=ld7b613[22];cob370a<=ld7b613[23];vx9b851<=ld7b613[24];endc28f<=ld7b613[25];xwe147d<=ld7b613[26];wya3eb<=ld7b613[27];en51f59<=ld7b613[28];qv8facc<=ld7b613[29];cm7d664<=ld7b613[30];tueb320<=ld7b613[31];qg59902<=ld7b613[32];mrcc810<=ld7b613[33];dz64085<=ld7b613[34];tw2042f<=ld7b613[35];sj217b<=ld7b613[36];sw10bdd<=ld7b613[37];yz85ee8<=ld7b613[38];pu2f745<=ld7b613[39];nr7ba2a<={yx4ee02>>1,ld7b613[40]};fndd156<={os77014>>1,ld7b613[41]};gbe8ab7<={lsb80a1>>1,ld7b613[42]};th455bc<={nec050a>>1,ld7b613[43]};xy2ade6<={cb2852>>1,ld7b613[44]};ay56f33<={ri14294>>1,ld7b613[45]};ngb7999<=ld7b613[46];ymbccca<=ld7b613[47];the6651<=ld7b613[48];oh3328e<=ld7b613[49];ls99475<=ld7b613[50];byca3ab<=ld7b613[51];sh51d5b<={rte97cd>>1,ld7b613[52]};zz8eadc<={gb4be6f>>1,ld7b613[53]};yx756e6<={dz5f37c>>1,ld7b613[54]};kfab734<={nrf9be6>>1,ld7b613[55]};yx5b9a4<={jpcdf37>>1,ld7b613[56]};czdcd25<={en6f9bf>>1,ld7b613[57]};fne692c<={fa7cdfd>>1,ld7b613[58]};ie34967<={xje6feb>>1,ld7b613[59]};qva4b39<={zz37f5f>>1,ld7b613[60]};pu259cc<={tjbfafe>>1,ld7b613[61]};ir2ce62<={alfd7f6>>1,ld7b613[62]};go67314<={dmebfb4>>1,ld7b613[63]};oh398a0<={zx5fda3>>1,ld7b613[64]};qtcc505<={jcfed1f>>1,ld7b613[65]};cm6282c<={zxf68fa>>1,ld7b613[66]};ls14161<={sjb47d6>>1,ld7b613[67]};zza0b0b<={mga3eb4>>1,ld7b613[68]};ie585e<={mg1f5a1>>1,ld7b613[69]};sj2c2f1<={eafad08>>1,ld7b613[70]};pf6178d<={kdd6840>>1,ld7b613[71]};lsbc6f<={qvb4205>>1,ld7b613[72]};qt5e37a<=ld7b613[73];lqf1bd4<=ld7b613[74];mg8dea3<=ld7b613[75];cz6f519<=ld7b613[76];mr7a8cc<=ld7b613[77];uid4664<={qv2ce64>>1,ld7b613[78]};qia3321<={su67324>>1,ld7b613[79]};rv19908<={gd39920>>1,ld7b613[80]};uvcc846<={encc905>>1,ld7b613[81]};pf64235<=ld7b613[82];ks211af<=ld7b613[83];yz8d79<=ld7b613[84];su46bcd<=ld7b613[85];pu35e68<=ld7b613[86];vxaf343<=ld7b613[87];ho79a1e<=ld7b613[88];end
always@* begin necf6c2[2047]<=ho79420;necf6c2[2046]<=cm72a72;necf6c2[2044]<=qv95390[0];necf6c2[2040]<=ksa9c85[0];necf6c2[2032]<=mtb4ec3;necf6c2[2016]<=yk78c4c;necf6c2[1985]<=shc6261;necf6c2[1950]<=ep850d2;necf6c2[1930]<=jea723e;necf6c2[1923]<=yz8514c;necf6c2[1909]<=wy2416e;necf6c2[1878]<=jpcdf37[0];necf6c2[1874]<=vv6e28e;necf6c2[1870]<=wl2cb39;necf6c2[1852]<=jr28694;necf6c2[1813]<=mt391f2;necf6c2[1799]<=nt28a64;necf6c2[1770]<=pu20b71;necf6c2[1708]<=en6f9bf[0];necf6c2[1700]<=jp71476;necf6c2[1693]<=qt659cc;necf6c2[1656]<=su434a7;necf6c2[1578]<=xjc8f94;necf6c2[1573]<=zx5fda3[0];necf6c2[1551]<=xj45326[0];necf6c2[1493]<=dz5f37c[0];necf6c2[1492]<=gq5b8a;necf6c2[1491]<=dz40b2c;necf6c2[1417]<=alfd7f6[0];necf6c2[1396]<=qvb4205[0];necf6c2[1378]<=zz37f5f[0];necf6c2[1368]<=fa7cdfd[0];necf6c2[1353]<=yx4ee02[0];necf6c2[1345]<=hqa7466;necf6c2[1339]<=qv2ce64[0];necf6c2[1316]<=lsb80a1[0];necf6c2[1285]<=sud1993;necf6c2[1265]<=sw1a539;necf6c2[1262]<=gd39920[0];necf6c2[1198]<=mg1f5a1[0];necf6c2[1169]<=cb2852[0];necf6c2[1163]<=yma51d;necf6c2[1117]<=wya3a5f;necf6c2[1108]<=lq47ca7;necf6c2[1098]<=jcfed1f[0];necf6c2[1054]<=ep29936;necf6c2[1045]<=qtc35d1;necf6c2[1023]<=fnddca9;necf6c2[975]<=jcd0a1a;necf6c2[965]<=nt94e47;necf6c2[954]<=rt6482d;necf6c2[939]<=nrf9be6[0];necf6c2[937]<=db2dc51;necf6c2[935]<=co5967;necf6c2[786]<=dmebfb4[0];necf6c2[746]<=gb4be6f[0];necf6c2[745]<=yza102c;necf6c2[708]<=tjbfafe[0];necf6c2[698]<=kdd6840[0];necf6c2[689]<=xje6feb[0];necf6c2[676]<=mg8d3b8;necf6c2[672]<=db94e8c;necf6c2[658]<=os77014[0];necf6c2[642]<=vk3a332;necf6c2[631]<=su67324[0];necf6c2[599]<=mga3eb4[0];necf6c2[584]<=nec050a[0];necf6c2[581]<=uxa14a3;necf6c2[558]<=lf9474b;necf6c2[522]<=lq664c3;necf6c2[487]<=mt36875[0];necf6c2[482]<=dzd29c8;necf6c2[477]<=encc905[0];necf6c2[373]<=rte97cd[0];necf6c2[349]<=eafad08[0];necf6c2[338]<=uid1a77;necf6c2[336]<=kdf29d1;necf6c2[299]<=sjb47d6[0];necf6c2[290]<=ri14294[0];necf6c2[279]<=tu528e9;necf6c2[243]<=cb26d0e[0];necf6c2[186]<=qv1d2f9;necf6c2[169]<=fpba34e;necf6c2[168]<=ks3e53a;necf6c2[149]<=zxf68fa[0];necf6c2[121]<=ld64da1;necf6c2[84]<=jpd7469;necf6c2[60]<=ay4c9b4;necf6c2[42]<=co1ae8d;end         assign suff972 = necf6c2,ld7b613 = cme5c87;   initial begin   jcc030e = $fopen(".fred");   $fdisplay( jcc030e, "%3h\n%3h", (thc27c7 >> 4) & fnc7fe5, (thc27c7 >> (mt9f1ff+4)) & fnc7fe5 );   $fclose(jcc030e);   $readmemh(".fred", qg721c0);   end   always @ (suff972) begin   ym8700c = qg721c0[1];       for (vk1872=0; vk1872<qgdb09f; vk1872=vk1872+1) begin           cme5c87[vk1872] = suff972[ym8700c];       rv38061  = ^(ym8700c & qg721c0[0]);       ym8700c =  {ym8700c, rv38061};       end   end
endmodule