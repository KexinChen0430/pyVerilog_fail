module fir_band_pass_st (clk,
              rst,
              data_in,
              clk_en,
              rdy_to_ld,
              done,
              fir_result);
parameter DATA_WIDTH  = 11;
parameter COEF_WIDTH  = 11;
parameter ACCUM_WIDTH = 24;
parameter MSB_RM = 0;
parameter LSB_RM = 8;
parameter WIDTH_SAT = ACCUM_WIDTH-LSB_RM;
input clk, rst;
input [DATA_WIDTH-1:0] data_in;
input clk_en;
output rdy_to_ld;
wire rdy_to_ld;
wire rdy_int;
wire data_ld;
output done;
wire done;
wire done_int;
output [ACCUM_WIDTH-MSB_RM-LSB_RM-1:0] fir_result;
wire addr_low;
assign addr_low = 1'b0;
wire inv_rst;
assign inv_rst = ~rst;
assign data_ld = rdy_int;
wire [10:0] tdl_0_n;
wire [10:0] tdl_1_n;
wire [10:0] tdl_2_n;
wire [10:0] tdl_3_n;
wire [10:0] tdl_4_n;
wire [10:0] tdl_5_n;
wire [10:0] tdl_6_n;
wire [10:0] tdl_7_n;
wire [10:0] tdl_8_n;
wire [10:0] tdl_9_n;
wire [10:0] tdl_10_n;
wire [10:0] tdl_11_n;
wire [10:0] tdl_12_n;
wire [10:0] tdl_13_n;
wire [10:0] tdl_14_n;
wire [10:0] tdl_15_n;
wire [10:0] tdl_16_n;
wire [10:0] tdl_17_n;
wire [10:0] tdl_18_n;
wire [10:0] tdl_19_n;
wire [10:0] tdl_20_n;
wire [10:0] tdl_21_n;
wire [10:0] tdl_22_n;
wire [10:0] tdl_23_n;
wire [10:0] tdl_24_n;
wire [10:0] tdl_25_n;
wire [10:0] tdl_26_n;
wire [10:0] tdl_27_n;
wire [10:0] tdl_28_n;
wire [10:0] tdl_29_n;
wire [10:0] tdl_30_n;
wire [10:0] tdl_31_n;
tdl_da_lc Utdldalc0n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(data_in), .data_out(tdl_0_n) );
defparam Utdldalc0n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc1n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_0_n), .data_out(tdl_1_n) );
defparam Utdldalc1n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc2n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_1_n), .data_out(tdl_2_n) );
defparam Utdldalc2n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc3n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_2_n), .data_out(tdl_3_n) );
defparam Utdldalc3n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc4n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_3_n), .data_out(tdl_4_n) );
defparam Utdldalc4n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc5n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_4_n), .data_out(tdl_5_n) );
defparam Utdldalc5n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc6n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_5_n), .data_out(tdl_6_n) );
defparam Utdldalc6n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc7n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_6_n), .data_out(tdl_7_n) );
defparam Utdldalc7n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc8n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_7_n), .data_out(tdl_8_n) );
defparam Utdldalc8n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc9n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_8_n), .data_out(tdl_9_n) );
defparam Utdldalc9n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc10n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_9_n), .data_out(tdl_10_n) );
defparam Utdldalc10n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc11n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_10_n), .data_out(tdl_11_n) );
defparam Utdldalc11n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc12n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_11_n), .data_out(tdl_12_n) );
defparam Utdldalc12n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc13n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_12_n), .data_out(tdl_13_n) );
defparam Utdldalc13n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc14n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_13_n), .data_out(tdl_14_n) );
defparam Utdldalc14n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc15n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_14_n), .data_out(tdl_15_n) );
defparam Utdldalc15n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc16n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_15_n), .data_out(tdl_16_n) );
defparam Utdldalc16n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc17n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_16_n), .data_out(tdl_17_n) );
defparam Utdldalc17n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc18n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_17_n), .data_out(tdl_18_n) );
defparam Utdldalc18n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc19n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_18_n), .data_out(tdl_19_n) );
defparam Utdldalc19n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc20n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_19_n), .data_out(tdl_20_n) );
defparam Utdldalc20n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc21n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_20_n), .data_out(tdl_21_n) );
defparam Utdldalc21n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc22n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_21_n), .data_out(tdl_22_n) );
defparam Utdldalc22n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc23n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_22_n), .data_out(tdl_23_n) );
defparam Utdldalc23n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc24n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_23_n), .data_out(tdl_24_n) );
defparam Utdldalc24n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc25n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_24_n), .data_out(tdl_25_n) );
defparam Utdldalc25n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc26n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_25_n), .data_out(tdl_26_n) );
defparam Utdldalc26n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc27n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_26_n), .data_out(tdl_27_n) );
defparam Utdldalc27n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc28n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_27_n), .data_out(tdl_28_n) );
defparam Utdldalc28n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc29n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_28_n), .data_out(tdl_29_n) );
defparam Utdldalc29n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc30n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_29_n), .data_out(tdl_30_n) );
defparam Utdldalc30n.WIDTH = DATA_WIDTH;
tdl_da_lc Utdldalc31n (.clk(clk), .clk_en(rdy_int & clk_en),.rst(rst),.data_in(tdl_30_n), .data_out(tdl_31_n) );
defparam Utdldalc31n.WIDTH = DATA_WIDTH;
// symmetrical adders ...
wire [11:0] sym_res_0_n;
sadd_cen U_0_sym_add (.clk(clk), .gclk_en(clk_en), .ain(tdl_0_n), .bin(tdl_31_n), .res(sym_res_0_n) );
defparam U_0_sym_add.IN_WIDTH = 11;
defparam U_0_sym_add.PIPE_DEPTH = 1;
wire [11:0] sym_res_1_n;
sadd_cen U_1_sym_add (.clk(clk), .gclk_en(clk_en), .ain(tdl_1_n), .bin(tdl_30_n), .res(sym_res_1_n) );
defparam U_1_sym_add.IN_WIDTH = 11;
defparam U_1_sym_add.PIPE_DEPTH = 1;
wire [11:0] sym_res_2_n;
sadd_cen U_2_sym_add (.clk(clk), .gclk_en(clk_en), .ain(tdl_2_n), .bin(tdl_29_n), .res(sym_res_2_n) );
defparam U_2_sym_add.IN_WIDTH = 11;
defparam U_2_sym_add.PIPE_DEPTH = 1;
wire [11:0] sym_res_3_n;
sadd_cen U_3_sym_add (.clk(clk), .gclk_en(clk_en), .ain(tdl_3_n), .bin(tdl_28_n), .res(sym_res_3_n) );
defparam U_3_sym_add.IN_WIDTH = 11;
defparam U_3_sym_add.PIPE_DEPTH = 1;
wire [11:0] sym_res_4_n;
sadd_cen U_4_sym_add (.clk(clk), .gclk_en(clk_en), .ain(tdl_4_n), .bin(tdl_27_n), .res(sym_res_4_n) );
defparam U_4_sym_add.IN_WIDTH = 11;
defparam U_4_sym_add.PIPE_DEPTH = 1;
wire [11:0] sym_res_5_n;
sadd_cen U_5_sym_add (.clk(clk), .gclk_en(clk_en), .ain(tdl_5_n), .bin(tdl_26_n), .res(sym_res_5_n) );
defparam U_5_sym_add.IN_WIDTH = 11;
defparam U_5_sym_add.PIPE_DEPTH = 1;
wire [11:0] sym_res_6_n;
sadd_cen U_6_sym_add (.clk(clk), .gclk_en(clk_en), .ain(tdl_6_n), .bin(tdl_25_n), .res(sym_res_6_n) );
defparam U_6_sym_add.IN_WIDTH = 11;
defparam U_6_sym_add.PIPE_DEPTH = 1;
wire [11:0] sym_res_7_n;
sadd_cen U_7_sym_add (.clk(clk), .gclk_en(clk_en), .ain(tdl_7_n), .bin(tdl_24_n), .res(sym_res_7_n) );
defparam U_7_sym_add.IN_WIDTH = 11;
defparam U_7_sym_add.PIPE_DEPTH = 1;
wire [11:0] sym_res_8_n;
sadd_cen U_8_sym_add (.clk(clk), .gclk_en(clk_en), .ain(tdl_8_n), .bin(tdl_23_n), .res(sym_res_8_n) );
defparam U_8_sym_add.IN_WIDTH = 11;
defparam U_8_sym_add.PIPE_DEPTH = 1;
wire [11:0] sym_res_9_n;
sadd_cen U_9_sym_add (.clk(clk), .gclk_en(clk_en), .ain(tdl_9_n), .bin(tdl_22_n), .res(sym_res_9_n) );
defparam U_9_sym_add.IN_WIDTH = 11;
defparam U_9_sym_add.PIPE_DEPTH = 1;
wire [11:0] sym_res_10_n;
sadd_cen U_10_sym_add (.clk(clk), .gclk_en(clk_en), .ain(tdl_10_n), .bin(tdl_21_n), .res(sym_res_10_n) );
defparam U_10_sym_add.IN_WIDTH = 11;
defparam U_10_sym_add.PIPE_DEPTH = 1;
wire [11:0] sym_res_11_n;
sadd_cen U_11_sym_add (.clk(clk), .gclk_en(clk_en), .ain(tdl_11_n), .bin(tdl_20_n), .res(sym_res_11_n) );
defparam U_11_sym_add.IN_WIDTH = 11;
defparam U_11_sym_add.PIPE_DEPTH = 1;
wire [11:0] sym_res_12_n;
sadd_cen U_12_sym_add (.clk(clk), .gclk_en(clk_en), .ain(tdl_12_n), .bin(tdl_19_n), .res(sym_res_12_n) );
defparam U_12_sym_add.IN_WIDTH = 11;
defparam U_12_sym_add.PIPE_DEPTH = 1;
wire [11:0] sym_res_13_n;
sadd_cen U_13_sym_add (.clk(clk), .gclk_en(clk_en), .ain(tdl_13_n), .bin(tdl_18_n), .res(sym_res_13_n) );
defparam U_13_sym_add.IN_WIDTH = 11;
defparam U_13_sym_add.PIPE_DEPTH = 1;
wire [11:0] sym_res_14_n;
sadd_cen U_14_sym_add (.clk(clk), .gclk_en(clk_en), .ain(tdl_14_n), .bin(tdl_17_n), .res(sym_res_14_n) );
defparam U_14_sym_add.IN_WIDTH = 11;
defparam U_14_sym_add.PIPE_DEPTH = 1;
wire [11:0] sym_res_15_n;
sadd_cen U_15_sym_add (.clk(clk), .gclk_en(clk_en), .ain(tdl_15_n), .bin(tdl_16_n), .res(sym_res_15_n) );
defparam U_15_sym_add.IN_WIDTH = 11;
defparam U_15_sym_add.PIPE_DEPTH = 1;
wire [10:0] lut_val_0_n_0_pp;
rom_lut_r_cen Ur0_n_0_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_4_n[0],sym_res_3_n[0],sym_res_2_n[0],sym_res_1_n[0] } ), .data_out( lut_val_0_n_0_pp[5:0]) ) ;
 defparam Ur0_n_0_pp.DATA_WIDTH = 6;
defparam Ur0_n_0_pp.C0 = 6'd                   0;
defparam Ur0_n_0_pp.C1 = 6'd                   1;
defparam Ur0_n_0_pp.C2 = 6'd                  59;
defparam Ur0_n_0_pp.C3 = 6'd                  60;
defparam Ur0_n_0_pp.C4 = 6'd                  50;
defparam Ur0_n_0_pp.C5 = 6'd                  51;
defparam Ur0_n_0_pp.C6 = 6'd                  45;
defparam Ur0_n_0_pp.C7 = 6'd                  46;
defparam Ur0_n_0_pp.C8 = 6'd                   2;
defparam Ur0_n_0_pp.C9 = 6'd                   3;
defparam Ur0_n_0_pp.CA = 6'd                  61;
defparam Ur0_n_0_pp.CB = 6'd                  62;
defparam Ur0_n_0_pp.CC = 6'd                  52;
defparam Ur0_n_0_pp.CD = 6'd                  53;
defparam Ur0_n_0_pp.CE = 6'd                  47;
defparam Ur0_n_0_pp.CF = 6'd                  48;
assign lut_val_0_n_0_pp[10] = lut_val_0_n_0_pp[5];
assign lut_val_0_n_0_pp[9] = lut_val_0_n_0_pp[5];
assign lut_val_0_n_0_pp[8] = lut_val_0_n_0_pp[5];
assign lut_val_0_n_0_pp[7] = lut_val_0_n_0_pp[5];
assign lut_val_0_n_0_pp[6] = lut_val_0_n_0_pp[5];
wire [10:0] lut_val_0_n_1_pp;
rom_lut_r_cen Ur0_n_1_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_4_n[1],sym_res_3_n[1],sym_res_2_n[1],sym_res_1_n[1] } ), .data_out( lut_val_0_n_1_pp[5:0]) ) ;
 defparam Ur0_n_1_pp.DATA_WIDTH = 6;
defparam Ur0_n_1_pp.C0 = 6'd                   0;
defparam Ur0_n_1_pp.C1 = 6'd                   1;
defparam Ur0_n_1_pp.C2 = 6'd                  59;
defparam Ur0_n_1_pp.C3 = 6'd                  60;
defparam Ur0_n_1_pp.C4 = 6'd                  50;
defparam Ur0_n_1_pp.C5 = 6'd                  51;
defparam Ur0_n_1_pp.C6 = 6'd                  45;
defparam Ur0_n_1_pp.C7 = 6'd                  46;
defparam Ur0_n_1_pp.C8 = 6'd                   2;
defparam Ur0_n_1_pp.C9 = 6'd                   3;
defparam Ur0_n_1_pp.CA = 6'd                  61;
defparam Ur0_n_1_pp.CB = 6'd                  62;
defparam Ur0_n_1_pp.CC = 6'd                  52;
defparam Ur0_n_1_pp.CD = 6'd                  53;
defparam Ur0_n_1_pp.CE = 6'd                  47;
defparam Ur0_n_1_pp.CF = 6'd                  48;
assign lut_val_0_n_1_pp[10] = lut_val_0_n_1_pp[5];
assign lut_val_0_n_1_pp[9] = lut_val_0_n_1_pp[5];
assign lut_val_0_n_1_pp[8] = lut_val_0_n_1_pp[5];
assign lut_val_0_n_1_pp[7] = lut_val_0_n_1_pp[5];
assign lut_val_0_n_1_pp[6] = lut_val_0_n_1_pp[5];
wire [10:0] lut_val_0_n_2_pp;
rom_lut_r_cen Ur0_n_2_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_4_n[2],sym_res_3_n[2],sym_res_2_n[2],sym_res_1_n[2] } ), .data_out( lut_val_0_n_2_pp[5:0]) ) ;
 defparam Ur0_n_2_pp.DATA_WIDTH = 6;
defparam Ur0_n_2_pp.C0 = 6'd                   0;
defparam Ur0_n_2_pp.C1 = 6'd                   1;
defparam Ur0_n_2_pp.C2 = 6'd                  59;
defparam Ur0_n_2_pp.C3 = 6'd                  60;
defparam Ur0_n_2_pp.C4 = 6'd                  50;
defparam Ur0_n_2_pp.C5 = 6'd                  51;
defparam Ur0_n_2_pp.C6 = 6'd                  45;
defparam Ur0_n_2_pp.C7 = 6'd                  46;
defparam Ur0_n_2_pp.C8 = 6'd                   2;
defparam Ur0_n_2_pp.C9 = 6'd                   3;
defparam Ur0_n_2_pp.CA = 6'd                  61;
defparam Ur0_n_2_pp.CB = 6'd                  62;
defparam Ur0_n_2_pp.CC = 6'd                  52;
defparam Ur0_n_2_pp.CD = 6'd                  53;
defparam Ur0_n_2_pp.CE = 6'd                  47;
defparam Ur0_n_2_pp.CF = 6'd                  48;
assign lut_val_0_n_2_pp[10] = lut_val_0_n_2_pp[5];
assign lut_val_0_n_2_pp[9] = lut_val_0_n_2_pp[5];
assign lut_val_0_n_2_pp[8] = lut_val_0_n_2_pp[5];
assign lut_val_0_n_2_pp[7] = lut_val_0_n_2_pp[5];
assign lut_val_0_n_2_pp[6] = lut_val_0_n_2_pp[5];
wire [10:0] lut_val_0_n_3_pp;
rom_lut_r_cen Ur0_n_3_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_4_n[3],sym_res_3_n[3],sym_res_2_n[3],sym_res_1_n[3] } ), .data_out( lut_val_0_n_3_pp[5:0]) ) ;
 defparam Ur0_n_3_pp.DATA_WIDTH = 6;
defparam Ur0_n_3_pp.C0 = 6'd                   0;
defparam Ur0_n_3_pp.C1 = 6'd                   1;
defparam Ur0_n_3_pp.C2 = 6'd                  59;
defparam Ur0_n_3_pp.C3 = 6'd                  60;
defparam Ur0_n_3_pp.C4 = 6'd                  50;
defparam Ur0_n_3_pp.C5 = 6'd                  51;
defparam Ur0_n_3_pp.C6 = 6'd                  45;
defparam Ur0_n_3_pp.C7 = 6'd                  46;
defparam Ur0_n_3_pp.C8 = 6'd                   2;
defparam Ur0_n_3_pp.C9 = 6'd                   3;
defparam Ur0_n_3_pp.CA = 6'd                  61;
defparam Ur0_n_3_pp.CB = 6'd                  62;
defparam Ur0_n_3_pp.CC = 6'd                  52;
defparam Ur0_n_3_pp.CD = 6'd                  53;
defparam Ur0_n_3_pp.CE = 6'd                  47;
defparam Ur0_n_3_pp.CF = 6'd                  48;
assign lut_val_0_n_3_pp[10] = lut_val_0_n_3_pp[5];
assign lut_val_0_n_3_pp[9] = lut_val_0_n_3_pp[5];
assign lut_val_0_n_3_pp[8] = lut_val_0_n_3_pp[5];
assign lut_val_0_n_3_pp[7] = lut_val_0_n_3_pp[5];
assign lut_val_0_n_3_pp[6] = lut_val_0_n_3_pp[5];
wire [10:0] lut_val_0_n_4_pp;
rom_lut_r_cen Ur0_n_4_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_4_n[4],sym_res_3_n[4],sym_res_2_n[4],sym_res_1_n[4] } ), .data_out( lut_val_0_n_4_pp[5:0]) ) ;
 defparam Ur0_n_4_pp.DATA_WIDTH = 6;
defparam Ur0_n_4_pp.C0 = 6'd                   0;
defparam Ur0_n_4_pp.C1 = 6'd                   1;
defparam Ur0_n_4_pp.C2 = 6'd                  59;
defparam Ur0_n_4_pp.C3 = 6'd                  60;
defparam Ur0_n_4_pp.C4 = 6'd                  50;
defparam Ur0_n_4_pp.C5 = 6'd                  51;
defparam Ur0_n_4_pp.C6 = 6'd                  45;
defparam Ur0_n_4_pp.C7 = 6'd                  46;
defparam Ur0_n_4_pp.C8 = 6'd                   2;
defparam Ur0_n_4_pp.C9 = 6'd                   3;
defparam Ur0_n_4_pp.CA = 6'd                  61;
defparam Ur0_n_4_pp.CB = 6'd                  62;
defparam Ur0_n_4_pp.CC = 6'd                  52;
defparam Ur0_n_4_pp.CD = 6'd                  53;
defparam Ur0_n_4_pp.CE = 6'd                  47;
defparam Ur0_n_4_pp.CF = 6'd                  48;
assign lut_val_0_n_4_pp[10] = lut_val_0_n_4_pp[5];
assign lut_val_0_n_4_pp[9] = lut_val_0_n_4_pp[5];
assign lut_val_0_n_4_pp[8] = lut_val_0_n_4_pp[5];
assign lut_val_0_n_4_pp[7] = lut_val_0_n_4_pp[5];
assign lut_val_0_n_4_pp[6] = lut_val_0_n_4_pp[5];
wire [10:0] lut_val_0_n_5_pp;
rom_lut_r_cen Ur0_n_5_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_4_n[5],sym_res_3_n[5],sym_res_2_n[5],sym_res_1_n[5] } ), .data_out( lut_val_0_n_5_pp[5:0]) ) ;
 defparam Ur0_n_5_pp.DATA_WIDTH = 6;
defparam Ur0_n_5_pp.C0 = 6'd                   0;
defparam Ur0_n_5_pp.C1 = 6'd                   1;
defparam Ur0_n_5_pp.C2 = 6'd                  59;
defparam Ur0_n_5_pp.C3 = 6'd                  60;
defparam Ur0_n_5_pp.C4 = 6'd                  50;
defparam Ur0_n_5_pp.C5 = 6'd                  51;
defparam Ur0_n_5_pp.C6 = 6'd                  45;
defparam Ur0_n_5_pp.C7 = 6'd                  46;
defparam Ur0_n_5_pp.C8 = 6'd                   2;
defparam Ur0_n_5_pp.C9 = 6'd                   3;
defparam Ur0_n_5_pp.CA = 6'd                  61;
defparam Ur0_n_5_pp.CB = 6'd                  62;
defparam Ur0_n_5_pp.CC = 6'd                  52;
defparam Ur0_n_5_pp.CD = 6'd                  53;
defparam Ur0_n_5_pp.CE = 6'd                  47;
defparam Ur0_n_5_pp.CF = 6'd                  48;
assign lut_val_0_n_5_pp[10] = lut_val_0_n_5_pp[5];
assign lut_val_0_n_5_pp[9] = lut_val_0_n_5_pp[5];
assign lut_val_0_n_5_pp[8] = lut_val_0_n_5_pp[5];
assign lut_val_0_n_5_pp[7] = lut_val_0_n_5_pp[5];
assign lut_val_0_n_5_pp[6] = lut_val_0_n_5_pp[5];
wire [10:0] lut_val_0_n_6_pp;
rom_lut_r_cen Ur0_n_6_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_4_n[6],sym_res_3_n[6],sym_res_2_n[6],sym_res_1_n[6] } ), .data_out( lut_val_0_n_6_pp[5:0]) ) ;
 defparam Ur0_n_6_pp.DATA_WIDTH = 6;
defparam Ur0_n_6_pp.C0 = 6'd                   0;
defparam Ur0_n_6_pp.C1 = 6'd                   1;
defparam Ur0_n_6_pp.C2 = 6'd                  59;
defparam Ur0_n_6_pp.C3 = 6'd                  60;
defparam Ur0_n_6_pp.C4 = 6'd                  50;
defparam Ur0_n_6_pp.C5 = 6'd                  51;
defparam Ur0_n_6_pp.C6 = 6'd                  45;
defparam Ur0_n_6_pp.C7 = 6'd                  46;
defparam Ur0_n_6_pp.C8 = 6'd                   2;
defparam Ur0_n_6_pp.C9 = 6'd                   3;
defparam Ur0_n_6_pp.CA = 6'd                  61;
defparam Ur0_n_6_pp.CB = 6'd                  62;
defparam Ur0_n_6_pp.CC = 6'd                  52;
defparam Ur0_n_6_pp.CD = 6'd                  53;
defparam Ur0_n_6_pp.CE = 6'd                  47;
defparam Ur0_n_6_pp.CF = 6'd                  48;
assign lut_val_0_n_6_pp[10] = lut_val_0_n_6_pp[5];
assign lut_val_0_n_6_pp[9] = lut_val_0_n_6_pp[5];
assign lut_val_0_n_6_pp[8] = lut_val_0_n_6_pp[5];
assign lut_val_0_n_6_pp[7] = lut_val_0_n_6_pp[5];
assign lut_val_0_n_6_pp[6] = lut_val_0_n_6_pp[5];
wire [10:0] lut_val_0_n_7_pp;
rom_lut_r_cen Ur0_n_7_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_4_n[7],sym_res_3_n[7],sym_res_2_n[7],sym_res_1_n[7] } ), .data_out( lut_val_0_n_7_pp[5:0]) ) ;
 defparam Ur0_n_7_pp.DATA_WIDTH = 6;
defparam Ur0_n_7_pp.C0 = 6'd                   0;
defparam Ur0_n_7_pp.C1 = 6'd                   1;
defparam Ur0_n_7_pp.C2 = 6'd                  59;
defparam Ur0_n_7_pp.C3 = 6'd                  60;
defparam Ur0_n_7_pp.C4 = 6'd                  50;
defparam Ur0_n_7_pp.C5 = 6'd                  51;
defparam Ur0_n_7_pp.C6 = 6'd                  45;
defparam Ur0_n_7_pp.C7 = 6'd                  46;
defparam Ur0_n_7_pp.C8 = 6'd                   2;
defparam Ur0_n_7_pp.C9 = 6'd                   3;
defparam Ur0_n_7_pp.CA = 6'd                  61;
defparam Ur0_n_7_pp.CB = 6'd                  62;
defparam Ur0_n_7_pp.CC = 6'd                  52;
defparam Ur0_n_7_pp.CD = 6'd                  53;
defparam Ur0_n_7_pp.CE = 6'd                  47;
defparam Ur0_n_7_pp.CF = 6'd                  48;
assign lut_val_0_n_7_pp[10] = lut_val_0_n_7_pp[5];
assign lut_val_0_n_7_pp[9] = lut_val_0_n_7_pp[5];
assign lut_val_0_n_7_pp[8] = lut_val_0_n_7_pp[5];
assign lut_val_0_n_7_pp[7] = lut_val_0_n_7_pp[5];
assign lut_val_0_n_7_pp[6] = lut_val_0_n_7_pp[5];
wire [10:0] lut_val_0_n_8_pp;
rom_lut_r_cen Ur0_n_8_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_4_n[8],sym_res_3_n[8],sym_res_2_n[8],sym_res_1_n[8] } ), .data_out( lut_val_0_n_8_pp[5:0]) ) ;
 defparam Ur0_n_8_pp.DATA_WIDTH = 6;
defparam Ur0_n_8_pp.C0 = 6'd                   0;
defparam Ur0_n_8_pp.C1 = 6'd                   1;
defparam Ur0_n_8_pp.C2 = 6'd                  59;
defparam Ur0_n_8_pp.C3 = 6'd                  60;
defparam Ur0_n_8_pp.C4 = 6'd                  50;
defparam Ur0_n_8_pp.C5 = 6'd                  51;
defparam Ur0_n_8_pp.C6 = 6'd                  45;
defparam Ur0_n_8_pp.C7 = 6'd                  46;
defparam Ur0_n_8_pp.C8 = 6'd                   2;
defparam Ur0_n_8_pp.C9 = 6'd                   3;
defparam Ur0_n_8_pp.CA = 6'd                  61;
defparam Ur0_n_8_pp.CB = 6'd                  62;
defparam Ur0_n_8_pp.CC = 6'd                  52;
defparam Ur0_n_8_pp.CD = 6'd                  53;
defparam Ur0_n_8_pp.CE = 6'd                  47;
defparam Ur0_n_8_pp.CF = 6'd                  48;
assign lut_val_0_n_8_pp[10] = lut_val_0_n_8_pp[5];
assign lut_val_0_n_8_pp[9] = lut_val_0_n_8_pp[5];
assign lut_val_0_n_8_pp[8] = lut_val_0_n_8_pp[5];
assign lut_val_0_n_8_pp[7] = lut_val_0_n_8_pp[5];
assign lut_val_0_n_8_pp[6] = lut_val_0_n_8_pp[5];
wire [10:0] lut_val_0_n_9_pp;
rom_lut_r_cen Ur0_n_9_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_4_n[9],sym_res_3_n[9],sym_res_2_n[9],sym_res_1_n[9] } ), .data_out( lut_val_0_n_9_pp[5:0]) ) ;
 defparam Ur0_n_9_pp.DATA_WIDTH = 6;
defparam Ur0_n_9_pp.C0 = 6'd                   0;
defparam Ur0_n_9_pp.C1 = 6'd                   1;
defparam Ur0_n_9_pp.C2 = 6'd                  59;
defparam Ur0_n_9_pp.C3 = 6'd                  60;
defparam Ur0_n_9_pp.C4 = 6'd                  50;
defparam Ur0_n_9_pp.C5 = 6'd                  51;
defparam Ur0_n_9_pp.C6 = 6'd                  45;
defparam Ur0_n_9_pp.C7 = 6'd                  46;
defparam Ur0_n_9_pp.C8 = 6'd                   2;
defparam Ur0_n_9_pp.C9 = 6'd                   3;
defparam Ur0_n_9_pp.CA = 6'd                  61;
defparam Ur0_n_9_pp.CB = 6'd                  62;
defparam Ur0_n_9_pp.CC = 6'd                  52;
defparam Ur0_n_9_pp.CD = 6'd                  53;
defparam Ur0_n_9_pp.CE = 6'd                  47;
defparam Ur0_n_9_pp.CF = 6'd                  48;
assign lut_val_0_n_9_pp[10] = lut_val_0_n_9_pp[5];
assign lut_val_0_n_9_pp[9] = lut_val_0_n_9_pp[5];
assign lut_val_0_n_9_pp[8] = lut_val_0_n_9_pp[5];
assign lut_val_0_n_9_pp[7] = lut_val_0_n_9_pp[5];
assign lut_val_0_n_9_pp[6] = lut_val_0_n_9_pp[5];
wire [10:0] lut_val_0_n_10_pp;
rom_lut_r_cen Ur0_n_10_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_4_n[10],sym_res_3_n[10],sym_res_2_n[10],sym_res_1_n[10] } ), .data_out( lut_val_0_n_10_pp[5:0]) ) ;
 defparam Ur0_n_10_pp.DATA_WIDTH = 6;
defparam Ur0_n_10_pp.C0 = 6'd                   0;
defparam Ur0_n_10_pp.C1 = 6'd                   1;
defparam Ur0_n_10_pp.C2 = 6'd                  59;
defparam Ur0_n_10_pp.C3 = 6'd                  60;
defparam Ur0_n_10_pp.C4 = 6'd                  50;
defparam Ur0_n_10_pp.C5 = 6'd                  51;
defparam Ur0_n_10_pp.C6 = 6'd                  45;
defparam Ur0_n_10_pp.C7 = 6'd                  46;
defparam Ur0_n_10_pp.C8 = 6'd                   2;
defparam Ur0_n_10_pp.C9 = 6'd                   3;
defparam Ur0_n_10_pp.CA = 6'd                  61;
defparam Ur0_n_10_pp.CB = 6'd                  62;
defparam Ur0_n_10_pp.CC = 6'd                  52;
defparam Ur0_n_10_pp.CD = 6'd                  53;
defparam Ur0_n_10_pp.CE = 6'd                  47;
defparam Ur0_n_10_pp.CF = 6'd                  48;
assign lut_val_0_n_10_pp[10] = lut_val_0_n_10_pp[5];
assign lut_val_0_n_10_pp[9] = lut_val_0_n_10_pp[5];
assign lut_val_0_n_10_pp[8] = lut_val_0_n_10_pp[5];
assign lut_val_0_n_10_pp[7] = lut_val_0_n_10_pp[5];
assign lut_val_0_n_10_pp[6] = lut_val_0_n_10_pp[5];
wire [10:0] lut_val_0_n_11_pp;
rom_lut_r_cen Ur0_n_11_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_4_n[11],sym_res_3_n[11],sym_res_2_n[11],sym_res_1_n[11] } ), .data_out( lut_val_0_n_11_pp[5:0]) ) ;
 defparam Ur0_n_11_pp.DATA_WIDTH = 6;
defparam Ur0_n_11_pp.C0 = 6'd                   0;
defparam Ur0_n_11_pp.C1 = 6'd                  63;
defparam Ur0_n_11_pp.C2 = 6'd                   5;
defparam Ur0_n_11_pp.C3 = 6'd                   4;
defparam Ur0_n_11_pp.C4 = 6'd                  14;
defparam Ur0_n_11_pp.C5 = 6'd                  13;
defparam Ur0_n_11_pp.C6 = 6'd                  19;
defparam Ur0_n_11_pp.C7 = 6'd                  18;
defparam Ur0_n_11_pp.C8 = 6'd                  62;
defparam Ur0_n_11_pp.C9 = 6'd                  61;
defparam Ur0_n_11_pp.CA = 6'd                   3;
defparam Ur0_n_11_pp.CB = 6'd                   2;
defparam Ur0_n_11_pp.CC = 6'd                  12;
defparam Ur0_n_11_pp.CD = 6'd                  11;
defparam Ur0_n_11_pp.CE = 6'd                  17;
defparam Ur0_n_11_pp.CF = 6'd                  16;
assign lut_val_0_n_11_pp[10] = lut_val_0_n_11_pp[5];
assign lut_val_0_n_11_pp[9] = lut_val_0_n_11_pp[5];
assign lut_val_0_n_11_pp[8] = lut_val_0_n_11_pp[5];
assign lut_val_0_n_11_pp[7] = lut_val_0_n_11_pp[5];
assign lut_val_0_n_11_pp[6] = lut_val_0_n_11_pp[5];
wire [10:0] lut_val_1_n_0_pp;
rom_lut_r_cen Ur1_n_0_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_9_n[0],sym_res_7_n[0],sym_res_6_n[0],sym_res_5_n[0] } ), .data_out( lut_val_1_n_0_pp[8:0]) ) ;
 defparam Ur1_n_0_pp.DATA_WIDTH = 9;
defparam Ur1_n_0_pp.C0 = 9'd                   0;
defparam Ur1_n_0_pp.C1 = 9'd                 486;
defparam Ur1_n_0_pp.C2 = 9'd                  14;
defparam Ur1_n_0_pp.C3 = 9'd                 500;
defparam Ur1_n_0_pp.C4 = 9'd                  70;
defparam Ur1_n_0_pp.C5 = 9'd                  44;
defparam Ur1_n_0_pp.C6 = 9'd                  84;
defparam Ur1_n_0_pp.C7 = 9'd                  58;
defparam Ur1_n_0_pp.C8 = 9'd                 127;
defparam Ur1_n_0_pp.C9 = 9'd                 101;
defparam Ur1_n_0_pp.CA = 9'd                 141;
defparam Ur1_n_0_pp.CB = 9'd                 115;
defparam Ur1_n_0_pp.CC = 9'd                 197;
defparam Ur1_n_0_pp.CD = 9'd                 171;
defparam Ur1_n_0_pp.CE = 9'd                 211;
defparam Ur1_n_0_pp.CF = 9'd                 185;
assign lut_val_1_n_0_pp[10] = lut_val_1_n_0_pp[8];
assign lut_val_1_n_0_pp[9] = lut_val_1_n_0_pp[8];
wire [10:0] lut_val_1_n_1_pp;
rom_lut_r_cen Ur1_n_1_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_9_n[1],sym_res_7_n[1],sym_res_6_n[1],sym_res_5_n[1] } ), .data_out( lut_val_1_n_1_pp[8:0]) ) ;
 defparam Ur1_n_1_pp.DATA_WIDTH = 9;
defparam Ur1_n_1_pp.C0 = 9'd                   0;
defparam Ur1_n_1_pp.C1 = 9'd                 486;
defparam Ur1_n_1_pp.C2 = 9'd                  14;
defparam Ur1_n_1_pp.C3 = 9'd                 500;
defparam Ur1_n_1_pp.C4 = 9'd                  70;
defparam Ur1_n_1_pp.C5 = 9'd                  44;
defparam Ur1_n_1_pp.C6 = 9'd                  84;
defparam Ur1_n_1_pp.C7 = 9'd                  58;
defparam Ur1_n_1_pp.C8 = 9'd                 127;
defparam Ur1_n_1_pp.C9 = 9'd                 101;
defparam Ur1_n_1_pp.CA = 9'd                 141;
defparam Ur1_n_1_pp.CB = 9'd                 115;
defparam Ur1_n_1_pp.CC = 9'd                 197;
defparam Ur1_n_1_pp.CD = 9'd                 171;
defparam Ur1_n_1_pp.CE = 9'd                 211;
defparam Ur1_n_1_pp.CF = 9'd                 185;
assign lut_val_1_n_1_pp[10] = lut_val_1_n_1_pp[8];
assign lut_val_1_n_1_pp[9] = lut_val_1_n_1_pp[8];
wire [10:0] lut_val_1_n_2_pp;
rom_lut_r_cen Ur1_n_2_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_9_n[2],sym_res_7_n[2],sym_res_6_n[2],sym_res_5_n[2] } ), .data_out( lut_val_1_n_2_pp[8:0]) ) ;
 defparam Ur1_n_2_pp.DATA_WIDTH = 9;
defparam Ur1_n_2_pp.C0 = 9'd                   0;
defparam Ur1_n_2_pp.C1 = 9'd                 486;
defparam Ur1_n_2_pp.C2 = 9'd                  14;
defparam Ur1_n_2_pp.C3 = 9'd                 500;
defparam Ur1_n_2_pp.C4 = 9'd                  70;
defparam Ur1_n_2_pp.C5 = 9'd                  44;
defparam Ur1_n_2_pp.C6 = 9'd                  84;
defparam Ur1_n_2_pp.C7 = 9'd                  58;
defparam Ur1_n_2_pp.C8 = 9'd                 127;
defparam Ur1_n_2_pp.C9 = 9'd                 101;
defparam Ur1_n_2_pp.CA = 9'd                 141;
defparam Ur1_n_2_pp.CB = 9'd                 115;
defparam Ur1_n_2_pp.CC = 9'd                 197;
defparam Ur1_n_2_pp.CD = 9'd                 171;
defparam Ur1_n_2_pp.CE = 9'd                 211;
defparam Ur1_n_2_pp.CF = 9'd                 185;
assign lut_val_1_n_2_pp[10] = lut_val_1_n_2_pp[8];
assign lut_val_1_n_2_pp[9] = lut_val_1_n_2_pp[8];
wire [10:0] lut_val_1_n_3_pp;
rom_lut_r_cen Ur1_n_3_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_9_n[3],sym_res_7_n[3],sym_res_6_n[3],sym_res_5_n[3] } ), .data_out( lut_val_1_n_3_pp[8:0]) ) ;
 defparam Ur1_n_3_pp.DATA_WIDTH = 9;
defparam Ur1_n_3_pp.C0 = 9'd                   0;
defparam Ur1_n_3_pp.C1 = 9'd                 486;
defparam Ur1_n_3_pp.C2 = 9'd                  14;
defparam Ur1_n_3_pp.C3 = 9'd                 500;
defparam Ur1_n_3_pp.C4 = 9'd                  70;
defparam Ur1_n_3_pp.C5 = 9'd                  44;
defparam Ur1_n_3_pp.C6 = 9'd                  84;
defparam Ur1_n_3_pp.C7 = 9'd                  58;
defparam Ur1_n_3_pp.C8 = 9'd                 127;
defparam Ur1_n_3_pp.C9 = 9'd                 101;
defparam Ur1_n_3_pp.CA = 9'd                 141;
defparam Ur1_n_3_pp.CB = 9'd                 115;
defparam Ur1_n_3_pp.CC = 9'd                 197;
defparam Ur1_n_3_pp.CD = 9'd                 171;
defparam Ur1_n_3_pp.CE = 9'd                 211;
defparam Ur1_n_3_pp.CF = 9'd                 185;
assign lut_val_1_n_3_pp[10] = lut_val_1_n_3_pp[8];
assign lut_val_1_n_3_pp[9] = lut_val_1_n_3_pp[8];
wire [10:0] lut_val_1_n_4_pp;
rom_lut_r_cen Ur1_n_4_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_9_n[4],sym_res_7_n[4],sym_res_6_n[4],sym_res_5_n[4] } ), .data_out( lut_val_1_n_4_pp[8:0]) ) ;
 defparam Ur1_n_4_pp.DATA_WIDTH = 9;
defparam Ur1_n_4_pp.C0 = 9'd                   0;
defparam Ur1_n_4_pp.C1 = 9'd                 486;
defparam Ur1_n_4_pp.C2 = 9'd                  14;
defparam Ur1_n_4_pp.C3 = 9'd                 500;
defparam Ur1_n_4_pp.C4 = 9'd                  70;
defparam Ur1_n_4_pp.C5 = 9'd                  44;
defparam Ur1_n_4_pp.C6 = 9'd                  84;
defparam Ur1_n_4_pp.C7 = 9'd                  58;
defparam Ur1_n_4_pp.C8 = 9'd                 127;
defparam Ur1_n_4_pp.C9 = 9'd                 101;
defparam Ur1_n_4_pp.CA = 9'd                 141;
defparam Ur1_n_4_pp.CB = 9'd                 115;
defparam Ur1_n_4_pp.CC = 9'd                 197;
defparam Ur1_n_4_pp.CD = 9'd                 171;
defparam Ur1_n_4_pp.CE = 9'd                 211;
defparam Ur1_n_4_pp.CF = 9'd                 185;
assign lut_val_1_n_4_pp[10] = lut_val_1_n_4_pp[8];
assign lut_val_1_n_4_pp[9] = lut_val_1_n_4_pp[8];
wire [10:0] lut_val_1_n_5_pp;
rom_lut_r_cen Ur1_n_5_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_9_n[5],sym_res_7_n[5],sym_res_6_n[5],sym_res_5_n[5] } ), .data_out( lut_val_1_n_5_pp[8:0]) ) ;
 defparam Ur1_n_5_pp.DATA_WIDTH = 9;
defparam Ur1_n_5_pp.C0 = 9'd                   0;
defparam Ur1_n_5_pp.C1 = 9'd                 486;
defparam Ur1_n_5_pp.C2 = 9'd                  14;
defparam Ur1_n_5_pp.C3 = 9'd                 500;
defparam Ur1_n_5_pp.C4 = 9'd                  70;
defparam Ur1_n_5_pp.C5 = 9'd                  44;
defparam Ur1_n_5_pp.C6 = 9'd                  84;
defparam Ur1_n_5_pp.C7 = 9'd                  58;
defparam Ur1_n_5_pp.C8 = 9'd                 127;
defparam Ur1_n_5_pp.C9 = 9'd                 101;
defparam Ur1_n_5_pp.CA = 9'd                 141;
defparam Ur1_n_5_pp.CB = 9'd                 115;
defparam Ur1_n_5_pp.CC = 9'd                 197;
defparam Ur1_n_5_pp.CD = 9'd                 171;
defparam Ur1_n_5_pp.CE = 9'd                 211;
defparam Ur1_n_5_pp.CF = 9'd                 185;
assign lut_val_1_n_5_pp[10] = lut_val_1_n_5_pp[8];
assign lut_val_1_n_5_pp[9] = lut_val_1_n_5_pp[8];
wire [10:0] lut_val_1_n_6_pp;
rom_lut_r_cen Ur1_n_6_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_9_n[6],sym_res_7_n[6],sym_res_6_n[6],sym_res_5_n[6] } ), .data_out( lut_val_1_n_6_pp[8:0]) ) ;
 defparam Ur1_n_6_pp.DATA_WIDTH = 9;
defparam Ur1_n_6_pp.C0 = 9'd                   0;
defparam Ur1_n_6_pp.C1 = 9'd                 486;
defparam Ur1_n_6_pp.C2 = 9'd                  14;
defparam Ur1_n_6_pp.C3 = 9'd                 500;
defparam Ur1_n_6_pp.C4 = 9'd                  70;
defparam Ur1_n_6_pp.C5 = 9'd                  44;
defparam Ur1_n_6_pp.C6 = 9'd                  84;
defparam Ur1_n_6_pp.C7 = 9'd                  58;
defparam Ur1_n_6_pp.C8 = 9'd                 127;
defparam Ur1_n_6_pp.C9 = 9'd                 101;
defparam Ur1_n_6_pp.CA = 9'd                 141;
defparam Ur1_n_6_pp.CB = 9'd                 115;
defparam Ur1_n_6_pp.CC = 9'd                 197;
defparam Ur1_n_6_pp.CD = 9'd                 171;
defparam Ur1_n_6_pp.CE = 9'd                 211;
defparam Ur1_n_6_pp.CF = 9'd                 185;
assign lut_val_1_n_6_pp[10] = lut_val_1_n_6_pp[8];
assign lut_val_1_n_6_pp[9] = lut_val_1_n_6_pp[8];
wire [10:0] lut_val_1_n_7_pp;
rom_lut_r_cen Ur1_n_7_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_9_n[7],sym_res_7_n[7],sym_res_6_n[7],sym_res_5_n[7] } ), .data_out( lut_val_1_n_7_pp[8:0]) ) ;
 defparam Ur1_n_7_pp.DATA_WIDTH = 9;
defparam Ur1_n_7_pp.C0 = 9'd                   0;
defparam Ur1_n_7_pp.C1 = 9'd                 486;
defparam Ur1_n_7_pp.C2 = 9'd                  14;
defparam Ur1_n_7_pp.C3 = 9'd                 500;
defparam Ur1_n_7_pp.C4 = 9'd                  70;
defparam Ur1_n_7_pp.C5 = 9'd                  44;
defparam Ur1_n_7_pp.C6 = 9'd                  84;
defparam Ur1_n_7_pp.C7 = 9'd                  58;
defparam Ur1_n_7_pp.C8 = 9'd                 127;
defparam Ur1_n_7_pp.C9 = 9'd                 101;
defparam Ur1_n_7_pp.CA = 9'd                 141;
defparam Ur1_n_7_pp.CB = 9'd                 115;
defparam Ur1_n_7_pp.CC = 9'd                 197;
defparam Ur1_n_7_pp.CD = 9'd                 171;
defparam Ur1_n_7_pp.CE = 9'd                 211;
defparam Ur1_n_7_pp.CF = 9'd                 185;
assign lut_val_1_n_7_pp[10] = lut_val_1_n_7_pp[8];
assign lut_val_1_n_7_pp[9] = lut_val_1_n_7_pp[8];
wire [10:0] lut_val_1_n_8_pp;
rom_lut_r_cen Ur1_n_8_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_9_n[8],sym_res_7_n[8],sym_res_6_n[8],sym_res_5_n[8] } ), .data_out( lut_val_1_n_8_pp[8:0]) ) ;
 defparam Ur1_n_8_pp.DATA_WIDTH = 9;
defparam Ur1_n_8_pp.C0 = 9'd                   0;
defparam Ur1_n_8_pp.C1 = 9'd                 486;
defparam Ur1_n_8_pp.C2 = 9'd                  14;
defparam Ur1_n_8_pp.C3 = 9'd                 500;
defparam Ur1_n_8_pp.C4 = 9'd                  70;
defparam Ur1_n_8_pp.C5 = 9'd                  44;
defparam Ur1_n_8_pp.C6 = 9'd                  84;
defparam Ur1_n_8_pp.C7 = 9'd                  58;
defparam Ur1_n_8_pp.C8 = 9'd                 127;
defparam Ur1_n_8_pp.C9 = 9'd                 101;
defparam Ur1_n_8_pp.CA = 9'd                 141;
defparam Ur1_n_8_pp.CB = 9'd                 115;
defparam Ur1_n_8_pp.CC = 9'd                 197;
defparam Ur1_n_8_pp.CD = 9'd                 171;
defparam Ur1_n_8_pp.CE = 9'd                 211;
defparam Ur1_n_8_pp.CF = 9'd                 185;
assign lut_val_1_n_8_pp[10] = lut_val_1_n_8_pp[8];
assign lut_val_1_n_8_pp[9] = lut_val_1_n_8_pp[8];
wire [10:0] lut_val_1_n_9_pp;
rom_lut_r_cen Ur1_n_9_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_9_n[9],sym_res_7_n[9],sym_res_6_n[9],sym_res_5_n[9] } ), .data_out( lut_val_1_n_9_pp[8:0]) ) ;
 defparam Ur1_n_9_pp.DATA_WIDTH = 9;
defparam Ur1_n_9_pp.C0 = 9'd                   0;
defparam Ur1_n_9_pp.C1 = 9'd                 486;
defparam Ur1_n_9_pp.C2 = 9'd                  14;
defparam Ur1_n_9_pp.C3 = 9'd                 500;
defparam Ur1_n_9_pp.C4 = 9'd                  70;
defparam Ur1_n_9_pp.C5 = 9'd                  44;
defparam Ur1_n_9_pp.C6 = 9'd                  84;
defparam Ur1_n_9_pp.C7 = 9'd                  58;
defparam Ur1_n_9_pp.C8 = 9'd                 127;
defparam Ur1_n_9_pp.C9 = 9'd                 101;
defparam Ur1_n_9_pp.CA = 9'd                 141;
defparam Ur1_n_9_pp.CB = 9'd                 115;
defparam Ur1_n_9_pp.CC = 9'd                 197;
defparam Ur1_n_9_pp.CD = 9'd                 171;
defparam Ur1_n_9_pp.CE = 9'd                 211;
defparam Ur1_n_9_pp.CF = 9'd                 185;
assign lut_val_1_n_9_pp[10] = lut_val_1_n_9_pp[8];
assign lut_val_1_n_9_pp[9] = lut_val_1_n_9_pp[8];
wire [10:0] lut_val_1_n_10_pp;
rom_lut_r_cen Ur1_n_10_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_9_n[10],sym_res_7_n[10],sym_res_6_n[10],sym_res_5_n[10] } ), .data_out( lut_val_1_n_10_pp[8:0]) ) ;
 defparam Ur1_n_10_pp.DATA_WIDTH = 9;
defparam Ur1_n_10_pp.C0 = 9'd                   0;
defparam Ur1_n_10_pp.C1 = 9'd                 486;
defparam Ur1_n_10_pp.C2 = 9'd                  14;
defparam Ur1_n_10_pp.C3 = 9'd                 500;
defparam Ur1_n_10_pp.C4 = 9'd                  70;
defparam Ur1_n_10_pp.C5 = 9'd                  44;
defparam Ur1_n_10_pp.C6 = 9'd                  84;
defparam Ur1_n_10_pp.C7 = 9'd                  58;
defparam Ur1_n_10_pp.C8 = 9'd                 127;
defparam Ur1_n_10_pp.C9 = 9'd                 101;
defparam Ur1_n_10_pp.CA = 9'd                 141;
defparam Ur1_n_10_pp.CB = 9'd                 115;
defparam Ur1_n_10_pp.CC = 9'd                 197;
defparam Ur1_n_10_pp.CD = 9'd                 171;
defparam Ur1_n_10_pp.CE = 9'd                 211;
defparam Ur1_n_10_pp.CF = 9'd                 185;
assign lut_val_1_n_10_pp[10] = lut_val_1_n_10_pp[8];
assign lut_val_1_n_10_pp[9] = lut_val_1_n_10_pp[8];
wire [10:0] lut_val_1_n_11_pp;
rom_lut_r_cen Ur1_n_11_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_9_n[11],sym_res_7_n[11],sym_res_6_n[11],sym_res_5_n[11] } ), .data_out( lut_val_1_n_11_pp[8:0]) ) ;
 defparam Ur1_n_11_pp.DATA_WIDTH = 9;
defparam Ur1_n_11_pp.C0 = 9'd                   0;
defparam Ur1_n_11_pp.C1 = 9'd                  26;
defparam Ur1_n_11_pp.C2 = 9'd                 498;
defparam Ur1_n_11_pp.C3 = 9'd                  12;
defparam Ur1_n_11_pp.C4 = 9'd                 442;
defparam Ur1_n_11_pp.C5 = 9'd                 468;
defparam Ur1_n_11_pp.C6 = 9'd                 428;
defparam Ur1_n_11_pp.C7 = 9'd                 454;
defparam Ur1_n_11_pp.C8 = 9'd                 385;
defparam Ur1_n_11_pp.C9 = 9'd                 411;
defparam Ur1_n_11_pp.CA = 9'd                 371;
defparam Ur1_n_11_pp.CB = 9'd                 397;
defparam Ur1_n_11_pp.CC = 9'd                 315;
defparam Ur1_n_11_pp.CD = 9'd                 341;
defparam Ur1_n_11_pp.CE = 9'd                 301;
defparam Ur1_n_11_pp.CF = 9'd                 327;
assign lut_val_1_n_11_pp[10] = lut_val_1_n_11_pp[8];
assign lut_val_1_n_11_pp[9] = lut_val_1_n_11_pp[8];
wire [10:0] lut_val_2_n_0_pp;
rom_lut_r_cen Ur2_n_0_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_13_n[0],sym_res_12_n[0],sym_res_11_n[0],sym_res_10_n[0] } ), .data_out( lut_val_2_n_0_pp[10:0]) ) ;
 defparam Ur2_n_0_pp.DATA_WIDTH = 11;
defparam Ur2_n_0_pp.C0 = 11'd                   0;
defparam Ur2_n_0_pp.C1 = 11'd                  47;
defparam Ur2_n_0_pp.C2 = 11'd                1874;
defparam Ur2_n_0_pp.C3 = 11'd                1921;
defparam Ur2_n_0_pp.C4 = 11'd                  36;
defparam Ur2_n_0_pp.C5 = 11'd                  83;
defparam Ur2_n_0_pp.C6 = 11'd                1910;
defparam Ur2_n_0_pp.C7 = 11'd                1957;
defparam Ur2_n_0_pp.C8 = 11'd                1568;
defparam Ur2_n_0_pp.C9 = 11'd                1615;
defparam Ur2_n_0_pp.CA = 11'd                1394;
defparam Ur2_n_0_pp.CB = 11'd                1441;
defparam Ur2_n_0_pp.CC = 11'd                1604;
defparam Ur2_n_0_pp.CD = 11'd                1651;
defparam Ur2_n_0_pp.CE = 11'd                1430;
defparam Ur2_n_0_pp.CF = 11'd                1477;
wire [10:0] lut_val_2_n_1_pp;
rom_lut_r_cen Ur2_n_1_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_13_n[1],sym_res_12_n[1],sym_res_11_n[1],sym_res_10_n[1] } ), .data_out( lut_val_2_n_1_pp[10:0]) ) ;
 defparam Ur2_n_1_pp.DATA_WIDTH = 11;
defparam Ur2_n_1_pp.C0 = 11'd                   0;
defparam Ur2_n_1_pp.C1 = 11'd                  47;
defparam Ur2_n_1_pp.C2 = 11'd                1874;
defparam Ur2_n_1_pp.C3 = 11'd                1921;
defparam Ur2_n_1_pp.C4 = 11'd                  36;
defparam Ur2_n_1_pp.C5 = 11'd                  83;
defparam Ur2_n_1_pp.C6 = 11'd                1910;
defparam Ur2_n_1_pp.C7 = 11'd                1957;
defparam Ur2_n_1_pp.C8 = 11'd                1568;
defparam Ur2_n_1_pp.C9 = 11'd                1615;
defparam Ur2_n_1_pp.CA = 11'd                1394;
defparam Ur2_n_1_pp.CB = 11'd                1441;
defparam Ur2_n_1_pp.CC = 11'd                1604;
defparam Ur2_n_1_pp.CD = 11'd                1651;
defparam Ur2_n_1_pp.CE = 11'd                1430;
defparam Ur2_n_1_pp.CF = 11'd                1477;
wire [10:0] lut_val_2_n_2_pp;
rom_lut_r_cen Ur2_n_2_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_13_n[2],sym_res_12_n[2],sym_res_11_n[2],sym_res_10_n[2] } ), .data_out( lut_val_2_n_2_pp[10:0]) ) ;
 defparam Ur2_n_2_pp.DATA_WIDTH = 11;
defparam Ur2_n_2_pp.C0 = 11'd                   0;
defparam Ur2_n_2_pp.C1 = 11'd                  47;
defparam Ur2_n_2_pp.C2 = 11'd                1874;
defparam Ur2_n_2_pp.C3 = 11'd                1921;
defparam Ur2_n_2_pp.C4 = 11'd                  36;
defparam Ur2_n_2_pp.C5 = 11'd                  83;
defparam Ur2_n_2_pp.C6 = 11'd                1910;
defparam Ur2_n_2_pp.C7 = 11'd                1957;
defparam Ur2_n_2_pp.C8 = 11'd                1568;
defparam Ur2_n_2_pp.C9 = 11'd                1615;
defparam Ur2_n_2_pp.CA = 11'd                1394;
defparam Ur2_n_2_pp.CB = 11'd                1441;
defparam Ur2_n_2_pp.CC = 11'd                1604;
defparam Ur2_n_2_pp.CD = 11'd                1651;
defparam Ur2_n_2_pp.CE = 11'd                1430;
defparam Ur2_n_2_pp.CF = 11'd                1477;
wire [10:0] lut_val_2_n_3_pp;
rom_lut_r_cen Ur2_n_3_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_13_n[3],sym_res_12_n[3],sym_res_11_n[3],sym_res_10_n[3] } ), .data_out( lut_val_2_n_3_pp[10:0]) ) ;
 defparam Ur2_n_3_pp.DATA_WIDTH = 11;
defparam Ur2_n_3_pp.C0 = 11'd                   0;
defparam Ur2_n_3_pp.C1 = 11'd                  47;
defparam Ur2_n_3_pp.C2 = 11'd                1874;
defparam Ur2_n_3_pp.C3 = 11'd                1921;
defparam Ur2_n_3_pp.C4 = 11'd                  36;
defparam Ur2_n_3_pp.C5 = 11'd                  83;
defparam Ur2_n_3_pp.C6 = 11'd                1910;
defparam Ur2_n_3_pp.C7 = 11'd                1957;
defparam Ur2_n_3_pp.C8 = 11'd                1568;
defparam Ur2_n_3_pp.C9 = 11'd                1615;
defparam Ur2_n_3_pp.CA = 11'd                1394;
defparam Ur2_n_3_pp.CB = 11'd                1441;
defparam Ur2_n_3_pp.CC = 11'd                1604;
defparam Ur2_n_3_pp.CD = 11'd                1651;
defparam Ur2_n_3_pp.CE = 11'd                1430;
defparam Ur2_n_3_pp.CF = 11'd                1477;
wire [10:0] lut_val_2_n_4_pp;
rom_lut_r_cen Ur2_n_4_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_13_n[4],sym_res_12_n[4],sym_res_11_n[4],sym_res_10_n[4] } ), .data_out( lut_val_2_n_4_pp[10:0]) ) ;
 defparam Ur2_n_4_pp.DATA_WIDTH = 11;
defparam Ur2_n_4_pp.C0 = 11'd                   0;
defparam Ur2_n_4_pp.C1 = 11'd                  47;
defparam Ur2_n_4_pp.C2 = 11'd                1874;
defparam Ur2_n_4_pp.C3 = 11'd                1921;
defparam Ur2_n_4_pp.C4 = 11'd                  36;
defparam Ur2_n_4_pp.C5 = 11'd                  83;
defparam Ur2_n_4_pp.C6 = 11'd                1910;
defparam Ur2_n_4_pp.C7 = 11'd                1957;
defparam Ur2_n_4_pp.C8 = 11'd                1568;
defparam Ur2_n_4_pp.C9 = 11'd                1615;
defparam Ur2_n_4_pp.CA = 11'd                1394;
defparam Ur2_n_4_pp.CB = 11'd                1441;
defparam Ur2_n_4_pp.CC = 11'd                1604;
defparam Ur2_n_4_pp.CD = 11'd                1651;
defparam Ur2_n_4_pp.CE = 11'd                1430;
defparam Ur2_n_4_pp.CF = 11'd                1477;
wire [10:0] lut_val_2_n_5_pp;
rom_lut_r_cen Ur2_n_5_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_13_n[5],sym_res_12_n[5],sym_res_11_n[5],sym_res_10_n[5] } ), .data_out( lut_val_2_n_5_pp[10:0]) ) ;
 defparam Ur2_n_5_pp.DATA_WIDTH = 11;
defparam Ur2_n_5_pp.C0 = 11'd                   0;
defparam Ur2_n_5_pp.C1 = 11'd                  47;
defparam Ur2_n_5_pp.C2 = 11'd                1874;
defparam Ur2_n_5_pp.C3 = 11'd                1921;
defparam Ur2_n_5_pp.C4 = 11'd                  36;
defparam Ur2_n_5_pp.C5 = 11'd                  83;
defparam Ur2_n_5_pp.C6 = 11'd                1910;
defparam Ur2_n_5_pp.C7 = 11'd                1957;
defparam Ur2_n_5_pp.C8 = 11'd                1568;
defparam Ur2_n_5_pp.C9 = 11'd                1615;
defparam Ur2_n_5_pp.CA = 11'd                1394;
defparam Ur2_n_5_pp.CB = 11'd                1441;
defparam Ur2_n_5_pp.CC = 11'd                1604;
defparam Ur2_n_5_pp.CD = 11'd                1651;
defparam Ur2_n_5_pp.CE = 11'd                1430;
defparam Ur2_n_5_pp.CF = 11'd                1477;
wire [10:0] lut_val_2_n_6_pp;
rom_lut_r_cen Ur2_n_6_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_13_n[6],sym_res_12_n[6],sym_res_11_n[6],sym_res_10_n[6] } ), .data_out( lut_val_2_n_6_pp[10:0]) ) ;
 defparam Ur2_n_6_pp.DATA_WIDTH = 11;
defparam Ur2_n_6_pp.C0 = 11'd                   0;
defparam Ur2_n_6_pp.C1 = 11'd                  47;
defparam Ur2_n_6_pp.C2 = 11'd                1874;
defparam Ur2_n_6_pp.C3 = 11'd                1921;
defparam Ur2_n_6_pp.C4 = 11'd                  36;
defparam Ur2_n_6_pp.C5 = 11'd                  83;
defparam Ur2_n_6_pp.C6 = 11'd                1910;
defparam Ur2_n_6_pp.C7 = 11'd                1957;
defparam Ur2_n_6_pp.C8 = 11'd                1568;
defparam Ur2_n_6_pp.C9 = 11'd                1615;
defparam Ur2_n_6_pp.CA = 11'd                1394;
defparam Ur2_n_6_pp.CB = 11'd                1441;
defparam Ur2_n_6_pp.CC = 11'd                1604;
defparam Ur2_n_6_pp.CD = 11'd                1651;
defparam Ur2_n_6_pp.CE = 11'd                1430;
defparam Ur2_n_6_pp.CF = 11'd                1477;
wire [10:0] lut_val_2_n_7_pp;
rom_lut_r_cen Ur2_n_7_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_13_n[7],sym_res_12_n[7],sym_res_11_n[7],sym_res_10_n[7] } ), .data_out( lut_val_2_n_7_pp[10:0]) ) ;
 defparam Ur2_n_7_pp.DATA_WIDTH = 11;
defparam Ur2_n_7_pp.C0 = 11'd                   0;
defparam Ur2_n_7_pp.C1 = 11'd                  47;
defparam Ur2_n_7_pp.C2 = 11'd                1874;
defparam Ur2_n_7_pp.C3 = 11'd                1921;
defparam Ur2_n_7_pp.C4 = 11'd                  36;
defparam Ur2_n_7_pp.C5 = 11'd                  83;
defparam Ur2_n_7_pp.C6 = 11'd                1910;
defparam Ur2_n_7_pp.C7 = 11'd                1957;
defparam Ur2_n_7_pp.C8 = 11'd                1568;
defparam Ur2_n_7_pp.C9 = 11'd                1615;
defparam Ur2_n_7_pp.CA = 11'd                1394;
defparam Ur2_n_7_pp.CB = 11'd                1441;
defparam Ur2_n_7_pp.CC = 11'd                1604;
defparam Ur2_n_7_pp.CD = 11'd                1651;
defparam Ur2_n_7_pp.CE = 11'd                1430;
defparam Ur2_n_7_pp.CF = 11'd                1477;
wire [10:0] lut_val_2_n_8_pp;
rom_lut_r_cen Ur2_n_8_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_13_n[8],sym_res_12_n[8],sym_res_11_n[8],sym_res_10_n[8] } ), .data_out( lut_val_2_n_8_pp[10:0]) ) ;
 defparam Ur2_n_8_pp.DATA_WIDTH = 11;
defparam Ur2_n_8_pp.C0 = 11'd                   0;
defparam Ur2_n_8_pp.C1 = 11'd                  47;
defparam Ur2_n_8_pp.C2 = 11'd                1874;
defparam Ur2_n_8_pp.C3 = 11'd                1921;
defparam Ur2_n_8_pp.C4 = 11'd                  36;
defparam Ur2_n_8_pp.C5 = 11'd                  83;
defparam Ur2_n_8_pp.C6 = 11'd                1910;
defparam Ur2_n_8_pp.C7 = 11'd                1957;
defparam Ur2_n_8_pp.C8 = 11'd                1568;
defparam Ur2_n_8_pp.C9 = 11'd                1615;
defparam Ur2_n_8_pp.CA = 11'd                1394;
defparam Ur2_n_8_pp.CB = 11'd                1441;
defparam Ur2_n_8_pp.CC = 11'd                1604;
defparam Ur2_n_8_pp.CD = 11'd                1651;
defparam Ur2_n_8_pp.CE = 11'd                1430;
defparam Ur2_n_8_pp.CF = 11'd                1477;
wire [10:0] lut_val_2_n_9_pp;
rom_lut_r_cen Ur2_n_9_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_13_n[9],sym_res_12_n[9],sym_res_11_n[9],sym_res_10_n[9] } ), .data_out( lut_val_2_n_9_pp[10:0]) ) ;
 defparam Ur2_n_9_pp.DATA_WIDTH = 11;
defparam Ur2_n_9_pp.C0 = 11'd                   0;
defparam Ur2_n_9_pp.C1 = 11'd                  47;
defparam Ur2_n_9_pp.C2 = 11'd                1874;
defparam Ur2_n_9_pp.C3 = 11'd                1921;
defparam Ur2_n_9_pp.C4 = 11'd                  36;
defparam Ur2_n_9_pp.C5 = 11'd                  83;
defparam Ur2_n_9_pp.C6 = 11'd                1910;
defparam Ur2_n_9_pp.C7 = 11'd                1957;
defparam Ur2_n_9_pp.C8 = 11'd                1568;
defparam Ur2_n_9_pp.C9 = 11'd                1615;
defparam Ur2_n_9_pp.CA = 11'd                1394;
defparam Ur2_n_9_pp.CB = 11'd                1441;
defparam Ur2_n_9_pp.CC = 11'd                1604;
defparam Ur2_n_9_pp.CD = 11'd                1651;
defparam Ur2_n_9_pp.CE = 11'd                1430;
defparam Ur2_n_9_pp.CF = 11'd                1477;
wire [10:0] lut_val_2_n_10_pp;
rom_lut_r_cen Ur2_n_10_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_13_n[10],sym_res_12_n[10],sym_res_11_n[10],sym_res_10_n[10] } ), .data_out( lut_val_2_n_10_pp[10:0]) ) ;
 defparam Ur2_n_10_pp.DATA_WIDTH = 11;
defparam Ur2_n_10_pp.C0 = 11'd                   0;
defparam Ur2_n_10_pp.C1 = 11'd                  47;
defparam Ur2_n_10_pp.C2 = 11'd                1874;
defparam Ur2_n_10_pp.C3 = 11'd                1921;
defparam Ur2_n_10_pp.C4 = 11'd                  36;
defparam Ur2_n_10_pp.C5 = 11'd                  83;
defparam Ur2_n_10_pp.C6 = 11'd                1910;
defparam Ur2_n_10_pp.C7 = 11'd                1957;
defparam Ur2_n_10_pp.C8 = 11'd                1568;
defparam Ur2_n_10_pp.C9 = 11'd                1615;
defparam Ur2_n_10_pp.CA = 11'd                1394;
defparam Ur2_n_10_pp.CB = 11'd                1441;
defparam Ur2_n_10_pp.CC = 11'd                1604;
defparam Ur2_n_10_pp.CD = 11'd                1651;
defparam Ur2_n_10_pp.CE = 11'd                1430;
defparam Ur2_n_10_pp.CF = 11'd                1477;
wire [10:0] lut_val_2_n_11_pp;
rom_lut_r_cen Ur2_n_11_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {sym_res_13_n[11],sym_res_12_n[11],sym_res_11_n[11],sym_res_10_n[11] } ), .data_out( lut_val_2_n_11_pp[10:0]) ) ;
 defparam Ur2_n_11_pp.DATA_WIDTH = 11;
defparam Ur2_n_11_pp.C0 = 11'd                   0;
defparam Ur2_n_11_pp.C1 = 11'd                2001;
defparam Ur2_n_11_pp.C2 = 11'd                 174;
defparam Ur2_n_11_pp.C3 = 11'd                 127;
defparam Ur2_n_11_pp.C4 = 11'd                2012;
defparam Ur2_n_11_pp.C5 = 11'd                1965;
defparam Ur2_n_11_pp.C6 = 11'd                 138;
defparam Ur2_n_11_pp.C7 = 11'd                  91;
defparam Ur2_n_11_pp.C8 = 11'd                 480;
defparam Ur2_n_11_pp.C9 = 11'd                 433;
defparam Ur2_n_11_pp.CA = 11'd                 654;
defparam Ur2_n_11_pp.CB = 11'd                 607;
defparam Ur2_n_11_pp.CC = 11'd                 444;
defparam Ur2_n_11_pp.CD = 11'd                 397;
defparam Ur2_n_11_pp.CE = 11'd                 618;
defparam Ur2_n_11_pp.CF = 11'd                 571;
wire [10:0] lut_val_3_n_0_pp;
rom_lut_r_cen Ur3_n_0_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {addr_low,addr_low,sym_res_15_n[0],sym_res_14_n[0] } ), .data_out( lut_val_3_n_0_pp[10:0]) ) ;
 defparam Ur3_n_0_pp.DATA_WIDTH = 11;
defparam Ur3_n_0_pp.C0 = 11'd                   0;
defparam Ur3_n_0_pp.C1 = 11'd                1429;
defparam Ur3_n_0_pp.C2 = 11'd                1023;
defparam Ur3_n_0_pp.C3 = 11'd                 404;
defparam Ur3_n_0_pp.C4 = 11'd                   0;
defparam Ur3_n_0_pp.C5 = 11'd                1429;
defparam Ur3_n_0_pp.C6 = 11'd                1023;
defparam Ur3_n_0_pp.C7 = 11'd                 404;
defparam Ur3_n_0_pp.C8 = 11'd                   0;
defparam Ur3_n_0_pp.C9 = 11'd                1429;
defparam Ur3_n_0_pp.CA = 11'd                1023;
defparam Ur3_n_0_pp.CB = 11'd                 404;
defparam Ur3_n_0_pp.CC = 11'd                   0;
defparam Ur3_n_0_pp.CD = 11'd                1429;
defparam Ur3_n_0_pp.CE = 11'd                1023;
defparam Ur3_n_0_pp.CF = 11'd                 404;
wire [10:0] lut_val_3_n_1_pp;
rom_lut_r_cen Ur3_n_1_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {addr_low,addr_low,sym_res_15_n[1],sym_res_14_n[1] } ), .data_out( lut_val_3_n_1_pp[10:0]) ) ;
 defparam Ur3_n_1_pp.DATA_WIDTH = 11;
defparam Ur3_n_1_pp.C0 = 11'd                   0;
defparam Ur3_n_1_pp.C1 = 11'd                1429;
defparam Ur3_n_1_pp.C2 = 11'd                1023;
defparam Ur3_n_1_pp.C3 = 11'd                 404;
defparam Ur3_n_1_pp.C4 = 11'd                   0;
defparam Ur3_n_1_pp.C5 = 11'd                1429;
defparam Ur3_n_1_pp.C6 = 11'd                1023;
defparam Ur3_n_1_pp.C7 = 11'd                 404;
defparam Ur3_n_1_pp.C8 = 11'd                   0;
defparam Ur3_n_1_pp.C9 = 11'd                1429;
defparam Ur3_n_1_pp.CA = 11'd                1023;
defparam Ur3_n_1_pp.CB = 11'd                 404;
defparam Ur3_n_1_pp.CC = 11'd                   0;
defparam Ur3_n_1_pp.CD = 11'd                1429;
defparam Ur3_n_1_pp.CE = 11'd                1023;
defparam Ur3_n_1_pp.CF = 11'd                 404;
wire [10:0] lut_val_3_n_2_pp;
rom_lut_r_cen Ur3_n_2_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {addr_low,addr_low,sym_res_15_n[2],sym_res_14_n[2] } ), .data_out( lut_val_3_n_2_pp[10:0]) ) ;
 defparam Ur3_n_2_pp.DATA_WIDTH = 11;
defparam Ur3_n_2_pp.C0 = 11'd                   0;
defparam Ur3_n_2_pp.C1 = 11'd                1429;
defparam Ur3_n_2_pp.C2 = 11'd                1023;
defparam Ur3_n_2_pp.C3 = 11'd                 404;
defparam Ur3_n_2_pp.C4 = 11'd                   0;
defparam Ur3_n_2_pp.C5 = 11'd                1429;
defparam Ur3_n_2_pp.C6 = 11'd                1023;
defparam Ur3_n_2_pp.C7 = 11'd                 404;
defparam Ur3_n_2_pp.C8 = 11'd                   0;
defparam Ur3_n_2_pp.C9 = 11'd                1429;
defparam Ur3_n_2_pp.CA = 11'd                1023;
defparam Ur3_n_2_pp.CB = 11'd                 404;
defparam Ur3_n_2_pp.CC = 11'd                   0;
defparam Ur3_n_2_pp.CD = 11'd                1429;
defparam Ur3_n_2_pp.CE = 11'd                1023;
defparam Ur3_n_2_pp.CF = 11'd                 404;
wire [10:0] lut_val_3_n_3_pp;
rom_lut_r_cen Ur3_n_3_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {addr_low,addr_low,sym_res_15_n[3],sym_res_14_n[3] } ), .data_out( lut_val_3_n_3_pp[10:0]) ) ;
 defparam Ur3_n_3_pp.DATA_WIDTH = 11;
defparam Ur3_n_3_pp.C0 = 11'd                   0;
defparam Ur3_n_3_pp.C1 = 11'd                1429;
defparam Ur3_n_3_pp.C2 = 11'd                1023;
defparam Ur3_n_3_pp.C3 = 11'd                 404;
defparam Ur3_n_3_pp.C4 = 11'd                   0;
defparam Ur3_n_3_pp.C5 = 11'd                1429;
defparam Ur3_n_3_pp.C6 = 11'd                1023;
defparam Ur3_n_3_pp.C7 = 11'd                 404;
defparam Ur3_n_3_pp.C8 = 11'd                   0;
defparam Ur3_n_3_pp.C9 = 11'd                1429;
defparam Ur3_n_3_pp.CA = 11'd                1023;
defparam Ur3_n_3_pp.CB = 11'd                 404;
defparam Ur3_n_3_pp.CC = 11'd                   0;
defparam Ur3_n_3_pp.CD = 11'd                1429;
defparam Ur3_n_3_pp.CE = 11'd                1023;
defparam Ur3_n_3_pp.CF = 11'd                 404;
wire [10:0] lut_val_3_n_4_pp;
rom_lut_r_cen Ur3_n_4_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {addr_low,addr_low,sym_res_15_n[4],sym_res_14_n[4] } ), .data_out( lut_val_3_n_4_pp[10:0]) ) ;
 defparam Ur3_n_4_pp.DATA_WIDTH = 11;
defparam Ur3_n_4_pp.C0 = 11'd                   0;
defparam Ur3_n_4_pp.C1 = 11'd                1429;
defparam Ur3_n_4_pp.C2 = 11'd                1023;
defparam Ur3_n_4_pp.C3 = 11'd                 404;
defparam Ur3_n_4_pp.C4 = 11'd                   0;
defparam Ur3_n_4_pp.C5 = 11'd                1429;
defparam Ur3_n_4_pp.C6 = 11'd                1023;
defparam Ur3_n_4_pp.C7 = 11'd                 404;
defparam Ur3_n_4_pp.C8 = 11'd                   0;
defparam Ur3_n_4_pp.C9 = 11'd                1429;
defparam Ur3_n_4_pp.CA = 11'd                1023;
defparam Ur3_n_4_pp.CB = 11'd                 404;
defparam Ur3_n_4_pp.CC = 11'd                   0;
defparam Ur3_n_4_pp.CD = 11'd                1429;
defparam Ur3_n_4_pp.CE = 11'd                1023;
defparam Ur3_n_4_pp.CF = 11'd                 404;
wire [10:0] lut_val_3_n_5_pp;
rom_lut_r_cen Ur3_n_5_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {addr_low,addr_low,sym_res_15_n[5],sym_res_14_n[5] } ), .data_out( lut_val_3_n_5_pp[10:0]) ) ;
 defparam Ur3_n_5_pp.DATA_WIDTH = 11;
defparam Ur3_n_5_pp.C0 = 11'd                   0;
defparam Ur3_n_5_pp.C1 = 11'd                1429;
defparam Ur3_n_5_pp.C2 = 11'd                1023;
defparam Ur3_n_5_pp.C3 = 11'd                 404;
defparam Ur3_n_5_pp.C4 = 11'd                   0;
defparam Ur3_n_5_pp.C5 = 11'd                1429;
defparam Ur3_n_5_pp.C6 = 11'd                1023;
defparam Ur3_n_5_pp.C7 = 11'd                 404;
defparam Ur3_n_5_pp.C8 = 11'd                   0;
defparam Ur3_n_5_pp.C9 = 11'd                1429;
defparam Ur3_n_5_pp.CA = 11'd                1023;
defparam Ur3_n_5_pp.CB = 11'd                 404;
defparam Ur3_n_5_pp.CC = 11'd                   0;
defparam Ur3_n_5_pp.CD = 11'd                1429;
defparam Ur3_n_5_pp.CE = 11'd                1023;
defparam Ur3_n_5_pp.CF = 11'd                 404;
wire [10:0] lut_val_3_n_6_pp;
rom_lut_r_cen Ur3_n_6_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {addr_low,addr_low,sym_res_15_n[6],sym_res_14_n[6] } ), .data_out( lut_val_3_n_6_pp[10:0]) ) ;
 defparam Ur3_n_6_pp.DATA_WIDTH = 11;
defparam Ur3_n_6_pp.C0 = 11'd                   0;
defparam Ur3_n_6_pp.C1 = 11'd                1429;
defparam Ur3_n_6_pp.C2 = 11'd                1023;
defparam Ur3_n_6_pp.C3 = 11'd                 404;
defparam Ur3_n_6_pp.C4 = 11'd                   0;
defparam Ur3_n_6_pp.C5 = 11'd                1429;
defparam Ur3_n_6_pp.C6 = 11'd                1023;
defparam Ur3_n_6_pp.C7 = 11'd                 404;
defparam Ur3_n_6_pp.C8 = 11'd                   0;
defparam Ur3_n_6_pp.C9 = 11'd                1429;
defparam Ur3_n_6_pp.CA = 11'd                1023;
defparam Ur3_n_6_pp.CB = 11'd                 404;
defparam Ur3_n_6_pp.CC = 11'd                   0;
defparam Ur3_n_6_pp.CD = 11'd                1429;
defparam Ur3_n_6_pp.CE = 11'd                1023;
defparam Ur3_n_6_pp.CF = 11'd                 404;
wire [10:0] lut_val_3_n_7_pp;
rom_lut_r_cen Ur3_n_7_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {addr_low,addr_low,sym_res_15_n[7],sym_res_14_n[7] } ), .data_out( lut_val_3_n_7_pp[10:0]) ) ;
 defparam Ur3_n_7_pp.DATA_WIDTH = 11;
defparam Ur3_n_7_pp.C0 = 11'd                   0;
defparam Ur3_n_7_pp.C1 = 11'd                1429;
defparam Ur3_n_7_pp.C2 = 11'd                1023;
defparam Ur3_n_7_pp.C3 = 11'd                 404;
defparam Ur3_n_7_pp.C4 = 11'd                   0;
defparam Ur3_n_7_pp.C5 = 11'd                1429;
defparam Ur3_n_7_pp.C6 = 11'd                1023;
defparam Ur3_n_7_pp.C7 = 11'd                 404;
defparam Ur3_n_7_pp.C8 = 11'd                   0;
defparam Ur3_n_7_pp.C9 = 11'd                1429;
defparam Ur3_n_7_pp.CA = 11'd                1023;
defparam Ur3_n_7_pp.CB = 11'd                 404;
defparam Ur3_n_7_pp.CC = 11'd                   0;
defparam Ur3_n_7_pp.CD = 11'd                1429;
defparam Ur3_n_7_pp.CE = 11'd                1023;
defparam Ur3_n_7_pp.CF = 11'd                 404;
wire [10:0] lut_val_3_n_8_pp;
rom_lut_r_cen Ur3_n_8_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {addr_low,addr_low,sym_res_15_n[8],sym_res_14_n[8] } ), .data_out( lut_val_3_n_8_pp[10:0]) ) ;
 defparam Ur3_n_8_pp.DATA_WIDTH = 11;
defparam Ur3_n_8_pp.C0 = 11'd                   0;
defparam Ur3_n_8_pp.C1 = 11'd                1429;
defparam Ur3_n_8_pp.C2 = 11'd                1023;
defparam Ur3_n_8_pp.C3 = 11'd                 404;
defparam Ur3_n_8_pp.C4 = 11'd                   0;
defparam Ur3_n_8_pp.C5 = 11'd                1429;
defparam Ur3_n_8_pp.C6 = 11'd                1023;
defparam Ur3_n_8_pp.C7 = 11'd                 404;
defparam Ur3_n_8_pp.C8 = 11'd                   0;
defparam Ur3_n_8_pp.C9 = 11'd                1429;
defparam Ur3_n_8_pp.CA = 11'd                1023;
defparam Ur3_n_8_pp.CB = 11'd                 404;
defparam Ur3_n_8_pp.CC = 11'd                   0;
defparam Ur3_n_8_pp.CD = 11'd                1429;
defparam Ur3_n_8_pp.CE = 11'd                1023;
defparam Ur3_n_8_pp.CF = 11'd                 404;
wire [10:0] lut_val_3_n_9_pp;
rom_lut_r_cen Ur3_n_9_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {addr_low,addr_low,sym_res_15_n[9],sym_res_14_n[9] } ), .data_out( lut_val_3_n_9_pp[10:0]) ) ;
 defparam Ur3_n_9_pp.DATA_WIDTH = 11;
defparam Ur3_n_9_pp.C0 = 11'd                   0;
defparam Ur3_n_9_pp.C1 = 11'd                1429;
defparam Ur3_n_9_pp.C2 = 11'd                1023;
defparam Ur3_n_9_pp.C3 = 11'd                 404;
defparam Ur3_n_9_pp.C4 = 11'd                   0;
defparam Ur3_n_9_pp.C5 = 11'd                1429;
defparam Ur3_n_9_pp.C6 = 11'd                1023;
defparam Ur3_n_9_pp.C7 = 11'd                 404;
defparam Ur3_n_9_pp.C8 = 11'd                   0;
defparam Ur3_n_9_pp.C9 = 11'd                1429;
defparam Ur3_n_9_pp.CA = 11'd                1023;
defparam Ur3_n_9_pp.CB = 11'd                 404;
defparam Ur3_n_9_pp.CC = 11'd                   0;
defparam Ur3_n_9_pp.CD = 11'd                1429;
defparam Ur3_n_9_pp.CE = 11'd                1023;
defparam Ur3_n_9_pp.CF = 11'd                 404;
wire [10:0] lut_val_3_n_10_pp;
rom_lut_r_cen Ur3_n_10_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {addr_low,addr_low,sym_res_15_n[10],sym_res_14_n[10] } ), .data_out( lut_val_3_n_10_pp[10:0]) ) ;
 defparam Ur3_n_10_pp.DATA_WIDTH = 11;
defparam Ur3_n_10_pp.C0 = 11'd                   0;
defparam Ur3_n_10_pp.C1 = 11'd                1429;
defparam Ur3_n_10_pp.C2 = 11'd                1023;
defparam Ur3_n_10_pp.C3 = 11'd                 404;
defparam Ur3_n_10_pp.C4 = 11'd                   0;
defparam Ur3_n_10_pp.C5 = 11'd                1429;
defparam Ur3_n_10_pp.C6 = 11'd                1023;
defparam Ur3_n_10_pp.C7 = 11'd                 404;
defparam Ur3_n_10_pp.C8 = 11'd                   0;
defparam Ur3_n_10_pp.C9 = 11'd                1429;
defparam Ur3_n_10_pp.CA = 11'd                1023;
defparam Ur3_n_10_pp.CB = 11'd                 404;
defparam Ur3_n_10_pp.CC = 11'd                   0;
defparam Ur3_n_10_pp.CD = 11'd                1429;
defparam Ur3_n_10_pp.CE = 11'd                1023;
defparam Ur3_n_10_pp.CF = 11'd                 404;
wire [10:0] lut_val_3_n_11_pp;
rom_lut_r_cen Ur3_n_11_pp (.clk(clk),.gclk_en(clk_en),.addr_in( {addr_low,addr_low,sym_res_15_n[11],sym_res_14_n[11] } ), .data_out( lut_val_3_n_11_pp[10:0]) ) ;
 defparam Ur3_n_11_pp.DATA_WIDTH = 11;
defparam Ur3_n_11_pp.C0 = 11'd                   0;
defparam Ur3_n_11_pp.C1 = 11'd                 619;
defparam Ur3_n_11_pp.C2 = 11'd                1025;
defparam Ur3_n_11_pp.C3 = 11'd                1644;
defparam Ur3_n_11_pp.C4 = 11'd                   0;
defparam Ur3_n_11_pp.C5 = 11'd                 619;
defparam Ur3_n_11_pp.C6 = 11'd                1025;
defparam Ur3_n_11_pp.C7 = 11'd                1644;
defparam Ur3_n_11_pp.C8 = 11'd                   0;
defparam Ur3_n_11_pp.C9 = 11'd                 619;
defparam Ur3_n_11_pp.CA = 11'd                1025;
defparam Ur3_n_11_pp.CB = 11'd                1644;
defparam Ur3_n_11_pp.CC = 11'd                   0;
defparam Ur3_n_11_pp.CD = 11'd                 619;
defparam Ur3_n_11_pp.CE = 11'd                1025;
defparam Ur3_n_11_pp.CF = 11'd                1644;
wire [21:0] lut_0_bit_0_fill;
wire [21:0] lut_0_bit_1_fill;
wire [21:0] lut_0_bit_2_fill;
wire [21:0] lut_0_bit_3_fill;
wire [21:0] lut_0_bit_4_fill;
wire [21:0] lut_0_bit_5_fill;
wire [21:0] lut_0_bit_6_fill;
wire [21:0] lut_0_bit_7_fill;
wire [21:0] lut_0_bit_8_fill;
wire [21:0] lut_0_bit_9_fill;
wire [21:0] lut_0_bit_10_fill;
wire [21:0] lut_0_bit_11_fill;
assign lut_0_bit_0_fill = {lut_val_0_n_0_pp[10], lut_val_0_n_0_pp[10], lut_val_0_n_0_pp[10], lut_val_0_n_0_pp[10], lut_val_0_n_0_pp[10], lut_val_0_n_0_pp[10], lut_val_0_n_0_pp[10], lut_val_0_n_0_pp[10], lut_val_0_n_0_pp[10], lut_val_0_n_0_pp[10], lut_val_0_n_0_pp[10],  lut_val_0_n_0_pp };
assign lut_0_bit_1_fill = {lut_val_0_n_1_pp[10], lut_val_0_n_1_pp[10], lut_val_0_n_1_pp[10], lut_val_0_n_1_pp[10], lut_val_0_n_1_pp[10], lut_val_0_n_1_pp[10], lut_val_0_n_1_pp[10], lut_val_0_n_1_pp[10], lut_val_0_n_1_pp[10], lut_val_0_n_1_pp[10],  lut_val_0_n_1_pp, 1'd0 };
assign lut_0_bit_2_fill = {lut_val_0_n_2_pp[10], lut_val_0_n_2_pp[10], lut_val_0_n_2_pp[10], lut_val_0_n_2_pp[10], lut_val_0_n_2_pp[10], lut_val_0_n_2_pp[10], lut_val_0_n_2_pp[10], lut_val_0_n_2_pp[10], lut_val_0_n_2_pp[10],  lut_val_0_n_2_pp, 2'd0 };
assign lut_0_bit_3_fill = {lut_val_0_n_3_pp[10], lut_val_0_n_3_pp[10], lut_val_0_n_3_pp[10], lut_val_0_n_3_pp[10], lut_val_0_n_3_pp[10], lut_val_0_n_3_pp[10], lut_val_0_n_3_pp[10], lut_val_0_n_3_pp[10],  lut_val_0_n_3_pp, 3'd0 };
assign lut_0_bit_4_fill = {lut_val_0_n_4_pp[10], lut_val_0_n_4_pp[10], lut_val_0_n_4_pp[10], lut_val_0_n_4_pp[10], lut_val_0_n_4_pp[10], lut_val_0_n_4_pp[10], lut_val_0_n_4_pp[10],  lut_val_0_n_4_pp, 4'd0 };
assign lut_0_bit_5_fill = {lut_val_0_n_5_pp[10], lut_val_0_n_5_pp[10], lut_val_0_n_5_pp[10], lut_val_0_n_5_pp[10], lut_val_0_n_5_pp[10], lut_val_0_n_5_pp[10],  lut_val_0_n_5_pp, 5'd0 };
assign lut_0_bit_6_fill = {lut_val_0_n_6_pp[10], lut_val_0_n_6_pp[10], lut_val_0_n_6_pp[10], lut_val_0_n_6_pp[10], lut_val_0_n_6_pp[10],  lut_val_0_n_6_pp, 6'd0 };
assign lut_0_bit_7_fill = {lut_val_0_n_7_pp[10], lut_val_0_n_7_pp[10], lut_val_0_n_7_pp[10], lut_val_0_n_7_pp[10],  lut_val_0_n_7_pp, 7'd0 };
assign lut_0_bit_8_fill = {lut_val_0_n_8_pp[10], lut_val_0_n_8_pp[10], lut_val_0_n_8_pp[10],  lut_val_0_n_8_pp, 8'd0 };
assign lut_0_bit_9_fill = {lut_val_0_n_9_pp[10], lut_val_0_n_9_pp[10],  lut_val_0_n_9_pp, 9'd0 };
assign lut_0_bit_10_fill = {lut_val_0_n_10_pp[10],  lut_val_0_n_10_pp, 10'd0 };
assign lut_0_bit_11_fill = { lut_val_0_n_11_pp, 11'd0 };
wire [22:0] tree_0_pp_l_0_n_0_n;
sadd_lpm_cen Uadd_0_lut_l_0_n_0_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_0_bit_0_fill), .bin(lut_0_bit_1_fill), .res(tree_0_pp_l_0_n_0_n) );
defparam Uadd_0_lut_l_0_n_0_n.IN_WIDTH = 22;
defparam Uadd_0_lut_l_0_n_0_n.PIPE_DEPTH = 3;
wire [22:0] tree_0_pp_l_0_n_1_n;
sadd_lpm_cen Uadd_0_lut_l_0_n_1_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_0_bit_2_fill), .bin(lut_0_bit_3_fill), .res(tree_0_pp_l_0_n_1_n) );
defparam Uadd_0_lut_l_0_n_1_n.IN_WIDTH = 22;
defparam Uadd_0_lut_l_0_n_1_n.PIPE_DEPTH = 3;
wire [22:0] tree_0_pp_l_0_n_2_n;
sadd_lpm_cen Uadd_0_lut_l_0_n_2_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_0_bit_4_fill), .bin(lut_0_bit_5_fill), .res(tree_0_pp_l_0_n_2_n) );
defparam Uadd_0_lut_l_0_n_2_n.IN_WIDTH = 22;
defparam Uadd_0_lut_l_0_n_2_n.PIPE_DEPTH = 3;
wire [22:0] tree_0_pp_l_0_n_3_n;
sadd_lpm_cen Uadd_0_lut_l_0_n_3_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_0_bit_6_fill), .bin(lut_0_bit_7_fill), .res(tree_0_pp_l_0_n_3_n) );
defparam Uadd_0_lut_l_0_n_3_n.IN_WIDTH = 22;
defparam Uadd_0_lut_l_0_n_3_n.PIPE_DEPTH = 3;
wire [22:0] tree_0_pp_l_0_n_4_n;
sadd_lpm_cen Uadd_0_lut_l_0_n_4_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_0_bit_8_fill), .bin(lut_0_bit_9_fill), .res(tree_0_pp_l_0_n_4_n) );
defparam Uadd_0_lut_l_0_n_4_n.IN_WIDTH = 22;
defparam Uadd_0_lut_l_0_n_4_n.PIPE_DEPTH = 3;
wire [22:0] tree_0_pp_l_0_n_5_n;
sadd_lpm_cen Uadd_0_lut_l_0_n_5_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_0_bit_10_fill), .bin(lut_0_bit_11_fill), .res(tree_0_pp_l_0_n_5_n) );
defparam Uadd_0_lut_l_0_n_5_n.IN_WIDTH = 22;
defparam Uadd_0_lut_l_0_n_5_n.PIPE_DEPTH = 3;
wire [23:0] tree_0_pp_l_1_n_0_n;
sadd_lpm_cen Uadd_0_lut_l_1_n_0_n (.clk(clk),  .gclk_en(clk_en), .ain(tree_0_pp_l_0_n_0_n), .bin(tree_0_pp_l_0_n_1_n), .res(tree_0_pp_l_1_n_0_n) );
defparam Uadd_0_lut_l_1_n_0_n.IN_WIDTH = 23;
defparam Uadd_0_lut_l_1_n_0_n.PIPE_DEPTH = 3;
wire [23:0] tree_0_pp_l_1_n_1_n;
sadd_lpm_cen Uadd_0_lut_l_1_n_1_n (.clk(clk),  .gclk_en(clk_en), .ain(tree_0_pp_l_0_n_2_n), .bin(tree_0_pp_l_0_n_3_n), .res(tree_0_pp_l_1_n_1_n) );
defparam Uadd_0_lut_l_1_n_1_n.IN_WIDTH = 23;
defparam Uadd_0_lut_l_1_n_1_n.PIPE_DEPTH = 3;
wire [23:0] tree_0_pp_l_1_n_2_n;
sadd_lpm_cen Uadd_0_lut_l_1_n_2_n (.clk(clk),  .gclk_en(clk_en), .ain(tree_0_pp_l_0_n_4_n), .bin(tree_0_pp_l_0_n_5_n), .res(tree_0_pp_l_1_n_2_n) );
defparam Uadd_0_lut_l_1_n_2_n.IN_WIDTH = 23;
defparam Uadd_0_lut_l_1_n_2_n.PIPE_DEPTH = 3;
wire [24:0] tree_0_pp_l_2_n_0_n;
sadd_lpm_cen Uadd_0_lut_l_2_n_0_n (.clk(clk),  .gclk_en(clk_en), .ain(tree_0_pp_l_1_n_0_n), .bin(tree_0_pp_l_1_n_1_n), .res(tree_0_pp_l_2_n_0_n) );
defparam Uadd_0_lut_l_2_n_0_n.IN_WIDTH = 24;
defparam Uadd_0_lut_l_2_n_0_n.PIPE_DEPTH = 3;
wire [24:0] tree_0_pp_l_2_n_1_n;
sadd_lpm_cen Uadd_0_lut_l_2_n_1_n (.clk(clk),  .gclk_en(clk_en), .ain(tree_0_pp_l_1_n_2_n), .bin(24'd0), .res(tree_0_pp_l_2_n_1_n) );
defparam Uadd_0_lut_l_2_n_1_n.IN_WIDTH = 24;
defparam Uadd_0_lut_l_2_n_1_n.PIPE_DEPTH = 3;
wire [25:0] tree_0_pp_l_3_n_0_n;
sadd_lpm_cen Uadd_0_lut_l_3_n_0_n (.clk(clk),  .gclk_en(clk_en), .ain(tree_0_pp_l_2_n_0_n), .bin(tree_0_pp_l_2_n_1_n), .res(tree_0_pp_l_3_n_0_n) );
defparam Uadd_0_lut_l_3_n_0_n.IN_WIDTH = 25;
defparam Uadd_0_lut_l_3_n_0_n.PIPE_DEPTH = 3;
wire [25:0] lut_val_0_n;
assign lut_val_0_n=tree_0_pp_l_3_n_0_n;
wire [21:0] lut_1_bit_0_fill;
wire [21:0] lut_1_bit_1_fill;
wire [21:0] lut_1_bit_2_fill;
wire [21:0] lut_1_bit_3_fill;
wire [21:0] lut_1_bit_4_fill;
wire [21:0] lut_1_bit_5_fill;
wire [21:0] lut_1_bit_6_fill;
wire [21:0] lut_1_bit_7_fill;
wire [21:0] lut_1_bit_8_fill;
wire [21:0] lut_1_bit_9_fill;
wire [21:0] lut_1_bit_10_fill;
wire [21:0] lut_1_bit_11_fill;
assign lut_1_bit_0_fill = {lut_val_1_n_0_pp[10], lut_val_1_n_0_pp[10], lut_val_1_n_0_pp[10], lut_val_1_n_0_pp[10], lut_val_1_n_0_pp[10], lut_val_1_n_0_pp[10], lut_val_1_n_0_pp[10], lut_val_1_n_0_pp[10], lut_val_1_n_0_pp[10], lut_val_1_n_0_pp[10], lut_val_1_n_0_pp[10],  lut_val_1_n_0_pp };
assign lut_1_bit_1_fill = {lut_val_1_n_1_pp[10], lut_val_1_n_1_pp[10], lut_val_1_n_1_pp[10], lut_val_1_n_1_pp[10], lut_val_1_n_1_pp[10], lut_val_1_n_1_pp[10], lut_val_1_n_1_pp[10], lut_val_1_n_1_pp[10], lut_val_1_n_1_pp[10], lut_val_1_n_1_pp[10],  lut_val_1_n_1_pp, 1'd0 };
assign lut_1_bit_2_fill = {lut_val_1_n_2_pp[10], lut_val_1_n_2_pp[10], lut_val_1_n_2_pp[10], lut_val_1_n_2_pp[10], lut_val_1_n_2_pp[10], lut_val_1_n_2_pp[10], lut_val_1_n_2_pp[10], lut_val_1_n_2_pp[10], lut_val_1_n_2_pp[10],  lut_val_1_n_2_pp, 2'd0 };
assign lut_1_bit_3_fill = {lut_val_1_n_3_pp[10], lut_val_1_n_3_pp[10], lut_val_1_n_3_pp[10], lut_val_1_n_3_pp[10], lut_val_1_n_3_pp[10], lut_val_1_n_3_pp[10], lut_val_1_n_3_pp[10], lut_val_1_n_3_pp[10],  lut_val_1_n_3_pp, 3'd0 };
assign lut_1_bit_4_fill = {lut_val_1_n_4_pp[10], lut_val_1_n_4_pp[10], lut_val_1_n_4_pp[10], lut_val_1_n_4_pp[10], lut_val_1_n_4_pp[10], lut_val_1_n_4_pp[10], lut_val_1_n_4_pp[10],  lut_val_1_n_4_pp, 4'd0 };
assign lut_1_bit_5_fill = {lut_val_1_n_5_pp[10], lut_val_1_n_5_pp[10], lut_val_1_n_5_pp[10], lut_val_1_n_5_pp[10], lut_val_1_n_5_pp[10], lut_val_1_n_5_pp[10],  lut_val_1_n_5_pp, 5'd0 };
assign lut_1_bit_6_fill = {lut_val_1_n_6_pp[10], lut_val_1_n_6_pp[10], lut_val_1_n_6_pp[10], lut_val_1_n_6_pp[10], lut_val_1_n_6_pp[10],  lut_val_1_n_6_pp, 6'd0 };
assign lut_1_bit_7_fill = {lut_val_1_n_7_pp[10], lut_val_1_n_7_pp[10], lut_val_1_n_7_pp[10], lut_val_1_n_7_pp[10],  lut_val_1_n_7_pp, 7'd0 };
assign lut_1_bit_8_fill = {lut_val_1_n_8_pp[10], lut_val_1_n_8_pp[10], lut_val_1_n_8_pp[10],  lut_val_1_n_8_pp, 8'd0 };
assign lut_1_bit_9_fill = {lut_val_1_n_9_pp[10], lut_val_1_n_9_pp[10],  lut_val_1_n_9_pp, 9'd0 };
assign lut_1_bit_10_fill = {lut_val_1_n_10_pp[10],  lut_val_1_n_10_pp, 10'd0 };
assign lut_1_bit_11_fill = { lut_val_1_n_11_pp, 11'd0 };
wire [22:0] tree_1_pp_l_0_n_0_n;
sadd_lpm_cen Uadd_1_lut_l_0_n_0_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_1_bit_0_fill), .bin(lut_1_bit_1_fill), .res(tree_1_pp_l_0_n_0_n) );
defparam Uadd_1_lut_l_0_n_0_n.IN_WIDTH = 22;
defparam Uadd_1_lut_l_0_n_0_n.PIPE_DEPTH = 3;
wire [22:0] tree_1_pp_l_0_n_1_n;
sadd_lpm_cen Uadd_1_lut_l_0_n_1_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_1_bit_2_fill), .bin(lut_1_bit_3_fill), .res(tree_1_pp_l_0_n_1_n) );
defparam Uadd_1_lut_l_0_n_1_n.IN_WIDTH = 22;
defparam Uadd_1_lut_l_0_n_1_n.PIPE_DEPTH = 3;
wire [22:0] tree_1_pp_l_0_n_2_n;
sadd_lpm_cen Uadd_1_lut_l_0_n_2_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_1_bit_4_fill), .bin(lut_1_bit_5_fill), .res(tree_1_pp_l_0_n_2_n) );
defparam Uadd_1_lut_l_0_n_2_n.IN_WIDTH = 22;
defparam Uadd_1_lut_l_0_n_2_n.PIPE_DEPTH = 3;
wire [22:0] tree_1_pp_l_0_n_3_n;
sadd_lpm_cen Uadd_1_lut_l_0_n_3_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_1_bit_6_fill), .bin(lut_1_bit_7_fill), .res(tree_1_pp_l_0_n_3_n) );
defparam Uadd_1_lut_l_0_n_3_n.IN_WIDTH = 22;
defparam Uadd_1_lut_l_0_n_3_n.PIPE_DEPTH = 3;
wire [22:0] tree_1_pp_l_0_n_4_n;
sadd_lpm_cen Uadd_1_lut_l_0_n_4_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_1_bit_8_fill), .bin(lut_1_bit_9_fill), .res(tree_1_pp_l_0_n_4_n) );
defparam Uadd_1_lut_l_0_n_4_n.IN_WIDTH = 22;
defparam Uadd_1_lut_l_0_n_4_n.PIPE_DEPTH = 3;
wire [22:0] tree_1_pp_l_0_n_5_n;
sadd_lpm_cen Uadd_1_lut_l_0_n_5_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_1_bit_10_fill), .bin(lut_1_bit_11_fill), .res(tree_1_pp_l_0_n_5_n) );
defparam Uadd_1_lut_l_0_n_5_n.IN_WIDTH = 22;
defparam Uadd_1_lut_l_0_n_5_n.PIPE_DEPTH = 3;
wire [23:0] tree_1_pp_l_1_n_0_n;
sadd_lpm_cen Uadd_1_lut_l_1_n_0_n (.clk(clk),  .gclk_en(clk_en), .ain(tree_1_pp_l_0_n_0_n), .bin(tree_1_pp_l_0_n_1_n), .res(tree_1_pp_l_1_n_0_n) );
defparam Uadd_1_lut_l_1_n_0_n.IN_WIDTH = 23;
defparam Uadd_1_lut_l_1_n_0_n.PIPE_DEPTH = 3;
wire [23:0] tree_1_pp_l_1_n_1_n;
sadd_lpm_cen Uadd_1_lut_l_1_n_1_n (.clk(clk),  .gclk_en(clk_en), .ain(tree_1_pp_l_0_n_2_n), .bin(tree_1_pp_l_0_n_3_n), .res(tree_1_pp_l_1_n_1_n) );
defparam Uadd_1_lut_l_1_n_1_n.IN_WIDTH = 23;
defparam Uadd_1_lut_l_1_n_1_n.PIPE_DEPTH = 3;
wire [23:0] tree_1_pp_l_1_n_2_n;
sadd_lpm_cen Uadd_1_lut_l_1_n_2_n (.clk(clk),  .gclk_en(clk_en), .ain(tree_1_pp_l_0_n_4_n), .bin(tree_1_pp_l_0_n_5_n), .res(tree_1_pp_l_1_n_2_n) );
defparam Uadd_1_lut_l_1_n_2_n.IN_WIDTH = 23;
defparam Uadd_1_lut_l_1_n_2_n.PIPE_DEPTH = 3;
wire [24:0] tree_1_pp_l_2_n_0_n;
sadd_lpm_cen Uadd_1_lut_l_2_n_0_n (.clk(clk),  .gclk_en(clk_en), .ain(tree_1_pp_l_1_n_0_n), .bin(tree_1_pp_l_1_n_1_n), .res(tree_1_pp_l_2_n_0_n) );
defparam Uadd_1_lut_l_2_n_0_n.IN_WIDTH = 24;
defparam Uadd_1_lut_l_2_n_0_n.PIPE_DEPTH = 3;
wire [24:0] tree_1_pp_l_2_n_1_n;
sadd_lpm_cen Uadd_1_lut_l_2_n_1_n (.clk(clk),  .gclk_en(clk_en), .ain(tree_1_pp_l_1_n_2_n), .bin(24'd0), .res(tree_1_pp_l_2_n_1_n) );
defparam Uadd_1_lut_l_2_n_1_n.IN_WIDTH = 24;
defparam Uadd_1_lut_l_2_n_1_n.PIPE_DEPTH = 3;
wire [25:0] tree_1_pp_l_3_n_0_n;
sadd_lpm_cen Uadd_1_lut_l_3_n_0_n (.clk(clk),  .gclk_en(clk_en), .ain(tree_1_pp_l_2_n_0_n), .bin(tree_1_pp_l_2_n_1_n), .res(tree_1_pp_l_3_n_0_n) );
defparam Uadd_1_lut_l_3_n_0_n.IN_WIDTH = 25;
defparam Uadd_1_lut_l_3_n_0_n.PIPE_DEPTH = 3;
wire [25:0] lut_val_1_n;
assign lut_val_1_n=tree_1_pp_l_3_n_0_n;
wire [21:0] lut_2_bit_0_fill;
wire [21:0] lut_2_bit_1_fill;
wire [21:0] lut_2_bit_2_fill;
wire [21:0] lut_2_bit_3_fill;
wire [21:0] lut_2_bit_4_fill;
wire [21:0] lut_2_bit_5_fill;
wire [21:0] lut_2_bit_6_fill;
wire [21:0] lut_2_bit_7_fill;
wire [21:0] lut_2_bit_8_fill;
wire [21:0] lut_2_bit_9_fill;
wire [21:0] lut_2_bit_10_fill;
wire [21:0] lut_2_bit_11_fill;
assign lut_2_bit_0_fill = {lut_val_2_n_0_pp[10], lut_val_2_n_0_pp[10], lut_val_2_n_0_pp[10], lut_val_2_n_0_pp[10], lut_val_2_n_0_pp[10], lut_val_2_n_0_pp[10], lut_val_2_n_0_pp[10], lut_val_2_n_0_pp[10], lut_val_2_n_0_pp[10], lut_val_2_n_0_pp[10], lut_val_2_n_0_pp[10],  lut_val_2_n_0_pp };
assign lut_2_bit_1_fill = {lut_val_2_n_1_pp[10], lut_val_2_n_1_pp[10], lut_val_2_n_1_pp[10], lut_val_2_n_1_pp[10], lut_val_2_n_1_pp[10], lut_val_2_n_1_pp[10], lut_val_2_n_1_pp[10], lut_val_2_n_1_pp[10], lut_val_2_n_1_pp[10], lut_val_2_n_1_pp[10],  lut_val_2_n_1_pp, 1'd0 };
assign lut_2_bit_2_fill = {lut_val_2_n_2_pp[10], lut_val_2_n_2_pp[10], lut_val_2_n_2_pp[10], lut_val_2_n_2_pp[10], lut_val_2_n_2_pp[10], lut_val_2_n_2_pp[10], lut_val_2_n_2_pp[10], lut_val_2_n_2_pp[10], lut_val_2_n_2_pp[10],  lut_val_2_n_2_pp, 2'd0 };
assign lut_2_bit_3_fill = {lut_val_2_n_3_pp[10], lut_val_2_n_3_pp[10], lut_val_2_n_3_pp[10], lut_val_2_n_3_pp[10], lut_val_2_n_3_pp[10], lut_val_2_n_3_pp[10], lut_val_2_n_3_pp[10], lut_val_2_n_3_pp[10],  lut_val_2_n_3_pp, 3'd0 };
assign lut_2_bit_4_fill = {lut_val_2_n_4_pp[10], lut_val_2_n_4_pp[10], lut_val_2_n_4_pp[10], lut_val_2_n_4_pp[10], lut_val_2_n_4_pp[10], lut_val_2_n_4_pp[10], lut_val_2_n_4_pp[10],  lut_val_2_n_4_pp, 4'd0 };
assign lut_2_bit_5_fill = {lut_val_2_n_5_pp[10], lut_val_2_n_5_pp[10], lut_val_2_n_5_pp[10], lut_val_2_n_5_pp[10], lut_val_2_n_5_pp[10], lut_val_2_n_5_pp[10],  lut_val_2_n_5_pp, 5'd0 };
assign lut_2_bit_6_fill = {lut_val_2_n_6_pp[10], lut_val_2_n_6_pp[10], lut_val_2_n_6_pp[10], lut_val_2_n_6_pp[10], lut_val_2_n_6_pp[10],  lut_val_2_n_6_pp, 6'd0 };
assign lut_2_bit_7_fill = {lut_val_2_n_7_pp[10], lut_val_2_n_7_pp[10], lut_val_2_n_7_pp[10], lut_val_2_n_7_pp[10],  lut_val_2_n_7_pp, 7'd0 };
assign lut_2_bit_8_fill = {lut_val_2_n_8_pp[10], lut_val_2_n_8_pp[10], lut_val_2_n_8_pp[10],  lut_val_2_n_8_pp, 8'd0 };
assign lut_2_bit_9_fill = {lut_val_2_n_9_pp[10], lut_val_2_n_9_pp[10],  lut_val_2_n_9_pp, 9'd0 };
assign lut_2_bit_10_fill = {lut_val_2_n_10_pp[10],  lut_val_2_n_10_pp, 10'd0 };
assign lut_2_bit_11_fill = { lut_val_2_n_11_pp, 11'd0 };
wire [22:0] tree_2_pp_l_0_n_0_n;
sadd_lpm_cen Uadd_2_lut_l_0_n_0_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_2_bit_0_fill), .bin(lut_2_bit_1_fill), .res(tree_2_pp_l_0_n_0_n) );
defparam Uadd_2_lut_l_0_n_0_n.IN_WIDTH = 22;
defparam Uadd_2_lut_l_0_n_0_n.PIPE_DEPTH = 3;
wire [22:0] tree_2_pp_l_0_n_1_n;
sadd_lpm_cen Uadd_2_lut_l_0_n_1_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_2_bit_2_fill), .bin(lut_2_bit_3_fill), .res(tree_2_pp_l_0_n_1_n) );
defparam Uadd_2_lut_l_0_n_1_n.IN_WIDTH = 22;
defparam Uadd_2_lut_l_0_n_1_n.PIPE_DEPTH = 3;
wire [22:0] tree_2_pp_l_0_n_2_n;
sadd_lpm_cen Uadd_2_lut_l_0_n_2_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_2_bit_4_fill), .bin(lut_2_bit_5_fill), .res(tree_2_pp_l_0_n_2_n) );
defparam Uadd_2_lut_l_0_n_2_n.IN_WIDTH = 22;
defparam Uadd_2_lut_l_0_n_2_n.PIPE_DEPTH = 3;
wire [22:0] tree_2_pp_l_0_n_3_n;
sadd_lpm_cen Uadd_2_lut_l_0_n_3_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_2_bit_6_fill), .bin(lut_2_bit_7_fill), .res(tree_2_pp_l_0_n_3_n) );
defparam Uadd_2_lut_l_0_n_3_n.IN_WIDTH = 22;
defparam Uadd_2_lut_l_0_n_3_n.PIPE_DEPTH = 3;
wire [22:0] tree_2_pp_l_0_n_4_n;
sadd_lpm_cen Uadd_2_lut_l_0_n_4_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_2_bit_8_fill), .bin(lut_2_bit_9_fill), .res(tree_2_pp_l_0_n_4_n) );
defparam Uadd_2_lut_l_0_n_4_n.IN_WIDTH = 22;
defparam Uadd_2_lut_l_0_n_4_n.PIPE_DEPTH = 3;
wire [22:0] tree_2_pp_l_0_n_5_n;
sadd_lpm_cen Uadd_2_lut_l_0_n_5_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_2_bit_10_fill), .bin(lut_2_bit_11_fill), .res(tree_2_pp_l_0_n_5_n) );
defparam Uadd_2_lut_l_0_n_5_n.IN_WIDTH = 22;
defparam Uadd_2_lut_l_0_n_5_n.PIPE_DEPTH = 3;
wire [23:0] tree_2_pp_l_1_n_0_n;
sadd_lpm_cen Uadd_2_lut_l_1_n_0_n (.clk(clk),  .gclk_en(clk_en), .ain(tree_2_pp_l_0_n_0_n), .bin(tree_2_pp_l_0_n_1_n), .res(tree_2_pp_l_1_n_0_n) );
defparam Uadd_2_lut_l_1_n_0_n.IN_WIDTH = 23;
defparam Uadd_2_lut_l_1_n_0_n.PIPE_DEPTH = 3;
wire [23:0] tree_2_pp_l_1_n_1_n;
sadd_lpm_cen Uadd_2_lut_l_1_n_1_n (.clk(clk),  .gclk_en(clk_en), .ain(tree_2_pp_l_0_n_2_n), .bin(tree_2_pp_l_0_n_3_n), .res(tree_2_pp_l_1_n_1_n) );
defparam Uadd_2_lut_l_1_n_1_n.IN_WIDTH = 23;
defparam Uadd_2_lut_l_1_n_1_n.PIPE_DEPTH = 3;
wire [23:0] tree_2_pp_l_1_n_2_n;
sadd_lpm_cen Uadd_2_lut_l_1_n_2_n (.clk(clk),  .gclk_en(clk_en), .ain(tree_2_pp_l_0_n_4_n), .bin(tree_2_pp_l_0_n_5_n), .res(tree_2_pp_l_1_n_2_n) );
defparam Uadd_2_lut_l_1_n_2_n.IN_WIDTH = 23;
defparam Uadd_2_lut_l_1_n_2_n.PIPE_DEPTH = 3;
wire [24:0] tree_2_pp_l_2_n_0_n;
sadd_lpm_cen Uadd_2_lut_l_2_n_0_n (.clk(clk),  .gclk_en(clk_en), .ain(tree_2_pp_l_1_n_0_n), .bin(tree_2_pp_l_1_n_1_n), .res(tree_2_pp_l_2_n_0_n) );
defparam Uadd_2_lut_l_2_n_0_n.IN_WIDTH = 24;
defparam Uadd_2_lut_l_2_n_0_n.PIPE_DEPTH = 3;
wire [24:0] tree_2_pp_l_2_n_1_n;
sadd_lpm_cen Uadd_2_lut_l_2_n_1_n (.clk(clk),  .gclk_en(clk_en), .ain(tree_2_pp_l_1_n_2_n), .bin(24'd0), .res(tree_2_pp_l_2_n_1_n) );
defparam Uadd_2_lut_l_2_n_1_n.IN_WIDTH = 24;
defparam Uadd_2_lut_l_2_n_1_n.PIPE_DEPTH = 3;
wire [25:0] tree_2_pp_l_3_n_0_n;
sadd_lpm_cen Uadd_2_lut_l_3_n_0_n (.clk(clk),  .gclk_en(clk_en), .ain(tree_2_pp_l_2_n_0_n), .bin(tree_2_pp_l_2_n_1_n), .res(tree_2_pp_l_3_n_0_n) );
defparam Uadd_2_lut_l_3_n_0_n.IN_WIDTH = 25;
defparam Uadd_2_lut_l_3_n_0_n.PIPE_DEPTH = 3;
wire [25:0] lut_val_2_n;
assign lut_val_2_n=tree_2_pp_l_3_n_0_n;
wire [21:0] lut_3_bit_0_fill;
wire [21:0] lut_3_bit_1_fill;
wire [21:0] lut_3_bit_2_fill;
wire [21:0] lut_3_bit_3_fill;
wire [21:0] lut_3_bit_4_fill;
wire [21:0] lut_3_bit_5_fill;
wire [21:0] lut_3_bit_6_fill;
wire [21:0] lut_3_bit_7_fill;
wire [21:0] lut_3_bit_8_fill;
wire [21:0] lut_3_bit_9_fill;
wire [21:0] lut_3_bit_10_fill;
wire [21:0] lut_3_bit_11_fill;
assign lut_3_bit_0_fill = {lut_val_3_n_0_pp[10], lut_val_3_n_0_pp[10], lut_val_3_n_0_pp[10], lut_val_3_n_0_pp[10], lut_val_3_n_0_pp[10], lut_val_3_n_0_pp[10], lut_val_3_n_0_pp[10], lut_val_3_n_0_pp[10], lut_val_3_n_0_pp[10], lut_val_3_n_0_pp[10], lut_val_3_n_0_pp[10],  lut_val_3_n_0_pp };
assign lut_3_bit_1_fill = {lut_val_3_n_1_pp[10], lut_val_3_n_1_pp[10], lut_val_3_n_1_pp[10], lut_val_3_n_1_pp[10], lut_val_3_n_1_pp[10], lut_val_3_n_1_pp[10], lut_val_3_n_1_pp[10], lut_val_3_n_1_pp[10], lut_val_3_n_1_pp[10], lut_val_3_n_1_pp[10],  lut_val_3_n_1_pp, 1'd0 };
assign lut_3_bit_2_fill = {lut_val_3_n_2_pp[10], lut_val_3_n_2_pp[10], lut_val_3_n_2_pp[10], lut_val_3_n_2_pp[10], lut_val_3_n_2_pp[10], lut_val_3_n_2_pp[10], lut_val_3_n_2_pp[10], lut_val_3_n_2_pp[10], lut_val_3_n_2_pp[10],  lut_val_3_n_2_pp, 2'd0 };
assign lut_3_bit_3_fill = {lut_val_3_n_3_pp[10], lut_val_3_n_3_pp[10], lut_val_3_n_3_pp[10], lut_val_3_n_3_pp[10], lut_val_3_n_3_pp[10], lut_val_3_n_3_pp[10], lut_val_3_n_3_pp[10], lut_val_3_n_3_pp[10],  lut_val_3_n_3_pp, 3'd0 };
assign lut_3_bit_4_fill = {lut_val_3_n_4_pp[10], lut_val_3_n_4_pp[10], lut_val_3_n_4_pp[10], lut_val_3_n_4_pp[10], lut_val_3_n_4_pp[10], lut_val_3_n_4_pp[10], lut_val_3_n_4_pp[10],  lut_val_3_n_4_pp, 4'd0 };
assign lut_3_bit_5_fill = {lut_val_3_n_5_pp[10], lut_val_3_n_5_pp[10], lut_val_3_n_5_pp[10], lut_val_3_n_5_pp[10], lut_val_3_n_5_pp[10], lut_val_3_n_5_pp[10],  lut_val_3_n_5_pp, 5'd0 };
assign lut_3_bit_6_fill = {lut_val_3_n_6_pp[10], lut_val_3_n_6_pp[10], lut_val_3_n_6_pp[10], lut_val_3_n_6_pp[10], lut_val_3_n_6_pp[10],  lut_val_3_n_6_pp, 6'd0 };
assign lut_3_bit_7_fill = {lut_val_3_n_7_pp[10], lut_val_3_n_7_pp[10], lut_val_3_n_7_pp[10], lut_val_3_n_7_pp[10],  lut_val_3_n_7_pp, 7'd0 };
assign lut_3_bit_8_fill = {lut_val_3_n_8_pp[10], lut_val_3_n_8_pp[10], lut_val_3_n_8_pp[10],  lut_val_3_n_8_pp, 8'd0 };
assign lut_3_bit_9_fill = {lut_val_3_n_9_pp[10], lut_val_3_n_9_pp[10],  lut_val_3_n_9_pp, 9'd0 };
assign lut_3_bit_10_fill = {lut_val_3_n_10_pp[10],  lut_val_3_n_10_pp, 10'd0 };
assign lut_3_bit_11_fill = { lut_val_3_n_11_pp, 11'd0 };
wire [22:0] tree_3_pp_l_0_n_0_n;
sadd_lpm_cen Uadd_3_lut_l_0_n_0_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_3_bit_0_fill), .bin(lut_3_bit_1_fill), .res(tree_3_pp_l_0_n_0_n) );
defparam Uadd_3_lut_l_0_n_0_n.IN_WIDTH = 22;
defparam Uadd_3_lut_l_0_n_0_n.PIPE_DEPTH = 3;
wire [22:0] tree_3_pp_l_0_n_1_n;
sadd_lpm_cen Uadd_3_lut_l_0_n_1_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_3_bit_2_fill), .bin(lut_3_bit_3_fill), .res(tree_3_pp_l_0_n_1_n) );
defparam Uadd_3_lut_l_0_n_1_n.IN_WIDTH = 22;
defparam Uadd_3_lut_l_0_n_1_n.PIPE_DEPTH = 3;
wire [22:0] tree_3_pp_l_0_n_2_n;
sadd_lpm_cen Uadd_3_lut_l_0_n_2_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_3_bit_4_fill), .bin(lut_3_bit_5_fill), .res(tree_3_pp_l_0_n_2_n) );
defparam Uadd_3_lut_l_0_n_2_n.IN_WIDTH = 22;
defparam Uadd_3_lut_l_0_n_2_n.PIPE_DEPTH = 3;
wire [22:0] tree_3_pp_l_0_n_3_n;
sadd_lpm_cen Uadd_3_lut_l_0_n_3_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_3_bit_6_fill), .bin(lut_3_bit_7_fill), .res(tree_3_pp_l_0_n_3_n) );
defparam Uadd_3_lut_l_0_n_3_n.IN_WIDTH = 22;
defparam Uadd_3_lut_l_0_n_3_n.PIPE_DEPTH = 3;
wire [22:0] tree_3_pp_l_0_n_4_n;
sadd_lpm_cen Uadd_3_lut_l_0_n_4_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_3_bit_8_fill), .bin(lut_3_bit_9_fill), .res(tree_3_pp_l_0_n_4_n) );
defparam Uadd_3_lut_l_0_n_4_n.IN_WIDTH = 22;
defparam Uadd_3_lut_l_0_n_4_n.PIPE_DEPTH = 3;
wire [22:0] tree_3_pp_l_0_n_5_n;
sadd_lpm_cen Uadd_3_lut_l_0_n_5_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_3_bit_10_fill), .bin(lut_3_bit_11_fill), .res(tree_3_pp_l_0_n_5_n) );
defparam Uadd_3_lut_l_0_n_5_n.IN_WIDTH = 22;
defparam Uadd_3_lut_l_0_n_5_n.PIPE_DEPTH = 3;
wire [23:0] tree_3_pp_l_1_n_0_n;
sadd_lpm_cen Uadd_3_lut_l_1_n_0_n (.clk(clk),  .gclk_en(clk_en), .ain(tree_3_pp_l_0_n_0_n), .bin(tree_3_pp_l_0_n_1_n), .res(tree_3_pp_l_1_n_0_n) );
defparam Uadd_3_lut_l_1_n_0_n.IN_WIDTH = 23;
defparam Uadd_3_lut_l_1_n_0_n.PIPE_DEPTH = 3;
wire [23:0] tree_3_pp_l_1_n_1_n;
sadd_lpm_cen Uadd_3_lut_l_1_n_1_n (.clk(clk),  .gclk_en(clk_en), .ain(tree_3_pp_l_0_n_2_n), .bin(tree_3_pp_l_0_n_3_n), .res(tree_3_pp_l_1_n_1_n) );
defparam Uadd_3_lut_l_1_n_1_n.IN_WIDTH = 23;
defparam Uadd_3_lut_l_1_n_1_n.PIPE_DEPTH = 3;
wire [23:0] tree_3_pp_l_1_n_2_n;
sadd_lpm_cen Uadd_3_lut_l_1_n_2_n (.clk(clk),  .gclk_en(clk_en), .ain(tree_3_pp_l_0_n_4_n), .bin(tree_3_pp_l_0_n_5_n), .res(tree_3_pp_l_1_n_2_n) );
defparam Uadd_3_lut_l_1_n_2_n.IN_WIDTH = 23;
defparam Uadd_3_lut_l_1_n_2_n.PIPE_DEPTH = 3;
wire [24:0] tree_3_pp_l_2_n_0_n;
sadd_lpm_cen Uadd_3_lut_l_2_n_0_n (.clk(clk),  .gclk_en(clk_en), .ain(tree_3_pp_l_1_n_0_n), .bin(tree_3_pp_l_1_n_1_n), .res(tree_3_pp_l_2_n_0_n) );
defparam Uadd_3_lut_l_2_n_0_n.IN_WIDTH = 24;
defparam Uadd_3_lut_l_2_n_0_n.PIPE_DEPTH = 3;
wire [24:0] tree_3_pp_l_2_n_1_n;
sadd_lpm_cen Uadd_3_lut_l_2_n_1_n (.clk(clk),  .gclk_en(clk_en), .ain(tree_3_pp_l_1_n_2_n), .bin(24'd0), .res(tree_3_pp_l_2_n_1_n) );
defparam Uadd_3_lut_l_2_n_1_n.IN_WIDTH = 24;
defparam Uadd_3_lut_l_2_n_1_n.PIPE_DEPTH = 3;
wire [25:0] tree_3_pp_l_3_n_0_n;
sadd_lpm_cen Uadd_3_lut_l_3_n_0_n (.clk(clk),  .gclk_en(clk_en), .ain(tree_3_pp_l_2_n_0_n), .bin(tree_3_pp_l_2_n_1_n), .res(tree_3_pp_l_3_n_0_n) );
defparam Uadd_3_lut_l_3_n_0_n.IN_WIDTH = 25;
defparam Uadd_3_lut_l_3_n_0_n.PIPE_DEPTH = 3;
wire [25:0] lut_val_3_n;
assign lut_val_3_n=tree_3_pp_l_3_n_0_n;
wire [26:0] fin_atree_l_0_n_0_n;
sadd_lpm_cen Uadd_cen_l_0_n_0_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_val_0_n), .bin(lut_val_1_n), .res(fin_atree_l_0_n_0_n) );
defparam Uadd_cen_l_0_n_0_n.IN_WIDTH = 26;
defparam Uadd_cen_l_0_n_0_n.PIPE_DEPTH = 3;
wire [26:0] fin_atree_l_0_n_1_n;
sadd_lpm_cen Uadd_cen_l_0_n_1_n (.clk(clk),  .gclk_en(clk_en), .ain(lut_val_2_n), .bin(lut_val_3_n), .res(fin_atree_l_0_n_1_n) );
defparam Uadd_cen_l_0_n_1_n.IN_WIDTH = 26;
defparam Uadd_cen_l_0_n_1_n.PIPE_DEPTH = 3;
wire [27:0] fin_atree_l_1_n_0_n;
sadd_lpm_cen Uadd_cen_l_1_n_0_n (.clk(clk),  .gclk_en(clk_en), .ain(fin_atree_l_0_n_0_n), .bin(fin_atree_l_0_n_1_n), .res(fin_atree_l_1_n_0_n) );
defparam Uadd_cen_l_1_n_0_n.IN_WIDTH = 27;
defparam Uadd_cen_l_1_n_0_n.PIPE_DEPTH = 3;
wire [27:0] mac_res;
assign mac_res=fin_atree_l_1_n_0_n;
wire [27:0] atree_res;
mac_tl Umtl (.clk(clk),
             .data_in(mac_res),
             .data_out(atree_res));
defparam Umtl.DATA_WIDTH = 28;
wire [23:0] fir_int_res;
assign fir_int_res = atree_res [23:0];
wire [23:0]fir_int_res_fill;
assign fir_int_res_fill =  fir_int_res[23 :0];
parameter TOT_WIDTH = ACCUM_WIDTH;
assign fir_result = fir_int_res_fill[TOT_WIDTH-MSB_RM-1:LSB_RM];
wire pre_rdy;
assign rdy_to_ld = pre_rdy;
assign done = done_int;
par_ctrl Uctrl(.rst(rst),
		.clk(clk),
		.clk_en(clk_en),
		.done(done_int),
		.rdy_int(rdy_int),
		.rdy_to_ld(pre_rdy));
defparam Uctrl.REG_LEN = 21;
defparam Uctrl.REG_BIT = 5;
defparam Uctrl.CH_WIDTH =0;
defparam Uctrl.NUM_CH =1;
endmodule