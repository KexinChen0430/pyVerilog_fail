module TOP(
	output N2_CAn_O,
	output N2_CBn_O,
	output N2_CCn_O,
	output N2_CDn_O,
	output N2_CEn_O,
	output N2_CFn_O,
	output N2_CGn_O,
	output N2_CDPn_O,
	output N2_AN0n_O,
	output N2_AN1n_O,
	output N2_AN2n_O,
	output N2_AN3n_O,
	output N2_HSYNC_O,
	output N2_VSYNC_O,
	output [2:0] N2_RED_O,
	output [2:0] N2_GRN_O,
	output [2:1] N2_BLU_O,
	input N2_PS2DAT_IO,
	input N2_PS2CLK_I,
	input N2_50MHZ_I,
	input N2_RST_I
);
	wire	[15:1]	cpu_adr;
	wire				cpu_we;
	wire				cpu_cyc;
	wire				cpu_stb;
	wire	[1:0]		cpu_sel;
	wire				cpu_vda;
	wire				cpu_vpa;
	wire	[15:0]	cpu_dat_o;
	wire	[7:0]		kia_dat_o;
	wire				kia_ack_o;
	wire	[15:0]	ram_dat_o;
	reg				ram_ack_o;
	reg				led_a;
	reg				led_b;
	reg				led_c;
	reg				led_d;
	reg				led_e;
	reg				led_f;
	reg				led_g;
	reg				led_dp;
	reg				led_anode_0;
	reg				led_anode_1;
	reg				led_anode_2;
	reg				led_anode_3;
	reg				vsync;
	reg				hsync;
	reg	[2:0]		red;
	reg	[2:0]		green;
	reg	[2:1]		blue;
	wire	bus_access				= cpu_cyc & cpu_stb;
	wire	kia_addressed 			= (cpu_adr[15:12] == 4'h2) & bus_access & cpu_sel[0];
	wire	ledport_addressed		= (cpu_adr[15:12] == 4'h1) & bus_access;
	wire	ram_addressed 			= (cpu_adr[15:12] == 4'h0) & bus_access;
	wire	[15:0]	cpu_dat_i 	= ({16{ram_addressed}} & ram_dat_o) | {8'h00, ({8{kia_addressed}} & kia_dat_o)};
	wire	cpu_ack_i				= ((ram_addressed | ledport_addressed ) & ram_ack_o) | (kia_addressed & kia_ack_o);
	STEAMER16X4 cpu(
		.clk_i(N2_50MHZ_I),
		.res_i(N2_RST_I),
		.adr_o(cpu_adr),
		.we_o (cpu_we),
		.cyc_o(cpu_cyc),
		.stb_o(cpu_stb),
		.sel_o(cpu_sel),
		.vda_o(cpu_vda),
		.vpa_o(cpu_vpa),
		.dat_o(cpu_dat_o),
		.ack_i(cpu_ack_i),
		.dat_i(cpu_dat_i)
	);
	wire	ram_even_en = ram_addressed & cpu_sel[0];
	wire	ram_odd_en  = ram_addressed & cpu_sel[1];
	RAMB16_S9 progmem_E(
		.CLK(N2_50MHZ_I),
		.WE(cpu_we),
		.EN(ram_even_en),
		.SSR(1'b0),
		.ADDR(cpu_adr[11:1]),
		.DI(cpu_dat_o[7:0]),
		.DO(ram_dat_o[7:0]),
		.DIP(1'b1)
	);
	RAMB16_S9 progmem_O(
		.CLK(N2_50MHZ_I),
		.WE(cpu_we),
		.EN(ram_odd_en),
		.SSR(1'b0),
		.ADDR(cpu_adr[11:1]),
		.DI(cpu_dat_o[15:8]),
		.DO(ram_dat_o[15:8]),
		.DIP(1'b1)
	);
	always @(posedge N2_50MHZ_I) begin
		if(N2_RST_I) begin
			ram_ack_o <= 0;
		end else begin
			ram_ack_o <= (~ram_ack_o) & (ram_addressed | ledport_addressed);
		end
	end
	KIA_M kia(
		.CLK_I(N2_50MHZ_I),
		.RES_I(N2_RST_I),
		.ADR_I(cpu_adr[1]),
		.WE_I(cpu_we),
		.CYC_I(cpu_cyc),
		.STB_I(kia_addressed),
		.ACK_O(kia_ack_o),
		.DAT_O(kia_dat_o[7:0]),
		.D_I(N2_PS2DAT_IO),
		.C_I(N2_PS2CLK_I)
	);
   assign N2_CAn_O = ~led_a;
   assign N2_CBn_O = ~led_b;
   assign N2_CCn_O = ~led_c;
   assign N2_CDn_O = ~led_d;
   assign N2_CEn_O = ~led_e;
   assign N2_CFn_O = ~led_f;
   assign N2_CGn_O = ~led_g;
   assign N2_CDPn_O = ~led_dp;
   assign N2_AN0n_O = ~led_anode_0;
   assign N2_AN1n_O = ~led_anode_1;
   assign N2_AN2n_O = ~led_anode_2;
   assign N2_AN3n_O = ~led_anode_3;
	assign N2_VSYNC_O = vsync;
	assign N2_HSYNC_O = hsync;
	assign N2_RED_O = red;
	assign N2_GRN_O = green;
	assign N2_BLU_O = blue;
	always @(posedge N2_50MHZ_I) begin
		if(N2_RST_I) begin
			led_a <= 1;				led_e <= 1;
			led_b <= 1;				led_f <= 1;
			led_c <= 1;				led_g <= 1;
			led_d <= 1;				led_dp <= 1;
			led_anode_0 <= 1;		led_anode_1 <= 1;
			led_anode_2 <= 1;		led_anode_3 <= 1;
			vsync <= 1;				hsync <= 1;
			red <= 3'b000;			green <= 3'b000;
			blue <= 2'b00;
		end
		else begin
			if(ledport_addressed & cpu_sel[0]) begin
				led_a <= cpu_dat_o[0];	led_e <= cpu_dat_o[4];
				led_b <= cpu_dat_o[1];	led_f <= cpu_dat_o[5];
				led_c <= cpu_dat_o[2];	led_g <= cpu_dat_o[6];
				led_d <= cpu_dat_o[3];	led_dp <= cpu_dat_o[7];
			end
			if(ledport_addressed & cpu_sel[1]) begin
				led_anode_0 <= cpu_dat_o[12];
				led_anode_1 <= cpu_dat_o[13];
				led_anode_2 <= cpu_dat_o[14];
				led_anode_3 <= cpu_dat_o[15];
			end
		end
	end
	defparam
progmem_E.INIT_00 = 256'h030202020202020202010101010101010100000000000000000000000000E200,
progmem_E.INIT_01 = 256'h0706060606060606060505050505050505040404040404040403030303030303,
progmem_E.INIT_02 = 256'h0B0A0A0A0A0A0A0A0A0909090909090909080808080808080807070707070707,
progmem_E.INIT_03 = 256'h0F0E0E0E0E0E0E0E0E0D0D0D0D0D0D0D0D0C0C0C0C0C0C0C0C0B0B0B0B0B0B0B,
progmem_E.INIT_04 = 256'h3A00001EE009081B0A091B0B0A1B1E00007939777F7D665B3F0F0F0F0F0F0F0F,
progmem_E.INIT_05 = 256'hE007000F06156E000054E03C6AE007B00E0614540000003A08B10E07142046E0,
progmem_E.INIT_06 = 256'h14B80000009E02128AB0E006021B9E000088E0709AE05694E08800006EE03C84,
progmem_E.INIT_07 = 256'hD600E00000000816EA0000D4E0BAE6E00C0030D40000B8E0BED01E0C0C12FF0C,
progmem_E.INIT_08 = 256'h163800001EE0D634E00000000A161E000004E0D61AE00000000916040000EAE0,
progmem_E.INIT_09 = 256'hE0EC7EE00678E02072E03A6CE06000000052001252000038E0D64EE00000000B,
progmem_E.INIT_0A = 256'h9CE0A20062B8E0A0B2E0B2008AA8E09C00000088011201001588000060E05484,
progmem_E.INIT_0B = 256'hFFFFBEFF00E0E09EF2E0C2ECE0E00000C0E00B001B0A000911000800B1C00000,
progmem_E.INIT_0C = 256'h3BBFDFFCE000BF6EFFFFFF162FFFF81DFFFDC2F8FB5E5DBEF9F7FBF1BBBFE2FF,
progmem_E.INIT_0D = 256'hBCE1FEFF241278FF972AFFFFFFFF6CFE2D2B7EFFFFC22CB216B2BFF8C003030E,
progmem_E.INIT_0E = 256'h5FC5FDFFFFFF7E2BFFCBC5C7FFFFFF5C92FFF2BFFFBFEF7EF0F87FBBBFBB5FC5,
progmem_E.INIT_0F = 256'hFFBFFB5FFD2FFF775F2D00000000200000000020BBFDC5FFE5E2EDE27EDF5FF9,
progmem_E.INIT_10 = 256'h97FFBFDFC5F7FFFFC57F8B26C4FEFFFBFFFFFFAF7FFFFFDDDFF1F7BDDF7FF2C5,
progmem_E.INIT_11 = 256'hE2FE7FE597F97E79F88BF8FFFF24F0F9FFE73FF297FF3F4949F1F1912CBDFDF9,
progmem_E.INIT_12 = 256'hFCFE5FE5FEFF7F5FF9BFFFABCBFFBF8500000000000048F2FFBFFFE2592E9716,
progmem_E.INIT_13 = 256'h5957E2FF97E6F1CCCC8CE5FCFFB6E2CB49FFD7D7FFF9FFFFFFFFF87F97F9FFFE,
progmem_E.INIT_14 = 256'h7CBFFFFFBF972FDB7BDFF97F5FFE2FFFEF6FF9FDF75BDF99F397D7E557FFFEFD,
progmem_E.INIT_15 = 256'hE2F9321244915FFF5FFFF998F9FF77F77FFBFF2FFCDFF1F2FD7B7F25F8E5975F,
progmem_E.INIT_16 = 256'hBFDFFF17FFFFF97F5F92BEFF8BBEFFC55FF2CBFFFFC57FFDFCFF452FFCE225FC,
progmem_E.INIT_17 = 256'hF8F876127D5B16CB49F75E0B4849249292CBF97FFD856619FDBF97FFFF655FCB,
progmem_E.INIT_18 = 256'hFFAFF797FFF2FFFFBFAF7C450402082021410410422110211020418108088484,
progmem_E.INIT_19 = 256'h5F5FFFDE7FBB1624482FF2E7F2FFFFFBBFFFFFFFFFDFFFE5FFFEFF92ED7F725B,
progmem_E.INIT_1A = 256'hFBFBFFF7FFEF7D7DFFFFFF8BFBEFFFF917EDFAFBFFFEED7FFF7D95F8FFFF7F7F,
progmem_E.INIT_1B = 256'hFFBFFEDF5BBFFFFFFB7FEFFFF7FFF67FBFFFE5FB7EF22BE589FFFFAFFF77927F,
progmem_E.INIT_1C = 256'hFFAF5FFF7FC27E080000209249248244BFFFF7FEDFFE7FAFFFFDFFFFFECBFF5F,
progmem_E.INIT_1D = 256'hFFF7CBBE81F81244E6FFFF5FF3FEFF3FE57FCFF95FF857FFFFC27F857EDFFFFB,
progmem_E.INIT_1E = 256'hEFFFFFEFFFFFF7EFFFDFFCF22FF8FFDBFFFFF1FFBFED8BFB5FE52FF2FEFF7FBC,
progmem_E.INIT_1F = 256'h5FBFFFFFFF5FFC2F85FFFFB51FFFFFF1FF62FFF1C28B8AFE7FFE7F6E25F7F7F2;
	defparam
progmem_O.INIT_00 = 256'h030202020202020202010101010101010100000000000000000000000000021E,
progmem_O.INIT_01 = 256'h0706060606060606060505050505050505040404040404040403030303030303,
progmem_O.INIT_02 = 256'h0B0A0A0A0A0A0A0A0A0909090909090909080808080808080807070707070707,
progmem_O.INIT_03 = 256'h0F0E0E0E0E0E0E0E0E0D0D0D0D0D0D0D0D0C0C0C0C0C0C0C0C0B0B0B0B0B0B0B,
progmem_O.INIT_04 = 256'h011300011200001A00001A00001A011300715E7C6F076D4F060F0F0F0F0F0F0F,
progmem_O.INIT_05 = 256'h11001B00001A011300011201011100A100001A0113002E0100A101001A010111,
progmem_O.INIT_06 = 256'h12011300E001201B01011100201A011300011201011101011101130001120101,
progmem_O.INIT_07 = 256'h010211101310001A01130001120101110040110113000112010117000013FF00,
progmem_O.INIT_08 = 256'h1A0213000212010211101340001A0213000212010211101320001A0213000112,
progmem_O.INIT_09 = 256'h11010211020211020211020211021300E0021013021300021201021110138000,
progmem_O.INIT_0A = 256'h0212021E0202110102110217020211021300E002001600201A02130002120202,
progmem_O.INIT_0B = 256'hFFFFFFED00021202021102021102130002120000B10000001B00000011021300,
progmem_O.INIT_0C = 256'hF0C083010E772FF8E1FF052FDF7FAFE58BFFFFBFFDFFF1FC7F17FF7DFEFDFCFB,
progmem_O.INIT_0D = 256'h5F63577F5E498959FFEFFEFFFFFF2FF9FF9757EF2FC5B2CB2CCB2C031DBFBFFC,
progmem_O.INIT_0E = 256'hCB7CEFFDF8E25F7F92FFEF7FFFDF975F49E4FFFF7FC5F300073B9DF7FFF38BFC,
progmem_O.INIT_0F = 256'hDFFFF777FCBBFFE2FFDE01000000000100000000FFF7BE2FFFFFFFDF2FF9FB7E,
progmem_O.INIT_10 = 256'hE5FFCBDCFBFF0BFFEFFFE12F0C2FBF7FBFFF8BFFF8F1C5F7BF7F7DC58B77EF7F,
progmem_O.INIT_11 = 256'hFF5FE579957F5DF959FFBFFFF2BF7E7FE1E22FFEF39F2F7F24227B7D48FAF87F,
progmem_O.INIT_12 = 256'h5D5FE5FE5FE5F2F97EFFFCFFFFFFF8FC25000000000082FC2ECBC5CB7FFCF35F,
progmem_O.INIT_13 = 256'h2596FE97FF2F7FCBCCCCF9AF155FF8FF652EEBE5AF77FFF22FF2B297F97F97FF,
progmem_O.INIT_14 = 256'hBE99FCF7FD8A97F7BFBF77EFF7FEFEFFEFFE25FF7DBE127F2FFFCB752B2E5FFF,
progmem_O.INIT_15 = 256'hF27FFF238922C8FC95FCCBBF7FFFF7FCFFBFEFC5BFF27DEFFFCBFFF9B1F2CB2F,
progmem_O.INIT_16 = 256'hF7FFE2BFBDFF7BFFE1E9A578FFC4FFBFDFFEFFFFFFF7E7F1BF7BFEF2BEFB8B91,
progmem_O.INIT_17 = 256'h88BF5F1689B1EC3B6E24E2DC9324924944E07EC1D98B2E8C7FCB7FDFF7FFE6DE,
progmem_O.INIT_18 = 256'hFEC5FCE5FF4BD7DFFFCC24FF2208128208041082100884084282080880442120,
progmem_O.INIT_19 = 256'hF1FCF9FFFBE52C89919249C5FFFFFFDFFFFED6FF2FFFFAFFD717EF57FDFFB9E5,
progmem_O.INIT_1A = 256'hF997FF7FBECAFFF1F1FFFFEFFFFF176FFFFFEFFFFF2FFFFAF9EFFFBFDEFBEDF9,
progmem_O.INIT_1B = 256'hFECB2496F29217BF7FDFCBDDF2DFFFCBF7FFFEFD5FFF77FF17FFFF729CE249BF,
progmem_O.INIT_1C = 256'h0BF7F8FCC5BF2FB1000000492492242495C2FFFFDF2EFFFFF8FF7FDF2BCBFFDF,
progmem_O.INIT_1D = 256'hEFFF2FA2F8572F89623FE5F3FE5F3FE5FFCFF97FF3B8C5BCE2BBFF7FFF85018B,
progmem_O.INIT_1E = 256'hFDFFEFFFFFEFFFFFBDEFB7FEFFAFFFFFC58B7FFFFFE2BEFDEBFCFFEC5D7ADEBF,
progmem_O.INIT_1F = 256'hFFBCFCFFFFFFBC0BFE17FFBFF8FE9F5FFFF7FF7FFFFFFF5F9549CBF9B9997FE5;
endmodule