module cpu_rom (Address, OutClock, OutClockEn, Reset, Q)/* synthesis NGD_DRC_MASK=1 */;
    input wire [7:0] Address;
    input wire OutClock;
    input wire OutClockEn;
    input wire Reset;
    output wire [15:0] Q;
    wire scuba_vhi;
    wire scuba_vlo;
    VHI scuba_vhi_inst (.Z(scuba_vhi));
    VLO scuba_vlo_inst (.Z(scuba_vlo));
    defparam cpu_rom_0_0_0.INIT_DATA = "STATIC" ;
    defparam cpu_rom_0_0_0.ASYNC_RESET_RELEASE = "SYNC" ;
    defparam cpu_rom_0_0_0.INITVAL_1F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam cpu_rom_0_0_0.INITVAL_1E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam cpu_rom_0_0_0.INITVAL_1D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam cpu_rom_0_0_0.INITVAL_1C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam cpu_rom_0_0_0.INITVAL_1B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam cpu_rom_0_0_0.INITVAL_1A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam cpu_rom_0_0_0.INITVAL_19 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam cpu_rom_0_0_0.INITVAL_18 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam cpu_rom_0_0_0.INITVAL_17 = "0x0FE7F0FE7F0FE7F0FE7F0FE7F0FE7F0FE7F0FE7F0FE7F0FE7F0FE7F0FE7F0FE7F0FE7F0FE7F0FE7F" ;
    defparam cpu_rom_0_0_0.INITVAL_16 = "0x0FE7F0FE7F0FE7F0FE7F0FE7F0FE7F0FE7F0FE7F0FE7F0FE7F0FE7F0FE7F0FE7F0FE7F0FE7F0FE7F" ;
    defparam cpu_rom_0_0_0.INITVAL_15 = "0x0FE7F0FE7F0FE7F0FE7F0FE7F0FE7F0FE7F0FE7F0FE7F0FE7F0FE7F0FE7F0FE7F0FE7F0FE7F0FE7F" ;
    defparam cpu_rom_0_0_0.INITVAL_14 = "0x0FE7F0FE7F0FE7F0FE7F0FE7F0FE7F0FE7F0FE7F0FE7F0FE7F0FE7F0FE7F0FE7F0FE7F0FE7F0FE7F" ;
    defparam cpu_rom_0_0_0.INITVAL_13 = "0x0FE7F0FE7F0FE7F0FE7F0FE7F0FE7F0FE7F0FE7F0FE7F0FE7F0FE7F0FE7F0FE7F0FE7F0FE7F0FE7F" ;
    defparam cpu_rom_0_0_0.INITVAL_12 = "0x0FE7F0FE7F0FE7F0FE7F0FE7F0FE7F0FE7F0FE7F0FE7F0FE7F0FE7F0FE7F0FE7F0FE7F0FE7F0FE7F" ;
    defparam cpu_rom_0_0_0.INITVAL_11 = "0x0FE7F0FE7F0FE7F0FE7F0FE7F0FE7F0FE050007F00E07008050060500C0300403002040040300C03" ;
    defparam cpu_rom_0_0_0.INITVAL_10 = "0x002010040300202006010000200A0600602002000040400602002020060200201000010020100201" ;
    defparam cpu_rom_0_0_0.INITVAL_0F = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam cpu_rom_0_0_0.INITVAL_0E = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam cpu_rom_0_0_0.INITVAL_0D = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam cpu_rom_0_0_0.INITVAL_0C = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam cpu_rom_0_0_0.INITVAL_0B = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam cpu_rom_0_0_0.INITVAL_0A = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam cpu_rom_0_0_0.INITVAL_09 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam cpu_rom_0_0_0.INITVAL_08 = "0x00000000000000000000000000000000000000000000000000000000000000000000000000000000" ;
    defparam cpu_rom_0_0_0.INITVAL_07 = "0x3FFFF3FFFF3FFFF3FFFF3FFFF3FFFF3FFFF3FFFF3FFFF3FFFF3FFFF3FFFF3FFFF3FFFF3FFFF3FFFF" ;
    defparam cpu_rom_0_0_0.INITVAL_06 = "0x3FFFF3FFFF3FFFF3FFFF3FFFF3FFFF3FFFF3FFFF3FFFF3FFFF3FFFF3FFFF3FFFF3FFFF3FFFF3FFFF" ;
    defparam cpu_rom_0_0_0.INITVAL_05 = "0x3FFFF3FFFF3FFFF3FFFF3FFFF3FFFF3FFFF3FFFF3FFFF3FFFF3FFFF3FFFF3FFFF3FFFF3FFFF3FFFF" ;
    defparam cpu_rom_0_0_0.INITVAL_04 = "0x3FFFF3FFFF3FFFF3FFFF3FFFF3FFFF3FFFF3FFFF3FFFF3FFFF3FFFF3FFFF3FFFF3FFFF3FFFF3FFFF" ;
    defparam cpu_rom_0_0_0.INITVAL_03 = "0x3FFFF3FFFF3FFFF3FFFF3FFFF3FFFF3FFFF3FFFF3FFFF3FFFF3FFFF3FFFF3FFFF3FFFF3FFFF3FFFF" ;
    defparam cpu_rom_0_0_0.INITVAL_02 = "0x3FFFF3FFFF3FFFF3FFFF3FFFF3FFFF3FFFF3FFFF3FFFF3FFFF3FFFF3FFFF3FFFF3FFFF3FFFF3FFFF" ;
    defparam cpu_rom_0_0_0.INITVAL_01 = "0x3FFFF3FFFF3FFFF3FFFF3FFFF3FFFF3FE0622100206632C13100A242007400212241100242120023" ;
    defparam cpu_rom_0_0_0.INITVAL_00 = "0x07110022122401102520224110321622500241120221022500240112250024071203100FE600BE41" ;
    defparam cpu_rom_0_0_0.CSDECODE_B = "0b000" ;
    defparam cpu_rom_0_0_0.CSDECODE_A = "0b000" ;
    defparam cpu_rom_0_0_0.WRITEMODE_B = "NORMAL" ;
    defparam cpu_rom_0_0_0.WRITEMODE_A = "NORMAL" ;
    defparam cpu_rom_0_0_0.GSR = "ENABLED" ;
    defparam cpu_rom_0_0_0.RESETMODE = "ASYNC" ;
    defparam cpu_rom_0_0_0.REGMODE_B = "OUTREG" ;
    defparam cpu_rom_0_0_0.REGMODE_A = "OUTREG" ;
    defparam cpu_rom_0_0_0.DATA_WIDTH_B = 9 ;
    defparam cpu_rom_0_0_0.DATA_WIDTH_A = 9 ;
    DP8KC cpu_rom_0_0_0 (.DIA8(scuba_vlo), .DIA7(scuba_vlo), .DIA6(scuba_vlo),
        .DIA5(scuba_vlo), .DIA4(scuba_vlo), .DIA3(scuba_vlo), .DIA2(scuba_vlo),
        .DIA1(scuba_vlo), .DIA0(scuba_vlo), .ADA12(scuba_vlo), .ADA11(scuba_vlo),
        .ADA10(Address[7]), .ADA9(Address[6]), .ADA8(Address[5]), .ADA7(Address[4]),
        .ADA6(Address[3]), .ADA5(Address[2]), .ADA4(Address[1]), .ADA3(Address[0]),
        .ADA2(scuba_vlo), .ADA1(scuba_vlo), .ADA0(scuba_vlo), .CEA(OutClockEn),
        .OCEA(OutClockEn), .CLKA(OutClock), .WEA(scuba_vlo), .CSA2(scuba_vlo),
        .CSA1(scuba_vlo), .CSA0(scuba_vlo), .RSTA(Reset), .DIB8(scuba_vlo),
        .DIB7(scuba_vlo), .DIB6(scuba_vlo), .DIB5(scuba_vlo), .DIB4(scuba_vlo),
        .DIB3(scuba_vlo), .DIB2(scuba_vlo), .DIB1(scuba_vlo), .DIB0(scuba_vlo),
        .ADB12(scuba_vhi), .ADB11(scuba_vlo), .ADB10(Address[7]), .ADB9(Address[6]),
        .ADB8(Address[5]), .ADB7(Address[4]), .ADB6(Address[3]), .ADB5(Address[2]),
        .ADB4(Address[1]), .ADB3(Address[0]), .ADB2(scuba_vlo), .ADB1(scuba_vlo),
        .ADB0(scuba_vlo), .CEB(OutClockEn), .OCEB(OutClockEn), .CLKB(OutClock),
        .WEB(scuba_vlo), .CSB2(scuba_vlo), .CSB1(scuba_vlo), .CSB0(scuba_vlo),
        .RSTB(Reset), .DOA8(Q[8]), .DOA7(Q[7]), .DOA6(Q[6]), .DOA5(Q[5]),
        .DOA4(Q[4]), .DOA3(Q[3]), .DOA2(Q[2]), .DOA1(Q[1]), .DOA0(Q[0]),
        .DOB8(), .DOB7(), .DOB6(Q[15]), .DOB5(Q[14]), .DOB4(Q[13]), .DOB3(Q[12]),
        .DOB2(Q[11]), .DOB1(Q[10]), .DOB0(Q[9]))
             /* synthesis MEM_LPC_FILE="cpu_rom.lpc" */
             /* synthesis MEM_INIT_FILE="cic_prog.mem" */;
    // exemplar begin
    // exemplar attribute cpu_rom_0_0_0 MEM_LPC_FILE cpu_rom.lpc
    // exemplar attribute cpu_rom_0_0_0 MEM_INIT_FILE cic_prog.mem
    // exemplar end
endmodule