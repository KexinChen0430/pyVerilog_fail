module
    // if port is stubbed
    ,.ready_i(ready_li)
    ,.my_x_i
    ,.my_y_i
    );
endmodule