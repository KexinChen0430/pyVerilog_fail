module tb;
	localparam [11:0] UPAE1 = 10;
	localparam [11:0] UPAF1 = 10;
	localparam [10:0] UPAE2 = 10;
	localparam [10:0] UPAF2 = 10;
	localparam [0:0] SPLIT = 0;
	localparam [0:0] SYNC_FIFO1 = 0;
	localparam [0:0] SYNC_FIFO2 = 0;
	localparam [0:0] FMODE1 = 1;
	localparam [0:0] POWERDN1 = 0;
	localparam [0:0] SLEEP1 = 0;
	localparam [0:0] PROTECT1 = 0;
	localparam [0:0] FMODE2 = 0;
	localparam [0:0] POWERDN2 = 0;
	localparam [0:0] SLEEP2 = 0;
	localparam [0:0] PROTECT2 = 0;
	localparam [2:0] RMODE_A1 = MODE_36;
	localparam [2:0] RMODE_B1 = MODE_36;
	localparam [2:0] WMODE_A1 = MODE_36;
	localparam [2:0] WMODE_B1 = MODE_36;
	localparam [2:0] RMODE_A2 = MODE_36;
	localparam [2:0] RMODE_B2 = MODE_36;
	localparam [2:0] WMODE_A2 = MODE_36;
	localparam [2:0] WMODE_B2 = MODE_36;
	localparam W_PERIOD = 30;
	localparam R_PERIOD = 29;
	reg WEN_A1;
	reg WEN_B1;
	reg REN_A1;
	reg REN_B1;
	reg CLK_A1;
	reg CLK_B1;
	reg [1:0] BE_A1;
	reg [1:0] BE_B1;
	reg [14:0] ADDR_A1;
	reg [14:0] ADDR_B1;
	reg [17:0] WDATA_A1;
	reg [17:0] WDATA_B1;
	wire [17:0] RDATA_A1;
	wire [17:0] RDATA_B1;
	wire UNDERRUN1;
	wire OVERRUN1;
	wire UNDERRUN2;
	wire OVERRUN2;
	wire EMPTY1;
	wire EPO1;
	wire EWM1;
	wire FULL1;
	wire FMO1;
	wire FWM1;
	reg FLUSH1;
	reg WEN_A2;
	reg WEN_B2;
	reg REN_A2;
	reg REN_B2;
	reg CLK_A2;
	reg CLK_B2;
	reg [1:0] BE_A2;
	reg [1:0] BE_B2;
	wire [13:0] ADDR_A2;
	wire [13:0] ADDR_B2;
	reg [17:0] WDATA_A2;
	reg [17:0] WDATA_B2;
	wire [17:0] RDATA_A2;
	wire [17:0] RDATA_B2;
	wire EMPTY2;
	wire EPO2;
	wire EWM2;
	wire FULL2;
	wire FMO2;
	wire FWM2;
	reg FLUSH2;
	wire [17:0] RDATA_A18;
	wire [17:0] RDATA_B18;
	wire [8:0] RDATA_A9;
	wire [8:0] RDATA_B9;
	wire [35:0] expected_data_a;
	wire [35:0] expected_data_b;
	wire [35:0] last_expected_a;
	wire [35:0] last_expected_b;
	wire [17:0] last_expected_a18;
	wire [17:0] last_expected_b18;
	wire [8:0] last_expected_a9;
	wire [8:0] last_expected_b9;
	wire [14:0] last_addr_a;
	wire [14:0] last_addr_b;
	wire valid_a;
	wire valid_b;
	wire [3:0] index4_a;
	wire [3:0] index4_b;
	wire [1:0] index2_a;
	wire [1:0] index2_b;
	wire index_a;
	wire index_b;
	reg last_empty1;
	wire last_empty2;
	wire [35:0] fifo_dout;
	wire [35:0] fifo_din;
	localparam MODE_36 = 3'b011;
	task fA_36x36;
		begin
			$display("%d: Fifo 36-bit write 36-bit read", $time);
			FLUSH1 = 1;
			@(posedge CLK_A1);
			@(posedge CLK_B1);
			FLUSH1 = 0;
		end
	endtask
	task fA_push36;
		input [35:0] data;
		begin
			@(negedge CLK_A1) begin
				WDATA_A2 = data[35:18];
				WDATA_A1 = data[17:0];
				WEN_A1 = 1;
			end
			@(posedge CLK_A1)
				#(2) WEN_A1 = 0;
		end
	endtask
	task fA_pop;
		input [35:0] expected;
		input [35:0] msk;
		begin
			if (last_empty1 || EMPTY1)
				while (EMPTY1 == 1) begin
					@(posedge CLK_B1);
				end
			if (({RDATA_B2, RDATA_B1} & msk) !== expected) begin
				$display("%d: POP FIFO ERROR: mismatch: expected = %9x mask = %5x, actuall = %9x", $time, expected, msk, {RDATA_B2, RDATA_B1});
				error_cnt = error_cnt + 1'b1;
			end
			@(negedge CLK_B1) REN_B1 = 1;
			@(posedge CLK_B1)
				#(2) REN_B1 = 0;
		end
	endtask
	integer wcount_a;
	integer rcount_a;
	integer state_a;
	integer wcount_b;
	integer rcount_b;
	integer state_b;
	integer error_cnt = 0;
	initial CLK_A1 = 0;
	initial CLK_B1 = 0;
	initial CLK_A2 = 0;
	initial CLK_B2 = 0;
	initial forever #(R_PERIOD) CLK_A1 = ~CLK_A1;
	initial forever #(W_PERIOD) CLK_B1 = ~CLK_B1;
	initial forever #(R_PERIOD) CLK_A2 = ~CLK_A2;
	initial forever #(W_PERIOD) CLK_B2 = ~CLK_B2;
	initial begin
		$dumpfile(`VCD_FILE);
		$dumpvars(0, tb);
	end
	initial #(1) begin
		WEN_A1 = 0;
		REN_A1 = 0;
		WEN_B1 = 0;
		REN_B1 = 0;
		BE_A1 = 2'b11;
		BE_A2 = 2'b11;
		BE_B1 = 2'b11;
		BE_B2 = 2'b11;
		ADDR_A1 = 14'b00000000000000;
		ADDR_B1 = 14'b00000000000000;
		WDATA_A1 = 18'b000000000000000000;
		WDATA_B1 = 18'h00000;
		wcount_a = 0;
		rcount_a = 0;
		state_a = 0;
		wcount_b = 0;
		rcount_b = 0;
		state_b = 0;
		WEN_A2 = 0;
		REN_A2 = 0;
		WEN_B2 = 0;
		REN_B2 = 0;
		FLUSH1 = 0;
		FLUSH2 = 0;
	end
	initial begin
		#(100)
		@(posedge CLK_A1);
		@(posedge CLK_B1);
	end
	assign fifo_dout = {RDATA_B2, RDATA_B1};
	assign fifo_din = {WDATA_A2, WDATA_A1};
	assign {EMPTY1, EPO1, EWM1, UNDERRUN1, FULL1, FMO1, FWM1, OVERRUN1} = RDATA_A1[7:0];
	assign {EMPTY2, EPO2, EWM2, UNDERRUN2, FULL2, FMO2, FWM2, OVERRUN2} = RDATA_A2[7:0];
	always @(posedge CLK_B1) last_empty1 <= EMPTY1;
	always @(*)
		case (state_a)
			0: begin
				fA_36x36;
				if (!EMPTY1) begin
					$display("%d: FIFO ERROR: EMPTY flag not set", $time);
					error_cnt = error_cnt + 1'b1;
				end
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				if (!EMPTY1) begin
					$display("%d: FIFO ERROR: EMPTY flag not set", $time);
					error_cnt = error_cnt + 1'b1;
				end
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				if (!EMPTY1) begin
					$display("%d: FIFO ERROR: EMPTY flag not set", $time);
					error_cnt = error_cnt + 1'b1;
				end
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				fA_push36(36'h0a5a5a5a5);
				fA_push36(36'h05a5a5a5a);
				if (!FULL1) begin
					$display("%d: FIFO ERROR: FULL flag not set", $time);
					error_cnt = error_cnt + 1'b1;
				end
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				fA_pop(36'h0a5a5a5a5, {36 {1'b1}});
				fA_pop(36'h05a5a5a5a, {36 {1'b1}});
				if (!EMPTY1) begin
					$display("%d: FIFO ERROR: EMPTY flag not set", $time);
					error_cnt = error_cnt + 1'b1;
				end
				@(posedge CLK_A1);
				@(posedge CLK_B1);
				@(posedge CLK_A1);
				@(posedge CLK_B1);
				@(posedge CLK_A1);
				@(posedge CLK_B1);
				@(posedge CLK_A1);
				@(posedge CLK_B1);
				@(posedge CLK_A1);
				@(posedge CLK_B1);
				@(posedge CLK_A1);
				@(posedge CLK_B1);
				$finish_and_return( (error_cnt == 0) ? 0 : -1 );
			end
		endcase
	TDP36K #(
		.MODE_BITS({SPLIT, UPAF2, UPAE2, PROTECT2, SLEEP2, POWERDN2, FMODE2, WMODE_B2, WMODE_A2, RMODE_B2, RMODE_A2, SYNC_FIFO2, UPAF1, UPAE1, PROTECT1, SLEEP1, POWERDN1, FMODE1, WMODE_B1, WMODE_A1, RMODE_B1, RMODE_A1, SYNC_FIFO1})
	)tdp36_1(
		.CLK_A1_i(CLK_A1),
		.CLK_B1_i(CLK_B1),
		.WEN_A1_i(WEN_A1),
		.WEN_B1_i(WEN_B1),
		.REN_A1_i(REN_A1),
		.REN_B1_i(REN_B1),
		.BE_A1_i(BE_A1),
		.BE_B1_i(BE_B1),
		.ADDR_A1_i(ADDR_A1),
		.ADDR_B1_i(ADDR_B1),
		.WDATA_A1_i(WDATA_A1),
		.WDATA_B1_i(WDATA_B1),
		.RDATA_A1_o(RDATA_A1),
		.RDATA_B1_o(RDATA_B1),
		.FLUSH1_i(FLUSH1),
		.CLK_A2_i(CLK_A2),
		.CLK_B2_i(CLK_B2),
		.WEN_A2_i(WEN_A2),
		.WEN_B2_i(WEN_B2),
		.REN_A2_i(REN_A2),
		.REN_B2_i(REN_B2),
		.BE_A2_i(BE_A2),
		.BE_B2_i(BE_B2),
		.ADDR_A2_i(ADDR_A2),
		.ADDR_B2_i(ADDR_B2),
		.WDATA_A2_i(WDATA_A2),
		.WDATA_B2_i(WDATA_B2),
		.RDATA_A2_o(RDATA_A2),
		.RDATA_B2_o(RDATA_B2),
		.FLUSH2_i(FLUSH2)
	);
endmodule