module header
	// Internal signals
	// Generated Signal List
	// End of Generated Signal List
	// %COMPILER_OPTS%
	// Generated Signal Assignments
	// Generated Instances and Port Mappings
		// Generated Instance Port Map for ebi_cs2_pad
		WYNA28SGA ebi_cs2_pad (
		);
		// End of Generated Instance Port Map for ebi_cs2_pad
		// Generated Instance Port Map for ebi_cs3_pad
		WYNA28SGA ebi_cs3_pad (
		);
		// End of Generated Instance Port Map for ebi_cs3_pad
		// Generated Instance Port Map for vgch_io_i
		vgch_io vgch_io_i (
		);
		// End of Generated Instance Port Map for vgch_io_i
endmodule