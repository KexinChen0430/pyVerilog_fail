module sky130_fd_sc_ms__udp_pwrgood_pp$G (
    UDP_OUT,
    UDP_IN ,
    VGND
);
    output UDP_OUT;
    input  UDP_IN ;
    input  VGND   ;
endmodule