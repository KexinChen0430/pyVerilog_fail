module shiftleft2_Testbench;
reg [31:0] inputA;
wire [31:0] result;
shiftleft2 UUT(inputA,result);
   initial begin
       #20 inputA = 32'b0000_0000_0000_0000_1010_1010_1010_1010;
       #40 inputA = 32'b0000_0000_0000_0000_1111_1111_1111_1111;
       #40 inputA = 32'b1110_1110_1110_1110_1110_1110_1110_1110;
       #40 inputA = 32'b1001_1001_1001_1001_0110_0110_0110_0110;
       #40 inputA = 32'b0000_1000_0001_0000_0100_0010_0010_0101;
       #40 inputA = 32'b0000_1111_0000_1111_0000_1111_0000_1111;
       #40 inputA = 32'b1111_0000_1111_0000_1111_0000_1111_0000;
       #40 inputA = 32'b0110_0011_1100_0110_0011_1100_0110_0011;
   end
   initial
       #340 $stop;
endmodule