module top ;
          wire  Net_14;
          wire  Net_12;
          wire  Net_24;
          wire  Net_10;
          wire  Net_23;
          wire  Net_22;
          wire  Net_21;
          wire  Net_20;
          wire  Net_19;
          wire  Net_18;
          wire  Net_17;
          wire  Net_16;
          wire  Net_15;
    TCPWM_P4_v1_10_0 PWM_1 (
        .stop(1'b0),
        .reload(1'b0),
        .start(1'b0),
        .count(1'b1),
        .capture(1'b0),
        .interrupt(Net_20),
        .ov(Net_21),
        .un(Net_22),
        .cc(Net_23),
        .line(Net_10),
        .line_n(Net_24),
        .clock(Net_12));
    defparam PWM_1.PWMCountMode = 3;
    defparam PWM_1.PWMReloadMode = 0;
    defparam PWM_1.PWMReloadPresent = 0;
    defparam PWM_1.PWMStartMode = 0;
    defparam PWM_1.PWMStopMode = 0;
    defparam PWM_1.PWMSwitchMode = 0;
    defparam PWM_1.QuadIndexMode = 0;
    defparam PWM_1.QuadPhiAMode = 3;
    defparam PWM_1.QuadPhiBMode = 3;
    defparam PWM_1.QuadStopMode = 0;
    defparam PWM_1.TCCaptureMode = 0;
    defparam PWM_1.TCCountMode = 3;
    defparam PWM_1.TCReloadMode = 0;
    defparam PWM_1.TCStartMode = 0;
    defparam PWM_1.TCStopMode = 0;
	cy_clock_v1_0
		#(.id("98c2df8a-317f-46c0-877f-ddd17972fb4c"),
		  .source_clock_id(""),
		  .divisor(0),
		  .period("1000000000"),
		  .is_direct(0),
		  .is_digital(0))
		servoClock
		 (.clock_out(Net_12));
	wire [0:0] tmpOE__Servo_net;
	wire [0:0] tmpFB_0__Servo_net;
	wire [0:0] tmpIO_0__Servo_net;
	wire [0:0] tmpINTERRUPT_0__Servo_net;
	electrical [0:0] tmpSIOVREF__Servo_net;
	cy_psoc3_pins_v1_10
		#(.id("0e0c9380-6965-4440-8709-ce08a91e474c"),
		  .drive_mode(3'b110),
		  .ibuf_enabled(1'b1),
		  .init_dr_st(1'b1),
		  .input_clk_en(0),
		  .input_sync(1'b1),
		  .input_sync_mode(1'b0),
		  .intr_mode(2'b00),
		  .invert_in_clock(0),
		  .invert_in_clock_en(0),
		  .invert_in_reset(0),
		  .invert_out_clock(0),
		  .invert_out_clock_en(0),
		  .invert_out_reset(0),
		  .io_voltage(""),
		  .layout_mode("CONTIGUOUS"),
		  .oe_conn(1'b0),
		  .oe_reset(0),
		  .oe_sync(1'b0),
		  .output_clk_en(0),
		  .output_clock_mode(1'b0),
		  .output_conn(1'b1),
		  .output_mode(1'b0),
		  .output_reset(0),
		  .output_sync(1'b0),
		  .pa_in_clock(-1),
		  .pa_in_clock_en(-1),
		  .pa_in_reset(-1),
		  .pa_out_clock(-1),
		  .pa_out_clock_en(-1),
		  .pa_out_reset(-1),
		  .pin_aliases(""),
		  .pin_mode("O"),
		  .por_state(4),
		  .sio_group_cnt(0),
		  .sio_hyst(1'b0),
		  .sio_ibuf(""),
		  .sio_info(2'b00),
		  .sio_obuf(""),
		  .sio_refsel(""),
		  .sio_vtrip(""),
		  .slew_rate(1'b0),
		  .spanning(0),
		  .use_annotation(1'b0),
		  .vtrip(2'b10),
		  .width(1))
		Servo
		 (.oe(tmpOE__Servo_net),
		  .y({Net_10}),
		  .fb({tmpFB_0__Servo_net[0:0]}),
		  .io({tmpIO_0__Servo_net[0:0]}),
		  .siovref(tmpSIOVREF__Servo_net),
		  .interrupt({tmpINTERRUPT_0__Servo_net[0:0]}),
		  .in_clock({1'b0}),
		  .in_clock_en({1'b1}),
		  .in_reset({1'b0}),
		  .out_clock({1'b0}),
		  .out_clock_en({1'b1}),
		  .out_reset({1'b0}));
	assign tmpOE__Servo_net = (`CYDEV_CHIP_MEMBER_USED == `CYDEV_CHIP_MEMBER_3A && `CYDEV_CHIP_REVISION_USED < `CYDEV_CHIP_REVISION_3A_ES3) ? ~{1'b1} : {1'b1};
endmodule