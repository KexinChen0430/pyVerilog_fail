module cell_with_typeparam;
   addr #(.PARAMTYPE(integer)) acell ();
endmodule